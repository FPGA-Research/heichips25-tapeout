magic
tech ihp-sg13g2
magscale 1 2
timestamp 1752757781
<< metal1 >>
rect 1152 41600 20452 41624
rect 1152 41560 4928 41600
rect 4968 41560 5010 41600
rect 5050 41560 5092 41600
rect 5132 41560 5174 41600
rect 5214 41560 5256 41600
rect 5296 41560 20048 41600
rect 20088 41560 20130 41600
rect 20170 41560 20212 41600
rect 20252 41560 20294 41600
rect 20334 41560 20376 41600
rect 20416 41560 20452 41600
rect 1152 41536 20452 41560
rect 2091 41432 2133 41441
rect 2091 41392 2092 41432
rect 2132 41392 2133 41432
rect 2091 41383 2133 41392
rect 5739 41432 5781 41441
rect 5739 41392 5740 41432
rect 5780 41392 5781 41432
rect 5739 41383 5781 41392
rect 6123 41432 6165 41441
rect 6123 41392 6124 41432
rect 6164 41392 6165 41432
rect 6123 41383 6165 41392
rect 9963 41432 10005 41441
rect 9963 41392 9964 41432
rect 10004 41392 10005 41432
rect 9963 41383 10005 41392
rect 10347 41432 10389 41441
rect 10347 41392 10348 41432
rect 10388 41392 10389 41432
rect 10347 41383 10389 41392
rect 13803 41432 13845 41441
rect 13803 41392 13804 41432
rect 13844 41392 13845 41432
rect 13803 41383 13845 41392
rect 15723 41432 15765 41441
rect 15723 41392 15724 41432
rect 15764 41392 15765 41432
rect 15723 41383 15765 41392
rect 16107 41432 16149 41441
rect 16107 41392 16108 41432
rect 16148 41392 16149 41432
rect 16107 41383 16149 41392
rect 17259 41432 17301 41441
rect 17259 41392 17260 41432
rect 17300 41392 17301 41432
rect 17259 41383 17301 41392
rect 17835 41432 17877 41441
rect 17835 41392 17836 41432
rect 17876 41392 17877 41432
rect 17835 41383 17877 41392
rect 18123 41432 18165 41441
rect 18123 41392 18124 41432
rect 18164 41392 18165 41432
rect 18123 41383 18165 41392
rect 18699 41432 18741 41441
rect 18699 41392 18700 41432
rect 18740 41392 18741 41432
rect 18699 41383 18741 41392
rect 19755 41432 19797 41441
rect 19755 41392 19756 41432
rect 19796 41392 19797 41432
rect 19755 41383 19797 41392
rect 2275 41264 2333 41265
rect 2275 41224 2284 41264
rect 2324 41224 2333 41264
rect 2275 41223 2333 41224
rect 3523 41264 3581 41265
rect 3523 41224 3532 41264
rect 3572 41224 3581 41264
rect 3523 41223 3581 41224
rect 4099 41264 4157 41265
rect 4099 41224 4108 41264
rect 4148 41224 4157 41264
rect 4099 41223 4157 41224
rect 5347 41264 5405 41265
rect 5347 41224 5356 41264
rect 5396 41224 5405 41264
rect 5347 41223 5405 41224
rect 6499 41264 6557 41265
rect 6499 41224 6508 41264
rect 6548 41224 6557 41264
rect 6499 41223 6557 41224
rect 7747 41264 7805 41265
rect 7747 41224 7756 41264
rect 7796 41224 7805 41264
rect 7747 41223 7805 41224
rect 8131 41264 8189 41265
rect 8131 41224 8140 41264
rect 8180 41224 8189 41264
rect 8131 41223 8189 41224
rect 9379 41264 9437 41265
rect 9379 41224 9388 41264
rect 9428 41224 9437 41264
rect 9379 41223 9437 41224
rect 11971 41264 12029 41265
rect 11971 41224 11980 41264
rect 12020 41224 12029 41264
rect 11971 41223 12029 41224
rect 13219 41264 13277 41265
rect 13219 41224 13228 41264
rect 13268 41224 13277 41264
rect 13219 41223 13277 41224
rect 1707 41180 1749 41189
rect 1707 41140 1708 41180
rect 1748 41140 1749 41180
rect 1707 41131 1749 41140
rect 1891 41180 1949 41181
rect 1891 41140 1900 41180
rect 1940 41140 1949 41180
rect 1891 41139 1949 41140
rect 5539 41180 5597 41181
rect 5539 41140 5548 41180
rect 5588 41140 5597 41180
rect 5539 41139 5597 41140
rect 5923 41180 5981 41181
rect 5923 41140 5932 41180
rect 5972 41140 5981 41180
rect 5923 41139 5981 41140
rect 9763 41180 9821 41181
rect 9763 41140 9772 41180
rect 9812 41140 9821 41180
rect 9763 41139 9821 41140
rect 10147 41180 10205 41181
rect 10147 41140 10156 41180
rect 10196 41140 10205 41180
rect 10147 41139 10205 41140
rect 10531 41180 10589 41181
rect 10531 41140 10540 41180
rect 10580 41140 10589 41180
rect 10531 41139 10589 41140
rect 11587 41180 11645 41181
rect 11587 41140 11596 41180
rect 11636 41140 11645 41180
rect 11587 41139 11645 41140
rect 13987 41180 14045 41181
rect 13987 41140 13996 41180
rect 14036 41140 14045 41180
rect 13987 41139 14045 41140
rect 14563 41180 14621 41181
rect 14563 41140 14572 41180
rect 14612 41140 14621 41180
rect 14563 41139 14621 41140
rect 14947 41180 15005 41181
rect 14947 41140 14956 41180
rect 14996 41140 15005 41180
rect 14947 41139 15005 41140
rect 15331 41180 15389 41181
rect 15331 41140 15340 41180
rect 15380 41140 15389 41180
rect 15331 41139 15389 41140
rect 15907 41180 15965 41181
rect 15907 41140 15916 41180
rect 15956 41140 15965 41180
rect 15907 41139 15965 41140
rect 16291 41180 16349 41181
rect 16291 41140 16300 41180
rect 16340 41140 16349 41180
rect 16291 41139 16349 41140
rect 16587 41180 16629 41189
rect 16587 41140 16588 41180
rect 16628 41140 16629 41180
rect 16587 41131 16629 41140
rect 16963 41180 17021 41181
rect 16963 41140 16972 41180
rect 17012 41140 17021 41180
rect 16963 41139 17021 41140
rect 17443 41180 17501 41181
rect 17443 41140 17452 41180
rect 17492 41140 17501 41180
rect 17443 41139 17501 41140
rect 17635 41180 17693 41181
rect 17635 41140 17644 41180
rect 17684 41140 17693 41180
rect 17635 41139 17693 41140
rect 18307 41180 18365 41181
rect 18307 41140 18316 41180
rect 18356 41140 18365 41180
rect 18307 41139 18365 41140
rect 18499 41180 18557 41181
rect 18499 41140 18508 41180
rect 18548 41140 18557 41180
rect 18499 41139 18557 41140
rect 19075 41180 19133 41181
rect 19075 41140 19084 41180
rect 19124 41140 19133 41180
rect 19075 41139 19133 41140
rect 19363 41180 19421 41181
rect 19363 41140 19372 41180
rect 19412 41140 19421 41180
rect 19363 41139 19421 41140
rect 19939 41180 19997 41181
rect 19939 41140 19948 41180
rect 19988 41140 19997 41180
rect 19939 41139 19997 41140
rect 1323 41096 1365 41105
rect 1323 41056 1324 41096
rect 1364 41056 1365 41096
rect 1323 41047 1365 41056
rect 3723 41096 3765 41105
rect 3723 41056 3724 41096
rect 3764 41056 3765 41096
rect 3723 41047 3765 41056
rect 9579 41096 9621 41105
rect 9579 41056 9580 41096
rect 9620 41056 9621 41096
rect 9579 41047 9621 41056
rect 11787 41096 11829 41105
rect 11787 41056 11788 41096
rect 11828 41056 11829 41096
rect 11787 41047 11829 41056
rect 16779 41096 16821 41105
rect 16779 41056 16780 41096
rect 16820 41056 16821 41096
rect 16779 41047 16821 41056
rect 18891 41096 18933 41105
rect 18891 41056 18892 41096
rect 18932 41056 18933 41096
rect 18891 41047 18933 41056
rect 3915 41012 3957 41021
rect 3915 40972 3916 41012
rect 3956 40972 3957 41012
rect 3915 40963 3957 40972
rect 6315 41012 6357 41021
rect 6315 40972 6316 41012
rect 6356 40972 6357 41012
rect 6315 40963 6357 40972
rect 7947 41012 7989 41021
rect 7947 40972 7948 41012
rect 7988 40972 7989 41012
rect 7947 40963 7989 40972
rect 13419 41012 13461 41021
rect 13419 40972 13420 41012
rect 13460 40972 13461 41012
rect 13419 40963 13461 40972
rect 14379 41012 14421 41021
rect 14379 40972 14380 41012
rect 14420 40972 14421 41012
rect 14379 40963 14421 40972
rect 14763 41012 14805 41021
rect 14763 40972 14764 41012
rect 14804 40972 14805 41012
rect 14763 40963 14805 40972
rect 15147 41012 15189 41021
rect 15147 40972 15148 41012
rect 15188 40972 15189 41012
rect 15147 40963 15189 40972
rect 19563 41012 19605 41021
rect 19563 40972 19564 41012
rect 19604 40972 19605 41012
rect 19563 40963 19605 40972
rect 1152 40844 20352 40868
rect 1152 40804 3688 40844
rect 3728 40804 3770 40844
rect 3810 40804 3852 40844
rect 3892 40804 3934 40844
rect 3974 40804 4016 40844
rect 4056 40804 18808 40844
rect 18848 40804 18890 40844
rect 18930 40804 18972 40844
rect 19012 40804 19054 40844
rect 19094 40804 19136 40844
rect 19176 40804 20352 40844
rect 1152 40780 20352 40804
rect 1707 40676 1749 40685
rect 1707 40636 1708 40676
rect 1748 40636 1749 40676
rect 1707 40627 1749 40636
rect 3051 40676 3093 40685
rect 3051 40636 3052 40676
rect 3092 40636 3093 40676
rect 3051 40627 3093 40636
rect 3435 40676 3477 40685
rect 3435 40636 3436 40676
rect 3476 40636 3477 40676
rect 3435 40627 3477 40636
rect 5451 40676 5493 40685
rect 5451 40636 5452 40676
rect 5492 40636 5493 40676
rect 5451 40627 5493 40636
rect 5835 40676 5877 40685
rect 5835 40636 5836 40676
rect 5876 40636 5877 40676
rect 5835 40627 5877 40636
rect 7947 40676 7989 40685
rect 7947 40636 7948 40676
rect 7988 40636 7989 40676
rect 7947 40627 7989 40636
rect 16203 40676 16245 40685
rect 16203 40636 16204 40676
rect 16244 40636 16245 40676
rect 16203 40627 16245 40636
rect 16587 40676 16629 40685
rect 16587 40636 16588 40676
rect 16628 40636 16629 40676
rect 16587 40627 16629 40636
rect 16971 40676 17013 40685
rect 16971 40636 16972 40676
rect 17012 40636 17013 40676
rect 16971 40627 17013 40636
rect 18123 40676 18165 40685
rect 18123 40636 18124 40676
rect 18164 40636 18165 40676
rect 18123 40627 18165 40636
rect 18507 40676 18549 40685
rect 18507 40636 18508 40676
rect 18548 40636 18549 40676
rect 18507 40627 18549 40636
rect 18891 40676 18933 40685
rect 18891 40636 18892 40676
rect 18932 40636 18933 40676
rect 18891 40627 18933 40636
rect 11971 40592 12029 40593
rect 11971 40552 11980 40592
rect 12020 40552 12029 40592
rect 11971 40551 12029 40552
rect 15819 40592 15861 40601
rect 15819 40552 15820 40592
rect 15860 40552 15861 40592
rect 15819 40543 15861 40552
rect 17931 40592 17973 40601
rect 17931 40552 17932 40592
rect 17972 40552 17973 40592
rect 17931 40543 17973 40552
rect 19563 40592 19605 40601
rect 19563 40552 19564 40592
rect 19604 40552 19605 40592
rect 19563 40543 19605 40552
rect 2851 40519 2909 40520
rect 1507 40508 1565 40509
rect 1507 40468 1516 40508
rect 1556 40468 1565 40508
rect 1507 40467 1565 40468
rect 2283 40508 2325 40517
rect 2283 40468 2284 40508
rect 2324 40468 2325 40508
rect 2851 40479 2860 40519
rect 2900 40479 2909 40519
rect 2851 40478 2909 40479
rect 3235 40508 3293 40509
rect 2283 40459 2325 40468
rect 3235 40468 3244 40508
rect 3284 40468 3293 40508
rect 3235 40467 3293 40468
rect 5251 40508 5309 40509
rect 5251 40468 5260 40508
rect 5300 40468 5309 40508
rect 5251 40467 5309 40468
rect 5635 40508 5693 40509
rect 5635 40468 5644 40508
rect 5684 40468 5693 40508
rect 5635 40467 5693 40468
rect 8131 40508 8189 40509
rect 8131 40468 8140 40508
rect 8180 40468 8189 40508
rect 8131 40467 8189 40468
rect 9003 40508 9045 40517
rect 9003 40468 9004 40508
rect 9044 40468 9045 40508
rect 9003 40459 9045 40468
rect 16003 40508 16061 40509
rect 16003 40468 16012 40508
rect 16052 40468 16061 40508
rect 16003 40467 16061 40468
rect 16387 40508 16445 40509
rect 16387 40468 16396 40508
rect 16436 40468 16445 40508
rect 16387 40467 16445 40468
rect 16771 40508 16829 40509
rect 16771 40468 16780 40508
rect 16820 40468 16829 40508
rect 16771 40467 16829 40468
rect 17155 40508 17213 40509
rect 17155 40468 17164 40508
rect 17204 40468 17213 40508
rect 17155 40467 17213 40468
rect 17731 40508 17789 40509
rect 17731 40468 17740 40508
rect 17780 40468 17789 40508
rect 17731 40467 17789 40468
rect 18307 40508 18365 40509
rect 18307 40468 18316 40508
rect 18356 40468 18365 40508
rect 18307 40467 18365 40468
rect 18691 40508 18749 40509
rect 18691 40468 18700 40508
rect 18740 40468 18749 40508
rect 18691 40467 18749 40468
rect 19075 40508 19133 40509
rect 19075 40468 19084 40508
rect 19124 40468 19133 40508
rect 19075 40467 19133 40468
rect 19363 40508 19421 40509
rect 19363 40468 19372 40508
rect 19412 40468 19421 40508
rect 19363 40467 19421 40468
rect 19843 40508 19901 40509
rect 19843 40468 19852 40508
rect 19892 40468 19901 40508
rect 19843 40467 19901 40468
rect 11587 40445 11645 40446
rect 3811 40424 3869 40425
rect 3811 40384 3820 40424
rect 3860 40384 3869 40424
rect 3811 40383 3869 40384
rect 5059 40424 5117 40425
rect 5059 40384 5068 40424
rect 5108 40384 5117 40424
rect 5059 40383 5117 40384
rect 6019 40424 6077 40425
rect 6019 40384 6028 40424
rect 6068 40384 6077 40424
rect 6019 40383 6077 40384
rect 7267 40424 7325 40425
rect 7267 40384 7276 40424
rect 7316 40384 7325 40424
rect 7267 40383 7325 40384
rect 8427 40424 8469 40433
rect 8427 40384 8428 40424
rect 8468 40384 8469 40424
rect 8427 40375 8469 40384
rect 8523 40424 8565 40433
rect 8523 40384 8524 40424
rect 8564 40384 8565 40424
rect 8523 40375 8565 40384
rect 8907 40424 8949 40433
rect 9963 40429 10005 40438
rect 8907 40384 8908 40424
rect 8948 40384 8949 40424
rect 8907 40375 8949 40384
rect 9475 40424 9533 40425
rect 9475 40384 9484 40424
rect 9524 40384 9533 40424
rect 9475 40383 9533 40384
rect 9963 40389 9964 40429
rect 10004 40389 10005 40429
rect 9963 40380 10005 40389
rect 10339 40424 10397 40425
rect 10339 40384 10348 40424
rect 10388 40384 10397 40424
rect 11587 40405 11596 40445
rect 11636 40405 11645 40445
rect 11587 40404 11645 40405
rect 11979 40424 12021 40433
rect 10339 40383 10397 40384
rect 11979 40384 11980 40424
rect 12020 40384 12021 40424
rect 11979 40375 12021 40384
rect 12075 40424 12117 40433
rect 12075 40384 12076 40424
rect 12116 40384 12117 40424
rect 12075 40375 12117 40384
rect 12267 40424 12309 40433
rect 12267 40384 12268 40424
rect 12308 40384 12309 40424
rect 12267 40375 12309 40384
rect 12547 40424 12605 40425
rect 12547 40384 12556 40424
rect 12596 40384 12605 40424
rect 12547 40383 12605 40384
rect 13795 40424 13853 40425
rect 13795 40384 13804 40424
rect 13844 40384 13853 40424
rect 13795 40383 13853 40384
rect 14371 40424 14429 40425
rect 14371 40384 14380 40424
rect 14420 40384 14429 40424
rect 14371 40383 14429 40384
rect 15619 40424 15677 40425
rect 15619 40384 15628 40424
rect 15668 40384 15677 40424
rect 15619 40383 15677 40384
rect 1899 40340 1941 40349
rect 1899 40300 1900 40340
rect 1940 40300 1941 40340
rect 1899 40291 1941 40300
rect 7467 40340 7509 40349
rect 7467 40300 7468 40340
rect 7508 40300 7509 40340
rect 7467 40291 7509 40300
rect 7659 40340 7701 40349
rect 7659 40300 7660 40340
rect 7700 40300 7701 40340
rect 7659 40291 7701 40300
rect 11787 40340 11829 40349
rect 11787 40300 11788 40340
rect 11828 40300 11829 40340
rect 11787 40291 11829 40300
rect 17547 40340 17589 40349
rect 17547 40300 17548 40340
rect 17588 40300 17589 40340
rect 17547 40291 17589 40300
rect 1227 40256 1269 40265
rect 1227 40216 1228 40256
rect 1268 40216 1269 40256
rect 1227 40207 1269 40216
rect 3627 40256 3669 40265
rect 3627 40216 3628 40256
rect 3668 40216 3669 40256
rect 3627 40207 3669 40216
rect 10155 40256 10197 40265
rect 10155 40216 10156 40256
rect 10196 40216 10197 40256
rect 10155 40207 10197 40216
rect 13995 40256 14037 40265
rect 13995 40216 13996 40256
rect 14036 40216 14037 40256
rect 13995 40207 14037 40216
rect 14187 40256 14229 40265
rect 14187 40216 14188 40256
rect 14228 40216 14229 40256
rect 14187 40207 14229 40216
rect 20043 40256 20085 40265
rect 20043 40216 20044 40256
rect 20084 40216 20085 40256
rect 20043 40207 20085 40216
rect 1152 40088 20452 40112
rect 1152 40048 4928 40088
rect 4968 40048 5010 40088
rect 5050 40048 5092 40088
rect 5132 40048 5174 40088
rect 5214 40048 5256 40088
rect 5296 40048 20048 40088
rect 20088 40048 20130 40088
rect 20170 40048 20212 40088
rect 20252 40048 20294 40088
rect 20334 40048 20376 40088
rect 20416 40048 20452 40088
rect 1152 40024 20452 40048
rect 1707 39920 1749 39929
rect 1707 39880 1708 39920
rect 1748 39880 1749 39920
rect 1707 39871 1749 39880
rect 8227 39920 8285 39921
rect 8227 39880 8236 39920
rect 8276 39880 8285 39920
rect 8227 39879 8285 39880
rect 9963 39920 10005 39929
rect 9963 39880 9964 39920
rect 10004 39880 10005 39920
rect 9963 39871 10005 39880
rect 12067 39920 12125 39921
rect 12067 39880 12076 39920
rect 12116 39880 12125 39920
rect 12067 39879 12125 39880
rect 12931 39920 12989 39921
rect 12931 39880 12940 39920
rect 12980 39880 12989 39920
rect 12931 39879 12989 39880
rect 18315 39920 18357 39929
rect 18315 39880 18316 39920
rect 18356 39880 18357 39920
rect 18315 39871 18357 39880
rect 18507 39920 18549 39929
rect 18507 39880 18508 39920
rect 18548 39880 18549 39920
rect 18507 39871 18549 39880
rect 18891 39920 18933 39929
rect 18891 39880 18892 39920
rect 18932 39880 18933 39920
rect 18891 39871 18933 39880
rect 3723 39836 3765 39845
rect 3723 39796 3724 39836
rect 3764 39796 3765 39836
rect 3723 39787 3765 39796
rect 8043 39836 8085 39845
rect 8043 39796 8044 39836
rect 8084 39796 8085 39836
rect 8043 39787 8085 39796
rect 11691 39836 11733 39845
rect 11691 39796 11692 39836
rect 11732 39796 11733 39836
rect 11691 39787 11733 39796
rect 15051 39836 15093 39845
rect 15051 39796 15052 39836
rect 15092 39796 15093 39836
rect 15051 39787 15093 39796
rect 1995 39752 2037 39761
rect 1995 39712 1996 39752
rect 2036 39712 2037 39752
rect 3043 39752 3101 39753
rect 1995 39703 2037 39712
rect 2091 39733 2133 39742
rect 2091 39693 2092 39733
rect 2132 39693 2133 39733
rect 3043 39712 3052 39752
rect 3092 39712 3101 39752
rect 4003 39752 4061 39753
rect 3043 39711 3101 39712
rect 3579 39742 3621 39751
rect 3579 39702 3580 39742
rect 3620 39702 3621 39742
rect 4003 39712 4012 39752
rect 4052 39712 4061 39752
rect 4003 39711 4061 39712
rect 5251 39752 5309 39753
rect 5251 39712 5260 39752
rect 5300 39712 5309 39752
rect 5251 39711 5309 39712
rect 6315 39752 6357 39761
rect 6315 39712 6316 39752
rect 6356 39712 6357 39752
rect 6315 39703 6357 39712
rect 6411 39752 6453 39761
rect 6411 39712 6412 39752
rect 6452 39712 6453 39752
rect 6411 39703 6453 39712
rect 7363 39752 7421 39753
rect 7363 39712 7372 39752
rect 7412 39712 7421 39752
rect 7363 39711 7421 39712
rect 7851 39747 7893 39756
rect 7851 39707 7852 39747
rect 7892 39707 7893 39747
rect 8515 39752 8573 39753
rect 8515 39712 8524 39752
rect 8564 39712 8573 39752
rect 8515 39711 8573 39712
rect 9763 39752 9821 39753
rect 9763 39712 9772 39752
rect 9812 39712 9821 39752
rect 9763 39711 9821 39712
rect 10243 39752 10301 39753
rect 10243 39712 10252 39752
rect 10292 39712 10301 39752
rect 10243 39711 10301 39712
rect 11491 39752 11549 39753
rect 11491 39712 11500 39752
rect 11540 39712 11549 39752
rect 11491 39711 11549 39712
rect 11875 39752 11933 39753
rect 11875 39712 11884 39752
rect 11924 39712 11933 39752
rect 11875 39711 11933 39712
rect 11971 39752 12029 39753
rect 11971 39712 11980 39752
rect 12020 39712 12029 39752
rect 11971 39711 12029 39712
rect 12171 39752 12213 39761
rect 12171 39712 12172 39752
rect 12212 39712 12213 39752
rect 3579 39693 3621 39702
rect 7851 39698 7893 39707
rect 12171 39703 12213 39712
rect 12267 39752 12309 39761
rect 12267 39712 12268 39752
rect 12308 39712 12309 39752
rect 12267 39703 12309 39712
rect 12360 39752 12418 39753
rect 12360 39712 12369 39752
rect 12409 39712 12418 39752
rect 12360 39711 12418 39712
rect 12651 39752 12693 39761
rect 12651 39712 12652 39752
rect 12692 39712 12693 39752
rect 12651 39703 12693 39712
rect 12747 39752 12789 39761
rect 12747 39712 12748 39752
rect 12788 39712 12789 39752
rect 12747 39703 12789 39712
rect 13323 39752 13365 39761
rect 13323 39712 13324 39752
rect 13364 39712 13365 39752
rect 13323 39703 13365 39712
rect 13419 39752 13461 39761
rect 13419 39712 13420 39752
rect 13460 39712 13461 39752
rect 13419 39703 13461 39712
rect 14371 39752 14429 39753
rect 14371 39712 14380 39752
rect 14420 39712 14429 39752
rect 14371 39711 14429 39712
rect 14859 39747 14901 39756
rect 14859 39707 14860 39747
rect 14900 39707 14901 39747
rect 15427 39752 15485 39753
rect 15427 39712 15436 39752
rect 15476 39712 15485 39752
rect 15427 39711 15485 39712
rect 16675 39752 16733 39753
rect 16675 39712 16684 39752
rect 16724 39712 16733 39752
rect 16675 39711 16733 39712
rect 16971 39752 17013 39761
rect 16971 39712 16972 39752
rect 17012 39712 17013 39752
rect 14859 39698 14901 39707
rect 16971 39703 17013 39712
rect 17163 39752 17205 39761
rect 17163 39712 17164 39752
rect 17204 39712 17205 39752
rect 17163 39703 17205 39712
rect 17251 39752 17309 39753
rect 17251 39712 17260 39752
rect 17300 39712 17309 39752
rect 17251 39711 17309 39712
rect 17547 39752 17589 39761
rect 17547 39712 17548 39752
rect 17588 39712 17589 39752
rect 17547 39703 17589 39712
rect 17643 39752 17685 39761
rect 17643 39712 17644 39752
rect 17684 39712 17685 39752
rect 17643 39703 17685 39712
rect 17739 39752 17781 39761
rect 17739 39712 17740 39752
rect 17780 39712 17781 39752
rect 17739 39703 17781 39712
rect 2091 39684 2133 39693
rect 1507 39668 1565 39669
rect 1507 39628 1516 39668
rect 1556 39628 1565 39668
rect 1507 39627 1565 39628
rect 2475 39668 2517 39677
rect 2475 39628 2476 39668
rect 2516 39628 2517 39668
rect 2475 39619 2517 39628
rect 2571 39668 2613 39677
rect 2571 39628 2572 39668
rect 2612 39628 2613 39668
rect 2571 39619 2613 39628
rect 5931 39668 5973 39677
rect 5931 39628 5932 39668
rect 5972 39628 5973 39668
rect 5931 39619 5973 39628
rect 6795 39668 6837 39677
rect 6795 39628 6796 39668
rect 6836 39628 6837 39668
rect 6795 39619 6837 39628
rect 6891 39668 6933 39677
rect 6891 39628 6892 39668
rect 6932 39628 6933 39668
rect 6891 39619 6933 39628
rect 13803 39668 13845 39677
rect 13803 39628 13804 39668
rect 13844 39628 13845 39668
rect 13803 39619 13845 39628
rect 13899 39668 13941 39677
rect 13899 39628 13900 39668
rect 13940 39628 13941 39668
rect 13899 39619 13941 39628
rect 18691 39668 18749 39669
rect 18691 39628 18700 39668
rect 18740 39628 18749 39668
rect 18691 39627 18749 39628
rect 19075 39668 19133 39669
rect 19075 39628 19084 39668
rect 19124 39628 19133 39668
rect 19075 39627 19133 39628
rect 19459 39668 19517 39669
rect 19459 39628 19468 39668
rect 19508 39628 19517 39668
rect 19459 39627 19517 39628
rect 20035 39668 20093 39669
rect 20035 39628 20044 39668
rect 20084 39628 20093 39668
rect 20035 39627 20093 39628
rect 1323 39584 1365 39593
rect 1323 39544 1324 39584
rect 1364 39544 1365 39584
rect 1323 39535 1365 39544
rect 5643 39584 5685 39593
rect 5643 39544 5644 39584
rect 5684 39544 5685 39584
rect 5643 39535 5685 39544
rect 18219 39584 18261 39593
rect 18219 39544 18220 39584
rect 18260 39544 18261 39584
rect 18219 39535 18261 39544
rect 5451 39500 5493 39509
rect 5451 39460 5452 39500
rect 5492 39460 5493 39500
rect 5451 39451 5493 39460
rect 15243 39500 15285 39509
rect 15243 39460 15244 39500
rect 15284 39460 15285 39500
rect 15243 39451 15285 39460
rect 16971 39500 17013 39509
rect 16971 39460 16972 39500
rect 17012 39460 17013 39500
rect 16971 39451 17013 39460
rect 17923 39500 17981 39501
rect 17923 39460 17932 39500
rect 17972 39460 17981 39500
rect 17923 39459 17981 39460
rect 19659 39500 19701 39509
rect 19659 39460 19660 39500
rect 19700 39460 19701 39500
rect 19659 39451 19701 39460
rect 20235 39500 20277 39509
rect 20235 39460 20236 39500
rect 20276 39460 20277 39500
rect 20235 39451 20277 39460
rect 1152 39332 20352 39356
rect 1152 39292 3688 39332
rect 3728 39292 3770 39332
rect 3810 39292 3852 39332
rect 3892 39292 3934 39332
rect 3974 39292 4016 39332
rect 4056 39292 18808 39332
rect 18848 39292 18890 39332
rect 18930 39292 18972 39332
rect 19012 39292 19054 39332
rect 19094 39292 19136 39332
rect 19176 39292 20352 39332
rect 1152 39268 20352 39292
rect 12459 39164 12501 39173
rect 12459 39124 12460 39164
rect 12500 39124 12501 39164
rect 12459 39115 12501 39124
rect 1515 39080 1557 39089
rect 1515 39040 1516 39080
rect 1556 39040 1557 39080
rect 1515 39031 1557 39040
rect 5355 39080 5397 39089
rect 5355 39040 5356 39080
rect 5396 39040 5397 39080
rect 5355 39031 5397 39040
rect 5835 39080 5877 39089
rect 5835 39040 5836 39080
rect 5876 39040 5877 39080
rect 5835 39031 5877 39040
rect 6219 39080 6261 39089
rect 6219 39040 6220 39080
rect 6260 39040 6261 39080
rect 6219 39031 6261 39040
rect 6603 39080 6645 39089
rect 6603 39040 6604 39080
rect 6644 39040 6645 39080
rect 6603 39031 6645 39040
rect 6795 39080 6837 39089
rect 6795 39040 6796 39080
rect 6836 39040 6837 39080
rect 6795 39031 6837 39040
rect 8619 39080 8661 39089
rect 8619 39040 8620 39080
rect 8660 39040 8661 39080
rect 8619 39031 8661 39040
rect 12843 39080 12885 39089
rect 12843 39040 12844 39080
rect 12884 39040 12885 39080
rect 12843 39031 12885 39040
rect 16299 39080 16341 39089
rect 16299 39040 16300 39080
rect 16340 39040 16341 39080
rect 16299 39031 16341 39040
rect 18603 39080 18645 39089
rect 18603 39040 18604 39080
rect 18644 39040 18645 39080
rect 18603 39031 18645 39040
rect 1315 38996 1373 38997
rect 1315 38956 1324 38996
rect 1364 38956 1373 38996
rect 1315 38955 1373 38956
rect 4963 38996 5021 38997
rect 4963 38956 4972 38996
rect 5012 38956 5021 38996
rect 4963 38955 5021 38956
rect 5539 38996 5597 38997
rect 5539 38956 5548 38996
rect 5588 38956 5597 38996
rect 5539 38955 5597 38956
rect 6019 38996 6077 38997
rect 6019 38956 6028 38996
rect 6068 38956 6077 38996
rect 6019 38955 6077 38956
rect 6403 38996 6461 38997
rect 6403 38956 6412 38996
rect 6452 38956 6461 38996
rect 6403 38955 6461 38956
rect 6979 38996 7037 38997
rect 6979 38956 6988 38996
rect 7028 38956 7037 38996
rect 6979 38955 7037 38956
rect 11115 38996 11157 39005
rect 11115 38956 11116 38996
rect 11156 38956 11157 38996
rect 11115 38947 11157 38956
rect 13027 38996 13085 38997
rect 13027 38956 13036 38996
rect 13076 38956 13085 38996
rect 13027 38955 13085 38956
rect 14571 38996 14613 39005
rect 14571 38956 14572 38996
rect 14612 38956 14613 38996
rect 14571 38947 14613 38956
rect 14667 38996 14709 39005
rect 14667 38956 14668 38996
rect 14708 38956 14709 38996
rect 14667 38947 14709 38956
rect 19267 38996 19325 38997
rect 19267 38956 19276 38996
rect 19316 38956 19325 38996
rect 19267 38955 19325 38956
rect 19651 38996 19709 38997
rect 19651 38956 19660 38996
rect 19700 38956 19709 38996
rect 19651 38955 19709 38956
rect 20035 38996 20093 38997
rect 20035 38956 20044 38996
rect 20084 38956 20093 38996
rect 20035 38955 20093 38956
rect 15627 38926 15669 38935
rect 1699 38912 1757 38913
rect 1699 38872 1708 38912
rect 1748 38872 1757 38912
rect 1699 38871 1757 38872
rect 2947 38912 3005 38913
rect 2947 38872 2956 38912
rect 2996 38872 3005 38912
rect 2947 38871 3005 38872
rect 3331 38912 3389 38913
rect 3331 38872 3340 38912
rect 3380 38872 3389 38912
rect 3331 38871 3389 38872
rect 4579 38912 4637 38913
rect 4579 38872 4588 38912
rect 4628 38872 4637 38912
rect 4579 38871 4637 38872
rect 7171 38912 7229 38913
rect 7171 38872 7180 38912
rect 7220 38872 7229 38912
rect 7171 38871 7229 38872
rect 8419 38912 8477 38913
rect 8419 38872 8428 38912
rect 8468 38872 8477 38912
rect 8419 38871 8477 38872
rect 8803 38912 8861 38913
rect 8803 38872 8812 38912
rect 8852 38872 8861 38912
rect 8803 38871 8861 38872
rect 10051 38912 10109 38913
rect 10051 38872 10060 38912
rect 10100 38872 10109 38912
rect 10051 38871 10109 38872
rect 10539 38912 10581 38921
rect 10539 38872 10540 38912
rect 10580 38872 10581 38912
rect 10539 38863 10581 38872
rect 10635 38912 10677 38921
rect 10635 38872 10636 38912
rect 10676 38872 10677 38912
rect 10635 38863 10677 38872
rect 11019 38912 11061 38921
rect 12075 38917 12117 38926
rect 11019 38872 11020 38912
rect 11060 38872 11061 38912
rect 11019 38863 11061 38872
rect 11587 38912 11645 38913
rect 11587 38872 11596 38912
rect 11636 38872 11645 38912
rect 11587 38871 11645 38872
rect 12075 38877 12076 38917
rect 12116 38877 12117 38917
rect 12075 38868 12117 38877
rect 12547 38912 12605 38913
rect 12547 38872 12556 38912
rect 12596 38872 12605 38912
rect 12547 38871 12605 38872
rect 14091 38912 14133 38921
rect 14091 38872 14092 38912
rect 14132 38872 14133 38912
rect 14091 38863 14133 38872
rect 14187 38912 14229 38921
rect 14187 38872 14188 38912
rect 14228 38872 14229 38912
rect 14187 38863 14229 38872
rect 15139 38912 15197 38913
rect 15139 38872 15148 38912
rect 15188 38872 15197 38912
rect 15627 38886 15628 38926
rect 15668 38886 15669 38926
rect 15627 38877 15669 38886
rect 16011 38912 16053 38921
rect 15139 38871 15197 38872
rect 16011 38872 16012 38912
rect 16052 38872 16053 38912
rect 16011 38863 16053 38872
rect 16299 38912 16341 38921
rect 16299 38872 16300 38912
rect 16340 38872 16341 38912
rect 16299 38863 16341 38872
rect 16483 38912 16541 38913
rect 16483 38872 16492 38912
rect 16532 38872 16541 38912
rect 16483 38871 16541 38872
rect 17731 38912 17789 38913
rect 17731 38872 17740 38912
rect 17780 38872 17789 38912
rect 17731 38871 17789 38872
rect 18795 38912 18837 38921
rect 18795 38872 18796 38912
rect 18836 38872 18837 38912
rect 18795 38863 18837 38872
rect 18891 38912 18933 38921
rect 18891 38872 18892 38912
rect 18932 38872 18933 38912
rect 18891 38863 18933 38872
rect 18987 38912 19029 38921
rect 18987 38872 18988 38912
rect 19028 38872 19029 38912
rect 18987 38863 19029 38872
rect 10251 38828 10293 38837
rect 10251 38788 10252 38828
rect 10292 38788 10293 38828
rect 10251 38779 10293 38788
rect 3147 38744 3189 38753
rect 3147 38704 3148 38744
rect 3188 38704 3189 38744
rect 3147 38695 3189 38704
rect 4779 38744 4821 38753
rect 4779 38704 4780 38744
rect 4820 38704 4821 38744
rect 4779 38695 4821 38704
rect 5163 38744 5205 38753
rect 5163 38704 5164 38744
rect 5204 38704 5205 38744
rect 5163 38695 5205 38704
rect 12267 38744 12309 38753
rect 12267 38704 12268 38744
rect 12308 38704 12309 38744
rect 12267 38695 12309 38704
rect 15819 38744 15861 38753
rect 15819 38704 15820 38744
rect 15860 38704 15861 38744
rect 15819 38695 15861 38704
rect 17931 38744 17973 38753
rect 17931 38704 17932 38744
rect 17972 38704 17973 38744
rect 17931 38695 17973 38704
rect 18115 38744 18173 38745
rect 18115 38704 18124 38744
rect 18164 38704 18173 38744
rect 18115 38703 18173 38704
rect 18499 38744 18557 38745
rect 18499 38704 18508 38744
rect 18548 38704 18557 38744
rect 18499 38703 18557 38704
rect 19075 38744 19133 38745
rect 19075 38704 19084 38744
rect 19124 38704 19133 38744
rect 19075 38703 19133 38704
rect 19467 38744 19509 38753
rect 19467 38704 19468 38744
rect 19508 38704 19509 38744
rect 19467 38695 19509 38704
rect 19851 38744 19893 38753
rect 19851 38704 19852 38744
rect 19892 38704 19893 38744
rect 19851 38695 19893 38704
rect 20235 38744 20277 38753
rect 20235 38704 20236 38744
rect 20276 38704 20277 38744
rect 20235 38695 20277 38704
rect 1152 38576 20452 38600
rect 1152 38536 4928 38576
rect 4968 38536 5010 38576
rect 5050 38536 5092 38576
rect 5132 38536 5174 38576
rect 5214 38536 5256 38576
rect 5296 38536 20048 38576
rect 20088 38536 20130 38576
rect 20170 38536 20212 38576
rect 20252 38536 20294 38576
rect 20334 38536 20376 38576
rect 20416 38536 20452 38576
rect 1152 38512 20452 38536
rect 3147 38408 3189 38417
rect 3147 38368 3148 38408
rect 3188 38368 3189 38408
rect 3147 38359 3189 38368
rect 3531 38408 3573 38417
rect 3531 38368 3532 38408
rect 3572 38368 3573 38408
rect 3531 38359 3573 38368
rect 4011 38408 4053 38417
rect 4011 38368 4012 38408
rect 4052 38368 4053 38408
rect 4011 38359 4053 38368
rect 8035 38408 8093 38409
rect 8035 38368 8044 38408
rect 8084 38368 8093 38408
rect 8035 38367 8093 38368
rect 12075 38408 12117 38417
rect 12075 38368 12076 38408
rect 12116 38368 12117 38408
rect 12075 38359 12117 38368
rect 16299 38408 16341 38417
rect 16299 38368 16300 38408
rect 16340 38368 16341 38408
rect 16299 38359 16341 38368
rect 18315 38324 18357 38333
rect 18315 38284 18316 38324
rect 18356 38284 18357 38324
rect 18315 38275 18357 38284
rect 18987 38324 19029 38333
rect 18987 38284 18988 38324
rect 19028 38284 19029 38324
rect 18987 38275 19029 38284
rect 1219 38240 1277 38241
rect 1219 38200 1228 38240
rect 1268 38200 1277 38240
rect 1219 38199 1277 38200
rect 2467 38240 2525 38241
rect 2467 38200 2476 38240
rect 2516 38200 2525 38240
rect 2467 38199 2525 38200
rect 4387 38240 4445 38241
rect 4387 38200 4396 38240
rect 4436 38200 4445 38240
rect 4387 38199 4445 38200
rect 5635 38240 5693 38241
rect 5635 38200 5644 38240
rect 5684 38200 5693 38240
rect 5635 38199 5693 38200
rect 6403 38240 6461 38241
rect 6403 38200 6412 38240
rect 6452 38200 6461 38240
rect 6403 38199 6461 38200
rect 7651 38240 7709 38241
rect 7651 38200 7660 38240
rect 7700 38200 7709 38240
rect 7651 38199 7709 38200
rect 8611 38240 8669 38241
rect 8611 38200 8620 38240
rect 8660 38200 8669 38240
rect 8611 38199 8669 38200
rect 9859 38240 9917 38241
rect 9859 38200 9868 38240
rect 9908 38200 9917 38240
rect 9859 38199 9917 38200
rect 10627 38240 10685 38241
rect 10627 38200 10636 38240
rect 10676 38200 10685 38240
rect 10627 38199 10685 38200
rect 11875 38240 11933 38241
rect 11875 38200 11884 38240
rect 11924 38200 11933 38240
rect 11875 38199 11933 38200
rect 12835 38240 12893 38241
rect 12835 38200 12844 38240
rect 12884 38200 12893 38240
rect 12835 38199 12893 38200
rect 14083 38240 14141 38241
rect 14083 38200 14092 38240
rect 14132 38200 14141 38240
rect 14083 38199 14141 38200
rect 14467 38240 14525 38241
rect 14467 38200 14476 38240
rect 14516 38200 14525 38240
rect 14467 38199 14525 38200
rect 15715 38240 15773 38241
rect 15715 38200 15724 38240
rect 15764 38200 15773 38240
rect 15715 38199 15773 38200
rect 16587 38240 16629 38249
rect 16587 38200 16588 38240
rect 16628 38200 16629 38240
rect 16587 38191 16629 38200
rect 16683 38240 16725 38249
rect 16683 38200 16684 38240
rect 16724 38200 16725 38240
rect 16683 38191 16725 38200
rect 17635 38240 17693 38241
rect 17635 38200 17644 38240
rect 17684 38200 17693 38240
rect 17635 38199 17693 38200
rect 18123 38235 18165 38244
rect 18123 38195 18124 38235
rect 18164 38195 18165 38235
rect 18595 38240 18653 38241
rect 18595 38200 18604 38240
rect 18644 38200 18653 38240
rect 18595 38199 18653 38200
rect 18891 38240 18933 38249
rect 18891 38200 18892 38240
rect 18932 38200 18933 38240
rect 18123 38186 18165 38195
rect 18891 38191 18933 38200
rect 19755 38240 19797 38249
rect 19755 38200 19756 38240
rect 19796 38200 19797 38240
rect 19755 38191 19797 38200
rect 19851 38240 19893 38249
rect 19851 38200 19852 38240
rect 19892 38200 19893 38240
rect 19851 38191 19893 38200
rect 20131 38240 20189 38241
rect 20131 38200 20140 38240
rect 20180 38200 20189 38240
rect 20131 38199 20189 38200
rect 2947 38156 3005 38157
rect 2947 38116 2956 38156
rect 2996 38116 3005 38156
rect 2947 38115 3005 38116
rect 3331 38156 3389 38157
rect 3331 38116 3340 38156
rect 3380 38116 3389 38156
rect 3331 38115 3389 38116
rect 3811 38156 3869 38157
rect 3811 38116 3820 38156
rect 3860 38116 3869 38156
rect 3811 38115 3869 38116
rect 16099 38156 16157 38157
rect 16099 38116 16108 38156
rect 16148 38116 16157 38156
rect 16099 38115 16157 38116
rect 17067 38156 17109 38165
rect 17067 38116 17068 38156
rect 17108 38116 17109 38156
rect 17067 38107 17109 38116
rect 17163 38156 17205 38165
rect 17163 38116 17164 38156
rect 17204 38116 17205 38156
rect 17163 38107 17205 38116
rect 6027 38072 6069 38081
rect 6027 38032 6028 38072
rect 6068 38032 6069 38072
rect 6027 38023 6069 38032
rect 8331 38072 8373 38081
rect 8331 38032 8332 38072
rect 8372 38032 8373 38072
rect 8331 38023 8373 38032
rect 19459 38072 19517 38073
rect 19459 38032 19468 38072
rect 19508 38032 19517 38072
rect 19459 38031 19517 38032
rect 2667 37988 2709 37997
rect 2667 37948 2668 37988
rect 2708 37948 2709 37988
rect 2667 37939 2709 37948
rect 4203 37988 4245 37997
rect 4203 37948 4204 37988
rect 4244 37948 4245 37988
rect 4203 37939 4245 37948
rect 7851 37988 7893 37997
rect 7851 37948 7852 37988
rect 7892 37948 7893 37988
rect 7851 37939 7893 37948
rect 10059 37988 10101 37997
rect 10059 37948 10060 37988
rect 10100 37948 10101 37988
rect 10059 37939 10101 37948
rect 14283 37988 14325 37997
rect 14283 37948 14284 37988
rect 14324 37948 14325 37988
rect 14283 37939 14325 37948
rect 15915 37988 15957 37997
rect 15915 37948 15916 37988
rect 15956 37948 15957 37988
rect 15915 37939 15957 37948
rect 19267 37988 19325 37989
rect 19267 37948 19276 37988
rect 19316 37948 19325 37988
rect 19267 37947 19325 37948
rect 1152 37820 20352 37844
rect 1152 37780 3688 37820
rect 3728 37780 3770 37820
rect 3810 37780 3852 37820
rect 3892 37780 3934 37820
rect 3974 37780 4016 37820
rect 4056 37780 18808 37820
rect 18848 37780 18890 37820
rect 18930 37780 18972 37820
rect 19012 37780 19054 37820
rect 19094 37780 19136 37820
rect 19176 37780 20352 37820
rect 1152 37756 20352 37780
rect 1611 37652 1653 37661
rect 1611 37612 1612 37652
rect 1652 37612 1653 37652
rect 1611 37603 1653 37612
rect 1995 37652 2037 37661
rect 1995 37612 1996 37652
rect 2036 37612 2037 37652
rect 1995 37603 2037 37612
rect 6987 37652 7029 37661
rect 6987 37612 6988 37652
rect 7028 37612 7029 37652
rect 6987 37603 7029 37612
rect 17643 37652 17685 37661
rect 17643 37612 17644 37652
rect 17684 37612 17685 37652
rect 17643 37603 17685 37612
rect 18315 37652 18357 37661
rect 18315 37612 18316 37652
rect 18356 37612 18357 37652
rect 18315 37603 18357 37612
rect 19179 37652 19221 37661
rect 19179 37612 19180 37652
rect 19220 37612 19221 37652
rect 19179 37603 19221 37612
rect 4395 37568 4437 37577
rect 4395 37528 4396 37568
rect 4436 37528 4437 37568
rect 4395 37519 4437 37528
rect 1411 37484 1469 37485
rect 1411 37444 1420 37484
rect 1460 37444 1469 37484
rect 1411 37443 1469 37444
rect 1795 37484 1853 37485
rect 1795 37444 1804 37484
rect 1844 37444 1853 37484
rect 1795 37443 1853 37444
rect 7171 37484 7229 37485
rect 7171 37444 7180 37484
rect 7220 37444 7229 37484
rect 7171 37443 7229 37444
rect 9003 37484 9045 37493
rect 9003 37444 9004 37484
rect 9044 37444 9045 37484
rect 18115 37484 18173 37485
rect 9003 37435 9045 37444
rect 15675 37442 15717 37451
rect 18115 37444 18124 37484
rect 18164 37444 18173 37484
rect 18115 37443 18173 37444
rect 20035 37484 20093 37485
rect 20035 37444 20044 37484
rect 20084 37444 20093 37484
rect 20035 37443 20093 37444
rect 3819 37414 3861 37423
rect 2283 37400 2325 37409
rect 2283 37360 2284 37400
rect 2324 37360 2325 37400
rect 2283 37351 2325 37360
rect 2379 37400 2421 37409
rect 2379 37360 2380 37400
rect 2420 37360 2421 37400
rect 2379 37351 2421 37360
rect 2763 37400 2805 37409
rect 2763 37360 2764 37400
rect 2804 37360 2805 37400
rect 2763 37351 2805 37360
rect 2859 37400 2901 37409
rect 2859 37360 2860 37400
rect 2900 37360 2901 37400
rect 2859 37351 2901 37360
rect 3331 37400 3389 37401
rect 3331 37360 3340 37400
rect 3380 37360 3389 37400
rect 3819 37374 3820 37414
rect 3860 37374 3861 37414
rect 6603 37414 6645 37423
rect 3819 37365 3861 37374
rect 5067 37400 5109 37409
rect 3331 37359 3389 37360
rect 5067 37360 5068 37400
rect 5108 37360 5109 37400
rect 5067 37351 5109 37360
rect 5163 37400 5205 37409
rect 5163 37360 5164 37400
rect 5204 37360 5205 37400
rect 5163 37351 5205 37360
rect 5547 37400 5589 37409
rect 5547 37360 5548 37400
rect 5588 37360 5589 37400
rect 5547 37351 5589 37360
rect 5643 37400 5685 37409
rect 5643 37360 5644 37400
rect 5684 37360 5685 37400
rect 5643 37351 5685 37360
rect 6115 37400 6173 37401
rect 6115 37360 6124 37400
rect 6164 37360 6173 37400
rect 6603 37374 6604 37414
rect 6644 37374 6645 37414
rect 9963 37414 10005 37423
rect 6603 37365 6645 37374
rect 7371 37400 7413 37409
rect 6115 37359 6173 37360
rect 7371 37360 7372 37400
rect 7412 37360 7413 37400
rect 7371 37351 7413 37360
rect 7659 37400 7701 37409
rect 7659 37360 7660 37400
rect 7700 37360 7701 37400
rect 7659 37351 7701 37360
rect 7939 37400 7997 37401
rect 7939 37360 7948 37400
rect 7988 37360 7997 37400
rect 7939 37359 7997 37360
rect 8427 37400 8469 37409
rect 8427 37360 8428 37400
rect 8468 37360 8469 37400
rect 8427 37351 8469 37360
rect 8523 37400 8565 37409
rect 8523 37360 8524 37400
rect 8564 37360 8565 37400
rect 8523 37351 8565 37360
rect 8907 37400 8949 37409
rect 8907 37360 8908 37400
rect 8948 37360 8949 37400
rect 8907 37351 8949 37360
rect 9475 37400 9533 37401
rect 9475 37360 9484 37400
rect 9524 37360 9533 37400
rect 9963 37374 9964 37414
rect 10004 37374 10005 37414
rect 9963 37365 10005 37374
rect 11491 37400 11549 37401
rect 9475 37359 9533 37360
rect 11491 37360 11500 37400
rect 11540 37360 11549 37400
rect 11491 37359 11549 37360
rect 12739 37400 12797 37401
rect 12739 37360 12748 37400
rect 12788 37360 12797 37400
rect 12739 37359 12797 37360
rect 14091 37400 14133 37409
rect 14091 37360 14092 37400
rect 14132 37360 14133 37400
rect 14091 37351 14133 37360
rect 14187 37400 14229 37409
rect 14187 37360 14188 37400
rect 14228 37360 14229 37400
rect 14187 37351 14229 37360
rect 14571 37400 14613 37409
rect 14571 37360 14572 37400
rect 14612 37360 14613 37400
rect 14571 37351 14613 37360
rect 14667 37400 14709 37409
rect 15675 37402 15676 37442
rect 15716 37402 15717 37442
rect 14667 37360 14668 37400
rect 14708 37360 14709 37400
rect 14667 37351 14709 37360
rect 15139 37400 15197 37401
rect 15139 37360 15148 37400
rect 15188 37360 15197 37400
rect 15675 37393 15717 37402
rect 16195 37400 16253 37401
rect 15139 37359 15197 37360
rect 16195 37360 16204 37400
rect 16244 37360 16253 37400
rect 16195 37359 16253 37360
rect 17443 37400 17501 37401
rect 17443 37360 17452 37400
rect 17492 37360 17501 37400
rect 17443 37359 17501 37360
rect 18987 37400 19029 37409
rect 18987 37360 18988 37400
rect 19028 37360 19029 37400
rect 18987 37351 19029 37360
rect 4011 37316 4053 37325
rect 4011 37276 4012 37316
rect 4052 37276 4053 37316
rect 4011 37267 4053 37276
rect 6795 37316 6837 37325
rect 6795 37276 6796 37316
rect 6836 37276 6837 37316
rect 6795 37267 6837 37276
rect 4675 37232 4733 37233
rect 4675 37192 4684 37232
rect 4724 37192 4733 37232
rect 4675 37191 4733 37192
rect 7467 37232 7509 37241
rect 7467 37192 7468 37232
rect 7508 37192 7509 37232
rect 7467 37183 7509 37192
rect 7843 37232 7901 37233
rect 7843 37192 7852 37232
rect 7892 37192 7901 37232
rect 7843 37191 7901 37192
rect 8131 37232 8189 37233
rect 8131 37192 8140 37232
rect 8180 37192 8189 37232
rect 8131 37191 8189 37192
rect 10155 37232 10197 37241
rect 10155 37192 10156 37232
rect 10196 37192 10197 37232
rect 10155 37183 10197 37192
rect 12939 37232 12981 37241
rect 12939 37192 12940 37232
rect 12980 37192 12981 37232
rect 12939 37183 12981 37192
rect 15819 37232 15861 37241
rect 15819 37192 15820 37232
rect 15860 37192 15861 37232
rect 15819 37183 15861 37192
rect 18499 37232 18557 37233
rect 18499 37192 18508 37232
rect 18548 37192 18557 37232
rect 18499 37191 18557 37192
rect 20235 37232 20277 37241
rect 20235 37192 20236 37232
rect 20276 37192 20277 37232
rect 20235 37183 20277 37192
rect 1152 37064 20452 37088
rect 1152 37024 4928 37064
rect 4968 37024 5010 37064
rect 5050 37024 5092 37064
rect 5132 37024 5174 37064
rect 5214 37024 5256 37064
rect 5296 37024 20048 37064
rect 20088 37024 20130 37064
rect 20170 37024 20212 37064
rect 20252 37024 20294 37064
rect 20334 37024 20376 37064
rect 20416 37024 20452 37064
rect 1152 37000 20452 37024
rect 8323 36896 8381 36897
rect 8323 36856 8332 36896
rect 8372 36856 8381 36896
rect 8323 36855 8381 36856
rect 16587 36896 16629 36905
rect 16587 36856 16588 36896
rect 16628 36856 16629 36896
rect 16587 36847 16629 36856
rect 18115 36896 18173 36897
rect 18115 36856 18124 36896
rect 18164 36856 18173 36896
rect 18115 36855 18173 36856
rect 18411 36896 18453 36905
rect 18411 36856 18412 36896
rect 18452 36856 18453 36896
rect 18411 36847 18453 36856
rect 6123 36812 6165 36821
rect 6123 36772 6124 36812
rect 6164 36772 6165 36812
rect 6123 36763 6165 36772
rect 8139 36812 8181 36821
rect 8139 36772 8140 36812
rect 8180 36772 8181 36812
rect 8139 36763 8181 36772
rect 12939 36812 12981 36821
rect 12939 36772 12940 36812
rect 12980 36772 12981 36812
rect 12939 36763 12981 36772
rect 1219 36728 1277 36729
rect 1219 36688 1228 36728
rect 1268 36688 1277 36728
rect 1219 36687 1277 36688
rect 2467 36728 2525 36729
rect 2467 36688 2476 36728
rect 2516 36688 2525 36728
rect 2467 36687 2525 36688
rect 4291 36728 4349 36729
rect 4291 36688 4300 36728
rect 4340 36688 4349 36728
rect 4291 36687 4349 36688
rect 4675 36728 4733 36729
rect 4675 36688 4684 36728
rect 4724 36688 4733 36728
rect 4675 36687 4733 36688
rect 5923 36728 5981 36729
rect 5923 36688 5932 36728
rect 5972 36688 5981 36728
rect 5923 36687 5981 36688
rect 6411 36728 6453 36737
rect 6411 36688 6412 36728
rect 6452 36688 6453 36728
rect 3043 36686 3101 36687
rect 3043 36646 3052 36686
rect 3092 36646 3101 36686
rect 6411 36679 6453 36688
rect 6507 36728 6549 36737
rect 6507 36688 6508 36728
rect 6548 36688 6549 36728
rect 6507 36679 6549 36688
rect 7459 36728 7517 36729
rect 7459 36688 7468 36728
rect 7508 36688 7517 36728
rect 8619 36728 8661 36737
rect 7459 36687 7517 36688
rect 7995 36686 8037 36695
rect 3043 36645 3101 36646
rect 6891 36644 6933 36653
rect 6891 36604 6892 36644
rect 6932 36604 6933 36644
rect 6891 36595 6933 36604
rect 6987 36644 7029 36653
rect 6987 36604 6988 36644
rect 7028 36604 7029 36644
rect 7995 36646 7996 36686
rect 8036 36646 8037 36686
rect 8619 36688 8620 36728
rect 8660 36688 8661 36728
rect 8619 36679 8661 36688
rect 8907 36728 8949 36737
rect 8907 36688 8908 36728
rect 8948 36688 8949 36728
rect 8907 36679 8949 36688
rect 9475 36728 9533 36729
rect 9475 36688 9484 36728
rect 9524 36688 9533 36728
rect 9475 36687 9533 36688
rect 10723 36728 10781 36729
rect 10723 36688 10732 36728
rect 10772 36688 10781 36728
rect 10723 36687 10781 36688
rect 11211 36728 11253 36737
rect 11211 36688 11212 36728
rect 11252 36688 11253 36728
rect 11211 36679 11253 36688
rect 11307 36728 11349 36737
rect 11307 36688 11308 36728
rect 11348 36688 11349 36728
rect 11307 36679 11349 36688
rect 12259 36728 12317 36729
rect 12259 36688 12268 36728
rect 12308 36688 12317 36728
rect 15139 36728 15197 36729
rect 12259 36687 12317 36688
rect 12795 36718 12837 36727
rect 12795 36678 12796 36718
rect 12836 36678 12837 36718
rect 15139 36688 15148 36728
rect 15188 36688 15197 36728
rect 15139 36687 15197 36688
rect 16387 36728 16445 36729
rect 16387 36688 16396 36728
rect 16436 36688 16445 36728
rect 16387 36687 16445 36688
rect 17347 36728 17405 36729
rect 17347 36688 17356 36728
rect 17396 36688 17405 36728
rect 17347 36687 17405 36688
rect 17451 36728 17493 36737
rect 17451 36688 17452 36728
rect 17492 36688 17493 36728
rect 17451 36679 17493 36688
rect 17643 36728 17685 36737
rect 17643 36688 17644 36728
rect 17684 36688 17685 36728
rect 17643 36679 17685 36688
rect 18595 36728 18653 36729
rect 18595 36688 18604 36728
rect 18644 36688 18653 36728
rect 18595 36687 18653 36688
rect 19843 36728 19901 36729
rect 19843 36688 19852 36728
rect 19892 36688 19901 36728
rect 19843 36687 19901 36688
rect 12795 36669 12837 36678
rect 7995 36637 8037 36646
rect 11691 36644 11733 36653
rect 6987 36595 7029 36604
rect 11691 36604 11692 36644
rect 11732 36604 11733 36644
rect 11691 36595 11733 36604
rect 11787 36644 11829 36653
rect 11787 36604 11788 36644
rect 11828 36604 11829 36644
rect 11787 36595 11829 36604
rect 16963 36644 17021 36645
rect 16963 36604 16972 36644
rect 17012 36604 17021 36644
rect 16963 36603 17021 36604
rect 20035 36644 20093 36645
rect 20035 36604 20044 36644
rect 20084 36604 20093 36644
rect 20035 36603 20093 36604
rect 8427 36560 8469 36569
rect 8427 36520 8428 36560
rect 8468 36520 8469 36560
rect 8427 36511 8469 36520
rect 17163 36560 17205 36569
rect 17163 36520 17164 36560
rect 17204 36520 17205 36560
rect 17163 36511 17205 36520
rect 17643 36560 17685 36569
rect 17643 36520 17644 36560
rect 17684 36520 17685 36560
rect 17643 36511 17685 36520
rect 18219 36560 18261 36569
rect 18219 36520 18220 36560
rect 18260 36520 18261 36560
rect 18219 36511 18261 36520
rect 2667 36476 2709 36485
rect 2667 36436 2668 36476
rect 2708 36436 2709 36476
rect 2667 36427 2709 36436
rect 4491 36476 4533 36485
rect 4491 36436 4492 36476
rect 4532 36436 4533 36476
rect 4491 36427 4533 36436
rect 8907 36476 8949 36485
rect 8907 36436 8908 36476
rect 8948 36436 8949 36476
rect 8907 36427 8949 36436
rect 10923 36476 10965 36485
rect 10923 36436 10924 36476
rect 10964 36436 10965 36476
rect 10923 36427 10965 36436
rect 20235 36476 20277 36485
rect 20235 36436 20236 36476
rect 20276 36436 20277 36476
rect 20235 36427 20277 36436
rect 1152 36308 20352 36332
rect 1152 36268 3688 36308
rect 3728 36268 3770 36308
rect 3810 36268 3852 36308
rect 3892 36268 3934 36308
rect 3974 36268 4016 36308
rect 4056 36268 18808 36308
rect 18848 36268 18890 36308
rect 18930 36268 18972 36308
rect 19012 36268 19054 36308
rect 19094 36268 19136 36308
rect 19176 36268 20352 36308
rect 1152 36244 20352 36268
rect 1611 36140 1653 36149
rect 1611 36100 1612 36140
rect 1652 36100 1653 36140
rect 1611 36091 1653 36100
rect 8235 36140 8277 36149
rect 8235 36100 8236 36140
rect 8276 36100 8277 36140
rect 8235 36091 8277 36100
rect 11019 36140 11061 36149
rect 11019 36100 11020 36140
rect 11060 36100 11061 36140
rect 11019 36091 11061 36100
rect 17451 36140 17493 36149
rect 17451 36100 17452 36140
rect 17492 36100 17493 36140
rect 17451 36091 17493 36100
rect 17835 36140 17877 36149
rect 17835 36100 17836 36140
rect 17876 36100 17877 36140
rect 17835 36091 17877 36100
rect 19467 36140 19509 36149
rect 19467 36100 19468 36140
rect 19508 36100 19509 36140
rect 19467 36091 19509 36100
rect 8427 36056 8469 36065
rect 8427 36016 8428 36056
rect 8468 36016 8469 36056
rect 8427 36007 8469 36016
rect 9195 36056 9237 36065
rect 9195 36016 9196 36056
rect 9236 36016 9237 36056
rect 9195 36007 9237 36016
rect 1411 35972 1469 35973
rect 1411 35932 1420 35972
rect 1460 35932 1469 35972
rect 1411 35931 1469 35932
rect 4971 35972 5013 35981
rect 4971 35932 4972 35972
rect 5012 35932 5013 35972
rect 4971 35923 5013 35932
rect 9099 35972 9141 35981
rect 9099 35932 9100 35972
rect 9140 35932 9141 35972
rect 9099 35923 9141 35932
rect 9291 35972 9333 35981
rect 9291 35932 9292 35972
rect 9332 35932 9333 35972
rect 17251 35972 17309 35973
rect 9291 35923 9333 35932
rect 11883 35930 11925 35939
rect 17251 35932 17260 35972
rect 17300 35932 17309 35972
rect 17251 35931 17309 35932
rect 17635 35972 17693 35973
rect 17635 35932 17644 35972
rect 17684 35932 17693 35972
rect 17635 35931 17693 35932
rect 3435 35902 3477 35911
rect 10819 35909 10877 35910
rect 1899 35888 1941 35897
rect 1899 35848 1900 35888
rect 1940 35848 1941 35888
rect 1899 35839 1941 35848
rect 1995 35888 2037 35897
rect 1995 35848 1996 35888
rect 2036 35848 2037 35888
rect 1995 35839 2037 35848
rect 2379 35888 2421 35897
rect 2379 35848 2380 35888
rect 2420 35848 2421 35888
rect 2379 35839 2421 35848
rect 2475 35888 2517 35897
rect 2475 35848 2476 35888
rect 2516 35848 2517 35888
rect 2475 35839 2517 35848
rect 2947 35888 3005 35889
rect 2947 35848 2956 35888
rect 2996 35848 3005 35888
rect 3435 35862 3436 35902
rect 3476 35862 3477 35902
rect 3435 35853 3477 35862
rect 4395 35888 4437 35897
rect 2947 35847 3005 35848
rect 4395 35848 4396 35888
rect 4436 35848 4437 35888
rect 4395 35839 4437 35848
rect 4491 35888 4533 35897
rect 4491 35848 4492 35888
rect 4532 35848 4533 35888
rect 4491 35839 4533 35848
rect 4875 35888 4917 35897
rect 5931 35893 5973 35902
rect 4875 35848 4876 35888
rect 4916 35848 4917 35888
rect 4875 35839 4917 35848
rect 5443 35888 5501 35889
rect 5443 35848 5452 35888
rect 5492 35848 5501 35888
rect 5443 35847 5501 35848
rect 5931 35853 5932 35893
rect 5972 35853 5973 35893
rect 5931 35844 5973 35853
rect 6411 35888 6453 35897
rect 6411 35848 6412 35888
rect 6452 35848 6453 35888
rect 6411 35839 6453 35848
rect 6507 35888 6549 35897
rect 6507 35848 6508 35888
rect 6548 35848 6549 35888
rect 6507 35839 6549 35848
rect 6603 35888 6645 35897
rect 6603 35848 6604 35888
rect 6644 35848 6645 35888
rect 6603 35839 6645 35848
rect 6787 35888 6845 35889
rect 6787 35848 6796 35888
rect 6836 35848 6845 35888
rect 6787 35847 6845 35848
rect 8035 35888 8093 35889
rect 8035 35848 8044 35888
rect 8084 35848 8093 35888
rect 8035 35847 8093 35848
rect 8995 35888 9053 35889
rect 8995 35848 9004 35888
rect 9044 35848 9053 35888
rect 8995 35847 9053 35848
rect 9387 35888 9429 35897
rect 9387 35848 9388 35888
rect 9428 35848 9429 35888
rect 9387 35839 9429 35848
rect 9571 35888 9629 35889
rect 9571 35848 9580 35888
rect 9620 35848 9629 35888
rect 10819 35869 10828 35909
rect 10868 35869 10877 35909
rect 10819 35868 10877 35869
rect 11307 35888 11349 35897
rect 9571 35847 9629 35848
rect 11307 35848 11308 35888
rect 11348 35848 11349 35888
rect 11307 35839 11349 35848
rect 11403 35888 11445 35897
rect 11403 35848 11404 35888
rect 11444 35848 11445 35888
rect 11403 35839 11445 35848
rect 11787 35888 11829 35897
rect 11787 35848 11788 35888
rect 11828 35848 11829 35888
rect 11883 35890 11884 35930
rect 11924 35890 11925 35930
rect 11883 35881 11925 35890
rect 12891 35897 12933 35906
rect 16923 35897 16965 35906
rect 12355 35888 12413 35889
rect 11787 35839 11829 35848
rect 12355 35848 12364 35888
rect 12404 35848 12413 35888
rect 12891 35857 12892 35897
rect 12932 35857 12933 35897
rect 12891 35848 12933 35857
rect 15339 35888 15381 35897
rect 15339 35848 15340 35888
rect 15380 35848 15381 35888
rect 12355 35847 12413 35848
rect 15339 35839 15381 35848
rect 15435 35888 15477 35897
rect 15435 35848 15436 35888
rect 15476 35848 15477 35888
rect 15435 35839 15477 35848
rect 15819 35888 15861 35897
rect 15819 35848 15820 35888
rect 15860 35848 15861 35888
rect 15819 35839 15861 35848
rect 15915 35888 15957 35897
rect 15915 35848 15916 35888
rect 15956 35848 15957 35888
rect 15915 35839 15957 35848
rect 16387 35888 16445 35889
rect 16387 35848 16396 35888
rect 16436 35848 16445 35888
rect 16923 35857 16924 35897
rect 16964 35857 16965 35897
rect 16923 35848 16965 35857
rect 18019 35888 18077 35889
rect 18019 35848 18028 35888
rect 18068 35848 18077 35888
rect 16387 35847 16445 35848
rect 18019 35847 18077 35848
rect 19267 35888 19325 35889
rect 19267 35848 19276 35888
rect 19316 35848 19325 35888
rect 19267 35847 19325 35848
rect 19755 35888 19797 35897
rect 19755 35848 19756 35888
rect 19796 35848 19797 35888
rect 19755 35839 19797 35848
rect 19851 35888 19893 35897
rect 19851 35848 19852 35888
rect 19892 35848 19893 35888
rect 19851 35839 19893 35848
rect 19947 35888 19989 35897
rect 19947 35848 19948 35888
rect 19988 35848 19989 35888
rect 19947 35839 19989 35848
rect 17067 35804 17109 35813
rect 17067 35764 17068 35804
rect 17108 35764 17109 35804
rect 17067 35755 17109 35764
rect 3627 35720 3669 35729
rect 3627 35680 3628 35720
rect 3668 35680 3669 35720
rect 3627 35671 3669 35680
rect 4003 35720 4061 35721
rect 4003 35680 4012 35720
rect 4052 35680 4061 35720
rect 4003 35679 4061 35680
rect 6123 35720 6165 35729
rect 6123 35680 6124 35720
rect 6164 35680 6165 35720
rect 6123 35671 6165 35680
rect 6307 35720 6365 35721
rect 6307 35680 6316 35720
rect 6356 35680 6365 35720
rect 6307 35679 6365 35680
rect 8523 35720 8565 35729
rect 8523 35680 8524 35720
rect 8564 35680 8565 35720
rect 8523 35671 8565 35680
rect 13035 35720 13077 35729
rect 13035 35680 13036 35720
rect 13076 35680 13077 35720
rect 13035 35671 13077 35680
rect 19467 35720 19509 35729
rect 19467 35680 19468 35720
rect 19508 35680 19509 35720
rect 19467 35671 19509 35680
rect 20139 35720 20181 35729
rect 20139 35680 20140 35720
rect 20180 35680 20181 35720
rect 20139 35671 20181 35680
rect 1152 35552 20452 35576
rect 1152 35512 4928 35552
rect 4968 35512 5010 35552
rect 5050 35512 5092 35552
rect 5132 35512 5174 35552
rect 5214 35512 5256 35552
rect 5296 35512 20048 35552
rect 20088 35512 20130 35552
rect 20170 35512 20212 35552
rect 20252 35512 20294 35552
rect 20334 35512 20376 35552
rect 20416 35512 20452 35552
rect 1152 35488 20452 35512
rect 5835 35384 5877 35393
rect 5835 35344 5836 35384
rect 5876 35344 5877 35384
rect 5835 35335 5877 35344
rect 7467 35384 7509 35393
rect 7467 35344 7468 35384
rect 7508 35344 7509 35384
rect 7467 35335 7509 35344
rect 10155 35388 10197 35397
rect 10155 35348 10156 35388
rect 10196 35348 10197 35388
rect 10155 35339 10197 35348
rect 13323 35384 13365 35393
rect 13323 35344 13324 35384
rect 13364 35344 13365 35384
rect 13323 35335 13365 35344
rect 15147 35384 15189 35393
rect 15147 35344 15148 35384
rect 15188 35344 15189 35384
rect 15147 35335 15189 35344
rect 8043 35300 8085 35309
rect 8043 35260 8044 35300
rect 8084 35260 8085 35300
rect 8043 35251 8085 35260
rect 10827 35300 10869 35309
rect 10827 35260 10828 35300
rect 10868 35260 10869 35300
rect 10827 35251 10869 35260
rect 17163 35300 17205 35309
rect 17163 35260 17164 35300
rect 17204 35260 17205 35300
rect 17163 35251 17205 35260
rect 19755 35300 19797 35309
rect 19755 35260 19756 35300
rect 19796 35260 19797 35300
rect 19755 35251 19797 35260
rect 20139 35237 20181 35246
rect 2083 35216 2141 35217
rect 2083 35176 2092 35216
rect 2132 35176 2141 35216
rect 2083 35175 2141 35176
rect 3331 35216 3389 35217
rect 3331 35176 3340 35216
rect 3380 35176 3389 35216
rect 3331 35175 3389 35176
rect 4387 35216 4445 35217
rect 4387 35176 4396 35216
rect 4436 35176 4445 35216
rect 4387 35175 4445 35176
rect 5635 35216 5693 35217
rect 5635 35176 5644 35216
rect 5684 35176 5693 35216
rect 5635 35175 5693 35176
rect 6019 35216 6077 35217
rect 6019 35176 6028 35216
rect 6068 35176 6077 35216
rect 6019 35175 6077 35176
rect 7267 35216 7325 35217
rect 7267 35176 7276 35216
rect 7316 35176 7325 35216
rect 7267 35175 7325 35176
rect 7947 35216 7989 35225
rect 7947 35176 7948 35216
rect 7988 35176 7989 35216
rect 7947 35167 7989 35176
rect 8139 35216 8181 35225
rect 8139 35176 8140 35216
rect 8180 35176 8181 35216
rect 8139 35167 8181 35176
rect 8227 35216 8285 35217
rect 8227 35176 8236 35216
rect 8276 35176 8285 35216
rect 8227 35175 8285 35176
rect 8811 35216 8853 35225
rect 8811 35176 8812 35216
rect 8852 35176 8853 35216
rect 8707 35174 8765 35175
rect 8707 35134 8716 35174
rect 8756 35134 8765 35174
rect 8811 35167 8853 35176
rect 9091 35216 9149 35217
rect 9091 35176 9100 35216
rect 9140 35176 9149 35216
rect 9091 35175 9149 35176
rect 9470 35216 9528 35217
rect 9470 35176 9479 35216
rect 9519 35176 9528 35216
rect 9470 35175 9528 35176
rect 9579 35216 9621 35225
rect 9579 35176 9580 35216
rect 9620 35176 9621 35216
rect 9579 35167 9621 35176
rect 9675 35216 9717 35225
rect 9675 35176 9676 35216
rect 9716 35176 9717 35216
rect 9675 35167 9717 35176
rect 9859 35216 9917 35217
rect 9859 35176 9868 35216
rect 9908 35176 9917 35216
rect 9859 35175 9917 35176
rect 9955 35216 10013 35217
rect 9955 35176 9964 35216
rect 10004 35176 10013 35216
rect 9955 35175 10013 35176
rect 10243 35216 10301 35217
rect 10243 35176 10252 35216
rect 10292 35176 10301 35216
rect 10243 35175 10301 35176
rect 10347 35216 10389 35225
rect 10347 35176 10348 35216
rect 10388 35176 10389 35216
rect 10347 35167 10389 35176
rect 11019 35216 11061 35225
rect 11019 35176 11020 35216
rect 11060 35176 11061 35216
rect 10915 35174 10973 35175
rect 8707 35133 8765 35134
rect 10915 35134 10924 35174
rect 10964 35134 10973 35174
rect 11019 35167 11061 35176
rect 11115 35216 11157 35225
rect 11115 35176 11116 35216
rect 11156 35176 11157 35216
rect 11115 35167 11157 35176
rect 11307 35216 11349 35225
rect 11307 35176 11308 35216
rect 11348 35176 11349 35216
rect 11307 35167 11349 35176
rect 11499 35216 11541 35225
rect 11499 35176 11500 35216
rect 11540 35176 11541 35216
rect 11499 35167 11541 35176
rect 11875 35216 11933 35217
rect 11875 35176 11884 35216
rect 11924 35176 11933 35216
rect 11875 35175 11933 35176
rect 13123 35216 13181 35217
rect 13123 35176 13132 35216
rect 13172 35176 13181 35216
rect 13123 35175 13181 35176
rect 13699 35216 13757 35217
rect 13699 35176 13708 35216
rect 13748 35176 13757 35216
rect 13699 35175 13757 35176
rect 14947 35216 15005 35217
rect 14947 35176 14956 35216
rect 14996 35176 15005 35216
rect 14947 35175 15005 35176
rect 15435 35216 15477 35225
rect 15435 35176 15436 35216
rect 15476 35176 15477 35216
rect 15435 35167 15477 35176
rect 15531 35216 15573 35225
rect 15531 35176 15532 35216
rect 15572 35176 15573 35216
rect 15531 35167 15573 35176
rect 16483 35216 16541 35217
rect 16483 35176 16492 35216
rect 16532 35176 16541 35216
rect 18027 35216 18069 35225
rect 16483 35175 16541 35176
rect 16971 35202 17013 35211
rect 16971 35162 16972 35202
rect 17012 35162 17013 35202
rect 18027 35176 18028 35216
rect 18068 35176 18069 35216
rect 18027 35167 18069 35176
rect 18123 35216 18165 35225
rect 18123 35176 18124 35216
rect 18164 35176 18165 35216
rect 18123 35167 18165 35176
rect 18507 35216 18549 35225
rect 18507 35176 18508 35216
rect 18548 35176 18549 35216
rect 18507 35167 18549 35176
rect 19075 35216 19133 35217
rect 19075 35176 19084 35216
rect 19124 35176 19133 35216
rect 19075 35175 19133 35176
rect 19563 35211 19605 35220
rect 19563 35171 19564 35211
rect 19604 35171 19605 35211
rect 19563 35162 19605 35171
rect 19947 35216 19989 35225
rect 19947 35176 19948 35216
rect 19988 35176 19989 35216
rect 19947 35167 19989 35176
rect 20043 35216 20085 35225
rect 20043 35176 20044 35216
rect 20084 35176 20085 35216
rect 20139 35197 20140 35237
rect 20180 35197 20181 35237
rect 20139 35188 20181 35197
rect 20235 35216 20277 35225
rect 20043 35167 20085 35176
rect 20235 35176 20236 35216
rect 20276 35176 20277 35216
rect 20235 35167 20277 35176
rect 16971 35153 17013 35162
rect 10915 35133 10973 35134
rect 1507 35132 1565 35133
rect 1507 35092 1516 35132
rect 1556 35092 1565 35132
rect 1507 35091 1565 35092
rect 4003 35132 4061 35133
rect 4003 35092 4012 35132
rect 4052 35092 4061 35132
rect 4003 35091 4061 35092
rect 11403 35132 11445 35141
rect 11403 35092 11404 35132
rect 11444 35092 11445 35132
rect 11403 35083 11445 35092
rect 15915 35132 15957 35141
rect 15915 35092 15916 35132
rect 15956 35092 15957 35132
rect 15915 35083 15957 35092
rect 16011 35132 16053 35141
rect 16011 35092 16012 35132
rect 16052 35092 16053 35132
rect 16011 35083 16053 35092
rect 18603 35132 18645 35141
rect 18603 35092 18604 35132
rect 18644 35092 18645 35132
rect 18603 35083 18645 35092
rect 1707 35048 1749 35057
rect 1707 35008 1708 35048
rect 1748 35008 1749 35048
rect 1707 34999 1749 35008
rect 3819 35048 3861 35057
rect 3819 35008 3820 35048
rect 3860 35008 3861 35048
rect 3819 34999 3861 35008
rect 8419 35048 8477 35049
rect 8419 35008 8428 35048
rect 8468 35008 8477 35048
rect 8419 35007 8477 35008
rect 17643 35048 17685 35057
rect 17643 35008 17644 35048
rect 17684 35008 17685 35048
rect 17643 34999 17685 35008
rect 1899 34964 1941 34973
rect 1899 34924 1900 34964
rect 1940 34924 1941 34964
rect 1899 34915 1941 34924
rect 9963 34964 10005 34973
rect 9963 34924 9964 34964
rect 10004 34924 10005 34964
rect 9963 34915 10005 34924
rect 10635 34922 10677 34931
rect 10635 34882 10636 34922
rect 10676 34882 10677 34922
rect 10635 34873 10677 34882
rect 1152 34796 20352 34820
rect 1152 34756 3688 34796
rect 3728 34756 3770 34796
rect 3810 34756 3852 34796
rect 3892 34756 3934 34796
rect 3974 34756 4016 34796
rect 4056 34756 18808 34796
rect 18848 34756 18890 34796
rect 18930 34756 18972 34796
rect 19012 34756 19054 34796
rect 19094 34756 19136 34796
rect 19176 34756 20352 34796
rect 1152 34732 20352 34756
rect 1707 34628 1749 34637
rect 1707 34588 1708 34628
rect 1748 34588 1749 34628
rect 1707 34579 1749 34588
rect 1899 34628 1941 34637
rect 1899 34588 1900 34628
rect 1940 34588 1941 34628
rect 1899 34579 1941 34588
rect 9771 34628 9813 34637
rect 9771 34588 9772 34628
rect 9812 34588 9813 34628
rect 9771 34579 9813 34588
rect 10059 34628 10101 34637
rect 10059 34588 10060 34628
rect 10100 34588 10101 34628
rect 10059 34579 10101 34588
rect 16971 34628 17013 34637
rect 16971 34588 16972 34628
rect 17012 34588 17013 34628
rect 16971 34579 17013 34588
rect 19755 34628 19797 34637
rect 19755 34588 19756 34628
rect 19796 34588 19797 34628
rect 19755 34579 19797 34588
rect 9571 34544 9629 34545
rect 9571 34504 9580 34544
rect 9620 34504 9629 34544
rect 9571 34503 9629 34504
rect 17643 34544 17685 34553
rect 17643 34504 17644 34544
rect 17684 34504 17685 34544
rect 17643 34495 17685 34504
rect 1507 34460 1565 34461
rect 1507 34420 1516 34460
rect 1556 34420 1565 34460
rect 1507 34419 1565 34420
rect 2083 34460 2141 34461
rect 2083 34420 2092 34460
rect 2132 34420 2141 34460
rect 2083 34419 2141 34420
rect 17443 34460 17501 34461
rect 17443 34420 17452 34460
rect 17492 34420 17501 34460
rect 17443 34419 17501 34420
rect 19939 34460 19997 34461
rect 19939 34420 19948 34460
rect 19988 34420 19997 34460
rect 19939 34419 19997 34420
rect 3963 34385 4005 34394
rect 15003 34385 15045 34394
rect 2379 34376 2421 34385
rect 2379 34336 2380 34376
rect 2420 34336 2421 34376
rect 2379 34327 2421 34336
rect 2475 34376 2517 34385
rect 2475 34336 2476 34376
rect 2516 34336 2517 34376
rect 2475 34327 2517 34336
rect 2859 34376 2901 34385
rect 2859 34336 2860 34376
rect 2900 34336 2901 34376
rect 2859 34327 2901 34336
rect 2955 34376 2997 34385
rect 2955 34336 2956 34376
rect 2996 34336 2997 34376
rect 2955 34327 2997 34336
rect 3427 34376 3485 34377
rect 3427 34336 3436 34376
rect 3476 34336 3485 34376
rect 3963 34345 3964 34385
rect 4004 34345 4005 34385
rect 3963 34336 4005 34345
rect 4483 34376 4541 34377
rect 4483 34336 4492 34376
rect 4532 34336 4541 34376
rect 3427 34335 3485 34336
rect 4483 34335 4541 34336
rect 5731 34376 5789 34377
rect 5731 34336 5740 34376
rect 5780 34336 5789 34376
rect 5731 34335 5789 34336
rect 6219 34376 6261 34385
rect 6219 34336 6220 34376
rect 6260 34336 6261 34376
rect 6219 34327 6261 34336
rect 6315 34376 6357 34385
rect 6315 34336 6316 34376
rect 6356 34336 6357 34376
rect 6315 34327 6357 34336
rect 6499 34376 6557 34377
rect 6499 34336 6508 34376
rect 6548 34336 6557 34376
rect 6499 34335 6557 34336
rect 7747 34376 7805 34377
rect 7747 34336 7756 34376
rect 7796 34336 7805 34376
rect 7747 34335 7805 34336
rect 8899 34376 8957 34377
rect 8899 34336 8908 34376
rect 8948 34336 8957 34376
rect 8899 34335 8957 34336
rect 9195 34376 9237 34385
rect 9195 34336 9196 34376
rect 9236 34336 9237 34376
rect 9195 34327 9237 34336
rect 9291 34376 9333 34385
rect 9291 34336 9292 34376
rect 9332 34336 9333 34376
rect 10243 34376 10301 34377
rect 9291 34327 9333 34336
rect 9859 34365 9917 34366
rect 9859 34325 9868 34365
rect 9908 34325 9917 34365
rect 10243 34336 10252 34376
rect 10292 34336 10301 34376
rect 10243 34335 10301 34336
rect 11491 34376 11549 34377
rect 11491 34336 11500 34376
rect 11540 34336 11549 34376
rect 11491 34335 11549 34336
rect 11683 34376 11741 34377
rect 11683 34336 11692 34376
rect 11732 34336 11741 34376
rect 11683 34335 11741 34336
rect 12931 34376 12989 34377
rect 12931 34336 12940 34376
rect 12980 34336 12989 34376
rect 12931 34335 12989 34336
rect 13419 34376 13461 34385
rect 13419 34336 13420 34376
rect 13460 34336 13461 34376
rect 13419 34327 13461 34336
rect 13515 34376 13557 34385
rect 13515 34336 13516 34376
rect 13556 34336 13557 34376
rect 13515 34327 13557 34336
rect 13899 34376 13941 34385
rect 13899 34336 13900 34376
rect 13940 34336 13941 34376
rect 13899 34327 13941 34336
rect 13995 34376 14037 34385
rect 13995 34336 13996 34376
rect 14036 34336 14037 34376
rect 13995 34327 14037 34336
rect 14467 34376 14525 34377
rect 14467 34336 14476 34376
rect 14516 34336 14525 34376
rect 15003 34345 15004 34385
rect 15044 34345 15045 34385
rect 15003 34336 15045 34345
rect 15523 34376 15581 34377
rect 15523 34336 15532 34376
rect 15572 34336 15581 34376
rect 14467 34335 14525 34336
rect 15523 34335 15581 34336
rect 16771 34376 16829 34377
rect 16771 34336 16780 34376
rect 16820 34336 16829 34376
rect 16771 34335 16829 34336
rect 17835 34376 17877 34385
rect 17835 34336 17836 34376
rect 17876 34336 17877 34376
rect 17835 34327 17877 34336
rect 18027 34376 18069 34385
rect 18027 34336 18028 34376
rect 18068 34336 18069 34376
rect 18027 34327 18069 34336
rect 18123 34376 18165 34385
rect 18123 34336 18124 34376
rect 18164 34336 18165 34376
rect 18123 34327 18165 34336
rect 18307 34376 18365 34377
rect 18307 34336 18316 34376
rect 18356 34336 18365 34376
rect 18307 34335 18365 34336
rect 19555 34376 19613 34377
rect 19555 34336 19564 34376
rect 19604 34336 19613 34376
rect 19555 34335 19613 34336
rect 9859 34324 9917 34325
rect 7947 34292 7989 34301
rect 7947 34252 7948 34292
rect 7988 34252 7989 34292
rect 7947 34243 7989 34252
rect 13131 34292 13173 34301
rect 13131 34252 13132 34292
rect 13172 34252 13173 34292
rect 13131 34243 13173 34252
rect 4107 34208 4149 34217
rect 4107 34168 4108 34208
rect 4148 34168 4149 34208
rect 4107 34159 4149 34168
rect 4299 34208 4341 34217
rect 4299 34168 4300 34208
rect 4340 34168 4341 34208
rect 4299 34159 4341 34168
rect 6019 34208 6077 34209
rect 6019 34168 6028 34208
rect 6068 34168 6077 34208
rect 6019 34167 6077 34168
rect 8523 34208 8565 34217
rect 8523 34168 8524 34208
rect 8564 34168 8565 34208
rect 8523 34159 8565 34168
rect 15147 34208 15189 34217
rect 15147 34168 15148 34208
rect 15188 34168 15189 34208
rect 15147 34159 15189 34168
rect 20139 34208 20181 34217
rect 20139 34168 20140 34208
rect 20180 34168 20181 34208
rect 20139 34159 20181 34168
rect 1152 34040 20452 34064
rect 1152 34000 4928 34040
rect 4968 34000 5010 34040
rect 5050 34000 5092 34040
rect 5132 34000 5174 34040
rect 5214 34000 5256 34040
rect 5296 34000 20048 34040
rect 20088 34000 20130 34040
rect 20170 34000 20212 34040
rect 20252 34000 20294 34040
rect 20334 34000 20376 34040
rect 20416 34000 20452 34040
rect 1152 33976 20452 34000
rect 13419 33914 13461 33923
rect 5739 33872 5781 33881
rect 5739 33832 5740 33872
rect 5780 33832 5781 33872
rect 13419 33874 13420 33914
rect 13460 33874 13461 33914
rect 13419 33865 13461 33874
rect 15051 33872 15093 33881
rect 5739 33823 5781 33832
rect 15051 33832 15052 33872
rect 15092 33832 15093 33872
rect 15051 33823 15093 33832
rect 11403 33788 11445 33797
rect 11403 33748 11404 33788
rect 11444 33748 11445 33788
rect 11403 33739 11445 33748
rect 16875 33788 16917 33797
rect 16875 33748 16876 33788
rect 16916 33748 16917 33788
rect 16875 33739 16917 33748
rect 1219 33704 1277 33705
rect 1219 33664 1228 33704
rect 1268 33664 1277 33704
rect 1219 33663 1277 33664
rect 2467 33704 2525 33705
rect 2467 33664 2476 33704
rect 2516 33664 2525 33704
rect 2467 33663 2525 33664
rect 3819 33704 3861 33713
rect 3819 33664 3820 33704
rect 3860 33664 3861 33704
rect 3819 33655 3861 33664
rect 4011 33704 4053 33713
rect 4011 33664 4012 33704
rect 4052 33664 4053 33704
rect 4011 33655 4053 33664
rect 4107 33704 4149 33713
rect 4107 33664 4108 33704
rect 4148 33664 4149 33704
rect 4107 33655 4149 33664
rect 4291 33704 4349 33705
rect 4291 33664 4300 33704
rect 4340 33664 4349 33704
rect 4291 33663 4349 33664
rect 5539 33704 5597 33705
rect 5539 33664 5548 33704
rect 5588 33664 5597 33704
rect 5539 33663 5597 33664
rect 5923 33704 5981 33705
rect 5923 33664 5932 33704
rect 5972 33664 5981 33704
rect 5923 33663 5981 33664
rect 7171 33704 7229 33705
rect 7171 33664 7180 33704
rect 7220 33664 7229 33704
rect 7843 33704 7901 33705
rect 7171 33663 7229 33664
rect 7651 33691 7709 33692
rect 7651 33651 7660 33691
rect 7700 33651 7709 33691
rect 7843 33664 7852 33704
rect 7892 33664 7901 33704
rect 7843 33663 7901 33664
rect 8235 33704 8277 33713
rect 8235 33664 8236 33704
rect 8276 33664 8277 33704
rect 8235 33655 8277 33664
rect 8515 33704 8573 33705
rect 8515 33664 8524 33704
rect 8564 33664 8573 33704
rect 8515 33663 8573 33664
rect 8811 33704 8853 33713
rect 8811 33664 8812 33704
rect 8852 33664 8853 33704
rect 8811 33655 8853 33664
rect 8907 33704 8949 33713
rect 8907 33664 8908 33704
rect 8948 33664 8949 33704
rect 8907 33655 8949 33664
rect 9387 33704 9429 33713
rect 9387 33664 9388 33704
rect 9428 33664 9429 33704
rect 9387 33655 9429 33664
rect 9763 33704 9821 33705
rect 9763 33664 9772 33704
rect 9812 33664 9821 33704
rect 9763 33663 9821 33664
rect 9955 33704 10013 33705
rect 9955 33664 9964 33704
rect 10004 33664 10013 33704
rect 9955 33663 10013 33664
rect 11203 33704 11261 33705
rect 11203 33664 11212 33704
rect 11252 33664 11261 33704
rect 11203 33663 11261 33664
rect 11691 33704 11733 33713
rect 11691 33664 11692 33704
rect 11732 33664 11733 33704
rect 11691 33655 11733 33664
rect 11787 33704 11829 33713
rect 11787 33664 11788 33704
rect 11828 33664 11829 33704
rect 11787 33655 11829 33664
rect 12739 33704 12797 33705
rect 12739 33664 12748 33704
rect 12788 33664 12797 33704
rect 13603 33704 13661 33705
rect 12739 33663 12797 33664
rect 13227 33690 13269 33699
rect 7651 33650 7709 33651
rect 13227 33650 13228 33690
rect 13268 33650 13269 33690
rect 13603 33664 13612 33704
rect 13652 33664 13661 33704
rect 13603 33663 13661 33664
rect 14851 33704 14909 33705
rect 14851 33664 14860 33704
rect 14900 33664 14909 33704
rect 14851 33663 14909 33664
rect 15427 33704 15485 33705
rect 15427 33664 15436 33704
rect 15476 33664 15485 33704
rect 15427 33663 15485 33664
rect 16675 33704 16733 33705
rect 16675 33664 16684 33704
rect 16724 33664 16733 33704
rect 16675 33663 16733 33664
rect 17155 33704 17213 33705
rect 17155 33664 17164 33704
rect 17204 33664 17213 33704
rect 17155 33663 17213 33664
rect 17451 33704 17493 33713
rect 17451 33664 17452 33704
rect 17492 33664 17493 33704
rect 17451 33655 17493 33664
rect 17547 33704 17589 33713
rect 17547 33664 17548 33704
rect 17588 33664 17589 33704
rect 17547 33655 17589 33664
rect 18307 33704 18365 33705
rect 18307 33664 18316 33704
rect 18356 33664 18365 33704
rect 18307 33663 18365 33664
rect 19555 33704 19613 33705
rect 19555 33664 19564 33704
rect 19604 33664 19613 33704
rect 19555 33663 19613 33664
rect 13227 33641 13269 33650
rect 7947 33620 7989 33629
rect 7947 33580 7948 33620
rect 7988 33580 7989 33620
rect 7947 33571 7989 33580
rect 8139 33620 8181 33629
rect 8139 33580 8140 33620
rect 8180 33580 8181 33620
rect 8139 33571 8181 33580
rect 9483 33620 9525 33629
rect 9483 33580 9484 33620
rect 9524 33580 9525 33620
rect 9483 33571 9525 33580
rect 9675 33620 9717 33629
rect 9675 33580 9676 33620
rect 9716 33580 9717 33620
rect 9675 33571 9717 33580
rect 12171 33620 12213 33629
rect 12171 33580 12172 33620
rect 12212 33580 12213 33620
rect 12171 33571 12213 33580
rect 12267 33620 12309 33629
rect 12267 33580 12268 33620
rect 12308 33580 12309 33620
rect 12267 33571 12309 33580
rect 19939 33620 19997 33621
rect 19939 33580 19948 33620
rect 19988 33580 19997 33620
rect 19939 33579 19997 33580
rect 4099 33536 4157 33537
rect 4099 33496 4108 33536
rect 4148 33496 4157 33536
rect 4099 33495 4157 33496
rect 8043 33536 8085 33545
rect 8043 33496 8044 33536
rect 8084 33496 8085 33536
rect 8043 33487 8085 33496
rect 9579 33536 9621 33545
rect 9579 33496 9580 33536
rect 9620 33496 9621 33536
rect 9579 33487 9621 33496
rect 2667 33452 2709 33461
rect 2667 33412 2668 33452
rect 2708 33412 2709 33452
rect 2667 33403 2709 33412
rect 5739 33452 5781 33461
rect 5739 33412 5740 33452
rect 5780 33412 5781 33452
rect 5739 33403 5781 33412
rect 7371 33452 7413 33461
rect 7371 33412 7372 33452
rect 7412 33412 7413 33452
rect 7371 33403 7413 33412
rect 7563 33452 7605 33461
rect 7563 33412 7564 33452
rect 7604 33412 7605 33452
rect 7563 33403 7605 33412
rect 9187 33452 9245 33453
rect 9187 33412 9196 33452
rect 9236 33412 9245 33452
rect 9187 33411 9245 33412
rect 17827 33452 17885 33453
rect 17827 33412 17836 33452
rect 17876 33412 17885 33452
rect 17827 33411 17885 33412
rect 19755 33452 19797 33461
rect 19755 33412 19756 33452
rect 19796 33412 19797 33452
rect 19755 33403 19797 33412
rect 20139 33452 20181 33461
rect 20139 33412 20140 33452
rect 20180 33412 20181 33452
rect 20139 33403 20181 33412
rect 1152 33284 20352 33308
rect 1152 33244 3688 33284
rect 3728 33244 3770 33284
rect 3810 33244 3852 33284
rect 3892 33244 3934 33284
rect 3974 33244 4016 33284
rect 4056 33244 18808 33284
rect 18848 33244 18890 33284
rect 18930 33244 18972 33284
rect 19012 33244 19054 33284
rect 19094 33244 19136 33284
rect 19176 33244 20352 33284
rect 1152 33220 20352 33244
rect 5835 33116 5877 33125
rect 5835 33076 5836 33116
rect 5876 33076 5877 33116
rect 5835 33067 5877 33076
rect 9291 33116 9333 33125
rect 9291 33076 9292 33116
rect 9332 33076 9333 33116
rect 9291 33067 9333 33076
rect 13323 33116 13365 33125
rect 13323 33076 13324 33116
rect 13364 33076 13365 33116
rect 13323 33067 13365 33076
rect 9483 33032 9525 33041
rect 9483 32992 9484 33032
rect 9524 32992 9525 33032
rect 9483 32983 9525 32992
rect 3147 32948 3189 32957
rect 3147 32908 3148 32948
rect 3188 32908 3189 32948
rect 3147 32899 3189 32908
rect 2139 32873 2181 32882
rect 2139 32833 2140 32873
rect 2180 32833 2181 32873
rect 2139 32824 2181 32833
rect 2659 32864 2717 32865
rect 2659 32824 2668 32864
rect 2708 32824 2717 32864
rect 2659 32823 2717 32824
rect 3243 32864 3285 32873
rect 3243 32824 3244 32864
rect 3284 32824 3285 32864
rect 3243 32815 3285 32824
rect 3627 32864 3669 32873
rect 3627 32824 3628 32864
rect 3668 32824 3669 32864
rect 3627 32815 3669 32824
rect 3723 32864 3765 32873
rect 3723 32824 3724 32864
rect 3764 32824 3765 32864
rect 3723 32815 3765 32824
rect 4387 32864 4445 32865
rect 4387 32824 4396 32864
rect 4436 32824 4445 32864
rect 4387 32823 4445 32824
rect 5635 32864 5693 32865
rect 5635 32824 5644 32864
rect 5684 32824 5693 32864
rect 5635 32823 5693 32824
rect 6115 32864 6173 32865
rect 6115 32824 6124 32864
rect 6164 32824 6173 32864
rect 6115 32823 6173 32824
rect 6211 32864 6269 32865
rect 6211 32824 6220 32864
rect 6260 32824 6269 32864
rect 6211 32823 6269 32824
rect 6411 32864 6453 32873
rect 6411 32824 6412 32864
rect 6452 32824 6453 32864
rect 6411 32815 6453 32824
rect 6507 32864 6549 32873
rect 6507 32824 6508 32864
rect 6548 32824 6549 32864
rect 6507 32815 6549 32824
rect 6600 32864 6658 32865
rect 6600 32824 6609 32864
rect 6649 32824 6658 32864
rect 6600 32823 6658 32824
rect 6979 32864 7037 32865
rect 6979 32824 6988 32864
rect 7028 32824 7037 32864
rect 6979 32823 7037 32824
rect 8227 32864 8285 32865
rect 8227 32824 8236 32864
rect 8276 32824 8285 32864
rect 8227 32823 8285 32824
rect 8707 32864 8765 32865
rect 8707 32824 8716 32864
rect 8756 32824 8765 32864
rect 8707 32823 8765 32824
rect 8811 32864 8853 32873
rect 8811 32824 8812 32864
rect 8852 32824 8853 32864
rect 8811 32815 8853 32824
rect 8995 32864 9053 32865
rect 8995 32824 9004 32864
rect 9044 32824 9053 32864
rect 8995 32823 9053 32824
rect 9099 32864 9141 32873
rect 9099 32824 9100 32864
rect 9140 32824 9141 32864
rect 9099 32815 9141 32824
rect 9291 32864 9333 32873
rect 9291 32824 9292 32864
rect 9332 32824 9333 32864
rect 9291 32815 9333 32824
rect 9483 32864 9525 32873
rect 9483 32824 9484 32864
rect 9524 32824 9525 32864
rect 9483 32815 9525 32824
rect 9675 32864 9717 32873
rect 9675 32824 9676 32864
rect 9716 32824 9717 32864
rect 9675 32815 9717 32824
rect 9763 32864 9821 32865
rect 9763 32824 9772 32864
rect 9812 32824 9821 32864
rect 9763 32823 9821 32824
rect 9963 32864 10005 32873
rect 9963 32824 9964 32864
rect 10004 32824 10005 32864
rect 9963 32815 10005 32824
rect 10147 32864 10205 32865
rect 10147 32824 10156 32864
rect 10196 32824 10205 32864
rect 10147 32823 10205 32824
rect 11875 32864 11933 32865
rect 11875 32824 11884 32864
rect 11924 32824 11933 32864
rect 11875 32823 11933 32824
rect 13123 32864 13181 32865
rect 13123 32824 13132 32864
rect 13172 32824 13181 32864
rect 13123 32823 13181 32824
rect 14083 32864 14141 32865
rect 14083 32824 14092 32864
rect 14132 32824 14141 32864
rect 14083 32823 14141 32824
rect 15331 32864 15389 32865
rect 15331 32824 15340 32864
rect 15380 32824 15389 32864
rect 15331 32823 15389 32824
rect 15819 32864 15861 32873
rect 15819 32824 15820 32864
rect 15860 32824 15861 32864
rect 15819 32815 15861 32824
rect 15915 32864 15957 32873
rect 15915 32824 15916 32864
rect 15956 32824 15957 32864
rect 15915 32815 15957 32824
rect 16299 32864 16341 32873
rect 16299 32824 16300 32864
rect 16340 32824 16341 32864
rect 16299 32815 16341 32824
rect 16395 32864 16437 32873
rect 17355 32869 17397 32878
rect 16395 32824 16396 32864
rect 16436 32824 16437 32864
rect 16395 32815 16437 32824
rect 16867 32864 16925 32865
rect 16867 32824 16876 32864
rect 16916 32824 16925 32864
rect 16867 32823 16925 32824
rect 17355 32829 17356 32869
rect 17396 32829 17397 32869
rect 17355 32820 17397 32829
rect 17923 32864 17981 32865
rect 17923 32824 17932 32864
rect 17972 32824 17981 32864
rect 17923 32823 17981 32824
rect 19171 32864 19229 32865
rect 19171 32824 19180 32864
rect 19220 32824 19229 32864
rect 19171 32823 19229 32824
rect 19459 32864 19517 32865
rect 19459 32824 19468 32864
rect 19508 32824 19517 32864
rect 19459 32823 19517 32824
rect 19755 32864 19797 32873
rect 19755 32824 19756 32864
rect 19796 32824 19797 32864
rect 19755 32815 19797 32824
rect 19851 32864 19893 32873
rect 19851 32824 19852 32864
rect 19892 32824 19893 32864
rect 19851 32815 19893 32824
rect 10059 32780 10101 32789
rect 10059 32740 10060 32780
rect 10100 32740 10101 32780
rect 10059 32731 10101 32740
rect 15531 32780 15573 32789
rect 15531 32740 15532 32780
rect 15572 32740 15573 32780
rect 15531 32731 15573 32740
rect 17739 32780 17781 32789
rect 17739 32740 17740 32780
rect 17780 32740 17781 32780
rect 17739 32731 17781 32740
rect 1995 32696 2037 32705
rect 1995 32656 1996 32696
rect 2036 32656 2037 32696
rect 1995 32647 2037 32656
rect 6595 32696 6653 32697
rect 6595 32656 6604 32696
rect 6644 32656 6653 32696
rect 6595 32655 6653 32656
rect 8427 32696 8469 32705
rect 8427 32656 8428 32696
rect 8468 32656 8469 32696
rect 8427 32647 8469 32656
rect 17547 32696 17589 32705
rect 17547 32656 17548 32696
rect 17588 32656 17589 32696
rect 17547 32647 17589 32656
rect 20139 32654 20181 32663
rect 20139 32614 20140 32654
rect 20180 32614 20181 32654
rect 20139 32605 20181 32614
rect 1152 32528 20452 32552
rect 1152 32488 4928 32528
rect 4968 32488 5010 32528
rect 5050 32488 5092 32528
rect 5132 32488 5174 32528
rect 5214 32488 5256 32528
rect 5296 32488 20048 32528
rect 20088 32488 20130 32528
rect 20170 32488 20212 32528
rect 20252 32488 20294 32528
rect 20334 32488 20376 32528
rect 20416 32488 20452 32528
rect 1152 32464 20452 32488
rect 6115 32360 6173 32361
rect 6115 32320 6124 32360
rect 6164 32320 6173 32360
rect 6115 32319 6173 32320
rect 8227 32360 8285 32361
rect 8227 32320 8236 32360
rect 8276 32320 8285 32360
rect 8227 32319 8285 32320
rect 17643 32360 17685 32369
rect 17643 32320 17644 32360
rect 17684 32320 17685 32360
rect 17643 32311 17685 32320
rect 2083 32192 2141 32193
rect 2083 32152 2092 32192
rect 2132 32152 2141 32192
rect 2083 32151 2141 32152
rect 3331 32192 3389 32193
rect 3331 32152 3340 32192
rect 3380 32152 3389 32192
rect 3331 32151 3389 32152
rect 4195 32192 4253 32193
rect 4195 32152 4204 32192
rect 4244 32152 4253 32192
rect 4195 32151 4253 32152
rect 5443 32192 5501 32193
rect 5443 32152 5452 32192
rect 5492 32152 5501 32192
rect 5443 32151 5501 32152
rect 5835 32192 5877 32201
rect 5835 32152 5836 32192
rect 5876 32152 5877 32192
rect 5835 32143 5877 32152
rect 5931 32192 5973 32201
rect 5931 32152 5932 32192
rect 5972 32152 5973 32192
rect 5931 32143 5973 32152
rect 6307 32192 6365 32193
rect 6307 32152 6316 32192
rect 6356 32152 6365 32192
rect 6307 32151 6365 32152
rect 7555 32192 7613 32193
rect 7555 32152 7564 32192
rect 7604 32152 7613 32192
rect 7555 32151 7613 32152
rect 7947 32192 7989 32201
rect 7947 32152 7948 32192
rect 7988 32152 7989 32192
rect 7947 32143 7989 32152
rect 8043 32192 8085 32201
rect 8043 32152 8044 32192
rect 8084 32152 8085 32192
rect 8043 32143 8085 32152
rect 8707 32192 8765 32193
rect 8707 32152 8716 32192
rect 8756 32152 8765 32192
rect 8707 32151 8765 32152
rect 9955 32192 10013 32193
rect 9955 32152 9964 32192
rect 10004 32152 10013 32192
rect 9955 32151 10013 32152
rect 12931 32192 12989 32193
rect 12931 32152 12940 32192
rect 12980 32152 12989 32192
rect 12931 32151 12989 32152
rect 14179 32192 14237 32193
rect 14179 32152 14188 32192
rect 14228 32152 14237 32192
rect 14179 32151 14237 32152
rect 14563 32192 14621 32193
rect 14563 32152 14572 32192
rect 14612 32152 14621 32192
rect 14563 32151 14621 32152
rect 15915 32192 15957 32201
rect 15915 32152 15916 32192
rect 15956 32152 15957 32192
rect 15915 32143 15957 32152
rect 16011 32192 16053 32201
rect 16011 32152 16012 32192
rect 16052 32152 16053 32192
rect 16011 32143 16053 32152
rect 16963 32192 17021 32193
rect 16963 32152 16972 32192
rect 17012 32152 17021 32192
rect 16963 32151 17021 32152
rect 17451 32187 17493 32196
rect 17451 32147 17452 32187
rect 17492 32147 17493 32187
rect 18115 32192 18173 32193
rect 18115 32152 18124 32192
rect 18164 32152 18173 32192
rect 18115 32151 18173 32152
rect 19075 32192 19133 32193
rect 19075 32152 19084 32192
rect 19124 32152 19133 32192
rect 19075 32151 19133 32152
rect 17451 32138 17493 32147
rect 16395 32108 16437 32117
rect 16395 32068 16396 32108
rect 16436 32068 16437 32108
rect 16395 32059 16437 32068
rect 16491 32108 16533 32117
rect 16491 32068 16492 32108
rect 16532 32068 16533 32108
rect 16491 32059 16533 32068
rect 19267 32108 19325 32109
rect 19267 32068 19276 32108
rect 19316 32068 19325 32108
rect 20035 32108 20093 32109
rect 19267 32067 19325 32068
rect 19651 32097 19709 32098
rect 19651 32057 19660 32097
rect 19700 32057 19709 32097
rect 20035 32068 20044 32108
rect 20084 32068 20093 32108
rect 20035 32067 20093 32068
rect 19651 32056 19709 32057
rect 19467 32024 19509 32033
rect 19467 31984 19468 32024
rect 19508 31984 19509 32024
rect 19467 31975 19509 31984
rect 19851 32024 19893 32033
rect 19851 31984 19852 32024
rect 19892 31984 19893 32024
rect 19851 31975 19893 31984
rect 3531 31940 3573 31949
rect 3531 31900 3532 31940
rect 3572 31900 3573 31940
rect 3531 31891 3573 31900
rect 5643 31940 5685 31949
rect 5643 31900 5644 31940
rect 5684 31900 5685 31940
rect 5643 31891 5685 31900
rect 7755 31940 7797 31949
rect 7755 31900 7756 31940
rect 7796 31900 7797 31940
rect 7755 31891 7797 31900
rect 10155 31940 10197 31949
rect 10155 31900 10156 31940
rect 10196 31900 10197 31940
rect 10155 31891 10197 31900
rect 14379 31940 14421 31949
rect 14379 31900 14380 31940
rect 14420 31900 14421 31940
rect 14379 31891 14421 31900
rect 14667 31940 14709 31949
rect 14667 31900 14668 31940
rect 14708 31900 14709 31940
rect 14667 31891 14709 31900
rect 20235 31940 20277 31949
rect 20235 31900 20236 31940
rect 20276 31900 20277 31940
rect 20235 31891 20277 31900
rect 1152 31772 20352 31796
rect 1152 31732 3688 31772
rect 3728 31732 3770 31772
rect 3810 31732 3852 31772
rect 3892 31732 3934 31772
rect 3974 31732 4016 31772
rect 4056 31732 18808 31772
rect 18848 31732 18890 31772
rect 18930 31732 18972 31772
rect 19012 31732 19054 31772
rect 19094 31732 19136 31772
rect 19176 31732 20352 31772
rect 1152 31708 20352 31732
rect 17163 31604 17205 31613
rect 17163 31564 17164 31604
rect 17204 31564 17205 31604
rect 17163 31555 17205 31564
rect 14187 31520 14229 31529
rect 14187 31480 14188 31520
rect 14228 31480 14229 31520
rect 14187 31471 14229 31480
rect 6507 31436 6549 31445
rect 6507 31396 6508 31436
rect 6548 31396 6549 31436
rect 8907 31436 8949 31445
rect 6507 31387 6549 31396
rect 6603 31394 6645 31403
rect 2659 31352 2717 31353
rect 2659 31312 2668 31352
rect 2708 31312 2717 31352
rect 2659 31311 2717 31312
rect 3907 31352 3965 31353
rect 3907 31312 3916 31352
rect 3956 31312 3965 31352
rect 3907 31311 3965 31312
rect 4291 31352 4349 31353
rect 4291 31312 4300 31352
rect 4340 31312 4349 31352
rect 4291 31311 4349 31312
rect 5539 31352 5597 31353
rect 5539 31312 5548 31352
rect 5588 31312 5597 31352
rect 5539 31311 5597 31312
rect 6027 31352 6069 31361
rect 6027 31312 6028 31352
rect 6068 31312 6069 31352
rect 6027 31303 6069 31312
rect 6123 31352 6165 31361
rect 6123 31312 6124 31352
rect 6164 31312 6165 31352
rect 6603 31354 6604 31394
rect 6644 31354 6645 31394
rect 8907 31396 8908 31436
rect 8948 31396 8949 31436
rect 10923 31436 10965 31445
rect 8907 31387 8949 31396
rect 9915 31394 9957 31403
rect 6603 31345 6645 31354
rect 7563 31357 7605 31366
rect 7075 31352 7133 31353
rect 6123 31303 6165 31312
rect 7075 31312 7084 31352
rect 7124 31312 7133 31352
rect 7075 31311 7133 31312
rect 7563 31317 7564 31357
rect 7604 31317 7605 31357
rect 7563 31308 7605 31317
rect 8331 31352 8373 31361
rect 8331 31312 8332 31352
rect 8372 31312 8373 31352
rect 8331 31303 8373 31312
rect 8427 31352 8469 31361
rect 8427 31312 8428 31352
rect 8468 31312 8469 31352
rect 8427 31303 8469 31312
rect 8811 31352 8853 31361
rect 9915 31354 9916 31394
rect 9956 31354 9957 31394
rect 10923 31396 10924 31436
rect 10964 31396 10965 31436
rect 10923 31387 10965 31396
rect 11019 31436 11061 31445
rect 11019 31396 11020 31436
rect 11060 31396 11061 31436
rect 11019 31387 11061 31396
rect 17635 31436 17693 31437
rect 17635 31396 17644 31436
rect 17684 31396 17693 31436
rect 17635 31395 17693 31396
rect 19651 31436 19709 31437
rect 19651 31396 19660 31436
rect 19700 31396 19709 31436
rect 19651 31395 19709 31396
rect 20035 31436 20093 31437
rect 20035 31396 20044 31436
rect 20084 31396 20093 31436
rect 20035 31395 20093 31396
rect 12027 31361 12069 31370
rect 8811 31312 8812 31352
rect 8852 31312 8853 31352
rect 8811 31303 8853 31312
rect 9379 31352 9437 31353
rect 9379 31312 9388 31352
rect 9428 31312 9437 31352
rect 9915 31345 9957 31354
rect 10443 31352 10485 31361
rect 9379 31311 9437 31312
rect 10443 31312 10444 31352
rect 10484 31312 10485 31352
rect 10443 31303 10485 31312
rect 10539 31352 10581 31361
rect 10539 31312 10540 31352
rect 10580 31312 10581 31352
rect 10539 31303 10581 31312
rect 11491 31352 11549 31353
rect 11491 31312 11500 31352
rect 11540 31312 11549 31352
rect 12027 31321 12028 31361
rect 12068 31321 12069 31361
rect 12027 31312 12069 31321
rect 12739 31352 12797 31353
rect 12739 31312 12748 31352
rect 12788 31312 12797 31352
rect 11491 31311 11549 31312
rect 12739 31311 12797 31312
rect 13987 31352 14045 31353
rect 13987 31312 13996 31352
rect 14036 31312 14045 31352
rect 13987 31311 14045 31312
rect 14371 31352 14429 31353
rect 14371 31312 14380 31352
rect 14420 31312 14429 31352
rect 14371 31311 14429 31312
rect 14467 31352 14525 31353
rect 14467 31312 14476 31352
rect 14516 31312 14525 31352
rect 14467 31311 14525 31312
rect 14667 31352 14709 31361
rect 14667 31312 14668 31352
rect 14708 31312 14709 31352
rect 14667 31303 14709 31312
rect 14763 31352 14805 31361
rect 14763 31312 14764 31352
rect 14804 31312 14805 31352
rect 14763 31303 14805 31312
rect 14856 31352 14914 31353
rect 14856 31312 14865 31352
rect 14905 31312 14914 31352
rect 14856 31311 14914 31312
rect 15147 31352 15189 31361
rect 15147 31312 15148 31352
rect 15188 31312 15189 31352
rect 15147 31303 15189 31312
rect 15243 31352 15285 31361
rect 15243 31312 15244 31352
rect 15284 31312 15285 31352
rect 15243 31303 15285 31312
rect 17163 31352 17205 31361
rect 17163 31312 17164 31352
rect 17204 31312 17205 31352
rect 17163 31303 17205 31312
rect 17355 31352 17397 31361
rect 17355 31312 17356 31352
rect 17396 31312 17397 31352
rect 17355 31303 17397 31312
rect 17443 31352 17501 31353
rect 17443 31312 17452 31352
rect 17492 31312 17501 31352
rect 17443 31311 17501 31312
rect 18123 31352 18165 31361
rect 18123 31312 18124 31352
rect 18164 31312 18165 31352
rect 18123 31303 18165 31312
rect 18219 31352 18261 31361
rect 18219 31312 18220 31352
rect 18260 31312 18261 31352
rect 18219 31303 18261 31312
rect 18315 31352 18357 31361
rect 18315 31312 18316 31352
rect 18356 31312 18357 31352
rect 18315 31303 18357 31312
rect 18699 31352 18741 31361
rect 18699 31312 18700 31352
rect 18740 31312 18741 31352
rect 18699 31303 18741 31312
rect 18795 31352 18837 31361
rect 18795 31312 18796 31352
rect 18836 31312 18837 31352
rect 18795 31303 18837 31312
rect 18891 31352 18933 31361
rect 18891 31312 18892 31352
rect 18932 31312 18933 31352
rect 18891 31303 18933 31312
rect 19179 31352 19221 31361
rect 19179 31312 19180 31352
rect 19220 31312 19221 31352
rect 19179 31303 19221 31312
rect 19275 31352 19317 31361
rect 19275 31312 19276 31352
rect 19316 31312 19317 31352
rect 19275 31303 19317 31312
rect 19371 31352 19413 31361
rect 19371 31312 19372 31352
rect 19412 31312 19413 31352
rect 19371 31303 19413 31312
rect 4107 31184 4149 31193
rect 4107 31144 4108 31184
rect 4148 31144 4149 31184
rect 4107 31135 4149 31144
rect 5739 31184 5781 31193
rect 5739 31144 5740 31184
rect 5780 31144 5781 31184
rect 5739 31135 5781 31144
rect 7755 31184 7797 31193
rect 7755 31144 7756 31184
rect 7796 31144 7797 31184
rect 7755 31135 7797 31144
rect 10059 31184 10101 31193
rect 10059 31144 10060 31184
rect 10100 31144 10101 31184
rect 10059 31135 10101 31144
rect 12171 31184 12213 31193
rect 12171 31144 12172 31184
rect 12212 31144 12213 31184
rect 12171 31135 12213 31144
rect 14851 31184 14909 31185
rect 14851 31144 14860 31184
rect 14900 31144 14909 31184
rect 14851 31143 14909 31144
rect 15427 31184 15485 31185
rect 15427 31144 15436 31184
rect 15476 31144 15485 31184
rect 15427 31143 15485 31144
rect 17835 31184 17877 31193
rect 17835 31144 17836 31184
rect 17876 31144 17877 31184
rect 17835 31135 17877 31144
rect 18507 31184 18549 31193
rect 18507 31144 18508 31184
rect 18548 31144 18549 31184
rect 18507 31135 18549 31144
rect 18979 31184 19037 31185
rect 18979 31144 18988 31184
rect 19028 31144 19037 31184
rect 18979 31143 19037 31144
rect 19459 31184 19517 31185
rect 19459 31144 19468 31184
rect 19508 31144 19517 31184
rect 19459 31143 19517 31144
rect 19851 31184 19893 31193
rect 19851 31144 19852 31184
rect 19892 31144 19893 31184
rect 19851 31135 19893 31144
rect 20235 31184 20277 31193
rect 20235 31144 20236 31184
rect 20276 31144 20277 31184
rect 20235 31135 20277 31144
rect 1152 31016 20452 31040
rect 1152 30976 4928 31016
rect 4968 30976 5010 31016
rect 5050 30976 5092 31016
rect 5132 30976 5174 31016
rect 5214 30976 5256 31016
rect 5296 30976 20048 31016
rect 20088 30976 20130 31016
rect 20170 30976 20212 31016
rect 20252 30976 20294 31016
rect 20334 30976 20376 31016
rect 20416 30976 20452 31016
rect 1152 30952 20452 30976
rect 4011 30848 4053 30857
rect 4011 30808 4012 30848
rect 4052 30808 4053 30848
rect 4011 30799 4053 30808
rect 6507 30848 6549 30857
rect 6507 30808 6508 30848
rect 6548 30808 6549 30848
rect 6507 30799 6549 30808
rect 8803 30848 8861 30849
rect 8803 30808 8812 30848
rect 8852 30808 8861 30848
rect 8803 30807 8861 30808
rect 10443 30848 10485 30857
rect 10443 30808 10444 30848
rect 10484 30808 10485 30848
rect 10443 30799 10485 30808
rect 12267 30848 12309 30857
rect 12267 30808 12268 30848
rect 12308 30808 12309 30848
rect 12267 30799 12309 30808
rect 16491 30848 16533 30857
rect 16491 30808 16492 30848
rect 16532 30808 16533 30848
rect 16491 30799 16533 30808
rect 18603 30764 18645 30773
rect 18603 30724 18604 30764
rect 18644 30724 18645 30764
rect 18603 30715 18645 30724
rect 2283 30680 2325 30689
rect 2283 30640 2284 30680
rect 2324 30640 2325 30680
rect 2283 30631 2325 30640
rect 2379 30680 2421 30689
rect 2379 30640 2380 30680
rect 2420 30640 2421 30680
rect 2379 30631 2421 30640
rect 3331 30680 3389 30681
rect 3331 30640 3340 30680
rect 3380 30640 3389 30680
rect 3331 30639 3389 30640
rect 3819 30675 3861 30684
rect 3819 30635 3820 30675
rect 3860 30635 3861 30675
rect 3819 30626 3861 30635
rect 4779 30680 4821 30689
rect 4779 30640 4780 30680
rect 4820 30640 4821 30680
rect 4779 30631 4821 30640
rect 4875 30680 4917 30689
rect 4875 30640 4876 30680
rect 4916 30640 4917 30680
rect 4875 30631 4917 30640
rect 5355 30680 5397 30689
rect 5355 30640 5356 30680
rect 5396 30640 5397 30680
rect 5355 30631 5397 30640
rect 5827 30680 5885 30681
rect 5827 30640 5836 30680
rect 5876 30640 5885 30680
rect 5827 30639 5885 30640
rect 6315 30675 6357 30684
rect 6315 30635 6316 30675
rect 6356 30635 6357 30675
rect 6315 30626 6357 30635
rect 8523 30680 8565 30689
rect 8523 30640 8524 30680
rect 8564 30640 8565 30680
rect 8523 30631 8565 30640
rect 8619 30680 8661 30689
rect 8619 30640 8620 30680
rect 8660 30640 8661 30680
rect 8619 30631 8661 30640
rect 8995 30680 9053 30681
rect 8995 30640 9004 30680
rect 9044 30640 9053 30680
rect 8995 30639 9053 30640
rect 10243 30680 10301 30681
rect 10243 30640 10252 30680
rect 10292 30640 10301 30680
rect 10243 30639 10301 30640
rect 10819 30680 10877 30681
rect 10819 30640 10828 30680
rect 10868 30640 10877 30680
rect 10819 30639 10877 30640
rect 12067 30680 12125 30681
rect 12067 30640 12076 30680
rect 12116 30640 12125 30680
rect 12067 30639 12125 30640
rect 12451 30680 12509 30681
rect 12451 30640 12460 30680
rect 12500 30640 12509 30680
rect 12451 30639 12509 30640
rect 13995 30680 14037 30689
rect 13995 30640 13996 30680
rect 14036 30640 14037 30680
rect 13995 30631 14037 30640
rect 14187 30680 14229 30689
rect 14187 30640 14188 30680
rect 14228 30640 14229 30680
rect 14187 30631 14229 30640
rect 14283 30680 14325 30689
rect 14283 30640 14284 30680
rect 14324 30640 14325 30680
rect 14283 30631 14325 30640
rect 14467 30680 14525 30681
rect 14467 30640 14476 30680
rect 14516 30640 14525 30680
rect 14467 30639 14525 30640
rect 15715 30680 15773 30681
rect 15715 30640 15724 30680
rect 15764 30640 15773 30680
rect 15715 30639 15773 30640
rect 16299 30680 16341 30689
rect 16299 30640 16300 30680
rect 16340 30640 16341 30680
rect 16299 30631 16341 30640
rect 16587 30680 16629 30689
rect 16587 30640 16588 30680
rect 16628 30640 16629 30680
rect 16587 30631 16629 30640
rect 16875 30680 16917 30689
rect 16875 30640 16876 30680
rect 16916 30640 16917 30680
rect 16875 30631 16917 30640
rect 16971 30680 17013 30689
rect 16971 30640 16972 30680
rect 17012 30640 17013 30680
rect 16971 30631 17013 30640
rect 17923 30680 17981 30681
rect 17923 30640 17932 30680
rect 17972 30640 17981 30680
rect 18787 30680 18845 30681
rect 17923 30639 17981 30640
rect 18411 30666 18453 30675
rect 18411 30626 18412 30666
rect 18452 30626 18453 30666
rect 18787 30640 18796 30680
rect 18836 30640 18845 30680
rect 18787 30639 18845 30640
rect 20035 30680 20093 30681
rect 20035 30640 20044 30680
rect 20084 30640 20093 30680
rect 20035 30639 20093 30640
rect 18411 30617 18453 30626
rect 2763 30596 2805 30605
rect 2763 30556 2764 30596
rect 2804 30556 2805 30596
rect 2763 30547 2805 30556
rect 2859 30596 2901 30605
rect 2859 30556 2860 30596
rect 2900 30556 2901 30596
rect 2859 30547 2901 30556
rect 5259 30596 5301 30605
rect 5259 30556 5260 30596
rect 5300 30556 5301 30596
rect 5259 30547 5301 30556
rect 17355 30596 17397 30605
rect 17355 30556 17356 30596
rect 17396 30556 17397 30596
rect 17355 30547 17397 30556
rect 17451 30596 17493 30605
rect 17451 30556 17452 30596
rect 17492 30556 17493 30596
rect 17451 30547 17493 30556
rect 14275 30512 14333 30513
rect 14275 30472 14284 30512
rect 14324 30472 14333 30512
rect 14275 30471 14333 30472
rect 12555 30428 12597 30437
rect 12555 30388 12556 30428
rect 12596 30388 12597 30428
rect 12555 30379 12597 30388
rect 15915 30428 15957 30437
rect 15915 30388 15916 30428
rect 15956 30388 15957 30428
rect 15915 30379 15957 30388
rect 20235 30428 20277 30437
rect 20235 30388 20236 30428
rect 20276 30388 20277 30428
rect 20235 30379 20277 30388
rect 1152 30260 20352 30284
rect 1152 30220 3688 30260
rect 3728 30220 3770 30260
rect 3810 30220 3852 30260
rect 3892 30220 3934 30260
rect 3974 30220 4016 30260
rect 4056 30220 18808 30260
rect 18848 30220 18890 30260
rect 18930 30220 18972 30260
rect 19012 30220 19054 30260
rect 19094 30220 19136 30260
rect 19176 30220 20352 30260
rect 1152 30196 20352 30220
rect 11883 30092 11925 30101
rect 11883 30052 11884 30092
rect 11924 30052 11925 30092
rect 11883 30043 11925 30052
rect 17163 30092 17205 30101
rect 17163 30052 17164 30092
rect 17204 30052 17205 30092
rect 17163 30043 17205 30052
rect 18891 30092 18933 30101
rect 18891 30052 18892 30092
rect 18932 30052 18933 30092
rect 18891 30043 18933 30052
rect 5931 30008 5973 30017
rect 5931 29968 5932 30008
rect 5972 29968 5973 30008
rect 5931 29959 5973 29968
rect 13515 30008 13557 30017
rect 13515 29968 13516 30008
rect 13556 29968 13557 30008
rect 13515 29959 13557 29968
rect 15339 29854 15381 29863
rect 1315 29840 1373 29841
rect 1315 29800 1324 29840
rect 1364 29800 1373 29840
rect 1315 29799 1373 29800
rect 2563 29840 2621 29841
rect 2563 29800 2572 29840
rect 2612 29800 2621 29840
rect 2563 29799 2621 29800
rect 3523 29840 3581 29841
rect 3523 29800 3532 29840
rect 3572 29800 3581 29840
rect 3523 29799 3581 29800
rect 4771 29840 4829 29841
rect 4771 29800 4780 29840
rect 4820 29800 4829 29840
rect 4771 29799 4829 29800
rect 5443 29840 5501 29841
rect 5443 29800 5452 29840
rect 5492 29800 5501 29840
rect 5443 29799 5501 29800
rect 5547 29840 5589 29849
rect 5547 29800 5548 29840
rect 5588 29800 5589 29840
rect 5547 29791 5589 29800
rect 5739 29840 5781 29849
rect 5739 29800 5740 29840
rect 5780 29800 5781 29840
rect 5739 29791 5781 29800
rect 5931 29840 5973 29849
rect 5931 29800 5932 29840
rect 5972 29800 5973 29840
rect 5931 29791 5973 29800
rect 6219 29840 6261 29849
rect 6219 29800 6220 29840
rect 6260 29800 6261 29840
rect 6219 29791 6261 29800
rect 6691 29840 6749 29841
rect 6691 29800 6700 29840
rect 6740 29800 6749 29840
rect 6691 29799 6749 29800
rect 7939 29840 7997 29841
rect 7939 29800 7948 29840
rect 7988 29800 7997 29840
rect 7939 29799 7997 29800
rect 8323 29840 8381 29841
rect 8323 29800 8332 29840
rect 8372 29800 8381 29840
rect 8323 29799 8381 29800
rect 8707 29840 8765 29841
rect 8707 29800 8716 29840
rect 8756 29800 8765 29840
rect 8707 29799 8765 29800
rect 8811 29840 8853 29849
rect 8811 29800 8812 29840
rect 8852 29800 8853 29840
rect 8811 29791 8853 29800
rect 9003 29840 9045 29849
rect 9003 29800 9004 29840
rect 9044 29800 9045 29840
rect 9003 29791 9045 29800
rect 9195 29840 9237 29849
rect 9195 29800 9196 29840
rect 9236 29800 9237 29840
rect 9195 29791 9237 29800
rect 9387 29840 9429 29849
rect 9387 29800 9388 29840
rect 9428 29800 9429 29840
rect 9387 29791 9429 29800
rect 9475 29840 9533 29841
rect 9475 29800 9484 29840
rect 9524 29800 9533 29840
rect 9475 29799 9533 29800
rect 10059 29840 10101 29849
rect 10059 29800 10060 29840
rect 10100 29800 10101 29840
rect 10059 29791 10101 29800
rect 10251 29840 10293 29849
rect 10251 29800 10252 29840
rect 10292 29800 10293 29840
rect 10251 29791 10293 29800
rect 10435 29840 10493 29841
rect 10435 29800 10444 29840
rect 10484 29800 10493 29840
rect 10435 29799 10493 29800
rect 11683 29840 11741 29841
rect 11683 29800 11692 29840
rect 11732 29800 11741 29840
rect 11683 29799 11741 29800
rect 12067 29840 12125 29841
rect 12067 29800 12076 29840
rect 12116 29800 12125 29840
rect 12067 29799 12125 29800
rect 13315 29840 13373 29841
rect 13315 29800 13324 29840
rect 13364 29800 13373 29840
rect 13315 29799 13373 29800
rect 13803 29840 13845 29849
rect 13803 29800 13804 29840
rect 13844 29800 13845 29840
rect 13803 29791 13845 29800
rect 13899 29840 13941 29849
rect 13899 29800 13900 29840
rect 13940 29800 13941 29840
rect 13899 29791 13941 29800
rect 14283 29840 14325 29849
rect 14283 29800 14284 29840
rect 14324 29800 14325 29840
rect 14283 29791 14325 29800
rect 14379 29840 14421 29849
rect 14379 29800 14380 29840
rect 14420 29800 14421 29840
rect 14379 29791 14421 29800
rect 14851 29840 14909 29841
rect 14851 29800 14860 29840
rect 14900 29800 14909 29840
rect 15339 29814 15340 29854
rect 15380 29814 15381 29854
rect 15339 29805 15381 29814
rect 15715 29840 15773 29841
rect 14851 29799 14909 29800
rect 15715 29800 15724 29840
rect 15764 29800 15773 29840
rect 15715 29799 15773 29800
rect 16963 29840 17021 29841
rect 16963 29800 16972 29840
rect 17012 29800 17021 29840
rect 16963 29799 17021 29800
rect 17443 29840 17501 29841
rect 17443 29800 17452 29840
rect 17492 29800 17501 29840
rect 17443 29799 17501 29800
rect 18691 29840 18749 29841
rect 18691 29800 18700 29840
rect 18740 29800 18749 29840
rect 18691 29799 18749 29800
rect 19275 29840 19317 29849
rect 19275 29800 19276 29840
rect 19316 29800 19317 29840
rect 19275 29791 19317 29800
rect 8139 29756 8181 29765
rect 8139 29716 8140 29756
rect 8180 29716 8181 29756
rect 8139 29707 8181 29716
rect 15531 29756 15573 29765
rect 15531 29716 15532 29756
rect 15572 29716 15573 29756
rect 15531 29707 15573 29716
rect 2763 29672 2805 29681
rect 2763 29632 2764 29672
rect 2804 29632 2805 29672
rect 2763 29623 2805 29632
rect 4971 29672 5013 29681
rect 4971 29632 4972 29672
rect 5012 29632 5013 29672
rect 4971 29623 5013 29632
rect 5635 29672 5693 29673
rect 5635 29632 5644 29672
rect 5684 29632 5693 29672
rect 5635 29631 5693 29632
rect 8427 29672 8469 29681
rect 8427 29632 8428 29672
rect 8468 29632 8469 29672
rect 8427 29623 8469 29632
rect 8899 29672 8957 29673
rect 8899 29632 8908 29672
rect 8948 29632 8957 29672
rect 8899 29631 8957 29632
rect 9283 29672 9341 29673
rect 9283 29632 9292 29672
rect 9332 29632 9341 29672
rect 9283 29631 9341 29632
rect 10155 29672 10197 29681
rect 10155 29632 10156 29672
rect 10196 29632 10197 29672
rect 10155 29623 10197 29632
rect 19659 29672 19701 29681
rect 19659 29632 19660 29672
rect 19700 29632 19701 29672
rect 19659 29623 19701 29632
rect 1152 29504 20452 29528
rect 1152 29464 4928 29504
rect 4968 29464 5010 29504
rect 5050 29464 5092 29504
rect 5132 29464 5174 29504
rect 5214 29464 5256 29504
rect 5296 29464 20048 29504
rect 20088 29464 20130 29504
rect 20170 29464 20212 29504
rect 20252 29464 20294 29504
rect 20334 29464 20376 29504
rect 20416 29464 20452 29504
rect 1152 29440 20452 29464
rect 8331 29340 8373 29349
rect 7651 29336 7709 29337
rect 7651 29296 7660 29336
rect 7700 29296 7709 29336
rect 7651 29295 7709 29296
rect 8331 29300 8332 29340
rect 8372 29300 8373 29340
rect 8331 29291 8373 29300
rect 8803 29336 8861 29337
rect 8803 29296 8812 29336
rect 8852 29296 8861 29336
rect 8803 29295 8861 29296
rect 18027 29336 18069 29345
rect 18027 29296 18028 29336
rect 18068 29296 18069 29336
rect 18027 29287 18069 29296
rect 18307 29336 18365 29337
rect 18307 29296 18316 29336
rect 18356 29296 18365 29336
rect 18307 29295 18365 29296
rect 18891 29336 18933 29345
rect 18891 29296 18892 29336
rect 18932 29296 18933 29336
rect 18891 29287 18933 29296
rect 13707 29252 13749 29261
rect 13707 29212 13708 29252
rect 13748 29212 13749 29252
rect 13707 29203 13749 29212
rect 15723 29252 15765 29261
rect 15723 29212 15724 29252
rect 15764 29212 15765 29252
rect 15723 29203 15765 29212
rect 19563 29252 19605 29261
rect 19563 29212 19564 29252
rect 19604 29212 19605 29252
rect 19563 29203 19605 29212
rect 13995 29188 14037 29197
rect 2083 29168 2141 29169
rect 2083 29128 2092 29168
rect 2132 29128 2141 29168
rect 2083 29127 2141 29128
rect 3331 29168 3389 29169
rect 3331 29128 3340 29168
rect 3380 29128 3389 29168
rect 3331 29127 3389 29128
rect 3907 29168 3965 29169
rect 3907 29128 3916 29168
rect 3956 29128 3965 29168
rect 3907 29127 3965 29128
rect 5155 29168 5213 29169
rect 5155 29128 5164 29168
rect 5204 29128 5213 29168
rect 5155 29127 5213 29128
rect 5643 29168 5685 29177
rect 5643 29128 5644 29168
rect 5684 29128 5685 29168
rect 5643 29119 5685 29128
rect 5739 29168 5781 29177
rect 5739 29128 5740 29168
rect 5780 29128 5781 29168
rect 5739 29119 5781 29128
rect 5835 29168 5877 29177
rect 5835 29128 5836 29168
rect 5876 29128 5877 29168
rect 5835 29119 5877 29128
rect 6219 29168 6261 29177
rect 6219 29128 6220 29168
rect 6260 29128 6261 29168
rect 6219 29119 6261 29128
rect 6315 29168 6357 29177
rect 6315 29128 6316 29168
rect 6356 29128 6357 29168
rect 6315 29119 6357 29128
rect 6411 29168 6453 29177
rect 6411 29128 6412 29168
rect 6452 29128 6453 29168
rect 6411 29119 6453 29128
rect 6507 29168 6549 29177
rect 6507 29128 6508 29168
rect 6548 29128 6549 29168
rect 6507 29119 6549 29128
rect 7371 29168 7413 29177
rect 7371 29128 7372 29168
rect 7412 29128 7413 29168
rect 7371 29119 7413 29128
rect 7467 29168 7509 29177
rect 7467 29128 7468 29168
rect 7508 29128 7509 29168
rect 7467 29119 7509 29128
rect 8139 29168 8181 29177
rect 8139 29128 8140 29168
rect 8180 29128 8181 29168
rect 8139 29119 8181 29128
rect 8227 29168 8285 29169
rect 8227 29128 8236 29168
rect 8276 29128 8285 29168
rect 8227 29127 8285 29128
rect 8515 29168 8573 29169
rect 8515 29128 8524 29168
rect 8564 29128 8573 29168
rect 8515 29127 8573 29128
rect 8611 29168 8669 29169
rect 8611 29128 8620 29168
rect 8660 29128 8669 29168
rect 8611 29127 8669 29128
rect 8811 29168 8853 29177
rect 8811 29128 8812 29168
rect 8852 29128 8853 29168
rect 8811 29119 8853 29128
rect 8907 29168 8949 29177
rect 8907 29128 8908 29168
rect 8948 29128 8949 29168
rect 8907 29119 8949 29128
rect 9000 29168 9058 29169
rect 9000 29128 9009 29168
rect 9049 29128 9058 29168
rect 9000 29127 9058 29128
rect 9667 29168 9725 29169
rect 9667 29128 9676 29168
rect 9716 29128 9725 29168
rect 9667 29127 9725 29128
rect 10915 29168 10973 29169
rect 10915 29128 10924 29168
rect 10964 29128 10973 29168
rect 10915 29127 10973 29128
rect 11299 29168 11357 29169
rect 11299 29128 11308 29168
rect 11348 29128 11357 29168
rect 11299 29127 11357 29128
rect 11595 29168 11637 29177
rect 11595 29128 11596 29168
rect 11636 29128 11637 29168
rect 11595 29119 11637 29128
rect 11691 29168 11733 29177
rect 11691 29128 11692 29168
rect 11732 29128 11733 29168
rect 11691 29119 11733 29128
rect 13507 29168 13565 29169
rect 13507 29128 13516 29168
rect 13556 29128 13565 29168
rect 13995 29148 13996 29188
rect 14036 29148 14037 29188
rect 13995 29139 14037 29148
rect 14091 29188 14133 29197
rect 14091 29148 14092 29188
rect 14132 29148 14133 29188
rect 14091 29139 14133 29148
rect 14475 29168 14517 29177
rect 13507 29127 13565 29128
rect 14475 29128 14476 29168
rect 14516 29128 14517 29168
rect 12259 29126 12317 29127
rect 12259 29086 12268 29126
rect 12308 29086 12317 29126
rect 14475 29119 14517 29128
rect 14571 29168 14613 29177
rect 14571 29128 14572 29168
rect 14612 29128 14613 29168
rect 14571 29119 14613 29128
rect 15043 29168 15101 29169
rect 15043 29128 15052 29168
rect 15092 29128 15101 29168
rect 16579 29168 16637 29169
rect 15043 29127 15101 29128
rect 15531 29154 15573 29163
rect 15531 29114 15532 29154
rect 15572 29114 15573 29154
rect 16579 29128 16588 29168
rect 16628 29128 16637 29168
rect 16579 29127 16637 29128
rect 17827 29168 17885 29169
rect 17827 29128 17836 29168
rect 17876 29128 17885 29168
rect 17827 29127 17885 29128
rect 18219 29168 18261 29177
rect 18219 29128 18220 29168
rect 18260 29128 18261 29168
rect 18219 29119 18261 29128
rect 18411 29168 18453 29177
rect 18411 29128 18412 29168
rect 18452 29128 18453 29168
rect 18411 29119 18453 29128
rect 18499 29168 18557 29169
rect 18499 29128 18508 29168
rect 18548 29128 18557 29168
rect 18499 29127 18557 29128
rect 19171 29168 19229 29169
rect 19171 29128 19180 29168
rect 19220 29128 19229 29168
rect 19171 29127 19229 29128
rect 19467 29168 19509 29177
rect 19467 29128 19468 29168
rect 19508 29128 19509 29168
rect 19467 29119 19509 29128
rect 15531 29105 15573 29114
rect 12259 29085 12317 29086
rect 18691 29084 18749 29085
rect 18691 29044 18700 29084
rect 18740 29044 18749 29084
rect 18691 29043 18749 29044
rect 20035 29084 20093 29085
rect 20035 29044 20044 29084
rect 20084 29044 20093 29084
rect 20035 29043 20093 29044
rect 6019 29000 6077 29001
rect 6019 28960 6028 29000
rect 6068 28960 6077 29000
rect 6019 28959 6077 28960
rect 7851 29000 7893 29009
rect 7851 28960 7852 29000
rect 7892 28960 7893 29000
rect 7851 28951 7893 28960
rect 19843 29000 19901 29001
rect 19843 28960 19852 29000
rect 19892 28960 19901 29000
rect 19843 28959 19901 28960
rect 3531 28916 3573 28925
rect 3531 28876 3532 28916
rect 3572 28876 3573 28916
rect 3531 28867 3573 28876
rect 5355 28916 5397 28925
rect 5355 28876 5356 28916
rect 5396 28876 5397 28916
rect 5355 28867 5397 28876
rect 9483 28916 9525 28925
rect 9483 28876 9484 28916
rect 9524 28876 9525 28916
rect 9483 28867 9525 28876
rect 11971 28916 12029 28917
rect 11971 28876 11980 28916
rect 12020 28876 12029 28916
rect 11971 28875 12029 28876
rect 18027 28916 18069 28925
rect 18027 28876 18028 28916
rect 18068 28876 18069 28916
rect 18027 28867 18069 28876
rect 20235 28916 20277 28925
rect 20235 28876 20236 28916
rect 20276 28876 20277 28916
rect 20235 28867 20277 28876
rect 1152 28748 20352 28772
rect 1152 28708 3688 28748
rect 3728 28708 3770 28748
rect 3810 28708 3852 28748
rect 3892 28708 3934 28748
rect 3974 28708 4016 28748
rect 4056 28708 18808 28748
rect 18848 28708 18890 28748
rect 18930 28708 18972 28748
rect 19012 28708 19054 28748
rect 19094 28708 19136 28748
rect 19176 28708 20352 28748
rect 1152 28684 20352 28708
rect 7179 28580 7221 28589
rect 7179 28540 7180 28580
rect 7220 28540 7221 28580
rect 7179 28531 7221 28540
rect 16107 28580 16149 28589
rect 16107 28540 16108 28580
rect 16148 28540 16149 28580
rect 16107 28531 16149 28540
rect 12171 28496 12213 28505
rect 12171 28456 12172 28496
rect 12212 28456 12213 28496
rect 12171 28447 12213 28456
rect 1995 28412 2037 28421
rect 1995 28372 1996 28412
rect 2036 28372 2037 28412
rect 1995 28363 2037 28372
rect 3915 28412 3957 28421
rect 3915 28372 3916 28412
rect 3956 28372 3957 28412
rect 3915 28363 3957 28372
rect 16971 28412 17013 28421
rect 16971 28372 16972 28412
rect 17012 28372 17013 28412
rect 6979 28370 7037 28371
rect 2955 28342 2997 28351
rect 1419 28328 1461 28337
rect 1419 28288 1420 28328
rect 1460 28288 1461 28328
rect 1419 28279 1461 28288
rect 1515 28328 1557 28337
rect 1515 28288 1516 28328
rect 1556 28288 1557 28328
rect 1515 28279 1557 28288
rect 1899 28328 1941 28337
rect 1899 28288 1900 28328
rect 1940 28288 1941 28328
rect 1899 28279 1941 28288
rect 2467 28328 2525 28329
rect 2467 28288 2476 28328
rect 2516 28288 2525 28328
rect 2955 28302 2956 28342
rect 2996 28302 2997 28342
rect 4971 28342 5013 28351
rect 2955 28293 2997 28302
rect 3435 28328 3477 28337
rect 2467 28287 2525 28288
rect 3435 28288 3436 28328
rect 3476 28288 3477 28328
rect 3435 28279 3477 28288
rect 3531 28328 3573 28337
rect 3531 28288 3532 28328
rect 3572 28288 3573 28328
rect 3531 28279 3573 28288
rect 4011 28328 4053 28337
rect 4011 28288 4012 28328
rect 4052 28288 4053 28328
rect 4011 28279 4053 28288
rect 4483 28328 4541 28329
rect 4483 28288 4492 28328
rect 4532 28288 4541 28328
rect 4971 28302 4972 28342
rect 5012 28302 5013 28342
rect 6979 28330 6988 28370
rect 7028 28330 7037 28370
rect 16971 28363 17013 28372
rect 17067 28412 17109 28421
rect 17067 28372 17068 28412
rect 17108 28372 17109 28412
rect 17067 28363 17109 28372
rect 6979 28329 7037 28330
rect 7467 28347 7509 28356
rect 4971 28293 5013 28302
rect 5731 28328 5789 28329
rect 4483 28287 4541 28288
rect 5731 28288 5740 28328
rect 5780 28288 5789 28328
rect 7467 28307 7468 28347
rect 7508 28307 7509 28347
rect 9003 28342 9045 28351
rect 18027 28342 18069 28351
rect 7467 28298 7509 28307
rect 7563 28328 7605 28337
rect 5731 28287 5789 28288
rect 7563 28288 7564 28328
rect 7604 28288 7605 28328
rect 7563 28279 7605 28288
rect 7947 28328 7989 28337
rect 7947 28288 7948 28328
rect 7988 28288 7989 28328
rect 7947 28279 7989 28288
rect 8043 28328 8085 28337
rect 8043 28288 8044 28328
rect 8084 28288 8085 28328
rect 8043 28279 8085 28288
rect 8515 28328 8573 28329
rect 8515 28288 8524 28328
rect 8564 28288 8573 28328
rect 9003 28302 9004 28342
rect 9044 28302 9045 28342
rect 9003 28293 9045 28302
rect 9483 28328 9525 28337
rect 8515 28287 8573 28288
rect 9483 28288 9484 28328
rect 9524 28288 9525 28328
rect 9483 28279 9525 28288
rect 9579 28328 9621 28337
rect 9579 28288 9580 28328
rect 9620 28288 9621 28328
rect 9579 28279 9621 28288
rect 9963 28328 10005 28337
rect 9963 28288 9964 28328
rect 10004 28288 10005 28328
rect 9963 28279 10005 28288
rect 10059 28328 10101 28337
rect 11019 28333 11061 28342
rect 10059 28288 10060 28328
rect 10100 28288 10101 28328
rect 10059 28279 10101 28288
rect 10531 28328 10589 28329
rect 10531 28288 10540 28328
rect 10580 28288 10589 28328
rect 10531 28287 10589 28288
rect 11019 28293 11020 28333
rect 11060 28293 11061 28333
rect 11019 28284 11061 28293
rect 11395 28328 11453 28329
rect 11395 28288 11404 28328
rect 11444 28288 11453 28328
rect 11395 28287 11453 28288
rect 11779 28328 11837 28329
rect 11779 28288 11788 28328
rect 11828 28288 11837 28328
rect 11779 28287 11837 28288
rect 11883 28328 11925 28337
rect 11883 28288 11884 28328
rect 11924 28288 11925 28328
rect 11883 28279 11925 28288
rect 12363 28328 12405 28337
rect 12363 28288 12364 28328
rect 12404 28288 12405 28328
rect 12363 28279 12405 28288
rect 12555 28328 12597 28337
rect 12555 28288 12556 28328
rect 12596 28288 12597 28328
rect 12555 28279 12597 28288
rect 12643 28328 12701 28329
rect 12643 28288 12652 28328
rect 12692 28288 12701 28328
rect 12643 28287 12701 28288
rect 12843 28328 12885 28337
rect 12843 28288 12844 28328
rect 12884 28288 12885 28328
rect 12843 28279 12885 28288
rect 13035 28328 13077 28337
rect 13035 28288 13036 28328
rect 13076 28288 13077 28328
rect 13035 28279 13077 28288
rect 13123 28328 13181 28329
rect 13123 28288 13132 28328
rect 13172 28288 13181 28328
rect 13123 28287 13181 28288
rect 14467 28328 14525 28329
rect 14467 28288 14476 28328
rect 14516 28288 14525 28328
rect 14467 28287 14525 28288
rect 14659 28328 14717 28329
rect 14659 28288 14668 28328
rect 14708 28288 14717 28328
rect 14659 28287 14717 28288
rect 15907 28328 15965 28329
rect 15907 28288 15916 28328
rect 15956 28288 15965 28328
rect 15907 28287 15965 28288
rect 16491 28328 16533 28337
rect 16491 28288 16492 28328
rect 16532 28288 16533 28328
rect 16491 28279 16533 28288
rect 16587 28328 16629 28337
rect 16587 28288 16588 28328
rect 16628 28288 16629 28328
rect 16587 28279 16629 28288
rect 17539 28328 17597 28329
rect 17539 28288 17548 28328
rect 17588 28288 17597 28328
rect 18027 28302 18028 28342
rect 18068 28302 18069 28342
rect 18027 28293 18069 28302
rect 18499 28328 18557 28329
rect 17539 28287 17597 28288
rect 18499 28288 18508 28328
rect 18548 28288 18557 28328
rect 18499 28287 18557 28288
rect 19747 28328 19805 28329
rect 19747 28288 19756 28328
rect 19796 28288 19805 28328
rect 19747 28287 19805 28288
rect 3147 28244 3189 28253
rect 3147 28204 3148 28244
rect 3188 28204 3189 28244
rect 3147 28195 3189 28204
rect 5163 28244 5205 28253
rect 5163 28204 5164 28244
rect 5204 28204 5205 28244
rect 5163 28195 5205 28204
rect 9195 28244 9237 28253
rect 9195 28204 9196 28244
rect 9236 28204 9237 28244
rect 9195 28195 9237 28204
rect 11211 28244 11253 28253
rect 11211 28204 11212 28244
rect 11252 28204 11253 28244
rect 11211 28195 11253 28204
rect 11499 28160 11541 28169
rect 11499 28120 11500 28160
rect 11540 28120 11541 28160
rect 11499 28111 11541 28120
rect 11691 28156 11733 28165
rect 11691 28116 11692 28156
rect 11732 28116 11733 28156
rect 12451 28160 12509 28161
rect 12451 28120 12460 28160
rect 12500 28120 12509 28160
rect 12451 28119 12509 28120
rect 12931 28160 12989 28161
rect 12931 28120 12940 28160
rect 12980 28120 12989 28160
rect 12931 28119 12989 28120
rect 14379 28160 14421 28169
rect 14379 28120 14380 28160
rect 14420 28120 14421 28160
rect 11691 28107 11733 28116
rect 14379 28111 14421 28120
rect 18219 28160 18261 28169
rect 18219 28120 18220 28160
rect 18260 28120 18261 28160
rect 18219 28111 18261 28120
rect 19947 28160 19989 28169
rect 19947 28120 19948 28160
rect 19988 28120 19989 28160
rect 19947 28111 19989 28120
rect 1152 27992 20452 28016
rect 1152 27952 4928 27992
rect 4968 27952 5010 27992
rect 5050 27952 5092 27992
rect 5132 27952 5174 27992
rect 5214 27952 5256 27992
rect 5296 27952 20048 27992
rect 20088 27952 20130 27992
rect 20170 27952 20212 27992
rect 20252 27952 20294 27992
rect 20334 27952 20376 27992
rect 20416 27952 20452 27992
rect 1152 27928 20452 27952
rect 3339 27824 3381 27833
rect 3339 27784 3340 27824
rect 3380 27784 3381 27824
rect 3339 27775 3381 27784
rect 11883 27824 11925 27833
rect 11883 27784 11884 27824
rect 11924 27784 11925 27824
rect 11883 27775 11925 27784
rect 12355 27824 12413 27825
rect 12355 27784 12364 27824
rect 12404 27784 12413 27824
rect 12355 27783 12413 27784
rect 18507 27824 18549 27833
rect 18507 27784 18508 27824
rect 18548 27784 18549 27824
rect 18507 27775 18549 27784
rect 5835 27740 5877 27749
rect 5835 27700 5836 27740
rect 5876 27700 5877 27740
rect 5835 27691 5877 27700
rect 9099 27740 9141 27749
rect 9099 27700 9100 27740
rect 9140 27700 9141 27740
rect 9099 27691 9141 27700
rect 17163 27740 17205 27749
rect 17163 27700 17164 27740
rect 17204 27700 17205 27740
rect 17163 27691 17205 27700
rect 19563 27740 19605 27749
rect 19563 27700 19564 27740
rect 19604 27700 19605 27740
rect 19563 27691 19605 27700
rect 1699 27656 1757 27657
rect 1699 27616 1708 27656
rect 1748 27616 1757 27656
rect 1699 27615 1757 27616
rect 2947 27656 3005 27657
rect 2947 27616 2956 27656
rect 2996 27616 3005 27656
rect 2947 27615 3005 27616
rect 3523 27656 3581 27657
rect 3523 27616 3532 27656
rect 3572 27616 3581 27656
rect 3523 27615 3581 27616
rect 4771 27656 4829 27657
rect 4771 27616 4780 27656
rect 4820 27616 4829 27656
rect 4771 27615 4829 27616
rect 5443 27656 5501 27657
rect 5443 27616 5452 27656
rect 5492 27616 5501 27656
rect 5443 27615 5501 27616
rect 5739 27656 5781 27665
rect 5739 27616 5740 27656
rect 5780 27616 5781 27656
rect 5739 27607 5781 27616
rect 6691 27656 6749 27657
rect 6691 27616 6700 27656
rect 6740 27616 6749 27656
rect 6691 27615 6749 27616
rect 7939 27656 7997 27657
rect 7939 27616 7948 27656
rect 7988 27616 7997 27656
rect 7939 27615 7997 27616
rect 8523 27656 8565 27665
rect 8523 27616 8524 27656
rect 8564 27616 8565 27656
rect 8523 27607 8565 27616
rect 8811 27656 8853 27665
rect 8811 27616 8812 27656
rect 8852 27616 8853 27656
rect 8811 27607 8853 27616
rect 8995 27656 9053 27657
rect 8995 27616 9004 27656
rect 9044 27616 9053 27656
rect 9579 27656 9621 27665
rect 8995 27615 9053 27616
rect 9387 27645 9429 27654
rect 9387 27605 9388 27645
rect 9428 27605 9429 27645
rect 9579 27616 9580 27656
rect 9620 27616 9621 27656
rect 9579 27607 9621 27616
rect 9667 27656 9725 27657
rect 9667 27616 9676 27656
rect 9716 27616 9725 27656
rect 9667 27615 9725 27616
rect 10435 27656 10493 27657
rect 10435 27616 10444 27656
rect 10484 27616 10493 27656
rect 10435 27615 10493 27616
rect 11683 27656 11741 27657
rect 11683 27616 11692 27656
rect 11732 27616 11741 27656
rect 11683 27615 11741 27616
rect 12075 27656 12117 27665
rect 12075 27616 12076 27656
rect 12116 27616 12117 27656
rect 12075 27607 12117 27616
rect 12171 27656 12213 27665
rect 12171 27616 12172 27656
rect 12212 27616 12213 27656
rect 12171 27607 12213 27616
rect 12267 27656 12309 27665
rect 12267 27616 12268 27656
rect 12308 27616 12309 27656
rect 12267 27607 12309 27616
rect 13507 27656 13565 27657
rect 13507 27616 13516 27656
rect 13556 27616 13565 27656
rect 13507 27615 13565 27616
rect 14755 27656 14813 27657
rect 14755 27616 14764 27656
rect 14804 27616 14813 27656
rect 14755 27615 14813 27616
rect 15147 27656 15189 27665
rect 15147 27616 15148 27656
rect 15188 27616 15189 27656
rect 15147 27607 15189 27616
rect 15243 27656 15285 27665
rect 15243 27616 15244 27656
rect 15284 27616 15285 27656
rect 15243 27607 15285 27616
rect 15339 27656 15381 27665
rect 15339 27616 15340 27656
rect 15380 27616 15381 27656
rect 15339 27607 15381 27616
rect 15435 27656 15477 27665
rect 15435 27616 15436 27656
rect 15476 27616 15477 27656
rect 15435 27607 15477 27616
rect 15715 27656 15773 27657
rect 15715 27616 15724 27656
rect 15764 27616 15773 27656
rect 15715 27615 15773 27616
rect 16963 27656 17021 27657
rect 16963 27616 16972 27656
rect 17012 27616 17021 27656
rect 16963 27615 17021 27616
rect 17547 27656 17589 27665
rect 17547 27616 17548 27656
rect 17588 27616 17589 27656
rect 17547 27607 17589 27616
rect 17835 27656 17877 27665
rect 17835 27616 17836 27656
rect 17876 27616 17877 27656
rect 17835 27607 17877 27616
rect 18123 27656 18165 27665
rect 18123 27616 18124 27656
rect 18164 27616 18165 27656
rect 18123 27607 18165 27616
rect 18219 27656 18261 27665
rect 18219 27616 18220 27656
rect 18260 27616 18261 27656
rect 18219 27607 18261 27616
rect 18315 27656 18357 27665
rect 18315 27616 18316 27656
rect 18356 27616 18357 27656
rect 18315 27607 18357 27616
rect 19171 27656 19229 27657
rect 19171 27616 19180 27656
rect 19220 27616 19229 27656
rect 19171 27615 19229 27616
rect 19467 27656 19509 27665
rect 19467 27616 19468 27656
rect 19508 27616 19509 27656
rect 19467 27607 19509 27616
rect 9387 27596 9429 27605
rect 18691 27572 18749 27573
rect 18691 27532 18700 27572
rect 18740 27532 18749 27572
rect 18691 27531 18749 27532
rect 6115 27488 6173 27489
rect 6115 27448 6124 27488
rect 6164 27448 6173 27488
rect 6115 27447 6173 27448
rect 8139 27488 8181 27497
rect 8139 27448 8140 27488
rect 8180 27448 8181 27488
rect 8139 27439 8181 27448
rect 8811 27488 8853 27497
rect 8811 27448 8812 27488
rect 8852 27448 8853 27488
rect 8811 27439 8853 27448
rect 17835 27488 17877 27497
rect 17835 27448 17836 27488
rect 17876 27448 17877 27488
rect 17835 27439 17877 27448
rect 18891 27488 18933 27497
rect 18891 27448 18892 27488
rect 18932 27448 18933 27488
rect 18891 27439 18933 27448
rect 3147 27404 3189 27413
rect 3147 27364 3148 27404
rect 3188 27364 3189 27404
rect 3147 27355 3189 27364
rect 9387 27404 9429 27413
rect 9387 27364 9388 27404
rect 9428 27364 9429 27404
rect 9387 27355 9429 27364
rect 14955 27404 14997 27413
rect 14955 27364 14956 27404
rect 14996 27364 14997 27404
rect 14955 27355 14997 27364
rect 19843 27404 19901 27405
rect 19843 27364 19852 27404
rect 19892 27364 19901 27404
rect 19843 27363 19901 27364
rect 1152 27236 20352 27260
rect 1152 27196 3688 27236
rect 3728 27196 3770 27236
rect 3810 27196 3852 27236
rect 3892 27196 3934 27236
rect 3974 27196 4016 27236
rect 4056 27196 18808 27236
rect 18848 27196 18890 27236
rect 18930 27196 18972 27236
rect 19012 27196 19054 27236
rect 19094 27196 19136 27236
rect 19176 27196 20352 27236
rect 1152 27172 20352 27196
rect 14187 27068 14229 27077
rect 14187 27028 14188 27068
rect 14228 27028 14229 27068
rect 14187 27019 14229 27028
rect 15915 27068 15957 27077
rect 15915 27028 15916 27068
rect 15956 27028 15957 27068
rect 15915 27019 15957 27028
rect 6211 26984 6269 26985
rect 6211 26944 6220 26984
rect 6260 26944 6269 26984
rect 6211 26943 6269 26944
rect 15139 26984 15197 26985
rect 15139 26944 15148 26984
rect 15188 26944 15197 26984
rect 15139 26943 15197 26944
rect 15531 26984 15573 26993
rect 15531 26944 15532 26984
rect 15572 26944 15573 26984
rect 15531 26935 15573 26944
rect 16107 26984 16149 26993
rect 16107 26944 16108 26984
rect 16148 26944 16149 26984
rect 16107 26935 16149 26944
rect 16395 26984 16437 26993
rect 16395 26944 16396 26984
rect 16436 26944 16437 26984
rect 16395 26935 16437 26944
rect 19947 26984 19989 26993
rect 19947 26944 19948 26984
rect 19988 26944 19989 26984
rect 19947 26935 19989 26944
rect 15428 26910 15486 26911
rect 11883 26900 11925 26909
rect 11883 26860 11884 26900
rect 11924 26860 11925 26900
rect 15428 26870 15437 26910
rect 15477 26870 15486 26910
rect 15428 26869 15486 26870
rect 15627 26900 15669 26909
rect 11883 26851 11925 26860
rect 15627 26860 15628 26900
rect 15668 26860 15669 26900
rect 19363 26900 19421 26901
rect 15627 26851 15669 26860
rect 15723 26858 15765 26867
rect 19363 26860 19372 26900
rect 19412 26860 19421 26900
rect 19363 26859 19421 26860
rect 19747 26900 19805 26901
rect 19747 26860 19756 26900
rect 19796 26860 19805 26900
rect 19747 26859 19805 26860
rect 1219 26816 1277 26817
rect 1219 26776 1228 26816
rect 1268 26776 1277 26816
rect 1219 26775 1277 26776
rect 2467 26816 2525 26817
rect 2467 26776 2476 26816
rect 2516 26776 2525 26816
rect 2467 26775 2525 26776
rect 3627 26816 3669 26825
rect 3627 26776 3628 26816
rect 3668 26776 3669 26816
rect 3627 26767 3669 26776
rect 3915 26816 3957 26825
rect 3915 26776 3916 26816
rect 3956 26776 3957 26816
rect 3915 26767 3957 26776
rect 4099 26816 4157 26817
rect 4099 26776 4108 26816
rect 4148 26776 4157 26816
rect 4099 26775 4157 26776
rect 5347 26816 5405 26817
rect 5347 26776 5356 26816
rect 5396 26776 5405 26816
rect 5347 26775 5405 26776
rect 5835 26816 5877 26825
rect 5835 26776 5836 26816
rect 5876 26776 5877 26816
rect 5835 26767 5877 26776
rect 5931 26816 5973 26825
rect 5931 26776 5932 26816
rect 5972 26776 5973 26816
rect 5931 26767 5973 26776
rect 6027 26816 6069 26825
rect 6027 26776 6028 26816
rect 6068 26776 6069 26816
rect 6027 26767 6069 26776
rect 6411 26816 6453 26825
rect 6411 26776 6412 26816
rect 6452 26776 6453 26816
rect 6411 26767 6453 26776
rect 6507 26816 6549 26825
rect 6507 26776 6508 26816
rect 6548 26776 6549 26816
rect 6507 26767 6549 26776
rect 6603 26816 6645 26825
rect 6603 26776 6604 26816
rect 6644 26776 6645 26816
rect 6603 26767 6645 26776
rect 7075 26816 7133 26817
rect 7075 26776 7084 26816
rect 7124 26776 7133 26816
rect 7075 26775 7133 26776
rect 8323 26816 8381 26817
rect 8323 26776 8332 26816
rect 8372 26776 8381 26816
rect 8323 26775 8381 26776
rect 8995 26816 9053 26817
rect 8995 26776 9004 26816
rect 9044 26776 9053 26816
rect 8995 26775 9053 26776
rect 10243 26816 10301 26817
rect 10243 26776 10252 26816
rect 10292 26776 10301 26816
rect 10243 26775 10301 26776
rect 10731 26816 10773 26825
rect 10731 26776 10732 26816
rect 10772 26776 10773 26816
rect 10731 26767 10773 26776
rect 10827 26816 10869 26825
rect 10827 26776 10828 26816
rect 10868 26776 10869 26816
rect 10827 26767 10869 26776
rect 10923 26816 10965 26825
rect 10923 26776 10924 26816
rect 10964 26776 10965 26816
rect 10923 26767 10965 26776
rect 11307 26816 11349 26825
rect 11307 26776 11308 26816
rect 11348 26776 11349 26816
rect 11307 26767 11349 26776
rect 11403 26816 11445 26825
rect 11403 26776 11404 26816
rect 11444 26776 11445 26816
rect 11403 26767 11445 26776
rect 11499 26816 11541 26825
rect 11499 26776 11500 26816
rect 11540 26776 11541 26816
rect 11499 26767 11541 26776
rect 11779 26816 11837 26817
rect 11779 26776 11788 26816
rect 11828 26776 11837 26816
rect 11779 26775 11837 26776
rect 12355 26816 12413 26817
rect 12355 26776 12364 26816
rect 12404 26776 12413 26816
rect 12355 26775 12413 26776
rect 13603 26816 13661 26817
rect 13603 26776 13612 26816
rect 13652 26776 13661 26816
rect 13603 26775 13661 26776
rect 14083 26816 14141 26817
rect 14083 26776 14092 26816
rect 14132 26776 14141 26816
rect 14083 26775 14141 26776
rect 14467 26816 14525 26817
rect 14467 26776 14476 26816
rect 14516 26776 14525 26816
rect 14467 26775 14525 26776
rect 14763 26816 14805 26825
rect 14763 26776 14764 26816
rect 14804 26776 14805 26816
rect 14763 26767 14805 26776
rect 14859 26816 14901 26825
rect 15723 26818 15724 26858
rect 15764 26818 15765 26858
rect 14859 26776 14860 26816
rect 14900 26776 14901 26816
rect 14859 26767 14901 26776
rect 15331 26816 15389 26817
rect 15331 26776 15340 26816
rect 15380 26776 15389 26816
rect 15723 26809 15765 26818
rect 16107 26816 16149 26825
rect 15331 26775 15389 26776
rect 16107 26776 16108 26816
rect 16148 26776 16149 26816
rect 16107 26767 16149 26776
rect 16395 26816 16437 26825
rect 16395 26776 16396 26816
rect 16436 26776 16437 26816
rect 16395 26767 16437 26776
rect 16587 26816 16629 26825
rect 16587 26776 16588 26816
rect 16628 26776 16629 26816
rect 16587 26767 16629 26776
rect 16675 26816 16733 26817
rect 16675 26776 16684 26816
rect 16724 26776 16733 26816
rect 16675 26775 16733 26776
rect 18411 26816 18453 26825
rect 18411 26776 18412 26816
rect 18452 26776 18453 26816
rect 18411 26767 18453 26776
rect 18595 26816 18653 26817
rect 18595 26776 18604 26816
rect 18644 26776 18653 26816
rect 18595 26775 18653 26776
rect 18795 26816 18837 26825
rect 18795 26776 18796 26816
rect 18836 26776 18837 26816
rect 18795 26767 18837 26776
rect 18891 26816 18933 26825
rect 18891 26776 18892 26816
rect 18932 26776 18933 26816
rect 18891 26767 18933 26776
rect 8523 26732 8565 26741
rect 8523 26692 8524 26732
rect 8564 26692 8565 26732
rect 8523 26683 8565 26692
rect 13803 26732 13845 26741
rect 13803 26692 13804 26732
rect 13844 26692 13845 26732
rect 13803 26683 13845 26692
rect 18507 26732 18549 26741
rect 18507 26692 18508 26732
rect 18548 26692 18549 26732
rect 18507 26683 18549 26692
rect 2667 26648 2709 26657
rect 2667 26608 2668 26648
rect 2708 26608 2709 26648
rect 2667 26599 2709 26608
rect 3819 26648 3861 26657
rect 3819 26608 3820 26648
rect 3860 26608 3861 26648
rect 3819 26599 3861 26608
rect 5547 26648 5589 26657
rect 5547 26608 5548 26648
rect 5588 26608 5589 26648
rect 5547 26599 5589 26608
rect 6691 26648 6749 26649
rect 6691 26608 6700 26648
rect 6740 26608 6749 26648
rect 6691 26607 6749 26608
rect 10443 26648 10485 26657
rect 10443 26608 10444 26648
rect 10484 26608 10485 26648
rect 10443 26599 10485 26608
rect 11115 26648 11157 26657
rect 11115 26608 11116 26648
rect 11156 26608 11157 26648
rect 11115 26599 11157 26608
rect 11587 26648 11645 26649
rect 11587 26608 11596 26648
rect 11636 26608 11645 26648
rect 11587 26607 11645 26608
rect 14187 26648 14229 26657
rect 14187 26608 14188 26648
rect 14228 26608 14229 26648
rect 14187 26599 14229 26608
rect 19075 26648 19133 26649
rect 19075 26608 19084 26648
rect 19124 26608 19133 26648
rect 19075 26607 19133 26608
rect 19563 26648 19605 26657
rect 19563 26608 19564 26648
rect 19604 26608 19605 26648
rect 19563 26599 19605 26608
rect 1152 26480 20452 26504
rect 1152 26440 4928 26480
rect 4968 26440 5010 26480
rect 5050 26440 5092 26480
rect 5132 26440 5174 26480
rect 5214 26440 5256 26480
rect 5296 26440 20048 26480
rect 20088 26440 20130 26480
rect 20170 26440 20212 26480
rect 20252 26440 20294 26480
rect 20334 26440 20376 26480
rect 20416 26440 20452 26480
rect 1152 26416 20452 26440
rect 4971 26312 5013 26321
rect 4971 26272 4972 26312
rect 5012 26272 5013 26312
rect 4971 26263 5013 26272
rect 13995 26312 14037 26321
rect 13995 26272 13996 26312
rect 14036 26272 14037 26312
rect 13995 26263 14037 26272
rect 14467 26312 14525 26313
rect 14467 26272 14476 26312
rect 14516 26272 14525 26312
rect 14467 26271 14525 26272
rect 15723 26312 15765 26321
rect 15723 26272 15724 26312
rect 15764 26272 15765 26312
rect 15723 26263 15765 26272
rect 18987 26312 19029 26321
rect 18987 26272 18988 26312
rect 19028 26272 19029 26312
rect 18987 26263 19029 26272
rect 6123 26228 6165 26237
rect 6123 26188 6124 26228
rect 6164 26188 6165 26228
rect 6123 26179 6165 26188
rect 10635 26228 10677 26237
rect 10635 26188 10636 26228
rect 10676 26188 10677 26228
rect 10635 26179 10677 26188
rect 1507 26144 1565 26145
rect 1507 26104 1516 26144
rect 1556 26104 1565 26144
rect 1507 26103 1565 26104
rect 2755 26144 2813 26145
rect 2755 26104 2764 26144
rect 2804 26104 2813 26144
rect 2755 26103 2813 26104
rect 3243 26144 3285 26153
rect 3243 26104 3244 26144
rect 3284 26104 3285 26144
rect 3243 26095 3285 26104
rect 3339 26144 3381 26153
rect 3339 26104 3340 26144
rect 3380 26104 3381 26144
rect 3339 26095 3381 26104
rect 3819 26144 3861 26153
rect 3819 26104 3820 26144
rect 3860 26104 3861 26144
rect 3819 26095 3861 26104
rect 4291 26144 4349 26145
rect 4291 26104 4300 26144
rect 4340 26104 4349 26144
rect 4291 26103 4349 26104
rect 4779 26139 4821 26148
rect 4779 26099 4780 26139
rect 4820 26099 4821 26139
rect 4779 26090 4821 26099
rect 5163 26144 5205 26153
rect 5163 26104 5164 26144
rect 5204 26104 5205 26144
rect 5163 26095 5205 26104
rect 5355 26144 5397 26153
rect 5355 26104 5356 26144
rect 5396 26104 5397 26144
rect 5355 26095 5397 26104
rect 5443 26144 5501 26145
rect 5443 26104 5452 26144
rect 5492 26104 5501 26144
rect 5443 26103 5501 26104
rect 5731 26144 5789 26145
rect 5731 26104 5740 26144
rect 5780 26104 5789 26144
rect 5731 26103 5789 26104
rect 6027 26144 6069 26153
rect 6027 26104 6028 26144
rect 6068 26104 6069 26144
rect 6027 26095 6069 26104
rect 8907 26144 8949 26153
rect 8907 26104 8908 26144
rect 8948 26104 8949 26144
rect 8907 26095 8949 26104
rect 9003 26144 9045 26153
rect 9003 26104 9004 26144
rect 9044 26104 9045 26144
rect 9003 26095 9045 26104
rect 9387 26144 9429 26153
rect 9387 26104 9388 26144
rect 9428 26104 9429 26144
rect 9387 26095 9429 26104
rect 9955 26144 10013 26145
rect 9955 26104 9964 26144
rect 10004 26104 10013 26144
rect 9955 26103 10013 26104
rect 10443 26139 10485 26148
rect 10443 26099 10444 26139
rect 10484 26099 10485 26139
rect 10819 26144 10877 26145
rect 10819 26104 10828 26144
rect 10868 26104 10877 26144
rect 10819 26103 10877 26104
rect 12067 26144 12125 26145
rect 12067 26104 12076 26144
rect 12116 26104 12125 26144
rect 12067 26103 12125 26104
rect 12547 26144 12605 26145
rect 12547 26104 12556 26144
rect 12596 26104 12605 26144
rect 12547 26103 12605 26104
rect 13795 26144 13853 26145
rect 13795 26104 13804 26144
rect 13844 26104 13853 26144
rect 13795 26103 13853 26104
rect 14187 26144 14229 26153
rect 14187 26104 14188 26144
rect 14228 26104 14229 26144
rect 10443 26090 10485 26099
rect 14187 26095 14229 26104
rect 14283 26144 14325 26153
rect 14283 26104 14284 26144
rect 14324 26104 14325 26144
rect 14283 26095 14325 26104
rect 14379 26144 14421 26153
rect 14379 26104 14380 26144
rect 14420 26104 14421 26144
rect 14379 26095 14421 26104
rect 14755 26144 14813 26145
rect 14755 26104 14764 26144
rect 14804 26104 14813 26144
rect 14755 26103 14813 26104
rect 15051 26144 15093 26153
rect 15051 26104 15052 26144
rect 15092 26104 15093 26144
rect 15051 26095 15093 26104
rect 15147 26144 15189 26153
rect 15147 26104 15148 26144
rect 15188 26104 15189 26144
rect 15147 26095 15189 26104
rect 15619 26144 15677 26145
rect 15619 26104 15628 26144
rect 15668 26104 15677 26144
rect 15619 26103 15677 26104
rect 15907 26144 15965 26145
rect 15907 26104 15916 26144
rect 15956 26104 15965 26144
rect 15907 26103 15965 26104
rect 17155 26144 17213 26145
rect 17155 26104 17164 26144
rect 17204 26104 17213 26144
rect 17155 26103 17213 26104
rect 17539 26144 17597 26145
rect 17539 26104 17548 26144
rect 17588 26104 17597 26144
rect 17539 26103 17597 26104
rect 18787 26144 18845 26145
rect 18787 26104 18796 26144
rect 18836 26104 18845 26144
rect 18787 26103 18845 26104
rect 19179 26144 19221 26153
rect 19179 26104 19180 26144
rect 19220 26104 19221 26144
rect 19179 26095 19221 26104
rect 19275 26144 19317 26153
rect 19275 26104 19276 26144
rect 19316 26104 19317 26144
rect 19275 26095 19317 26104
rect 19371 26144 19413 26153
rect 19371 26104 19372 26144
rect 19412 26104 19413 26144
rect 19371 26095 19413 26104
rect 19467 26144 19509 26153
rect 19467 26104 19468 26144
rect 19508 26104 19509 26144
rect 19467 26095 19509 26104
rect 3723 26060 3765 26069
rect 3723 26020 3724 26060
rect 3764 26020 3765 26060
rect 3723 26011 3765 26020
rect 9483 26060 9525 26069
rect 9483 26020 9484 26060
rect 9524 26020 9525 26060
rect 9483 26011 9525 26020
rect 19651 26060 19709 26061
rect 19651 26020 19660 26060
rect 19700 26020 19709 26060
rect 19651 26019 19709 26020
rect 20035 26060 20093 26061
rect 20035 26020 20044 26060
rect 20084 26020 20093 26060
rect 20035 26019 20093 26020
rect 5163 25976 5205 25985
rect 5163 25936 5164 25976
rect 5204 25936 5205 25976
rect 5163 25927 5205 25936
rect 20235 25976 20277 25985
rect 20235 25936 20236 25976
rect 20276 25936 20277 25976
rect 20235 25927 20277 25936
rect 2955 25892 2997 25901
rect 2955 25852 2956 25892
rect 2996 25852 2997 25892
rect 2955 25843 2997 25852
rect 6403 25892 6461 25893
rect 6403 25852 6412 25892
rect 6452 25852 6461 25892
rect 6403 25851 6461 25852
rect 12267 25892 12309 25901
rect 12267 25852 12268 25892
rect 12308 25852 12309 25892
rect 12267 25843 12309 25852
rect 15427 25892 15485 25893
rect 15427 25852 15436 25892
rect 15476 25852 15485 25892
rect 15427 25851 15485 25852
rect 17355 25892 17397 25901
rect 17355 25852 17356 25892
rect 17396 25852 17397 25892
rect 17355 25843 17397 25852
rect 19851 25892 19893 25901
rect 19851 25852 19852 25892
rect 19892 25852 19893 25892
rect 19851 25843 19893 25852
rect 1152 25724 20352 25748
rect 1152 25684 3688 25724
rect 3728 25684 3770 25724
rect 3810 25684 3852 25724
rect 3892 25684 3934 25724
rect 3974 25684 4016 25724
rect 4056 25684 18808 25724
rect 18848 25684 18890 25724
rect 18930 25684 18972 25724
rect 19012 25684 19054 25724
rect 19094 25684 19136 25724
rect 19176 25684 20352 25724
rect 1152 25660 20352 25684
rect 5835 25556 5877 25565
rect 5835 25516 5836 25556
rect 5876 25516 5877 25556
rect 5835 25507 5877 25516
rect 14091 25556 14133 25565
rect 14091 25516 14092 25556
rect 14132 25516 14133 25556
rect 14091 25507 14133 25516
rect 15531 25556 15573 25565
rect 15531 25516 15532 25556
rect 15572 25516 15573 25556
rect 15531 25507 15573 25516
rect 19555 25556 19613 25557
rect 19555 25516 19564 25556
rect 19604 25516 19613 25556
rect 19555 25515 19613 25516
rect 9579 25472 9621 25481
rect 9579 25432 9580 25472
rect 9620 25432 9621 25472
rect 9579 25423 9621 25432
rect 12259 25472 12317 25473
rect 12259 25432 12268 25472
rect 12308 25432 12317 25472
rect 12259 25431 12317 25432
rect 2763 25388 2805 25397
rect 2763 25348 2764 25388
rect 2804 25348 2805 25388
rect 2763 25339 2805 25348
rect 17355 25388 17397 25397
rect 17355 25348 17356 25388
rect 17396 25348 17397 25388
rect 17355 25339 17397 25348
rect 3819 25318 3861 25327
rect 2283 25304 2325 25313
rect 2283 25264 2284 25304
rect 2324 25264 2325 25304
rect 2283 25255 2325 25264
rect 2379 25304 2421 25313
rect 2379 25264 2380 25304
rect 2420 25264 2421 25304
rect 2379 25255 2421 25264
rect 2859 25304 2901 25313
rect 2859 25264 2860 25304
rect 2900 25264 2901 25304
rect 2859 25255 2901 25264
rect 3331 25304 3389 25305
rect 3331 25264 3340 25304
rect 3380 25264 3389 25304
rect 3819 25278 3820 25318
rect 3860 25278 3861 25318
rect 18411 25318 18453 25327
rect 3819 25269 3861 25278
rect 4387 25304 4445 25305
rect 3331 25263 3389 25264
rect 4387 25264 4396 25304
rect 4436 25264 4445 25304
rect 4387 25263 4445 25264
rect 5635 25304 5693 25305
rect 5635 25264 5644 25304
rect 5684 25264 5693 25304
rect 5635 25263 5693 25264
rect 6019 25304 6077 25305
rect 6019 25264 6028 25304
rect 6068 25264 6077 25304
rect 6019 25263 6077 25264
rect 7267 25304 7325 25305
rect 7267 25264 7276 25304
rect 7316 25264 7325 25304
rect 7267 25263 7325 25264
rect 7651 25304 7709 25305
rect 7651 25264 7660 25304
rect 7700 25264 7709 25304
rect 7651 25263 7709 25264
rect 8899 25304 8957 25305
rect 8899 25264 8908 25304
rect 8948 25264 8957 25304
rect 8899 25263 8957 25264
rect 9291 25304 9333 25313
rect 9291 25264 9292 25304
rect 9332 25264 9333 25304
rect 9291 25255 9333 25264
rect 9579 25304 9621 25313
rect 9579 25264 9580 25304
rect 9620 25264 9621 25304
rect 9579 25255 9621 25264
rect 9867 25304 9909 25313
rect 9867 25264 9868 25304
rect 9908 25264 9909 25304
rect 9867 25255 9909 25264
rect 10059 25304 10101 25313
rect 10059 25264 10060 25304
rect 10100 25264 10101 25304
rect 10059 25255 10101 25264
rect 10147 25304 10205 25305
rect 10147 25264 10156 25304
rect 10196 25264 10205 25304
rect 10147 25263 10205 25264
rect 10443 25304 10485 25313
rect 10443 25264 10444 25304
rect 10484 25264 10485 25304
rect 10443 25255 10485 25264
rect 10539 25304 10581 25313
rect 10539 25264 10540 25304
rect 10580 25264 10581 25304
rect 10539 25255 10581 25264
rect 10635 25304 10677 25313
rect 10635 25264 10636 25304
rect 10676 25264 10677 25304
rect 10635 25255 10677 25264
rect 11587 25304 11645 25305
rect 11587 25264 11596 25304
rect 11636 25264 11645 25304
rect 11587 25263 11645 25264
rect 11883 25304 11925 25313
rect 11883 25264 11884 25304
rect 11924 25264 11925 25304
rect 11883 25255 11925 25264
rect 11979 25304 12021 25313
rect 11979 25264 11980 25304
rect 12020 25264 12021 25304
rect 11979 25255 12021 25264
rect 13507 25304 13565 25305
rect 13507 25264 13516 25304
rect 13556 25264 13565 25304
rect 13507 25263 13565 25264
rect 13795 25304 13853 25305
rect 13795 25264 13804 25304
rect 13844 25264 13853 25304
rect 14091 25304 14133 25313
rect 13795 25263 13853 25264
rect 13899 25262 13941 25271
rect 4011 25220 4053 25229
rect 4011 25180 4012 25220
rect 4052 25180 4053 25220
rect 4011 25171 4053 25180
rect 13611 25220 13653 25229
rect 13611 25180 13612 25220
rect 13652 25180 13653 25220
rect 13899 25222 13900 25262
rect 13940 25222 13941 25262
rect 14091 25264 14092 25304
rect 14132 25264 14133 25304
rect 14091 25255 14133 25264
rect 14283 25304 14325 25313
rect 14283 25264 14284 25304
rect 14324 25264 14325 25304
rect 14283 25255 14325 25264
rect 14475 25304 14517 25313
rect 14475 25264 14476 25304
rect 14516 25264 14517 25304
rect 14475 25255 14517 25264
rect 14563 25304 14621 25305
rect 14563 25264 14572 25304
rect 14612 25264 14621 25304
rect 14563 25263 14621 25264
rect 14763 25304 14805 25313
rect 14763 25264 14764 25304
rect 14804 25264 14805 25304
rect 14763 25255 14805 25264
rect 14859 25304 14901 25313
rect 14859 25264 14860 25304
rect 14900 25264 14901 25304
rect 14859 25255 14901 25264
rect 14955 25304 14997 25313
rect 14955 25264 14956 25304
rect 14996 25264 14997 25304
rect 14955 25255 14997 25264
rect 15235 25304 15293 25305
rect 15235 25264 15244 25304
rect 15284 25264 15293 25304
rect 15235 25263 15293 25264
rect 15339 25304 15381 25313
rect 15339 25264 15340 25304
rect 15380 25264 15381 25304
rect 15339 25255 15381 25264
rect 15531 25304 15573 25313
rect 15531 25264 15532 25304
rect 15572 25264 15573 25304
rect 15531 25255 15573 25264
rect 16875 25304 16917 25313
rect 16875 25264 16876 25304
rect 16916 25264 16917 25304
rect 16875 25255 16917 25264
rect 16971 25304 17013 25313
rect 16971 25264 16972 25304
rect 17012 25264 17013 25304
rect 16971 25255 17013 25264
rect 17451 25304 17493 25313
rect 17451 25264 17452 25304
rect 17492 25264 17493 25304
rect 17451 25255 17493 25264
rect 17923 25304 17981 25305
rect 17923 25264 17932 25304
rect 17972 25264 17981 25304
rect 18411 25278 18412 25318
rect 18452 25278 18453 25318
rect 18411 25269 18453 25278
rect 18883 25304 18941 25305
rect 17923 25263 17981 25264
rect 18883 25264 18892 25304
rect 18932 25264 18941 25304
rect 18883 25263 18941 25264
rect 19179 25304 19221 25313
rect 19179 25264 19180 25304
rect 19220 25264 19221 25304
rect 19179 25255 19221 25264
rect 19275 25304 19317 25313
rect 19275 25264 19276 25304
rect 19316 25264 19317 25304
rect 19275 25255 19317 25264
rect 19755 25304 19797 25313
rect 19755 25264 19756 25304
rect 19796 25264 19797 25304
rect 19755 25255 19797 25264
rect 19851 25304 19893 25313
rect 19851 25264 19852 25304
rect 19892 25264 19893 25304
rect 19851 25255 19893 25264
rect 13899 25213 13941 25222
rect 14379 25220 14421 25229
rect 13611 25171 13653 25180
rect 14379 25180 14380 25220
rect 14420 25180 14421 25220
rect 14379 25171 14421 25180
rect 15051 25220 15093 25229
rect 15051 25180 15052 25220
rect 15092 25180 15093 25220
rect 15051 25171 15093 25180
rect 18603 25220 18645 25229
rect 18603 25180 18604 25220
rect 18644 25180 18645 25220
rect 18603 25171 18645 25180
rect 7467 25136 7509 25145
rect 7467 25096 7468 25136
rect 7508 25096 7509 25136
rect 7467 25087 7509 25096
rect 9099 25136 9141 25145
rect 9099 25096 9100 25136
rect 9140 25096 9141 25136
rect 9099 25087 9141 25096
rect 9955 25136 10013 25137
rect 9955 25096 9964 25136
rect 10004 25096 10013 25136
rect 9955 25095 10013 25096
rect 10827 25136 10869 25145
rect 10827 25096 10828 25136
rect 10868 25096 10869 25136
rect 10827 25087 10869 25096
rect 20035 25136 20093 25137
rect 20035 25096 20044 25136
rect 20084 25096 20093 25136
rect 20035 25095 20093 25096
rect 1152 24968 20452 24992
rect 1152 24928 4928 24968
rect 4968 24928 5010 24968
rect 5050 24928 5092 24968
rect 5132 24928 5174 24968
rect 5214 24928 5256 24968
rect 5296 24928 20048 24968
rect 20088 24928 20130 24968
rect 20170 24928 20212 24968
rect 20252 24928 20294 24968
rect 20334 24928 20376 24968
rect 20416 24928 20452 24968
rect 1152 24904 20452 24928
rect 18507 24842 18549 24851
rect 14379 24800 14421 24809
rect 14379 24760 14380 24800
rect 14420 24760 14421 24800
rect 14379 24751 14421 24760
rect 18027 24800 18069 24809
rect 18027 24760 18028 24800
rect 18068 24760 18069 24800
rect 18507 24802 18508 24842
rect 18548 24802 18549 24842
rect 18507 24793 18549 24802
rect 20235 24800 20277 24809
rect 18027 24751 18069 24760
rect 20235 24760 20236 24800
rect 20276 24760 20277 24800
rect 20235 24751 20277 24760
rect 10731 24716 10773 24725
rect 10731 24676 10732 24716
rect 10772 24676 10773 24716
rect 10731 24667 10773 24676
rect 15627 24716 15669 24725
rect 15627 24676 15628 24716
rect 15668 24676 15669 24716
rect 15627 24667 15669 24676
rect 11019 24653 11061 24662
rect 3331 24632 3389 24633
rect 3331 24592 3340 24632
rect 3380 24592 3389 24632
rect 3331 24591 3389 24592
rect 3435 24632 3477 24641
rect 3435 24592 3436 24632
rect 3476 24592 3477 24632
rect 3435 24583 3477 24592
rect 3627 24632 3669 24641
rect 3627 24592 3628 24632
rect 3668 24592 3669 24632
rect 3627 24583 3669 24592
rect 4771 24632 4829 24633
rect 4771 24592 4780 24632
rect 4820 24592 4829 24632
rect 4771 24591 4829 24592
rect 6019 24632 6077 24633
rect 6019 24592 6028 24632
rect 6068 24592 6077 24632
rect 6019 24591 6077 24592
rect 6603 24632 6645 24641
rect 6603 24592 6604 24632
rect 6644 24592 6645 24632
rect 6603 24583 6645 24592
rect 6699 24632 6741 24641
rect 6699 24592 6700 24632
rect 6740 24592 6741 24632
rect 6699 24583 6741 24592
rect 6795 24632 6837 24641
rect 6795 24592 6796 24632
rect 6836 24592 6837 24632
rect 6795 24583 6837 24592
rect 7651 24632 7709 24633
rect 7651 24592 7660 24632
rect 7700 24592 7709 24632
rect 7651 24591 7709 24592
rect 7947 24632 7989 24641
rect 7947 24592 7948 24632
rect 7988 24592 7989 24632
rect 7947 24583 7989 24592
rect 8043 24632 8085 24641
rect 8043 24592 8044 24632
rect 8084 24592 8085 24632
rect 8043 24583 8085 24592
rect 9003 24632 9045 24641
rect 9003 24592 9004 24632
rect 9044 24592 9045 24632
rect 9003 24583 9045 24592
rect 9099 24632 9141 24641
rect 9099 24592 9100 24632
rect 9140 24592 9141 24632
rect 9099 24583 9141 24592
rect 10051 24632 10109 24633
rect 10051 24592 10060 24632
rect 10100 24592 10109 24632
rect 10051 24591 10109 24592
rect 10539 24622 10581 24631
rect 10539 24582 10540 24622
rect 10580 24582 10581 24622
rect 11019 24613 11020 24653
rect 11060 24613 11061 24653
rect 11019 24604 11061 24613
rect 11115 24632 11157 24641
rect 10539 24573 10581 24582
rect 10923 24587 10965 24596
rect 9483 24548 9525 24557
rect 9483 24508 9484 24548
rect 9524 24508 9525 24548
rect 9483 24499 9525 24508
rect 9579 24548 9621 24557
rect 9579 24508 9580 24548
rect 9620 24508 9621 24548
rect 10923 24547 10924 24587
rect 10964 24547 10965 24587
rect 11115 24592 11116 24632
rect 11156 24592 11157 24632
rect 11115 24583 11157 24592
rect 11211 24632 11253 24641
rect 11211 24592 11212 24632
rect 11252 24592 11253 24632
rect 11211 24583 11253 24592
rect 11491 24632 11549 24633
rect 11491 24592 11500 24632
rect 11540 24592 11549 24632
rect 11491 24591 11549 24592
rect 11787 24632 11829 24641
rect 11787 24592 11788 24632
rect 11828 24592 11829 24632
rect 11787 24583 11829 24592
rect 11883 24632 11925 24641
rect 11883 24592 11884 24632
rect 11924 24592 11925 24632
rect 11883 24583 11925 24592
rect 12643 24632 12701 24633
rect 12643 24592 12652 24632
rect 12692 24592 12701 24632
rect 12643 24591 12701 24592
rect 13891 24632 13949 24633
rect 13891 24592 13900 24632
rect 13940 24592 13949 24632
rect 13891 24591 13949 24592
rect 14283 24632 14325 24641
rect 14283 24592 14284 24632
rect 14324 24592 14325 24632
rect 14283 24583 14325 24592
rect 14571 24632 14613 24641
rect 14571 24592 14572 24632
rect 14612 24592 14613 24632
rect 14955 24632 14997 24641
rect 14571 24583 14613 24592
rect 14763 24619 14805 24628
rect 14763 24579 14764 24619
rect 14804 24579 14805 24619
rect 14955 24592 14956 24632
rect 14996 24592 14997 24632
rect 14955 24583 14997 24592
rect 15235 24632 15293 24633
rect 15235 24592 15244 24632
rect 15284 24592 15293 24632
rect 15235 24591 15293 24592
rect 15531 24632 15573 24641
rect 15531 24592 15532 24632
rect 15572 24592 15573 24632
rect 15531 24583 15573 24592
rect 16579 24632 16637 24633
rect 16579 24592 16588 24632
rect 16628 24592 16637 24632
rect 16579 24591 16637 24592
rect 17827 24632 17885 24633
rect 17827 24592 17836 24632
rect 17876 24592 17885 24632
rect 17827 24591 17885 24592
rect 18699 24632 18741 24641
rect 18699 24592 18700 24632
rect 18740 24592 18741 24632
rect 18699 24583 18741 24592
rect 18795 24632 18837 24641
rect 18795 24592 18796 24632
rect 18836 24592 18837 24632
rect 18795 24583 18837 24592
rect 19179 24632 19221 24641
rect 19179 24592 19180 24632
rect 19220 24592 19221 24632
rect 19179 24583 19221 24592
rect 19275 24632 19317 24641
rect 19275 24592 19276 24632
rect 19316 24592 19317 24632
rect 19275 24583 19317 24592
rect 19371 24632 19413 24641
rect 19371 24592 19372 24632
rect 19412 24592 19413 24632
rect 19371 24583 19413 24592
rect 19467 24632 19509 24641
rect 19467 24592 19468 24632
rect 19508 24592 19509 24632
rect 19467 24583 19509 24592
rect 14763 24570 14805 24579
rect 10923 24538 10965 24547
rect 14859 24548 14901 24557
rect 9579 24499 9621 24508
rect 14859 24508 14860 24548
rect 14900 24508 14901 24548
rect 14859 24499 14901 24508
rect 19651 24548 19709 24549
rect 19651 24508 19660 24548
rect 19700 24508 19709 24548
rect 19651 24507 19709 24508
rect 20035 24548 20093 24549
rect 20035 24508 20044 24548
rect 20084 24508 20093 24548
rect 20035 24507 20093 24508
rect 6219 24464 6261 24473
rect 6219 24424 6220 24464
rect 6260 24424 6261 24464
rect 6219 24415 6261 24424
rect 18987 24464 19029 24473
rect 18987 24424 18988 24464
rect 19028 24424 19029 24464
rect 18987 24415 19029 24424
rect 19851 24464 19893 24473
rect 19851 24424 19852 24464
rect 19892 24424 19893 24464
rect 19851 24415 19893 24424
rect 3627 24380 3669 24389
rect 3627 24340 3628 24380
rect 3668 24340 3669 24380
rect 3627 24331 3669 24340
rect 6979 24380 7037 24381
rect 6979 24340 6988 24380
rect 7028 24340 7037 24380
rect 6979 24339 7037 24340
rect 8323 24380 8381 24381
rect 8323 24340 8332 24380
rect 8372 24340 8381 24380
rect 8323 24339 8381 24340
rect 12163 24380 12221 24381
rect 12163 24340 12172 24380
rect 12212 24340 12221 24380
rect 12163 24339 12221 24340
rect 14091 24380 14133 24389
rect 14091 24340 14092 24380
rect 14132 24340 14133 24380
rect 14091 24331 14133 24340
rect 15907 24380 15965 24381
rect 15907 24340 15916 24380
rect 15956 24340 15965 24380
rect 15907 24339 15965 24340
rect 1152 24212 20352 24236
rect 1152 24172 3688 24212
rect 3728 24172 3770 24212
rect 3810 24172 3852 24212
rect 3892 24172 3934 24212
rect 3974 24172 4016 24212
rect 4056 24172 18808 24212
rect 18848 24172 18890 24212
rect 18930 24172 18972 24212
rect 19012 24172 19054 24212
rect 19094 24172 19136 24212
rect 19176 24172 20352 24212
rect 1152 24148 20352 24172
rect 10827 24044 10869 24053
rect 10827 24004 10828 24044
rect 10868 24004 10869 24044
rect 10827 23995 10869 24004
rect 5259 23960 5301 23969
rect 5259 23920 5260 23960
rect 5300 23920 5301 23960
rect 5259 23911 5301 23920
rect 12843 23960 12885 23969
rect 12843 23920 12844 23960
rect 12884 23920 12885 23960
rect 12843 23911 12885 23920
rect 15043 23960 15101 23961
rect 15043 23920 15052 23960
rect 15092 23920 15101 23960
rect 15043 23919 15101 23920
rect 19267 23960 19325 23961
rect 19267 23920 19276 23960
rect 19316 23920 19325 23960
rect 19267 23919 19325 23920
rect 6507 23876 6549 23885
rect 6507 23836 6508 23876
rect 6548 23836 6549 23876
rect 6507 23827 6549 23836
rect 13707 23876 13749 23885
rect 13707 23836 13708 23876
rect 13748 23836 13749 23876
rect 13707 23827 13749 23836
rect 19939 23876 19997 23877
rect 19939 23836 19948 23876
rect 19988 23836 19997 23876
rect 19939 23835 19997 23836
rect 1219 23792 1277 23793
rect 1219 23752 1228 23792
rect 1268 23752 1277 23792
rect 1219 23751 1277 23752
rect 2467 23792 2525 23793
rect 2467 23752 2476 23792
rect 2516 23752 2525 23792
rect 2467 23751 2525 23752
rect 3051 23792 3093 23801
rect 3051 23752 3052 23792
rect 3092 23752 3093 23792
rect 3051 23743 3093 23752
rect 3147 23792 3189 23801
rect 3147 23752 3148 23792
rect 3188 23752 3189 23792
rect 3147 23743 3189 23752
rect 3531 23792 3573 23801
rect 3531 23752 3532 23792
rect 3572 23752 3573 23792
rect 3531 23743 3573 23752
rect 3627 23792 3669 23801
rect 4587 23797 4629 23806
rect 3627 23752 3628 23792
rect 3668 23752 3669 23792
rect 3627 23743 3669 23752
rect 4099 23792 4157 23793
rect 4099 23752 4108 23792
rect 4148 23752 4157 23792
rect 4099 23751 4157 23752
rect 4587 23757 4588 23797
rect 4628 23757 4629 23797
rect 4587 23748 4629 23757
rect 4971 23792 5013 23801
rect 4971 23752 4972 23792
rect 5012 23752 5013 23792
rect 4971 23743 5013 23752
rect 5259 23792 5301 23801
rect 5259 23752 5260 23792
rect 5300 23752 5301 23792
rect 5259 23743 5301 23752
rect 5451 23792 5493 23801
rect 5451 23752 5452 23792
rect 5492 23752 5493 23792
rect 5451 23743 5493 23752
rect 5643 23792 5685 23801
rect 5643 23752 5644 23792
rect 5684 23752 5685 23792
rect 5643 23743 5685 23752
rect 5731 23792 5789 23793
rect 5731 23752 5740 23792
rect 5780 23752 5789 23792
rect 5731 23751 5789 23752
rect 6027 23792 6069 23801
rect 6027 23752 6028 23792
rect 6068 23752 6069 23792
rect 6027 23743 6069 23752
rect 6123 23792 6165 23801
rect 6123 23752 6124 23792
rect 6164 23752 6165 23792
rect 6123 23743 6165 23752
rect 6603 23792 6645 23801
rect 7563 23797 7605 23806
rect 6603 23752 6604 23792
rect 6644 23752 6645 23792
rect 6603 23743 6645 23752
rect 7075 23792 7133 23793
rect 7075 23752 7084 23792
rect 7124 23752 7133 23792
rect 7075 23751 7133 23752
rect 7563 23757 7564 23797
rect 7604 23757 7605 23797
rect 7563 23748 7605 23757
rect 7947 23792 7989 23801
rect 7947 23752 7948 23792
rect 7988 23752 7989 23792
rect 7947 23743 7989 23752
rect 8043 23792 8085 23801
rect 8043 23752 8044 23792
rect 8084 23752 8085 23792
rect 8043 23743 8085 23752
rect 8139 23792 8181 23801
rect 8139 23752 8140 23792
rect 8180 23752 8181 23792
rect 8139 23743 8181 23752
rect 8235 23792 8277 23801
rect 8235 23752 8236 23792
rect 8276 23752 8277 23792
rect 8235 23743 8277 23752
rect 9379 23792 9437 23793
rect 9379 23752 9388 23792
rect 9428 23752 9437 23792
rect 9379 23751 9437 23752
rect 10627 23792 10685 23793
rect 10627 23752 10636 23792
rect 10676 23752 10685 23792
rect 10627 23751 10685 23752
rect 11395 23792 11453 23793
rect 11395 23752 11404 23792
rect 11444 23752 11453 23792
rect 11395 23751 11453 23752
rect 12643 23792 12701 23793
rect 12643 23752 12652 23792
rect 12692 23752 12701 23792
rect 12643 23751 12701 23752
rect 13131 23792 13173 23801
rect 13131 23752 13132 23792
rect 13172 23752 13173 23792
rect 13131 23743 13173 23752
rect 13227 23792 13269 23801
rect 13227 23752 13228 23792
rect 13268 23752 13269 23792
rect 13227 23743 13269 23752
rect 13611 23792 13653 23801
rect 14667 23797 14709 23806
rect 13611 23752 13612 23792
rect 13652 23752 13653 23792
rect 13611 23743 13653 23752
rect 14179 23792 14237 23793
rect 14179 23752 14188 23792
rect 14228 23752 14237 23792
rect 14179 23751 14237 23752
rect 14667 23757 14668 23797
rect 14708 23757 14709 23797
rect 14667 23748 14709 23757
rect 15243 23792 15285 23801
rect 15243 23752 15244 23792
rect 15284 23752 15285 23792
rect 15243 23743 15285 23752
rect 15339 23792 15381 23801
rect 15339 23752 15340 23792
rect 15380 23752 15381 23792
rect 15339 23743 15381 23752
rect 15435 23792 15477 23801
rect 15435 23752 15436 23792
rect 15476 23752 15477 23792
rect 15435 23743 15477 23752
rect 15715 23792 15773 23793
rect 15715 23752 15724 23792
rect 15764 23752 15773 23792
rect 15715 23751 15773 23752
rect 16963 23792 17021 23793
rect 16963 23752 16972 23792
rect 17012 23752 17021 23792
rect 16963 23751 17021 23752
rect 17355 23792 17397 23801
rect 17355 23752 17356 23792
rect 17396 23752 17397 23792
rect 17355 23743 17397 23752
rect 17451 23792 17493 23801
rect 17451 23752 17452 23792
rect 17492 23752 17493 23792
rect 17451 23743 17493 23752
rect 17547 23792 17589 23801
rect 17547 23752 17548 23792
rect 17588 23752 17589 23792
rect 17547 23743 17589 23752
rect 18315 23792 18357 23801
rect 18315 23752 18316 23792
rect 18356 23752 18357 23792
rect 18315 23743 18357 23752
rect 18507 23792 18549 23801
rect 18507 23752 18508 23792
rect 18548 23752 18549 23792
rect 18507 23743 18549 23752
rect 18595 23792 18653 23793
rect 18595 23752 18604 23792
rect 18644 23752 18653 23792
rect 18595 23751 18653 23752
rect 18891 23792 18933 23801
rect 18891 23752 18892 23792
rect 18932 23752 18933 23792
rect 18891 23743 18933 23752
rect 18987 23792 19029 23801
rect 18987 23752 18988 23792
rect 19028 23752 19029 23792
rect 18987 23743 19029 23752
rect 19083 23792 19125 23801
rect 19083 23752 19084 23792
rect 19124 23752 19125 23792
rect 19083 23743 19125 23752
rect 19467 23792 19509 23801
rect 19467 23752 19468 23792
rect 19508 23752 19509 23792
rect 19467 23743 19509 23752
rect 19563 23792 19605 23801
rect 19563 23752 19564 23792
rect 19604 23752 19605 23792
rect 19563 23743 19605 23752
rect 19659 23792 19701 23801
rect 19659 23752 19660 23792
rect 19700 23752 19701 23792
rect 19659 23743 19701 23752
rect 4779 23708 4821 23717
rect 4779 23668 4780 23708
rect 4820 23668 4821 23708
rect 4779 23659 4821 23668
rect 5547 23708 5589 23717
rect 5547 23668 5548 23708
rect 5588 23668 5589 23708
rect 5547 23659 5589 23668
rect 7755 23708 7797 23717
rect 7755 23668 7756 23708
rect 7796 23668 7797 23708
rect 7755 23659 7797 23668
rect 14859 23708 14901 23717
rect 14859 23668 14860 23708
rect 14900 23668 14901 23708
rect 14859 23659 14901 23668
rect 18411 23708 18453 23717
rect 18411 23668 18412 23708
rect 18452 23668 18453 23708
rect 18411 23659 18453 23668
rect 2667 23624 2709 23633
rect 2667 23584 2668 23624
rect 2708 23584 2709 23624
rect 2667 23575 2709 23584
rect 17163 23624 17205 23633
rect 17163 23584 17164 23624
rect 17204 23584 17205 23624
rect 17163 23575 17205 23584
rect 17635 23624 17693 23625
rect 17635 23584 17644 23624
rect 17684 23584 17693 23624
rect 17635 23583 17693 23584
rect 19747 23624 19805 23625
rect 19747 23584 19756 23624
rect 19796 23584 19805 23624
rect 19747 23583 19805 23584
rect 20139 23624 20181 23633
rect 20139 23584 20140 23624
rect 20180 23584 20181 23624
rect 20139 23575 20181 23584
rect 1152 23456 20452 23480
rect 1152 23416 4928 23456
rect 4968 23416 5010 23456
rect 5050 23416 5092 23456
rect 5132 23416 5174 23456
rect 5214 23416 5256 23456
rect 5296 23416 20048 23456
rect 20088 23416 20130 23456
rect 20170 23416 20212 23456
rect 20252 23416 20294 23456
rect 20334 23416 20376 23456
rect 20416 23416 20452 23456
rect 1152 23392 20452 23416
rect 2667 23288 2709 23297
rect 2667 23248 2668 23288
rect 2708 23248 2709 23288
rect 2667 23239 2709 23248
rect 4491 23288 4533 23297
rect 4491 23248 4492 23288
rect 4532 23248 4533 23288
rect 4491 23239 4533 23248
rect 6411 23288 6453 23297
rect 6411 23248 6412 23288
rect 6452 23248 6453 23288
rect 6411 23239 6453 23248
rect 12075 23288 12117 23297
rect 12075 23248 12076 23288
rect 12116 23248 12117 23288
rect 12075 23239 12117 23248
rect 15339 23288 15381 23297
rect 15339 23248 15340 23288
rect 15380 23248 15381 23288
rect 15339 23239 15381 23248
rect 17347 23288 17405 23289
rect 17347 23248 17356 23288
rect 17396 23248 17405 23288
rect 17347 23247 17405 23248
rect 18115 23288 18173 23289
rect 18115 23248 18124 23288
rect 18164 23248 18173 23288
rect 18115 23247 18173 23248
rect 18411 23288 18453 23297
rect 18411 23248 18412 23288
rect 18452 23248 18453 23288
rect 18411 23239 18453 23248
rect 9963 23132 10005 23141
rect 1219 23120 1277 23121
rect 1219 23080 1228 23120
rect 1268 23080 1277 23120
rect 1219 23079 1277 23080
rect 2467 23120 2525 23121
rect 2467 23080 2476 23120
rect 2516 23080 2525 23120
rect 2467 23079 2525 23080
rect 3043 23120 3101 23121
rect 3043 23080 3052 23120
rect 3092 23080 3101 23120
rect 3043 23079 3101 23080
rect 4291 23120 4349 23121
rect 4291 23080 4300 23120
rect 4340 23080 4349 23120
rect 4291 23079 4349 23080
rect 4675 23120 4733 23121
rect 4675 23080 4684 23120
rect 4724 23080 4733 23120
rect 4675 23079 4733 23080
rect 4963 23120 5021 23121
rect 4963 23080 4972 23120
rect 5012 23080 5021 23120
rect 4963 23079 5021 23080
rect 6211 23120 6269 23121
rect 6211 23080 6220 23120
rect 6260 23080 6269 23120
rect 6211 23079 6269 23080
rect 6603 23120 6645 23129
rect 6603 23080 6604 23120
rect 6644 23080 6645 23120
rect 6603 23071 6645 23080
rect 6699 23120 6741 23129
rect 6699 23080 6700 23120
rect 6740 23080 6741 23120
rect 6699 23071 6741 23080
rect 6795 23120 6837 23129
rect 6795 23080 6796 23120
rect 6836 23080 6837 23120
rect 6795 23071 6837 23080
rect 6891 23120 6933 23129
rect 6891 23080 6892 23120
rect 6932 23080 6933 23120
rect 6891 23071 6933 23080
rect 7179 23120 7221 23129
rect 7179 23080 7180 23120
rect 7220 23080 7221 23120
rect 7179 23071 7221 23080
rect 7467 23120 7509 23129
rect 7467 23080 7468 23120
rect 7508 23080 7509 23120
rect 7467 23071 7509 23080
rect 7659 23120 7701 23129
rect 7659 23080 7660 23120
rect 7700 23080 7701 23120
rect 7659 23071 7701 23080
rect 7851 23120 7893 23129
rect 7851 23080 7852 23120
rect 7892 23080 7893 23120
rect 7851 23071 7893 23080
rect 7939 23120 7997 23121
rect 7939 23080 7948 23120
rect 7988 23080 7997 23120
rect 7939 23079 7997 23080
rect 8131 23120 8189 23121
rect 8131 23080 8140 23120
rect 8180 23080 8189 23120
rect 8131 23079 8189 23080
rect 9379 23120 9437 23121
rect 9379 23080 9388 23120
rect 9428 23080 9437 23120
rect 9963 23092 9964 23132
rect 10004 23092 10005 23132
rect 9963 23083 10005 23092
rect 10059 23120 10101 23129
rect 9379 23079 9437 23080
rect 10059 23080 10060 23120
rect 10100 23080 10101 23120
rect 10059 23071 10101 23080
rect 10155 23120 10197 23129
rect 10155 23080 10156 23120
rect 10196 23080 10197 23120
rect 10155 23071 10197 23080
rect 10627 23120 10685 23121
rect 10627 23080 10636 23120
rect 10676 23080 10685 23120
rect 10627 23079 10685 23080
rect 11875 23120 11933 23121
rect 11875 23080 11884 23120
rect 11924 23080 11933 23120
rect 11875 23079 11933 23080
rect 13891 23120 13949 23121
rect 13891 23080 13900 23120
rect 13940 23080 13949 23120
rect 15715 23120 15773 23121
rect 13891 23079 13949 23080
rect 15139 23099 15197 23100
rect 15139 23059 15148 23099
rect 15188 23059 15197 23099
rect 15715 23080 15724 23120
rect 15764 23080 15773 23120
rect 15715 23079 15773 23080
rect 16963 23120 17021 23121
rect 16963 23080 16972 23120
rect 17012 23080 17021 23120
rect 16963 23079 17021 23080
rect 17547 23120 17589 23129
rect 17547 23080 17548 23120
rect 17588 23080 17589 23120
rect 17547 23071 17589 23080
rect 17643 23120 17685 23129
rect 17643 23080 17644 23120
rect 17684 23080 17685 23120
rect 17643 23071 17685 23080
rect 17835 23120 17877 23129
rect 17835 23080 17836 23120
rect 17876 23080 17877 23120
rect 17835 23071 17877 23080
rect 17931 23120 17973 23129
rect 17931 23080 17932 23120
rect 17972 23080 17973 23120
rect 17931 23071 17973 23080
rect 18027 23120 18069 23129
rect 18027 23080 18028 23120
rect 18068 23080 18069 23120
rect 19843 23120 19901 23121
rect 18027 23071 18069 23080
rect 18595 23099 18653 23100
rect 15139 23058 15197 23059
rect 18595 23059 18604 23099
rect 18644 23059 18653 23099
rect 19843 23080 19852 23120
rect 19892 23080 19901 23120
rect 19843 23079 19901 23080
rect 18595 23058 18653 23059
rect 7467 22952 7509 22961
rect 7467 22912 7468 22952
rect 7508 22912 7509 22952
rect 7467 22903 7509 22912
rect 17163 22952 17205 22961
rect 17163 22912 17164 22952
rect 17204 22912 17205 22952
rect 17163 22903 17205 22912
rect 4779 22868 4821 22877
rect 4779 22828 4780 22868
rect 4820 22828 4821 22868
rect 4779 22819 4821 22828
rect 7659 22868 7701 22877
rect 7659 22828 7660 22868
rect 7700 22828 7701 22868
rect 7659 22819 7701 22828
rect 9579 22868 9621 22877
rect 9579 22828 9580 22868
rect 9620 22828 9621 22868
rect 9579 22819 9621 22828
rect 9763 22868 9821 22869
rect 9763 22828 9772 22868
rect 9812 22828 9821 22868
rect 9763 22827 9821 22828
rect 1152 22700 20352 22724
rect 1152 22660 3688 22700
rect 3728 22660 3770 22700
rect 3810 22660 3852 22700
rect 3892 22660 3934 22700
rect 3974 22660 4016 22700
rect 4056 22660 18808 22700
rect 18848 22660 18890 22700
rect 18930 22660 18972 22700
rect 19012 22660 19054 22700
rect 19094 22660 19136 22700
rect 19176 22660 20352 22700
rect 1152 22636 20352 22660
rect 3139 22532 3197 22533
rect 3139 22492 3148 22532
rect 3188 22492 3197 22532
rect 3139 22491 3197 22492
rect 3331 22448 3389 22449
rect 3331 22408 3340 22448
rect 3380 22408 3389 22448
rect 3331 22407 3389 22408
rect 4299 22448 4341 22457
rect 4299 22408 4300 22448
rect 4340 22408 4341 22448
rect 4299 22399 4341 22408
rect 6507 22448 6549 22457
rect 6507 22408 6508 22448
rect 6548 22408 6549 22448
rect 6507 22399 6549 22408
rect 7459 22448 7517 22449
rect 7459 22408 7468 22448
rect 7508 22408 7517 22448
rect 7459 22407 7517 22408
rect 12355 22448 12413 22449
rect 12355 22408 12364 22448
rect 12404 22408 12413 22448
rect 12355 22407 12413 22408
rect 19843 22448 19901 22449
rect 19843 22408 19852 22448
rect 19892 22408 19901 22448
rect 19843 22407 19901 22408
rect 8523 22364 8565 22373
rect 8523 22324 8524 22364
rect 8564 22324 8565 22364
rect 8523 22315 8565 22324
rect 13707 22364 13749 22373
rect 13707 22324 13708 22364
rect 13748 22324 13749 22364
rect 13707 22315 13749 22324
rect 18699 22294 18741 22303
rect 2467 22280 2525 22281
rect 2467 22240 2476 22280
rect 2516 22240 2525 22280
rect 2467 22239 2525 22240
rect 2763 22280 2805 22289
rect 2763 22240 2764 22280
rect 2804 22240 2805 22280
rect 2763 22231 2805 22240
rect 2859 22280 2901 22289
rect 2859 22240 2860 22280
rect 2900 22240 2901 22280
rect 2859 22231 2901 22240
rect 3723 22280 3765 22289
rect 3723 22240 3724 22280
rect 3764 22240 3765 22280
rect 3723 22231 3765 22240
rect 4003 22280 4061 22281
rect 4003 22240 4012 22280
rect 4052 22240 4061 22280
rect 4003 22239 4061 22240
rect 4587 22280 4629 22289
rect 4587 22240 4588 22280
rect 4628 22240 4629 22280
rect 4587 22231 4629 22240
rect 4675 22280 4733 22281
rect 4675 22240 4684 22280
rect 4724 22240 4733 22280
rect 4675 22239 4733 22240
rect 5059 22280 5117 22281
rect 5059 22240 5068 22280
rect 5108 22240 5117 22280
rect 5059 22239 5117 22240
rect 6307 22280 6365 22281
rect 6307 22240 6316 22280
rect 6356 22240 6365 22280
rect 6307 22239 6365 22240
rect 6787 22280 6845 22281
rect 6787 22240 6796 22280
rect 6836 22240 6845 22280
rect 6787 22239 6845 22240
rect 7083 22280 7125 22289
rect 7083 22240 7084 22280
rect 7124 22240 7125 22280
rect 7083 22231 7125 22240
rect 8043 22280 8085 22289
rect 8043 22240 8044 22280
rect 8084 22240 8085 22280
rect 8043 22231 8085 22240
rect 8139 22280 8181 22289
rect 8139 22240 8140 22280
rect 8180 22240 8181 22280
rect 8139 22231 8181 22240
rect 8619 22280 8661 22289
rect 9579 22285 9621 22294
rect 8619 22240 8620 22280
rect 8660 22240 8661 22280
rect 8619 22231 8661 22240
rect 9091 22280 9149 22281
rect 9091 22240 9100 22280
rect 9140 22240 9149 22280
rect 9091 22239 9149 22240
rect 9579 22245 9580 22285
rect 9620 22245 9621 22285
rect 9579 22236 9621 22245
rect 9955 22280 10013 22281
rect 9955 22240 9964 22280
rect 10004 22240 10013 22280
rect 9955 22239 10013 22240
rect 11203 22280 11261 22281
rect 11203 22240 11212 22280
rect 11252 22240 11261 22280
rect 11203 22239 11261 22240
rect 11683 22280 11741 22281
rect 11683 22240 11692 22280
rect 11732 22240 11741 22280
rect 11683 22239 11741 22240
rect 11979 22280 12021 22289
rect 11979 22240 11980 22280
rect 12020 22240 12021 22280
rect 11979 22231 12021 22240
rect 13227 22280 13269 22289
rect 13227 22240 13228 22280
rect 13268 22240 13269 22280
rect 13227 22231 13269 22240
rect 13323 22280 13365 22289
rect 13323 22240 13324 22280
rect 13364 22240 13365 22280
rect 13323 22231 13365 22240
rect 13803 22280 13845 22289
rect 14763 22285 14805 22294
rect 13803 22240 13804 22280
rect 13844 22240 13845 22280
rect 13803 22231 13845 22240
rect 14275 22280 14333 22281
rect 14275 22240 14284 22280
rect 14324 22240 14333 22280
rect 14275 22239 14333 22240
rect 14763 22245 14764 22285
rect 14804 22245 14805 22285
rect 14763 22236 14805 22245
rect 15243 22280 15285 22289
rect 15243 22240 15244 22280
rect 15284 22240 15285 22280
rect 15243 22231 15285 22240
rect 15339 22280 15381 22289
rect 15339 22240 15340 22280
rect 15380 22240 15381 22280
rect 15339 22231 15381 22240
rect 15435 22280 15477 22289
rect 15435 22240 15436 22280
rect 15476 22240 15477 22280
rect 15435 22231 15477 22240
rect 15819 22280 15861 22289
rect 15819 22240 15820 22280
rect 15860 22240 15861 22280
rect 15819 22231 15861 22240
rect 15915 22280 15957 22289
rect 15915 22240 15916 22280
rect 15956 22240 15957 22280
rect 15915 22231 15957 22240
rect 16011 22280 16053 22289
rect 16011 22240 16012 22280
rect 16052 22240 16053 22280
rect 16011 22231 16053 22240
rect 17163 22280 17205 22289
rect 17163 22240 17164 22280
rect 17204 22240 17205 22280
rect 17163 22231 17205 22240
rect 17259 22280 17301 22289
rect 17259 22240 17260 22280
rect 17300 22240 17301 22280
rect 17259 22231 17301 22240
rect 17643 22280 17685 22289
rect 17643 22240 17644 22280
rect 17684 22240 17685 22280
rect 17643 22231 17685 22240
rect 17739 22280 17781 22289
rect 17739 22240 17740 22280
rect 17780 22240 17781 22280
rect 17739 22231 17781 22240
rect 18211 22280 18269 22281
rect 18211 22240 18220 22280
rect 18260 22240 18269 22280
rect 18699 22254 18700 22294
rect 18740 22254 18741 22294
rect 18699 22245 18741 22254
rect 19171 22280 19229 22281
rect 18211 22239 18269 22240
rect 19171 22240 19180 22280
rect 19220 22240 19229 22280
rect 19171 22239 19229 22240
rect 19467 22280 19509 22289
rect 19467 22240 19468 22280
rect 19508 22240 19509 22280
rect 19467 22231 19509 22240
rect 19563 22280 19605 22289
rect 19563 22240 19564 22280
rect 19604 22240 19605 22280
rect 19563 22231 19605 22240
rect 3627 22196 3669 22205
rect 3627 22156 3628 22196
rect 3668 22156 3669 22196
rect 3627 22147 3669 22156
rect 7179 22196 7221 22205
rect 7179 22156 7180 22196
rect 7220 22156 7221 22196
rect 7179 22147 7221 22156
rect 11403 22196 11445 22205
rect 11403 22156 11404 22196
rect 11444 22156 11445 22196
rect 11403 22147 11445 22156
rect 12075 22196 12117 22205
rect 12075 22156 12076 22196
rect 12116 22156 12117 22196
rect 12075 22147 12117 22156
rect 18891 22196 18933 22205
rect 18891 22156 18892 22196
rect 18932 22156 18933 22196
rect 18891 22147 18933 22156
rect 14955 22112 14997 22121
rect 9771 22070 9813 22079
rect 4779 22054 4821 22063
rect 4779 22014 4780 22054
rect 4820 22014 4821 22054
rect 9771 22030 9772 22070
rect 9812 22030 9813 22070
rect 14955 22072 14956 22112
rect 14996 22072 14997 22112
rect 14955 22063 14997 22072
rect 15627 22112 15669 22121
rect 15627 22072 15628 22112
rect 15668 22072 15669 22112
rect 15627 22063 15669 22072
rect 16099 22112 16157 22113
rect 16099 22072 16108 22112
rect 16148 22072 16157 22112
rect 16099 22071 16157 22072
rect 9771 22021 9813 22030
rect 4779 22005 4821 22014
rect 1152 21944 20452 21968
rect 1152 21904 4928 21944
rect 4968 21904 5010 21944
rect 5050 21904 5092 21944
rect 5132 21904 5174 21944
rect 5214 21904 5256 21944
rect 5296 21904 20048 21944
rect 20088 21904 20130 21944
rect 20170 21904 20212 21944
rect 20252 21904 20294 21944
rect 20334 21904 20376 21944
rect 20416 21904 20452 21944
rect 1152 21880 20452 21904
rect 3243 21834 3285 21843
rect 3243 21794 3244 21834
rect 3284 21794 3285 21834
rect 3243 21785 3285 21794
rect 3051 21776 3093 21785
rect 3051 21736 3052 21776
rect 3092 21736 3093 21776
rect 3051 21727 3093 21736
rect 4483 21776 4541 21777
rect 4483 21736 4492 21776
rect 4532 21736 4541 21776
rect 4483 21735 4541 21736
rect 7563 21776 7605 21785
rect 7563 21736 7564 21776
rect 7604 21736 7605 21776
rect 7563 21727 7605 21736
rect 14379 21776 14421 21785
rect 14379 21736 14380 21776
rect 14420 21736 14421 21776
rect 14379 21727 14421 21736
rect 18315 21776 18357 21785
rect 18315 21736 18316 21776
rect 18356 21736 18357 21776
rect 18315 21727 18357 21736
rect 20139 21776 20181 21785
rect 20139 21736 20140 21776
rect 20180 21736 20181 21776
rect 20139 21727 20181 21736
rect 2667 21692 2709 21701
rect 2667 21652 2668 21692
rect 2708 21652 2709 21692
rect 2667 21643 2709 21652
rect 10731 21692 10773 21701
rect 10731 21652 10732 21692
rect 10772 21652 10773 21692
rect 10731 21643 10773 21652
rect 12747 21692 12789 21701
rect 12747 21652 12748 21692
rect 12788 21652 12789 21692
rect 12747 21643 12789 21652
rect 15627 21692 15669 21701
rect 15627 21652 15628 21692
rect 15668 21652 15669 21692
rect 15627 21643 15669 21652
rect 17547 21692 17589 21701
rect 17547 21652 17548 21692
rect 17588 21652 17589 21692
rect 17547 21643 17589 21652
rect 1219 21608 1277 21609
rect 1219 21568 1228 21608
rect 1268 21568 1277 21608
rect 1219 21567 1277 21568
rect 2467 21608 2525 21609
rect 2467 21568 2476 21608
rect 2516 21568 2525 21608
rect 2467 21567 2525 21568
rect 2947 21608 3005 21609
rect 2947 21568 2956 21608
rect 2996 21568 3005 21608
rect 2947 21567 3005 21568
rect 3435 21608 3477 21617
rect 3435 21568 3436 21608
rect 3476 21568 3477 21608
rect 3331 21566 3389 21567
rect 3331 21526 3340 21566
rect 3380 21526 3389 21566
rect 3435 21559 3477 21568
rect 3915 21608 3957 21617
rect 3915 21568 3916 21608
rect 3956 21568 3957 21608
rect 3915 21559 3957 21568
rect 4291 21608 4349 21609
rect 4291 21568 4300 21608
rect 4340 21568 4349 21608
rect 4291 21567 4349 21568
rect 4587 21608 4629 21617
rect 4587 21568 4588 21608
rect 4628 21568 4629 21608
rect 4587 21559 4629 21568
rect 4779 21608 4821 21617
rect 4779 21568 4780 21608
rect 4820 21568 4821 21608
rect 4675 21566 4733 21567
rect 3331 21525 3389 21526
rect 4011 21524 4053 21533
rect 4011 21484 4012 21524
rect 4052 21484 4053 21524
rect 4011 21475 4053 21484
rect 4203 21524 4245 21533
rect 4675 21526 4684 21566
rect 4724 21526 4733 21566
rect 4779 21559 4821 21568
rect 5059 21608 5117 21609
rect 5059 21568 5068 21608
rect 5108 21568 5117 21608
rect 5059 21567 5117 21568
rect 6307 21608 6365 21609
rect 6307 21568 6316 21608
rect 6356 21568 6365 21608
rect 6307 21567 6365 21568
rect 6691 21608 6749 21609
rect 6691 21568 6700 21608
rect 6740 21568 6749 21608
rect 6691 21567 6749 21568
rect 7083 21608 7125 21617
rect 7083 21568 7084 21608
rect 7124 21568 7125 21608
rect 7083 21559 7125 21568
rect 7267 21608 7325 21609
rect 7267 21568 7276 21608
rect 7316 21568 7325 21608
rect 7267 21567 7325 21568
rect 7747 21608 7805 21609
rect 7747 21568 7756 21608
rect 7796 21568 7805 21608
rect 7747 21567 7805 21568
rect 8995 21608 9053 21609
rect 8995 21568 9004 21608
rect 9044 21568 9053 21608
rect 8995 21567 9053 21568
rect 9283 21608 9341 21609
rect 9283 21568 9292 21608
rect 9332 21568 9341 21608
rect 9283 21567 9341 21568
rect 10531 21608 10589 21609
rect 10531 21568 10540 21608
rect 10580 21568 10589 21608
rect 10531 21567 10589 21568
rect 11019 21608 11061 21617
rect 11019 21568 11020 21608
rect 11060 21568 11061 21608
rect 11019 21559 11061 21568
rect 11115 21608 11157 21617
rect 11115 21568 11116 21608
rect 11156 21568 11157 21608
rect 11115 21559 11157 21568
rect 11499 21608 11541 21617
rect 11499 21568 11500 21608
rect 11540 21568 11541 21608
rect 11499 21559 11541 21568
rect 11595 21608 11637 21617
rect 11595 21568 11596 21608
rect 11636 21568 11637 21608
rect 11595 21559 11637 21568
rect 12067 21608 12125 21609
rect 12067 21568 12076 21608
rect 12116 21568 12125 21608
rect 12931 21608 12989 21609
rect 12067 21567 12125 21568
rect 12603 21566 12645 21575
rect 12931 21568 12940 21608
rect 12980 21568 12989 21608
rect 12931 21567 12989 21568
rect 14179 21608 14237 21609
rect 14179 21568 14188 21608
rect 14228 21568 14237 21608
rect 14179 21567 14237 21568
rect 14571 21608 14613 21617
rect 14571 21568 14572 21608
rect 14612 21568 14613 21608
rect 4675 21525 4733 21526
rect 4203 21484 4204 21524
rect 4244 21484 4245 21524
rect 4203 21475 4245 21484
rect 6795 21524 6837 21533
rect 6795 21484 6796 21524
rect 6836 21484 6837 21524
rect 6795 21475 6837 21484
rect 6987 21524 7029 21533
rect 6987 21484 6988 21524
rect 7028 21484 7029 21524
rect 12603 21526 12604 21566
rect 12644 21526 12645 21566
rect 14571 21559 14613 21568
rect 14859 21608 14901 21617
rect 14859 21568 14860 21608
rect 14900 21568 14901 21608
rect 14859 21559 14901 21568
rect 15235 21608 15293 21609
rect 15235 21568 15244 21608
rect 15284 21568 15293 21608
rect 15235 21567 15293 21568
rect 15531 21608 15573 21617
rect 15531 21568 15532 21608
rect 15572 21568 15573 21608
rect 15531 21559 15573 21568
rect 16099 21608 16157 21609
rect 16099 21568 16108 21608
rect 16148 21568 16157 21608
rect 16099 21567 16157 21568
rect 17347 21608 17405 21609
rect 17347 21568 17356 21608
rect 17396 21568 17405 21608
rect 17347 21567 17405 21568
rect 18123 21608 18165 21617
rect 18123 21568 18124 21608
rect 18164 21568 18165 21608
rect 18123 21559 18165 21568
rect 18411 21608 18453 21617
rect 18411 21568 18412 21608
rect 18452 21568 18453 21608
rect 18411 21559 18453 21568
rect 18691 21608 18749 21609
rect 18691 21568 18700 21608
rect 18740 21568 18749 21608
rect 18691 21567 18749 21568
rect 19939 21608 19997 21609
rect 19939 21568 19948 21608
rect 19988 21568 19997 21608
rect 19939 21567 19997 21568
rect 12603 21517 12645 21526
rect 6987 21475 7029 21484
rect 3723 21440 3765 21449
rect 3723 21400 3724 21440
rect 3764 21400 3765 21440
rect 3723 21391 3765 21400
rect 4107 21440 4149 21449
rect 4107 21400 4108 21440
rect 4148 21400 4149 21440
rect 4107 21391 4149 21400
rect 6507 21440 6549 21449
rect 6507 21400 6508 21440
rect 6548 21400 6549 21440
rect 6507 21391 6549 21400
rect 6891 21440 6933 21449
rect 6891 21400 6892 21440
rect 6932 21400 6933 21440
rect 6891 21391 6933 21400
rect 15907 21440 15965 21441
rect 15907 21400 15916 21440
rect 15956 21400 15965 21440
rect 15907 21399 15965 21400
rect 3051 21356 3093 21365
rect 3051 21316 3052 21356
rect 3092 21316 3093 21356
rect 3051 21307 3093 21316
rect 7371 21356 7413 21365
rect 7371 21316 7372 21356
rect 7412 21316 7413 21356
rect 7371 21307 7413 21316
rect 14859 21356 14901 21365
rect 14859 21316 14860 21356
rect 14900 21316 14901 21356
rect 14859 21307 14901 21316
rect 1152 21188 20352 21212
rect 1152 21148 3688 21188
rect 3728 21148 3770 21188
rect 3810 21148 3852 21188
rect 3892 21148 3934 21188
rect 3974 21148 4016 21188
rect 4056 21148 18808 21188
rect 18848 21148 18890 21188
rect 18930 21148 18972 21188
rect 19012 21148 19054 21188
rect 19094 21148 19136 21188
rect 19176 21148 20352 21188
rect 1152 21124 20352 21148
rect 2667 21020 2709 21029
rect 2667 20980 2668 21020
rect 2708 20980 2709 21020
rect 2667 20971 2709 20980
rect 4971 21020 5013 21029
rect 4971 20980 4972 21020
rect 5012 20980 5013 21020
rect 4971 20971 5013 20980
rect 6411 21020 6453 21029
rect 6411 20980 6412 21020
rect 6452 20980 6453 21020
rect 6411 20971 6453 20980
rect 7851 21020 7893 21029
rect 7851 20980 7852 21020
rect 7892 20980 7893 21020
rect 7851 20971 7893 20980
rect 12747 21020 12789 21029
rect 12747 20980 12748 21020
rect 12788 20980 12789 21020
rect 12747 20971 12789 20980
rect 14763 21020 14805 21029
rect 14763 20980 14764 21020
rect 14804 20980 14805 21020
rect 14763 20971 14805 20980
rect 14955 21020 14997 21029
rect 14955 20980 14956 21020
rect 14996 20980 14997 21020
rect 14955 20971 14997 20980
rect 4107 20936 4149 20945
rect 4107 20896 4108 20936
rect 4148 20896 4149 20936
rect 4107 20887 4149 20896
rect 4299 20936 4341 20945
rect 4299 20896 4300 20936
rect 4340 20896 4341 20936
rect 4299 20887 4341 20896
rect 7363 20936 7421 20937
rect 7363 20896 7372 20936
rect 7412 20896 7421 20936
rect 7363 20895 7421 20896
rect 17835 20852 17877 20861
rect 17835 20812 17836 20852
rect 17876 20812 17877 20852
rect 17835 20803 17877 20812
rect 17931 20852 17973 20861
rect 17931 20812 17932 20852
rect 17972 20812 17973 20852
rect 17931 20803 17973 20812
rect 18939 20777 18981 20786
rect 1219 20768 1277 20769
rect 1219 20728 1228 20768
rect 1268 20728 1277 20768
rect 1219 20727 1277 20728
rect 2467 20768 2525 20769
rect 2467 20728 2476 20768
rect 2516 20728 2525 20768
rect 2467 20727 2525 20728
rect 2955 20768 2997 20777
rect 2955 20728 2956 20768
rect 2996 20728 2997 20768
rect 2955 20719 2997 20728
rect 3051 20768 3093 20777
rect 3051 20728 3052 20768
rect 3092 20728 3093 20768
rect 3051 20719 3093 20728
rect 3147 20768 3189 20777
rect 3147 20728 3148 20768
rect 3188 20728 3189 20768
rect 3147 20719 3189 20728
rect 3243 20768 3285 20777
rect 3243 20728 3244 20768
rect 3284 20728 3285 20768
rect 3243 20719 3285 20728
rect 3523 20768 3581 20769
rect 3523 20728 3532 20768
rect 3572 20728 3581 20768
rect 3523 20727 3581 20728
rect 3627 20768 3669 20777
rect 3627 20728 3628 20768
rect 3668 20728 3669 20768
rect 3627 20719 3669 20728
rect 3819 20768 3861 20777
rect 3819 20728 3820 20768
rect 3860 20728 3861 20768
rect 3819 20719 3861 20728
rect 4107 20768 4149 20777
rect 4107 20728 4108 20768
rect 4148 20728 4149 20768
rect 4107 20719 4149 20728
rect 4587 20768 4629 20777
rect 4587 20728 4588 20768
rect 4628 20728 4629 20768
rect 4587 20719 4629 20728
rect 4683 20768 4725 20777
rect 4683 20728 4684 20768
rect 4724 20728 4725 20768
rect 4683 20719 4725 20728
rect 4779 20768 4821 20777
rect 4779 20728 4780 20768
rect 4820 20728 4821 20768
rect 4779 20719 4821 20728
rect 5059 20768 5117 20769
rect 5059 20728 5068 20768
rect 5108 20728 5117 20768
rect 5059 20727 5117 20728
rect 5547 20768 5589 20777
rect 5547 20728 5548 20768
rect 5588 20728 5589 20768
rect 5547 20719 5589 20728
rect 5643 20768 5685 20777
rect 5643 20728 5644 20768
rect 5684 20728 5685 20768
rect 5643 20719 5685 20728
rect 5739 20768 5781 20777
rect 5739 20728 5740 20768
rect 5780 20728 5781 20768
rect 5739 20719 5781 20728
rect 6019 20768 6077 20769
rect 6019 20728 6028 20768
rect 6068 20728 6077 20768
rect 6019 20727 6077 20728
rect 6123 20768 6165 20777
rect 6123 20728 6124 20768
rect 6164 20728 6165 20768
rect 6123 20719 6165 20728
rect 6691 20768 6749 20769
rect 6691 20728 6700 20768
rect 6740 20728 6749 20768
rect 6691 20727 6749 20728
rect 6987 20768 7029 20777
rect 6987 20728 6988 20768
rect 7028 20728 7029 20768
rect 6987 20719 7029 20728
rect 7083 20768 7125 20777
rect 7083 20728 7084 20768
rect 7124 20728 7125 20768
rect 7083 20719 7125 20728
rect 7555 20768 7613 20769
rect 7555 20728 7564 20768
rect 7604 20728 7613 20768
rect 7555 20727 7613 20728
rect 7659 20768 7701 20777
rect 7659 20728 7660 20768
rect 7700 20728 7701 20768
rect 7659 20719 7701 20728
rect 7851 20768 7893 20777
rect 7851 20728 7852 20768
rect 7892 20728 7893 20768
rect 7851 20719 7893 20728
rect 9387 20768 9429 20777
rect 9387 20728 9388 20768
rect 9428 20728 9429 20768
rect 9387 20719 9429 20728
rect 9483 20768 9525 20777
rect 9483 20728 9484 20768
rect 9524 20728 9525 20768
rect 9483 20719 9525 20728
rect 9579 20768 9621 20777
rect 9579 20728 9580 20768
rect 9620 20728 9621 20768
rect 9579 20719 9621 20728
rect 11299 20768 11357 20769
rect 11299 20728 11308 20768
rect 11348 20728 11357 20768
rect 11299 20727 11357 20728
rect 12547 20768 12605 20769
rect 12547 20728 12556 20768
rect 12596 20728 12605 20768
rect 12547 20727 12605 20728
rect 13315 20768 13373 20769
rect 13315 20728 13324 20768
rect 13364 20728 13373 20768
rect 13315 20727 13373 20728
rect 14563 20768 14621 20769
rect 14563 20728 14572 20768
rect 14612 20728 14621 20768
rect 14563 20727 14621 20728
rect 15139 20768 15197 20769
rect 15139 20728 15148 20768
rect 15188 20728 15197 20768
rect 15139 20727 15197 20728
rect 16387 20768 16445 20769
rect 16387 20728 16396 20768
rect 16436 20728 16445 20768
rect 16387 20727 16445 20728
rect 17355 20768 17397 20777
rect 17355 20728 17356 20768
rect 17396 20728 17397 20768
rect 17355 20719 17397 20728
rect 17451 20768 17493 20777
rect 17451 20728 17452 20768
rect 17492 20728 17493 20768
rect 17451 20719 17493 20728
rect 18403 20768 18461 20769
rect 18403 20728 18412 20768
rect 18452 20728 18461 20768
rect 18939 20737 18940 20777
rect 18980 20737 18981 20777
rect 18939 20728 18981 20737
rect 19371 20768 19413 20777
rect 19371 20728 19372 20768
rect 19412 20728 19413 20768
rect 18403 20727 18461 20728
rect 19371 20719 19413 20728
rect 19467 20768 19509 20777
rect 19467 20728 19468 20768
rect 19508 20728 19509 20768
rect 19467 20719 19509 20728
rect 19563 20768 19605 20777
rect 19563 20728 19564 20768
rect 19604 20728 19605 20768
rect 19563 20719 19605 20728
rect 19947 20768 19989 20777
rect 19947 20728 19948 20768
rect 19988 20728 19989 20768
rect 19947 20719 19989 20728
rect 20043 20768 20085 20777
rect 20043 20728 20044 20768
rect 20084 20728 20085 20768
rect 20043 20719 20085 20728
rect 20139 20747 20181 20756
rect 20139 20707 20140 20747
rect 20180 20707 20181 20747
rect 20139 20698 20181 20707
rect 3723 20684 3765 20693
rect 3723 20644 3724 20684
rect 3764 20644 3765 20684
rect 3723 20635 3765 20644
rect 4483 20600 4541 20601
rect 4483 20560 4492 20600
rect 4532 20560 4541 20600
rect 4483 20559 4541 20560
rect 5443 20600 5501 20601
rect 5443 20560 5452 20600
rect 5492 20560 5501 20600
rect 5443 20559 5501 20560
rect 5931 20596 5973 20605
rect 5931 20556 5932 20596
rect 5972 20556 5973 20596
rect 9667 20600 9725 20601
rect 9667 20560 9676 20600
rect 9716 20560 9725 20600
rect 9667 20559 9725 20560
rect 14763 20600 14805 20609
rect 14763 20560 14764 20600
rect 14804 20560 14805 20600
rect 5931 20547 5973 20556
rect 14763 20551 14805 20560
rect 19083 20600 19125 20609
rect 19083 20560 19084 20600
rect 19124 20560 19125 20600
rect 19083 20551 19125 20560
rect 19755 20600 19797 20609
rect 19755 20560 19756 20600
rect 19796 20560 19797 20600
rect 19755 20551 19797 20560
rect 20227 20600 20285 20601
rect 20227 20560 20236 20600
rect 20276 20560 20285 20600
rect 20227 20559 20285 20560
rect 1152 20432 20452 20456
rect 1152 20392 4928 20432
rect 4968 20392 5010 20432
rect 5050 20392 5092 20432
rect 5132 20392 5174 20432
rect 5214 20392 5256 20432
rect 5296 20392 20048 20432
rect 20088 20392 20130 20432
rect 20170 20392 20212 20432
rect 20252 20392 20294 20432
rect 20334 20392 20376 20432
rect 20416 20392 20452 20432
rect 1152 20368 20452 20392
rect 2667 20264 2709 20273
rect 2667 20224 2668 20264
rect 2708 20224 2709 20264
rect 2667 20215 2709 20224
rect 6603 20268 6645 20277
rect 6603 20228 6604 20268
rect 6644 20228 6645 20268
rect 6603 20219 6645 20228
rect 7851 20264 7893 20273
rect 7851 20224 7852 20264
rect 7892 20224 7893 20264
rect 7851 20215 7893 20224
rect 6411 20180 6453 20189
rect 6411 20140 6412 20180
rect 6452 20140 6453 20180
rect 6411 20131 6453 20140
rect 10731 20180 10773 20189
rect 10731 20140 10732 20180
rect 10772 20140 10773 20180
rect 10731 20131 10773 20140
rect 12747 20180 12789 20189
rect 12747 20140 12748 20180
rect 12788 20140 12789 20180
rect 12747 20131 12789 20140
rect 15051 20180 15093 20189
rect 15051 20140 15052 20180
rect 15092 20140 15093 20180
rect 15051 20131 15093 20140
rect 1219 20096 1277 20097
rect 1219 20056 1228 20096
rect 1268 20056 1277 20096
rect 1219 20055 1277 20056
rect 2467 20096 2525 20097
rect 2467 20056 2476 20096
rect 2516 20056 2525 20096
rect 2467 20055 2525 20056
rect 2851 20096 2909 20097
rect 2851 20056 2860 20096
rect 2900 20056 2909 20096
rect 2851 20055 2909 20056
rect 4099 20096 4157 20097
rect 4099 20056 4108 20096
rect 4148 20056 4157 20096
rect 4099 20055 4157 20056
rect 4579 20096 4637 20097
rect 4579 20056 4588 20096
rect 4628 20056 4637 20096
rect 4579 20055 4637 20056
rect 4963 20096 5021 20097
rect 4963 20056 4972 20096
rect 5012 20056 5021 20096
rect 4963 20055 5021 20056
rect 5259 20096 5301 20105
rect 5259 20056 5260 20096
rect 5300 20056 5301 20096
rect 5259 20047 5301 20056
rect 5355 20096 5397 20105
rect 5355 20056 5356 20096
rect 5396 20056 5397 20096
rect 5355 20047 5397 20056
rect 5827 20096 5885 20097
rect 5827 20056 5836 20096
rect 5876 20056 5885 20096
rect 5827 20055 5885 20056
rect 6307 20096 6365 20097
rect 6307 20056 6316 20096
rect 6356 20056 6365 20096
rect 6307 20055 6365 20056
rect 6691 20096 6749 20097
rect 6691 20056 6700 20096
rect 6740 20056 6749 20096
rect 6691 20055 6749 20056
rect 6795 20096 6837 20105
rect 6795 20056 6796 20096
rect 6836 20056 6837 20096
rect 6795 20047 6837 20056
rect 7275 20096 7317 20105
rect 7275 20056 7276 20096
rect 7316 20056 7317 20096
rect 7275 20047 7317 20056
rect 7467 20096 7509 20105
rect 7467 20056 7468 20096
rect 7508 20056 7509 20096
rect 7467 20047 7509 20056
rect 7555 20096 7613 20097
rect 7555 20056 7564 20096
rect 7604 20056 7613 20096
rect 7555 20055 7613 20056
rect 7747 20096 7805 20097
rect 7747 20056 7756 20096
rect 7796 20056 7805 20096
rect 7747 20055 7805 20056
rect 9283 20096 9341 20097
rect 9283 20056 9292 20096
rect 9332 20056 9341 20096
rect 9283 20055 9341 20056
rect 10531 20096 10589 20097
rect 10531 20056 10540 20096
rect 10580 20056 10589 20096
rect 10531 20055 10589 20056
rect 11019 20096 11061 20105
rect 11019 20056 11020 20096
rect 11060 20056 11061 20096
rect 11019 20047 11061 20056
rect 11115 20096 11157 20105
rect 11115 20056 11116 20096
rect 11156 20056 11157 20096
rect 11115 20047 11157 20056
rect 11595 20096 11637 20105
rect 11595 20056 11596 20096
rect 11636 20056 11637 20096
rect 11595 20047 11637 20056
rect 12067 20096 12125 20097
rect 12067 20056 12076 20096
rect 12116 20056 12125 20096
rect 12931 20096 12989 20097
rect 12067 20055 12125 20056
rect 12555 20082 12597 20091
rect 12555 20042 12556 20082
rect 12596 20042 12597 20082
rect 12931 20056 12940 20096
rect 12980 20056 12989 20096
rect 12931 20055 12989 20056
rect 14179 20096 14237 20097
rect 14179 20056 14188 20096
rect 14228 20056 14237 20096
rect 14179 20055 14237 20056
rect 14955 20096 14997 20105
rect 14955 20056 14956 20096
rect 14996 20056 14997 20096
rect 14955 20047 14997 20056
rect 15147 20096 15189 20105
rect 15147 20056 15148 20096
rect 15188 20056 15189 20096
rect 15147 20047 15189 20056
rect 15235 20096 15293 20097
rect 15235 20056 15244 20096
rect 15284 20056 15293 20096
rect 15235 20055 15293 20056
rect 16483 20096 16541 20097
rect 16483 20056 16492 20096
rect 16532 20056 16541 20096
rect 16483 20055 16541 20056
rect 17731 20096 17789 20097
rect 17731 20056 17740 20096
rect 17780 20056 17789 20096
rect 17731 20055 17789 20056
rect 18123 20096 18165 20105
rect 18123 20056 18124 20096
rect 18164 20056 18165 20096
rect 18123 20047 18165 20056
rect 18411 20096 18453 20105
rect 18411 20056 18412 20096
rect 18452 20056 18453 20096
rect 18411 20047 18453 20056
rect 18691 20096 18749 20097
rect 18691 20056 18700 20096
rect 18740 20056 18749 20096
rect 18691 20055 18749 20056
rect 19939 20096 19997 20097
rect 19939 20056 19948 20096
rect 19988 20056 19997 20096
rect 19939 20055 19997 20056
rect 12555 20033 12597 20042
rect 4491 20012 4533 20021
rect 4491 19972 4492 20012
rect 4532 19972 4533 20012
rect 4491 19963 4533 19972
rect 11499 20012 11541 20021
rect 11499 19972 11500 20012
rect 11540 19972 11541 20012
rect 11499 19963 11541 19972
rect 7083 19928 7125 19937
rect 7083 19888 7084 19928
rect 7124 19888 7125 19928
rect 7083 19879 7125 19888
rect 7275 19928 7317 19937
rect 7275 19888 7276 19928
rect 7316 19888 7317 19928
rect 7275 19879 7317 19888
rect 17931 19928 17973 19937
rect 17931 19888 17932 19928
rect 17972 19888 17973 19928
rect 17931 19879 17973 19888
rect 2667 19844 2709 19853
rect 2667 19804 2668 19844
rect 2708 19804 2709 19844
rect 2667 19795 2709 19804
rect 4299 19844 4341 19853
rect 4299 19804 4300 19844
rect 4340 19804 4341 19844
rect 4299 19795 4341 19804
rect 5635 19844 5693 19845
rect 5635 19804 5644 19844
rect 5684 19804 5693 19844
rect 5635 19803 5693 19804
rect 5931 19844 5973 19853
rect 5931 19804 5932 19844
rect 5972 19804 5973 19844
rect 5931 19795 5973 19804
rect 14379 19844 14421 19853
rect 14379 19804 14380 19844
rect 14420 19804 14421 19844
rect 14379 19795 14421 19804
rect 18411 19844 18453 19853
rect 18411 19804 18412 19844
rect 18452 19804 18453 19844
rect 18411 19795 18453 19804
rect 20139 19844 20181 19853
rect 20139 19804 20140 19844
rect 20180 19804 20181 19844
rect 20139 19795 20181 19804
rect 1152 19676 20352 19700
rect 1152 19636 3688 19676
rect 3728 19636 3770 19676
rect 3810 19636 3852 19676
rect 3892 19636 3934 19676
rect 3974 19636 4016 19676
rect 4056 19636 18808 19676
rect 18848 19636 18890 19676
rect 18930 19636 18972 19676
rect 19012 19636 19054 19676
rect 19094 19636 19136 19676
rect 19176 19636 20352 19676
rect 1152 19612 20352 19636
rect 4395 19508 4437 19517
rect 4395 19468 4396 19508
rect 4436 19468 4437 19508
rect 4395 19459 4437 19468
rect 12555 19508 12597 19517
rect 12555 19468 12556 19508
rect 12596 19468 12597 19508
rect 12555 19459 12597 19468
rect 15915 19508 15957 19517
rect 15915 19468 15916 19508
rect 15956 19468 15957 19508
rect 15915 19459 15957 19468
rect 19275 19508 19317 19517
rect 19275 19468 19276 19508
rect 19316 19468 19317 19508
rect 19275 19459 19317 19468
rect 1995 19424 2037 19433
rect 1995 19384 1996 19424
rect 2036 19384 2037 19424
rect 1995 19375 2037 19384
rect 20227 19424 20285 19425
rect 20227 19384 20236 19424
rect 20276 19384 20285 19424
rect 20227 19383 20285 19384
rect 8715 19340 8757 19349
rect 8715 19300 8716 19340
rect 8756 19300 8757 19340
rect 8715 19291 8757 19300
rect 16099 19298 16157 19299
rect 4059 19265 4101 19274
rect 9819 19265 9861 19274
rect 1995 19256 2037 19265
rect 1995 19216 1996 19256
rect 2036 19216 2037 19256
rect 1995 19207 2037 19216
rect 2475 19256 2517 19265
rect 2475 19216 2476 19256
rect 2516 19216 2517 19256
rect 2475 19207 2517 19216
rect 2571 19256 2613 19265
rect 2571 19216 2572 19256
rect 2612 19216 2613 19256
rect 2571 19207 2613 19216
rect 2955 19256 2997 19265
rect 2955 19216 2956 19256
rect 2996 19216 2997 19256
rect 2955 19207 2997 19216
rect 3051 19256 3093 19265
rect 3051 19216 3052 19256
rect 3092 19216 3093 19256
rect 3051 19207 3093 19216
rect 3523 19256 3581 19257
rect 3523 19216 3532 19256
rect 3572 19216 3581 19256
rect 4059 19225 4060 19265
rect 4100 19225 4101 19265
rect 4059 19216 4101 19225
rect 4579 19256 4637 19257
rect 4579 19216 4588 19256
rect 4628 19216 4637 19256
rect 3523 19215 3581 19216
rect 4579 19215 4637 19216
rect 5827 19256 5885 19257
rect 5827 19216 5836 19256
rect 5876 19216 5885 19256
rect 5827 19215 5885 19216
rect 6499 19256 6557 19257
rect 6499 19216 6508 19256
rect 6548 19216 6557 19256
rect 6499 19215 6557 19216
rect 7747 19256 7805 19257
rect 7747 19216 7756 19256
rect 7796 19216 7805 19256
rect 7747 19215 7805 19216
rect 8235 19255 8277 19264
rect 8235 19215 8236 19255
rect 8276 19215 8277 19255
rect 8235 19206 8277 19215
rect 8331 19256 8373 19265
rect 8331 19216 8332 19256
rect 8372 19216 8373 19256
rect 8331 19207 8373 19216
rect 8811 19256 8853 19265
rect 8811 19216 8812 19256
rect 8852 19216 8853 19256
rect 8811 19207 8853 19216
rect 9283 19256 9341 19257
rect 9283 19216 9292 19256
rect 9332 19216 9341 19256
rect 9819 19225 9820 19265
rect 9860 19225 9861 19265
rect 9819 19216 9861 19225
rect 11107 19256 11165 19257
rect 11107 19216 11116 19256
rect 11156 19216 11165 19256
rect 9283 19215 9341 19216
rect 11107 19215 11165 19216
rect 12355 19256 12413 19257
rect 12355 19216 12364 19256
rect 12404 19216 12413 19256
rect 12355 19215 12413 19216
rect 13995 19256 14037 19265
rect 13995 19216 13996 19256
rect 14036 19216 14037 19256
rect 13995 19207 14037 19216
rect 14091 19256 14133 19265
rect 14091 19216 14092 19256
rect 14132 19216 14133 19256
rect 14091 19207 14133 19216
rect 14475 19256 14517 19265
rect 14475 19216 14476 19256
rect 14516 19216 14517 19256
rect 14475 19207 14517 19216
rect 14571 19256 14613 19265
rect 15531 19261 15573 19270
rect 14571 19216 14572 19256
rect 14612 19216 14613 19256
rect 14571 19207 14613 19216
rect 15043 19256 15101 19257
rect 15043 19216 15052 19256
rect 15092 19216 15101 19256
rect 15043 19215 15101 19216
rect 15531 19221 15532 19261
rect 15572 19221 15573 19261
rect 16099 19258 16108 19298
rect 16148 19258 16157 19298
rect 16099 19257 16157 19258
rect 15531 19212 15573 19221
rect 17347 19256 17405 19257
rect 17347 19216 17356 19256
rect 17396 19216 17405 19256
rect 17347 19215 17405 19216
rect 17827 19256 17885 19257
rect 17827 19216 17836 19256
rect 17876 19216 17885 19256
rect 17827 19215 17885 19216
rect 19075 19256 19133 19257
rect 19075 19216 19084 19256
rect 19124 19216 19133 19256
rect 19075 19215 19133 19216
rect 19555 19256 19613 19257
rect 19555 19216 19564 19256
rect 19604 19216 19613 19256
rect 19555 19215 19613 19216
rect 19851 19256 19893 19265
rect 19851 19216 19852 19256
rect 19892 19216 19893 19256
rect 19851 19207 19893 19216
rect 19947 19256 19989 19265
rect 19947 19216 19948 19256
rect 19988 19216 19989 19256
rect 19947 19207 19989 19216
rect 4203 19172 4245 19181
rect 4203 19132 4204 19172
rect 4244 19132 4245 19172
rect 4203 19123 4245 19132
rect 7947 19172 7989 19181
rect 7947 19132 7948 19172
rect 7988 19132 7989 19172
rect 7947 19123 7989 19132
rect 2187 19088 2229 19097
rect 2187 19048 2188 19088
rect 2228 19048 2229 19088
rect 2187 19039 2229 19048
rect 9963 19088 10005 19097
rect 9963 19048 9964 19088
rect 10004 19048 10005 19088
rect 19275 19088 19317 19097
rect 9963 19039 10005 19048
rect 15723 19046 15765 19055
rect 15723 19006 15724 19046
rect 15764 19006 15765 19046
rect 19275 19048 19276 19088
rect 19316 19048 19317 19088
rect 19275 19039 19317 19048
rect 15723 18997 15765 19006
rect 1152 18920 20452 18944
rect 1152 18880 4928 18920
rect 4968 18880 5010 18920
rect 5050 18880 5092 18920
rect 5132 18880 5174 18920
rect 5214 18880 5256 18920
rect 5296 18880 20048 18920
rect 20088 18880 20130 18920
rect 20170 18880 20212 18920
rect 20252 18880 20294 18920
rect 20334 18880 20376 18920
rect 20416 18880 20452 18920
rect 1152 18856 20452 18880
rect 4867 18752 4925 18753
rect 4867 18712 4876 18752
rect 4916 18712 4925 18752
rect 4867 18711 4925 18712
rect 7083 18752 7125 18761
rect 7083 18712 7084 18752
rect 7124 18712 7125 18752
rect 7083 18703 7125 18712
rect 9867 18752 9909 18761
rect 9867 18712 9868 18752
rect 9908 18712 9909 18752
rect 9867 18703 9909 18712
rect 16299 18752 16341 18761
rect 16299 18712 16300 18752
rect 16340 18712 16341 18752
rect 16299 18703 16341 18712
rect 16491 18752 16533 18761
rect 16491 18712 16492 18752
rect 16532 18712 16533 18752
rect 16491 18703 16533 18712
rect 18883 18752 18941 18753
rect 18883 18712 18892 18752
rect 18932 18712 18941 18752
rect 18883 18711 18941 18712
rect 3435 18668 3477 18677
rect 3435 18628 3436 18668
rect 3476 18628 3477 18668
rect 3435 18619 3477 18628
rect 13515 18668 13557 18677
rect 13515 18628 13516 18668
rect 13556 18628 13557 18668
rect 13515 18619 13557 18628
rect 15531 18668 15573 18677
rect 15531 18628 15532 18668
rect 15572 18628 15573 18668
rect 15531 18619 15573 18628
rect 1707 18584 1749 18593
rect 1707 18544 1708 18584
rect 1748 18544 1749 18584
rect 1707 18535 1749 18544
rect 1803 18584 1845 18593
rect 1803 18544 1804 18584
rect 1844 18544 1845 18584
rect 1803 18535 1845 18544
rect 2187 18584 2229 18593
rect 2187 18544 2188 18584
rect 2228 18544 2229 18584
rect 2187 18535 2229 18544
rect 2283 18584 2325 18593
rect 2283 18544 2284 18584
rect 2324 18544 2325 18584
rect 2283 18535 2325 18544
rect 2755 18584 2813 18585
rect 2755 18544 2764 18584
rect 2804 18544 2813 18584
rect 3619 18584 3677 18585
rect 2755 18543 2813 18544
rect 3243 18570 3285 18579
rect 3243 18530 3244 18570
rect 3284 18530 3285 18570
rect 3619 18544 3628 18584
rect 3668 18544 3677 18584
rect 3619 18543 3677 18544
rect 3819 18584 3861 18593
rect 3819 18544 3820 18584
rect 3860 18544 3861 18584
rect 3819 18535 3861 18544
rect 3907 18584 3965 18585
rect 3907 18544 3916 18584
rect 3956 18544 3965 18584
rect 3907 18543 3965 18544
rect 4099 18584 4157 18585
rect 4099 18544 4108 18584
rect 4148 18544 4157 18584
rect 4099 18543 4157 18544
rect 4203 18584 4245 18593
rect 4203 18544 4204 18584
rect 4244 18544 4245 18584
rect 4203 18535 4245 18544
rect 4387 18584 4445 18585
rect 4387 18544 4396 18584
rect 4436 18544 4445 18584
rect 4387 18543 4445 18544
rect 4587 18584 4629 18593
rect 4587 18544 4588 18584
rect 4628 18544 4629 18584
rect 4587 18535 4629 18544
rect 4683 18584 4725 18593
rect 4683 18544 4684 18584
rect 4724 18544 4725 18584
rect 4683 18535 4725 18544
rect 4779 18584 4821 18593
rect 4779 18544 4780 18584
rect 4820 18544 4821 18584
rect 4779 18535 4821 18544
rect 5635 18584 5693 18585
rect 5635 18544 5644 18584
rect 5684 18544 5693 18584
rect 5635 18543 5693 18544
rect 6883 18584 6941 18585
rect 6883 18544 6892 18584
rect 6932 18544 6941 18584
rect 6883 18543 6941 18544
rect 8419 18584 8477 18585
rect 8419 18544 8428 18584
rect 8468 18544 8477 18584
rect 8419 18543 8477 18544
rect 9667 18584 9725 18585
rect 9667 18544 9676 18584
rect 9716 18544 9725 18584
rect 9667 18543 9725 18544
rect 10051 18584 10109 18585
rect 10051 18544 10060 18584
rect 10100 18544 10109 18584
rect 10051 18543 10109 18544
rect 11299 18584 11357 18585
rect 11299 18544 11308 18584
rect 11348 18544 11357 18584
rect 11299 18543 11357 18544
rect 12067 18584 12125 18585
rect 12067 18544 12076 18584
rect 12116 18544 12125 18584
rect 12067 18543 12125 18544
rect 13315 18584 13373 18585
rect 13315 18544 13324 18584
rect 13364 18544 13373 18584
rect 13315 18543 13373 18544
rect 13803 18584 13845 18593
rect 13803 18544 13804 18584
rect 13844 18544 13845 18584
rect 13803 18535 13845 18544
rect 13899 18584 13941 18593
rect 13899 18544 13900 18584
rect 13940 18544 13941 18584
rect 13899 18535 13941 18544
rect 14851 18584 14909 18585
rect 14851 18544 14860 18584
rect 14900 18544 14909 18584
rect 17155 18584 17213 18585
rect 14851 18543 14909 18544
rect 15387 18542 15429 18551
rect 17155 18544 17164 18584
rect 17204 18544 17213 18584
rect 17155 18543 17213 18544
rect 18403 18584 18461 18585
rect 18403 18544 18412 18584
rect 18452 18544 18461 18584
rect 18403 18543 18461 18544
rect 18795 18584 18837 18593
rect 18795 18544 18796 18584
rect 18836 18544 18837 18584
rect 3243 18521 3285 18530
rect 14283 18500 14325 18509
rect 14283 18460 14284 18500
rect 14324 18460 14325 18500
rect 14283 18451 14325 18460
rect 14379 18500 14421 18509
rect 14379 18460 14380 18500
rect 14420 18460 14421 18500
rect 15387 18502 15388 18542
rect 15428 18502 15429 18542
rect 18795 18535 18837 18544
rect 18987 18584 19029 18593
rect 18987 18544 18988 18584
rect 19028 18544 19029 18584
rect 18987 18535 19029 18544
rect 19075 18584 19133 18585
rect 19075 18544 19084 18584
rect 19124 18544 19133 18584
rect 19075 18543 19133 18544
rect 15387 18493 15429 18502
rect 16099 18500 16157 18501
rect 14379 18451 14421 18460
rect 16099 18460 16108 18500
rect 16148 18460 16157 18500
rect 16099 18459 16157 18460
rect 16675 18500 16733 18501
rect 16675 18460 16684 18500
rect 16724 18460 16733 18500
rect 16675 18459 16733 18460
rect 3627 18332 3669 18341
rect 3627 18292 3628 18332
rect 3668 18292 3669 18332
rect 3627 18283 3669 18292
rect 4203 18332 4245 18341
rect 4203 18292 4204 18332
rect 4244 18292 4245 18332
rect 4203 18283 4245 18292
rect 11499 18332 11541 18341
rect 11499 18292 11500 18332
rect 11540 18292 11541 18332
rect 11499 18283 11541 18292
rect 18603 18332 18645 18341
rect 18603 18292 18604 18332
rect 18644 18292 18645 18332
rect 18603 18283 18645 18292
rect 1152 18164 20352 18188
rect 1152 18124 3688 18164
rect 3728 18124 3770 18164
rect 3810 18124 3852 18164
rect 3892 18124 3934 18164
rect 3974 18124 4016 18164
rect 4056 18124 18808 18164
rect 18848 18124 18890 18164
rect 18930 18124 18972 18164
rect 19012 18124 19054 18164
rect 19094 18124 19136 18164
rect 19176 18124 20352 18164
rect 1152 18100 20352 18124
rect 3627 17996 3669 18005
rect 3627 17956 3628 17996
rect 3668 17956 3669 17996
rect 3627 17947 3669 17956
rect 15627 17996 15669 18005
rect 15627 17956 15628 17996
rect 15668 17956 15669 17996
rect 15627 17947 15669 17956
rect 7659 17828 7701 17837
rect 7659 17788 7660 17828
rect 7700 17788 7701 17828
rect 7659 17779 7701 17788
rect 10251 17828 10293 17837
rect 10251 17788 10252 17828
rect 10292 17788 10293 17828
rect 10251 17779 10293 17788
rect 11259 17786 11301 17795
rect 1219 17744 1277 17745
rect 1219 17704 1228 17744
rect 1268 17704 1277 17744
rect 1219 17703 1277 17704
rect 2467 17744 2525 17745
rect 2467 17704 2476 17744
rect 2516 17704 2525 17744
rect 2467 17703 2525 17704
rect 3147 17744 3189 17753
rect 3147 17704 3148 17744
rect 3188 17704 3189 17744
rect 3147 17695 3189 17704
rect 3243 17744 3285 17753
rect 3243 17704 3244 17744
rect 3284 17704 3285 17744
rect 3243 17695 3285 17704
rect 3339 17744 3381 17753
rect 3339 17704 3340 17744
rect 3380 17704 3381 17744
rect 3339 17695 3381 17704
rect 3523 17744 3581 17745
rect 3523 17704 3532 17744
rect 3572 17704 3581 17744
rect 3523 17703 3581 17704
rect 3811 17744 3869 17745
rect 3811 17704 3820 17744
rect 3860 17704 3869 17744
rect 3811 17703 3869 17704
rect 5059 17744 5117 17745
rect 5059 17704 5068 17744
rect 5108 17704 5117 17744
rect 5059 17703 5117 17704
rect 5443 17744 5501 17745
rect 5443 17704 5452 17744
rect 5492 17704 5501 17744
rect 5443 17703 5501 17704
rect 6691 17744 6749 17745
rect 6691 17704 6700 17744
rect 6740 17704 6749 17744
rect 6691 17703 6749 17704
rect 7179 17744 7221 17753
rect 7179 17704 7180 17744
rect 7220 17704 7221 17744
rect 7179 17695 7221 17704
rect 7275 17744 7317 17753
rect 7275 17704 7276 17744
rect 7316 17704 7317 17744
rect 7275 17695 7317 17704
rect 7755 17744 7797 17753
rect 8715 17749 8757 17758
rect 7755 17704 7756 17744
rect 7796 17704 7797 17744
rect 7755 17695 7797 17704
rect 8227 17744 8285 17745
rect 8227 17704 8236 17744
rect 8276 17704 8285 17744
rect 8227 17703 8285 17704
rect 8715 17709 8716 17749
rect 8756 17709 8757 17749
rect 8715 17700 8757 17709
rect 9675 17744 9717 17753
rect 9675 17704 9676 17744
rect 9716 17704 9717 17744
rect 9675 17695 9717 17704
rect 9771 17744 9813 17753
rect 9771 17704 9772 17744
rect 9812 17704 9813 17744
rect 9771 17695 9813 17704
rect 10155 17744 10197 17753
rect 11259 17746 11260 17786
rect 11300 17746 11301 17786
rect 18459 17786 18501 17795
rect 10155 17704 10156 17744
rect 10196 17704 10197 17744
rect 10155 17695 10197 17704
rect 10723 17744 10781 17745
rect 10723 17704 10732 17744
rect 10772 17704 10781 17744
rect 11259 17737 11301 17746
rect 12075 17744 12117 17753
rect 10723 17703 10781 17704
rect 12075 17704 12076 17744
rect 12116 17704 12117 17744
rect 12075 17695 12117 17704
rect 12171 17744 12213 17753
rect 12171 17704 12172 17744
rect 12212 17704 12213 17744
rect 12171 17695 12213 17704
rect 12555 17744 12597 17753
rect 12555 17704 12556 17744
rect 12596 17704 12597 17744
rect 12555 17695 12597 17704
rect 12651 17744 12693 17753
rect 13611 17749 13653 17758
rect 12651 17704 12652 17744
rect 12692 17704 12693 17744
rect 12651 17695 12693 17704
rect 13123 17744 13181 17745
rect 13123 17704 13132 17744
rect 13172 17704 13181 17744
rect 13123 17703 13181 17704
rect 13611 17709 13612 17749
rect 13652 17709 13653 17749
rect 13611 17700 13653 17709
rect 14179 17744 14237 17745
rect 14179 17704 14188 17744
rect 14228 17704 14237 17744
rect 14179 17703 14237 17704
rect 15427 17744 15485 17745
rect 15427 17704 15436 17744
rect 15476 17704 15485 17744
rect 15427 17703 15485 17704
rect 16875 17744 16917 17753
rect 16875 17704 16876 17744
rect 16916 17704 16917 17744
rect 17355 17744 17397 17753
rect 16875 17695 16917 17704
rect 16971 17724 17013 17733
rect 16971 17684 16972 17724
rect 17012 17684 17013 17724
rect 17355 17704 17356 17744
rect 17396 17704 17397 17744
rect 17355 17695 17397 17704
rect 17451 17744 17493 17753
rect 18459 17746 18460 17786
rect 18500 17746 18501 17786
rect 17451 17704 17452 17744
rect 17492 17704 17493 17744
rect 17451 17695 17493 17704
rect 17923 17744 17981 17745
rect 17923 17704 17932 17744
rect 17972 17704 17981 17744
rect 18459 17737 18501 17746
rect 18979 17744 19037 17745
rect 17923 17703 17981 17704
rect 18979 17704 18988 17744
rect 19028 17704 19037 17744
rect 18979 17703 19037 17704
rect 20227 17744 20285 17745
rect 20227 17704 20236 17744
rect 20276 17704 20285 17744
rect 20227 17703 20285 17704
rect 16971 17675 17013 17684
rect 2667 17660 2709 17669
rect 2667 17620 2668 17660
rect 2708 17620 2709 17660
rect 2667 17611 2709 17620
rect 5259 17660 5301 17669
rect 5259 17620 5260 17660
rect 5300 17620 5301 17660
rect 5259 17611 5301 17620
rect 6891 17660 6933 17669
rect 6891 17620 6892 17660
rect 6932 17620 6933 17660
rect 6891 17611 6933 17620
rect 8907 17660 8949 17669
rect 8907 17620 8908 17660
rect 8948 17620 8949 17660
rect 8907 17611 8949 17620
rect 11403 17660 11445 17669
rect 11403 17620 11404 17660
rect 11444 17620 11445 17660
rect 11403 17611 11445 17620
rect 13803 17660 13845 17669
rect 13803 17620 13804 17660
rect 13844 17620 13845 17660
rect 13803 17611 13845 17620
rect 3043 17576 3101 17577
rect 3043 17536 3052 17576
rect 3092 17536 3101 17576
rect 3043 17535 3101 17536
rect 18603 17576 18645 17585
rect 18603 17536 18604 17576
rect 18644 17536 18645 17576
rect 18603 17527 18645 17536
rect 18795 17576 18837 17585
rect 18795 17536 18796 17576
rect 18836 17536 18837 17576
rect 18795 17527 18837 17536
rect 1152 17408 20452 17432
rect 1152 17368 4928 17408
rect 4968 17368 5010 17408
rect 5050 17368 5092 17408
rect 5132 17368 5174 17408
rect 5214 17368 5256 17408
rect 5296 17368 20048 17408
rect 20088 17368 20130 17408
rect 20170 17368 20212 17408
rect 20252 17368 20294 17408
rect 20334 17368 20376 17408
rect 20416 17368 20452 17408
rect 1152 17344 20452 17368
rect 2763 17240 2805 17249
rect 2763 17200 2764 17240
rect 2804 17200 2805 17240
rect 2763 17191 2805 17200
rect 9771 17240 9813 17249
rect 9771 17200 9772 17240
rect 9812 17200 9813 17240
rect 9771 17191 9813 17200
rect 11883 17240 11925 17249
rect 11883 17200 11884 17240
rect 11924 17200 11925 17240
rect 11883 17191 11925 17200
rect 13515 17240 13557 17249
rect 13515 17200 13516 17240
rect 13556 17200 13557 17240
rect 13515 17191 13557 17200
rect 16971 17240 17013 17249
rect 16971 17200 16972 17240
rect 17012 17200 17013 17240
rect 16971 17191 17013 17200
rect 4587 17156 4629 17165
rect 4587 17116 4588 17156
rect 4628 17116 4629 17156
rect 4587 17107 4629 17116
rect 6603 17156 6645 17165
rect 6603 17116 6604 17156
rect 6644 17116 6645 17156
rect 6603 17107 6645 17116
rect 18411 17156 18453 17165
rect 18411 17116 18412 17156
rect 18452 17116 18453 17156
rect 18411 17107 18453 17116
rect 1315 17072 1373 17073
rect 1315 17032 1324 17072
rect 1364 17032 1373 17072
rect 3139 17072 3197 17073
rect 1315 17031 1373 17032
rect 2563 17051 2621 17052
rect 2563 17011 2572 17051
rect 2612 17011 2621 17051
rect 3139 17032 3148 17072
rect 3188 17032 3197 17072
rect 3139 17031 3197 17032
rect 4387 17072 4445 17073
rect 4387 17032 4396 17072
rect 4436 17032 4445 17072
rect 4387 17031 4445 17032
rect 4875 17072 4917 17081
rect 4875 17032 4876 17072
rect 4916 17032 4917 17072
rect 4875 17023 4917 17032
rect 4971 17072 5013 17081
rect 4971 17032 4972 17072
rect 5012 17032 5013 17072
rect 4971 17023 5013 17032
rect 5355 17072 5397 17081
rect 5355 17032 5356 17072
rect 5396 17032 5397 17072
rect 5355 17023 5397 17032
rect 5923 17072 5981 17073
rect 5923 17032 5932 17072
rect 5972 17032 5981 17072
rect 5923 17031 5981 17032
rect 6411 17067 6453 17076
rect 6411 17027 6412 17067
rect 6452 17027 6453 17067
rect 8323 17072 8381 17073
rect 8323 17032 8332 17072
rect 8372 17032 8381 17072
rect 8323 17031 8381 17032
rect 9571 17072 9629 17073
rect 9571 17032 9580 17072
rect 9620 17032 9629 17072
rect 9571 17031 9629 17032
rect 10435 17072 10493 17073
rect 10435 17032 10444 17072
rect 10484 17032 10493 17072
rect 10435 17031 10493 17032
rect 12067 17072 12125 17073
rect 12067 17032 12076 17072
rect 12116 17032 12125 17072
rect 12067 17031 12125 17032
rect 13315 17072 13373 17073
rect 13315 17032 13324 17072
rect 13364 17032 13373 17072
rect 13315 17031 13373 17032
rect 15523 17072 15581 17073
rect 15523 17032 15532 17072
rect 15572 17032 15581 17072
rect 15523 17031 15581 17032
rect 16771 17072 16829 17073
rect 16771 17032 16780 17072
rect 16820 17032 16829 17072
rect 16771 17031 16829 17032
rect 18603 17067 18645 17076
rect 6411 17018 6453 17027
rect 11683 17030 11741 17031
rect 2563 17010 2621 17011
rect 5451 16988 5493 16997
rect 11683 16990 11692 17030
rect 11732 16990 11741 17030
rect 18603 17027 18604 17067
rect 18644 17027 18645 17067
rect 19075 17072 19133 17073
rect 19075 17032 19084 17072
rect 19124 17032 19133 17072
rect 19075 17031 19133 17032
rect 20043 17072 20085 17081
rect 20043 17032 20044 17072
rect 20084 17032 20085 17072
rect 18603 17018 18645 17027
rect 20043 17023 20085 17032
rect 20139 17053 20181 17062
rect 20139 17013 20140 17053
rect 20180 17013 20181 17053
rect 20139 17004 20181 17013
rect 11683 16989 11741 16990
rect 5451 16948 5452 16988
rect 5492 16948 5493 16988
rect 5451 16939 5493 16948
rect 18211 16988 18269 16989
rect 18211 16948 18220 16988
rect 18260 16948 18269 16988
rect 18211 16947 18269 16948
rect 19563 16988 19605 16997
rect 19563 16948 19564 16988
rect 19604 16948 19605 16988
rect 19563 16939 19605 16948
rect 19659 16988 19701 16997
rect 19659 16948 19660 16988
rect 19700 16948 19701 16988
rect 19659 16939 19701 16948
rect 2763 16820 2805 16829
rect 2763 16780 2764 16820
rect 2804 16780 2805 16820
rect 2763 16771 2805 16780
rect 18027 16820 18069 16829
rect 18027 16780 18028 16820
rect 18068 16780 18069 16820
rect 18027 16771 18069 16780
rect 1152 16652 20352 16676
rect 1152 16612 3688 16652
rect 3728 16612 3770 16652
rect 3810 16612 3852 16652
rect 3892 16612 3934 16652
rect 3974 16612 4016 16652
rect 4056 16612 18808 16652
rect 18848 16612 18890 16652
rect 18930 16612 18972 16652
rect 19012 16612 19054 16652
rect 19094 16612 19136 16652
rect 19176 16612 20352 16652
rect 1152 16588 20352 16612
rect 8811 16484 8853 16493
rect 8811 16444 8812 16484
rect 8852 16444 8853 16484
rect 8811 16435 8853 16444
rect 20235 16484 20277 16493
rect 20235 16444 20236 16484
rect 20276 16444 20277 16484
rect 20235 16435 20277 16444
rect 2955 16400 2997 16409
rect 2955 16360 2956 16400
rect 2996 16360 2997 16400
rect 2955 16351 2997 16360
rect 3907 16400 3965 16401
rect 3907 16360 3916 16400
rect 3956 16360 3965 16400
rect 3907 16359 3965 16360
rect 14187 16316 14229 16325
rect 14187 16276 14188 16316
rect 14228 16276 14229 16316
rect 14187 16267 14229 16276
rect 11163 16241 11205 16250
rect 15195 16241 15237 16250
rect 1507 16232 1565 16233
rect 1507 16192 1516 16232
rect 1556 16192 1565 16232
rect 1507 16191 1565 16192
rect 2755 16232 2813 16233
rect 2755 16192 2764 16232
rect 2804 16192 2813 16232
rect 2755 16191 2813 16192
rect 3235 16232 3293 16233
rect 3235 16192 3244 16232
rect 3284 16192 3293 16232
rect 3235 16191 3293 16192
rect 3531 16232 3573 16241
rect 3531 16192 3532 16232
rect 3572 16192 3573 16232
rect 3531 16183 3573 16192
rect 4291 16232 4349 16233
rect 4291 16192 4300 16232
rect 4340 16192 4349 16232
rect 4291 16191 4349 16192
rect 5539 16232 5597 16233
rect 5539 16192 5548 16232
rect 5588 16192 5597 16232
rect 5539 16191 5597 16192
rect 5931 16232 5973 16241
rect 5931 16192 5932 16232
rect 5972 16192 5973 16232
rect 5931 16183 5973 16192
rect 6027 16232 6069 16241
rect 6027 16192 6028 16232
rect 6068 16192 6069 16232
rect 6027 16183 6069 16192
rect 6499 16232 6557 16233
rect 6499 16192 6508 16232
rect 6548 16192 6557 16232
rect 6499 16191 6557 16192
rect 7363 16232 7421 16233
rect 7363 16192 7372 16232
rect 7412 16192 7421 16232
rect 7363 16191 7421 16192
rect 8611 16232 8669 16233
rect 8611 16192 8620 16232
rect 8660 16192 8669 16232
rect 8611 16191 8669 16192
rect 9579 16232 9621 16241
rect 9579 16192 9580 16232
rect 9620 16192 9621 16232
rect 9579 16183 9621 16192
rect 9675 16232 9717 16241
rect 9675 16192 9676 16232
rect 9716 16192 9717 16232
rect 9675 16183 9717 16192
rect 10059 16232 10101 16241
rect 10059 16192 10060 16232
rect 10100 16192 10101 16232
rect 10059 16183 10101 16192
rect 10155 16232 10197 16241
rect 10155 16192 10156 16232
rect 10196 16192 10197 16232
rect 10155 16183 10197 16192
rect 10627 16232 10685 16233
rect 10627 16192 10636 16232
rect 10676 16192 10685 16232
rect 11163 16201 11164 16241
rect 11204 16201 11205 16241
rect 11163 16192 11205 16201
rect 11875 16232 11933 16233
rect 11875 16192 11884 16232
rect 11924 16192 11933 16232
rect 10627 16191 10685 16192
rect 11875 16191 11933 16192
rect 13123 16232 13181 16233
rect 13123 16192 13132 16232
rect 13172 16192 13181 16232
rect 13123 16191 13181 16192
rect 13611 16232 13653 16241
rect 13611 16192 13612 16232
rect 13652 16192 13653 16232
rect 13611 16183 13653 16192
rect 13707 16232 13749 16241
rect 13707 16192 13708 16232
rect 13748 16192 13749 16232
rect 13707 16183 13749 16192
rect 14091 16232 14133 16241
rect 14091 16192 14092 16232
rect 14132 16192 14133 16232
rect 14091 16183 14133 16192
rect 14659 16232 14717 16233
rect 14659 16192 14668 16232
rect 14708 16192 14717 16232
rect 15195 16201 15196 16241
rect 15236 16201 15237 16241
rect 15195 16192 15237 16201
rect 15523 16232 15581 16233
rect 15523 16192 15532 16232
rect 15572 16192 15581 16232
rect 14659 16191 14717 16192
rect 15523 16191 15581 16192
rect 16771 16232 16829 16233
rect 16771 16192 16780 16232
rect 16820 16192 16829 16232
rect 16771 16191 16829 16192
rect 17347 16232 17405 16233
rect 17347 16192 17356 16232
rect 17396 16192 17405 16232
rect 17347 16191 17405 16192
rect 18595 16232 18653 16233
rect 18595 16192 18604 16232
rect 18644 16192 18653 16232
rect 18595 16191 18653 16192
rect 18787 16232 18845 16233
rect 18787 16192 18796 16232
rect 18836 16192 18845 16232
rect 18787 16191 18845 16192
rect 20035 16232 20093 16233
rect 20035 16192 20044 16232
rect 20084 16192 20093 16232
rect 20035 16191 20093 16192
rect 3627 16148 3669 16157
rect 3627 16108 3628 16148
rect 3668 16108 3669 16148
rect 3627 16099 3669 16108
rect 5739 16148 5781 16157
rect 5739 16108 5740 16148
rect 5780 16108 5781 16148
rect 5739 16099 5781 16108
rect 11307 16148 11349 16157
rect 11307 16108 11308 16148
rect 11348 16108 11349 16148
rect 11307 16099 11349 16108
rect 13323 16148 13365 16157
rect 13323 16108 13324 16148
rect 13364 16108 13365 16148
rect 13323 16099 13365 16108
rect 15339 16148 15381 16157
rect 15339 16108 15340 16148
rect 15380 16108 15381 16148
rect 15339 16099 15381 16108
rect 17163 16148 17205 16157
rect 17163 16108 17164 16148
rect 17204 16108 17205 16148
rect 17163 16099 17205 16108
rect 6211 16064 6269 16065
rect 6211 16024 6220 16064
rect 6260 16024 6269 16064
rect 6211 16023 6269 16024
rect 6411 16064 6453 16073
rect 6411 16024 6412 16064
rect 6452 16024 6453 16064
rect 6411 16015 6453 16024
rect 16971 16064 17013 16073
rect 16971 16024 16972 16064
rect 17012 16024 17013 16064
rect 16971 16015 17013 16024
rect 1152 15896 20452 15920
rect 1152 15856 4928 15896
rect 4968 15856 5010 15896
rect 5050 15856 5092 15896
rect 5132 15856 5174 15896
rect 5214 15856 5256 15896
rect 5296 15856 20048 15896
rect 20088 15856 20130 15896
rect 20170 15856 20212 15896
rect 20252 15856 20294 15896
rect 20334 15856 20376 15896
rect 20416 15856 20452 15896
rect 1152 15832 20452 15856
rect 3427 15728 3485 15729
rect 3427 15688 3436 15728
rect 3476 15688 3485 15728
rect 3427 15687 3485 15688
rect 5259 15728 5301 15737
rect 5259 15688 5260 15728
rect 5300 15688 5301 15728
rect 5259 15679 5301 15688
rect 8907 15728 8949 15737
rect 8907 15688 8908 15728
rect 8948 15688 8949 15728
rect 8907 15679 8949 15688
rect 11211 15728 11253 15737
rect 11211 15688 11212 15728
rect 11252 15688 11253 15728
rect 11211 15679 11253 15688
rect 15339 15728 15381 15737
rect 15339 15688 15340 15728
rect 15380 15688 15381 15728
rect 15339 15679 15381 15688
rect 6891 15644 6933 15653
rect 6891 15604 6892 15644
rect 6932 15604 6933 15644
rect 6891 15595 6933 15604
rect 18027 15644 18069 15653
rect 18027 15604 18028 15644
rect 18068 15604 18069 15644
rect 18027 15595 18069 15604
rect 7179 15580 7221 15589
rect 1219 15560 1277 15561
rect 1219 15520 1228 15560
rect 1268 15520 1277 15560
rect 1219 15519 1277 15520
rect 2467 15560 2525 15561
rect 2467 15520 2476 15560
rect 2516 15520 2525 15560
rect 2467 15519 2525 15520
rect 3147 15560 3189 15569
rect 3147 15520 3148 15560
rect 3188 15520 3189 15560
rect 3147 15511 3189 15520
rect 3243 15560 3285 15569
rect 3243 15520 3244 15560
rect 3284 15520 3285 15560
rect 3243 15511 3285 15520
rect 3339 15560 3381 15569
rect 3339 15520 3340 15560
rect 3380 15520 3381 15560
rect 3339 15511 3381 15520
rect 3811 15560 3869 15561
rect 3811 15520 3820 15560
rect 3860 15520 3869 15560
rect 3811 15519 3869 15520
rect 5059 15560 5117 15561
rect 5059 15520 5068 15560
rect 5108 15520 5117 15560
rect 5059 15519 5117 15520
rect 5443 15560 5501 15561
rect 5443 15520 5452 15560
rect 5492 15520 5501 15560
rect 5443 15519 5501 15520
rect 6691 15560 6749 15561
rect 6691 15520 6700 15560
rect 6740 15520 6749 15560
rect 7179 15540 7180 15580
rect 7220 15540 7221 15580
rect 7179 15531 7221 15540
rect 7275 15560 7317 15569
rect 6691 15519 6749 15520
rect 7275 15520 7276 15560
rect 7316 15520 7317 15560
rect 7275 15511 7317 15520
rect 7755 15560 7797 15569
rect 7755 15520 7756 15560
rect 7796 15520 7797 15560
rect 7755 15511 7797 15520
rect 8227 15560 8285 15561
rect 8227 15520 8236 15560
rect 8276 15520 8285 15560
rect 9763 15560 9821 15561
rect 8227 15519 8285 15520
rect 8715 15546 8757 15555
rect 8715 15506 8716 15546
rect 8756 15506 8757 15546
rect 9763 15520 9772 15560
rect 9812 15520 9821 15560
rect 9763 15519 9821 15520
rect 11011 15560 11069 15561
rect 11011 15520 11020 15560
rect 11060 15520 11069 15560
rect 11011 15519 11069 15520
rect 11587 15560 11645 15561
rect 11587 15520 11596 15560
rect 11636 15520 11645 15560
rect 11587 15519 11645 15520
rect 12835 15560 12893 15561
rect 12835 15520 12844 15560
rect 12884 15520 12893 15560
rect 12835 15519 12893 15520
rect 13891 15560 13949 15561
rect 13891 15520 13900 15560
rect 13940 15520 13949 15560
rect 13891 15519 13949 15520
rect 15139 15560 15197 15561
rect 15139 15520 15148 15560
rect 15188 15520 15197 15560
rect 15139 15519 15197 15520
rect 16299 15560 16341 15569
rect 16299 15520 16300 15560
rect 16340 15520 16341 15560
rect 16299 15511 16341 15520
rect 16395 15560 16437 15569
rect 16395 15520 16396 15560
rect 16436 15520 16437 15560
rect 16395 15511 16437 15520
rect 16779 15560 16821 15569
rect 16779 15520 16780 15560
rect 16820 15520 16821 15560
rect 16779 15511 16821 15520
rect 17347 15560 17405 15561
rect 17347 15520 17356 15560
rect 17396 15520 17405 15560
rect 17347 15519 17405 15520
rect 17835 15555 17877 15564
rect 17835 15515 17836 15555
rect 17876 15515 17877 15555
rect 18499 15560 18557 15561
rect 18499 15520 18508 15560
rect 18548 15520 18557 15560
rect 18499 15519 18557 15520
rect 19747 15560 19805 15561
rect 19747 15520 19756 15560
rect 19796 15520 19805 15560
rect 19747 15519 19805 15520
rect 17835 15506 17877 15515
rect 8715 15497 8757 15506
rect 7659 15476 7701 15485
rect 7659 15436 7660 15476
rect 7700 15436 7701 15476
rect 7659 15427 7701 15436
rect 16875 15476 16917 15485
rect 16875 15436 16876 15476
rect 16916 15436 16917 15476
rect 16875 15427 16917 15436
rect 2667 15308 2709 15317
rect 2667 15268 2668 15308
rect 2708 15268 2709 15308
rect 2667 15259 2709 15268
rect 5259 15308 5301 15317
rect 5259 15268 5260 15308
rect 5300 15268 5301 15308
rect 5259 15259 5301 15268
rect 11403 15308 11445 15317
rect 11403 15268 11404 15308
rect 11444 15268 11445 15308
rect 11403 15259 11445 15268
rect 19947 15308 19989 15317
rect 19947 15268 19948 15308
rect 19988 15268 19989 15308
rect 19947 15259 19989 15268
rect 1152 15140 20352 15164
rect 1152 15100 3688 15140
rect 3728 15100 3770 15140
rect 3810 15100 3852 15140
rect 3892 15100 3934 15140
rect 3974 15100 4016 15140
rect 4056 15100 18808 15140
rect 18848 15100 18890 15140
rect 18930 15100 18972 15140
rect 19012 15100 19054 15140
rect 19094 15100 19136 15140
rect 19176 15100 20352 15140
rect 1152 15076 20352 15100
rect 1515 14972 1557 14981
rect 1515 14932 1516 14972
rect 1556 14932 1557 14972
rect 1515 14923 1557 14932
rect 1899 14972 1941 14981
rect 1899 14932 1900 14972
rect 1940 14932 1941 14972
rect 1899 14923 1941 14932
rect 7947 14972 7989 14981
rect 7947 14932 7948 14972
rect 7988 14932 7989 14972
rect 7947 14923 7989 14932
rect 9579 14972 9621 14981
rect 9579 14932 9580 14972
rect 9620 14932 9621 14972
rect 9579 14923 9621 14932
rect 5347 14888 5405 14889
rect 5347 14848 5356 14888
rect 5396 14848 5405 14888
rect 5347 14847 5405 14848
rect 1699 14804 1757 14805
rect 1699 14764 1708 14804
rect 1748 14764 1757 14804
rect 1699 14763 1757 14764
rect 2083 14804 2141 14805
rect 2083 14764 2092 14804
rect 2132 14764 2141 14804
rect 2083 14763 2141 14764
rect 10731 14804 10773 14813
rect 10731 14764 10732 14804
rect 10772 14764 10773 14804
rect 10731 14755 10773 14764
rect 14091 14804 14133 14813
rect 14091 14764 14092 14804
rect 14132 14764 14133 14804
rect 14091 14755 14133 14764
rect 14187 14804 14229 14813
rect 14187 14764 14188 14804
rect 14228 14764 14229 14804
rect 14187 14755 14229 14764
rect 18891 14804 18933 14813
rect 18891 14764 18892 14804
rect 18932 14764 18933 14804
rect 18891 14755 18933 14764
rect 11691 14734 11733 14743
rect 2667 14720 2709 14729
rect 2667 14680 2668 14720
rect 2708 14680 2709 14720
rect 2667 14671 2709 14680
rect 2763 14720 2805 14729
rect 2763 14680 2764 14720
rect 2804 14680 2805 14720
rect 2763 14671 2805 14680
rect 3147 14720 3189 14729
rect 3147 14680 3148 14720
rect 3188 14680 3189 14720
rect 3147 14671 3189 14680
rect 3243 14720 3285 14729
rect 4203 14725 4245 14734
rect 3243 14680 3244 14720
rect 3284 14680 3285 14720
rect 3243 14671 3285 14680
rect 3715 14720 3773 14721
rect 3715 14680 3724 14720
rect 3764 14680 3773 14720
rect 3715 14679 3773 14680
rect 4203 14685 4204 14725
rect 4244 14685 4245 14725
rect 4203 14676 4245 14685
rect 5067 14720 5109 14729
rect 5067 14680 5068 14720
rect 5108 14680 5109 14720
rect 5067 14671 5109 14680
rect 5259 14720 5301 14729
rect 5259 14680 5260 14720
rect 5300 14680 5301 14720
rect 5259 14671 5301 14680
rect 5355 14720 5397 14729
rect 5355 14680 5356 14720
rect 5396 14680 5397 14720
rect 5355 14671 5397 14680
rect 5539 14720 5597 14721
rect 5539 14680 5548 14720
rect 5588 14680 5597 14720
rect 5539 14679 5597 14680
rect 5635 14720 5693 14721
rect 5635 14680 5644 14720
rect 5684 14680 5693 14720
rect 5635 14679 5693 14680
rect 5835 14720 5877 14729
rect 5835 14680 5836 14720
rect 5876 14680 5877 14720
rect 5835 14671 5877 14680
rect 5931 14720 5973 14729
rect 5931 14680 5932 14720
rect 5972 14680 5973 14720
rect 5931 14671 5973 14680
rect 6024 14720 6082 14721
rect 6024 14680 6033 14720
rect 6073 14680 6082 14720
rect 6024 14679 6082 14680
rect 6499 14720 6557 14721
rect 6499 14680 6508 14720
rect 6548 14680 6557 14720
rect 6499 14679 6557 14680
rect 7747 14720 7805 14721
rect 7747 14680 7756 14720
rect 7796 14680 7805 14720
rect 7747 14679 7805 14680
rect 8131 14720 8189 14721
rect 8131 14680 8140 14720
rect 8180 14680 8189 14720
rect 8131 14679 8189 14680
rect 9379 14720 9437 14721
rect 9379 14680 9388 14720
rect 9428 14680 9437 14720
rect 9379 14679 9437 14680
rect 10155 14720 10197 14729
rect 10155 14680 10156 14720
rect 10196 14680 10197 14720
rect 10155 14671 10197 14680
rect 10251 14720 10293 14729
rect 10251 14680 10252 14720
rect 10292 14680 10293 14720
rect 10251 14671 10293 14680
rect 10635 14720 10677 14729
rect 10635 14680 10636 14720
rect 10676 14680 10677 14720
rect 10635 14671 10677 14680
rect 11203 14720 11261 14721
rect 11203 14680 11212 14720
rect 11252 14680 11261 14720
rect 11691 14694 11692 14734
rect 11732 14694 11733 14734
rect 15195 14729 15237 14738
rect 19851 14734 19893 14743
rect 11691 14685 11733 14694
rect 13611 14720 13653 14729
rect 11203 14679 11261 14680
rect 13611 14680 13612 14720
rect 13652 14680 13653 14720
rect 13611 14671 13653 14680
rect 13707 14720 13749 14729
rect 13707 14680 13708 14720
rect 13748 14680 13749 14720
rect 13707 14671 13749 14680
rect 14659 14720 14717 14721
rect 14659 14680 14668 14720
rect 14708 14680 14717 14720
rect 15195 14689 15196 14729
rect 15236 14689 15237 14729
rect 15195 14680 15237 14689
rect 16099 14720 16157 14721
rect 16099 14680 16108 14720
rect 16148 14680 16157 14720
rect 14659 14679 14717 14680
rect 16099 14679 16157 14680
rect 17347 14720 17405 14721
rect 17347 14680 17356 14720
rect 17396 14680 17405 14720
rect 18411 14720 18453 14729
rect 17347 14679 17405 14680
rect 18315 14700 18357 14709
rect 18315 14660 18316 14700
rect 18356 14660 18357 14700
rect 18411 14680 18412 14720
rect 18452 14680 18453 14720
rect 18411 14671 18453 14680
rect 18795 14720 18837 14729
rect 18795 14680 18796 14720
rect 18836 14680 18837 14720
rect 18795 14671 18837 14680
rect 19363 14720 19421 14721
rect 19363 14680 19372 14720
rect 19412 14680 19421 14720
rect 19851 14694 19852 14734
rect 19892 14694 19893 14734
rect 19851 14685 19893 14694
rect 19363 14679 19421 14680
rect 18315 14651 18357 14660
rect 4395 14636 4437 14645
rect 4395 14596 4396 14636
rect 4436 14596 4437 14636
rect 4395 14587 4437 14596
rect 11883 14636 11925 14645
rect 11883 14596 11884 14636
rect 11924 14596 11925 14636
rect 11883 14587 11925 14596
rect 5731 14552 5789 14553
rect 5731 14512 5740 14552
rect 5780 14512 5789 14552
rect 5731 14511 5789 14512
rect 15339 14552 15381 14561
rect 15339 14512 15340 14552
rect 15380 14512 15381 14552
rect 15339 14503 15381 14512
rect 15915 14552 15957 14561
rect 15915 14512 15916 14552
rect 15956 14512 15957 14552
rect 15915 14503 15957 14512
rect 20043 14552 20085 14561
rect 20043 14512 20044 14552
rect 20084 14512 20085 14552
rect 20043 14503 20085 14512
rect 1152 14384 20452 14408
rect 1152 14344 4928 14384
rect 4968 14344 5010 14384
rect 5050 14344 5092 14384
rect 5132 14344 5174 14384
rect 5214 14344 5256 14384
rect 5296 14344 20048 14384
rect 20088 14344 20130 14384
rect 20170 14344 20212 14384
rect 20252 14344 20294 14384
rect 20334 14344 20376 14384
rect 20416 14344 20452 14384
rect 1152 14320 20452 14344
rect 1515 14216 1557 14225
rect 1515 14176 1516 14216
rect 1556 14176 1557 14216
rect 1515 14167 1557 14176
rect 2283 14216 2325 14225
rect 2283 14176 2284 14216
rect 2324 14176 2325 14216
rect 2283 14167 2325 14176
rect 4107 14216 4149 14225
rect 4107 14176 4108 14216
rect 4148 14176 4149 14216
rect 4107 14167 4149 14176
rect 11883 14216 11925 14225
rect 11883 14176 11884 14216
rect 11924 14176 11925 14216
rect 11883 14167 11925 14176
rect 13611 14216 13653 14225
rect 13611 14176 13612 14216
rect 13652 14176 13653 14216
rect 13611 14167 13653 14176
rect 15243 14216 15285 14225
rect 15243 14176 15244 14216
rect 15284 14176 15285 14216
rect 15243 14167 15285 14176
rect 17643 14216 17685 14225
rect 17643 14176 17644 14216
rect 17684 14176 17685 14216
rect 17643 14167 17685 14176
rect 6507 14132 6549 14141
rect 6507 14092 6508 14132
rect 6548 14092 6549 14132
rect 6507 14083 6549 14092
rect 8523 14132 8565 14141
rect 8523 14092 8524 14132
rect 8564 14092 8565 14132
rect 8523 14083 8565 14092
rect 15627 14132 15669 14141
rect 15627 14092 15628 14132
rect 15668 14092 15669 14132
rect 15627 14083 15669 14092
rect 2659 14048 2717 14049
rect 2659 14008 2668 14048
rect 2708 14008 2717 14048
rect 2659 14007 2717 14008
rect 3907 14048 3965 14049
rect 3907 14008 3916 14048
rect 3956 14008 3965 14048
rect 3907 14007 3965 14008
rect 5059 14048 5117 14049
rect 5059 14008 5068 14048
rect 5108 14008 5117 14048
rect 5059 14007 5117 14008
rect 6307 14048 6365 14049
rect 6307 14008 6316 14048
rect 6356 14008 6365 14048
rect 6307 14007 6365 14008
rect 6795 14048 6837 14057
rect 6795 14008 6796 14048
rect 6836 14008 6837 14048
rect 6795 13999 6837 14008
rect 6891 14048 6933 14057
rect 6891 14008 6892 14048
rect 6932 14008 6933 14048
rect 6891 13999 6933 14008
rect 7275 14048 7317 14057
rect 7275 14008 7276 14048
rect 7316 14008 7317 14048
rect 7275 13999 7317 14008
rect 7371 14048 7413 14057
rect 7371 14008 7372 14048
rect 7412 14008 7413 14048
rect 7371 13999 7413 14008
rect 7843 14048 7901 14049
rect 7843 14008 7852 14048
rect 7892 14008 7901 14048
rect 10155 14048 10197 14057
rect 7843 14007 7901 14008
rect 8379 14006 8421 14015
rect 8379 13966 8380 14006
rect 8420 13966 8421 14006
rect 10155 14008 10156 14048
rect 10196 14008 10197 14048
rect 10155 13999 10197 14008
rect 10251 14048 10293 14057
rect 10251 14008 10252 14048
rect 10292 14008 10293 14048
rect 10251 13999 10293 14008
rect 10635 14048 10677 14057
rect 10635 14008 10636 14048
rect 10676 14008 10677 14048
rect 10635 13999 10677 14008
rect 10731 14048 10773 14057
rect 10731 14008 10732 14048
rect 10772 14008 10773 14048
rect 10731 13999 10773 14008
rect 11203 14048 11261 14049
rect 11203 14008 11212 14048
rect 11252 14008 11261 14048
rect 11203 14007 11261 14008
rect 11691 14043 11733 14052
rect 11691 14003 11692 14043
rect 11732 14003 11733 14043
rect 12163 14048 12221 14049
rect 12163 14008 12172 14048
rect 12212 14008 12221 14048
rect 12163 14007 12221 14008
rect 13411 14048 13469 14049
rect 13411 14008 13420 14048
rect 13460 14008 13469 14048
rect 13411 14007 13469 14008
rect 13795 14048 13853 14049
rect 13795 14008 13804 14048
rect 13844 14008 13853 14048
rect 13795 14007 13853 14008
rect 15043 14048 15101 14049
rect 15043 14008 15052 14048
rect 15092 14008 15101 14048
rect 15043 14007 15101 14008
rect 15819 14043 15861 14052
rect 11691 13994 11733 14003
rect 15819 14003 15820 14043
rect 15860 14003 15861 14043
rect 16291 14048 16349 14049
rect 16291 14008 16300 14048
rect 16340 14008 16349 14048
rect 16291 14007 16349 14008
rect 16779 14048 16821 14057
rect 16779 14008 16780 14048
rect 16820 14008 16821 14048
rect 15819 13994 15861 14003
rect 16779 13999 16821 14008
rect 17259 14048 17301 14057
rect 17259 14008 17260 14048
rect 17300 14008 17301 14048
rect 17259 13999 17301 14008
rect 17355 14048 17397 14057
rect 17355 14008 17356 14048
rect 17396 14008 17397 14048
rect 17355 13999 17397 14008
rect 17827 14048 17885 14049
rect 17827 14008 17836 14048
rect 17876 14008 17885 14048
rect 17827 14007 17885 14008
rect 19075 14048 19133 14049
rect 19075 14008 19084 14048
rect 19124 14008 19133 14048
rect 19075 14007 19133 14008
rect 1699 13964 1757 13965
rect 1699 13924 1708 13964
rect 1748 13924 1757 13964
rect 1699 13923 1757 13924
rect 2083 13964 2141 13965
rect 2083 13924 2092 13964
rect 2132 13924 2141 13964
rect 2083 13923 2141 13924
rect 2467 13964 2525 13965
rect 2467 13924 2476 13964
rect 2516 13924 2525 13964
rect 8379 13957 8421 13966
rect 16875 13964 16917 13973
rect 2467 13923 2525 13924
rect 16875 13924 16876 13964
rect 16916 13924 16917 13964
rect 16875 13915 16917 13924
rect 1899 13880 1941 13889
rect 1899 13840 1900 13880
rect 1940 13840 1941 13880
rect 1899 13831 1941 13840
rect 1152 13628 20352 13652
rect 1152 13588 3688 13628
rect 3728 13588 3770 13628
rect 3810 13588 3852 13628
rect 3892 13588 3934 13628
rect 3974 13588 4016 13628
rect 4056 13588 18808 13628
rect 18848 13588 18890 13628
rect 18930 13588 18972 13628
rect 19012 13588 19054 13628
rect 19094 13588 19136 13628
rect 19176 13588 20352 13628
rect 1152 13564 20352 13588
rect 1323 13460 1365 13469
rect 1323 13420 1324 13460
rect 1364 13420 1365 13460
rect 1323 13411 1365 13420
rect 8427 13460 8469 13469
rect 8427 13420 8428 13460
rect 8468 13420 8469 13460
rect 8427 13411 8469 13420
rect 10155 13460 10197 13469
rect 10155 13420 10156 13460
rect 10196 13420 10197 13460
rect 10155 13411 10197 13420
rect 12363 13460 12405 13469
rect 12363 13420 12364 13460
rect 12404 13420 12405 13460
rect 12363 13411 12405 13420
rect 16395 13460 16437 13469
rect 16395 13420 16396 13460
rect 16436 13420 16437 13460
rect 16395 13411 16437 13420
rect 1507 13292 1565 13293
rect 1507 13252 1516 13292
rect 1556 13252 1565 13292
rect 1507 13251 1565 13252
rect 1891 13292 1949 13293
rect 1891 13252 1900 13292
rect 1940 13252 1949 13292
rect 1891 13251 1949 13252
rect 13515 13292 13557 13301
rect 13515 13252 13516 13292
rect 13556 13252 13557 13292
rect 13515 13243 13557 13252
rect 18891 13292 18933 13301
rect 18891 13252 18892 13292
rect 18932 13252 18933 13292
rect 18891 13243 18933 13252
rect 18987 13292 19029 13301
rect 18987 13252 18988 13292
rect 19028 13252 19029 13292
rect 18987 13243 19029 13252
rect 5403 13217 5445 13226
rect 14619 13217 14661 13226
rect 2083 13208 2141 13209
rect 2083 13168 2092 13208
rect 2132 13168 2141 13208
rect 2083 13167 2141 13168
rect 3331 13208 3389 13209
rect 3331 13168 3340 13208
rect 3380 13168 3389 13208
rect 3331 13167 3389 13168
rect 3819 13208 3861 13217
rect 3819 13168 3820 13208
rect 3860 13168 3861 13208
rect 3819 13159 3861 13168
rect 3915 13208 3957 13217
rect 3915 13168 3916 13208
rect 3956 13168 3957 13208
rect 3915 13159 3957 13168
rect 4299 13208 4341 13217
rect 4299 13168 4300 13208
rect 4340 13168 4341 13208
rect 4299 13159 4341 13168
rect 4395 13208 4437 13217
rect 4395 13168 4396 13208
rect 4436 13168 4437 13208
rect 4395 13159 4437 13168
rect 4867 13208 4925 13209
rect 4867 13168 4876 13208
rect 4916 13168 4925 13208
rect 5403 13177 5404 13217
rect 5444 13177 5445 13217
rect 5403 13168 5445 13177
rect 6979 13208 7037 13209
rect 6979 13168 6988 13208
rect 7028 13168 7037 13208
rect 4867 13167 4925 13168
rect 6979 13167 7037 13168
rect 8227 13208 8285 13209
rect 8227 13168 8236 13208
rect 8276 13168 8285 13208
rect 8227 13167 8285 13168
rect 8707 13208 8765 13209
rect 8707 13168 8716 13208
rect 8756 13168 8765 13208
rect 8707 13167 8765 13168
rect 9955 13208 10013 13209
rect 9955 13168 9964 13208
rect 10004 13168 10013 13208
rect 9955 13167 10013 13168
rect 10915 13208 10973 13209
rect 10915 13168 10924 13208
rect 10964 13168 10973 13208
rect 10915 13167 10973 13168
rect 12163 13208 12221 13209
rect 12163 13168 12172 13208
rect 12212 13168 12221 13208
rect 12163 13167 12221 13168
rect 13035 13208 13077 13217
rect 13035 13168 13036 13208
rect 13076 13168 13077 13208
rect 13035 13159 13077 13168
rect 13131 13208 13173 13217
rect 13131 13168 13132 13208
rect 13172 13168 13173 13208
rect 13131 13159 13173 13168
rect 13611 13208 13653 13217
rect 13611 13168 13612 13208
rect 13652 13168 13653 13208
rect 13611 13159 13653 13168
rect 14083 13208 14141 13209
rect 14083 13168 14092 13208
rect 14132 13168 14141 13208
rect 14619 13177 14620 13217
rect 14660 13177 14661 13217
rect 14619 13168 14661 13177
rect 14947 13208 15005 13209
rect 14947 13168 14956 13208
rect 14996 13168 15005 13208
rect 14083 13167 14141 13168
rect 14947 13167 15005 13168
rect 16195 13208 16253 13209
rect 16195 13168 16204 13208
rect 16244 13168 16253 13208
rect 16195 13167 16253 13168
rect 16675 13208 16733 13209
rect 16675 13168 16684 13208
rect 16724 13168 16733 13208
rect 16675 13167 16733 13168
rect 17923 13208 17981 13209
rect 17923 13168 17932 13208
rect 17972 13168 17981 13208
rect 17923 13167 17981 13168
rect 18411 13208 18453 13217
rect 18411 13168 18412 13208
rect 18452 13168 18453 13208
rect 18411 13159 18453 13168
rect 18507 13208 18549 13217
rect 19947 13213 19989 13222
rect 18507 13168 18508 13208
rect 18548 13168 18549 13208
rect 18507 13159 18549 13168
rect 19459 13208 19517 13209
rect 19459 13168 19468 13208
rect 19508 13168 19517 13208
rect 19459 13167 19517 13168
rect 19947 13173 19948 13213
rect 19988 13173 19989 13213
rect 19947 13164 19989 13173
rect 3531 13124 3573 13133
rect 3531 13084 3532 13124
rect 3572 13084 3573 13124
rect 3531 13075 3573 13084
rect 5547 13124 5589 13133
rect 5547 13084 5548 13124
rect 5588 13084 5589 13124
rect 5547 13075 5589 13084
rect 18123 13124 18165 13133
rect 18123 13084 18124 13124
rect 18164 13084 18165 13124
rect 18123 13075 18165 13084
rect 1707 13040 1749 13049
rect 1707 13000 1708 13040
rect 1748 13000 1749 13040
rect 1707 12991 1749 13000
rect 14763 13040 14805 13049
rect 14763 13000 14764 13040
rect 14804 13000 14805 13040
rect 14763 12991 14805 13000
rect 20139 13040 20181 13049
rect 20139 13000 20140 13040
rect 20180 13000 20181 13040
rect 20139 12991 20181 13000
rect 1152 12872 20452 12896
rect 1152 12832 4928 12872
rect 4968 12832 5010 12872
rect 5050 12832 5092 12872
rect 5132 12832 5174 12872
rect 5214 12832 5256 12872
rect 5296 12832 20048 12872
rect 20088 12832 20130 12872
rect 20170 12832 20212 12872
rect 20252 12832 20294 12872
rect 20334 12832 20376 12872
rect 20416 12832 20452 12872
rect 1152 12808 20452 12832
rect 5547 12704 5589 12713
rect 5547 12664 5548 12704
rect 5588 12664 5589 12704
rect 5547 12655 5589 12664
rect 10923 12704 10965 12713
rect 10923 12664 10924 12704
rect 10964 12664 10965 12704
rect 10923 12655 10965 12664
rect 13035 12704 13077 12713
rect 13035 12664 13036 12704
rect 13076 12664 13077 12704
rect 13035 12655 13077 12664
rect 14667 12704 14709 12713
rect 14667 12664 14668 12704
rect 14708 12664 14709 12704
rect 14667 12655 14709 12664
rect 20139 12704 20181 12713
rect 20139 12664 20140 12704
rect 20180 12664 20181 12704
rect 20139 12655 20181 12664
rect 8907 12620 8949 12629
rect 8907 12580 8908 12620
rect 8948 12580 8949 12620
rect 8907 12571 8949 12580
rect 17067 12620 17109 12629
rect 17067 12580 17068 12620
rect 17108 12580 17109 12620
rect 17067 12571 17109 12580
rect 2467 12536 2525 12537
rect 2467 12496 2476 12536
rect 2516 12496 2525 12536
rect 2467 12495 2525 12496
rect 3715 12536 3773 12537
rect 3715 12496 3724 12536
rect 3764 12496 3773 12536
rect 3715 12495 3773 12496
rect 4099 12536 4157 12537
rect 4099 12496 4108 12536
rect 4148 12496 4157 12536
rect 4099 12495 4157 12496
rect 5347 12536 5405 12537
rect 5347 12496 5356 12536
rect 5396 12496 5405 12536
rect 5347 12495 5405 12496
rect 8707 12536 8765 12537
rect 8707 12496 8716 12536
rect 8756 12496 8765 12536
rect 8707 12495 8765 12496
rect 9195 12536 9237 12545
rect 9195 12496 9196 12536
rect 9236 12496 9237 12536
rect 7459 12494 7517 12495
rect 7459 12454 7468 12494
rect 7508 12454 7517 12494
rect 9195 12487 9237 12496
rect 9291 12536 9333 12545
rect 9291 12496 9292 12536
rect 9332 12496 9333 12536
rect 9291 12487 9333 12496
rect 9675 12536 9717 12545
rect 9675 12496 9676 12536
rect 9716 12496 9717 12536
rect 9675 12487 9717 12496
rect 10243 12536 10301 12537
rect 10243 12496 10252 12536
rect 10292 12496 10301 12536
rect 11587 12536 11645 12537
rect 10243 12495 10301 12496
rect 10779 12526 10821 12535
rect 10779 12486 10780 12526
rect 10820 12486 10821 12526
rect 11587 12496 11596 12536
rect 11636 12496 11645 12536
rect 11587 12495 11645 12496
rect 12835 12536 12893 12537
rect 12835 12496 12844 12536
rect 12884 12496 12893 12536
rect 12835 12495 12893 12496
rect 13219 12536 13277 12537
rect 13219 12496 13228 12536
rect 13268 12496 13277 12536
rect 13219 12495 13277 12496
rect 14467 12536 14525 12537
rect 14467 12496 14476 12536
rect 14516 12496 14525 12536
rect 14467 12495 14525 12496
rect 15339 12536 15381 12545
rect 15339 12496 15340 12536
rect 15380 12496 15381 12536
rect 15339 12487 15381 12496
rect 15435 12536 15477 12545
rect 15435 12496 15436 12536
rect 15476 12496 15477 12536
rect 15435 12487 15477 12496
rect 15819 12536 15861 12545
rect 15819 12496 15820 12536
rect 15860 12496 15861 12536
rect 15819 12487 15861 12496
rect 15915 12536 15957 12545
rect 15915 12496 15916 12536
rect 15956 12496 15957 12536
rect 15915 12487 15957 12496
rect 16387 12536 16445 12537
rect 16387 12496 16396 12536
rect 16436 12496 16445 12536
rect 18691 12536 18749 12537
rect 16387 12495 16445 12496
rect 16875 12522 16917 12531
rect 10779 12477 10821 12486
rect 16875 12482 16876 12522
rect 16916 12482 16917 12522
rect 18691 12496 18700 12536
rect 18740 12496 18749 12536
rect 18691 12495 18749 12496
rect 19939 12536 19997 12537
rect 19939 12496 19948 12536
rect 19988 12496 19997 12536
rect 19939 12495 19997 12496
rect 16875 12473 16917 12482
rect 7459 12453 7517 12454
rect 1699 12452 1757 12453
rect 1699 12412 1708 12452
rect 1748 12412 1757 12452
rect 1699 12411 1757 12412
rect 2083 12452 2141 12453
rect 2083 12412 2092 12452
rect 2132 12412 2141 12452
rect 2083 12411 2141 12412
rect 9771 12452 9813 12461
rect 9771 12412 9772 12452
rect 9812 12412 9813 12452
rect 9771 12403 9813 12412
rect 1515 12368 1557 12377
rect 1515 12328 1516 12368
rect 1556 12328 1557 12368
rect 1515 12319 1557 12328
rect 1899 12368 1941 12377
rect 1899 12328 1900 12368
rect 1940 12328 1941 12368
rect 1899 12319 1941 12328
rect 3915 12284 3957 12293
rect 3915 12244 3916 12284
rect 3956 12244 3957 12284
rect 3915 12235 3957 12244
rect 1152 12116 20352 12140
rect 1152 12076 3688 12116
rect 3728 12076 3770 12116
rect 3810 12076 3852 12116
rect 3892 12076 3934 12116
rect 3974 12076 4016 12116
rect 4056 12076 18808 12116
rect 18848 12076 18890 12116
rect 18930 12076 18972 12116
rect 19012 12076 19054 12116
rect 19094 12076 19136 12116
rect 19176 12076 20352 12116
rect 1152 12052 20352 12076
rect 1515 11948 1557 11957
rect 1515 11908 1516 11948
rect 1556 11908 1557 11948
rect 1515 11899 1557 11908
rect 1899 11948 1941 11957
rect 1899 11908 1900 11948
rect 1940 11908 1941 11948
rect 1899 11899 1941 11908
rect 10155 11948 10197 11957
rect 10155 11908 10156 11948
rect 10196 11908 10197 11948
rect 10155 11899 10197 11908
rect 15339 11948 15381 11957
rect 15339 11908 15340 11948
rect 15380 11908 15381 11948
rect 15339 11899 15381 11908
rect 17259 11948 17301 11957
rect 17259 11908 17260 11948
rect 17300 11908 17301 11948
rect 17259 11899 17301 11908
rect 1699 11780 1757 11781
rect 1699 11740 1708 11780
rect 1748 11740 1757 11780
rect 1699 11739 1757 11740
rect 2083 11780 2141 11781
rect 2083 11740 2092 11780
rect 2132 11740 2141 11780
rect 2083 11739 2141 11740
rect 3147 11780 3189 11789
rect 3147 11740 3148 11780
rect 3188 11740 3189 11780
rect 3147 11731 3189 11740
rect 7275 11780 7317 11789
rect 7275 11740 7276 11780
rect 7316 11740 7317 11780
rect 7275 11731 7317 11740
rect 18891 11780 18933 11789
rect 18891 11740 18892 11780
rect 18932 11740 18933 11780
rect 9955 11738 10013 11739
rect 4203 11710 4245 11719
rect 2667 11696 2709 11705
rect 2667 11656 2668 11696
rect 2708 11656 2709 11696
rect 2667 11647 2709 11656
rect 2763 11696 2805 11705
rect 2763 11656 2764 11696
rect 2804 11656 2805 11696
rect 2763 11647 2805 11656
rect 3243 11696 3285 11705
rect 3243 11656 3244 11696
rect 3284 11656 3285 11696
rect 3243 11647 3285 11656
rect 3715 11696 3773 11697
rect 3715 11656 3724 11696
rect 3764 11656 3773 11696
rect 4203 11670 4204 11710
rect 4244 11670 4245 11710
rect 4203 11661 4245 11670
rect 5059 11696 5117 11697
rect 3715 11655 3773 11656
rect 5059 11656 5068 11696
rect 5108 11656 5117 11696
rect 5059 11655 5117 11656
rect 6307 11696 6365 11697
rect 6307 11656 6316 11696
rect 6356 11656 6365 11696
rect 6307 11655 6365 11656
rect 6795 11696 6837 11705
rect 6795 11656 6796 11696
rect 6836 11656 6837 11696
rect 6795 11647 6837 11656
rect 6891 11696 6933 11705
rect 6891 11656 6892 11696
rect 6932 11656 6933 11696
rect 6891 11647 6933 11656
rect 7371 11696 7413 11705
rect 8331 11701 8373 11710
rect 7371 11656 7372 11696
rect 7412 11656 7413 11696
rect 7371 11647 7413 11656
rect 7843 11696 7901 11697
rect 7843 11656 7852 11696
rect 7892 11656 7901 11696
rect 7843 11655 7901 11656
rect 8331 11661 8332 11701
rect 8372 11661 8373 11701
rect 9955 11698 9964 11738
rect 10004 11698 10013 11738
rect 18891 11731 18933 11740
rect 18987 11780 19029 11789
rect 18987 11740 18988 11780
rect 19028 11740 19029 11780
rect 18987 11731 19029 11740
rect 9955 11697 10013 11698
rect 8331 11652 8373 11661
rect 8707 11696 8765 11697
rect 8707 11656 8716 11696
rect 8756 11656 8765 11696
rect 8707 11655 8765 11656
rect 10339 11696 10397 11697
rect 10339 11656 10348 11696
rect 10388 11656 10397 11696
rect 10339 11655 10397 11656
rect 11587 11696 11645 11697
rect 11587 11656 11596 11696
rect 11636 11656 11645 11696
rect 11587 11655 11645 11656
rect 13891 11696 13949 11697
rect 13891 11656 13900 11696
rect 13940 11656 13949 11696
rect 13891 11655 13949 11656
rect 15139 11696 15197 11697
rect 15139 11656 15148 11696
rect 15188 11656 15197 11696
rect 15139 11655 15197 11656
rect 15811 11696 15869 11697
rect 15811 11656 15820 11696
rect 15860 11656 15869 11696
rect 15811 11655 15869 11656
rect 17059 11696 17117 11697
rect 17059 11656 17068 11696
rect 17108 11656 17117 11696
rect 17059 11655 17117 11656
rect 18411 11696 18453 11705
rect 18411 11656 18412 11696
rect 18452 11656 18453 11696
rect 18411 11647 18453 11656
rect 18507 11696 18549 11705
rect 19947 11701 19989 11710
rect 18507 11656 18508 11696
rect 18548 11656 18549 11696
rect 18507 11647 18549 11656
rect 19459 11696 19517 11697
rect 19459 11656 19468 11696
rect 19508 11656 19517 11696
rect 19459 11655 19517 11656
rect 19947 11661 19948 11701
rect 19988 11661 19989 11701
rect 19947 11652 19989 11661
rect 6507 11612 6549 11621
rect 6507 11572 6508 11612
rect 6548 11572 6549 11612
rect 6507 11563 6549 11572
rect 8523 11612 8565 11621
rect 8523 11572 8524 11612
rect 8564 11572 8565 11612
rect 8523 11563 8565 11572
rect 4395 11528 4437 11537
rect 4395 11488 4396 11528
rect 4436 11488 4437 11528
rect 4395 11479 4437 11488
rect 11787 11528 11829 11537
rect 11787 11488 11788 11528
rect 11828 11488 11829 11528
rect 11787 11479 11829 11488
rect 20139 11528 20181 11537
rect 20139 11488 20140 11528
rect 20180 11488 20181 11528
rect 20139 11479 20181 11488
rect 1152 11360 20452 11384
rect 1152 11320 4928 11360
rect 4968 11320 5010 11360
rect 5050 11320 5092 11360
rect 5132 11320 5174 11360
rect 5214 11320 5256 11360
rect 5296 11320 20048 11360
rect 20088 11320 20130 11360
rect 20170 11320 20212 11360
rect 20252 11320 20294 11360
rect 20334 11320 20376 11360
rect 20416 11320 20452 11360
rect 1152 11296 20452 11320
rect 2667 11192 2709 11201
rect 2667 11152 2668 11192
rect 2708 11152 2709 11192
rect 2667 11143 2709 11152
rect 7371 11192 7413 11201
rect 7371 11152 7372 11192
rect 7412 11152 7413 11192
rect 7371 11143 7413 11152
rect 9003 11192 9045 11201
rect 9003 11152 9004 11192
rect 9044 11152 9045 11192
rect 9003 11143 9045 11152
rect 11019 11192 11061 11201
rect 11019 11152 11020 11192
rect 11060 11152 11061 11192
rect 11019 11143 11061 11152
rect 16011 11192 16053 11201
rect 16011 11152 16012 11192
rect 16052 11152 16053 11192
rect 16011 11143 16053 11152
rect 18507 11192 18549 11201
rect 18507 11152 18508 11192
rect 18548 11152 18549 11192
rect 18507 11143 18549 11152
rect 20139 11192 20181 11201
rect 20139 11152 20140 11192
rect 20180 11152 20181 11192
rect 20139 11143 20181 11152
rect 5355 11108 5397 11117
rect 5355 11068 5356 11108
rect 5396 11068 5397 11108
rect 5355 11059 5397 11068
rect 1219 11024 1277 11025
rect 1219 10984 1228 11024
rect 1268 10984 1277 11024
rect 1219 10983 1277 10984
rect 2467 11024 2525 11025
rect 2467 10984 2476 11024
rect 2516 10984 2525 11024
rect 2467 10983 2525 10984
rect 3907 11024 3965 11025
rect 3907 10984 3916 11024
rect 3956 10984 3965 11024
rect 3907 10983 3965 10984
rect 5155 11024 5213 11025
rect 5155 10984 5164 11024
rect 5204 10984 5213 11024
rect 5155 10983 5213 10984
rect 5643 11024 5685 11033
rect 5643 10984 5644 11024
rect 5684 10984 5685 11024
rect 5643 10975 5685 10984
rect 5739 11024 5781 11033
rect 5739 10984 5740 11024
rect 5780 10984 5781 11024
rect 5739 10975 5781 10984
rect 6219 11024 6261 11033
rect 6219 10984 6220 11024
rect 6260 10984 6261 11024
rect 6219 10975 6261 10984
rect 6691 11024 6749 11025
rect 6691 10984 6700 11024
rect 6740 10984 6749 11024
rect 7555 11024 7613 11025
rect 6691 10983 6749 10984
rect 7179 11010 7221 11019
rect 7179 10970 7180 11010
rect 7220 10970 7221 11010
rect 7555 10984 7564 11024
rect 7604 10984 7613 11024
rect 7555 10983 7613 10984
rect 8803 11024 8861 11025
rect 8803 10984 8812 11024
rect 8852 10984 8861 11024
rect 8803 10983 8861 10984
rect 9571 11024 9629 11025
rect 9571 10984 9580 11024
rect 9620 10984 9629 11024
rect 9571 10983 9629 10984
rect 10819 11024 10877 11025
rect 10819 10984 10828 11024
rect 10868 10984 10877 11024
rect 10819 10983 10877 10984
rect 11587 11024 11645 11025
rect 11587 10984 11596 11024
rect 11636 10984 11645 11024
rect 11587 10983 11645 10984
rect 12835 11024 12893 11025
rect 12835 10984 12844 11024
rect 12884 10984 12893 11024
rect 12835 10983 12893 10984
rect 14283 11024 14325 11033
rect 14283 10984 14284 11024
rect 14324 10984 14325 11024
rect 14283 10975 14325 10984
rect 14379 11024 14421 11033
rect 14379 10984 14380 11024
rect 14420 10984 14421 11024
rect 14379 10975 14421 10984
rect 14859 11024 14901 11033
rect 14859 10984 14860 11024
rect 14900 10984 14901 11024
rect 14859 10975 14901 10984
rect 15331 11024 15389 11025
rect 15331 10984 15340 11024
rect 15380 10984 15389 11024
rect 17059 11024 17117 11025
rect 15331 10983 15389 10984
rect 15819 11010 15861 11019
rect 7179 10961 7221 10970
rect 15819 10970 15820 11010
rect 15860 10970 15861 11010
rect 17059 10984 17068 11024
rect 17108 10984 17117 11024
rect 17059 10983 17117 10984
rect 18307 11024 18365 11025
rect 18307 10984 18316 11024
rect 18356 10984 18365 11024
rect 18307 10983 18365 10984
rect 18691 11024 18749 11025
rect 18691 10984 18700 11024
rect 18740 10984 18749 11024
rect 18691 10983 18749 10984
rect 19939 11024 19997 11025
rect 19939 10984 19948 11024
rect 19988 10984 19997 11024
rect 19939 10983 19997 10984
rect 15819 10961 15861 10970
rect 3043 10940 3101 10941
rect 3043 10900 3052 10940
rect 3092 10900 3101 10940
rect 3043 10899 3101 10900
rect 6123 10940 6165 10949
rect 6123 10900 6124 10940
rect 6164 10900 6165 10940
rect 6123 10891 6165 10900
rect 14763 10940 14805 10949
rect 14763 10900 14764 10940
rect 14804 10900 14805 10940
rect 14763 10891 14805 10900
rect 2859 10772 2901 10781
rect 2859 10732 2860 10772
rect 2900 10732 2901 10772
rect 2859 10723 2901 10732
rect 13035 10772 13077 10781
rect 13035 10732 13036 10772
rect 13076 10732 13077 10772
rect 13035 10723 13077 10732
rect 1152 10604 20352 10628
rect 1152 10564 3688 10604
rect 3728 10564 3770 10604
rect 3810 10564 3852 10604
rect 3892 10564 3934 10604
rect 3974 10564 4016 10604
rect 4056 10564 18808 10604
rect 18848 10564 18890 10604
rect 18930 10564 18972 10604
rect 19012 10564 19054 10604
rect 19094 10564 19136 10604
rect 19176 10564 20352 10604
rect 1152 10540 20352 10564
rect 6987 10352 7029 10361
rect 6987 10312 6988 10352
rect 7028 10312 7029 10352
rect 6987 10303 7029 10312
rect 8619 10352 8661 10361
rect 8619 10312 8620 10352
rect 8660 10312 8661 10352
rect 8619 10303 8661 10312
rect 17451 10352 17493 10361
rect 17451 10312 17452 10352
rect 17492 10312 17493 10352
rect 17451 10303 17493 10312
rect 3819 10268 3861 10277
rect 3819 10228 3820 10268
rect 3860 10228 3861 10268
rect 3819 10219 3861 10228
rect 9387 10268 9429 10277
rect 9387 10228 9388 10268
rect 9428 10228 9429 10268
rect 9387 10219 9429 10228
rect 11691 10268 11733 10277
rect 11691 10228 11692 10268
rect 11732 10228 11733 10268
rect 16011 10268 16053 10277
rect 11691 10219 11733 10228
rect 12795 10226 12837 10235
rect 16011 10228 16012 10268
rect 16052 10228 16053 10268
rect 1507 10184 1565 10185
rect 1507 10144 1516 10184
rect 1556 10144 1565 10184
rect 1507 10143 1565 10144
rect 2755 10184 2813 10185
rect 2755 10144 2764 10184
rect 2804 10144 2813 10184
rect 2755 10143 2813 10144
rect 3243 10184 3285 10193
rect 3243 10144 3244 10184
rect 3284 10144 3285 10184
rect 3243 10135 3285 10144
rect 3339 10184 3381 10193
rect 3339 10144 3340 10184
rect 3380 10144 3381 10184
rect 3339 10135 3381 10144
rect 3723 10184 3765 10193
rect 4779 10189 4821 10198
rect 10491 10193 10533 10202
rect 3723 10144 3724 10184
rect 3764 10144 3765 10184
rect 3723 10135 3765 10144
rect 4291 10184 4349 10185
rect 4291 10144 4300 10184
rect 4340 10144 4349 10184
rect 4291 10143 4349 10144
rect 4779 10149 4780 10189
rect 4820 10149 4821 10189
rect 4779 10140 4821 10149
rect 5539 10184 5597 10185
rect 5539 10144 5548 10184
rect 5588 10144 5597 10184
rect 5539 10143 5597 10144
rect 6787 10184 6845 10185
rect 6787 10144 6796 10184
rect 6836 10144 6845 10184
rect 6787 10143 6845 10144
rect 7171 10184 7229 10185
rect 7171 10144 7180 10184
rect 7220 10144 7229 10184
rect 7171 10143 7229 10144
rect 8419 10184 8477 10185
rect 8419 10144 8428 10184
rect 8468 10144 8477 10184
rect 8419 10143 8477 10144
rect 8907 10184 8949 10193
rect 8907 10144 8908 10184
rect 8948 10144 8949 10184
rect 8907 10135 8949 10144
rect 9003 10184 9045 10193
rect 9003 10144 9004 10184
rect 9044 10144 9045 10184
rect 9003 10135 9045 10144
rect 9483 10184 9525 10193
rect 9483 10144 9484 10184
rect 9524 10144 9525 10184
rect 9483 10135 9525 10144
rect 9955 10184 10013 10185
rect 9955 10144 9964 10184
rect 10004 10144 10013 10184
rect 10491 10153 10492 10193
rect 10532 10153 10533 10193
rect 10491 10144 10533 10153
rect 11211 10184 11253 10193
rect 11211 10144 11212 10184
rect 11252 10144 11253 10184
rect 9955 10143 10013 10144
rect 11211 10135 11253 10144
rect 11307 10184 11349 10193
rect 11307 10144 11308 10184
rect 11348 10144 11349 10184
rect 11307 10135 11349 10144
rect 11787 10184 11829 10193
rect 12795 10186 12796 10226
rect 12836 10186 12837 10226
rect 11787 10144 11788 10184
rect 11828 10144 11829 10184
rect 11787 10135 11829 10144
rect 12259 10184 12317 10185
rect 12259 10144 12268 10184
rect 12308 10144 12317 10184
rect 12795 10177 12837 10186
rect 14371 10226 14429 10227
rect 14371 10186 14380 10226
rect 14420 10186 14429 10226
rect 16011 10219 16053 10228
rect 16107 10268 16149 10277
rect 16107 10228 16108 10268
rect 16148 10228 16149 10268
rect 16107 10219 16149 10228
rect 17635 10268 17693 10269
rect 17635 10228 17644 10268
rect 17684 10228 17693 10268
rect 17635 10227 17693 10228
rect 19179 10268 19221 10277
rect 19179 10228 19180 10268
rect 19220 10228 19221 10268
rect 19179 10219 19221 10228
rect 19275 10268 19317 10277
rect 19275 10228 19276 10268
rect 19316 10228 19317 10268
rect 19275 10219 19317 10228
rect 17115 10193 17157 10202
rect 14371 10185 14429 10186
rect 13123 10184 13181 10185
rect 12259 10143 12317 10144
rect 13123 10144 13132 10184
rect 13172 10144 13181 10184
rect 13123 10143 13181 10144
rect 15531 10184 15573 10193
rect 15531 10144 15532 10184
rect 15572 10144 15573 10184
rect 15531 10135 15573 10144
rect 15627 10184 15669 10193
rect 15627 10144 15628 10184
rect 15668 10144 15669 10184
rect 15627 10135 15669 10144
rect 16579 10184 16637 10185
rect 16579 10144 16588 10184
rect 16628 10144 16637 10184
rect 17115 10153 17116 10193
rect 17156 10153 17157 10193
rect 17115 10144 17157 10153
rect 18219 10189 18261 10198
rect 18219 10149 18220 10189
rect 18260 10149 18261 10189
rect 16579 10143 16637 10144
rect 18219 10140 18261 10149
rect 18691 10184 18749 10185
rect 18691 10144 18700 10184
rect 18740 10144 18749 10184
rect 18691 10143 18749 10144
rect 19659 10184 19701 10193
rect 19659 10144 19660 10184
rect 19700 10144 19701 10184
rect 19659 10135 19701 10144
rect 19755 10184 19797 10193
rect 19755 10144 19756 10184
rect 19796 10144 19797 10184
rect 19755 10135 19797 10144
rect 2955 10100 2997 10109
rect 2955 10060 2956 10100
rect 2996 10060 2997 10100
rect 2955 10051 2997 10060
rect 4971 10100 5013 10109
rect 4971 10060 4972 10100
rect 5012 10060 5013 10100
rect 4971 10051 5013 10060
rect 12939 10100 12981 10109
rect 12939 10060 12940 10100
rect 12980 10060 12981 10100
rect 12939 10051 12981 10060
rect 14571 10100 14613 10109
rect 14571 10060 14572 10100
rect 14612 10060 14613 10100
rect 14571 10051 14613 10060
rect 17259 10100 17301 10109
rect 17259 10060 17260 10100
rect 17300 10060 17301 10100
rect 17259 10051 17301 10060
rect 18027 10100 18069 10109
rect 18027 10060 18028 10100
rect 18068 10060 18069 10100
rect 18027 10051 18069 10060
rect 10635 10016 10677 10025
rect 10635 9976 10636 10016
rect 10676 9976 10677 10016
rect 10635 9967 10677 9976
rect 1152 9848 20452 9872
rect 1152 9808 4928 9848
rect 4968 9808 5010 9848
rect 5050 9808 5092 9848
rect 5132 9808 5174 9848
rect 5214 9808 5256 9848
rect 5296 9808 20048 9848
rect 20088 9808 20130 9848
rect 20170 9808 20212 9848
rect 20252 9808 20294 9848
rect 20334 9808 20376 9848
rect 20416 9808 20452 9848
rect 1152 9784 20452 9808
rect 1515 9680 1557 9689
rect 1515 9640 1516 9680
rect 1556 9640 1557 9680
rect 1515 9631 1557 9640
rect 3339 9680 3381 9689
rect 3339 9640 3340 9680
rect 3380 9640 3381 9680
rect 3339 9631 3381 9640
rect 7179 9680 7221 9689
rect 7179 9640 7180 9680
rect 7220 9640 7221 9680
rect 7179 9631 7221 9640
rect 10635 9680 10677 9689
rect 10635 9640 10636 9680
rect 10676 9640 10677 9680
rect 10635 9631 10677 9640
rect 15723 9680 15765 9689
rect 15723 9640 15724 9680
rect 15764 9640 15765 9680
rect 15723 9631 15765 9640
rect 17451 9680 17493 9689
rect 17451 9640 17452 9680
rect 17492 9640 17493 9680
rect 17451 9631 17493 9640
rect 19083 9680 19125 9689
rect 19083 9640 19084 9680
rect 19124 9640 19125 9680
rect 19083 9631 19125 9640
rect 5451 9596 5493 9605
rect 5451 9556 5452 9596
rect 5492 9556 5493 9596
rect 5451 9547 5493 9556
rect 12747 9596 12789 9605
rect 12747 9556 12748 9596
rect 12788 9556 12789 9596
rect 12747 9547 12789 9556
rect 1891 9512 1949 9513
rect 1891 9472 1900 9512
rect 1940 9472 1949 9512
rect 1891 9471 1949 9472
rect 3139 9512 3197 9513
rect 3139 9472 3148 9512
rect 3188 9472 3197 9512
rect 3139 9471 3197 9472
rect 3723 9512 3765 9521
rect 3723 9472 3724 9512
rect 3764 9472 3765 9512
rect 3723 9463 3765 9472
rect 3819 9512 3861 9521
rect 3819 9472 3820 9512
rect 3860 9472 3861 9512
rect 3819 9463 3861 9472
rect 4771 9512 4829 9513
rect 4771 9472 4780 9512
rect 4820 9472 4829 9512
rect 7843 9512 7901 9513
rect 7371 9498 7413 9507
rect 4771 9471 4829 9472
rect 5307 9470 5349 9479
rect 1699 9428 1757 9429
rect 1699 9388 1708 9428
rect 1748 9388 1757 9428
rect 1699 9387 1757 9388
rect 4203 9428 4245 9437
rect 4203 9388 4204 9428
rect 4244 9388 4245 9428
rect 4203 9379 4245 9388
rect 4299 9428 4341 9437
rect 4299 9388 4300 9428
rect 4340 9388 4341 9428
rect 5307 9430 5308 9470
rect 5348 9430 5349 9470
rect 7371 9458 7372 9498
rect 7412 9458 7413 9498
rect 7843 9472 7852 9512
rect 7892 9472 7901 9512
rect 7843 9471 7901 9472
rect 8331 9512 8373 9521
rect 8331 9472 8332 9512
rect 8372 9472 8373 9512
rect 8331 9463 8373 9472
rect 8427 9512 8469 9521
rect 8427 9472 8428 9512
rect 8468 9472 8469 9512
rect 8427 9463 8469 9472
rect 8811 9512 8853 9521
rect 8811 9472 8812 9512
rect 8852 9472 8853 9512
rect 8811 9463 8853 9472
rect 8907 9512 8949 9521
rect 8907 9472 8908 9512
rect 8948 9472 8949 9512
rect 8907 9463 8949 9472
rect 9187 9512 9245 9513
rect 9187 9472 9196 9512
rect 9236 9472 9245 9512
rect 9187 9471 9245 9472
rect 10435 9512 10493 9513
rect 10435 9472 10444 9512
rect 10484 9472 10493 9512
rect 10435 9471 10493 9472
rect 11019 9512 11061 9521
rect 11019 9472 11020 9512
rect 11060 9472 11061 9512
rect 11019 9463 11061 9472
rect 11115 9512 11157 9521
rect 11115 9472 11116 9512
rect 11156 9472 11157 9512
rect 11115 9463 11157 9472
rect 11595 9512 11637 9521
rect 11595 9472 11596 9512
rect 11636 9472 11637 9512
rect 11595 9463 11637 9472
rect 12067 9512 12125 9513
rect 12067 9472 12076 9512
rect 12116 9472 12125 9512
rect 14275 9512 14333 9513
rect 12067 9471 12125 9472
rect 12555 9498 12597 9507
rect 7371 9449 7413 9458
rect 12555 9458 12556 9498
rect 12596 9458 12597 9498
rect 14275 9472 14284 9512
rect 14324 9472 14333 9512
rect 14275 9471 14333 9472
rect 15523 9512 15581 9513
rect 15523 9472 15532 9512
rect 15572 9472 15581 9512
rect 15523 9471 15581 9472
rect 16003 9512 16061 9513
rect 16003 9472 16012 9512
rect 16052 9472 16061 9512
rect 16003 9471 16061 9472
rect 17251 9512 17309 9513
rect 17251 9472 17260 9512
rect 17300 9472 17309 9512
rect 17251 9471 17309 9472
rect 17635 9512 17693 9513
rect 17635 9472 17644 9512
rect 17684 9472 17693 9512
rect 17635 9471 17693 9472
rect 18883 9512 18941 9513
rect 18883 9472 18892 9512
rect 18932 9472 18941 9512
rect 18883 9471 18941 9472
rect 12555 9449 12597 9458
rect 5307 9421 5349 9430
rect 11499 9428 11541 9437
rect 4299 9379 4341 9388
rect 11499 9388 11500 9428
rect 11540 9388 11541 9428
rect 11499 9379 11541 9388
rect 19555 9428 19613 9429
rect 19555 9388 19564 9428
rect 19604 9388 19613 9428
rect 19555 9387 19613 9388
rect 19371 9260 19413 9269
rect 19371 9220 19372 9260
rect 19412 9220 19413 9260
rect 19371 9211 19413 9220
rect 1152 9092 20352 9116
rect 1152 9052 3688 9092
rect 3728 9052 3770 9092
rect 3810 9052 3852 9092
rect 3892 9052 3934 9092
rect 3974 9052 4016 9092
rect 4056 9052 18808 9092
rect 18848 9052 18890 9092
rect 18930 9052 18972 9092
rect 19012 9052 19054 9092
rect 19094 9052 19136 9092
rect 19176 9052 20352 9092
rect 1152 9028 20352 9052
rect 7275 8924 7317 8933
rect 7275 8884 7276 8924
rect 7316 8884 7317 8924
rect 7275 8875 7317 8884
rect 11211 8924 11253 8933
rect 11211 8884 11212 8924
rect 11252 8884 11253 8924
rect 11211 8875 11253 8884
rect 20139 8924 20181 8933
rect 20139 8884 20140 8924
rect 20180 8884 20181 8924
rect 20139 8875 20181 8884
rect 1515 8840 1557 8849
rect 1515 8800 1516 8840
rect 1556 8800 1557 8840
rect 1515 8791 1557 8800
rect 1899 8840 1941 8849
rect 1899 8800 1900 8840
rect 1940 8800 1941 8840
rect 1899 8791 1941 8800
rect 2283 8840 2325 8849
rect 2283 8800 2284 8840
rect 2324 8800 2325 8840
rect 2283 8791 2325 8800
rect 2667 8840 2709 8849
rect 2667 8800 2668 8840
rect 2708 8800 2709 8840
rect 2667 8791 2709 8800
rect 4971 8840 5013 8849
rect 4971 8800 4972 8840
rect 5012 8800 5013 8840
rect 4971 8791 5013 8800
rect 7083 8840 7125 8849
rect 7083 8800 7084 8840
rect 7124 8800 7125 8840
rect 7083 8791 7125 8800
rect 13035 8840 13077 8849
rect 13035 8800 13036 8840
rect 13076 8800 13077 8840
rect 13035 8791 13077 8800
rect 14859 8840 14901 8849
rect 14859 8800 14860 8840
rect 14900 8800 14901 8840
rect 14859 8791 14901 8800
rect 17067 8840 17109 8849
rect 17067 8800 17068 8840
rect 17108 8800 17109 8840
rect 17067 8791 17109 8800
rect 1699 8756 1757 8757
rect 1699 8716 1708 8756
rect 1748 8716 1757 8756
rect 1699 8715 1757 8716
rect 2083 8756 2141 8757
rect 2083 8716 2092 8756
rect 2132 8716 2141 8756
rect 2083 8715 2141 8716
rect 2467 8756 2525 8757
rect 2467 8716 2476 8756
rect 2516 8716 2525 8756
rect 2467 8715 2525 8716
rect 2851 8756 2909 8757
rect 2851 8716 2860 8756
rect 2900 8716 2909 8756
rect 2851 8715 2909 8716
rect 15627 8756 15669 8765
rect 15627 8716 15628 8756
rect 15668 8716 15669 8756
rect 15627 8707 15669 8716
rect 15723 8756 15765 8765
rect 15723 8716 15724 8756
rect 15764 8716 15765 8756
rect 15723 8707 15765 8716
rect 16683 8686 16725 8695
rect 3523 8672 3581 8673
rect 3523 8632 3532 8672
rect 3572 8632 3581 8672
rect 3523 8631 3581 8632
rect 4771 8672 4829 8673
rect 4771 8632 4780 8672
rect 4820 8632 4829 8672
rect 4771 8631 4829 8632
rect 5635 8672 5693 8673
rect 5635 8632 5644 8672
rect 5684 8632 5693 8672
rect 5635 8631 5693 8632
rect 6883 8672 6941 8673
rect 6883 8632 6892 8672
rect 6932 8632 6941 8672
rect 6883 8631 6941 8632
rect 7459 8672 7517 8673
rect 7459 8632 7468 8672
rect 7508 8632 7517 8672
rect 7459 8631 7517 8632
rect 8707 8672 8765 8673
rect 8707 8632 8716 8672
rect 8756 8632 8765 8672
rect 8707 8631 8765 8632
rect 9763 8672 9821 8673
rect 9763 8632 9772 8672
rect 9812 8632 9821 8672
rect 9763 8631 9821 8632
rect 11011 8672 11069 8673
rect 11011 8632 11020 8672
rect 11060 8632 11069 8672
rect 11011 8631 11069 8632
rect 11587 8672 11645 8673
rect 11587 8632 11596 8672
rect 11636 8632 11645 8672
rect 11587 8631 11645 8632
rect 12835 8672 12893 8673
rect 12835 8632 12844 8672
rect 12884 8632 12893 8672
rect 12835 8631 12893 8632
rect 13411 8672 13469 8673
rect 13411 8632 13420 8672
rect 13460 8632 13469 8672
rect 13411 8631 13469 8632
rect 14659 8672 14717 8673
rect 14659 8632 14668 8672
rect 14708 8632 14717 8672
rect 14659 8631 14717 8632
rect 15147 8672 15189 8681
rect 15147 8632 15148 8672
rect 15188 8632 15189 8672
rect 15147 8623 15189 8632
rect 15243 8672 15285 8681
rect 15243 8632 15244 8672
rect 15284 8632 15285 8672
rect 15243 8623 15285 8632
rect 16195 8672 16253 8673
rect 16195 8632 16204 8672
rect 16244 8632 16253 8672
rect 16683 8646 16684 8686
rect 16724 8646 16725 8686
rect 16683 8637 16725 8646
rect 17251 8672 17309 8673
rect 16195 8631 16253 8632
rect 17251 8632 17260 8672
rect 17300 8632 17309 8672
rect 17251 8631 17309 8632
rect 18499 8672 18557 8673
rect 18499 8632 18508 8672
rect 18548 8632 18557 8672
rect 18499 8631 18557 8632
rect 18691 8672 18749 8673
rect 18691 8632 18700 8672
rect 18740 8632 18749 8672
rect 18691 8631 18749 8632
rect 19939 8672 19997 8673
rect 19939 8632 19948 8672
rect 19988 8632 19997 8672
rect 19939 8631 19997 8632
rect 16875 8504 16917 8513
rect 16875 8464 16876 8504
rect 16916 8464 16917 8504
rect 16875 8455 16917 8464
rect 1152 8336 20452 8360
rect 1152 8296 4928 8336
rect 4968 8296 5010 8336
rect 5050 8296 5092 8336
rect 5132 8296 5174 8336
rect 5214 8296 5256 8336
rect 5296 8296 20048 8336
rect 20088 8296 20130 8336
rect 20170 8296 20212 8336
rect 20252 8296 20294 8336
rect 20334 8296 20376 8336
rect 20416 8296 20452 8336
rect 1152 8272 20452 8296
rect 1419 8168 1461 8177
rect 1419 8128 1420 8168
rect 1460 8128 1461 8168
rect 1419 8119 1461 8128
rect 1803 8168 1845 8177
rect 1803 8128 1804 8168
rect 1844 8128 1845 8168
rect 1803 8119 1845 8128
rect 5643 8168 5685 8177
rect 5643 8128 5644 8168
rect 5684 8128 5685 8168
rect 5643 8119 5685 8128
rect 15051 8168 15093 8177
rect 15051 8128 15052 8168
rect 15092 8128 15093 8168
rect 15051 8119 15093 8128
rect 10827 8084 10869 8093
rect 10827 8044 10828 8084
rect 10868 8044 10869 8084
rect 4195 8042 4253 8043
rect 4195 8002 4204 8042
rect 4244 8002 4253 8042
rect 10827 8035 10869 8044
rect 12843 8084 12885 8093
rect 12843 8044 12844 8084
rect 12884 8044 12885 8084
rect 12843 8035 12885 8044
rect 19947 8084 19989 8093
rect 19947 8044 19948 8084
rect 19988 8044 19989 8084
rect 19947 8035 19989 8044
rect 4195 8001 4253 8002
rect 2179 8000 2237 8001
rect 2179 7960 2188 8000
rect 2228 7960 2237 8000
rect 2179 7959 2237 7960
rect 3427 8000 3485 8001
rect 3427 7960 3436 8000
rect 3476 7960 3485 8000
rect 3427 7959 3485 7960
rect 5443 8000 5501 8001
rect 5443 7960 5452 8000
rect 5492 7960 5501 8000
rect 5443 7959 5501 7960
rect 6115 8000 6173 8001
rect 6115 7960 6124 8000
rect 6164 7960 6173 8000
rect 6115 7959 6173 7960
rect 7363 8000 7421 8001
rect 7363 7960 7372 8000
rect 7412 7960 7421 8000
rect 7363 7959 7421 7960
rect 7747 8000 7805 8001
rect 7747 7960 7756 8000
rect 7796 7960 7805 8000
rect 7747 7959 7805 7960
rect 8995 8000 9053 8001
rect 8995 7960 9004 8000
rect 9044 7960 9053 8000
rect 8995 7959 9053 7960
rect 9379 8000 9437 8001
rect 9379 7960 9388 8000
rect 9428 7960 9437 8000
rect 9379 7959 9437 7960
rect 10627 8000 10685 8001
rect 10627 7960 10636 8000
rect 10676 7960 10685 8000
rect 10627 7959 10685 7960
rect 11115 8000 11157 8009
rect 11115 7960 11116 8000
rect 11156 7960 11157 8000
rect 11115 7951 11157 7960
rect 11211 8000 11253 8009
rect 11211 7960 11212 8000
rect 11252 7960 11253 8000
rect 11211 7951 11253 7960
rect 11595 8000 11637 8009
rect 11595 7960 11596 8000
rect 11636 7960 11637 8000
rect 11595 7951 11637 7960
rect 11691 8000 11733 8009
rect 11691 7960 11692 8000
rect 11732 7960 11733 8000
rect 11691 7951 11733 7960
rect 12163 8000 12221 8001
rect 12163 7960 12172 8000
rect 12212 7960 12221 8000
rect 13603 8000 13661 8001
rect 12163 7959 12221 7960
rect 12699 7958 12741 7967
rect 13603 7960 13612 8000
rect 13652 7960 13661 8000
rect 13603 7959 13661 7960
rect 14851 8000 14909 8001
rect 14851 7960 14860 8000
rect 14900 7960 14909 8000
rect 14851 7959 14909 7960
rect 15427 8000 15485 8001
rect 15427 7960 15436 8000
rect 15476 7960 15485 8000
rect 15427 7959 15485 7960
rect 16675 8000 16733 8001
rect 16675 7960 16684 8000
rect 16724 7960 16733 8000
rect 18315 8000 18357 8009
rect 16675 7959 16733 7960
rect 18219 7981 18261 7990
rect 12699 7918 12700 7958
rect 12740 7918 12741 7958
rect 18219 7941 18220 7981
rect 18260 7941 18261 7981
rect 18315 7960 18316 8000
rect 18356 7960 18357 8000
rect 18315 7951 18357 7960
rect 18699 8000 18741 8009
rect 18699 7960 18700 8000
rect 18740 7960 18741 8000
rect 18699 7951 18741 7960
rect 19267 8000 19325 8001
rect 19267 7960 19276 8000
rect 19316 7960 19325 8000
rect 19267 7959 19325 7960
rect 19755 7986 19797 7995
rect 18219 7932 18261 7941
rect 19755 7946 19756 7986
rect 19796 7946 19797 7986
rect 19755 7937 19797 7946
rect 1603 7916 1661 7917
rect 1603 7876 1612 7916
rect 1652 7876 1661 7916
rect 1603 7875 1661 7876
rect 1987 7916 2045 7917
rect 1987 7876 1996 7916
rect 2036 7876 2045 7916
rect 12699 7909 12741 7918
rect 18795 7916 18837 7925
rect 1987 7875 2045 7876
rect 18795 7876 18796 7916
rect 18836 7876 18837 7916
rect 18795 7867 18837 7876
rect 3627 7748 3669 7757
rect 3627 7708 3628 7748
rect 3668 7708 3669 7748
rect 3627 7699 3669 7708
rect 7563 7748 7605 7757
rect 7563 7708 7564 7748
rect 7604 7708 7605 7748
rect 7563 7699 7605 7708
rect 9195 7748 9237 7757
rect 9195 7708 9196 7748
rect 9236 7708 9237 7748
rect 9195 7699 9237 7708
rect 15243 7748 15285 7757
rect 15243 7708 15244 7748
rect 15284 7708 15285 7748
rect 15243 7699 15285 7708
rect 1152 7580 20352 7604
rect 1152 7540 3688 7580
rect 3728 7540 3770 7580
rect 3810 7540 3852 7580
rect 3892 7540 3934 7580
rect 3974 7540 4016 7580
rect 4056 7540 18808 7580
rect 18848 7540 18890 7580
rect 18930 7540 18972 7580
rect 19012 7540 19054 7580
rect 19094 7540 19136 7580
rect 19176 7540 20352 7580
rect 1152 7516 20352 7540
rect 1419 7412 1461 7421
rect 1419 7372 1420 7412
rect 1460 7372 1461 7412
rect 1419 7363 1461 7372
rect 1803 7412 1845 7421
rect 1803 7372 1804 7412
rect 1844 7372 1845 7412
rect 1803 7363 1845 7372
rect 13035 7412 13077 7421
rect 13035 7372 13036 7412
rect 13076 7372 13077 7412
rect 13035 7363 13077 7372
rect 17931 7412 17973 7421
rect 17931 7372 17932 7412
rect 17972 7372 17973 7412
rect 17931 7363 17973 7372
rect 1603 7244 1661 7245
rect 1603 7204 1612 7244
rect 1652 7204 1661 7244
rect 1603 7203 1661 7204
rect 1987 7244 2045 7245
rect 1987 7204 1996 7244
rect 2036 7204 2045 7244
rect 1987 7203 2045 7204
rect 4395 7244 4437 7253
rect 4395 7204 4396 7244
rect 4436 7204 4437 7244
rect 4395 7195 4437 7204
rect 4491 7244 4533 7253
rect 4491 7204 4492 7244
rect 4532 7204 4533 7244
rect 4491 7195 4533 7204
rect 6699 7244 6741 7253
rect 6699 7204 6700 7244
rect 6740 7204 6741 7244
rect 6699 7195 6741 7204
rect 6795 7244 6837 7253
rect 6795 7204 6796 7244
rect 6836 7204 6837 7244
rect 6795 7195 6837 7204
rect 9387 7244 9429 7253
rect 9387 7204 9388 7244
rect 9428 7204 9429 7244
rect 8899 7202 8957 7203
rect 5499 7169 5541 7178
rect 8427 7174 8469 7183
rect 2371 7160 2429 7161
rect 2371 7120 2380 7160
rect 2420 7120 2429 7160
rect 2371 7119 2429 7120
rect 3619 7160 3677 7161
rect 3619 7120 3628 7160
rect 3668 7120 3677 7160
rect 3619 7119 3677 7120
rect 3915 7160 3957 7169
rect 3915 7120 3916 7160
rect 3956 7120 3957 7160
rect 3915 7111 3957 7120
rect 4011 7160 4053 7169
rect 4011 7120 4012 7160
rect 4052 7120 4053 7160
rect 4011 7111 4053 7120
rect 4963 7160 5021 7161
rect 4963 7120 4972 7160
rect 5012 7120 5021 7160
rect 5499 7129 5500 7169
rect 5540 7129 5541 7169
rect 5499 7120 5541 7129
rect 6219 7160 6261 7169
rect 6219 7120 6220 7160
rect 6260 7120 6261 7160
rect 4963 7119 5021 7120
rect 6219 7111 6261 7120
rect 6315 7160 6357 7169
rect 7755 7165 7797 7174
rect 6315 7120 6316 7160
rect 6356 7120 6357 7160
rect 6315 7111 6357 7120
rect 7267 7160 7325 7161
rect 7267 7120 7276 7160
rect 7316 7120 7325 7160
rect 7267 7119 7325 7120
rect 7755 7125 7756 7165
rect 7796 7125 7797 7165
rect 8427 7134 8428 7174
rect 8468 7134 8469 7174
rect 8899 7162 8908 7202
rect 8948 7162 8957 7202
rect 9387 7195 9429 7204
rect 15051 7244 15093 7253
rect 15051 7204 15052 7244
rect 15092 7204 15093 7244
rect 15051 7195 15093 7204
rect 16491 7244 16533 7253
rect 16491 7204 16492 7244
rect 16532 7204 16533 7244
rect 16491 7195 16533 7204
rect 16587 7244 16629 7253
rect 16587 7204 16588 7244
rect 16628 7204 16629 7244
rect 16587 7195 16629 7204
rect 19747 7244 19805 7245
rect 19747 7204 19756 7244
rect 19796 7204 19805 7244
rect 19747 7203 19805 7204
rect 14091 7174 14133 7183
rect 8899 7161 8957 7162
rect 8427 7125 8469 7134
rect 9483 7160 9525 7169
rect 7755 7116 7797 7125
rect 9483 7120 9484 7160
rect 9524 7120 9525 7160
rect 9483 7111 9525 7120
rect 9867 7160 9909 7169
rect 9867 7120 9868 7160
rect 9908 7120 9909 7160
rect 9867 7111 9909 7120
rect 9963 7160 10005 7169
rect 9963 7120 9964 7160
rect 10004 7120 10005 7160
rect 9963 7111 10005 7120
rect 11587 7160 11645 7161
rect 11587 7120 11596 7160
rect 11636 7120 11645 7160
rect 11587 7119 11645 7120
rect 12835 7160 12893 7161
rect 12835 7120 12844 7160
rect 12884 7120 12893 7160
rect 14091 7134 14092 7174
rect 14132 7134 14133 7174
rect 14091 7125 14133 7134
rect 14563 7160 14621 7161
rect 12835 7119 12893 7120
rect 14563 7120 14572 7160
rect 14612 7120 14621 7160
rect 14563 7119 14621 7120
rect 15147 7160 15189 7169
rect 15147 7120 15148 7160
rect 15188 7120 15189 7160
rect 15147 7111 15189 7120
rect 15531 7160 15573 7169
rect 15531 7120 15532 7160
rect 15572 7120 15573 7160
rect 16011 7160 16053 7169
rect 15531 7111 15573 7120
rect 15627 7140 15669 7149
rect 15627 7100 15628 7140
rect 15668 7100 15669 7140
rect 16011 7120 16012 7160
rect 16052 7120 16053 7160
rect 16011 7111 16053 7120
rect 16107 7160 16149 7169
rect 17547 7165 17589 7174
rect 16107 7120 16108 7160
rect 16148 7120 16149 7160
rect 16107 7111 16149 7120
rect 17059 7160 17117 7161
rect 17059 7120 17068 7160
rect 17108 7120 17117 7160
rect 17059 7119 17117 7120
rect 17547 7125 17548 7165
rect 17588 7125 17589 7165
rect 17547 7116 17589 7125
rect 18115 7160 18173 7161
rect 18115 7120 18124 7160
rect 18164 7120 18173 7160
rect 18115 7119 18173 7120
rect 19363 7160 19421 7161
rect 19363 7120 19372 7160
rect 19412 7120 19421 7160
rect 19363 7119 19421 7120
rect 15627 7091 15669 7100
rect 7947 7076 7989 7085
rect 7947 7036 7948 7076
rect 7988 7036 7989 7076
rect 7947 7027 7989 7036
rect 2187 6992 2229 7001
rect 2187 6952 2188 6992
rect 2228 6952 2229 6992
rect 2187 6943 2229 6952
rect 5643 6992 5685 7001
rect 5643 6952 5644 6992
rect 5684 6952 5685 6992
rect 5643 6943 5685 6952
rect 8235 6992 8277 7001
rect 8235 6952 8236 6992
rect 8276 6952 8277 6992
rect 8235 6943 8277 6952
rect 13899 6992 13941 7001
rect 13899 6952 13900 6992
rect 13940 6952 13941 6992
rect 13899 6943 13941 6952
rect 17739 6992 17781 7001
rect 17739 6952 17740 6992
rect 17780 6952 17781 6992
rect 17739 6943 17781 6952
rect 19563 6992 19605 7001
rect 19563 6952 19564 6992
rect 19604 6952 19605 6992
rect 19563 6943 19605 6952
rect 1152 6824 20452 6848
rect 1152 6784 4928 6824
rect 4968 6784 5010 6824
rect 5050 6784 5092 6824
rect 5132 6784 5174 6824
rect 5214 6784 5256 6824
rect 5296 6784 20048 6824
rect 20088 6784 20130 6824
rect 20170 6784 20212 6824
rect 20252 6784 20294 6824
rect 20334 6784 20376 6824
rect 20416 6784 20452 6824
rect 1152 6760 20452 6784
rect 1515 6656 1557 6665
rect 1515 6616 1516 6656
rect 1556 6616 1557 6656
rect 1515 6607 1557 6616
rect 1899 6656 1941 6665
rect 1899 6616 1900 6656
rect 1940 6616 1941 6656
rect 1899 6607 1941 6616
rect 6123 6656 6165 6665
rect 6123 6616 6124 6656
rect 6164 6616 6165 6656
rect 6123 6607 6165 6616
rect 7755 6656 7797 6665
rect 7755 6616 7756 6656
rect 7796 6616 7797 6656
rect 7755 6607 7797 6616
rect 8427 6656 8469 6665
rect 8427 6616 8428 6656
rect 8468 6616 8469 6656
rect 8427 6607 8469 6616
rect 14667 6656 14709 6665
rect 14667 6616 14668 6656
rect 14708 6616 14709 6656
rect 14667 6607 14709 6616
rect 17259 6656 17301 6665
rect 17259 6616 17260 6656
rect 17300 6616 17301 6656
rect 17259 6607 17301 6616
rect 19755 6656 19797 6665
rect 19755 6616 19756 6656
rect 19796 6616 19797 6656
rect 19755 6607 19797 6616
rect 2667 6572 2709 6581
rect 2667 6532 2668 6572
rect 2708 6532 2709 6572
rect 2667 6523 2709 6532
rect 13035 6572 13077 6581
rect 13035 6532 13036 6572
rect 13076 6532 13077 6572
rect 13035 6523 13077 6532
rect 2859 6483 2901 6492
rect 2859 6443 2860 6483
rect 2900 6443 2901 6483
rect 3331 6488 3389 6489
rect 3331 6448 3340 6488
rect 3380 6448 3389 6488
rect 3331 6447 3389 6448
rect 3819 6488 3861 6497
rect 3819 6448 3820 6488
rect 3860 6448 3861 6488
rect 2859 6434 2901 6443
rect 3819 6439 3861 6448
rect 3915 6488 3957 6497
rect 3915 6448 3916 6488
rect 3956 6448 3957 6488
rect 3915 6439 3957 6448
rect 4299 6488 4341 6497
rect 4299 6448 4300 6488
rect 4340 6448 4341 6488
rect 4299 6439 4341 6448
rect 4395 6488 4437 6497
rect 4395 6448 4396 6488
rect 4436 6448 4437 6488
rect 4395 6439 4437 6448
rect 4675 6488 4733 6489
rect 4675 6448 4684 6488
rect 4724 6448 4733 6488
rect 4675 6447 4733 6448
rect 5923 6488 5981 6489
rect 5923 6448 5932 6488
rect 5972 6448 5981 6488
rect 5923 6447 5981 6448
rect 7555 6488 7613 6489
rect 7555 6448 7564 6488
rect 7604 6448 7613 6488
rect 9091 6488 9149 6489
rect 7555 6447 7613 6448
rect 6307 6446 6365 6447
rect 6307 6406 6316 6446
rect 6356 6406 6365 6446
rect 6307 6405 6365 6406
rect 8571 6446 8613 6455
rect 9091 6448 9100 6488
rect 9140 6448 9149 6488
rect 9091 6447 9149 6448
rect 9675 6488 9717 6497
rect 9675 6448 9676 6488
rect 9716 6448 9717 6488
rect 8571 6406 8572 6446
rect 8612 6406 8613 6446
rect 9675 6439 9717 6448
rect 10059 6488 10101 6497
rect 10059 6448 10060 6488
rect 10100 6448 10101 6488
rect 10059 6439 10101 6448
rect 10155 6488 10197 6497
rect 10155 6448 10156 6488
rect 10196 6448 10197 6488
rect 10155 6439 10197 6448
rect 11307 6488 11349 6497
rect 11307 6448 11308 6488
rect 11348 6448 11349 6488
rect 11307 6439 11349 6448
rect 11403 6488 11445 6497
rect 11403 6448 11404 6488
rect 11444 6448 11445 6488
rect 11403 6439 11445 6448
rect 11883 6488 11925 6497
rect 11883 6448 11884 6488
rect 11924 6448 11925 6488
rect 11883 6439 11925 6448
rect 12355 6488 12413 6489
rect 12355 6448 12364 6488
rect 12404 6448 12413 6488
rect 13219 6488 13277 6489
rect 12355 6447 12413 6448
rect 12891 6446 12933 6455
rect 13219 6448 13228 6488
rect 13268 6448 13277 6488
rect 13219 6447 13277 6448
rect 14467 6488 14525 6489
rect 14467 6448 14476 6488
rect 14516 6448 14525 6488
rect 14467 6447 14525 6448
rect 15811 6488 15869 6489
rect 15811 6448 15820 6488
rect 15860 6448 15869 6488
rect 15811 6447 15869 6448
rect 17059 6488 17117 6489
rect 17059 6448 17068 6488
rect 17108 6448 17117 6488
rect 17059 6447 17117 6448
rect 18027 6488 18069 6497
rect 18027 6448 18028 6488
rect 18068 6448 18069 6488
rect 1699 6404 1757 6405
rect 1699 6364 1708 6404
rect 1748 6364 1757 6404
rect 1699 6363 1757 6364
rect 2083 6404 2141 6405
rect 2083 6364 2092 6404
rect 2132 6364 2141 6404
rect 8571 6397 8613 6406
rect 9579 6404 9621 6413
rect 2083 6363 2141 6364
rect 2467 6393 2525 6394
rect 2467 6353 2476 6393
rect 2516 6353 2525 6393
rect 9579 6364 9580 6404
rect 9620 6364 9621 6404
rect 9579 6355 9621 6364
rect 11787 6404 11829 6413
rect 11787 6364 11788 6404
rect 11828 6364 11829 6404
rect 12891 6406 12892 6446
rect 12932 6406 12933 6446
rect 18027 6439 18069 6448
rect 18123 6488 18165 6497
rect 18123 6448 18124 6488
rect 18164 6448 18165 6488
rect 18123 6439 18165 6448
rect 18507 6488 18549 6497
rect 18507 6448 18508 6488
rect 18548 6448 18549 6488
rect 18507 6439 18549 6448
rect 18603 6488 18645 6497
rect 18603 6448 18604 6488
rect 18644 6448 18645 6488
rect 18603 6439 18645 6448
rect 19075 6488 19133 6489
rect 19075 6448 19084 6488
rect 19124 6448 19133 6488
rect 19075 6447 19133 6448
rect 19563 6474 19605 6483
rect 19563 6434 19564 6474
rect 19604 6434 19605 6474
rect 19563 6425 19605 6434
rect 12891 6397 12933 6406
rect 20120 6401 20162 6410
rect 11787 6355 11829 6364
rect 20120 6361 20121 6401
rect 20161 6361 20162 6401
rect 2467 6352 2525 6353
rect 20120 6352 20162 6361
rect 19947 6320 19989 6329
rect 19947 6280 19948 6320
rect 19988 6280 19989 6320
rect 19947 6271 19989 6280
rect 2283 6236 2325 6245
rect 2283 6196 2284 6236
rect 2324 6196 2325 6236
rect 2283 6187 2325 6196
rect 1152 6068 20352 6092
rect 1152 6028 3688 6068
rect 3728 6028 3770 6068
rect 3810 6028 3852 6068
rect 3892 6028 3934 6068
rect 3974 6028 4016 6068
rect 4056 6028 18808 6068
rect 18848 6028 18890 6068
rect 18930 6028 18972 6068
rect 19012 6028 19054 6068
rect 19094 6028 19136 6068
rect 19176 6028 20352 6068
rect 1152 6004 20352 6028
rect 2667 5900 2709 5909
rect 2667 5860 2668 5900
rect 2708 5860 2709 5900
rect 2667 5851 2709 5860
rect 2859 5900 2901 5909
rect 2859 5860 2860 5900
rect 2900 5860 2901 5900
rect 2859 5851 2901 5860
rect 5931 5900 5973 5909
rect 5931 5860 5932 5900
rect 5972 5860 5973 5900
rect 5931 5851 5973 5860
rect 8139 5900 8181 5909
rect 8139 5860 8140 5900
rect 8180 5860 8181 5900
rect 8139 5851 8181 5860
rect 8331 5900 8373 5909
rect 8331 5860 8332 5900
rect 8372 5860 8373 5900
rect 8331 5851 8373 5860
rect 11403 5900 11445 5909
rect 11403 5860 11404 5900
rect 11444 5860 11445 5900
rect 11403 5851 11445 5860
rect 13131 5900 13173 5909
rect 13131 5860 13132 5900
rect 13172 5860 13173 5900
rect 13131 5851 13173 5860
rect 15435 5900 15477 5909
rect 15435 5860 15436 5900
rect 15476 5860 15477 5900
rect 15435 5851 15477 5860
rect 17739 5900 17781 5909
rect 17739 5860 17740 5900
rect 17780 5860 17781 5900
rect 17739 5851 17781 5860
rect 20131 5743 20189 5744
rect 3043 5732 3101 5733
rect 3043 5692 3052 5732
rect 3092 5692 3101 5732
rect 3043 5691 3101 5692
rect 3427 5732 3485 5733
rect 3427 5692 3436 5732
rect 3476 5692 3485 5732
rect 3427 5691 3485 5692
rect 18507 5732 18549 5741
rect 18507 5692 18508 5732
rect 18548 5692 18549 5732
rect 20131 5703 20140 5743
rect 20180 5703 20189 5743
rect 20131 5702 20189 5703
rect 18507 5683 18549 5692
rect 1219 5648 1277 5649
rect 1219 5608 1228 5648
rect 1268 5608 1277 5648
rect 1219 5607 1277 5608
rect 2467 5648 2525 5649
rect 2467 5608 2476 5648
rect 2516 5608 2525 5648
rect 2467 5607 2525 5608
rect 4483 5648 4541 5649
rect 4483 5608 4492 5648
rect 4532 5608 4541 5648
rect 4483 5607 4541 5608
rect 5731 5648 5789 5649
rect 5731 5608 5740 5648
rect 5780 5608 5789 5648
rect 5731 5607 5789 5608
rect 6691 5648 6749 5649
rect 6691 5608 6700 5648
rect 6740 5608 6749 5648
rect 6691 5607 6749 5608
rect 7939 5648 7997 5649
rect 7939 5608 7948 5648
rect 7988 5608 7997 5648
rect 7939 5607 7997 5608
rect 8515 5648 8573 5649
rect 8515 5608 8524 5648
rect 8564 5608 8573 5648
rect 8515 5607 8573 5608
rect 9763 5648 9821 5649
rect 9763 5608 9772 5648
rect 9812 5608 9821 5648
rect 9763 5607 9821 5608
rect 9955 5648 10013 5649
rect 9955 5608 9964 5648
rect 10004 5608 10013 5648
rect 9955 5607 10013 5608
rect 11203 5648 11261 5649
rect 11203 5608 11212 5648
rect 11252 5608 11261 5648
rect 11203 5607 11261 5608
rect 11683 5648 11741 5649
rect 11683 5608 11692 5648
rect 11732 5608 11741 5648
rect 11683 5607 11741 5608
rect 12931 5648 12989 5649
rect 12931 5608 12940 5648
rect 12980 5608 12989 5648
rect 12931 5607 12989 5608
rect 13987 5648 14045 5649
rect 13987 5608 13996 5648
rect 14036 5608 14045 5648
rect 13987 5607 14045 5608
rect 15235 5648 15293 5649
rect 15235 5608 15244 5648
rect 15284 5608 15293 5648
rect 15235 5607 15293 5608
rect 16291 5648 16349 5649
rect 16291 5608 16300 5648
rect 16340 5608 16349 5648
rect 16291 5607 16349 5608
rect 17539 5648 17597 5649
rect 17539 5608 17548 5648
rect 17588 5608 17597 5648
rect 17539 5607 17597 5608
rect 18027 5648 18069 5657
rect 18027 5608 18028 5648
rect 18068 5608 18069 5648
rect 18027 5599 18069 5608
rect 18123 5648 18165 5657
rect 18123 5608 18124 5648
rect 18164 5608 18165 5648
rect 18123 5599 18165 5608
rect 18603 5648 18645 5657
rect 19563 5653 19605 5662
rect 18603 5608 18604 5648
rect 18644 5608 18645 5648
rect 18603 5599 18645 5608
rect 19075 5648 19133 5649
rect 19075 5608 19084 5648
rect 19124 5608 19133 5648
rect 19075 5607 19133 5608
rect 19563 5613 19564 5653
rect 19604 5613 19605 5653
rect 19563 5604 19605 5613
rect 19755 5564 19797 5573
rect 19755 5524 19756 5564
rect 19796 5524 19797 5564
rect 19755 5515 19797 5524
rect 3243 5480 3285 5489
rect 3243 5440 3244 5480
rect 3284 5440 3285 5480
rect 3243 5431 3285 5440
rect 19947 5480 19989 5489
rect 19947 5440 19948 5480
rect 19988 5440 19989 5480
rect 19947 5431 19989 5440
rect 1152 5312 20452 5336
rect 1152 5272 4928 5312
rect 4968 5272 5010 5312
rect 5050 5272 5092 5312
rect 5132 5272 5174 5312
rect 5214 5272 5256 5312
rect 5296 5272 20048 5312
rect 20088 5272 20130 5312
rect 20170 5272 20212 5312
rect 20252 5272 20294 5312
rect 20334 5272 20376 5312
rect 20416 5272 20452 5312
rect 1152 5248 20452 5272
rect 7755 5144 7797 5153
rect 7755 5104 7756 5144
rect 7796 5104 7797 5144
rect 7755 5095 7797 5104
rect 18315 5144 18357 5153
rect 18315 5104 18316 5144
rect 18356 5104 18357 5144
rect 18315 5095 18357 5104
rect 3531 5060 3573 5069
rect 3531 5020 3532 5060
rect 3572 5020 3573 5060
rect 3531 5011 3573 5020
rect 5643 5060 5685 5069
rect 5643 5020 5644 5060
rect 5684 5020 5685 5060
rect 5643 5011 5685 5020
rect 13035 5060 13077 5069
rect 13035 5020 13036 5060
rect 13076 5020 13077 5060
rect 13035 5011 13077 5020
rect 15051 5060 15093 5069
rect 15051 5020 15052 5060
rect 15092 5020 15093 5060
rect 15051 5011 15093 5020
rect 20043 5060 20085 5069
rect 20043 5020 20044 5060
rect 20084 5020 20085 5060
rect 20043 5011 20085 5020
rect 2083 4976 2141 4977
rect 2083 4936 2092 4976
rect 2132 4936 2141 4976
rect 2083 4935 2141 4936
rect 3331 4976 3389 4977
rect 3331 4936 3340 4976
rect 3380 4936 3389 4976
rect 3331 4935 3389 4936
rect 3915 4976 3957 4985
rect 3915 4936 3916 4976
rect 3956 4936 3957 4976
rect 3915 4927 3957 4936
rect 4011 4976 4053 4985
rect 4011 4936 4012 4976
rect 4052 4936 4053 4976
rect 4011 4927 4053 4936
rect 4395 4976 4437 4985
rect 4395 4936 4396 4976
rect 4436 4936 4437 4976
rect 4395 4927 4437 4936
rect 4491 4976 4533 4985
rect 4491 4936 4492 4976
rect 4532 4936 4533 4976
rect 4491 4927 4533 4936
rect 4963 4976 5021 4977
rect 4963 4936 4972 4976
rect 5012 4936 5021 4976
rect 6027 4976 6069 4985
rect 4963 4935 5021 4936
rect 5451 4962 5493 4971
rect 5451 4922 5452 4962
rect 5492 4922 5493 4962
rect 6027 4936 6028 4976
rect 6068 4936 6069 4976
rect 6027 4927 6069 4936
rect 6123 4976 6165 4985
rect 6123 4936 6124 4976
rect 6164 4936 6165 4976
rect 6123 4927 6165 4936
rect 6507 4976 6549 4985
rect 6507 4936 6508 4976
rect 6548 4936 6549 4976
rect 6507 4927 6549 4936
rect 6603 4976 6645 4985
rect 6603 4936 6604 4976
rect 6644 4936 6645 4976
rect 6603 4927 6645 4936
rect 7075 4976 7133 4977
rect 7075 4936 7084 4976
rect 7124 4936 7133 4976
rect 8323 4976 8381 4977
rect 7075 4935 7133 4936
rect 7563 4962 7605 4971
rect 5451 4913 5493 4922
rect 7563 4922 7564 4962
rect 7604 4922 7605 4962
rect 8323 4936 8332 4976
rect 8372 4936 8381 4976
rect 8323 4935 8381 4936
rect 9571 4976 9629 4977
rect 9571 4936 9580 4976
rect 9620 4936 9629 4976
rect 9571 4935 9629 4936
rect 9955 4976 10013 4977
rect 9955 4936 9964 4976
rect 10004 4936 10013 4976
rect 9955 4935 10013 4936
rect 11203 4976 11261 4977
rect 11203 4936 11212 4976
rect 11252 4936 11261 4976
rect 11203 4935 11261 4936
rect 11587 4976 11645 4977
rect 11587 4936 11596 4976
rect 11636 4936 11645 4976
rect 11587 4935 11645 4936
rect 12835 4976 12893 4977
rect 12835 4936 12844 4976
rect 12884 4936 12893 4976
rect 13419 4976 13461 4985
rect 12835 4935 12893 4936
rect 13323 4957 13365 4966
rect 7563 4913 7605 4922
rect 13323 4917 13324 4957
rect 13364 4917 13365 4957
rect 13419 4936 13420 4976
rect 13460 4936 13461 4976
rect 13419 4927 13461 4936
rect 13803 4976 13845 4985
rect 13803 4936 13804 4976
rect 13844 4936 13845 4976
rect 13803 4927 13845 4936
rect 14371 4976 14429 4977
rect 14371 4936 14380 4976
rect 14420 4936 14429 4976
rect 15235 4976 15293 4977
rect 14371 4935 14429 4936
rect 14859 4962 14901 4971
rect 13323 4908 13365 4917
rect 14859 4922 14860 4962
rect 14900 4922 14901 4962
rect 15235 4936 15244 4976
rect 15284 4936 15293 4976
rect 15235 4935 15293 4936
rect 16483 4976 16541 4977
rect 16483 4936 16492 4976
rect 16532 4936 16541 4976
rect 16483 4935 16541 4936
rect 16867 4976 16925 4977
rect 16867 4936 16876 4976
rect 16916 4936 16925 4976
rect 16867 4935 16925 4936
rect 18115 4976 18173 4977
rect 18115 4936 18124 4976
rect 18164 4936 18173 4976
rect 18115 4935 18173 4936
rect 18595 4976 18653 4977
rect 18595 4936 18604 4976
rect 18644 4936 18653 4976
rect 18595 4935 18653 4936
rect 19843 4976 19901 4977
rect 19843 4936 19852 4976
rect 19892 4936 19901 4976
rect 19843 4935 19901 4936
rect 14859 4913 14901 4922
rect 1507 4892 1565 4893
rect 1507 4852 1516 4892
rect 1556 4852 1565 4892
rect 1507 4851 1565 4852
rect 1891 4892 1949 4893
rect 1891 4852 1900 4892
rect 1940 4852 1949 4892
rect 1891 4851 1949 4852
rect 13899 4892 13941 4901
rect 13899 4852 13900 4892
rect 13940 4852 13941 4892
rect 13899 4843 13941 4852
rect 1323 4808 1365 4817
rect 1323 4768 1324 4808
rect 1364 4768 1365 4808
rect 1323 4759 1365 4768
rect 1707 4808 1749 4817
rect 1707 4768 1708 4808
rect 1748 4768 1749 4808
rect 1707 4759 1749 4768
rect 9771 4724 9813 4733
rect 9771 4684 9772 4724
rect 9812 4684 9813 4724
rect 9771 4675 9813 4684
rect 11403 4724 11445 4733
rect 11403 4684 11404 4724
rect 11444 4684 11445 4724
rect 11403 4675 11445 4684
rect 16683 4724 16725 4733
rect 16683 4684 16684 4724
rect 16724 4684 16725 4724
rect 16683 4675 16725 4684
rect 1152 4556 20352 4580
rect 1152 4516 3688 4556
rect 3728 4516 3770 4556
rect 3810 4516 3852 4556
rect 3892 4516 3934 4556
rect 3974 4516 4016 4556
rect 4056 4516 18808 4556
rect 18848 4516 18890 4556
rect 18930 4516 18972 4556
rect 19012 4516 19054 4556
rect 19094 4516 19136 4556
rect 19176 4516 20352 4556
rect 1152 4492 20352 4516
rect 7083 4388 7125 4397
rect 7083 4348 7084 4388
rect 7124 4348 7125 4388
rect 7083 4339 7125 4348
rect 14667 4388 14709 4397
rect 14667 4348 14668 4388
rect 14708 4348 14709 4388
rect 14667 4339 14709 4348
rect 17355 4388 17397 4397
rect 17355 4348 17356 4388
rect 17396 4348 17397 4388
rect 17355 4339 17397 4348
rect 17739 4388 17781 4397
rect 17739 4348 17740 4388
rect 17780 4348 17781 4388
rect 17739 4339 17781 4348
rect 4011 4220 4053 4229
rect 4011 4180 4012 4220
rect 4052 4180 4053 4220
rect 4011 4171 4053 4180
rect 4107 4220 4149 4229
rect 4107 4180 4108 4220
rect 4148 4180 4149 4220
rect 4107 4171 4149 4180
rect 5059 4220 5117 4221
rect 5059 4180 5068 4220
rect 5108 4180 5117 4220
rect 5059 4179 5117 4180
rect 7851 4220 7893 4229
rect 7851 4180 7852 4220
rect 7892 4180 7893 4220
rect 7851 4171 7893 4180
rect 7947 4220 7989 4229
rect 7947 4180 7948 4220
rect 7988 4180 7989 4220
rect 7947 4171 7989 4180
rect 10635 4220 10677 4229
rect 10635 4180 10636 4220
rect 10676 4180 10677 4220
rect 10635 4171 10677 4180
rect 10731 4220 10773 4229
rect 10731 4180 10732 4220
rect 10772 4180 10773 4220
rect 10731 4171 10773 4180
rect 15531 4220 15573 4229
rect 15531 4180 15532 4220
rect 15572 4180 15573 4220
rect 15531 4171 15573 4180
rect 17539 4220 17597 4221
rect 17539 4180 17548 4220
rect 17588 4180 17597 4220
rect 17539 4179 17597 4180
rect 17923 4220 17981 4221
rect 17923 4180 17932 4220
rect 17972 4180 17981 4220
rect 17923 4179 17981 4180
rect 18699 4220 18741 4229
rect 18699 4180 18700 4220
rect 18740 4180 18741 4220
rect 18699 4171 18741 4180
rect 18795 4220 18837 4229
rect 18795 4180 18796 4220
rect 18836 4180 18837 4220
rect 18795 4171 18837 4180
rect 3003 4145 3045 4154
rect 8955 4145 8997 4154
rect 11691 4150 11733 4159
rect 1219 4136 1277 4137
rect 1219 4096 1228 4136
rect 1268 4096 1277 4136
rect 1219 4095 1277 4096
rect 2467 4136 2525 4137
rect 2467 4096 2476 4136
rect 2516 4096 2525 4136
rect 3003 4105 3004 4145
rect 3044 4105 3045 4145
rect 3003 4096 3045 4105
rect 3523 4136 3581 4137
rect 3523 4096 3532 4136
rect 3572 4096 3581 4136
rect 2467 4095 2525 4096
rect 3523 4095 3581 4096
rect 4491 4136 4533 4145
rect 4491 4096 4492 4136
rect 4532 4096 4533 4136
rect 4491 4087 4533 4096
rect 4587 4136 4629 4145
rect 4587 4096 4588 4136
rect 4628 4096 4629 4136
rect 4587 4087 4629 4096
rect 5635 4136 5693 4137
rect 5635 4096 5644 4136
rect 5684 4096 5693 4136
rect 5635 4095 5693 4096
rect 6883 4136 6941 4137
rect 6883 4096 6892 4136
rect 6932 4096 6941 4136
rect 6883 4095 6941 4096
rect 7371 4136 7413 4145
rect 7371 4096 7372 4136
rect 7412 4096 7413 4136
rect 7371 4087 7413 4096
rect 7467 4136 7509 4145
rect 7467 4096 7468 4136
rect 7508 4096 7509 4136
rect 7467 4087 7509 4096
rect 8419 4136 8477 4137
rect 8419 4096 8428 4136
rect 8468 4096 8477 4136
rect 8955 4105 8956 4145
rect 8996 4105 8997 4145
rect 8955 4096 8997 4105
rect 10155 4136 10197 4145
rect 10155 4096 10156 4136
rect 10196 4096 10197 4136
rect 8419 4095 8477 4096
rect 10155 4087 10197 4096
rect 10251 4136 10293 4145
rect 10251 4096 10252 4136
rect 10292 4096 10293 4136
rect 10251 4087 10293 4096
rect 11203 4136 11261 4137
rect 11203 4096 11212 4136
rect 11252 4096 11261 4136
rect 11691 4110 11692 4150
rect 11732 4110 11733 4150
rect 16491 4150 16533 4159
rect 11691 4101 11733 4110
rect 13219 4136 13277 4137
rect 11203 4095 11261 4096
rect 13219 4096 13228 4136
rect 13268 4096 13277 4136
rect 13219 4095 13277 4096
rect 14467 4136 14525 4137
rect 14467 4096 14476 4136
rect 14516 4096 14525 4136
rect 14467 4095 14525 4096
rect 14955 4136 14997 4145
rect 14955 4096 14956 4136
rect 14996 4096 14997 4136
rect 14955 4087 14997 4096
rect 15051 4136 15093 4145
rect 15051 4096 15052 4136
rect 15092 4096 15093 4136
rect 15051 4087 15093 4096
rect 15435 4136 15477 4145
rect 15435 4096 15436 4136
rect 15476 4096 15477 4136
rect 15435 4087 15477 4096
rect 16003 4136 16061 4137
rect 16003 4096 16012 4136
rect 16052 4096 16061 4136
rect 16491 4110 16492 4150
rect 16532 4110 16533 4150
rect 16491 4101 16533 4110
rect 18219 4136 18261 4145
rect 16003 4095 16061 4096
rect 18219 4096 18220 4136
rect 18260 4096 18261 4136
rect 18219 4087 18261 4096
rect 18315 4136 18357 4145
rect 19755 4141 19797 4150
rect 18315 4096 18316 4136
rect 18356 4096 18357 4136
rect 18315 4087 18357 4096
rect 19267 4136 19325 4137
rect 19267 4096 19276 4136
rect 19316 4096 19325 4136
rect 19267 4095 19325 4096
rect 19755 4101 19756 4141
rect 19796 4101 19797 4141
rect 19755 4092 19797 4101
rect 2667 4052 2709 4061
rect 2667 4012 2668 4052
rect 2708 4012 2709 4052
rect 2667 4003 2709 4012
rect 11883 4052 11925 4061
rect 11883 4012 11884 4052
rect 11924 4012 11925 4052
rect 11883 4003 11925 4012
rect 19947 4052 19989 4061
rect 19947 4012 19948 4052
rect 19988 4012 19989 4052
rect 19947 4003 19989 4012
rect 2859 3968 2901 3977
rect 2859 3928 2860 3968
rect 2900 3928 2901 3968
rect 2859 3919 2901 3928
rect 4875 3968 4917 3977
rect 4875 3928 4876 3968
rect 4916 3928 4917 3968
rect 4875 3919 4917 3928
rect 9099 3968 9141 3977
rect 9099 3928 9100 3968
rect 9140 3928 9141 3968
rect 9099 3919 9141 3928
rect 16683 3968 16725 3977
rect 16683 3928 16684 3968
rect 16724 3928 16725 3968
rect 16683 3919 16725 3928
rect 1152 3800 20452 3824
rect 1152 3760 4928 3800
rect 4968 3760 5010 3800
rect 5050 3760 5092 3800
rect 5132 3760 5174 3800
rect 5214 3760 5256 3800
rect 5296 3760 20048 3800
rect 20088 3760 20130 3800
rect 20170 3760 20212 3800
rect 20252 3760 20294 3800
rect 20334 3760 20376 3800
rect 20416 3760 20452 3800
rect 1152 3736 20452 3760
rect 1899 3632 1941 3641
rect 1899 3592 1900 3632
rect 1940 3592 1941 3632
rect 1899 3583 1941 3592
rect 2667 3632 2709 3641
rect 2667 3592 2668 3632
rect 2708 3592 2709 3632
rect 2667 3583 2709 3592
rect 5739 3632 5781 3641
rect 5739 3592 5740 3632
rect 5780 3592 5781 3632
rect 5739 3583 5781 3592
rect 7467 3632 7509 3641
rect 7467 3592 7468 3632
rect 7508 3592 7509 3632
rect 7467 3583 7509 3592
rect 9195 3632 9237 3641
rect 9195 3592 9196 3632
rect 9236 3592 9237 3632
rect 9195 3583 9237 3592
rect 14955 3632 14997 3641
rect 14955 3592 14956 3632
rect 14996 3592 14997 3632
rect 14955 3583 14997 3592
rect 20043 3632 20085 3641
rect 20043 3592 20044 3632
rect 20084 3592 20085 3632
rect 20043 3583 20085 3592
rect 11019 3548 11061 3557
rect 11019 3508 11020 3548
rect 11060 3508 11061 3548
rect 11019 3499 11061 3508
rect 13035 3548 13077 3557
rect 13035 3508 13036 3548
rect 13076 3508 13077 3548
rect 13035 3499 13077 3508
rect 18411 3548 18453 3557
rect 18411 3508 18412 3548
rect 18452 3508 18453 3548
rect 18411 3499 18453 3508
rect 2851 3464 2909 3465
rect 2851 3424 2860 3464
rect 2900 3424 2909 3464
rect 2851 3423 2909 3424
rect 4099 3464 4157 3465
rect 4099 3424 4108 3464
rect 4148 3424 4157 3464
rect 4099 3423 4157 3424
rect 4291 3464 4349 3465
rect 4291 3424 4300 3464
rect 4340 3424 4349 3464
rect 4291 3423 4349 3424
rect 5539 3464 5597 3465
rect 5539 3424 5548 3464
rect 5588 3424 5597 3464
rect 5539 3423 5597 3424
rect 6019 3464 6077 3465
rect 6019 3424 6028 3464
rect 6068 3424 6077 3464
rect 6019 3423 6077 3424
rect 7267 3464 7325 3465
rect 7267 3424 7276 3464
rect 7316 3424 7325 3464
rect 7267 3423 7325 3424
rect 7747 3464 7805 3465
rect 7747 3424 7756 3464
rect 7796 3424 7805 3464
rect 7747 3423 7805 3424
rect 8995 3464 9053 3465
rect 8995 3424 9004 3464
rect 9044 3424 9053 3464
rect 8995 3423 9053 3424
rect 9571 3464 9629 3465
rect 9571 3424 9580 3464
rect 9620 3424 9629 3464
rect 9571 3423 9629 3424
rect 10819 3464 10877 3465
rect 10819 3424 10828 3464
rect 10868 3424 10877 3464
rect 10819 3423 10877 3424
rect 11307 3464 11349 3473
rect 11307 3424 11308 3464
rect 11348 3424 11349 3464
rect 11307 3415 11349 3424
rect 11403 3464 11445 3473
rect 11403 3424 11404 3464
rect 11444 3424 11445 3464
rect 11403 3415 11445 3424
rect 11787 3464 11829 3473
rect 11787 3424 11788 3464
rect 11828 3424 11829 3464
rect 11787 3415 11829 3424
rect 11883 3464 11925 3473
rect 11883 3424 11884 3464
rect 11924 3424 11925 3464
rect 11883 3415 11925 3424
rect 12355 3464 12413 3465
rect 12355 3424 12364 3464
rect 12404 3424 12413 3464
rect 13507 3464 13565 3465
rect 12355 3423 12413 3424
rect 12891 3454 12933 3463
rect 12891 3414 12892 3454
rect 12932 3414 12933 3454
rect 13507 3424 13516 3464
rect 13556 3424 13565 3464
rect 13507 3423 13565 3424
rect 14755 3464 14813 3465
rect 14755 3424 14764 3464
rect 14804 3424 14813 3464
rect 14755 3423 14813 3424
rect 16683 3464 16725 3473
rect 16683 3424 16684 3464
rect 16724 3424 16725 3464
rect 16683 3415 16725 3424
rect 16779 3464 16821 3473
rect 16779 3424 16780 3464
rect 16820 3424 16821 3464
rect 16779 3415 16821 3424
rect 17163 3464 17205 3473
rect 17163 3424 17164 3464
rect 17204 3424 17205 3464
rect 17163 3415 17205 3424
rect 17259 3464 17301 3473
rect 17259 3424 17260 3464
rect 17300 3424 17301 3464
rect 17259 3415 17301 3424
rect 17731 3464 17789 3465
rect 17731 3424 17740 3464
rect 17780 3424 17789 3464
rect 18595 3464 18653 3465
rect 17731 3423 17789 3424
rect 18267 3422 18309 3431
rect 18595 3424 18604 3464
rect 18644 3424 18653 3464
rect 18595 3423 18653 3424
rect 19843 3464 19901 3465
rect 19843 3424 19852 3464
rect 19892 3424 19901 3464
rect 19843 3423 19901 3424
rect 12891 3405 12933 3414
rect 18267 3382 18268 3422
rect 18308 3382 18309 3422
rect 1699 3380 1757 3381
rect 1699 3340 1708 3380
rect 1748 3340 1757 3380
rect 1699 3339 1757 3340
rect 2083 3380 2141 3381
rect 2083 3340 2092 3380
rect 2132 3340 2141 3380
rect 2083 3339 2141 3340
rect 2467 3380 2525 3381
rect 2467 3340 2476 3380
rect 2516 3340 2525 3380
rect 2467 3339 2525 3340
rect 15427 3380 15485 3381
rect 15427 3340 15436 3380
rect 15476 3340 15485 3380
rect 18267 3373 18309 3382
rect 15427 3339 15485 3340
rect 2283 3296 2325 3305
rect 2283 3256 2284 3296
rect 2324 3256 2325 3296
rect 2283 3247 2325 3256
rect 1515 3212 1557 3221
rect 1515 3172 1516 3212
rect 1556 3172 1557 3212
rect 1515 3163 1557 3172
rect 15243 3212 15285 3221
rect 15243 3172 15244 3212
rect 15284 3172 15285 3212
rect 15243 3163 15285 3172
rect 1152 3044 20352 3068
rect 1152 3004 3688 3044
rect 3728 3004 3770 3044
rect 3810 3004 3852 3044
rect 3892 3004 3934 3044
rect 3974 3004 4016 3044
rect 4056 3004 18808 3044
rect 18848 3004 18890 3044
rect 18930 3004 18972 3044
rect 19012 3004 19054 3044
rect 19094 3004 19136 3044
rect 19176 3004 20352 3044
rect 1152 2980 20352 3004
rect 2283 2876 2325 2885
rect 2283 2836 2284 2876
rect 2324 2836 2325 2876
rect 2283 2827 2325 2836
rect 7659 2876 7701 2885
rect 7659 2836 7660 2876
rect 7700 2836 7701 2876
rect 7659 2827 7701 2836
rect 8043 2876 8085 2885
rect 8043 2836 8044 2876
rect 8084 2836 8085 2876
rect 8043 2827 8085 2836
rect 13323 2876 13365 2885
rect 13323 2836 13324 2876
rect 13364 2836 13365 2876
rect 13323 2827 13365 2836
rect 16779 2876 16821 2885
rect 16779 2836 16780 2876
rect 16820 2836 16821 2876
rect 16779 2827 16821 2836
rect 18411 2876 18453 2885
rect 18411 2836 18412 2876
rect 18452 2836 18453 2876
rect 18411 2827 18453 2836
rect 20043 2876 20085 2885
rect 20043 2836 20044 2876
rect 20084 2836 20085 2876
rect 20043 2827 20085 2836
rect 1899 2792 1941 2801
rect 1899 2752 1900 2792
rect 1940 2752 1941 2792
rect 1899 2743 1941 2752
rect 8419 2719 8477 2720
rect 1699 2708 1757 2709
rect 1699 2668 1708 2708
rect 1748 2668 1757 2708
rect 1699 2667 1757 2668
rect 2083 2708 2141 2709
rect 2083 2668 2092 2708
rect 2132 2668 2141 2708
rect 2083 2667 2141 2668
rect 2467 2708 2525 2709
rect 2467 2668 2476 2708
rect 2516 2668 2525 2708
rect 2467 2667 2525 2668
rect 5155 2708 5213 2709
rect 5155 2668 5164 2708
rect 5204 2668 5213 2708
rect 5155 2667 5213 2668
rect 5931 2708 5973 2717
rect 5931 2668 5932 2708
rect 5972 2668 5973 2708
rect 5931 2659 5973 2668
rect 6027 2708 6069 2717
rect 6027 2668 6028 2708
rect 6068 2668 6069 2708
rect 6027 2659 6069 2668
rect 7843 2708 7901 2709
rect 7843 2668 7852 2708
rect 7892 2668 7901 2708
rect 7843 2667 7901 2668
rect 8227 2708 8285 2709
rect 8227 2668 8236 2708
rect 8276 2668 8285 2708
rect 8419 2679 8428 2719
rect 8468 2679 8477 2719
rect 8419 2678 8477 2679
rect 9379 2708 9437 2709
rect 8227 2667 8285 2668
rect 9379 2668 9388 2708
rect 9428 2668 9437 2708
rect 9379 2667 9437 2668
rect 9763 2708 9821 2709
rect 9763 2668 9772 2708
rect 9812 2668 9821 2708
rect 9763 2667 9821 2668
rect 10147 2708 10205 2709
rect 10147 2668 10156 2708
rect 10196 2668 10205 2708
rect 10147 2667 10205 2668
rect 11107 2708 11165 2709
rect 11107 2668 11116 2708
rect 11156 2668 11165 2708
rect 11107 2667 11165 2668
rect 13699 2708 13757 2709
rect 13699 2668 13708 2708
rect 13748 2668 13757 2708
rect 13699 2667 13757 2668
rect 14083 2708 14141 2709
rect 14083 2668 14092 2708
rect 14132 2668 14141 2708
rect 14083 2667 14141 2668
rect 14467 2708 14525 2709
rect 14467 2668 14476 2708
rect 14516 2668 14525 2708
rect 14467 2667 14525 2668
rect 14851 2708 14909 2709
rect 14851 2668 14860 2708
rect 14900 2668 14909 2708
rect 14851 2667 14909 2668
rect 16579 2645 16637 2646
rect 3051 2624 3093 2633
rect 3051 2584 3052 2624
rect 3092 2584 3093 2624
rect 3051 2575 3093 2584
rect 3147 2624 3189 2633
rect 3147 2584 3148 2624
rect 3188 2584 3189 2624
rect 3147 2575 3189 2584
rect 3531 2624 3573 2633
rect 3531 2584 3532 2624
rect 3572 2584 3573 2624
rect 3531 2575 3573 2584
rect 3627 2624 3669 2633
rect 4587 2629 4629 2638
rect 3627 2584 3628 2624
rect 3668 2584 3669 2624
rect 3627 2575 3669 2584
rect 4099 2624 4157 2625
rect 4099 2584 4108 2624
rect 4148 2584 4157 2624
rect 4099 2583 4157 2584
rect 4587 2589 4588 2629
rect 4628 2589 4629 2629
rect 4587 2580 4629 2589
rect 5451 2624 5493 2633
rect 5451 2584 5452 2624
rect 5492 2584 5493 2624
rect 5451 2575 5493 2584
rect 5547 2624 5589 2633
rect 6987 2629 7029 2638
rect 5547 2584 5548 2624
rect 5588 2584 5589 2624
rect 5547 2575 5589 2584
rect 6499 2624 6557 2625
rect 6499 2584 6508 2624
rect 6548 2584 6557 2624
rect 6499 2583 6557 2584
rect 6987 2589 6988 2629
rect 7028 2589 7029 2629
rect 6987 2580 7029 2589
rect 11875 2624 11933 2625
rect 11875 2584 11884 2624
rect 11924 2584 11933 2624
rect 11875 2583 11933 2584
rect 13123 2624 13181 2625
rect 13123 2584 13132 2624
rect 13172 2584 13181 2624
rect 13123 2583 13181 2584
rect 15331 2624 15389 2625
rect 15331 2584 15340 2624
rect 15380 2584 15389 2624
rect 16579 2605 16588 2645
rect 16628 2605 16637 2645
rect 16579 2604 16637 2605
rect 16963 2624 17021 2625
rect 15331 2583 15389 2584
rect 16963 2584 16972 2624
rect 17012 2584 17021 2624
rect 16963 2583 17021 2584
rect 18211 2624 18269 2625
rect 18211 2584 18220 2624
rect 18260 2584 18269 2624
rect 18211 2583 18269 2584
rect 18595 2624 18653 2625
rect 18595 2584 18604 2624
rect 18644 2584 18653 2624
rect 18595 2583 18653 2584
rect 19843 2624 19901 2625
rect 19843 2584 19852 2624
rect 19892 2584 19901 2624
rect 19843 2583 19901 2584
rect 4779 2540 4821 2549
rect 4779 2500 4780 2540
rect 4820 2500 4821 2540
rect 4779 2491 4821 2500
rect 7179 2540 7221 2549
rect 7179 2500 7180 2540
rect 7220 2500 7221 2540
rect 7179 2491 7221 2500
rect 1515 2456 1557 2465
rect 1515 2416 1516 2456
rect 1556 2416 1557 2456
rect 1515 2407 1557 2416
rect 4971 2456 5013 2465
rect 4971 2416 4972 2456
rect 5012 2416 5013 2456
rect 4971 2407 5013 2416
rect 8619 2456 8661 2465
rect 8619 2416 8620 2456
rect 8660 2416 8661 2456
rect 8619 2407 8661 2416
rect 9579 2456 9621 2465
rect 9579 2416 9580 2456
rect 9620 2416 9621 2456
rect 9579 2407 9621 2416
rect 9963 2456 10005 2465
rect 9963 2416 9964 2456
rect 10004 2416 10005 2456
rect 9963 2407 10005 2416
rect 10347 2456 10389 2465
rect 10347 2416 10348 2456
rect 10388 2416 10389 2456
rect 10347 2407 10389 2416
rect 10923 2456 10965 2465
rect 10923 2416 10924 2456
rect 10964 2416 10965 2456
rect 10923 2407 10965 2416
rect 13515 2456 13557 2465
rect 13515 2416 13516 2456
rect 13556 2416 13557 2456
rect 13515 2407 13557 2416
rect 13899 2456 13941 2465
rect 13899 2416 13900 2456
rect 13940 2416 13941 2456
rect 13899 2407 13941 2416
rect 14283 2456 14325 2465
rect 14283 2416 14284 2456
rect 14324 2416 14325 2456
rect 14283 2407 14325 2416
rect 14667 2456 14709 2465
rect 14667 2416 14668 2456
rect 14708 2416 14709 2456
rect 14667 2407 14709 2416
rect 1152 2288 20452 2312
rect 1152 2248 4928 2288
rect 4968 2248 5010 2288
rect 5050 2248 5092 2288
rect 5132 2248 5174 2288
rect 5214 2248 5256 2288
rect 5296 2248 20048 2288
rect 20088 2248 20130 2288
rect 20170 2248 20212 2288
rect 20252 2248 20294 2288
rect 20334 2248 20376 2288
rect 20416 2248 20452 2288
rect 1152 2224 20452 2248
rect 2859 2120 2901 2129
rect 2859 2080 2860 2120
rect 2900 2080 2901 2120
rect 2859 2071 2901 2080
rect 4491 2120 4533 2129
rect 4491 2080 4492 2120
rect 4532 2080 4533 2120
rect 4491 2071 4533 2080
rect 6123 2120 6165 2129
rect 6123 2080 6124 2120
rect 6164 2080 6165 2120
rect 6123 2071 6165 2080
rect 9867 2120 9909 2129
rect 9867 2080 9868 2120
rect 9908 2080 9909 2120
rect 9867 2071 9909 2080
rect 18219 2120 18261 2129
rect 18219 2080 18220 2120
rect 18260 2080 18261 2120
rect 18219 2071 18261 2080
rect 19947 2120 19989 2129
rect 19947 2080 19948 2120
rect 19988 2080 19989 2120
rect 19947 2071 19989 2080
rect 7851 2036 7893 2045
rect 7851 1996 7852 2036
rect 7892 1996 7893 2036
rect 3043 1994 3101 1995
rect 3043 1954 3052 1994
rect 3092 1954 3101 1994
rect 7851 1987 7893 1996
rect 16587 2036 16629 2045
rect 16587 1996 16588 2036
rect 16628 1996 16629 2036
rect 16587 1987 16629 1996
rect 3043 1953 3101 1954
rect 1411 1952 1469 1953
rect 1411 1912 1420 1952
rect 1460 1912 1469 1952
rect 1411 1911 1469 1912
rect 2659 1952 2717 1953
rect 2659 1912 2668 1952
rect 2708 1912 2717 1952
rect 2659 1911 2717 1912
rect 4291 1952 4349 1953
rect 4291 1912 4300 1952
rect 4340 1912 4349 1952
rect 4291 1911 4349 1912
rect 4675 1952 4733 1953
rect 4675 1912 4684 1952
rect 4724 1912 4733 1952
rect 4675 1911 4733 1912
rect 5923 1952 5981 1953
rect 5923 1912 5932 1952
rect 5972 1912 5981 1952
rect 5923 1911 5981 1912
rect 6403 1952 6461 1953
rect 6403 1912 6412 1952
rect 6452 1912 6461 1952
rect 6403 1911 6461 1912
rect 7651 1952 7709 1953
rect 7651 1912 7660 1952
rect 7700 1912 7709 1952
rect 7651 1911 7709 1912
rect 8139 1952 8181 1961
rect 8139 1912 8140 1952
rect 8180 1912 8181 1952
rect 8139 1903 8181 1912
rect 8235 1952 8277 1961
rect 8235 1912 8236 1952
rect 8276 1912 8277 1952
rect 8235 1903 8277 1912
rect 8715 1952 8757 1961
rect 8715 1912 8716 1952
rect 8756 1912 8757 1952
rect 8715 1903 8757 1912
rect 9187 1952 9245 1953
rect 9187 1912 9196 1952
rect 9236 1912 9245 1952
rect 12451 1952 12509 1953
rect 9187 1911 9245 1912
rect 9675 1938 9717 1947
rect 9675 1898 9676 1938
rect 9716 1898 9717 1938
rect 12451 1912 12460 1952
rect 12500 1912 12509 1952
rect 12451 1911 12509 1912
rect 13699 1952 13757 1953
rect 13699 1912 13708 1952
rect 13748 1912 13757 1952
rect 13699 1911 13757 1912
rect 14859 1952 14901 1961
rect 14859 1912 14860 1952
rect 14900 1912 14901 1952
rect 14859 1903 14901 1912
rect 14955 1952 14997 1961
rect 14955 1912 14956 1952
rect 14996 1912 14997 1952
rect 14955 1903 14997 1912
rect 15339 1952 15381 1961
rect 15339 1912 15340 1952
rect 15380 1912 15381 1952
rect 15339 1903 15381 1912
rect 15435 1952 15477 1961
rect 15435 1912 15436 1952
rect 15476 1912 15477 1952
rect 15435 1903 15477 1912
rect 15907 1952 15965 1953
rect 15907 1912 15916 1952
rect 15956 1912 15965 1952
rect 16771 1952 16829 1953
rect 15907 1911 15965 1912
rect 16395 1938 16437 1947
rect 9675 1889 9717 1898
rect 16395 1898 16396 1938
rect 16436 1898 16437 1938
rect 16771 1912 16780 1952
rect 16820 1912 16829 1952
rect 16771 1911 16829 1912
rect 18019 1952 18077 1953
rect 18019 1912 18028 1952
rect 18068 1912 18077 1952
rect 18019 1911 18077 1912
rect 18499 1952 18557 1953
rect 18499 1912 18508 1952
rect 18548 1912 18557 1952
rect 18499 1911 18557 1912
rect 19747 1952 19805 1953
rect 19747 1912 19756 1952
rect 19796 1912 19805 1952
rect 19747 1911 19805 1912
rect 16395 1889 16437 1898
rect 8619 1868 8661 1877
rect 8619 1828 8620 1868
rect 8660 1828 8661 1868
rect 8619 1819 8661 1828
rect 10051 1868 10109 1869
rect 10051 1828 10060 1868
rect 10100 1828 10109 1868
rect 10051 1827 10109 1828
rect 10435 1868 10493 1869
rect 10435 1828 10444 1868
rect 10484 1828 10493 1868
rect 10435 1827 10493 1828
rect 11011 1868 11069 1869
rect 11011 1828 11020 1868
rect 11060 1828 11069 1868
rect 11011 1827 11069 1828
rect 11203 1868 11261 1869
rect 11203 1828 11212 1868
rect 11252 1828 11261 1868
rect 11203 1827 11261 1828
rect 11587 1868 11645 1869
rect 11587 1828 11596 1868
rect 11636 1828 11645 1868
rect 11587 1827 11645 1828
rect 12259 1868 12317 1869
rect 12259 1828 12268 1868
rect 12308 1828 12317 1868
rect 12259 1827 12317 1828
rect 14091 1868 14133 1877
rect 14091 1828 14092 1868
rect 14132 1828 14133 1868
rect 14091 1819 14133 1828
rect 14371 1868 14429 1869
rect 14371 1828 14380 1868
rect 14420 1828 14429 1868
rect 14371 1827 14429 1828
rect 13899 1784 13941 1793
rect 13899 1744 13900 1784
rect 13940 1744 13941 1784
rect 13899 1735 13941 1744
rect 10251 1700 10293 1709
rect 10251 1660 10252 1700
rect 10292 1660 10293 1700
rect 10251 1651 10293 1660
rect 10635 1700 10677 1709
rect 10635 1660 10636 1700
rect 10676 1660 10677 1700
rect 10635 1651 10677 1660
rect 10827 1700 10869 1709
rect 10827 1660 10828 1700
rect 10868 1660 10869 1700
rect 10827 1651 10869 1660
rect 11403 1700 11445 1709
rect 11403 1660 11404 1700
rect 11444 1660 11445 1700
rect 11403 1651 11445 1660
rect 11787 1700 11829 1709
rect 11787 1660 11788 1700
rect 11828 1660 11829 1700
rect 11787 1651 11829 1660
rect 12075 1700 12117 1709
rect 12075 1660 12076 1700
rect 12116 1660 12117 1700
rect 12075 1651 12117 1660
rect 14571 1700 14613 1709
rect 14571 1660 14572 1700
rect 14612 1660 14613 1700
rect 14571 1651 14613 1660
rect 1152 1532 20352 1556
rect 1152 1492 3688 1532
rect 3728 1492 3770 1532
rect 3810 1492 3852 1532
rect 3892 1492 3934 1532
rect 3974 1492 4016 1532
rect 4056 1492 18808 1532
rect 18848 1492 18890 1532
rect 18930 1492 18972 1532
rect 19012 1492 19054 1532
rect 19094 1492 19136 1532
rect 19176 1492 20352 1532
rect 1152 1468 20352 1492
rect 9675 1364 9717 1373
rect 9675 1324 9676 1364
rect 9716 1324 9717 1364
rect 9675 1315 9717 1324
rect 16875 1364 16917 1373
rect 16875 1324 16876 1364
rect 16916 1324 16917 1364
rect 16875 1315 16917 1324
rect 1515 1280 1557 1289
rect 1515 1240 1516 1280
rect 1556 1240 1557 1280
rect 1515 1231 1557 1240
rect 1899 1280 1941 1289
rect 1899 1240 1900 1280
rect 1940 1240 1941 1280
rect 1899 1231 1941 1240
rect 2283 1280 2325 1289
rect 2283 1240 2284 1280
rect 2324 1240 2325 1280
rect 2283 1231 2325 1240
rect 4683 1280 4725 1289
rect 4683 1240 4684 1280
rect 4724 1240 4725 1280
rect 4683 1231 4725 1240
rect 6795 1280 6837 1289
rect 6795 1240 6796 1280
rect 6836 1240 6837 1280
rect 6795 1231 6837 1240
rect 7851 1280 7893 1289
rect 7851 1240 7852 1280
rect 7892 1240 7893 1280
rect 7851 1231 7893 1240
rect 1699 1196 1757 1197
rect 1699 1156 1708 1196
rect 1748 1156 1757 1196
rect 1699 1155 1757 1156
rect 2083 1196 2141 1197
rect 2083 1156 2092 1196
rect 2132 1156 2141 1196
rect 2083 1155 2141 1156
rect 2467 1196 2525 1197
rect 2467 1156 2476 1196
rect 2516 1156 2525 1196
rect 2467 1155 2525 1156
rect 2851 1196 2909 1197
rect 2851 1156 2860 1196
rect 2900 1156 2909 1196
rect 2851 1155 2909 1156
rect 4867 1196 4925 1197
rect 4867 1156 4876 1196
rect 4916 1156 4925 1196
rect 4867 1155 4925 1156
rect 7459 1196 7517 1197
rect 7459 1156 7468 1196
rect 7508 1156 7517 1196
rect 7459 1155 7517 1156
rect 8035 1196 8093 1197
rect 8035 1156 8044 1196
rect 8084 1156 8093 1196
rect 8035 1155 8093 1156
rect 10051 1196 10109 1197
rect 10051 1156 10060 1196
rect 10100 1156 10109 1196
rect 10051 1155 10109 1156
rect 10435 1196 10493 1197
rect 10435 1156 10444 1196
rect 10484 1156 10493 1196
rect 10435 1155 10493 1156
rect 10819 1196 10877 1197
rect 10819 1156 10828 1196
rect 10868 1156 10877 1196
rect 10819 1155 10877 1156
rect 11203 1196 11261 1197
rect 11203 1156 11212 1196
rect 11252 1156 11261 1196
rect 11203 1155 11261 1156
rect 12643 1196 12701 1197
rect 12643 1156 12652 1196
rect 12692 1156 12701 1196
rect 12643 1155 12701 1156
rect 13027 1196 13085 1197
rect 13027 1156 13036 1196
rect 13076 1156 13085 1196
rect 13027 1155 13085 1156
rect 13411 1196 13469 1197
rect 13411 1156 13420 1196
rect 13460 1156 13469 1196
rect 13411 1155 13469 1156
rect 13795 1196 13853 1197
rect 13795 1156 13804 1196
rect 13844 1156 13853 1196
rect 13795 1155 13853 1156
rect 14275 1196 14333 1197
rect 14275 1156 14284 1196
rect 14324 1156 14333 1196
rect 14275 1155 14333 1156
rect 14659 1196 14717 1197
rect 14659 1156 14668 1196
rect 14708 1156 14717 1196
rect 14659 1155 14717 1156
rect 15043 1196 15101 1197
rect 15043 1156 15052 1196
rect 15092 1156 15101 1196
rect 15043 1155 15101 1156
rect 17347 1196 17405 1197
rect 17347 1156 17356 1196
rect 17396 1156 17405 1196
rect 17347 1155 17405 1156
rect 18403 1196 18461 1197
rect 18403 1156 18412 1196
rect 18452 1156 18461 1196
rect 18403 1155 18461 1156
rect 3235 1112 3293 1113
rect 3235 1072 3244 1112
rect 3284 1072 3293 1112
rect 3235 1071 3293 1072
rect 4483 1112 4541 1113
rect 4483 1072 4492 1112
rect 4532 1072 4541 1112
rect 4483 1071 4541 1072
rect 5347 1112 5405 1113
rect 5347 1072 5356 1112
rect 5396 1072 5405 1112
rect 5347 1071 5405 1072
rect 6595 1112 6653 1113
rect 6595 1072 6604 1112
rect 6644 1072 6653 1112
rect 6595 1071 6653 1072
rect 8227 1112 8285 1113
rect 8227 1072 8236 1112
rect 8276 1072 8285 1112
rect 8227 1071 8285 1072
rect 9475 1112 9533 1113
rect 9475 1072 9484 1112
rect 9524 1072 9533 1112
rect 9475 1071 9533 1072
rect 15427 1112 15485 1113
rect 15427 1072 15436 1112
rect 15476 1072 15485 1112
rect 15427 1071 15485 1072
rect 16675 1112 16733 1113
rect 16675 1072 16684 1112
rect 16724 1072 16733 1112
rect 16675 1071 16733 1072
rect 2667 944 2709 953
rect 2667 904 2668 944
rect 2708 904 2709 944
rect 2667 895 2709 904
rect 5067 944 5109 953
rect 5067 904 5068 944
rect 5108 904 5109 944
rect 5067 895 5109 904
rect 7659 944 7701 953
rect 7659 904 7660 944
rect 7700 904 7701 944
rect 7659 895 7701 904
rect 10251 944 10293 953
rect 10251 904 10252 944
rect 10292 904 10293 944
rect 10251 895 10293 904
rect 10635 944 10677 953
rect 10635 904 10636 944
rect 10676 904 10677 944
rect 10635 895 10677 904
rect 11019 944 11061 953
rect 11019 904 11020 944
rect 11060 904 11061 944
rect 11019 895 11061 904
rect 11403 944 11445 953
rect 11403 904 11404 944
rect 11444 904 11445 944
rect 11403 895 11445 904
rect 12459 944 12501 953
rect 12459 904 12460 944
rect 12500 904 12501 944
rect 12459 895 12501 904
rect 12843 944 12885 953
rect 12843 904 12844 944
rect 12884 904 12885 944
rect 12843 895 12885 904
rect 13227 944 13269 953
rect 13227 904 13228 944
rect 13268 904 13269 944
rect 13227 895 13269 904
rect 13611 944 13653 953
rect 13611 904 13612 944
rect 13652 904 13653 944
rect 13611 895 13653 904
rect 14091 944 14133 953
rect 14091 904 14092 944
rect 14132 904 14133 944
rect 14091 895 14133 904
rect 14475 944 14517 953
rect 14475 904 14476 944
rect 14516 904 14517 944
rect 14475 895 14517 904
rect 14859 944 14901 953
rect 14859 904 14860 944
rect 14900 904 14901 944
rect 14859 895 14901 904
rect 17163 944 17205 953
rect 17163 904 17164 944
rect 17204 904 17205 944
rect 17163 895 17205 904
rect 18219 944 18261 953
rect 18219 904 18220 944
rect 18260 904 18261 944
rect 18219 895 18261 904
rect 1152 776 20452 800
rect 1152 736 4928 776
rect 4968 736 5010 776
rect 5050 736 5092 776
rect 5132 736 5174 776
rect 5214 736 5256 776
rect 5296 736 20048 776
rect 20088 736 20130 776
rect 20170 736 20212 776
rect 20252 736 20294 776
rect 20334 736 20376 776
rect 20416 736 20452 776
rect 1152 712 20452 736
<< via1 >>
rect 4928 41560 4968 41600
rect 5010 41560 5050 41600
rect 5092 41560 5132 41600
rect 5174 41560 5214 41600
rect 5256 41560 5296 41600
rect 20048 41560 20088 41600
rect 20130 41560 20170 41600
rect 20212 41560 20252 41600
rect 20294 41560 20334 41600
rect 20376 41560 20416 41600
rect 2092 41392 2132 41432
rect 5740 41392 5780 41432
rect 6124 41392 6164 41432
rect 9964 41392 10004 41432
rect 10348 41392 10388 41432
rect 13804 41392 13844 41432
rect 15724 41392 15764 41432
rect 16108 41392 16148 41432
rect 17260 41392 17300 41432
rect 17836 41392 17876 41432
rect 18124 41392 18164 41432
rect 18700 41392 18740 41432
rect 19756 41392 19796 41432
rect 2284 41224 2324 41264
rect 3532 41224 3572 41264
rect 4108 41224 4148 41264
rect 5356 41224 5396 41264
rect 6508 41224 6548 41264
rect 7756 41224 7796 41264
rect 8140 41224 8180 41264
rect 9388 41224 9428 41264
rect 11980 41224 12020 41264
rect 13228 41224 13268 41264
rect 1708 41140 1748 41180
rect 1900 41140 1940 41180
rect 5548 41140 5588 41180
rect 5932 41140 5972 41180
rect 9772 41140 9812 41180
rect 10156 41140 10196 41180
rect 10540 41140 10580 41180
rect 11596 41140 11636 41180
rect 13996 41140 14036 41180
rect 14572 41140 14612 41180
rect 14956 41140 14996 41180
rect 15340 41140 15380 41180
rect 15916 41140 15956 41180
rect 16300 41140 16340 41180
rect 16588 41140 16628 41180
rect 16972 41140 17012 41180
rect 17452 41140 17492 41180
rect 17644 41140 17684 41180
rect 18316 41140 18356 41180
rect 18508 41140 18548 41180
rect 19084 41140 19124 41180
rect 19372 41140 19412 41180
rect 19948 41140 19988 41180
rect 1324 41056 1364 41096
rect 3724 41056 3764 41096
rect 9580 41056 9620 41096
rect 11788 41056 11828 41096
rect 16780 41056 16820 41096
rect 18892 41056 18932 41096
rect 3916 40972 3956 41012
rect 6316 40972 6356 41012
rect 7948 40972 7988 41012
rect 13420 40972 13460 41012
rect 14380 40972 14420 41012
rect 14764 40972 14804 41012
rect 15148 40972 15188 41012
rect 19564 40972 19604 41012
rect 3688 40804 3728 40844
rect 3770 40804 3810 40844
rect 3852 40804 3892 40844
rect 3934 40804 3974 40844
rect 4016 40804 4056 40844
rect 18808 40804 18848 40844
rect 18890 40804 18930 40844
rect 18972 40804 19012 40844
rect 19054 40804 19094 40844
rect 19136 40804 19176 40844
rect 1708 40636 1748 40676
rect 3052 40636 3092 40676
rect 3436 40636 3476 40676
rect 5452 40636 5492 40676
rect 5836 40636 5876 40676
rect 7948 40636 7988 40676
rect 16204 40636 16244 40676
rect 16588 40636 16628 40676
rect 16972 40636 17012 40676
rect 18124 40636 18164 40676
rect 18508 40636 18548 40676
rect 18892 40636 18932 40676
rect 11980 40552 12020 40592
rect 15820 40552 15860 40592
rect 17932 40552 17972 40592
rect 19564 40552 19604 40592
rect 1516 40468 1556 40508
rect 2284 40468 2324 40508
rect 2860 40479 2900 40519
rect 3244 40468 3284 40508
rect 5260 40468 5300 40508
rect 5644 40468 5684 40508
rect 8140 40468 8180 40508
rect 9004 40468 9044 40508
rect 16012 40468 16052 40508
rect 16396 40468 16436 40508
rect 16780 40468 16820 40508
rect 17164 40468 17204 40508
rect 17740 40468 17780 40508
rect 18316 40468 18356 40508
rect 18700 40468 18740 40508
rect 19084 40468 19124 40508
rect 19372 40468 19412 40508
rect 19852 40468 19892 40508
rect 3820 40384 3860 40424
rect 5068 40384 5108 40424
rect 6028 40384 6068 40424
rect 7276 40384 7316 40424
rect 8428 40384 8468 40424
rect 8524 40384 8564 40424
rect 8908 40384 8948 40424
rect 9484 40384 9524 40424
rect 9964 40389 10004 40429
rect 10348 40384 10388 40424
rect 11596 40405 11636 40445
rect 11980 40384 12020 40424
rect 12076 40384 12116 40424
rect 12268 40384 12308 40424
rect 12556 40384 12596 40424
rect 13804 40384 13844 40424
rect 14380 40384 14420 40424
rect 15628 40384 15668 40424
rect 1900 40300 1940 40340
rect 7468 40300 7508 40340
rect 7660 40300 7700 40340
rect 11788 40300 11828 40340
rect 17548 40300 17588 40340
rect 1228 40216 1268 40256
rect 3628 40216 3668 40256
rect 10156 40216 10196 40256
rect 13996 40216 14036 40256
rect 14188 40216 14228 40256
rect 20044 40216 20084 40256
rect 4928 40048 4968 40088
rect 5010 40048 5050 40088
rect 5092 40048 5132 40088
rect 5174 40048 5214 40088
rect 5256 40048 5296 40088
rect 20048 40048 20088 40088
rect 20130 40048 20170 40088
rect 20212 40048 20252 40088
rect 20294 40048 20334 40088
rect 20376 40048 20416 40088
rect 1708 39880 1748 39920
rect 8236 39880 8276 39920
rect 9964 39880 10004 39920
rect 12076 39880 12116 39920
rect 12940 39880 12980 39920
rect 18316 39880 18356 39920
rect 18508 39880 18548 39920
rect 18892 39880 18932 39920
rect 3724 39796 3764 39836
rect 8044 39796 8084 39836
rect 11692 39796 11732 39836
rect 15052 39796 15092 39836
rect 1996 39712 2036 39752
rect 2092 39693 2132 39733
rect 3052 39712 3092 39752
rect 3580 39702 3620 39742
rect 4012 39712 4052 39752
rect 5260 39712 5300 39752
rect 6316 39712 6356 39752
rect 6412 39712 6452 39752
rect 7372 39712 7412 39752
rect 7852 39707 7892 39747
rect 8524 39712 8564 39752
rect 9772 39712 9812 39752
rect 10252 39712 10292 39752
rect 11500 39712 11540 39752
rect 11884 39712 11924 39752
rect 11980 39712 12020 39752
rect 12172 39712 12212 39752
rect 12268 39712 12308 39752
rect 12369 39712 12409 39752
rect 12652 39712 12692 39752
rect 12748 39712 12788 39752
rect 13324 39712 13364 39752
rect 13420 39712 13460 39752
rect 14380 39712 14420 39752
rect 14860 39707 14900 39747
rect 15436 39712 15476 39752
rect 16684 39712 16724 39752
rect 16972 39712 17012 39752
rect 17164 39712 17204 39752
rect 17260 39712 17300 39752
rect 17548 39712 17588 39752
rect 17644 39712 17684 39752
rect 17740 39712 17780 39752
rect 1516 39628 1556 39668
rect 2476 39628 2516 39668
rect 2572 39628 2612 39668
rect 5932 39628 5972 39668
rect 6796 39628 6836 39668
rect 6892 39628 6932 39668
rect 13804 39628 13844 39668
rect 13900 39628 13940 39668
rect 18700 39628 18740 39668
rect 19084 39628 19124 39668
rect 19468 39628 19508 39668
rect 20044 39628 20084 39668
rect 1324 39544 1364 39584
rect 5644 39544 5684 39584
rect 18220 39544 18260 39584
rect 5452 39460 5492 39500
rect 15244 39460 15284 39500
rect 16972 39460 17012 39500
rect 17932 39460 17972 39500
rect 19660 39460 19700 39500
rect 20236 39460 20276 39500
rect 3688 39292 3728 39332
rect 3770 39292 3810 39332
rect 3852 39292 3892 39332
rect 3934 39292 3974 39332
rect 4016 39292 4056 39332
rect 18808 39292 18848 39332
rect 18890 39292 18930 39332
rect 18972 39292 19012 39332
rect 19054 39292 19094 39332
rect 19136 39292 19176 39332
rect 12460 39124 12500 39164
rect 1516 39040 1556 39080
rect 5356 39040 5396 39080
rect 5836 39040 5876 39080
rect 6220 39040 6260 39080
rect 6604 39040 6644 39080
rect 6796 39040 6836 39080
rect 8620 39040 8660 39080
rect 12844 39040 12884 39080
rect 16300 39040 16340 39080
rect 18604 39040 18644 39080
rect 1324 38956 1364 38996
rect 4972 38956 5012 38996
rect 5548 38956 5588 38996
rect 6028 38956 6068 38996
rect 6412 38956 6452 38996
rect 6988 38956 7028 38996
rect 11116 38956 11156 38996
rect 13036 38956 13076 38996
rect 14572 38956 14612 38996
rect 14668 38956 14708 38996
rect 19276 38956 19316 38996
rect 19660 38956 19700 38996
rect 20044 38956 20084 38996
rect 1708 38872 1748 38912
rect 2956 38872 2996 38912
rect 3340 38872 3380 38912
rect 4588 38872 4628 38912
rect 7180 38872 7220 38912
rect 8428 38872 8468 38912
rect 8812 38872 8852 38912
rect 10060 38872 10100 38912
rect 10540 38872 10580 38912
rect 10636 38872 10676 38912
rect 11020 38872 11060 38912
rect 11596 38872 11636 38912
rect 12076 38877 12116 38917
rect 12556 38872 12596 38912
rect 14092 38872 14132 38912
rect 14188 38872 14228 38912
rect 15148 38872 15188 38912
rect 15628 38886 15668 38926
rect 16012 38872 16052 38912
rect 16300 38872 16340 38912
rect 16492 38872 16532 38912
rect 17740 38872 17780 38912
rect 18796 38872 18836 38912
rect 18892 38872 18932 38912
rect 18988 38872 19028 38912
rect 10252 38788 10292 38828
rect 3148 38704 3188 38744
rect 4780 38704 4820 38744
rect 5164 38704 5204 38744
rect 12268 38704 12308 38744
rect 15820 38704 15860 38744
rect 17932 38704 17972 38744
rect 18124 38704 18164 38744
rect 18508 38704 18548 38744
rect 19084 38704 19124 38744
rect 19468 38704 19508 38744
rect 19852 38704 19892 38744
rect 20236 38704 20276 38744
rect 4928 38536 4968 38576
rect 5010 38536 5050 38576
rect 5092 38536 5132 38576
rect 5174 38536 5214 38576
rect 5256 38536 5296 38576
rect 20048 38536 20088 38576
rect 20130 38536 20170 38576
rect 20212 38536 20252 38576
rect 20294 38536 20334 38576
rect 20376 38536 20416 38576
rect 3148 38368 3188 38408
rect 3532 38368 3572 38408
rect 4012 38368 4052 38408
rect 8044 38368 8084 38408
rect 12076 38368 12116 38408
rect 16300 38368 16340 38408
rect 18316 38284 18356 38324
rect 18988 38284 19028 38324
rect 1228 38200 1268 38240
rect 2476 38200 2516 38240
rect 4396 38200 4436 38240
rect 5644 38200 5684 38240
rect 6412 38200 6452 38240
rect 7660 38200 7700 38240
rect 8620 38200 8660 38240
rect 9868 38200 9908 38240
rect 10636 38200 10676 38240
rect 11884 38200 11924 38240
rect 12844 38200 12884 38240
rect 14092 38200 14132 38240
rect 14476 38200 14516 38240
rect 15724 38200 15764 38240
rect 16588 38200 16628 38240
rect 16684 38200 16724 38240
rect 17644 38200 17684 38240
rect 18124 38195 18164 38235
rect 18604 38200 18644 38240
rect 18892 38200 18932 38240
rect 19756 38200 19796 38240
rect 19852 38200 19892 38240
rect 20140 38200 20180 38240
rect 2956 38116 2996 38156
rect 3340 38116 3380 38156
rect 3820 38116 3860 38156
rect 16108 38116 16148 38156
rect 17068 38116 17108 38156
rect 17164 38116 17204 38156
rect 6028 38032 6068 38072
rect 8332 38032 8372 38072
rect 19468 38032 19508 38072
rect 2668 37948 2708 37988
rect 4204 37948 4244 37988
rect 7852 37948 7892 37988
rect 10060 37948 10100 37988
rect 14284 37948 14324 37988
rect 15916 37948 15956 37988
rect 19276 37948 19316 37988
rect 3688 37780 3728 37820
rect 3770 37780 3810 37820
rect 3852 37780 3892 37820
rect 3934 37780 3974 37820
rect 4016 37780 4056 37820
rect 18808 37780 18848 37820
rect 18890 37780 18930 37820
rect 18972 37780 19012 37820
rect 19054 37780 19094 37820
rect 19136 37780 19176 37820
rect 1612 37612 1652 37652
rect 1996 37612 2036 37652
rect 6988 37612 7028 37652
rect 17644 37612 17684 37652
rect 18316 37612 18356 37652
rect 19180 37612 19220 37652
rect 4396 37528 4436 37568
rect 1420 37444 1460 37484
rect 1804 37444 1844 37484
rect 7180 37444 7220 37484
rect 9004 37444 9044 37484
rect 18124 37444 18164 37484
rect 20044 37444 20084 37484
rect 2284 37360 2324 37400
rect 2380 37360 2420 37400
rect 2764 37360 2804 37400
rect 2860 37360 2900 37400
rect 3340 37360 3380 37400
rect 3820 37374 3860 37414
rect 5068 37360 5108 37400
rect 5164 37360 5204 37400
rect 5548 37360 5588 37400
rect 5644 37360 5684 37400
rect 6124 37360 6164 37400
rect 6604 37374 6644 37414
rect 7372 37360 7412 37400
rect 7660 37360 7700 37400
rect 7948 37360 7988 37400
rect 8428 37360 8468 37400
rect 8524 37360 8564 37400
rect 8908 37360 8948 37400
rect 9484 37360 9524 37400
rect 9964 37374 10004 37414
rect 11500 37360 11540 37400
rect 12748 37360 12788 37400
rect 14092 37360 14132 37400
rect 14188 37360 14228 37400
rect 14572 37360 14612 37400
rect 15676 37402 15716 37442
rect 14668 37360 14708 37400
rect 15148 37360 15188 37400
rect 16204 37360 16244 37400
rect 17452 37360 17492 37400
rect 18988 37360 19028 37400
rect 4012 37276 4052 37316
rect 6796 37276 6836 37316
rect 4684 37192 4724 37232
rect 7468 37192 7508 37232
rect 7852 37192 7892 37232
rect 8140 37192 8180 37232
rect 10156 37192 10196 37232
rect 12940 37192 12980 37232
rect 15820 37192 15860 37232
rect 18508 37192 18548 37232
rect 20236 37192 20276 37232
rect 4928 37024 4968 37064
rect 5010 37024 5050 37064
rect 5092 37024 5132 37064
rect 5174 37024 5214 37064
rect 5256 37024 5296 37064
rect 20048 37024 20088 37064
rect 20130 37024 20170 37064
rect 20212 37024 20252 37064
rect 20294 37024 20334 37064
rect 20376 37024 20416 37064
rect 8332 36856 8372 36896
rect 16588 36856 16628 36896
rect 18124 36856 18164 36896
rect 18412 36856 18452 36896
rect 6124 36772 6164 36812
rect 8140 36772 8180 36812
rect 12940 36772 12980 36812
rect 1228 36688 1268 36728
rect 2476 36688 2516 36728
rect 4300 36688 4340 36728
rect 4684 36688 4724 36728
rect 5932 36688 5972 36728
rect 6412 36688 6452 36728
rect 3052 36646 3092 36686
rect 6508 36688 6548 36728
rect 7468 36688 7508 36728
rect 6892 36604 6932 36644
rect 6988 36604 7028 36644
rect 7996 36646 8036 36686
rect 8620 36688 8660 36728
rect 8908 36688 8948 36728
rect 9484 36688 9524 36728
rect 10732 36688 10772 36728
rect 11212 36688 11252 36728
rect 11308 36688 11348 36728
rect 12268 36688 12308 36728
rect 12796 36678 12836 36718
rect 15148 36688 15188 36728
rect 16396 36688 16436 36728
rect 17356 36688 17396 36728
rect 17452 36688 17492 36728
rect 17644 36688 17684 36728
rect 18604 36688 18644 36728
rect 19852 36688 19892 36728
rect 11692 36604 11732 36644
rect 11788 36604 11828 36644
rect 16972 36604 17012 36644
rect 20044 36604 20084 36644
rect 8428 36520 8468 36560
rect 17164 36520 17204 36560
rect 17644 36520 17684 36560
rect 18220 36520 18260 36560
rect 2668 36436 2708 36476
rect 4492 36436 4532 36476
rect 8908 36436 8948 36476
rect 10924 36436 10964 36476
rect 20236 36436 20276 36476
rect 3688 36268 3728 36308
rect 3770 36268 3810 36308
rect 3852 36268 3892 36308
rect 3934 36268 3974 36308
rect 4016 36268 4056 36308
rect 18808 36268 18848 36308
rect 18890 36268 18930 36308
rect 18972 36268 19012 36308
rect 19054 36268 19094 36308
rect 19136 36268 19176 36308
rect 1612 36100 1652 36140
rect 8236 36100 8276 36140
rect 11020 36100 11060 36140
rect 17452 36100 17492 36140
rect 17836 36100 17876 36140
rect 19468 36100 19508 36140
rect 8428 36016 8468 36056
rect 9196 36016 9236 36056
rect 1420 35932 1460 35972
rect 4972 35932 5012 35972
rect 9100 35932 9140 35972
rect 9292 35932 9332 35972
rect 17260 35932 17300 35972
rect 17644 35932 17684 35972
rect 1900 35848 1940 35888
rect 1996 35848 2036 35888
rect 2380 35848 2420 35888
rect 2476 35848 2516 35888
rect 2956 35848 2996 35888
rect 3436 35862 3476 35902
rect 4396 35848 4436 35888
rect 4492 35848 4532 35888
rect 4876 35848 4916 35888
rect 5452 35848 5492 35888
rect 5932 35853 5972 35893
rect 6412 35848 6452 35888
rect 6508 35848 6548 35888
rect 6604 35848 6644 35888
rect 6796 35848 6836 35888
rect 8044 35848 8084 35888
rect 9004 35848 9044 35888
rect 9388 35848 9428 35888
rect 9580 35848 9620 35888
rect 10828 35869 10868 35909
rect 11308 35848 11348 35888
rect 11404 35848 11444 35888
rect 11788 35848 11828 35888
rect 11884 35890 11924 35930
rect 12364 35848 12404 35888
rect 12892 35857 12932 35897
rect 15340 35848 15380 35888
rect 15436 35848 15476 35888
rect 15820 35848 15860 35888
rect 15916 35848 15956 35888
rect 16396 35848 16436 35888
rect 16924 35857 16964 35897
rect 18028 35848 18068 35888
rect 19276 35848 19316 35888
rect 19756 35848 19796 35888
rect 19852 35848 19892 35888
rect 19948 35848 19988 35888
rect 17068 35764 17108 35804
rect 3628 35680 3668 35720
rect 4012 35680 4052 35720
rect 6124 35680 6164 35720
rect 6316 35680 6356 35720
rect 8524 35680 8564 35720
rect 13036 35680 13076 35720
rect 19468 35680 19508 35720
rect 20140 35680 20180 35720
rect 4928 35512 4968 35552
rect 5010 35512 5050 35552
rect 5092 35512 5132 35552
rect 5174 35512 5214 35552
rect 5256 35512 5296 35552
rect 20048 35512 20088 35552
rect 20130 35512 20170 35552
rect 20212 35512 20252 35552
rect 20294 35512 20334 35552
rect 20376 35512 20416 35552
rect 5836 35344 5876 35384
rect 7468 35344 7508 35384
rect 10156 35348 10196 35388
rect 13324 35344 13364 35384
rect 15148 35344 15188 35384
rect 8044 35260 8084 35300
rect 10828 35260 10868 35300
rect 17164 35260 17204 35300
rect 19756 35260 19796 35300
rect 2092 35176 2132 35216
rect 3340 35176 3380 35216
rect 4396 35176 4436 35216
rect 5644 35176 5684 35216
rect 6028 35176 6068 35216
rect 7276 35176 7316 35216
rect 7948 35176 7988 35216
rect 8140 35176 8180 35216
rect 8236 35176 8276 35216
rect 8812 35176 8852 35216
rect 8716 35134 8756 35174
rect 9100 35176 9140 35216
rect 9479 35176 9519 35216
rect 9580 35176 9620 35216
rect 9676 35176 9716 35216
rect 9868 35176 9908 35216
rect 9964 35176 10004 35216
rect 10252 35176 10292 35216
rect 10348 35176 10388 35216
rect 11020 35176 11060 35216
rect 10924 35134 10964 35174
rect 11116 35176 11156 35216
rect 11308 35176 11348 35216
rect 11500 35176 11540 35216
rect 11884 35176 11924 35216
rect 13132 35176 13172 35216
rect 13708 35176 13748 35216
rect 14956 35176 14996 35216
rect 15436 35176 15476 35216
rect 15532 35176 15572 35216
rect 16492 35176 16532 35216
rect 16972 35162 17012 35202
rect 18028 35176 18068 35216
rect 18124 35176 18164 35216
rect 18508 35176 18548 35216
rect 19084 35176 19124 35216
rect 19564 35171 19604 35211
rect 19948 35176 19988 35216
rect 20044 35176 20084 35216
rect 20140 35197 20180 35237
rect 20236 35176 20276 35216
rect 1516 35092 1556 35132
rect 4012 35092 4052 35132
rect 11404 35092 11444 35132
rect 15916 35092 15956 35132
rect 16012 35092 16052 35132
rect 18604 35092 18644 35132
rect 1708 35008 1748 35048
rect 3820 35008 3860 35048
rect 8428 35008 8468 35048
rect 17644 35008 17684 35048
rect 1900 34924 1940 34964
rect 9964 34924 10004 34964
rect 10636 34882 10676 34922
rect 3688 34756 3728 34796
rect 3770 34756 3810 34796
rect 3852 34756 3892 34796
rect 3934 34756 3974 34796
rect 4016 34756 4056 34796
rect 18808 34756 18848 34796
rect 18890 34756 18930 34796
rect 18972 34756 19012 34796
rect 19054 34756 19094 34796
rect 19136 34756 19176 34796
rect 1708 34588 1748 34628
rect 1900 34588 1940 34628
rect 9772 34588 9812 34628
rect 10060 34588 10100 34628
rect 16972 34588 17012 34628
rect 19756 34588 19796 34628
rect 9580 34504 9620 34544
rect 17644 34504 17684 34544
rect 1516 34420 1556 34460
rect 2092 34420 2132 34460
rect 17452 34420 17492 34460
rect 19948 34420 19988 34460
rect 2380 34336 2420 34376
rect 2476 34336 2516 34376
rect 2860 34336 2900 34376
rect 2956 34336 2996 34376
rect 3436 34336 3476 34376
rect 3964 34345 4004 34385
rect 4492 34336 4532 34376
rect 5740 34336 5780 34376
rect 6220 34336 6260 34376
rect 6316 34336 6356 34376
rect 6508 34336 6548 34376
rect 7756 34336 7796 34376
rect 8908 34336 8948 34376
rect 9196 34336 9236 34376
rect 9292 34336 9332 34376
rect 9868 34325 9908 34365
rect 10252 34336 10292 34376
rect 11500 34336 11540 34376
rect 11692 34336 11732 34376
rect 12940 34336 12980 34376
rect 13420 34336 13460 34376
rect 13516 34336 13556 34376
rect 13900 34336 13940 34376
rect 13996 34336 14036 34376
rect 14476 34336 14516 34376
rect 15004 34345 15044 34385
rect 15532 34336 15572 34376
rect 16780 34336 16820 34376
rect 17836 34336 17876 34376
rect 18028 34336 18068 34376
rect 18124 34336 18164 34376
rect 18316 34336 18356 34376
rect 19564 34336 19604 34376
rect 7948 34252 7988 34292
rect 13132 34252 13172 34292
rect 4108 34168 4148 34208
rect 4300 34168 4340 34208
rect 6028 34168 6068 34208
rect 8524 34168 8564 34208
rect 15148 34168 15188 34208
rect 20140 34168 20180 34208
rect 4928 34000 4968 34040
rect 5010 34000 5050 34040
rect 5092 34000 5132 34040
rect 5174 34000 5214 34040
rect 5256 34000 5296 34040
rect 20048 34000 20088 34040
rect 20130 34000 20170 34040
rect 20212 34000 20252 34040
rect 20294 34000 20334 34040
rect 20376 34000 20416 34040
rect 5740 33832 5780 33872
rect 13420 33874 13460 33914
rect 15052 33832 15092 33872
rect 11404 33748 11444 33788
rect 16876 33748 16916 33788
rect 1228 33664 1268 33704
rect 2476 33664 2516 33704
rect 3820 33664 3860 33704
rect 4012 33664 4052 33704
rect 4108 33664 4148 33704
rect 4300 33664 4340 33704
rect 5548 33664 5588 33704
rect 5932 33664 5972 33704
rect 7180 33664 7220 33704
rect 7660 33651 7700 33691
rect 7852 33664 7892 33704
rect 8236 33664 8276 33704
rect 8524 33664 8564 33704
rect 8812 33664 8852 33704
rect 8908 33664 8948 33704
rect 9388 33664 9428 33704
rect 9772 33664 9812 33704
rect 9964 33664 10004 33704
rect 11212 33664 11252 33704
rect 11692 33664 11732 33704
rect 11788 33664 11828 33704
rect 12748 33664 12788 33704
rect 13228 33650 13268 33690
rect 13612 33664 13652 33704
rect 14860 33664 14900 33704
rect 15436 33664 15476 33704
rect 16684 33664 16724 33704
rect 17164 33664 17204 33704
rect 17452 33664 17492 33704
rect 17548 33664 17588 33704
rect 18316 33664 18356 33704
rect 19564 33664 19604 33704
rect 7948 33580 7988 33620
rect 8140 33580 8180 33620
rect 9484 33580 9524 33620
rect 9676 33580 9716 33620
rect 12172 33580 12212 33620
rect 12268 33580 12308 33620
rect 19948 33580 19988 33620
rect 4108 33496 4148 33536
rect 8044 33496 8084 33536
rect 9580 33496 9620 33536
rect 2668 33412 2708 33452
rect 5740 33412 5780 33452
rect 7372 33412 7412 33452
rect 7564 33412 7604 33452
rect 9196 33412 9236 33452
rect 17836 33412 17876 33452
rect 19756 33412 19796 33452
rect 20140 33412 20180 33452
rect 3688 33244 3728 33284
rect 3770 33244 3810 33284
rect 3852 33244 3892 33284
rect 3934 33244 3974 33284
rect 4016 33244 4056 33284
rect 18808 33244 18848 33284
rect 18890 33244 18930 33284
rect 18972 33244 19012 33284
rect 19054 33244 19094 33284
rect 19136 33244 19176 33284
rect 5836 33076 5876 33116
rect 9292 33076 9332 33116
rect 13324 33076 13364 33116
rect 9484 32992 9524 33032
rect 3148 32908 3188 32948
rect 2140 32833 2180 32873
rect 2668 32824 2708 32864
rect 3244 32824 3284 32864
rect 3628 32824 3668 32864
rect 3724 32824 3764 32864
rect 4396 32824 4436 32864
rect 5644 32824 5684 32864
rect 6124 32824 6164 32864
rect 6220 32824 6260 32864
rect 6412 32824 6452 32864
rect 6508 32824 6548 32864
rect 6609 32824 6649 32864
rect 6988 32824 7028 32864
rect 8236 32824 8276 32864
rect 8716 32824 8756 32864
rect 8812 32824 8852 32864
rect 9004 32824 9044 32864
rect 9100 32824 9140 32864
rect 9292 32824 9332 32864
rect 9484 32824 9524 32864
rect 9676 32824 9716 32864
rect 9772 32824 9812 32864
rect 9964 32824 10004 32864
rect 10156 32824 10196 32864
rect 11884 32824 11924 32864
rect 13132 32824 13172 32864
rect 14092 32824 14132 32864
rect 15340 32824 15380 32864
rect 15820 32824 15860 32864
rect 15916 32824 15956 32864
rect 16300 32824 16340 32864
rect 16396 32824 16436 32864
rect 16876 32824 16916 32864
rect 17356 32829 17396 32869
rect 17932 32824 17972 32864
rect 19180 32824 19220 32864
rect 19468 32824 19508 32864
rect 19756 32824 19796 32864
rect 19852 32824 19892 32864
rect 10060 32740 10100 32780
rect 15532 32740 15572 32780
rect 17740 32740 17780 32780
rect 1996 32656 2036 32696
rect 6604 32656 6644 32696
rect 8428 32656 8468 32696
rect 17548 32656 17588 32696
rect 20140 32614 20180 32654
rect 4928 32488 4968 32528
rect 5010 32488 5050 32528
rect 5092 32488 5132 32528
rect 5174 32488 5214 32528
rect 5256 32488 5296 32528
rect 20048 32488 20088 32528
rect 20130 32488 20170 32528
rect 20212 32488 20252 32528
rect 20294 32488 20334 32528
rect 20376 32488 20416 32528
rect 6124 32320 6164 32360
rect 8236 32320 8276 32360
rect 17644 32320 17684 32360
rect 2092 32152 2132 32192
rect 3340 32152 3380 32192
rect 4204 32152 4244 32192
rect 5452 32152 5492 32192
rect 5836 32152 5876 32192
rect 5932 32152 5972 32192
rect 6316 32152 6356 32192
rect 7564 32152 7604 32192
rect 7948 32152 7988 32192
rect 8044 32152 8084 32192
rect 8716 32152 8756 32192
rect 9964 32152 10004 32192
rect 12940 32152 12980 32192
rect 14188 32152 14228 32192
rect 14572 32152 14612 32192
rect 15916 32152 15956 32192
rect 16012 32152 16052 32192
rect 16972 32152 17012 32192
rect 17452 32147 17492 32187
rect 18124 32152 18164 32192
rect 19084 32152 19124 32192
rect 16396 32068 16436 32108
rect 16492 32068 16532 32108
rect 19276 32068 19316 32108
rect 19660 32057 19700 32097
rect 20044 32068 20084 32108
rect 19468 31984 19508 32024
rect 19852 31984 19892 32024
rect 3532 31900 3572 31940
rect 5644 31900 5684 31940
rect 7756 31900 7796 31940
rect 10156 31900 10196 31940
rect 14380 31900 14420 31940
rect 14668 31900 14708 31940
rect 20236 31900 20276 31940
rect 3688 31732 3728 31772
rect 3770 31732 3810 31772
rect 3852 31732 3892 31772
rect 3934 31732 3974 31772
rect 4016 31732 4056 31772
rect 18808 31732 18848 31772
rect 18890 31732 18930 31772
rect 18972 31732 19012 31772
rect 19054 31732 19094 31772
rect 19136 31732 19176 31772
rect 17164 31564 17204 31604
rect 14188 31480 14228 31520
rect 6508 31396 6548 31436
rect 2668 31312 2708 31352
rect 3916 31312 3956 31352
rect 4300 31312 4340 31352
rect 5548 31312 5588 31352
rect 6028 31312 6068 31352
rect 6124 31312 6164 31352
rect 6604 31354 6644 31394
rect 8908 31396 8948 31436
rect 7084 31312 7124 31352
rect 7564 31317 7604 31357
rect 8332 31312 8372 31352
rect 8428 31312 8468 31352
rect 9916 31354 9956 31394
rect 10924 31396 10964 31436
rect 11020 31396 11060 31436
rect 17644 31396 17684 31436
rect 19660 31396 19700 31436
rect 20044 31396 20084 31436
rect 8812 31312 8852 31352
rect 9388 31312 9428 31352
rect 10444 31312 10484 31352
rect 10540 31312 10580 31352
rect 11500 31312 11540 31352
rect 12028 31321 12068 31361
rect 12748 31312 12788 31352
rect 13996 31312 14036 31352
rect 14380 31312 14420 31352
rect 14476 31312 14516 31352
rect 14668 31312 14708 31352
rect 14764 31312 14804 31352
rect 14865 31312 14905 31352
rect 15148 31312 15188 31352
rect 15244 31312 15284 31352
rect 17164 31312 17204 31352
rect 17356 31312 17396 31352
rect 17452 31312 17492 31352
rect 18124 31312 18164 31352
rect 18220 31312 18260 31352
rect 18316 31312 18356 31352
rect 18700 31312 18740 31352
rect 18796 31312 18836 31352
rect 18892 31312 18932 31352
rect 19180 31312 19220 31352
rect 19276 31312 19316 31352
rect 19372 31312 19412 31352
rect 4108 31144 4148 31184
rect 5740 31144 5780 31184
rect 7756 31144 7796 31184
rect 10060 31144 10100 31184
rect 12172 31144 12212 31184
rect 14860 31144 14900 31184
rect 15436 31144 15476 31184
rect 17836 31144 17876 31184
rect 18508 31144 18548 31184
rect 18988 31144 19028 31184
rect 19468 31144 19508 31184
rect 19852 31144 19892 31184
rect 20236 31144 20276 31184
rect 4928 30976 4968 31016
rect 5010 30976 5050 31016
rect 5092 30976 5132 31016
rect 5174 30976 5214 31016
rect 5256 30976 5296 31016
rect 20048 30976 20088 31016
rect 20130 30976 20170 31016
rect 20212 30976 20252 31016
rect 20294 30976 20334 31016
rect 20376 30976 20416 31016
rect 4012 30808 4052 30848
rect 6508 30808 6548 30848
rect 8812 30808 8852 30848
rect 10444 30808 10484 30848
rect 12268 30808 12308 30848
rect 16492 30808 16532 30848
rect 18604 30724 18644 30764
rect 2284 30640 2324 30680
rect 2380 30640 2420 30680
rect 3340 30640 3380 30680
rect 3820 30635 3860 30675
rect 4780 30640 4820 30680
rect 4876 30640 4916 30680
rect 5356 30640 5396 30680
rect 5836 30640 5876 30680
rect 6316 30635 6356 30675
rect 8524 30640 8564 30680
rect 8620 30640 8660 30680
rect 9004 30640 9044 30680
rect 10252 30640 10292 30680
rect 10828 30640 10868 30680
rect 12076 30640 12116 30680
rect 12460 30640 12500 30680
rect 13996 30640 14036 30680
rect 14188 30640 14228 30680
rect 14284 30640 14324 30680
rect 14476 30640 14516 30680
rect 15724 30640 15764 30680
rect 16300 30640 16340 30680
rect 16588 30640 16628 30680
rect 16876 30640 16916 30680
rect 16972 30640 17012 30680
rect 17932 30640 17972 30680
rect 18412 30626 18452 30666
rect 18796 30640 18836 30680
rect 20044 30640 20084 30680
rect 2764 30556 2804 30596
rect 2860 30556 2900 30596
rect 5260 30556 5300 30596
rect 17356 30556 17396 30596
rect 17452 30556 17492 30596
rect 14284 30472 14324 30512
rect 12556 30388 12596 30428
rect 15916 30388 15956 30428
rect 20236 30388 20276 30428
rect 3688 30220 3728 30260
rect 3770 30220 3810 30260
rect 3852 30220 3892 30260
rect 3934 30220 3974 30260
rect 4016 30220 4056 30260
rect 18808 30220 18848 30260
rect 18890 30220 18930 30260
rect 18972 30220 19012 30260
rect 19054 30220 19094 30260
rect 19136 30220 19176 30260
rect 11884 30052 11924 30092
rect 17164 30052 17204 30092
rect 18892 30052 18932 30092
rect 5932 29968 5972 30008
rect 13516 29968 13556 30008
rect 1324 29800 1364 29840
rect 2572 29800 2612 29840
rect 3532 29800 3572 29840
rect 4780 29800 4820 29840
rect 5452 29800 5492 29840
rect 5548 29800 5588 29840
rect 5740 29800 5780 29840
rect 5932 29800 5972 29840
rect 6220 29800 6260 29840
rect 6700 29800 6740 29840
rect 7948 29800 7988 29840
rect 8332 29800 8372 29840
rect 8716 29800 8756 29840
rect 8812 29800 8852 29840
rect 9004 29800 9044 29840
rect 9196 29800 9236 29840
rect 9388 29800 9428 29840
rect 9484 29800 9524 29840
rect 10060 29800 10100 29840
rect 10252 29800 10292 29840
rect 10444 29800 10484 29840
rect 11692 29800 11732 29840
rect 12076 29800 12116 29840
rect 13324 29800 13364 29840
rect 13804 29800 13844 29840
rect 13900 29800 13940 29840
rect 14284 29800 14324 29840
rect 14380 29800 14420 29840
rect 14860 29800 14900 29840
rect 15340 29814 15380 29854
rect 15724 29800 15764 29840
rect 16972 29800 17012 29840
rect 17452 29800 17492 29840
rect 18700 29800 18740 29840
rect 19276 29800 19316 29840
rect 8140 29716 8180 29756
rect 15532 29716 15572 29756
rect 2764 29632 2804 29672
rect 4972 29632 5012 29672
rect 5644 29632 5684 29672
rect 8428 29632 8468 29672
rect 8908 29632 8948 29672
rect 9292 29632 9332 29672
rect 10156 29632 10196 29672
rect 19660 29632 19700 29672
rect 4928 29464 4968 29504
rect 5010 29464 5050 29504
rect 5092 29464 5132 29504
rect 5174 29464 5214 29504
rect 5256 29464 5296 29504
rect 20048 29464 20088 29504
rect 20130 29464 20170 29504
rect 20212 29464 20252 29504
rect 20294 29464 20334 29504
rect 20376 29464 20416 29504
rect 7660 29296 7700 29336
rect 8332 29300 8372 29340
rect 8812 29296 8852 29336
rect 18028 29296 18068 29336
rect 18316 29296 18356 29336
rect 18892 29296 18932 29336
rect 13708 29212 13748 29252
rect 15724 29212 15764 29252
rect 19564 29212 19604 29252
rect 2092 29128 2132 29168
rect 3340 29128 3380 29168
rect 3916 29128 3956 29168
rect 5164 29128 5204 29168
rect 5644 29128 5684 29168
rect 5740 29128 5780 29168
rect 5836 29128 5876 29168
rect 6220 29128 6260 29168
rect 6316 29128 6356 29168
rect 6412 29128 6452 29168
rect 6508 29128 6548 29168
rect 7372 29128 7412 29168
rect 7468 29128 7508 29168
rect 8140 29128 8180 29168
rect 8236 29128 8276 29168
rect 8524 29128 8564 29168
rect 8620 29128 8660 29168
rect 8812 29128 8852 29168
rect 8908 29128 8948 29168
rect 9009 29128 9049 29168
rect 9676 29128 9716 29168
rect 10924 29128 10964 29168
rect 11308 29128 11348 29168
rect 11596 29128 11636 29168
rect 11692 29128 11732 29168
rect 13516 29128 13556 29168
rect 13996 29148 14036 29188
rect 14092 29148 14132 29188
rect 14476 29128 14516 29168
rect 12268 29086 12308 29126
rect 14572 29128 14612 29168
rect 15052 29128 15092 29168
rect 15532 29114 15572 29154
rect 16588 29128 16628 29168
rect 17836 29128 17876 29168
rect 18220 29128 18260 29168
rect 18412 29128 18452 29168
rect 18508 29128 18548 29168
rect 19180 29128 19220 29168
rect 19468 29128 19508 29168
rect 18700 29044 18740 29084
rect 20044 29044 20084 29084
rect 6028 28960 6068 29000
rect 7852 28960 7892 29000
rect 19852 28960 19892 29000
rect 3532 28876 3572 28916
rect 5356 28876 5396 28916
rect 9484 28876 9524 28916
rect 11980 28876 12020 28916
rect 18028 28876 18068 28916
rect 20236 28876 20276 28916
rect 3688 28708 3728 28748
rect 3770 28708 3810 28748
rect 3852 28708 3892 28748
rect 3934 28708 3974 28748
rect 4016 28708 4056 28748
rect 18808 28708 18848 28748
rect 18890 28708 18930 28748
rect 18972 28708 19012 28748
rect 19054 28708 19094 28748
rect 19136 28708 19176 28748
rect 7180 28540 7220 28580
rect 16108 28540 16148 28580
rect 12172 28456 12212 28496
rect 1996 28372 2036 28412
rect 3916 28372 3956 28412
rect 16972 28372 17012 28412
rect 1420 28288 1460 28328
rect 1516 28288 1556 28328
rect 1900 28288 1940 28328
rect 2476 28288 2516 28328
rect 2956 28302 2996 28342
rect 3436 28288 3476 28328
rect 3532 28288 3572 28328
rect 4012 28288 4052 28328
rect 4492 28288 4532 28328
rect 4972 28302 5012 28342
rect 6988 28330 7028 28370
rect 17068 28372 17108 28412
rect 5740 28288 5780 28328
rect 7468 28307 7508 28347
rect 7564 28288 7604 28328
rect 7948 28288 7988 28328
rect 8044 28288 8084 28328
rect 8524 28288 8564 28328
rect 9004 28302 9044 28342
rect 9484 28288 9524 28328
rect 9580 28288 9620 28328
rect 9964 28288 10004 28328
rect 10060 28288 10100 28328
rect 10540 28288 10580 28328
rect 11020 28293 11060 28333
rect 11404 28288 11444 28328
rect 11788 28288 11828 28328
rect 11884 28288 11924 28328
rect 12364 28288 12404 28328
rect 12556 28288 12596 28328
rect 12652 28288 12692 28328
rect 12844 28288 12884 28328
rect 13036 28288 13076 28328
rect 13132 28288 13172 28328
rect 14476 28288 14516 28328
rect 14668 28288 14708 28328
rect 15916 28288 15956 28328
rect 16492 28288 16532 28328
rect 16588 28288 16628 28328
rect 17548 28288 17588 28328
rect 18028 28302 18068 28342
rect 18508 28288 18548 28328
rect 19756 28288 19796 28328
rect 3148 28204 3188 28244
rect 5164 28204 5204 28244
rect 9196 28204 9236 28244
rect 11212 28204 11252 28244
rect 11500 28120 11540 28160
rect 11692 28116 11732 28156
rect 12460 28120 12500 28160
rect 12940 28120 12980 28160
rect 14380 28120 14420 28160
rect 18220 28120 18260 28160
rect 19948 28120 19988 28160
rect 4928 27952 4968 27992
rect 5010 27952 5050 27992
rect 5092 27952 5132 27992
rect 5174 27952 5214 27992
rect 5256 27952 5296 27992
rect 20048 27952 20088 27992
rect 20130 27952 20170 27992
rect 20212 27952 20252 27992
rect 20294 27952 20334 27992
rect 20376 27952 20416 27992
rect 3340 27784 3380 27824
rect 11884 27784 11924 27824
rect 12364 27784 12404 27824
rect 18508 27784 18548 27824
rect 5836 27700 5876 27740
rect 9100 27700 9140 27740
rect 17164 27700 17204 27740
rect 19564 27700 19604 27740
rect 1708 27616 1748 27656
rect 2956 27616 2996 27656
rect 3532 27616 3572 27656
rect 4780 27616 4820 27656
rect 5452 27616 5492 27656
rect 5740 27616 5780 27656
rect 6700 27616 6740 27656
rect 7948 27616 7988 27656
rect 8524 27616 8564 27656
rect 8812 27616 8852 27656
rect 9004 27616 9044 27656
rect 9388 27605 9428 27645
rect 9580 27616 9620 27656
rect 9676 27616 9716 27656
rect 10444 27616 10484 27656
rect 11692 27616 11732 27656
rect 12076 27616 12116 27656
rect 12172 27616 12212 27656
rect 12268 27616 12308 27656
rect 13516 27616 13556 27656
rect 14764 27616 14804 27656
rect 15148 27616 15188 27656
rect 15244 27616 15284 27656
rect 15340 27616 15380 27656
rect 15436 27616 15476 27656
rect 15724 27616 15764 27656
rect 16972 27616 17012 27656
rect 17548 27616 17588 27656
rect 17836 27616 17876 27656
rect 18124 27616 18164 27656
rect 18220 27616 18260 27656
rect 18316 27616 18356 27656
rect 19180 27616 19220 27656
rect 19468 27616 19508 27656
rect 18700 27532 18740 27572
rect 6124 27448 6164 27488
rect 8140 27448 8180 27488
rect 8812 27448 8852 27488
rect 17836 27448 17876 27488
rect 18892 27448 18932 27488
rect 3148 27364 3188 27404
rect 9388 27364 9428 27404
rect 14956 27364 14996 27404
rect 19852 27364 19892 27404
rect 3688 27196 3728 27236
rect 3770 27196 3810 27236
rect 3852 27196 3892 27236
rect 3934 27196 3974 27236
rect 4016 27196 4056 27236
rect 18808 27196 18848 27236
rect 18890 27196 18930 27236
rect 18972 27196 19012 27236
rect 19054 27196 19094 27236
rect 19136 27196 19176 27236
rect 14188 27028 14228 27068
rect 15916 27028 15956 27068
rect 6220 26944 6260 26984
rect 15148 26944 15188 26984
rect 15532 26944 15572 26984
rect 16108 26944 16148 26984
rect 16396 26944 16436 26984
rect 19948 26944 19988 26984
rect 11884 26860 11924 26900
rect 15437 26870 15477 26910
rect 15628 26860 15668 26900
rect 19372 26860 19412 26900
rect 19756 26860 19796 26900
rect 1228 26776 1268 26816
rect 2476 26776 2516 26816
rect 3628 26776 3668 26816
rect 3916 26776 3956 26816
rect 4108 26776 4148 26816
rect 5356 26776 5396 26816
rect 5836 26776 5876 26816
rect 5932 26776 5972 26816
rect 6028 26776 6068 26816
rect 6412 26776 6452 26816
rect 6508 26776 6548 26816
rect 6604 26776 6644 26816
rect 7084 26776 7124 26816
rect 8332 26776 8372 26816
rect 9004 26776 9044 26816
rect 10252 26776 10292 26816
rect 10732 26776 10772 26816
rect 10828 26776 10868 26816
rect 10924 26776 10964 26816
rect 11308 26776 11348 26816
rect 11404 26776 11444 26816
rect 11500 26776 11540 26816
rect 11788 26776 11828 26816
rect 12364 26776 12404 26816
rect 13612 26776 13652 26816
rect 14092 26776 14132 26816
rect 14476 26776 14516 26816
rect 14764 26776 14804 26816
rect 15724 26818 15764 26858
rect 14860 26776 14900 26816
rect 15340 26776 15380 26816
rect 16108 26776 16148 26816
rect 16396 26776 16436 26816
rect 16588 26776 16628 26816
rect 16684 26776 16724 26816
rect 18412 26776 18452 26816
rect 18604 26776 18644 26816
rect 18796 26776 18836 26816
rect 18892 26776 18932 26816
rect 8524 26692 8564 26732
rect 13804 26692 13844 26732
rect 18508 26692 18548 26732
rect 2668 26608 2708 26648
rect 3820 26608 3860 26648
rect 5548 26608 5588 26648
rect 6700 26608 6740 26648
rect 10444 26608 10484 26648
rect 11116 26608 11156 26648
rect 11596 26608 11636 26648
rect 14188 26608 14228 26648
rect 19084 26608 19124 26648
rect 19564 26608 19604 26648
rect 4928 26440 4968 26480
rect 5010 26440 5050 26480
rect 5092 26440 5132 26480
rect 5174 26440 5214 26480
rect 5256 26440 5296 26480
rect 20048 26440 20088 26480
rect 20130 26440 20170 26480
rect 20212 26440 20252 26480
rect 20294 26440 20334 26480
rect 20376 26440 20416 26480
rect 4972 26272 5012 26312
rect 13996 26272 14036 26312
rect 14476 26272 14516 26312
rect 15724 26272 15764 26312
rect 18988 26272 19028 26312
rect 6124 26188 6164 26228
rect 10636 26188 10676 26228
rect 1516 26104 1556 26144
rect 2764 26104 2804 26144
rect 3244 26104 3284 26144
rect 3340 26104 3380 26144
rect 3820 26104 3860 26144
rect 4300 26104 4340 26144
rect 4780 26099 4820 26139
rect 5164 26104 5204 26144
rect 5356 26104 5396 26144
rect 5452 26104 5492 26144
rect 5740 26104 5780 26144
rect 6028 26104 6068 26144
rect 8908 26104 8948 26144
rect 9004 26104 9044 26144
rect 9388 26104 9428 26144
rect 9964 26104 10004 26144
rect 10444 26099 10484 26139
rect 10828 26104 10868 26144
rect 12076 26104 12116 26144
rect 12556 26104 12596 26144
rect 13804 26104 13844 26144
rect 14188 26104 14228 26144
rect 14284 26104 14324 26144
rect 14380 26104 14420 26144
rect 14764 26104 14804 26144
rect 15052 26104 15092 26144
rect 15148 26104 15188 26144
rect 15628 26104 15668 26144
rect 15916 26104 15956 26144
rect 17164 26104 17204 26144
rect 17548 26104 17588 26144
rect 18796 26104 18836 26144
rect 19180 26104 19220 26144
rect 19276 26104 19316 26144
rect 19372 26104 19412 26144
rect 19468 26104 19508 26144
rect 3724 26020 3764 26060
rect 9484 26020 9524 26060
rect 19660 26020 19700 26060
rect 20044 26020 20084 26060
rect 5164 25936 5204 25976
rect 20236 25936 20276 25976
rect 2956 25852 2996 25892
rect 6412 25852 6452 25892
rect 12268 25852 12308 25892
rect 15436 25852 15476 25892
rect 17356 25852 17396 25892
rect 19852 25852 19892 25892
rect 3688 25684 3728 25724
rect 3770 25684 3810 25724
rect 3852 25684 3892 25724
rect 3934 25684 3974 25724
rect 4016 25684 4056 25724
rect 18808 25684 18848 25724
rect 18890 25684 18930 25724
rect 18972 25684 19012 25724
rect 19054 25684 19094 25724
rect 19136 25684 19176 25724
rect 5836 25516 5876 25556
rect 14092 25516 14132 25556
rect 15532 25516 15572 25556
rect 19564 25516 19604 25556
rect 9580 25432 9620 25472
rect 12268 25432 12308 25472
rect 2764 25348 2804 25388
rect 17356 25348 17396 25388
rect 2284 25264 2324 25304
rect 2380 25264 2420 25304
rect 2860 25264 2900 25304
rect 3340 25264 3380 25304
rect 3820 25278 3860 25318
rect 4396 25264 4436 25304
rect 5644 25264 5684 25304
rect 6028 25264 6068 25304
rect 7276 25264 7316 25304
rect 7660 25264 7700 25304
rect 8908 25264 8948 25304
rect 9292 25264 9332 25304
rect 9580 25264 9620 25304
rect 9868 25264 9908 25304
rect 10060 25264 10100 25304
rect 10156 25264 10196 25304
rect 10444 25264 10484 25304
rect 10540 25264 10580 25304
rect 10636 25264 10676 25304
rect 11596 25264 11636 25304
rect 11884 25264 11924 25304
rect 11980 25264 12020 25304
rect 13516 25264 13556 25304
rect 13804 25264 13844 25304
rect 4012 25180 4052 25220
rect 13612 25180 13652 25220
rect 13900 25222 13940 25262
rect 14092 25264 14132 25304
rect 14284 25264 14324 25304
rect 14476 25264 14516 25304
rect 14572 25264 14612 25304
rect 14764 25264 14804 25304
rect 14860 25264 14900 25304
rect 14956 25264 14996 25304
rect 15244 25264 15284 25304
rect 15340 25264 15380 25304
rect 15532 25264 15572 25304
rect 16876 25264 16916 25304
rect 16972 25264 17012 25304
rect 17452 25264 17492 25304
rect 17932 25264 17972 25304
rect 18412 25278 18452 25318
rect 18892 25264 18932 25304
rect 19180 25264 19220 25304
rect 19276 25264 19316 25304
rect 19756 25264 19796 25304
rect 19852 25264 19892 25304
rect 14380 25180 14420 25220
rect 15052 25180 15092 25220
rect 18604 25180 18644 25220
rect 7468 25096 7508 25136
rect 9100 25096 9140 25136
rect 9964 25096 10004 25136
rect 10828 25096 10868 25136
rect 20044 25096 20084 25136
rect 4928 24928 4968 24968
rect 5010 24928 5050 24968
rect 5092 24928 5132 24968
rect 5174 24928 5214 24968
rect 5256 24928 5296 24968
rect 20048 24928 20088 24968
rect 20130 24928 20170 24968
rect 20212 24928 20252 24968
rect 20294 24928 20334 24968
rect 20376 24928 20416 24968
rect 14380 24760 14420 24800
rect 18028 24760 18068 24800
rect 18508 24802 18548 24842
rect 20236 24760 20276 24800
rect 10732 24676 10772 24716
rect 15628 24676 15668 24716
rect 3340 24592 3380 24632
rect 3436 24592 3476 24632
rect 3628 24592 3668 24632
rect 4780 24592 4820 24632
rect 6028 24592 6068 24632
rect 6604 24592 6644 24632
rect 6700 24592 6740 24632
rect 6796 24592 6836 24632
rect 7660 24592 7700 24632
rect 7948 24592 7988 24632
rect 8044 24592 8084 24632
rect 9004 24592 9044 24632
rect 9100 24592 9140 24632
rect 10060 24592 10100 24632
rect 10540 24582 10580 24622
rect 11020 24613 11060 24653
rect 9484 24508 9524 24548
rect 9580 24508 9620 24548
rect 10924 24547 10964 24587
rect 11116 24592 11156 24632
rect 11212 24592 11252 24632
rect 11500 24592 11540 24632
rect 11788 24592 11828 24632
rect 11884 24592 11924 24632
rect 12652 24592 12692 24632
rect 13900 24592 13940 24632
rect 14284 24592 14324 24632
rect 14572 24592 14612 24632
rect 14764 24579 14804 24619
rect 14956 24592 14996 24632
rect 15244 24592 15284 24632
rect 15532 24592 15572 24632
rect 16588 24592 16628 24632
rect 17836 24592 17876 24632
rect 18700 24592 18740 24632
rect 18796 24592 18836 24632
rect 19180 24592 19220 24632
rect 19276 24592 19316 24632
rect 19372 24592 19412 24632
rect 19468 24592 19508 24632
rect 14860 24508 14900 24548
rect 19660 24508 19700 24548
rect 20044 24508 20084 24548
rect 6220 24424 6260 24464
rect 18988 24424 19028 24464
rect 19852 24424 19892 24464
rect 3628 24340 3668 24380
rect 6988 24340 7028 24380
rect 8332 24340 8372 24380
rect 12172 24340 12212 24380
rect 14092 24340 14132 24380
rect 15916 24340 15956 24380
rect 3688 24172 3728 24212
rect 3770 24172 3810 24212
rect 3852 24172 3892 24212
rect 3934 24172 3974 24212
rect 4016 24172 4056 24212
rect 18808 24172 18848 24212
rect 18890 24172 18930 24212
rect 18972 24172 19012 24212
rect 19054 24172 19094 24212
rect 19136 24172 19176 24212
rect 10828 24004 10868 24044
rect 5260 23920 5300 23960
rect 12844 23920 12884 23960
rect 15052 23920 15092 23960
rect 19276 23920 19316 23960
rect 6508 23836 6548 23876
rect 13708 23836 13748 23876
rect 19948 23836 19988 23876
rect 1228 23752 1268 23792
rect 2476 23752 2516 23792
rect 3052 23752 3092 23792
rect 3148 23752 3188 23792
rect 3532 23752 3572 23792
rect 3628 23752 3668 23792
rect 4108 23752 4148 23792
rect 4588 23757 4628 23797
rect 4972 23752 5012 23792
rect 5260 23752 5300 23792
rect 5452 23752 5492 23792
rect 5644 23752 5684 23792
rect 5740 23752 5780 23792
rect 6028 23752 6068 23792
rect 6124 23752 6164 23792
rect 6604 23752 6644 23792
rect 7084 23752 7124 23792
rect 7564 23757 7604 23797
rect 7948 23752 7988 23792
rect 8044 23752 8084 23792
rect 8140 23752 8180 23792
rect 8236 23752 8276 23792
rect 9388 23752 9428 23792
rect 10636 23752 10676 23792
rect 11404 23752 11444 23792
rect 12652 23752 12692 23792
rect 13132 23752 13172 23792
rect 13228 23752 13268 23792
rect 13612 23752 13652 23792
rect 14188 23752 14228 23792
rect 14668 23757 14708 23797
rect 15244 23752 15284 23792
rect 15340 23752 15380 23792
rect 15436 23752 15476 23792
rect 15724 23752 15764 23792
rect 16972 23752 17012 23792
rect 17356 23752 17396 23792
rect 17452 23752 17492 23792
rect 17548 23752 17588 23792
rect 18316 23752 18356 23792
rect 18508 23752 18548 23792
rect 18604 23752 18644 23792
rect 18892 23752 18932 23792
rect 18988 23752 19028 23792
rect 19084 23752 19124 23792
rect 19468 23752 19508 23792
rect 19564 23752 19604 23792
rect 19660 23752 19700 23792
rect 4780 23668 4820 23708
rect 5548 23668 5588 23708
rect 7756 23668 7796 23708
rect 14860 23668 14900 23708
rect 18412 23668 18452 23708
rect 2668 23584 2708 23624
rect 17164 23584 17204 23624
rect 17644 23584 17684 23624
rect 19756 23584 19796 23624
rect 20140 23584 20180 23624
rect 4928 23416 4968 23456
rect 5010 23416 5050 23456
rect 5092 23416 5132 23456
rect 5174 23416 5214 23456
rect 5256 23416 5296 23456
rect 20048 23416 20088 23456
rect 20130 23416 20170 23456
rect 20212 23416 20252 23456
rect 20294 23416 20334 23456
rect 20376 23416 20416 23456
rect 2668 23248 2708 23288
rect 4492 23248 4532 23288
rect 6412 23248 6452 23288
rect 12076 23248 12116 23288
rect 15340 23248 15380 23288
rect 17356 23248 17396 23288
rect 18124 23248 18164 23288
rect 18412 23248 18452 23288
rect 1228 23080 1268 23120
rect 2476 23080 2516 23120
rect 3052 23080 3092 23120
rect 4300 23080 4340 23120
rect 4684 23080 4724 23120
rect 4972 23080 5012 23120
rect 6220 23080 6260 23120
rect 6604 23080 6644 23120
rect 6700 23080 6740 23120
rect 6796 23080 6836 23120
rect 6892 23080 6932 23120
rect 7180 23080 7220 23120
rect 7468 23080 7508 23120
rect 7660 23080 7700 23120
rect 7852 23080 7892 23120
rect 7948 23080 7988 23120
rect 8140 23080 8180 23120
rect 9388 23080 9428 23120
rect 9964 23092 10004 23132
rect 10060 23080 10100 23120
rect 10156 23080 10196 23120
rect 10636 23080 10676 23120
rect 11884 23080 11924 23120
rect 13900 23080 13940 23120
rect 15148 23059 15188 23099
rect 15724 23080 15764 23120
rect 16972 23080 17012 23120
rect 17548 23080 17588 23120
rect 17644 23080 17684 23120
rect 17836 23080 17876 23120
rect 17932 23080 17972 23120
rect 18028 23080 18068 23120
rect 18604 23059 18644 23099
rect 19852 23080 19892 23120
rect 7468 22912 7508 22952
rect 17164 22912 17204 22952
rect 4780 22828 4820 22868
rect 7660 22828 7700 22868
rect 9580 22828 9620 22868
rect 9772 22828 9812 22868
rect 3688 22660 3728 22700
rect 3770 22660 3810 22700
rect 3852 22660 3892 22700
rect 3934 22660 3974 22700
rect 4016 22660 4056 22700
rect 18808 22660 18848 22700
rect 18890 22660 18930 22700
rect 18972 22660 19012 22700
rect 19054 22660 19094 22700
rect 19136 22660 19176 22700
rect 3148 22492 3188 22532
rect 3340 22408 3380 22448
rect 4300 22408 4340 22448
rect 6508 22408 6548 22448
rect 7468 22408 7508 22448
rect 12364 22408 12404 22448
rect 19852 22408 19892 22448
rect 8524 22324 8564 22364
rect 13708 22324 13748 22364
rect 2476 22240 2516 22280
rect 2764 22240 2804 22280
rect 2860 22240 2900 22280
rect 3724 22240 3764 22280
rect 4012 22240 4052 22280
rect 4588 22240 4628 22280
rect 4684 22240 4724 22280
rect 5068 22240 5108 22280
rect 6316 22240 6356 22280
rect 6796 22240 6836 22280
rect 7084 22240 7124 22280
rect 8044 22240 8084 22280
rect 8140 22240 8180 22280
rect 8620 22240 8660 22280
rect 9100 22240 9140 22280
rect 9580 22245 9620 22285
rect 9964 22240 10004 22280
rect 11212 22240 11252 22280
rect 11692 22240 11732 22280
rect 11980 22240 12020 22280
rect 13228 22240 13268 22280
rect 13324 22240 13364 22280
rect 13804 22240 13844 22280
rect 14284 22240 14324 22280
rect 14764 22245 14804 22285
rect 15244 22240 15284 22280
rect 15340 22240 15380 22280
rect 15436 22240 15476 22280
rect 15820 22240 15860 22280
rect 15916 22240 15956 22280
rect 16012 22240 16052 22280
rect 17164 22240 17204 22280
rect 17260 22240 17300 22280
rect 17644 22240 17684 22280
rect 17740 22240 17780 22280
rect 18220 22240 18260 22280
rect 18700 22254 18740 22294
rect 19180 22240 19220 22280
rect 19468 22240 19508 22280
rect 19564 22240 19604 22280
rect 3628 22156 3668 22196
rect 7180 22156 7220 22196
rect 11404 22156 11444 22196
rect 12076 22156 12116 22196
rect 18892 22156 18932 22196
rect 4780 22014 4820 22054
rect 9772 22030 9812 22070
rect 14956 22072 14996 22112
rect 15628 22072 15668 22112
rect 16108 22072 16148 22112
rect 4928 21904 4968 21944
rect 5010 21904 5050 21944
rect 5092 21904 5132 21944
rect 5174 21904 5214 21944
rect 5256 21904 5296 21944
rect 20048 21904 20088 21944
rect 20130 21904 20170 21944
rect 20212 21904 20252 21944
rect 20294 21904 20334 21944
rect 20376 21904 20416 21944
rect 3244 21794 3284 21834
rect 3052 21736 3092 21776
rect 4492 21736 4532 21776
rect 7564 21736 7604 21776
rect 14380 21736 14420 21776
rect 18316 21736 18356 21776
rect 20140 21736 20180 21776
rect 2668 21652 2708 21692
rect 10732 21652 10772 21692
rect 12748 21652 12788 21692
rect 15628 21652 15668 21692
rect 17548 21652 17588 21692
rect 1228 21568 1268 21608
rect 2476 21568 2516 21608
rect 2956 21568 2996 21608
rect 3436 21568 3476 21608
rect 3340 21526 3380 21566
rect 3916 21568 3956 21608
rect 4300 21568 4340 21608
rect 4588 21568 4628 21608
rect 4780 21568 4820 21608
rect 4012 21484 4052 21524
rect 4684 21526 4724 21566
rect 5068 21568 5108 21608
rect 6316 21568 6356 21608
rect 6700 21568 6740 21608
rect 7084 21568 7124 21608
rect 7276 21568 7316 21608
rect 7756 21568 7796 21608
rect 9004 21568 9044 21608
rect 9292 21568 9332 21608
rect 10540 21568 10580 21608
rect 11020 21568 11060 21608
rect 11116 21568 11156 21608
rect 11500 21568 11540 21608
rect 11596 21568 11636 21608
rect 12076 21568 12116 21608
rect 12940 21568 12980 21608
rect 14188 21568 14228 21608
rect 14572 21568 14612 21608
rect 4204 21484 4244 21524
rect 6796 21484 6836 21524
rect 6988 21484 7028 21524
rect 12604 21526 12644 21566
rect 14860 21568 14900 21608
rect 15244 21568 15284 21608
rect 15532 21568 15572 21608
rect 16108 21568 16148 21608
rect 17356 21568 17396 21608
rect 18124 21568 18164 21608
rect 18412 21568 18452 21608
rect 18700 21568 18740 21608
rect 19948 21568 19988 21608
rect 3724 21400 3764 21440
rect 4108 21400 4148 21440
rect 6508 21400 6548 21440
rect 6892 21400 6932 21440
rect 15916 21400 15956 21440
rect 3052 21316 3092 21356
rect 7372 21316 7412 21356
rect 14860 21316 14900 21356
rect 3688 21148 3728 21188
rect 3770 21148 3810 21188
rect 3852 21148 3892 21188
rect 3934 21148 3974 21188
rect 4016 21148 4056 21188
rect 18808 21148 18848 21188
rect 18890 21148 18930 21188
rect 18972 21148 19012 21188
rect 19054 21148 19094 21188
rect 19136 21148 19176 21188
rect 2668 20980 2708 21020
rect 4972 20980 5012 21020
rect 6412 20980 6452 21020
rect 7852 20980 7892 21020
rect 12748 20980 12788 21020
rect 14764 20980 14804 21020
rect 14956 20980 14996 21020
rect 4108 20896 4148 20936
rect 4300 20896 4340 20936
rect 7372 20896 7412 20936
rect 17836 20812 17876 20852
rect 17932 20812 17972 20852
rect 1228 20728 1268 20768
rect 2476 20728 2516 20768
rect 2956 20728 2996 20768
rect 3052 20728 3092 20768
rect 3148 20728 3188 20768
rect 3244 20728 3284 20768
rect 3532 20728 3572 20768
rect 3628 20728 3668 20768
rect 3820 20728 3860 20768
rect 4108 20728 4148 20768
rect 4588 20728 4628 20768
rect 4684 20728 4724 20768
rect 4780 20728 4820 20768
rect 5068 20728 5108 20768
rect 5548 20728 5588 20768
rect 5644 20728 5684 20768
rect 5740 20728 5780 20768
rect 6028 20728 6068 20768
rect 6124 20728 6164 20768
rect 6700 20728 6740 20768
rect 6988 20728 7028 20768
rect 7084 20728 7124 20768
rect 7564 20728 7604 20768
rect 7660 20728 7700 20768
rect 7852 20728 7892 20768
rect 9388 20728 9428 20768
rect 9484 20728 9524 20768
rect 9580 20728 9620 20768
rect 11308 20728 11348 20768
rect 12556 20728 12596 20768
rect 13324 20728 13364 20768
rect 14572 20728 14612 20768
rect 15148 20728 15188 20768
rect 16396 20728 16436 20768
rect 17356 20728 17396 20768
rect 17452 20728 17492 20768
rect 18412 20728 18452 20768
rect 18940 20737 18980 20777
rect 19372 20728 19412 20768
rect 19468 20728 19508 20768
rect 19564 20728 19604 20768
rect 19948 20728 19988 20768
rect 20044 20728 20084 20768
rect 20140 20707 20180 20747
rect 3724 20644 3764 20684
rect 4492 20560 4532 20600
rect 5452 20560 5492 20600
rect 5932 20556 5972 20596
rect 9676 20560 9716 20600
rect 14764 20560 14804 20600
rect 19084 20560 19124 20600
rect 19756 20560 19796 20600
rect 20236 20560 20276 20600
rect 4928 20392 4968 20432
rect 5010 20392 5050 20432
rect 5092 20392 5132 20432
rect 5174 20392 5214 20432
rect 5256 20392 5296 20432
rect 20048 20392 20088 20432
rect 20130 20392 20170 20432
rect 20212 20392 20252 20432
rect 20294 20392 20334 20432
rect 20376 20392 20416 20432
rect 2668 20224 2708 20264
rect 6604 20228 6644 20268
rect 7852 20224 7892 20264
rect 6412 20140 6452 20180
rect 10732 20140 10772 20180
rect 12748 20140 12788 20180
rect 15052 20140 15092 20180
rect 1228 20056 1268 20096
rect 2476 20056 2516 20096
rect 2860 20056 2900 20096
rect 4108 20056 4148 20096
rect 4588 20056 4628 20096
rect 4972 20056 5012 20096
rect 5260 20056 5300 20096
rect 5356 20056 5396 20096
rect 5836 20056 5876 20096
rect 6316 20056 6356 20096
rect 6700 20056 6740 20096
rect 6796 20056 6836 20096
rect 7276 20056 7316 20096
rect 7468 20056 7508 20096
rect 7564 20056 7604 20096
rect 7756 20056 7796 20096
rect 9292 20056 9332 20096
rect 10540 20056 10580 20096
rect 11020 20056 11060 20096
rect 11116 20056 11156 20096
rect 11596 20056 11636 20096
rect 12076 20056 12116 20096
rect 12556 20042 12596 20082
rect 12940 20056 12980 20096
rect 14188 20056 14228 20096
rect 14956 20056 14996 20096
rect 15148 20056 15188 20096
rect 15244 20056 15284 20096
rect 16492 20056 16532 20096
rect 17740 20056 17780 20096
rect 18124 20056 18164 20096
rect 18412 20056 18452 20096
rect 18700 20056 18740 20096
rect 19948 20056 19988 20096
rect 4492 19972 4532 20012
rect 11500 19972 11540 20012
rect 7084 19888 7124 19928
rect 7276 19888 7316 19928
rect 17932 19888 17972 19928
rect 2668 19804 2708 19844
rect 4300 19804 4340 19844
rect 5644 19804 5684 19844
rect 5932 19804 5972 19844
rect 14380 19804 14420 19844
rect 18412 19804 18452 19844
rect 20140 19804 20180 19844
rect 3688 19636 3728 19676
rect 3770 19636 3810 19676
rect 3852 19636 3892 19676
rect 3934 19636 3974 19676
rect 4016 19636 4056 19676
rect 18808 19636 18848 19676
rect 18890 19636 18930 19676
rect 18972 19636 19012 19676
rect 19054 19636 19094 19676
rect 19136 19636 19176 19676
rect 4396 19468 4436 19508
rect 12556 19468 12596 19508
rect 15916 19468 15956 19508
rect 19276 19468 19316 19508
rect 1996 19384 2036 19424
rect 20236 19384 20276 19424
rect 8716 19300 8756 19340
rect 1996 19216 2036 19256
rect 2476 19216 2516 19256
rect 2572 19216 2612 19256
rect 2956 19216 2996 19256
rect 3052 19216 3092 19256
rect 3532 19216 3572 19256
rect 4060 19225 4100 19265
rect 4588 19216 4628 19256
rect 5836 19216 5876 19256
rect 6508 19216 6548 19256
rect 7756 19216 7796 19256
rect 8236 19215 8276 19255
rect 8332 19216 8372 19256
rect 8812 19216 8852 19256
rect 9292 19216 9332 19256
rect 9820 19225 9860 19265
rect 11116 19216 11156 19256
rect 12364 19216 12404 19256
rect 13996 19216 14036 19256
rect 14092 19216 14132 19256
rect 14476 19216 14516 19256
rect 14572 19216 14612 19256
rect 15052 19216 15092 19256
rect 15532 19221 15572 19261
rect 16108 19258 16148 19298
rect 17356 19216 17396 19256
rect 17836 19216 17876 19256
rect 19084 19216 19124 19256
rect 19564 19216 19604 19256
rect 19852 19216 19892 19256
rect 19948 19216 19988 19256
rect 4204 19132 4244 19172
rect 7948 19132 7988 19172
rect 2188 19048 2228 19088
rect 9964 19048 10004 19088
rect 15724 19006 15764 19046
rect 19276 19048 19316 19088
rect 4928 18880 4968 18920
rect 5010 18880 5050 18920
rect 5092 18880 5132 18920
rect 5174 18880 5214 18920
rect 5256 18880 5296 18920
rect 20048 18880 20088 18920
rect 20130 18880 20170 18920
rect 20212 18880 20252 18920
rect 20294 18880 20334 18920
rect 20376 18880 20416 18920
rect 4876 18712 4916 18752
rect 7084 18712 7124 18752
rect 9868 18712 9908 18752
rect 16300 18712 16340 18752
rect 16492 18712 16532 18752
rect 18892 18712 18932 18752
rect 3436 18628 3476 18668
rect 13516 18628 13556 18668
rect 15532 18628 15572 18668
rect 1708 18544 1748 18584
rect 1804 18544 1844 18584
rect 2188 18544 2228 18584
rect 2284 18544 2324 18584
rect 2764 18544 2804 18584
rect 3244 18530 3284 18570
rect 3628 18544 3668 18584
rect 3820 18544 3860 18584
rect 3916 18544 3956 18584
rect 4108 18544 4148 18584
rect 4204 18544 4244 18584
rect 4396 18544 4436 18584
rect 4588 18544 4628 18584
rect 4684 18544 4724 18584
rect 4780 18544 4820 18584
rect 5644 18544 5684 18584
rect 6892 18544 6932 18584
rect 8428 18544 8468 18584
rect 9676 18544 9716 18584
rect 10060 18544 10100 18584
rect 11308 18544 11348 18584
rect 12076 18544 12116 18584
rect 13324 18544 13364 18584
rect 13804 18544 13844 18584
rect 13900 18544 13940 18584
rect 14860 18544 14900 18584
rect 17164 18544 17204 18584
rect 18412 18544 18452 18584
rect 18796 18544 18836 18584
rect 14284 18460 14324 18500
rect 14380 18460 14420 18500
rect 15388 18502 15428 18542
rect 18988 18544 19028 18584
rect 19084 18544 19124 18584
rect 16108 18460 16148 18500
rect 16684 18460 16724 18500
rect 3628 18292 3668 18332
rect 4204 18292 4244 18332
rect 11500 18292 11540 18332
rect 18604 18292 18644 18332
rect 3688 18124 3728 18164
rect 3770 18124 3810 18164
rect 3852 18124 3892 18164
rect 3934 18124 3974 18164
rect 4016 18124 4056 18164
rect 18808 18124 18848 18164
rect 18890 18124 18930 18164
rect 18972 18124 19012 18164
rect 19054 18124 19094 18164
rect 19136 18124 19176 18164
rect 3628 17956 3668 17996
rect 15628 17956 15668 17996
rect 7660 17788 7700 17828
rect 10252 17788 10292 17828
rect 1228 17704 1268 17744
rect 2476 17704 2516 17744
rect 3148 17704 3188 17744
rect 3244 17704 3284 17744
rect 3340 17704 3380 17744
rect 3532 17704 3572 17744
rect 3820 17704 3860 17744
rect 5068 17704 5108 17744
rect 5452 17704 5492 17744
rect 6700 17704 6740 17744
rect 7180 17704 7220 17744
rect 7276 17704 7316 17744
rect 7756 17704 7796 17744
rect 8236 17704 8276 17744
rect 8716 17709 8756 17749
rect 9676 17704 9716 17744
rect 9772 17704 9812 17744
rect 11260 17746 11300 17786
rect 10156 17704 10196 17744
rect 10732 17704 10772 17744
rect 12076 17704 12116 17744
rect 12172 17704 12212 17744
rect 12556 17704 12596 17744
rect 12652 17704 12692 17744
rect 13132 17704 13172 17744
rect 13612 17709 13652 17749
rect 14188 17704 14228 17744
rect 15436 17704 15476 17744
rect 16876 17704 16916 17744
rect 16972 17684 17012 17724
rect 17356 17704 17396 17744
rect 18460 17746 18500 17786
rect 17452 17704 17492 17744
rect 17932 17704 17972 17744
rect 18988 17704 19028 17744
rect 20236 17704 20276 17744
rect 2668 17620 2708 17660
rect 5260 17620 5300 17660
rect 6892 17620 6932 17660
rect 8908 17620 8948 17660
rect 11404 17620 11444 17660
rect 13804 17620 13844 17660
rect 3052 17536 3092 17576
rect 18604 17536 18644 17576
rect 18796 17536 18836 17576
rect 4928 17368 4968 17408
rect 5010 17368 5050 17408
rect 5092 17368 5132 17408
rect 5174 17368 5214 17408
rect 5256 17368 5296 17408
rect 20048 17368 20088 17408
rect 20130 17368 20170 17408
rect 20212 17368 20252 17408
rect 20294 17368 20334 17408
rect 20376 17368 20416 17408
rect 2764 17200 2804 17240
rect 9772 17200 9812 17240
rect 11884 17200 11924 17240
rect 13516 17200 13556 17240
rect 16972 17200 17012 17240
rect 4588 17116 4628 17156
rect 6604 17116 6644 17156
rect 18412 17116 18452 17156
rect 1324 17032 1364 17072
rect 2572 17011 2612 17051
rect 3148 17032 3188 17072
rect 4396 17032 4436 17072
rect 4876 17032 4916 17072
rect 4972 17032 5012 17072
rect 5356 17032 5396 17072
rect 5932 17032 5972 17072
rect 6412 17027 6452 17067
rect 8332 17032 8372 17072
rect 9580 17032 9620 17072
rect 10444 17032 10484 17072
rect 12076 17032 12116 17072
rect 13324 17032 13364 17072
rect 15532 17032 15572 17072
rect 16780 17032 16820 17072
rect 11692 16990 11732 17030
rect 18604 17027 18644 17067
rect 19084 17032 19124 17072
rect 20044 17032 20084 17072
rect 20140 17013 20180 17053
rect 5452 16948 5492 16988
rect 18220 16948 18260 16988
rect 19564 16948 19604 16988
rect 19660 16948 19700 16988
rect 2764 16780 2804 16820
rect 18028 16780 18068 16820
rect 3688 16612 3728 16652
rect 3770 16612 3810 16652
rect 3852 16612 3892 16652
rect 3934 16612 3974 16652
rect 4016 16612 4056 16652
rect 18808 16612 18848 16652
rect 18890 16612 18930 16652
rect 18972 16612 19012 16652
rect 19054 16612 19094 16652
rect 19136 16612 19176 16652
rect 8812 16444 8852 16484
rect 20236 16444 20276 16484
rect 2956 16360 2996 16400
rect 3916 16360 3956 16400
rect 14188 16276 14228 16316
rect 1516 16192 1556 16232
rect 2764 16192 2804 16232
rect 3244 16192 3284 16232
rect 3532 16192 3572 16232
rect 4300 16192 4340 16232
rect 5548 16192 5588 16232
rect 5932 16192 5972 16232
rect 6028 16192 6068 16232
rect 6508 16192 6548 16232
rect 7372 16192 7412 16232
rect 8620 16192 8660 16232
rect 9580 16192 9620 16232
rect 9676 16192 9716 16232
rect 10060 16192 10100 16232
rect 10156 16192 10196 16232
rect 10636 16192 10676 16232
rect 11164 16201 11204 16241
rect 11884 16192 11924 16232
rect 13132 16192 13172 16232
rect 13612 16192 13652 16232
rect 13708 16192 13748 16232
rect 14092 16192 14132 16232
rect 14668 16192 14708 16232
rect 15196 16201 15236 16241
rect 15532 16192 15572 16232
rect 16780 16192 16820 16232
rect 17356 16192 17396 16232
rect 18604 16192 18644 16232
rect 18796 16192 18836 16232
rect 20044 16192 20084 16232
rect 3628 16108 3668 16148
rect 5740 16108 5780 16148
rect 11308 16108 11348 16148
rect 13324 16108 13364 16148
rect 15340 16108 15380 16148
rect 17164 16108 17204 16148
rect 6220 16024 6260 16064
rect 6412 16024 6452 16064
rect 16972 16024 17012 16064
rect 4928 15856 4968 15896
rect 5010 15856 5050 15896
rect 5092 15856 5132 15896
rect 5174 15856 5214 15896
rect 5256 15856 5296 15896
rect 20048 15856 20088 15896
rect 20130 15856 20170 15896
rect 20212 15856 20252 15896
rect 20294 15856 20334 15896
rect 20376 15856 20416 15896
rect 3436 15688 3476 15728
rect 5260 15688 5300 15728
rect 8908 15688 8948 15728
rect 11212 15688 11252 15728
rect 15340 15688 15380 15728
rect 6892 15604 6932 15644
rect 18028 15604 18068 15644
rect 1228 15520 1268 15560
rect 2476 15520 2516 15560
rect 3148 15520 3188 15560
rect 3244 15520 3284 15560
rect 3340 15520 3380 15560
rect 3820 15520 3860 15560
rect 5068 15520 5108 15560
rect 5452 15520 5492 15560
rect 6700 15520 6740 15560
rect 7180 15540 7220 15580
rect 7276 15520 7316 15560
rect 7756 15520 7796 15560
rect 8236 15520 8276 15560
rect 8716 15506 8756 15546
rect 9772 15520 9812 15560
rect 11020 15520 11060 15560
rect 11596 15520 11636 15560
rect 12844 15520 12884 15560
rect 13900 15520 13940 15560
rect 15148 15520 15188 15560
rect 16300 15520 16340 15560
rect 16396 15520 16436 15560
rect 16780 15520 16820 15560
rect 17356 15520 17396 15560
rect 17836 15515 17876 15555
rect 18508 15520 18548 15560
rect 19756 15520 19796 15560
rect 7660 15436 7700 15476
rect 16876 15436 16916 15476
rect 2668 15268 2708 15308
rect 5260 15268 5300 15308
rect 11404 15268 11444 15308
rect 19948 15268 19988 15308
rect 3688 15100 3728 15140
rect 3770 15100 3810 15140
rect 3852 15100 3892 15140
rect 3934 15100 3974 15140
rect 4016 15100 4056 15140
rect 18808 15100 18848 15140
rect 18890 15100 18930 15140
rect 18972 15100 19012 15140
rect 19054 15100 19094 15140
rect 19136 15100 19176 15140
rect 1516 14932 1556 14972
rect 1900 14932 1940 14972
rect 7948 14932 7988 14972
rect 9580 14932 9620 14972
rect 5356 14848 5396 14888
rect 1708 14764 1748 14804
rect 2092 14764 2132 14804
rect 10732 14764 10772 14804
rect 14092 14764 14132 14804
rect 14188 14764 14228 14804
rect 18892 14764 18932 14804
rect 2668 14680 2708 14720
rect 2764 14680 2804 14720
rect 3148 14680 3188 14720
rect 3244 14680 3284 14720
rect 3724 14680 3764 14720
rect 4204 14685 4244 14725
rect 5068 14680 5108 14720
rect 5260 14680 5300 14720
rect 5356 14680 5396 14720
rect 5548 14680 5588 14720
rect 5644 14680 5684 14720
rect 5836 14680 5876 14720
rect 5932 14680 5972 14720
rect 6033 14680 6073 14720
rect 6508 14680 6548 14720
rect 7756 14680 7796 14720
rect 8140 14680 8180 14720
rect 9388 14680 9428 14720
rect 10156 14680 10196 14720
rect 10252 14680 10292 14720
rect 10636 14680 10676 14720
rect 11212 14680 11252 14720
rect 11692 14694 11732 14734
rect 13612 14680 13652 14720
rect 13708 14680 13748 14720
rect 14668 14680 14708 14720
rect 15196 14689 15236 14729
rect 16108 14680 16148 14720
rect 17356 14680 17396 14720
rect 18316 14660 18356 14700
rect 18412 14680 18452 14720
rect 18796 14680 18836 14720
rect 19372 14680 19412 14720
rect 19852 14694 19892 14734
rect 4396 14596 4436 14636
rect 11884 14596 11924 14636
rect 5740 14512 5780 14552
rect 15340 14512 15380 14552
rect 15916 14512 15956 14552
rect 20044 14512 20084 14552
rect 4928 14344 4968 14384
rect 5010 14344 5050 14384
rect 5092 14344 5132 14384
rect 5174 14344 5214 14384
rect 5256 14344 5296 14384
rect 20048 14344 20088 14384
rect 20130 14344 20170 14384
rect 20212 14344 20252 14384
rect 20294 14344 20334 14384
rect 20376 14344 20416 14384
rect 1516 14176 1556 14216
rect 2284 14176 2324 14216
rect 4108 14176 4148 14216
rect 11884 14176 11924 14216
rect 13612 14176 13652 14216
rect 15244 14176 15284 14216
rect 17644 14176 17684 14216
rect 6508 14092 6548 14132
rect 8524 14092 8564 14132
rect 15628 14092 15668 14132
rect 2668 14008 2708 14048
rect 3916 14008 3956 14048
rect 5068 14008 5108 14048
rect 6316 14008 6356 14048
rect 6796 14008 6836 14048
rect 6892 14008 6932 14048
rect 7276 14008 7316 14048
rect 7372 14008 7412 14048
rect 7852 14008 7892 14048
rect 8380 13966 8420 14006
rect 10156 14008 10196 14048
rect 10252 14008 10292 14048
rect 10636 14008 10676 14048
rect 10732 14008 10772 14048
rect 11212 14008 11252 14048
rect 11692 14003 11732 14043
rect 12172 14008 12212 14048
rect 13420 14008 13460 14048
rect 13804 14008 13844 14048
rect 15052 14008 15092 14048
rect 15820 14003 15860 14043
rect 16300 14008 16340 14048
rect 16780 14008 16820 14048
rect 17260 14008 17300 14048
rect 17356 14008 17396 14048
rect 17836 14008 17876 14048
rect 19084 14008 19124 14048
rect 1708 13924 1748 13964
rect 2092 13924 2132 13964
rect 2476 13924 2516 13964
rect 16876 13924 16916 13964
rect 1900 13840 1940 13880
rect 3688 13588 3728 13628
rect 3770 13588 3810 13628
rect 3852 13588 3892 13628
rect 3934 13588 3974 13628
rect 4016 13588 4056 13628
rect 18808 13588 18848 13628
rect 18890 13588 18930 13628
rect 18972 13588 19012 13628
rect 19054 13588 19094 13628
rect 19136 13588 19176 13628
rect 1324 13420 1364 13460
rect 8428 13420 8468 13460
rect 10156 13420 10196 13460
rect 12364 13420 12404 13460
rect 16396 13420 16436 13460
rect 1516 13252 1556 13292
rect 1900 13252 1940 13292
rect 13516 13252 13556 13292
rect 18892 13252 18932 13292
rect 18988 13252 19028 13292
rect 2092 13168 2132 13208
rect 3340 13168 3380 13208
rect 3820 13168 3860 13208
rect 3916 13168 3956 13208
rect 4300 13168 4340 13208
rect 4396 13168 4436 13208
rect 4876 13168 4916 13208
rect 5404 13177 5444 13217
rect 6988 13168 7028 13208
rect 8236 13168 8276 13208
rect 8716 13168 8756 13208
rect 9964 13168 10004 13208
rect 10924 13168 10964 13208
rect 12172 13168 12212 13208
rect 13036 13168 13076 13208
rect 13132 13168 13172 13208
rect 13612 13168 13652 13208
rect 14092 13168 14132 13208
rect 14620 13177 14660 13217
rect 14956 13168 14996 13208
rect 16204 13168 16244 13208
rect 16684 13168 16724 13208
rect 17932 13168 17972 13208
rect 18412 13168 18452 13208
rect 18508 13168 18548 13208
rect 19468 13168 19508 13208
rect 19948 13173 19988 13213
rect 3532 13084 3572 13124
rect 5548 13084 5588 13124
rect 18124 13084 18164 13124
rect 1708 13000 1748 13040
rect 14764 13000 14804 13040
rect 20140 13000 20180 13040
rect 4928 12832 4968 12872
rect 5010 12832 5050 12872
rect 5092 12832 5132 12872
rect 5174 12832 5214 12872
rect 5256 12832 5296 12872
rect 20048 12832 20088 12872
rect 20130 12832 20170 12872
rect 20212 12832 20252 12872
rect 20294 12832 20334 12872
rect 20376 12832 20416 12872
rect 5548 12664 5588 12704
rect 10924 12664 10964 12704
rect 13036 12664 13076 12704
rect 14668 12664 14708 12704
rect 20140 12664 20180 12704
rect 8908 12580 8948 12620
rect 17068 12580 17108 12620
rect 2476 12496 2516 12536
rect 3724 12496 3764 12536
rect 4108 12496 4148 12536
rect 5356 12496 5396 12536
rect 8716 12496 8756 12536
rect 9196 12496 9236 12536
rect 7468 12454 7508 12494
rect 9292 12496 9332 12536
rect 9676 12496 9716 12536
rect 10252 12496 10292 12536
rect 10780 12486 10820 12526
rect 11596 12496 11636 12536
rect 12844 12496 12884 12536
rect 13228 12496 13268 12536
rect 14476 12496 14516 12536
rect 15340 12496 15380 12536
rect 15436 12496 15476 12536
rect 15820 12496 15860 12536
rect 15916 12496 15956 12536
rect 16396 12496 16436 12536
rect 16876 12482 16916 12522
rect 18700 12496 18740 12536
rect 19948 12496 19988 12536
rect 1708 12412 1748 12452
rect 2092 12412 2132 12452
rect 9772 12412 9812 12452
rect 1516 12328 1556 12368
rect 1900 12328 1940 12368
rect 3916 12244 3956 12284
rect 3688 12076 3728 12116
rect 3770 12076 3810 12116
rect 3852 12076 3892 12116
rect 3934 12076 3974 12116
rect 4016 12076 4056 12116
rect 18808 12076 18848 12116
rect 18890 12076 18930 12116
rect 18972 12076 19012 12116
rect 19054 12076 19094 12116
rect 19136 12076 19176 12116
rect 1516 11908 1556 11948
rect 1900 11908 1940 11948
rect 10156 11908 10196 11948
rect 15340 11908 15380 11948
rect 17260 11908 17300 11948
rect 1708 11740 1748 11780
rect 2092 11740 2132 11780
rect 3148 11740 3188 11780
rect 7276 11740 7316 11780
rect 18892 11740 18932 11780
rect 2668 11656 2708 11696
rect 2764 11656 2804 11696
rect 3244 11656 3284 11696
rect 3724 11656 3764 11696
rect 4204 11670 4244 11710
rect 5068 11656 5108 11696
rect 6316 11656 6356 11696
rect 6796 11656 6836 11696
rect 6892 11656 6932 11696
rect 7372 11656 7412 11696
rect 7852 11656 7892 11696
rect 8332 11661 8372 11701
rect 9964 11698 10004 11738
rect 18988 11740 19028 11780
rect 8716 11656 8756 11696
rect 10348 11656 10388 11696
rect 11596 11656 11636 11696
rect 13900 11656 13940 11696
rect 15148 11656 15188 11696
rect 15820 11656 15860 11696
rect 17068 11656 17108 11696
rect 18412 11656 18452 11696
rect 18508 11656 18548 11696
rect 19468 11656 19508 11696
rect 19948 11661 19988 11701
rect 6508 11572 6548 11612
rect 8524 11572 8564 11612
rect 4396 11488 4436 11528
rect 11788 11488 11828 11528
rect 20140 11488 20180 11528
rect 4928 11320 4968 11360
rect 5010 11320 5050 11360
rect 5092 11320 5132 11360
rect 5174 11320 5214 11360
rect 5256 11320 5296 11360
rect 20048 11320 20088 11360
rect 20130 11320 20170 11360
rect 20212 11320 20252 11360
rect 20294 11320 20334 11360
rect 20376 11320 20416 11360
rect 2668 11152 2708 11192
rect 7372 11152 7412 11192
rect 9004 11152 9044 11192
rect 11020 11152 11060 11192
rect 16012 11152 16052 11192
rect 18508 11152 18548 11192
rect 20140 11152 20180 11192
rect 5356 11068 5396 11108
rect 1228 10984 1268 11024
rect 2476 10984 2516 11024
rect 3916 10984 3956 11024
rect 5164 10984 5204 11024
rect 5644 10984 5684 11024
rect 5740 10984 5780 11024
rect 6220 10984 6260 11024
rect 6700 10984 6740 11024
rect 7180 10970 7220 11010
rect 7564 10984 7604 11024
rect 8812 10984 8852 11024
rect 9580 10984 9620 11024
rect 10828 10984 10868 11024
rect 11596 10984 11636 11024
rect 12844 10984 12884 11024
rect 14284 10984 14324 11024
rect 14380 10984 14420 11024
rect 14860 10984 14900 11024
rect 15340 10984 15380 11024
rect 15820 10970 15860 11010
rect 17068 10984 17108 11024
rect 18316 10984 18356 11024
rect 18700 10984 18740 11024
rect 19948 10984 19988 11024
rect 3052 10900 3092 10940
rect 6124 10900 6164 10940
rect 14764 10900 14804 10940
rect 2860 10732 2900 10772
rect 13036 10732 13076 10772
rect 3688 10564 3728 10604
rect 3770 10564 3810 10604
rect 3852 10564 3892 10604
rect 3934 10564 3974 10604
rect 4016 10564 4056 10604
rect 18808 10564 18848 10604
rect 18890 10564 18930 10604
rect 18972 10564 19012 10604
rect 19054 10564 19094 10604
rect 19136 10564 19176 10604
rect 6988 10312 7028 10352
rect 8620 10312 8660 10352
rect 17452 10312 17492 10352
rect 3820 10228 3860 10268
rect 9388 10228 9428 10268
rect 11692 10228 11732 10268
rect 16012 10228 16052 10268
rect 1516 10144 1556 10184
rect 2764 10144 2804 10184
rect 3244 10144 3284 10184
rect 3340 10144 3380 10184
rect 3724 10144 3764 10184
rect 4300 10144 4340 10184
rect 4780 10149 4820 10189
rect 5548 10144 5588 10184
rect 6796 10144 6836 10184
rect 7180 10144 7220 10184
rect 8428 10144 8468 10184
rect 8908 10144 8948 10184
rect 9004 10144 9044 10184
rect 9484 10144 9524 10184
rect 9964 10144 10004 10184
rect 10492 10153 10532 10193
rect 11212 10144 11252 10184
rect 11308 10144 11348 10184
rect 12796 10186 12836 10226
rect 11788 10144 11828 10184
rect 12268 10144 12308 10184
rect 14380 10186 14420 10226
rect 16108 10228 16148 10268
rect 17644 10228 17684 10268
rect 19180 10228 19220 10268
rect 19276 10228 19316 10268
rect 13132 10144 13172 10184
rect 15532 10144 15572 10184
rect 15628 10144 15668 10184
rect 16588 10144 16628 10184
rect 17116 10153 17156 10193
rect 18220 10149 18260 10189
rect 18700 10144 18740 10184
rect 19660 10144 19700 10184
rect 19756 10144 19796 10184
rect 2956 10060 2996 10100
rect 4972 10060 5012 10100
rect 12940 10060 12980 10100
rect 14572 10060 14612 10100
rect 17260 10060 17300 10100
rect 18028 10060 18068 10100
rect 10636 9976 10676 10016
rect 4928 9808 4968 9848
rect 5010 9808 5050 9848
rect 5092 9808 5132 9848
rect 5174 9808 5214 9848
rect 5256 9808 5296 9848
rect 20048 9808 20088 9848
rect 20130 9808 20170 9848
rect 20212 9808 20252 9848
rect 20294 9808 20334 9848
rect 20376 9808 20416 9848
rect 1516 9640 1556 9680
rect 3340 9640 3380 9680
rect 7180 9640 7220 9680
rect 10636 9640 10676 9680
rect 15724 9640 15764 9680
rect 17452 9640 17492 9680
rect 19084 9640 19124 9680
rect 5452 9556 5492 9596
rect 12748 9556 12788 9596
rect 1900 9472 1940 9512
rect 3148 9472 3188 9512
rect 3724 9472 3764 9512
rect 3820 9472 3860 9512
rect 4780 9472 4820 9512
rect 1708 9388 1748 9428
rect 4204 9388 4244 9428
rect 4300 9388 4340 9428
rect 5308 9430 5348 9470
rect 7372 9458 7412 9498
rect 7852 9472 7892 9512
rect 8332 9472 8372 9512
rect 8428 9472 8468 9512
rect 8812 9472 8852 9512
rect 8908 9472 8948 9512
rect 9196 9472 9236 9512
rect 10444 9472 10484 9512
rect 11020 9472 11060 9512
rect 11116 9472 11156 9512
rect 11596 9472 11636 9512
rect 12076 9472 12116 9512
rect 12556 9458 12596 9498
rect 14284 9472 14324 9512
rect 15532 9472 15572 9512
rect 16012 9472 16052 9512
rect 17260 9472 17300 9512
rect 17644 9472 17684 9512
rect 18892 9472 18932 9512
rect 11500 9388 11540 9428
rect 19564 9388 19604 9428
rect 19372 9220 19412 9260
rect 3688 9052 3728 9092
rect 3770 9052 3810 9092
rect 3852 9052 3892 9092
rect 3934 9052 3974 9092
rect 4016 9052 4056 9092
rect 18808 9052 18848 9092
rect 18890 9052 18930 9092
rect 18972 9052 19012 9092
rect 19054 9052 19094 9092
rect 19136 9052 19176 9092
rect 7276 8884 7316 8924
rect 11212 8884 11252 8924
rect 20140 8884 20180 8924
rect 1516 8800 1556 8840
rect 1900 8800 1940 8840
rect 2284 8800 2324 8840
rect 2668 8800 2708 8840
rect 4972 8800 5012 8840
rect 7084 8800 7124 8840
rect 13036 8800 13076 8840
rect 14860 8800 14900 8840
rect 17068 8800 17108 8840
rect 1708 8716 1748 8756
rect 2092 8716 2132 8756
rect 2476 8716 2516 8756
rect 2860 8716 2900 8756
rect 15628 8716 15668 8756
rect 15724 8716 15764 8756
rect 3532 8632 3572 8672
rect 4780 8632 4820 8672
rect 5644 8632 5684 8672
rect 6892 8632 6932 8672
rect 7468 8632 7508 8672
rect 8716 8632 8756 8672
rect 9772 8632 9812 8672
rect 11020 8632 11060 8672
rect 11596 8632 11636 8672
rect 12844 8632 12884 8672
rect 13420 8632 13460 8672
rect 14668 8632 14708 8672
rect 15148 8632 15188 8672
rect 15244 8632 15284 8672
rect 16204 8632 16244 8672
rect 16684 8646 16724 8686
rect 17260 8632 17300 8672
rect 18508 8632 18548 8672
rect 18700 8632 18740 8672
rect 19948 8632 19988 8672
rect 16876 8464 16916 8504
rect 4928 8296 4968 8336
rect 5010 8296 5050 8336
rect 5092 8296 5132 8336
rect 5174 8296 5214 8336
rect 5256 8296 5296 8336
rect 20048 8296 20088 8336
rect 20130 8296 20170 8336
rect 20212 8296 20252 8336
rect 20294 8296 20334 8336
rect 20376 8296 20416 8336
rect 1420 8128 1460 8168
rect 1804 8128 1844 8168
rect 5644 8128 5684 8168
rect 15052 8128 15092 8168
rect 10828 8044 10868 8084
rect 4204 8002 4244 8042
rect 12844 8044 12884 8084
rect 19948 8044 19988 8084
rect 2188 7960 2228 8000
rect 3436 7960 3476 8000
rect 5452 7960 5492 8000
rect 6124 7960 6164 8000
rect 7372 7960 7412 8000
rect 7756 7960 7796 8000
rect 9004 7960 9044 8000
rect 9388 7960 9428 8000
rect 10636 7960 10676 8000
rect 11116 7960 11156 8000
rect 11212 7960 11252 8000
rect 11596 7960 11636 8000
rect 11692 7960 11732 8000
rect 12172 7960 12212 8000
rect 13612 7960 13652 8000
rect 14860 7960 14900 8000
rect 15436 7960 15476 8000
rect 16684 7960 16724 8000
rect 12700 7918 12740 7958
rect 18220 7941 18260 7981
rect 18316 7960 18356 8000
rect 18700 7960 18740 8000
rect 19276 7960 19316 8000
rect 19756 7946 19796 7986
rect 1612 7876 1652 7916
rect 1996 7876 2036 7916
rect 18796 7876 18836 7916
rect 3628 7708 3668 7748
rect 7564 7708 7604 7748
rect 9196 7708 9236 7748
rect 15244 7708 15284 7748
rect 3688 7540 3728 7580
rect 3770 7540 3810 7580
rect 3852 7540 3892 7580
rect 3934 7540 3974 7580
rect 4016 7540 4056 7580
rect 18808 7540 18848 7580
rect 18890 7540 18930 7580
rect 18972 7540 19012 7580
rect 19054 7540 19094 7580
rect 19136 7540 19176 7580
rect 1420 7372 1460 7412
rect 1804 7372 1844 7412
rect 13036 7372 13076 7412
rect 17932 7372 17972 7412
rect 1612 7204 1652 7244
rect 1996 7204 2036 7244
rect 4396 7204 4436 7244
rect 4492 7204 4532 7244
rect 6700 7204 6740 7244
rect 6796 7204 6836 7244
rect 9388 7204 9428 7244
rect 2380 7120 2420 7160
rect 3628 7120 3668 7160
rect 3916 7120 3956 7160
rect 4012 7120 4052 7160
rect 4972 7120 5012 7160
rect 5500 7129 5540 7169
rect 6220 7120 6260 7160
rect 6316 7120 6356 7160
rect 7276 7120 7316 7160
rect 7756 7125 7796 7165
rect 8428 7134 8468 7174
rect 8908 7162 8948 7202
rect 15052 7204 15092 7244
rect 16492 7204 16532 7244
rect 16588 7204 16628 7244
rect 19756 7204 19796 7244
rect 9484 7120 9524 7160
rect 9868 7120 9908 7160
rect 9964 7120 10004 7160
rect 11596 7120 11636 7160
rect 12844 7120 12884 7160
rect 14092 7134 14132 7174
rect 14572 7120 14612 7160
rect 15148 7120 15188 7160
rect 15532 7120 15572 7160
rect 15628 7100 15668 7140
rect 16012 7120 16052 7160
rect 16108 7120 16148 7160
rect 17068 7120 17108 7160
rect 17548 7125 17588 7165
rect 18124 7120 18164 7160
rect 19372 7120 19412 7160
rect 7948 7036 7988 7076
rect 2188 6952 2228 6992
rect 5644 6952 5684 6992
rect 8236 6952 8276 6992
rect 13900 6952 13940 6992
rect 17740 6952 17780 6992
rect 19564 6952 19604 6992
rect 4928 6784 4968 6824
rect 5010 6784 5050 6824
rect 5092 6784 5132 6824
rect 5174 6784 5214 6824
rect 5256 6784 5296 6824
rect 20048 6784 20088 6824
rect 20130 6784 20170 6824
rect 20212 6784 20252 6824
rect 20294 6784 20334 6824
rect 20376 6784 20416 6824
rect 1516 6616 1556 6656
rect 1900 6616 1940 6656
rect 6124 6616 6164 6656
rect 7756 6616 7796 6656
rect 8428 6616 8468 6656
rect 14668 6616 14708 6656
rect 17260 6616 17300 6656
rect 19756 6616 19796 6656
rect 2668 6532 2708 6572
rect 13036 6532 13076 6572
rect 2860 6443 2900 6483
rect 3340 6448 3380 6488
rect 3820 6448 3860 6488
rect 3916 6448 3956 6488
rect 4300 6448 4340 6488
rect 4396 6448 4436 6488
rect 4684 6448 4724 6488
rect 5932 6448 5972 6488
rect 7564 6448 7604 6488
rect 6316 6406 6356 6446
rect 9100 6448 9140 6488
rect 9676 6448 9716 6488
rect 8572 6406 8612 6446
rect 10060 6448 10100 6488
rect 10156 6448 10196 6488
rect 11308 6448 11348 6488
rect 11404 6448 11444 6488
rect 11884 6448 11924 6488
rect 12364 6448 12404 6488
rect 13228 6448 13268 6488
rect 14476 6448 14516 6488
rect 15820 6448 15860 6488
rect 17068 6448 17108 6488
rect 18028 6448 18068 6488
rect 1708 6364 1748 6404
rect 2092 6364 2132 6404
rect 2476 6353 2516 6393
rect 9580 6364 9620 6404
rect 11788 6364 11828 6404
rect 12892 6406 12932 6446
rect 18124 6448 18164 6488
rect 18508 6448 18548 6488
rect 18604 6448 18644 6488
rect 19084 6448 19124 6488
rect 19564 6434 19604 6474
rect 20121 6361 20161 6401
rect 19948 6280 19988 6320
rect 2284 6196 2324 6236
rect 3688 6028 3728 6068
rect 3770 6028 3810 6068
rect 3852 6028 3892 6068
rect 3934 6028 3974 6068
rect 4016 6028 4056 6068
rect 18808 6028 18848 6068
rect 18890 6028 18930 6068
rect 18972 6028 19012 6068
rect 19054 6028 19094 6068
rect 19136 6028 19176 6068
rect 2668 5860 2708 5900
rect 2860 5860 2900 5900
rect 5932 5860 5972 5900
rect 8140 5860 8180 5900
rect 8332 5860 8372 5900
rect 11404 5860 11444 5900
rect 13132 5860 13172 5900
rect 15436 5860 15476 5900
rect 17740 5860 17780 5900
rect 3052 5692 3092 5732
rect 3436 5692 3476 5732
rect 18508 5692 18548 5732
rect 20140 5703 20180 5743
rect 1228 5608 1268 5648
rect 2476 5608 2516 5648
rect 4492 5608 4532 5648
rect 5740 5608 5780 5648
rect 6700 5608 6740 5648
rect 7948 5608 7988 5648
rect 8524 5608 8564 5648
rect 9772 5608 9812 5648
rect 9964 5608 10004 5648
rect 11212 5608 11252 5648
rect 11692 5608 11732 5648
rect 12940 5608 12980 5648
rect 13996 5608 14036 5648
rect 15244 5608 15284 5648
rect 16300 5608 16340 5648
rect 17548 5608 17588 5648
rect 18028 5608 18068 5648
rect 18124 5608 18164 5648
rect 18604 5608 18644 5648
rect 19084 5608 19124 5648
rect 19564 5613 19604 5653
rect 19756 5524 19796 5564
rect 3244 5440 3284 5480
rect 19948 5440 19988 5480
rect 4928 5272 4968 5312
rect 5010 5272 5050 5312
rect 5092 5272 5132 5312
rect 5174 5272 5214 5312
rect 5256 5272 5296 5312
rect 20048 5272 20088 5312
rect 20130 5272 20170 5312
rect 20212 5272 20252 5312
rect 20294 5272 20334 5312
rect 20376 5272 20416 5312
rect 7756 5104 7796 5144
rect 18316 5104 18356 5144
rect 3532 5020 3572 5060
rect 5644 5020 5684 5060
rect 13036 5020 13076 5060
rect 15052 5020 15092 5060
rect 20044 5020 20084 5060
rect 2092 4936 2132 4976
rect 3340 4936 3380 4976
rect 3916 4936 3956 4976
rect 4012 4936 4052 4976
rect 4396 4936 4436 4976
rect 4492 4936 4532 4976
rect 4972 4936 5012 4976
rect 5452 4922 5492 4962
rect 6028 4936 6068 4976
rect 6124 4936 6164 4976
rect 6508 4936 6548 4976
rect 6604 4936 6644 4976
rect 7084 4936 7124 4976
rect 7564 4922 7604 4962
rect 8332 4936 8372 4976
rect 9580 4936 9620 4976
rect 9964 4936 10004 4976
rect 11212 4936 11252 4976
rect 11596 4936 11636 4976
rect 12844 4936 12884 4976
rect 13324 4917 13364 4957
rect 13420 4936 13460 4976
rect 13804 4936 13844 4976
rect 14380 4936 14420 4976
rect 14860 4922 14900 4962
rect 15244 4936 15284 4976
rect 16492 4936 16532 4976
rect 16876 4936 16916 4976
rect 18124 4936 18164 4976
rect 18604 4936 18644 4976
rect 19852 4936 19892 4976
rect 1516 4852 1556 4892
rect 1900 4852 1940 4892
rect 13900 4852 13940 4892
rect 1324 4768 1364 4808
rect 1708 4768 1748 4808
rect 9772 4684 9812 4724
rect 11404 4684 11444 4724
rect 16684 4684 16724 4724
rect 3688 4516 3728 4556
rect 3770 4516 3810 4556
rect 3852 4516 3892 4556
rect 3934 4516 3974 4556
rect 4016 4516 4056 4556
rect 18808 4516 18848 4556
rect 18890 4516 18930 4556
rect 18972 4516 19012 4556
rect 19054 4516 19094 4556
rect 19136 4516 19176 4556
rect 7084 4348 7124 4388
rect 14668 4348 14708 4388
rect 17356 4348 17396 4388
rect 17740 4348 17780 4388
rect 4012 4180 4052 4220
rect 4108 4180 4148 4220
rect 5068 4180 5108 4220
rect 7852 4180 7892 4220
rect 7948 4180 7988 4220
rect 10636 4180 10676 4220
rect 10732 4180 10772 4220
rect 15532 4180 15572 4220
rect 17548 4180 17588 4220
rect 17932 4180 17972 4220
rect 18700 4180 18740 4220
rect 18796 4180 18836 4220
rect 1228 4096 1268 4136
rect 2476 4096 2516 4136
rect 3004 4105 3044 4145
rect 3532 4096 3572 4136
rect 4492 4096 4532 4136
rect 4588 4096 4628 4136
rect 5644 4096 5684 4136
rect 6892 4096 6932 4136
rect 7372 4096 7412 4136
rect 7468 4096 7508 4136
rect 8428 4096 8468 4136
rect 8956 4105 8996 4145
rect 10156 4096 10196 4136
rect 10252 4096 10292 4136
rect 11212 4096 11252 4136
rect 11692 4110 11732 4150
rect 13228 4096 13268 4136
rect 14476 4096 14516 4136
rect 14956 4096 14996 4136
rect 15052 4096 15092 4136
rect 15436 4096 15476 4136
rect 16012 4096 16052 4136
rect 16492 4110 16532 4150
rect 18220 4096 18260 4136
rect 18316 4096 18356 4136
rect 19276 4096 19316 4136
rect 19756 4101 19796 4141
rect 2668 4012 2708 4052
rect 11884 4012 11924 4052
rect 19948 4012 19988 4052
rect 2860 3928 2900 3968
rect 4876 3928 4916 3968
rect 9100 3928 9140 3968
rect 16684 3928 16724 3968
rect 4928 3760 4968 3800
rect 5010 3760 5050 3800
rect 5092 3760 5132 3800
rect 5174 3760 5214 3800
rect 5256 3760 5296 3800
rect 20048 3760 20088 3800
rect 20130 3760 20170 3800
rect 20212 3760 20252 3800
rect 20294 3760 20334 3800
rect 20376 3760 20416 3800
rect 1900 3592 1940 3632
rect 2668 3592 2708 3632
rect 5740 3592 5780 3632
rect 7468 3592 7508 3632
rect 9196 3592 9236 3632
rect 14956 3592 14996 3632
rect 20044 3592 20084 3632
rect 11020 3508 11060 3548
rect 13036 3508 13076 3548
rect 18412 3508 18452 3548
rect 2860 3424 2900 3464
rect 4108 3424 4148 3464
rect 4300 3424 4340 3464
rect 5548 3424 5588 3464
rect 6028 3424 6068 3464
rect 7276 3424 7316 3464
rect 7756 3424 7796 3464
rect 9004 3424 9044 3464
rect 9580 3424 9620 3464
rect 10828 3424 10868 3464
rect 11308 3424 11348 3464
rect 11404 3424 11444 3464
rect 11788 3424 11828 3464
rect 11884 3424 11924 3464
rect 12364 3424 12404 3464
rect 12892 3414 12932 3454
rect 13516 3424 13556 3464
rect 14764 3424 14804 3464
rect 16684 3424 16724 3464
rect 16780 3424 16820 3464
rect 17164 3424 17204 3464
rect 17260 3424 17300 3464
rect 17740 3424 17780 3464
rect 18604 3424 18644 3464
rect 19852 3424 19892 3464
rect 18268 3382 18308 3422
rect 1708 3340 1748 3380
rect 2092 3340 2132 3380
rect 2476 3340 2516 3380
rect 15436 3340 15476 3380
rect 2284 3256 2324 3296
rect 1516 3172 1556 3212
rect 15244 3172 15284 3212
rect 3688 3004 3728 3044
rect 3770 3004 3810 3044
rect 3852 3004 3892 3044
rect 3934 3004 3974 3044
rect 4016 3004 4056 3044
rect 18808 3004 18848 3044
rect 18890 3004 18930 3044
rect 18972 3004 19012 3044
rect 19054 3004 19094 3044
rect 19136 3004 19176 3044
rect 2284 2836 2324 2876
rect 7660 2836 7700 2876
rect 8044 2836 8084 2876
rect 13324 2836 13364 2876
rect 16780 2836 16820 2876
rect 18412 2836 18452 2876
rect 20044 2836 20084 2876
rect 1900 2752 1940 2792
rect 1708 2668 1748 2708
rect 2092 2668 2132 2708
rect 2476 2668 2516 2708
rect 5164 2668 5204 2708
rect 5932 2668 5972 2708
rect 6028 2668 6068 2708
rect 7852 2668 7892 2708
rect 8236 2668 8276 2708
rect 8428 2679 8468 2719
rect 9388 2668 9428 2708
rect 9772 2668 9812 2708
rect 10156 2668 10196 2708
rect 11116 2668 11156 2708
rect 13708 2668 13748 2708
rect 14092 2668 14132 2708
rect 14476 2668 14516 2708
rect 14860 2668 14900 2708
rect 3052 2584 3092 2624
rect 3148 2584 3188 2624
rect 3532 2584 3572 2624
rect 3628 2584 3668 2624
rect 4108 2584 4148 2624
rect 4588 2589 4628 2629
rect 5452 2584 5492 2624
rect 5548 2584 5588 2624
rect 6508 2584 6548 2624
rect 6988 2589 7028 2629
rect 11884 2584 11924 2624
rect 13132 2584 13172 2624
rect 15340 2584 15380 2624
rect 16588 2605 16628 2645
rect 16972 2584 17012 2624
rect 18220 2584 18260 2624
rect 18604 2584 18644 2624
rect 19852 2584 19892 2624
rect 4780 2500 4820 2540
rect 7180 2500 7220 2540
rect 1516 2416 1556 2456
rect 4972 2416 5012 2456
rect 8620 2416 8660 2456
rect 9580 2416 9620 2456
rect 9964 2416 10004 2456
rect 10348 2416 10388 2456
rect 10924 2416 10964 2456
rect 13516 2416 13556 2456
rect 13900 2416 13940 2456
rect 14284 2416 14324 2456
rect 14668 2416 14708 2456
rect 4928 2248 4968 2288
rect 5010 2248 5050 2288
rect 5092 2248 5132 2288
rect 5174 2248 5214 2288
rect 5256 2248 5296 2288
rect 20048 2248 20088 2288
rect 20130 2248 20170 2288
rect 20212 2248 20252 2288
rect 20294 2248 20334 2288
rect 20376 2248 20416 2288
rect 2860 2080 2900 2120
rect 4492 2080 4532 2120
rect 6124 2080 6164 2120
rect 9868 2080 9908 2120
rect 18220 2080 18260 2120
rect 19948 2080 19988 2120
rect 7852 1996 7892 2036
rect 3052 1954 3092 1994
rect 16588 1996 16628 2036
rect 1420 1912 1460 1952
rect 2668 1912 2708 1952
rect 4300 1912 4340 1952
rect 4684 1912 4724 1952
rect 5932 1912 5972 1952
rect 6412 1912 6452 1952
rect 7660 1912 7700 1952
rect 8140 1912 8180 1952
rect 8236 1912 8276 1952
rect 8716 1912 8756 1952
rect 9196 1912 9236 1952
rect 9676 1898 9716 1938
rect 12460 1912 12500 1952
rect 13708 1912 13748 1952
rect 14860 1912 14900 1952
rect 14956 1912 14996 1952
rect 15340 1912 15380 1952
rect 15436 1912 15476 1952
rect 15916 1912 15956 1952
rect 16396 1898 16436 1938
rect 16780 1912 16820 1952
rect 18028 1912 18068 1952
rect 18508 1912 18548 1952
rect 19756 1912 19796 1952
rect 8620 1828 8660 1868
rect 10060 1828 10100 1868
rect 10444 1828 10484 1868
rect 11020 1828 11060 1868
rect 11212 1828 11252 1868
rect 11596 1828 11636 1868
rect 12268 1828 12308 1868
rect 14092 1828 14132 1868
rect 14380 1828 14420 1868
rect 13900 1744 13940 1784
rect 10252 1660 10292 1700
rect 10636 1660 10676 1700
rect 10828 1660 10868 1700
rect 11404 1660 11444 1700
rect 11788 1660 11828 1700
rect 12076 1660 12116 1700
rect 14572 1660 14612 1700
rect 3688 1492 3728 1532
rect 3770 1492 3810 1532
rect 3852 1492 3892 1532
rect 3934 1492 3974 1532
rect 4016 1492 4056 1532
rect 18808 1492 18848 1532
rect 18890 1492 18930 1532
rect 18972 1492 19012 1532
rect 19054 1492 19094 1532
rect 19136 1492 19176 1532
rect 9676 1324 9716 1364
rect 16876 1324 16916 1364
rect 1516 1240 1556 1280
rect 1900 1240 1940 1280
rect 2284 1240 2324 1280
rect 4684 1240 4724 1280
rect 6796 1240 6836 1280
rect 7852 1240 7892 1280
rect 1708 1156 1748 1196
rect 2092 1156 2132 1196
rect 2476 1156 2516 1196
rect 2860 1156 2900 1196
rect 4876 1156 4916 1196
rect 7468 1156 7508 1196
rect 8044 1156 8084 1196
rect 10060 1156 10100 1196
rect 10444 1156 10484 1196
rect 10828 1156 10868 1196
rect 11212 1156 11252 1196
rect 12652 1156 12692 1196
rect 13036 1156 13076 1196
rect 13420 1156 13460 1196
rect 13804 1156 13844 1196
rect 14284 1156 14324 1196
rect 14668 1156 14708 1196
rect 15052 1156 15092 1196
rect 17356 1156 17396 1196
rect 18412 1156 18452 1196
rect 3244 1072 3284 1112
rect 4492 1072 4532 1112
rect 5356 1072 5396 1112
rect 6604 1072 6644 1112
rect 8236 1072 8276 1112
rect 9484 1072 9524 1112
rect 15436 1072 15476 1112
rect 16684 1072 16724 1112
rect 2668 904 2708 944
rect 5068 904 5108 944
rect 7660 904 7700 944
rect 10252 904 10292 944
rect 10636 904 10676 944
rect 11020 904 11060 944
rect 11404 904 11444 944
rect 12460 904 12500 944
rect 12844 904 12884 944
rect 13228 904 13268 944
rect 13612 904 13652 944
rect 14092 904 14132 944
rect 14476 904 14516 944
rect 14860 904 14900 944
rect 17164 904 17204 944
rect 18220 904 18260 944
rect 4928 736 4968 776
rect 5010 736 5050 776
rect 5092 736 5132 776
rect 5174 736 5214 776
rect 5256 736 5296 776
rect 20048 736 20088 776
rect 20130 736 20170 776
rect 20212 736 20252 776
rect 20294 736 20334 776
rect 20376 736 20416 776
<< metal2 >>
rect 1420 42953 1652 42988
rect 1420 42948 1653 42953
rect 1324 41096 1364 41107
rect 1324 41021 1364 41056
rect 1323 41012 1365 41021
rect 1323 40972 1324 41012
rect 1364 40972 1365 41012
rect 1323 40963 1365 40972
rect 1323 40760 1365 40769
rect 1323 40720 1324 40760
rect 1364 40720 1365 40760
rect 1323 40711 1365 40720
rect 1324 40349 1364 40711
rect 1323 40340 1365 40349
rect 1323 40300 1324 40340
rect 1364 40300 1365 40340
rect 1323 40291 1365 40300
rect 1228 40256 1268 40265
rect 1228 40172 1268 40216
rect 1228 40132 1364 40172
rect 1324 39593 1364 40132
rect 1323 39584 1365 39593
rect 1323 39544 1324 39584
rect 1364 39544 1365 39584
rect 1323 39535 1365 39544
rect 1131 39500 1173 39509
rect 1131 39460 1132 39500
rect 1172 39460 1173 39500
rect 1131 39451 1173 39460
rect 1132 39089 1172 39451
rect 1324 39450 1364 39535
rect 1131 39080 1173 39089
rect 1131 39040 1132 39080
rect 1172 39040 1173 39080
rect 1131 39031 1173 39040
rect 1323 38996 1365 39005
rect 1323 38956 1324 38996
rect 1364 38956 1365 38996
rect 1323 38947 1365 38956
rect 1324 38862 1364 38947
rect 1323 38492 1365 38501
rect 1323 38452 1324 38492
rect 1364 38452 1365 38492
rect 1323 38443 1365 38452
rect 1228 38240 1268 38249
rect 1324 38240 1364 38443
rect 1268 38200 1364 38240
rect 1228 38191 1268 38200
rect 1420 37904 1460 42948
rect 1611 42944 1653 42948
rect 1611 42904 1612 42944
rect 1652 42904 1653 42944
rect 1784 42944 1864 43008
rect 1784 42928 1804 42944
rect 1611 42895 1653 42904
rect 1803 42904 1804 42928
rect 1844 42928 1864 42944
rect 1976 42928 2056 43008
rect 2168 42928 2248 43008
rect 2360 42928 2440 43008
rect 2552 42928 2632 43008
rect 2744 42928 2824 43008
rect 2936 42928 3016 43008
rect 3128 42928 3208 43008
rect 3320 42928 3400 43008
rect 3512 42928 3592 43008
rect 3704 42928 3784 43008
rect 3896 42928 3976 43008
rect 4088 42928 4168 43008
rect 4280 42928 4360 43008
rect 4472 42928 4552 43008
rect 4664 42928 4744 43008
rect 4856 42928 4936 43008
rect 5048 42928 5128 43008
rect 5240 42928 5320 43008
rect 5432 42928 5512 43008
rect 5624 42928 5704 43008
rect 5816 42928 5896 43008
rect 6008 42928 6088 43008
rect 6200 42928 6280 43008
rect 6392 42928 6472 43008
rect 6584 42928 6664 43008
rect 6776 42928 6856 43008
rect 6968 42928 7048 43008
rect 7160 42928 7240 43008
rect 7352 42928 7432 43008
rect 7544 42928 7624 43008
rect 7736 42928 7816 43008
rect 7928 42928 8008 43008
rect 8120 42928 8200 43008
rect 8312 42928 8392 43008
rect 8504 42928 8584 43008
rect 8696 42928 8776 43008
rect 8888 42928 8968 43008
rect 9080 42928 9160 43008
rect 9272 42928 9352 43008
rect 9464 42928 9544 43008
rect 9656 42928 9736 43008
rect 9848 42928 9928 43008
rect 10040 42928 10120 43008
rect 10232 42928 10312 43008
rect 10424 42928 10504 43008
rect 10616 42928 10696 43008
rect 10808 42928 10888 43008
rect 11000 42928 11080 43008
rect 11192 42928 11272 43008
rect 11384 42928 11464 43008
rect 11576 42928 11656 43008
rect 11768 42928 11848 43008
rect 11960 42928 12040 43008
rect 12152 42928 12232 43008
rect 12344 42928 12424 43008
rect 12536 42928 12616 43008
rect 12728 42928 12808 43008
rect 12920 42928 13000 43008
rect 13112 42928 13192 43008
rect 13304 42928 13384 43008
rect 13496 42928 13576 43008
rect 13688 42928 13768 43008
rect 13880 42928 13960 43008
rect 14072 42928 14152 43008
rect 14264 42928 14344 43008
rect 14456 42928 14536 43008
rect 14648 42928 14728 43008
rect 14840 42928 14920 43008
rect 15032 42928 15112 43008
rect 15224 42928 15304 43008
rect 15416 42928 15496 43008
rect 15608 42928 15688 43008
rect 15800 42928 15880 43008
rect 15992 42928 16072 43008
rect 16184 42928 16264 43008
rect 16376 42928 16456 43008
rect 16568 42928 16648 43008
rect 16760 42928 16840 43008
rect 16952 42928 17032 43008
rect 17144 42928 17224 43008
rect 17336 42928 17416 43008
rect 17528 42928 17608 43008
rect 17720 42928 17800 43008
rect 17912 42928 17992 43008
rect 18104 42928 18184 43008
rect 18296 42928 18376 43008
rect 18488 42928 18568 43008
rect 18680 42928 18760 43008
rect 18872 42928 18952 43008
rect 19064 42928 19144 43008
rect 19256 42928 19336 43008
rect 19448 42928 19528 43008
rect 1844 42904 1845 42928
rect 1803 42895 1845 42904
rect 1803 42356 1845 42365
rect 1803 42316 1804 42356
rect 1844 42316 1845 42356
rect 1803 42307 1845 42316
rect 1611 42272 1653 42281
rect 1611 42232 1612 42272
rect 1652 42232 1653 42272
rect 1611 42223 1653 42232
rect 1515 41012 1557 41021
rect 1515 40972 1516 41012
rect 1556 40972 1557 41012
rect 1515 40963 1557 40972
rect 1516 40517 1556 40963
rect 1515 40508 1557 40517
rect 1515 40468 1516 40508
rect 1556 40468 1557 40508
rect 1515 40459 1557 40468
rect 1515 40340 1557 40349
rect 1515 40300 1516 40340
rect 1556 40300 1557 40340
rect 1515 40291 1557 40300
rect 1516 39836 1556 40291
rect 1612 39920 1652 42223
rect 1707 41180 1749 41189
rect 1707 41140 1708 41180
rect 1748 41140 1749 41180
rect 1707 41131 1749 41140
rect 1708 41046 1748 41131
rect 1708 40676 1748 40685
rect 1804 40676 1844 42307
rect 1899 41180 1941 41189
rect 1899 41140 1900 41180
rect 1940 41140 1941 41180
rect 1899 41131 1941 41140
rect 1748 40636 1844 40676
rect 1708 40627 1748 40636
rect 1803 40424 1845 40433
rect 1803 40384 1804 40424
rect 1844 40384 1845 40424
rect 1803 40375 1845 40384
rect 1708 39920 1748 39929
rect 1612 39880 1708 39920
rect 1708 39871 1748 39880
rect 1516 39796 1652 39836
rect 1516 39668 1556 39679
rect 1516 39593 1556 39628
rect 1515 39584 1557 39593
rect 1515 39544 1516 39584
rect 1556 39544 1557 39584
rect 1515 39535 1557 39544
rect 1515 39080 1557 39089
rect 1515 39040 1516 39080
rect 1556 39040 1557 39080
rect 1515 39031 1557 39040
rect 1516 38946 1556 39031
rect 1612 38501 1652 39796
rect 1708 38912 1748 38921
rect 1708 38753 1748 38872
rect 1707 38744 1749 38753
rect 1707 38704 1708 38744
rect 1748 38704 1749 38744
rect 1707 38695 1749 38704
rect 1611 38492 1653 38501
rect 1611 38452 1612 38492
rect 1652 38452 1653 38492
rect 1611 38443 1653 38452
rect 1708 38417 1748 38695
rect 1707 38408 1749 38417
rect 1707 38368 1708 38408
rect 1748 38368 1749 38408
rect 1707 38359 1749 38368
rect 1804 38240 1844 40375
rect 1900 40349 1940 41131
rect 1899 40340 1941 40349
rect 1899 40300 1900 40340
rect 1940 40300 1941 40340
rect 1899 40291 1941 40300
rect 1900 40206 1940 40291
rect 1996 39920 2036 42928
rect 2092 41432 2132 41443
rect 2092 41357 2132 41392
rect 2091 41348 2133 41357
rect 2091 41308 2092 41348
rect 2132 41308 2133 41348
rect 2091 41299 2133 41308
rect 2091 40844 2133 40853
rect 2091 40804 2092 40844
rect 2132 40804 2133 40844
rect 2091 40795 2133 40804
rect 1708 38200 1844 38240
rect 1900 39880 2036 39920
rect 1420 37864 1556 37904
rect 1420 37484 1460 37493
rect 1324 37444 1420 37484
rect 1131 37064 1173 37073
rect 1131 37024 1132 37064
rect 1172 37024 1173 37064
rect 1131 37015 1173 37024
rect 1132 36233 1172 37015
rect 1228 36728 1268 36737
rect 1228 36569 1268 36688
rect 1227 36560 1269 36569
rect 1227 36520 1228 36560
rect 1268 36520 1269 36560
rect 1227 36511 1269 36520
rect 1131 36224 1173 36233
rect 1131 36184 1132 36224
rect 1172 36184 1173 36224
rect 1131 36175 1173 36184
rect 1324 34301 1364 37444
rect 1420 37435 1460 37444
rect 1420 35972 1460 35981
rect 1420 35477 1460 35932
rect 1516 35552 1556 37864
rect 1611 37736 1653 37745
rect 1611 37696 1612 37736
rect 1652 37696 1653 37736
rect 1611 37687 1653 37696
rect 1612 37652 1652 37687
rect 1612 37601 1652 37612
rect 1611 36140 1653 36149
rect 1611 36100 1612 36140
rect 1652 36100 1653 36140
rect 1611 36091 1653 36100
rect 1612 36006 1652 36091
rect 1516 35512 1652 35552
rect 1419 35468 1461 35477
rect 1419 35428 1420 35468
rect 1460 35428 1461 35468
rect 1419 35419 1461 35428
rect 1419 35300 1461 35309
rect 1419 35260 1420 35300
rect 1460 35260 1461 35300
rect 1419 35251 1461 35260
rect 1420 34469 1460 35251
rect 1516 35132 1556 35141
rect 1516 34721 1556 35092
rect 1515 34712 1557 34721
rect 1515 34672 1516 34712
rect 1556 34672 1557 34712
rect 1515 34663 1557 34672
rect 1612 34628 1652 35512
rect 1708 35048 1748 38200
rect 1804 37484 1844 37493
rect 1804 37157 1844 37444
rect 1803 37148 1845 37157
rect 1803 37108 1804 37148
rect 1844 37108 1845 37148
rect 1803 37099 1845 37108
rect 1900 36140 1940 39880
rect 2092 39836 2132 40795
rect 2188 40433 2228 42928
rect 2284 41264 2324 41273
rect 2284 40685 2324 41224
rect 2283 40676 2325 40685
rect 2283 40636 2284 40676
rect 2324 40636 2325 40676
rect 2283 40627 2325 40636
rect 2283 40508 2325 40517
rect 2283 40468 2284 40508
rect 2324 40468 2325 40508
rect 2283 40459 2325 40468
rect 2187 40424 2229 40433
rect 2187 40384 2188 40424
rect 2228 40384 2229 40424
rect 2187 40375 2229 40384
rect 2284 40374 2324 40459
rect 2283 39920 2325 39929
rect 2283 39880 2284 39920
rect 2324 39880 2325 39920
rect 2283 39871 2325 39880
rect 1996 39796 2132 39836
rect 1996 39752 2036 39796
rect 1996 39703 2036 39712
rect 2092 39733 2132 39742
rect 2092 39584 2132 39693
rect 1996 39544 2132 39584
rect 1996 39173 2036 39544
rect 2091 39416 2133 39425
rect 2091 39376 2092 39416
rect 2132 39376 2133 39416
rect 2091 39367 2133 39376
rect 1995 39164 2037 39173
rect 1995 39124 1996 39164
rect 2036 39124 2037 39164
rect 1995 39115 2037 39124
rect 1995 38996 2037 39005
rect 1995 38956 1996 38996
rect 2036 38956 2037 38996
rect 1995 38947 2037 38956
rect 1996 37820 2036 38947
rect 2092 38333 2132 39367
rect 2187 38576 2229 38585
rect 2187 38536 2188 38576
rect 2228 38536 2229 38576
rect 2187 38527 2229 38536
rect 2091 38324 2133 38333
rect 2091 38284 2092 38324
rect 2132 38284 2133 38324
rect 2091 38275 2133 38284
rect 1996 37780 2132 37820
rect 1995 37652 2037 37661
rect 1995 37612 1996 37652
rect 2036 37612 2037 37652
rect 1995 37603 2037 37612
rect 1996 37518 2036 37603
rect 1995 37064 2037 37073
rect 1995 37024 1996 37064
rect 2036 37024 2037 37064
rect 1995 37015 2037 37024
rect 1708 34999 1748 35008
rect 1804 36100 1940 36140
rect 1708 34628 1748 34637
rect 1612 34588 1708 34628
rect 1804 34628 1844 36100
rect 1996 36056 2036 37015
rect 2092 36569 2132 37780
rect 2091 36560 2133 36569
rect 2091 36520 2092 36560
rect 2132 36520 2133 36560
rect 2091 36511 2133 36520
rect 2091 36308 2133 36317
rect 2091 36268 2092 36308
rect 2132 36268 2133 36308
rect 2091 36259 2133 36268
rect 1900 36016 2036 36056
rect 1900 35888 1940 36016
rect 1900 35839 1940 35848
rect 1995 35888 2037 35897
rect 1995 35848 1996 35888
rect 2036 35848 2037 35888
rect 1995 35839 2037 35848
rect 1996 35754 2036 35839
rect 1899 35636 1941 35645
rect 1899 35596 1900 35636
rect 1940 35596 1941 35636
rect 1899 35587 1941 35596
rect 1900 35309 1940 35587
rect 2092 35561 2132 36259
rect 2188 36149 2228 38527
rect 2284 37400 2324 39871
rect 2380 38744 2420 42928
rect 2572 41861 2612 42928
rect 2571 41852 2613 41861
rect 2571 41812 2572 41852
rect 2612 41812 2613 41852
rect 2571 41803 2613 41812
rect 2667 41684 2709 41693
rect 2667 41644 2668 41684
rect 2708 41644 2709 41684
rect 2667 41635 2709 41644
rect 2572 39677 2612 39762
rect 2476 39668 2516 39677
rect 2476 39257 2516 39628
rect 2571 39668 2613 39677
rect 2571 39628 2572 39668
rect 2612 39628 2613 39668
rect 2571 39619 2613 39628
rect 2571 39416 2613 39425
rect 2571 39376 2572 39416
rect 2612 39376 2613 39416
rect 2571 39367 2613 39376
rect 2475 39248 2517 39257
rect 2475 39208 2476 39248
rect 2516 39208 2517 39248
rect 2475 39199 2517 39208
rect 2380 38704 2516 38744
rect 2476 38585 2516 38704
rect 2475 38576 2517 38585
rect 2475 38536 2476 38576
rect 2516 38536 2517 38576
rect 2475 38527 2517 38536
rect 2476 38249 2516 38334
rect 2475 38240 2517 38249
rect 2380 38200 2476 38240
rect 2516 38200 2517 38240
rect 2380 37568 2420 38200
rect 2475 38191 2517 38200
rect 2572 38072 2612 39367
rect 2668 38165 2708 41635
rect 2764 38240 2804 42928
rect 2859 40676 2901 40685
rect 2859 40636 2860 40676
rect 2900 40636 2901 40676
rect 2859 40627 2901 40636
rect 2860 40519 2900 40627
rect 2860 40470 2900 40479
rect 2956 40340 2996 42928
rect 3051 42440 3093 42449
rect 3051 42400 3052 42440
rect 3092 42400 3093 42440
rect 3051 42391 3093 42400
rect 3052 40676 3092 42391
rect 3148 41693 3188 42928
rect 3147 41684 3189 41693
rect 3147 41644 3148 41684
rect 3188 41644 3189 41684
rect 3147 41635 3189 41644
rect 3340 41516 3380 42928
rect 3435 42188 3477 42197
rect 3435 42148 3436 42188
rect 3476 42148 3477 42188
rect 3435 42139 3477 42148
rect 3052 40627 3092 40636
rect 3148 41476 3380 41516
rect 2860 40300 2996 40340
rect 2860 39425 2900 40300
rect 2955 39836 2997 39845
rect 2955 39796 2956 39836
rect 2996 39796 2997 39836
rect 2955 39787 2997 39796
rect 2859 39416 2901 39425
rect 2859 39376 2860 39416
rect 2900 39376 2901 39416
rect 2859 39367 2901 39376
rect 2956 39248 2996 39787
rect 3051 39752 3093 39761
rect 3051 39712 3052 39752
rect 3092 39712 3093 39752
rect 3051 39703 3093 39712
rect 3052 39618 3092 39703
rect 2860 39208 2996 39248
rect 2860 38417 2900 39208
rect 2955 38912 2997 38921
rect 3148 38912 3188 41476
rect 3339 41180 3381 41189
rect 3339 41140 3340 41180
rect 3380 41140 3381 41180
rect 3339 41131 3381 41140
rect 3244 40508 3284 40517
rect 3244 40349 3284 40468
rect 3243 40340 3285 40349
rect 3243 40300 3244 40340
rect 3284 40300 3285 40340
rect 3243 40291 3285 40300
rect 3340 39584 3380 41131
rect 3436 40676 3476 42139
rect 3532 41516 3572 42928
rect 3724 42533 3764 42928
rect 3723 42524 3765 42533
rect 3723 42484 3724 42524
rect 3764 42484 3765 42524
rect 3723 42475 3765 42484
rect 3532 41476 3668 41516
rect 3436 40627 3476 40636
rect 3532 41264 3572 41273
rect 3532 40433 3572 41224
rect 3628 41189 3668 41476
rect 3916 41264 3956 42928
rect 4108 41936 4148 42928
rect 4300 42281 4340 42928
rect 4492 42365 4532 42928
rect 4491 42356 4533 42365
rect 4491 42316 4492 42356
rect 4532 42316 4533 42356
rect 4491 42307 4533 42316
rect 4299 42272 4341 42281
rect 4299 42232 4300 42272
rect 4340 42232 4341 42272
rect 4299 42223 4341 42232
rect 4108 41896 4436 41936
rect 4203 41768 4245 41777
rect 4203 41728 4204 41768
rect 4244 41728 4245 41768
rect 4203 41719 4245 41728
rect 4107 41516 4149 41525
rect 4107 41476 4108 41516
rect 4148 41476 4149 41516
rect 4107 41467 4149 41476
rect 4108 41264 4148 41467
rect 3916 41224 4052 41264
rect 3627 41180 3669 41189
rect 3627 41140 3628 41180
rect 3668 41140 3669 41180
rect 3627 41131 3669 41140
rect 3724 41105 3764 41190
rect 3723 41096 3765 41105
rect 3723 41056 3724 41096
rect 3764 41056 3765 41096
rect 3723 41047 3765 41056
rect 3916 41021 3956 41106
rect 4012 41096 4052 41224
rect 4108 41215 4148 41224
rect 4012 41056 4148 41096
rect 3915 41012 3957 41021
rect 3915 40972 3916 41012
rect 3956 40972 3957 41012
rect 3915 40963 3957 40972
rect 3688 40844 4056 40853
rect 3728 40804 3770 40844
rect 3810 40804 3852 40844
rect 3892 40804 3934 40844
rect 3974 40804 4016 40844
rect 3688 40795 4056 40804
rect 3531 40424 3573 40433
rect 3531 40384 3532 40424
rect 3572 40384 3573 40424
rect 3531 40375 3573 40384
rect 3819 40424 3861 40433
rect 3819 40384 3820 40424
rect 3860 40384 3861 40424
rect 3819 40375 3861 40384
rect 3820 40290 3860 40375
rect 3628 40256 3668 40265
rect 3628 39752 3668 40216
rect 3580 39742 3668 39752
rect 3620 39712 3668 39742
rect 3724 39836 3764 39845
rect 3580 39693 3620 39702
rect 3340 39544 3572 39584
rect 3435 39416 3477 39425
rect 3435 39376 3436 39416
rect 3476 39376 3477 39416
rect 3435 39367 3477 39376
rect 3340 38912 3380 38921
rect 2955 38872 2956 38912
rect 2996 38872 2997 38912
rect 2955 38863 2997 38872
rect 3052 38872 3188 38912
rect 3244 38872 3340 38912
rect 2956 38778 2996 38863
rect 2859 38408 2901 38417
rect 2859 38368 2860 38408
rect 2900 38368 2901 38408
rect 3052 38408 3092 38872
rect 3147 38744 3189 38753
rect 3147 38704 3148 38744
rect 3188 38704 3189 38744
rect 3147 38695 3189 38704
rect 3148 38610 3188 38695
rect 3148 38408 3188 38417
rect 3052 38368 3148 38408
rect 2859 38359 2901 38368
rect 3148 38359 3188 38368
rect 2764 38200 2900 38240
rect 2667 38156 2709 38165
rect 2667 38116 2668 38156
rect 2708 38116 2709 38156
rect 2667 38107 2709 38116
rect 2476 38032 2612 38072
rect 2476 37745 2516 38032
rect 2668 37988 2708 37997
rect 2668 37820 2708 37948
rect 2572 37780 2708 37820
rect 2763 37820 2805 37829
rect 2763 37780 2764 37820
rect 2804 37780 2805 37820
rect 2860 37820 2900 38200
rect 2955 38156 2997 38165
rect 2955 38116 2956 38156
rect 2996 38116 2997 38156
rect 2955 38107 2997 38116
rect 2956 38022 2996 38107
rect 3244 37988 3284 38872
rect 3340 38863 3380 38872
rect 3340 38156 3380 38165
rect 3436 38156 3476 39367
rect 3532 38408 3572 39544
rect 3724 39509 3764 39796
rect 4012 39752 4052 39763
rect 4012 39677 4052 39712
rect 4011 39668 4053 39677
rect 4011 39628 4012 39668
rect 4052 39628 4053 39668
rect 4011 39619 4053 39628
rect 3723 39500 3765 39509
rect 3723 39460 3724 39500
rect 3764 39460 3765 39500
rect 3723 39451 3765 39460
rect 3688 39332 4056 39341
rect 3728 39292 3770 39332
rect 3810 39292 3852 39332
rect 3892 39292 3934 39332
rect 3974 39292 4016 39332
rect 3688 39283 4056 39292
rect 4108 39173 4148 41056
rect 4107 39164 4149 39173
rect 4107 39124 4108 39164
rect 4148 39124 4149 39164
rect 4107 39115 4149 39124
rect 3627 39080 3669 39089
rect 3627 39040 3628 39080
rect 3668 39040 3669 39080
rect 3627 39031 3669 39040
rect 3628 38753 3668 39031
rect 3627 38744 3669 38753
rect 3627 38704 3628 38744
rect 3668 38704 3669 38744
rect 3627 38695 3669 38704
rect 3532 38359 3572 38368
rect 3627 38408 3669 38417
rect 3627 38368 3628 38408
rect 3668 38368 3669 38408
rect 3627 38359 3669 38368
rect 4012 38408 4052 38417
rect 4204 38408 4244 41719
rect 4299 39668 4341 39677
rect 4299 39628 4300 39668
rect 4340 39628 4341 39668
rect 4299 39619 4341 39628
rect 4052 38368 4244 38408
rect 4012 38359 4052 38368
rect 3380 38116 3476 38156
rect 3340 38107 3380 38116
rect 3628 37997 3668 38359
rect 3820 38156 3860 38165
rect 3820 37997 3860 38116
rect 4107 38156 4149 38165
rect 4107 38116 4108 38156
rect 4148 38116 4149 38156
rect 4107 38107 4149 38116
rect 3627 37988 3669 37997
rect 3244 37948 3572 37988
rect 3243 37820 3285 37829
rect 2860 37780 2996 37820
rect 2475 37736 2517 37745
rect 2475 37696 2476 37736
rect 2516 37696 2517 37736
rect 2475 37687 2517 37696
rect 2380 37528 2516 37568
rect 2284 37351 2324 37360
rect 2380 37400 2420 37409
rect 2380 36989 2420 37360
rect 2379 36980 2421 36989
rect 2379 36940 2380 36980
rect 2420 36940 2421 36980
rect 2379 36931 2421 36940
rect 2476 36728 2516 37528
rect 2476 36317 2516 36688
rect 2475 36308 2517 36317
rect 2475 36268 2476 36308
rect 2516 36268 2517 36308
rect 2475 36259 2517 36268
rect 2187 36140 2229 36149
rect 2187 36100 2188 36140
rect 2228 36100 2229 36140
rect 2187 36091 2229 36100
rect 2380 35888 2420 35897
rect 2284 35848 2380 35888
rect 2091 35552 2133 35561
rect 2091 35512 2092 35552
rect 2132 35512 2133 35552
rect 2091 35503 2133 35512
rect 1899 35300 1941 35309
rect 1899 35260 1900 35300
rect 1940 35260 1941 35300
rect 1899 35251 1941 35260
rect 2092 35216 2132 35503
rect 2092 35167 2132 35176
rect 1900 34964 1940 34973
rect 1940 34924 2036 34964
rect 1900 34915 1940 34924
rect 1900 34628 1940 34637
rect 1804 34588 1900 34628
rect 1708 34579 1748 34588
rect 1900 34579 1940 34588
rect 1419 34460 1461 34469
rect 1419 34420 1420 34460
rect 1460 34420 1461 34460
rect 1419 34411 1461 34420
rect 1516 34460 1556 34469
rect 1323 34292 1365 34301
rect 1323 34252 1324 34292
rect 1364 34252 1365 34292
rect 1323 34243 1365 34252
rect 1228 33704 1268 33713
rect 1268 33664 1460 33704
rect 1228 33655 1268 33664
rect 939 33032 981 33041
rect 939 32992 940 33032
rect 980 32992 981 33032
rect 939 32983 981 32992
rect 171 31856 213 31865
rect 171 31816 172 31856
rect 212 31816 213 31856
rect 171 31807 213 31816
rect 172 23960 212 31807
rect 76 23920 212 23960
rect 76 23633 116 23920
rect 75 23624 117 23633
rect 75 23584 76 23624
rect 116 23584 117 23624
rect 75 23575 117 23584
rect 940 21617 980 32983
rect 1420 32369 1460 33664
rect 1419 32360 1461 32369
rect 1419 32320 1420 32360
rect 1460 32320 1461 32360
rect 1419 32311 1461 32320
rect 1035 32108 1077 32117
rect 1035 32068 1036 32108
rect 1076 32068 1077 32108
rect 1035 32059 1077 32068
rect 1036 26321 1076 32059
rect 1323 31520 1365 31529
rect 1323 31480 1324 31520
rect 1364 31480 1365 31520
rect 1323 31471 1365 31480
rect 1324 30353 1364 31471
rect 1323 30344 1365 30353
rect 1323 30304 1324 30344
rect 1364 30304 1365 30344
rect 1323 30295 1365 30304
rect 1323 29840 1365 29849
rect 1323 29800 1324 29840
rect 1364 29800 1365 29840
rect 1323 29791 1365 29800
rect 1324 29706 1364 29791
rect 1420 28496 1460 32311
rect 1516 28505 1556 34420
rect 1611 34460 1653 34469
rect 1611 34420 1612 34460
rect 1652 34420 1653 34460
rect 1611 34411 1653 34420
rect 1899 34460 1941 34469
rect 1899 34420 1900 34460
rect 1940 34420 1941 34460
rect 1899 34411 1941 34420
rect 1612 31529 1652 34411
rect 1803 34292 1845 34301
rect 1803 34252 1804 34292
rect 1844 34252 1845 34292
rect 1803 34243 1845 34252
rect 1804 32780 1844 34243
rect 1900 33377 1940 34411
rect 1899 33368 1941 33377
rect 1899 33328 1900 33368
rect 1940 33328 1941 33368
rect 1899 33319 1941 33328
rect 1996 32864 2036 34924
rect 2092 34460 2132 34469
rect 2092 33032 2132 34420
rect 2284 33209 2324 35848
rect 2380 35839 2420 35848
rect 2476 35888 2516 35897
rect 2476 35645 2516 35848
rect 2475 35636 2517 35645
rect 2475 35596 2476 35636
rect 2516 35596 2517 35636
rect 2475 35587 2517 35596
rect 2572 35300 2612 37780
rect 2763 37771 2805 37780
rect 2764 37661 2804 37771
rect 2763 37652 2805 37661
rect 2763 37612 2764 37652
rect 2804 37612 2805 37652
rect 2763 37603 2805 37612
rect 2764 37400 2804 37409
rect 2764 36653 2804 37360
rect 2860 37400 2900 37409
rect 2763 36644 2805 36653
rect 2763 36604 2764 36644
rect 2804 36604 2805 36644
rect 2763 36595 2805 36604
rect 2668 36476 2708 36485
rect 2708 36436 2804 36476
rect 2668 36427 2708 36436
rect 2380 35260 2612 35300
rect 2380 34376 2420 35260
rect 2380 34327 2420 34336
rect 2476 34376 2516 34385
rect 2476 33872 2516 34336
rect 2380 33832 2516 33872
rect 2283 33200 2325 33209
rect 2283 33160 2284 33200
rect 2324 33160 2325 33200
rect 2283 33151 2325 33160
rect 2092 32992 2324 33032
rect 2140 32873 2180 32882
rect 1996 32833 2140 32864
rect 1996 32824 2180 32833
rect 1804 32740 2036 32780
rect 1996 32696 2036 32740
rect 1996 32647 2036 32656
rect 2091 32696 2133 32705
rect 2091 32656 2092 32696
rect 2132 32656 2133 32696
rect 2091 32647 2133 32656
rect 1803 32192 1845 32201
rect 1803 32152 1804 32192
rect 1844 32152 1845 32192
rect 1803 32143 1845 32152
rect 2092 32192 2132 32647
rect 2284 32369 2324 32992
rect 2283 32360 2325 32369
rect 2283 32320 2284 32360
rect 2324 32320 2325 32360
rect 2283 32311 2325 32320
rect 2380 32201 2420 33832
rect 2475 33704 2517 33713
rect 2475 33664 2476 33704
rect 2516 33664 2517 33704
rect 2475 33655 2517 33664
rect 2476 33570 2516 33655
rect 2668 33452 2708 33461
rect 2572 33412 2668 33452
rect 2475 33368 2517 33377
rect 2475 33328 2476 33368
rect 2516 33328 2517 33368
rect 2475 33319 2517 33328
rect 1611 31520 1653 31529
rect 1611 31480 1612 31520
rect 1652 31480 1653 31520
rect 1611 31471 1653 31480
rect 1707 30680 1749 30689
rect 1707 30640 1708 30680
rect 1748 30640 1749 30680
rect 1707 30631 1749 30640
rect 1611 30596 1653 30605
rect 1611 30556 1612 30596
rect 1652 30556 1653 30596
rect 1611 30547 1653 30556
rect 1324 28456 1460 28496
rect 1515 28496 1557 28505
rect 1515 28456 1516 28496
rect 1556 28456 1557 28496
rect 1227 27068 1269 27077
rect 1227 27028 1228 27068
rect 1268 27028 1269 27068
rect 1227 27019 1269 27028
rect 1228 26816 1268 27019
rect 1324 26909 1364 28456
rect 1515 28447 1557 28456
rect 1420 28328 1460 28337
rect 1420 27917 1460 28288
rect 1516 28328 1556 28339
rect 1612 28337 1652 30547
rect 1708 28421 1748 30631
rect 1707 28412 1749 28421
rect 1707 28372 1708 28412
rect 1748 28372 1749 28412
rect 1707 28363 1749 28372
rect 1516 28253 1556 28288
rect 1611 28328 1653 28337
rect 1611 28288 1612 28328
rect 1652 28288 1653 28328
rect 1611 28279 1653 28288
rect 1515 28244 1557 28253
rect 1515 28204 1516 28244
rect 1556 28204 1557 28244
rect 1515 28195 1557 28204
rect 1419 27908 1461 27917
rect 1419 27868 1420 27908
rect 1460 27868 1461 27908
rect 1419 27859 1461 27868
rect 1612 27833 1652 28279
rect 1611 27824 1653 27833
rect 1611 27784 1612 27824
rect 1652 27784 1653 27824
rect 1611 27775 1653 27784
rect 1707 27656 1749 27665
rect 1707 27616 1708 27656
rect 1748 27616 1749 27656
rect 1707 27607 1749 27616
rect 1419 27572 1461 27581
rect 1419 27532 1420 27572
rect 1460 27532 1461 27572
rect 1419 27523 1461 27532
rect 1323 26900 1365 26909
rect 1323 26860 1324 26900
rect 1364 26860 1365 26900
rect 1323 26851 1365 26860
rect 1228 26767 1268 26776
rect 1035 26312 1077 26321
rect 1035 26272 1036 26312
rect 1076 26272 1077 26312
rect 1035 26263 1077 26272
rect 1035 25640 1077 25649
rect 1035 25600 1036 25640
rect 1076 25600 1077 25640
rect 1035 25591 1077 25600
rect 939 21608 981 21617
rect 939 21568 940 21608
rect 980 21568 981 21608
rect 939 21559 981 21568
rect 1036 18929 1076 25591
rect 1228 23792 1268 23801
rect 1323 23792 1365 23801
rect 1268 23752 1324 23792
rect 1364 23752 1365 23792
rect 1228 23743 1268 23752
rect 1323 23743 1365 23752
rect 1228 23120 1268 23129
rect 1268 23080 1364 23120
rect 1228 23071 1268 23080
rect 1131 22952 1173 22961
rect 1131 22912 1132 22952
rect 1172 22912 1173 22952
rect 1131 22903 1173 22912
rect 1132 20861 1172 22903
rect 1227 21608 1269 21617
rect 1227 21568 1228 21608
rect 1268 21568 1269 21608
rect 1227 21559 1269 21568
rect 1228 21029 1268 21559
rect 1227 21020 1269 21029
rect 1227 20980 1228 21020
rect 1268 20980 1269 21020
rect 1227 20971 1269 20980
rect 1131 20852 1173 20861
rect 1131 20812 1132 20852
rect 1172 20812 1173 20852
rect 1131 20803 1173 20812
rect 1227 20768 1269 20777
rect 1227 20728 1228 20768
rect 1268 20728 1269 20768
rect 1227 20719 1269 20728
rect 1228 20634 1268 20719
rect 1131 20180 1173 20189
rect 1131 20140 1132 20180
rect 1172 20140 1173 20180
rect 1131 20131 1173 20140
rect 1132 19601 1172 20131
rect 1228 20096 1268 20105
rect 1324 20096 1364 23080
rect 1268 20056 1364 20096
rect 1228 19685 1268 20056
rect 1227 19676 1269 19685
rect 1227 19636 1228 19676
rect 1268 19636 1269 19676
rect 1227 19627 1269 19636
rect 1131 19592 1173 19601
rect 1131 19552 1132 19592
rect 1172 19552 1173 19592
rect 1131 19543 1173 19552
rect 1035 18920 1077 18929
rect 1035 18880 1036 18920
rect 1076 18880 1077 18920
rect 1035 18871 1077 18880
rect 1323 18248 1365 18257
rect 1323 18208 1324 18248
rect 1364 18208 1365 18248
rect 1323 18199 1365 18208
rect 1228 17744 1268 17753
rect 1324 17744 1364 18199
rect 1268 17704 1364 17744
rect 1228 17695 1268 17704
rect 1323 17072 1365 17081
rect 1323 17032 1324 17072
rect 1364 17032 1365 17072
rect 1323 17023 1365 17032
rect 1324 16938 1364 17023
rect 1228 15560 1268 15569
rect 1420 15560 1460 27523
rect 1708 27522 1748 27607
rect 1804 26480 1844 32143
rect 2092 31268 2132 32152
rect 2379 32192 2421 32201
rect 2379 32152 2380 32192
rect 2420 32152 2421 32192
rect 2379 32143 2421 32152
rect 2476 31856 2516 33319
rect 2380 31816 2516 31856
rect 2380 31772 2420 31816
rect 1996 31228 2132 31268
rect 2188 31732 2420 31772
rect 1996 28832 2036 31228
rect 2092 29168 2132 29177
rect 2188 29168 2228 31732
rect 2572 31688 2612 33412
rect 2668 33403 2708 33412
rect 2667 33200 2709 33209
rect 2667 33160 2668 33200
rect 2708 33160 2709 33200
rect 2667 33151 2709 33160
rect 2668 32864 2708 33151
rect 2764 32873 2804 36436
rect 2860 34553 2900 37360
rect 2956 36056 2996 37780
rect 3243 37780 3244 37820
rect 3284 37780 3285 37820
rect 3243 37771 3285 37780
rect 3435 37820 3477 37829
rect 3435 37780 3436 37820
rect 3476 37780 3477 37820
rect 3435 37771 3477 37780
rect 3051 36728 3093 36737
rect 3051 36688 3052 36728
rect 3092 36688 3093 36728
rect 3051 36686 3093 36688
rect 3051 36679 3052 36686
rect 3092 36679 3093 36686
rect 3052 36140 3092 36646
rect 3052 36100 3188 36140
rect 2956 36016 3092 36056
rect 2956 35888 2996 35897
rect 2956 35225 2996 35848
rect 2955 35216 2997 35225
rect 2955 35176 2956 35216
rect 2996 35176 2997 35216
rect 2955 35167 2997 35176
rect 3052 35057 3092 36016
rect 3148 35729 3188 36100
rect 3147 35720 3189 35729
rect 3147 35680 3148 35720
rect 3188 35680 3189 35720
rect 3147 35671 3189 35680
rect 3147 35300 3189 35309
rect 3147 35260 3148 35300
rect 3188 35260 3189 35300
rect 3244 35300 3284 37771
rect 3339 37400 3381 37409
rect 3339 37360 3340 37400
rect 3380 37360 3381 37400
rect 3339 37351 3381 37360
rect 3340 37266 3380 37351
rect 3436 35902 3476 37771
rect 3532 37745 3572 37948
rect 3627 37948 3628 37988
rect 3668 37948 3669 37988
rect 3627 37939 3669 37948
rect 3819 37988 3861 37997
rect 3819 37948 3820 37988
rect 3860 37948 3861 37988
rect 3819 37939 3861 37948
rect 3688 37820 4056 37829
rect 3728 37780 3770 37820
rect 3810 37780 3852 37820
rect 3892 37780 3934 37820
rect 3974 37780 4016 37820
rect 3688 37771 4056 37780
rect 3531 37736 3573 37745
rect 3531 37696 3532 37736
rect 3572 37696 3573 37736
rect 3531 37687 3573 37696
rect 3436 35853 3476 35862
rect 3435 35300 3477 35309
rect 3532 35300 3572 37687
rect 3819 37652 3861 37661
rect 3819 37612 3820 37652
rect 3860 37612 3861 37652
rect 3819 37603 3861 37612
rect 3820 37414 3860 37603
rect 3820 37365 3860 37374
rect 4012 37316 4052 37325
rect 4108 37316 4148 38107
rect 4300 38081 4340 39619
rect 4396 38921 4436 41896
rect 4684 41693 4724 42928
rect 4876 42113 4916 42928
rect 4875 42104 4917 42113
rect 4875 42064 4876 42104
rect 4916 42064 4917 42104
rect 4875 42055 4917 42064
rect 5068 41768 5108 42928
rect 5260 41777 5300 42928
rect 5355 42020 5397 42029
rect 5355 41980 5356 42020
rect 5396 41980 5397 42020
rect 5355 41971 5397 41980
rect 4780 41728 5108 41768
rect 5259 41768 5301 41777
rect 5259 41728 5260 41768
rect 5300 41728 5301 41768
rect 4683 41684 4725 41693
rect 4683 41644 4684 41684
rect 4724 41644 4725 41684
rect 4683 41635 4725 41644
rect 4587 41600 4629 41609
rect 4587 41560 4588 41600
rect 4628 41560 4629 41600
rect 4587 41551 4629 41560
rect 4491 41516 4533 41525
rect 4491 41476 4492 41516
rect 4532 41476 4533 41516
rect 4491 41467 4533 41476
rect 4492 40433 4532 41467
rect 4588 41180 4628 41551
rect 4780 41357 4820 41728
rect 5259 41719 5301 41728
rect 4928 41600 5296 41609
rect 4968 41560 5010 41600
rect 5050 41560 5092 41600
rect 5132 41560 5174 41600
rect 5214 41560 5256 41600
rect 4928 41551 5296 41560
rect 4779 41348 4821 41357
rect 4779 41308 4780 41348
rect 4820 41308 4821 41348
rect 4779 41299 4821 41308
rect 5356 41264 5396 41971
rect 4588 41140 5108 41180
rect 4491 40424 4533 40433
rect 4491 40384 4492 40424
rect 4532 40384 4533 40424
rect 4491 40375 4533 40384
rect 5068 40424 5108 41140
rect 5356 41021 5396 41224
rect 5355 41012 5397 41021
rect 5355 40972 5356 41012
rect 5396 40972 5397 41012
rect 5355 40963 5397 40972
rect 5452 40844 5492 42928
rect 5644 42449 5684 42928
rect 5643 42440 5685 42449
rect 5643 42400 5644 42440
rect 5684 42400 5685 42440
rect 5643 42391 5685 42400
rect 5836 42104 5876 42928
rect 6028 42197 6068 42928
rect 6027 42188 6069 42197
rect 6027 42148 6028 42188
rect 6068 42148 6069 42188
rect 6027 42139 6069 42148
rect 5644 42064 5876 42104
rect 5547 41180 5589 41189
rect 5547 41140 5548 41180
rect 5588 41140 5589 41180
rect 5547 41131 5589 41140
rect 5548 41046 5588 41131
rect 5356 40804 5492 40844
rect 4395 38912 4437 38921
rect 4395 38872 4396 38912
rect 4436 38872 4437 38912
rect 4395 38863 4437 38872
rect 4395 38240 4437 38249
rect 4492 38240 4532 40375
rect 5068 40265 5108 40384
rect 5260 40508 5300 40517
rect 5260 40349 5300 40468
rect 5259 40340 5301 40349
rect 5259 40300 5260 40340
rect 5300 40300 5301 40340
rect 5259 40291 5301 40300
rect 5067 40256 5109 40265
rect 5067 40216 5068 40256
rect 5108 40216 5109 40256
rect 5067 40207 5109 40216
rect 4928 40088 5296 40097
rect 4968 40048 5010 40088
rect 5050 40048 5092 40088
rect 5132 40048 5174 40088
rect 5214 40048 5256 40088
rect 4928 40039 5296 40048
rect 5260 39752 5300 39761
rect 5260 39593 5300 39712
rect 4587 39584 4629 39593
rect 4587 39544 4588 39584
rect 4628 39544 4629 39584
rect 4587 39535 4629 39544
rect 5259 39584 5301 39593
rect 5259 39544 5260 39584
rect 5300 39544 5301 39584
rect 5259 39535 5301 39544
rect 4588 38912 4628 39535
rect 5356 39080 5396 40804
rect 5451 40676 5493 40685
rect 5644 40676 5684 42064
rect 6220 42020 6260 42928
rect 5740 41980 6260 42020
rect 5740 41432 5780 41980
rect 6412 41600 6452 42928
rect 6220 41560 6452 41600
rect 6507 41600 6549 41609
rect 6507 41560 6508 41600
rect 6548 41560 6549 41600
rect 6123 41516 6165 41525
rect 6123 41476 6124 41516
rect 6164 41476 6165 41516
rect 6123 41467 6165 41476
rect 5740 41383 5780 41392
rect 6124 41432 6164 41467
rect 6124 41381 6164 41392
rect 5835 41180 5877 41189
rect 5835 41140 5836 41180
rect 5876 41140 5877 41180
rect 5835 41131 5877 41140
rect 5932 41180 5972 41189
rect 5451 40636 5452 40676
rect 5492 40636 5493 40676
rect 5451 40627 5493 40636
rect 5548 40636 5684 40676
rect 5836 40676 5876 41131
rect 5452 40542 5492 40627
rect 5451 39500 5493 39509
rect 5451 39460 5452 39500
rect 5492 39460 5493 39500
rect 5451 39451 5493 39460
rect 5452 39366 5492 39451
rect 5548 39248 5588 40636
rect 5836 40627 5876 40636
rect 5644 40508 5684 40517
rect 5684 40468 5780 40508
rect 5644 40459 5684 40468
rect 5643 40340 5685 40349
rect 5643 40300 5644 40340
rect 5684 40300 5685 40340
rect 5643 40291 5685 40300
rect 5644 39593 5684 40291
rect 5643 39584 5685 39593
rect 5643 39544 5644 39584
rect 5684 39544 5685 39584
rect 5643 39535 5685 39544
rect 5643 39416 5685 39425
rect 5643 39376 5644 39416
rect 5684 39376 5685 39416
rect 5643 39367 5685 39376
rect 5356 39031 5396 39040
rect 5452 39208 5588 39248
rect 4971 38996 5013 39005
rect 4971 38956 4972 38996
rect 5012 38956 5013 38996
rect 4971 38947 5013 38956
rect 4588 38837 4628 38872
rect 4972 38862 5012 38947
rect 4587 38828 4629 38837
rect 4587 38788 4588 38828
rect 4628 38788 4629 38828
rect 4587 38779 4629 38788
rect 4395 38200 4396 38240
rect 4436 38200 4532 38240
rect 4395 38191 4437 38200
rect 4396 38106 4436 38191
rect 4299 38072 4341 38081
rect 4299 38032 4300 38072
rect 4340 38032 4341 38072
rect 4299 38023 4341 38032
rect 4491 38072 4533 38081
rect 4491 38032 4492 38072
rect 4532 38032 4533 38072
rect 4491 38023 4533 38032
rect 4052 37276 4148 37316
rect 4204 37988 4244 37997
rect 4012 37267 4052 37276
rect 4107 37148 4149 37157
rect 4107 37108 4108 37148
rect 4148 37108 4149 37148
rect 4107 37099 4149 37108
rect 3688 36308 4056 36317
rect 3728 36268 3770 36308
rect 3810 36268 3852 36308
rect 3892 36268 3934 36308
rect 3974 36268 4016 36308
rect 3688 36259 4056 36268
rect 3628 35720 3668 35729
rect 3628 35309 3668 35680
rect 4011 35720 4053 35729
rect 4011 35680 4012 35720
rect 4052 35680 4053 35720
rect 4011 35671 4053 35680
rect 4012 35586 4052 35671
rect 3244 35260 3380 35300
rect 3147 35251 3189 35260
rect 3051 35048 3093 35057
rect 3051 35008 3052 35048
rect 3092 35008 3093 35048
rect 3051 34999 3093 35008
rect 2859 34544 2901 34553
rect 2859 34504 2860 34544
rect 2900 34504 2901 34544
rect 2859 34495 2901 34504
rect 2860 34376 2900 34385
rect 2668 32815 2708 32824
rect 2763 32864 2805 32873
rect 2763 32824 2764 32864
rect 2804 32824 2805 32864
rect 2763 32815 2805 32824
rect 2284 31648 2612 31688
rect 2284 30680 2324 31648
rect 2379 31520 2421 31529
rect 2379 31480 2380 31520
rect 2420 31480 2421 31520
rect 2379 31471 2421 31480
rect 2284 30631 2324 30640
rect 2380 30680 2420 31471
rect 2667 31352 2709 31361
rect 2572 31312 2668 31352
rect 2708 31312 2709 31352
rect 2475 31268 2517 31277
rect 2475 31228 2476 31268
rect 2516 31228 2517 31268
rect 2475 31219 2517 31228
rect 2283 30260 2325 30269
rect 2283 30220 2284 30260
rect 2324 30220 2325 30260
rect 2283 30211 2325 30220
rect 2132 29128 2228 29168
rect 2092 29119 2132 29128
rect 1996 28792 2132 28832
rect 1995 28412 2037 28421
rect 1995 28372 1996 28412
rect 2036 28372 2037 28412
rect 1995 28363 2037 28372
rect 1899 28328 1941 28337
rect 1899 28288 1900 28328
rect 1940 28288 1941 28328
rect 1899 28279 1941 28288
rect 1900 28194 1940 28279
rect 1996 28278 2036 28363
rect 1899 28076 1941 28085
rect 1899 28036 1900 28076
rect 1940 28036 1941 28076
rect 1899 28027 1941 28036
rect 1708 26440 1844 26480
rect 1515 26144 1557 26153
rect 1515 26104 1516 26144
rect 1556 26104 1557 26144
rect 1515 26095 1557 26104
rect 1516 25817 1556 26095
rect 1515 25808 1557 25817
rect 1515 25768 1516 25808
rect 1556 25768 1557 25808
rect 1515 25759 1557 25768
rect 1708 23549 1748 26440
rect 1900 23960 1940 28027
rect 1995 27824 2037 27833
rect 1995 27784 1996 27824
rect 2036 27784 2037 27824
rect 1995 27775 2037 27784
rect 1804 23920 1940 23960
rect 1707 23540 1749 23549
rect 1707 23500 1708 23540
rect 1748 23500 1749 23540
rect 1707 23491 1749 23500
rect 1611 20768 1653 20777
rect 1611 20728 1612 20768
rect 1652 20728 1653 20768
rect 1611 20719 1653 20728
rect 1515 16232 1557 16241
rect 1515 16192 1516 16232
rect 1556 16192 1557 16232
rect 1515 16183 1557 16192
rect 1516 16098 1556 16183
rect 1612 15653 1652 20719
rect 1708 19013 1748 23491
rect 1804 19265 1844 23920
rect 1996 19424 2036 27775
rect 2092 25649 2132 28792
rect 2187 28580 2229 28589
rect 2187 28540 2188 28580
rect 2228 28540 2229 28580
rect 2187 28531 2229 28540
rect 2188 28085 2228 28531
rect 2187 28076 2229 28085
rect 2187 28036 2188 28076
rect 2228 28036 2229 28076
rect 2187 28027 2229 28036
rect 2284 27236 2324 30211
rect 2380 28832 2420 30640
rect 2476 29840 2516 31219
rect 2572 30101 2612 31312
rect 2667 31303 2709 31312
rect 2668 31218 2708 31303
rect 2667 31016 2709 31025
rect 2667 30976 2668 31016
rect 2708 30976 2709 31016
rect 2667 30967 2709 30976
rect 2571 30092 2613 30101
rect 2571 30052 2572 30092
rect 2612 30052 2613 30092
rect 2571 30043 2613 30052
rect 2572 29840 2612 29849
rect 2476 29800 2572 29840
rect 2380 28792 2516 28832
rect 2476 28589 2516 28792
rect 2475 28580 2517 28589
rect 2475 28540 2476 28580
rect 2516 28540 2517 28580
rect 2475 28531 2517 28540
rect 2476 28328 2516 28337
rect 2379 28244 2421 28253
rect 2379 28204 2380 28244
rect 2420 28204 2421 28244
rect 2379 28195 2421 28204
rect 2188 27196 2324 27236
rect 2091 25640 2133 25649
rect 2091 25600 2092 25640
rect 2132 25600 2133 25640
rect 2091 25591 2133 25600
rect 2188 20264 2228 27196
rect 2380 25985 2420 28195
rect 2476 26984 2516 28288
rect 2572 27749 2612 29800
rect 2571 27740 2613 27749
rect 2571 27700 2572 27740
rect 2612 27700 2613 27740
rect 2571 27691 2613 27700
rect 2668 27161 2708 30967
rect 2860 30764 2900 34336
rect 2956 34376 2996 34385
rect 2956 34133 2996 34336
rect 2955 34124 2997 34133
rect 2955 34084 2956 34124
rect 2996 34084 2997 34124
rect 2955 34075 2997 34084
rect 3148 33956 3188 35251
rect 3340 35216 3380 35260
rect 3435 35260 3436 35300
rect 3476 35260 3572 35300
rect 3627 35300 3669 35309
rect 3627 35260 3628 35300
rect 3668 35260 3669 35300
rect 3435 35251 3477 35260
rect 3627 35251 3669 35260
rect 4011 35300 4053 35309
rect 4011 35260 4012 35300
rect 4052 35260 4053 35300
rect 4011 35251 4053 35260
rect 3340 34805 3380 35176
rect 3531 35132 3573 35141
rect 3531 35092 3532 35132
rect 3572 35092 3573 35132
rect 3531 35083 3573 35092
rect 4012 35132 4052 35251
rect 4012 35083 4052 35092
rect 3435 34964 3477 34973
rect 3435 34924 3436 34964
rect 3476 34924 3477 34964
rect 3435 34915 3477 34924
rect 3339 34796 3381 34805
rect 3339 34756 3340 34796
rect 3380 34756 3381 34796
rect 3339 34747 3381 34756
rect 3243 34544 3285 34553
rect 3243 34504 3244 34544
rect 3284 34504 3285 34544
rect 3243 34495 3285 34504
rect 2956 33916 3188 33956
rect 2956 31361 2996 33916
rect 3244 33116 3284 34495
rect 3436 34376 3476 34915
rect 3436 34327 3476 34336
rect 3339 33704 3381 33713
rect 3339 33664 3340 33704
rect 3380 33664 3381 33704
rect 3339 33655 3381 33664
rect 3052 33076 3284 33116
rect 3052 32621 3092 33076
rect 3147 32948 3189 32957
rect 3147 32908 3148 32948
rect 3188 32908 3189 32948
rect 3147 32899 3189 32908
rect 3148 32814 3188 32899
rect 3244 32864 3284 32873
rect 3147 32696 3189 32705
rect 3147 32656 3148 32696
rect 3188 32656 3189 32696
rect 3147 32647 3189 32656
rect 3051 32612 3093 32621
rect 3051 32572 3052 32612
rect 3092 32572 3093 32612
rect 3051 32563 3093 32572
rect 2955 31352 2997 31361
rect 2955 31312 2956 31352
rect 2996 31312 2997 31352
rect 2955 31303 2997 31312
rect 2860 30724 2996 30764
rect 2764 30596 2804 30605
rect 2764 30269 2804 30556
rect 2859 30596 2901 30605
rect 2859 30556 2860 30596
rect 2900 30556 2901 30596
rect 2859 30547 2901 30556
rect 2860 30462 2900 30547
rect 2956 30344 2996 30724
rect 2860 30304 2996 30344
rect 2763 30260 2805 30269
rect 2763 30220 2764 30260
rect 2804 30220 2805 30260
rect 2763 30211 2805 30220
rect 2763 29672 2805 29681
rect 2763 29632 2764 29672
rect 2804 29632 2805 29672
rect 2763 29623 2805 29632
rect 2764 29538 2804 29623
rect 2860 29513 2900 30304
rect 2955 29672 2997 29681
rect 2955 29632 2956 29672
rect 2996 29632 2997 29672
rect 2955 29623 2997 29632
rect 2859 29504 2901 29513
rect 2859 29464 2860 29504
rect 2900 29464 2901 29504
rect 2859 29455 2901 29464
rect 2667 27152 2709 27161
rect 2667 27112 2668 27152
rect 2708 27112 2709 27152
rect 2667 27103 2709 27112
rect 2476 26944 2804 26984
rect 2476 26816 2516 26825
rect 2476 26153 2516 26776
rect 2668 26648 2708 26657
rect 2571 26480 2613 26489
rect 2571 26440 2572 26480
rect 2612 26440 2613 26480
rect 2571 26431 2613 26440
rect 2475 26144 2517 26153
rect 2475 26104 2476 26144
rect 2516 26104 2517 26144
rect 2475 26095 2517 26104
rect 2379 25976 2421 25985
rect 2379 25936 2380 25976
rect 2420 25936 2421 25976
rect 2379 25927 2421 25936
rect 2380 25481 2420 25927
rect 2379 25472 2421 25481
rect 2379 25432 2380 25472
rect 2420 25432 2421 25472
rect 2379 25423 2421 25432
rect 2283 25304 2325 25313
rect 2283 25264 2284 25304
rect 2324 25264 2325 25304
rect 2283 25255 2325 25264
rect 2380 25304 2420 25423
rect 2380 25255 2420 25264
rect 2284 25170 2324 25255
rect 2476 23792 2516 26095
rect 2380 23752 2476 23792
rect 2380 21608 2420 23752
rect 2476 23743 2516 23752
rect 2572 23129 2612 26431
rect 2668 25313 2708 26608
rect 2764 26312 2804 26944
rect 2860 26489 2900 29455
rect 2956 28342 2996 29623
rect 3052 29345 3092 32563
rect 3148 30185 3188 32647
rect 3147 30176 3189 30185
rect 3147 30136 3148 30176
rect 3188 30136 3189 30176
rect 3147 30127 3189 30136
rect 3244 30017 3284 32824
rect 3340 32453 3380 33655
rect 3532 32705 3572 35083
rect 3819 35048 3861 35057
rect 3819 35008 3820 35048
rect 3860 35008 3861 35048
rect 3819 34999 3861 35008
rect 3820 34914 3860 34999
rect 3688 34796 4056 34805
rect 3728 34756 3770 34796
rect 3810 34756 3852 34796
rect 3892 34756 3934 34796
rect 3974 34756 4016 34796
rect 3688 34747 4056 34756
rect 3964 34385 4004 34394
rect 4004 34345 4052 34376
rect 3964 34336 4052 34345
rect 4012 34040 4052 34336
rect 4108 34208 4148 37099
rect 4204 37073 4244 37948
rect 4395 37568 4437 37577
rect 4395 37528 4396 37568
rect 4436 37528 4437 37568
rect 4395 37519 4437 37528
rect 4396 37434 4436 37519
rect 4299 37148 4341 37157
rect 4299 37108 4300 37148
rect 4340 37108 4341 37148
rect 4299 37099 4341 37108
rect 4203 37064 4245 37073
rect 4203 37024 4204 37064
rect 4244 37024 4245 37064
rect 4203 37015 4245 37024
rect 4300 36728 4340 37099
rect 4300 36679 4340 36688
rect 4492 36644 4532 38023
rect 4588 37157 4628 38779
rect 4780 38744 4820 38753
rect 4780 37820 4820 38704
rect 5164 38744 5204 38753
rect 5452 38744 5492 39208
rect 5548 38996 5588 39005
rect 5548 38837 5588 38956
rect 5547 38828 5589 38837
rect 5547 38788 5548 38828
rect 5588 38788 5589 38828
rect 5547 38779 5589 38788
rect 5644 38753 5684 39367
rect 5740 38912 5780 40468
rect 5932 39845 5972 41140
rect 6028 40424 6068 40433
rect 6028 40013 6068 40384
rect 6027 40004 6069 40013
rect 6027 39964 6028 40004
rect 6068 39964 6069 40004
rect 6027 39955 6069 39964
rect 5931 39836 5973 39845
rect 5931 39796 5932 39836
rect 5972 39796 5973 39836
rect 5931 39787 5973 39796
rect 5931 39668 5973 39677
rect 5931 39628 5932 39668
rect 5972 39628 5973 39668
rect 5931 39619 5973 39628
rect 5932 39534 5972 39619
rect 6028 39341 6068 39955
rect 6027 39332 6069 39341
rect 6027 39292 6028 39332
rect 6068 39292 6069 39332
rect 6027 39283 6069 39292
rect 5836 39080 5876 39089
rect 5836 38996 5876 39040
rect 6220 39080 6260 41560
rect 6507 41551 6549 41560
rect 6508 41357 6548 41551
rect 6507 41348 6549 41357
rect 6507 41308 6508 41348
rect 6548 41308 6549 41348
rect 6507 41299 6549 41308
rect 6508 41264 6548 41299
rect 6508 41214 6548 41224
rect 6604 41096 6644 42928
rect 6508 41056 6644 41096
rect 6316 41012 6356 41021
rect 6316 39929 6356 40972
rect 6508 40685 6548 41056
rect 6507 40676 6549 40685
rect 6796 40676 6836 42928
rect 6988 41945 7028 42928
rect 6987 41936 7029 41945
rect 6987 41896 6988 41936
rect 7028 41896 7029 41936
rect 6987 41887 7029 41896
rect 7083 41684 7125 41693
rect 7083 41644 7084 41684
rect 7124 41644 7125 41684
rect 7083 41635 7125 41644
rect 6987 41012 7029 41021
rect 6987 40972 6988 41012
rect 7028 40972 7029 41012
rect 6987 40963 7029 40972
rect 6507 40636 6508 40676
rect 6548 40636 6549 40676
rect 6507 40627 6549 40636
rect 6604 40636 6836 40676
rect 6315 39920 6357 39929
rect 6315 39880 6316 39920
rect 6356 39880 6357 39920
rect 6315 39871 6357 39880
rect 6316 39752 6356 39761
rect 6316 39089 6356 39712
rect 6412 39752 6452 39763
rect 6412 39677 6452 39712
rect 6411 39668 6453 39677
rect 6411 39628 6412 39668
rect 6452 39628 6453 39668
rect 6411 39619 6453 39628
rect 6220 39031 6260 39040
rect 6315 39080 6357 39089
rect 6315 39040 6316 39080
rect 6356 39040 6357 39080
rect 6315 39031 6357 39040
rect 6604 39080 6644 40636
rect 6988 40601 7028 40963
rect 6987 40592 7029 40601
rect 6987 40552 6988 40592
rect 7028 40552 7029 40592
rect 6987 40543 7029 40552
rect 6795 39668 6837 39677
rect 6795 39628 6796 39668
rect 6836 39628 6837 39668
rect 6795 39619 6837 39628
rect 6892 39668 6932 39679
rect 6796 39534 6836 39619
rect 6892 39593 6932 39628
rect 6891 39584 6933 39593
rect 6891 39544 6892 39584
rect 6932 39544 6933 39584
rect 6891 39535 6933 39544
rect 6988 39416 7028 40543
rect 6892 39376 7028 39416
rect 6604 39031 6644 39040
rect 6796 39080 6836 39089
rect 6028 38996 6068 39005
rect 5836 38956 6028 38996
rect 5740 38872 5876 38912
rect 5204 38704 5492 38744
rect 5643 38744 5685 38753
rect 5643 38704 5644 38744
rect 5684 38704 5685 38744
rect 5164 38695 5204 38704
rect 5643 38695 5685 38704
rect 4928 38576 5296 38585
rect 4968 38536 5010 38576
rect 5050 38536 5092 38576
rect 5132 38536 5174 38576
rect 5214 38536 5256 38576
rect 4928 38527 5296 38536
rect 5643 38576 5685 38585
rect 5643 38536 5644 38576
rect 5684 38536 5685 38576
rect 5643 38527 5685 38536
rect 5644 38240 5684 38527
rect 5644 38165 5684 38200
rect 5643 38156 5685 38165
rect 5643 38116 5644 38156
rect 5684 38116 5685 38156
rect 5643 38107 5685 38116
rect 5644 38076 5684 38107
rect 5836 37820 5876 38872
rect 6028 38081 6068 38956
rect 6411 38996 6453 39005
rect 6411 38956 6412 38996
rect 6452 38956 6453 38996
rect 6411 38947 6453 38956
rect 6412 38862 6452 38947
rect 6796 38921 6836 39040
rect 6795 38912 6837 38921
rect 6795 38872 6796 38912
rect 6836 38872 6837 38912
rect 6795 38863 6837 38872
rect 6603 38744 6645 38753
rect 6603 38704 6604 38744
rect 6644 38704 6645 38744
rect 6603 38695 6645 38704
rect 6795 38744 6837 38753
rect 6795 38704 6796 38744
rect 6836 38704 6837 38744
rect 6795 38695 6837 38704
rect 6412 38240 6452 38249
rect 6452 38200 6548 38240
rect 6412 38191 6452 38200
rect 6027 38072 6069 38081
rect 6027 38032 6028 38072
rect 6068 38032 6069 38072
rect 6027 38023 6069 38032
rect 6028 37938 6068 38023
rect 6508 37913 6548 38200
rect 6507 37904 6549 37913
rect 6507 37864 6508 37904
rect 6548 37864 6549 37904
rect 6507 37855 6549 37864
rect 4780 37780 5108 37820
rect 4779 37484 4821 37493
rect 4779 37444 4780 37484
rect 4820 37444 4821 37484
rect 4779 37435 4821 37444
rect 4683 37232 4725 37241
rect 4683 37192 4684 37232
rect 4724 37192 4725 37232
rect 4683 37183 4725 37192
rect 4587 37148 4629 37157
rect 4587 37108 4588 37148
rect 4628 37108 4629 37148
rect 4587 37099 4629 37108
rect 4684 37098 4724 37183
rect 4684 36728 4724 36737
rect 4780 36728 4820 37435
rect 5068 37400 5108 37780
rect 5740 37780 5876 37820
rect 5931 37820 5973 37829
rect 5931 37780 5932 37820
rect 5972 37780 5973 37820
rect 5068 37351 5108 37360
rect 5164 37400 5204 37409
rect 5164 37241 5204 37360
rect 5547 37400 5589 37409
rect 5547 37360 5548 37400
rect 5588 37360 5589 37400
rect 5547 37351 5589 37360
rect 5644 37400 5684 37409
rect 5548 37266 5588 37351
rect 5163 37232 5205 37241
rect 5163 37192 5164 37232
rect 5204 37192 5205 37232
rect 5163 37183 5205 37192
rect 5644 37157 5684 37360
rect 5643 37148 5685 37157
rect 5643 37108 5644 37148
rect 5684 37108 5685 37148
rect 5643 37099 5685 37108
rect 4928 37064 5296 37073
rect 4968 37024 5010 37064
rect 5050 37024 5092 37064
rect 5132 37024 5174 37064
rect 5214 37024 5256 37064
rect 4928 37015 5296 37024
rect 5547 37064 5589 37073
rect 5547 37024 5548 37064
rect 5588 37024 5589 37064
rect 5547 37015 5589 37024
rect 4724 36688 4820 36728
rect 4684 36679 4724 36688
rect 4492 36604 4628 36644
rect 4203 36560 4245 36569
rect 4203 36520 4204 36560
rect 4244 36520 4245 36560
rect 4203 36511 4245 36520
rect 4204 34460 4244 36511
rect 4492 36476 4532 36485
rect 4396 36436 4492 36476
rect 4299 36056 4341 36065
rect 4299 36016 4300 36056
rect 4340 36016 4341 36056
rect 4299 36007 4341 36016
rect 4300 35300 4340 36007
rect 4396 35888 4436 36436
rect 4492 36427 4532 36436
rect 4396 35839 4436 35848
rect 4492 35888 4532 35897
rect 4492 35729 4532 35848
rect 4491 35720 4533 35729
rect 4491 35680 4492 35720
rect 4532 35680 4533 35720
rect 4491 35671 4533 35680
rect 4491 35552 4533 35561
rect 4491 35512 4492 35552
rect 4532 35512 4533 35552
rect 4491 35503 4533 35512
rect 4395 35300 4437 35309
rect 4300 35260 4396 35300
rect 4436 35260 4437 35300
rect 4395 35251 4437 35260
rect 4396 35216 4436 35251
rect 4396 35165 4436 35176
rect 4204 34420 4436 34460
rect 4300 34208 4340 34217
rect 4108 34159 4148 34168
rect 4204 34168 4300 34208
rect 4204 34040 4244 34168
rect 4300 34159 4340 34168
rect 4012 34000 4244 34040
rect 4107 33872 4149 33881
rect 4107 33832 4108 33872
rect 4148 33832 4149 33872
rect 4107 33823 4149 33832
rect 3820 33704 3860 33713
rect 3820 33545 3860 33664
rect 4011 33704 4053 33713
rect 4011 33664 4012 33704
rect 4052 33664 4053 33704
rect 4011 33655 4053 33664
rect 4108 33704 4148 33823
rect 4299 33788 4341 33797
rect 4299 33748 4300 33788
rect 4340 33748 4341 33788
rect 4299 33739 4341 33748
rect 4108 33655 4148 33664
rect 4300 33704 4340 33739
rect 4012 33570 4052 33655
rect 4300 33653 4340 33664
rect 3819 33536 3861 33545
rect 3819 33496 3820 33536
rect 3860 33496 3861 33536
rect 3819 33487 3861 33496
rect 4108 33536 4148 33545
rect 3688 33284 4056 33293
rect 3728 33244 3770 33284
rect 3810 33244 3852 33284
rect 3892 33244 3934 33284
rect 3974 33244 4016 33284
rect 3688 33235 4056 33244
rect 4108 32873 4148 33496
rect 4396 33032 4436 34420
rect 4492 34385 4532 35503
rect 4491 34376 4533 34385
rect 4491 34336 4492 34376
rect 4532 34336 4533 34376
rect 4491 34327 4533 34336
rect 4492 34242 4532 34327
rect 4300 32992 4436 33032
rect 3628 32864 3668 32873
rect 3531 32696 3573 32705
rect 3531 32656 3532 32696
rect 3572 32656 3573 32696
rect 3531 32647 3573 32656
rect 3339 32444 3381 32453
rect 3339 32404 3340 32444
rect 3380 32404 3381 32444
rect 3339 32395 3381 32404
rect 3340 32192 3380 32395
rect 3340 32143 3380 32152
rect 3628 31949 3668 32824
rect 3723 32864 3765 32873
rect 3723 32824 3724 32864
rect 3764 32824 3765 32864
rect 3723 32815 3765 32824
rect 4107 32864 4149 32873
rect 4107 32824 4108 32864
rect 4148 32824 4149 32864
rect 4107 32815 4149 32824
rect 3724 32730 3764 32815
rect 4203 32192 4245 32201
rect 4203 32152 4204 32192
rect 4244 32152 4245 32192
rect 4203 32143 4245 32152
rect 4204 32058 4244 32143
rect 3339 31940 3381 31949
rect 3339 31900 3340 31940
rect 3380 31900 3381 31940
rect 3339 31891 3381 31900
rect 3532 31940 3572 31949
rect 3340 31109 3380 31891
rect 3532 31604 3572 31900
rect 3627 31940 3669 31949
rect 3627 31900 3628 31940
rect 3668 31900 3669 31940
rect 3627 31891 3669 31900
rect 3688 31772 4056 31781
rect 3728 31732 3770 31772
rect 3810 31732 3852 31772
rect 3892 31732 3934 31772
rect 3974 31732 4016 31772
rect 3688 31723 4056 31732
rect 4300 31604 4340 32992
rect 4396 32864 4436 32875
rect 4396 32789 4436 32824
rect 4395 32780 4437 32789
rect 4395 32740 4396 32780
rect 4436 32740 4437 32780
rect 4395 32731 4437 32740
rect 3532 31564 3860 31604
rect 3339 31100 3381 31109
rect 3339 31060 3340 31100
rect 3380 31060 3381 31100
rect 3339 31051 3381 31060
rect 3340 30680 3380 30689
rect 3380 30640 3476 30680
rect 3340 30631 3380 30640
rect 3243 30008 3285 30017
rect 3243 29968 3244 30008
rect 3284 29968 3285 30008
rect 3243 29959 3285 29968
rect 3339 29420 3381 29429
rect 3339 29380 3340 29420
rect 3380 29380 3381 29420
rect 3339 29371 3381 29380
rect 3051 29336 3093 29345
rect 3051 29296 3052 29336
rect 3092 29296 3093 29336
rect 3051 29287 3093 29296
rect 3340 29168 3380 29371
rect 3244 29128 3340 29168
rect 3147 28580 3189 28589
rect 3147 28540 3148 28580
rect 3188 28540 3189 28580
rect 3147 28531 3189 28540
rect 2956 28293 2996 28302
rect 3148 28244 3188 28531
rect 3148 28195 3188 28204
rect 2956 27656 2996 27665
rect 3244 27656 3284 29128
rect 3340 29119 3380 29128
rect 3436 29093 3476 30640
rect 3820 30675 3860 31564
rect 4012 31564 4340 31604
rect 3916 31352 3956 31363
rect 3916 31277 3956 31312
rect 3915 31268 3957 31277
rect 3915 31228 3916 31268
rect 3956 31228 3957 31268
rect 3915 31219 3957 31228
rect 4012 30848 4052 31564
rect 4300 31352 4340 31361
rect 4588 31352 4628 36604
rect 5451 36308 5493 36317
rect 5451 36268 5452 36308
rect 5492 36268 5493 36308
rect 5451 36259 5493 36268
rect 4971 36140 5013 36149
rect 4971 36100 4972 36140
rect 5012 36100 5013 36140
rect 4971 36091 5013 36100
rect 4972 35972 5012 36091
rect 4972 35923 5012 35932
rect 4875 35888 4917 35897
rect 4875 35848 4876 35888
rect 4916 35848 4917 35888
rect 4875 35839 4917 35848
rect 5452 35888 5492 36259
rect 5452 35839 5492 35848
rect 4876 35754 4916 35839
rect 5548 35729 5588 37015
rect 5547 35720 5589 35729
rect 5547 35680 5548 35720
rect 5588 35680 5589 35720
rect 5547 35671 5589 35680
rect 4928 35552 5296 35561
rect 4968 35512 5010 35552
rect 5050 35512 5092 35552
rect 5132 35512 5174 35552
rect 5214 35512 5256 35552
rect 4928 35503 5296 35512
rect 4683 35300 4725 35309
rect 4683 35260 4684 35300
rect 4724 35260 4725 35300
rect 5548 35300 5588 35671
rect 5548 35260 5684 35300
rect 4683 35251 4725 35260
rect 4204 31312 4300 31352
rect 4340 31312 4628 31352
rect 4107 31184 4149 31193
rect 4107 31144 4108 31184
rect 4148 31144 4149 31184
rect 4107 31135 4149 31144
rect 4108 31050 4148 31135
rect 4012 30799 4052 30808
rect 3820 30626 3860 30635
rect 3688 30260 4056 30269
rect 3728 30220 3770 30260
rect 3810 30220 3852 30260
rect 3892 30220 3934 30260
rect 3974 30220 4016 30260
rect 3688 30211 4056 30220
rect 3531 30176 3573 30185
rect 3531 30136 3532 30176
rect 3572 30136 3573 30176
rect 3531 30127 3573 30136
rect 3532 29840 3572 30127
rect 3532 29791 3572 29800
rect 3915 29168 3957 29177
rect 3915 29128 3916 29168
rect 3956 29128 3957 29168
rect 3915 29119 3957 29128
rect 3435 29084 3477 29093
rect 3435 29044 3436 29084
rect 3476 29044 3477 29084
rect 3435 29035 3477 29044
rect 3916 29034 3956 29119
rect 4204 29000 4244 31312
rect 4300 31303 4340 31312
rect 4684 31268 4724 35251
rect 5644 35216 5684 35260
rect 5548 35176 5644 35216
rect 5740 35216 5780 37780
rect 5931 37771 5973 37780
rect 5932 37073 5972 37771
rect 6123 37568 6165 37577
rect 6123 37528 6124 37568
rect 6164 37528 6165 37568
rect 6123 37519 6165 37528
rect 6124 37400 6164 37519
rect 6124 37351 6164 37360
rect 5931 37064 5973 37073
rect 5931 37024 5932 37064
rect 5972 37024 5973 37064
rect 5931 37015 5973 37024
rect 5932 36728 5972 37015
rect 6508 36905 6548 37855
rect 6604 37414 6644 38695
rect 6699 38660 6741 38669
rect 6699 38620 6700 38660
rect 6740 38620 6741 38660
rect 6699 38611 6741 38620
rect 6700 38333 6740 38611
rect 6796 38417 6836 38695
rect 6795 38408 6837 38417
rect 6795 38368 6796 38408
rect 6836 38368 6837 38408
rect 6795 38359 6837 38368
rect 6699 38324 6741 38333
rect 6699 38284 6700 38324
rect 6740 38284 6741 38324
rect 6699 38275 6741 38284
rect 6604 37365 6644 37374
rect 6796 37325 6836 37410
rect 6795 37316 6837 37325
rect 6795 37276 6796 37316
rect 6836 37276 6837 37316
rect 6795 37267 6837 37276
rect 6796 37064 6836 37267
rect 6700 37024 6836 37064
rect 6507 36896 6549 36905
rect 6507 36856 6508 36896
rect 6548 36856 6549 36896
rect 6507 36847 6549 36856
rect 6124 36812 6164 36821
rect 6164 36772 6452 36812
rect 6124 36763 6164 36772
rect 5932 36679 5972 36688
rect 6412 36728 6452 36772
rect 6412 36679 6452 36688
rect 6507 36728 6549 36737
rect 6507 36688 6508 36728
rect 6548 36688 6549 36728
rect 6507 36679 6549 36688
rect 6508 36594 6548 36679
rect 6603 35972 6645 35981
rect 6603 35932 6604 35972
rect 6644 35932 6645 35972
rect 6603 35923 6645 35932
rect 5932 35893 5972 35902
rect 5836 35384 5876 35393
rect 5932 35384 5972 35853
rect 6412 35888 6452 35897
rect 5876 35344 5972 35384
rect 6124 35720 6164 35729
rect 5836 35335 5876 35344
rect 6028 35216 6068 35227
rect 6124 35225 6164 35680
rect 6316 35720 6356 35729
rect 5740 35176 5876 35216
rect 5355 35132 5397 35141
rect 5355 35092 5356 35132
rect 5396 35092 5397 35132
rect 5355 35083 5397 35092
rect 5356 34217 5396 35083
rect 5355 34208 5397 34217
rect 5355 34168 5356 34208
rect 5396 34168 5397 34208
rect 5355 34159 5397 34168
rect 4928 34040 5296 34049
rect 4968 34000 5010 34040
rect 5050 34000 5092 34040
rect 5132 34000 5174 34040
rect 5214 34000 5256 34040
rect 4928 33991 5296 34000
rect 4928 32528 5296 32537
rect 4968 32488 5010 32528
rect 5050 32488 5092 32528
rect 5132 32488 5174 32528
rect 5214 32488 5256 32528
rect 4928 32479 5296 32488
rect 5356 32024 5396 34159
rect 5548 33704 5588 35176
rect 5644 35167 5684 35176
rect 5740 34376 5780 34385
rect 5740 34217 5780 34336
rect 5739 34208 5781 34217
rect 5739 34168 5740 34208
rect 5780 34168 5781 34208
rect 5739 34159 5781 34168
rect 5836 34040 5876 35176
rect 6028 35141 6068 35176
rect 6123 35216 6165 35225
rect 6123 35176 6124 35216
rect 6164 35176 6165 35216
rect 6123 35167 6165 35176
rect 6027 35132 6069 35141
rect 6027 35092 6028 35132
rect 6068 35092 6069 35132
rect 6027 35083 6069 35092
rect 6027 34796 6069 34805
rect 6027 34756 6028 34796
rect 6068 34756 6069 34796
rect 6027 34747 6069 34756
rect 6028 34208 6068 34747
rect 6124 34553 6164 35167
rect 6123 34544 6165 34553
rect 6123 34504 6124 34544
rect 6164 34504 6165 34544
rect 6123 34495 6165 34504
rect 6219 34376 6261 34385
rect 6219 34336 6220 34376
rect 6260 34336 6261 34376
rect 6219 34327 6261 34336
rect 6316 34376 6356 35680
rect 6412 35309 6452 35848
rect 6508 35888 6548 35897
rect 6411 35300 6453 35309
rect 6411 35260 6412 35300
rect 6452 35260 6453 35300
rect 6411 35251 6453 35260
rect 6508 35057 6548 35848
rect 6604 35888 6644 35923
rect 6604 35837 6644 35848
rect 6700 35636 6740 37024
rect 6795 36896 6837 36905
rect 6795 36856 6796 36896
rect 6836 36856 6837 36896
rect 6892 36896 6932 39376
rect 6987 38996 7029 39005
rect 6987 38956 6988 38996
rect 7028 38956 7029 38996
rect 6987 38947 7029 38956
rect 6988 38862 7028 38947
rect 6988 37652 7028 37661
rect 7084 37652 7124 41635
rect 7180 40685 7220 42928
rect 7372 41609 7412 42928
rect 7564 41693 7604 42928
rect 7756 41777 7796 42928
rect 7755 41768 7797 41777
rect 7755 41728 7756 41768
rect 7796 41728 7797 41768
rect 7755 41719 7797 41728
rect 7563 41684 7605 41693
rect 7563 41644 7564 41684
rect 7604 41644 7605 41684
rect 7563 41635 7605 41644
rect 7371 41600 7413 41609
rect 7371 41560 7372 41600
rect 7412 41560 7413 41600
rect 7371 41551 7413 41560
rect 7755 41264 7797 41273
rect 7755 41224 7756 41264
rect 7796 41224 7797 41264
rect 7755 41215 7797 41224
rect 7756 41130 7796 41215
rect 7948 41189 7988 42928
rect 8140 41609 8180 42928
rect 8139 41600 8181 41609
rect 8139 41560 8140 41600
rect 8180 41560 8181 41600
rect 8139 41551 8181 41560
rect 8139 41348 8181 41357
rect 8139 41308 8140 41348
rect 8180 41308 8181 41348
rect 8139 41299 8181 41308
rect 8043 41264 8085 41273
rect 8043 41224 8044 41264
rect 8084 41224 8085 41264
rect 8043 41215 8085 41224
rect 8140 41264 8180 41299
rect 7947 41180 7989 41189
rect 7947 41140 7948 41180
rect 7988 41140 7989 41180
rect 7947 41131 7989 41140
rect 7948 41012 7988 41021
rect 7756 40972 7948 41012
rect 7371 40928 7413 40937
rect 7371 40888 7372 40928
rect 7412 40888 7413 40928
rect 7371 40879 7413 40888
rect 7179 40676 7221 40685
rect 7179 40636 7180 40676
rect 7220 40636 7221 40676
rect 7179 40627 7221 40636
rect 7276 40424 7316 40433
rect 7276 40097 7316 40384
rect 7275 40088 7317 40097
rect 7275 40048 7276 40088
rect 7316 40048 7317 40088
rect 7275 40039 7317 40048
rect 7275 39836 7317 39845
rect 7275 39796 7276 39836
rect 7316 39796 7317 39836
rect 7275 39787 7317 39796
rect 7180 38912 7220 38921
rect 7180 38753 7220 38872
rect 7179 38744 7221 38753
rect 7179 38704 7180 38744
rect 7220 38704 7221 38744
rect 7179 38695 7221 38704
rect 7028 37612 7124 37652
rect 6988 37603 7028 37612
rect 7180 37484 7220 37493
rect 6892 36856 7124 36896
rect 6795 36847 6837 36856
rect 6796 36476 6836 36847
rect 6892 36653 6932 36738
rect 6891 36644 6933 36653
rect 6891 36604 6892 36644
rect 6932 36604 6933 36644
rect 6891 36595 6933 36604
rect 6988 36644 7028 36653
rect 6796 36436 6932 36476
rect 6795 36224 6837 36233
rect 6795 36184 6796 36224
rect 6836 36184 6837 36224
rect 6795 36175 6837 36184
rect 6796 35897 6836 36175
rect 6795 35888 6837 35897
rect 6795 35848 6796 35888
rect 6836 35848 6837 35888
rect 6795 35839 6837 35848
rect 6796 35754 6836 35839
rect 6700 35596 6836 35636
rect 6699 35468 6741 35477
rect 6699 35428 6700 35468
rect 6740 35428 6741 35468
rect 6699 35419 6741 35428
rect 6507 35048 6549 35057
rect 6507 35008 6508 35048
rect 6548 35008 6549 35048
rect 6507 34999 6549 35008
rect 6316 34327 6356 34336
rect 6508 34376 6548 34387
rect 6220 34242 6260 34327
rect 6508 34301 6548 34336
rect 6507 34292 6549 34301
rect 6507 34252 6508 34292
rect 6548 34252 6549 34292
rect 6507 34243 6549 34252
rect 6028 34159 6068 34168
rect 5836 34000 6068 34040
rect 5739 33872 5781 33881
rect 5739 33832 5740 33872
rect 5780 33832 5781 33872
rect 5739 33823 5781 33832
rect 5931 33872 5973 33881
rect 5931 33832 5932 33872
rect 5972 33832 5973 33872
rect 5931 33823 5973 33832
rect 5740 33738 5780 33823
rect 5835 33704 5877 33713
rect 5588 33664 5684 33704
rect 5548 33655 5588 33664
rect 5644 32864 5684 33664
rect 5835 33664 5836 33704
rect 5876 33664 5877 33704
rect 5835 33655 5877 33664
rect 5932 33704 5972 33823
rect 5932 33655 5972 33664
rect 5740 33452 5780 33461
rect 5740 32957 5780 33412
rect 5836 33125 5876 33655
rect 5835 33116 5877 33125
rect 5835 33076 5836 33116
rect 5876 33076 5877 33116
rect 5835 33067 5877 33076
rect 5836 32982 5876 33067
rect 5739 32948 5781 32957
rect 5739 32908 5740 32948
rect 5780 32908 5781 32948
rect 5739 32899 5781 32908
rect 5644 32815 5684 32824
rect 5451 32444 5493 32453
rect 5451 32404 5452 32444
rect 5492 32404 5493 32444
rect 5451 32395 5493 32404
rect 5452 32192 5492 32395
rect 5740 32192 5780 32899
rect 5931 32612 5973 32621
rect 5931 32572 5932 32612
rect 5972 32572 5973 32612
rect 5931 32563 5973 32572
rect 5836 32192 5876 32201
rect 5740 32152 5836 32192
rect 5452 32143 5492 32152
rect 5836 32143 5876 32152
rect 5932 32192 5972 32563
rect 6028 32192 6068 34000
rect 6219 33116 6261 33125
rect 6219 33076 6220 33116
rect 6260 33076 6261 33116
rect 6219 33067 6261 33076
rect 6123 32864 6165 32873
rect 6123 32824 6124 32864
rect 6164 32824 6165 32864
rect 6123 32815 6165 32824
rect 6220 32864 6260 33067
rect 6608 32948 6650 32957
rect 6608 32908 6609 32948
rect 6649 32908 6650 32948
rect 6608 32899 6650 32908
rect 6220 32815 6260 32824
rect 6412 32864 6452 32873
rect 6124 32730 6164 32815
rect 6412 32528 6452 32824
rect 6507 32864 6549 32873
rect 6507 32824 6508 32864
rect 6548 32824 6549 32864
rect 6507 32815 6549 32824
rect 6609 32864 6649 32899
rect 6508 32730 6548 32815
rect 6609 32813 6649 32824
rect 6220 32488 6452 32528
rect 6604 32696 6644 32705
rect 6124 32360 6164 32369
rect 6220 32360 6260 32488
rect 6164 32320 6260 32360
rect 6124 32311 6164 32320
rect 6316 32192 6356 32203
rect 6028 32152 6260 32192
rect 5356 31984 5492 32024
rect 4492 31228 4724 31268
rect 4492 29000 4532 31228
rect 4779 31184 4821 31193
rect 4779 31144 4780 31184
rect 4820 31144 4821 31184
rect 4779 31135 4821 31144
rect 4780 30680 4820 31135
rect 4928 31016 5296 31025
rect 4968 30976 5010 31016
rect 5050 30976 5092 31016
rect 5132 30976 5174 31016
rect 5214 30976 5256 31016
rect 4928 30967 5296 30976
rect 5355 30764 5397 30773
rect 5355 30724 5356 30764
rect 5396 30724 5397 30764
rect 5355 30715 5397 30724
rect 4780 30631 4820 30640
rect 4875 30680 4917 30689
rect 4875 30640 4876 30680
rect 4916 30640 4917 30680
rect 4875 30631 4917 30640
rect 5356 30680 5396 30715
rect 4876 30344 4916 30631
rect 5356 30629 5396 30640
rect 5259 30596 5301 30605
rect 5259 30556 5260 30596
rect 5300 30556 5301 30596
rect 5259 30547 5301 30556
rect 4684 30304 4916 30344
rect 4587 29840 4629 29849
rect 4587 29800 4588 29840
rect 4628 29800 4629 29840
rect 4587 29791 4629 29800
rect 4588 29429 4628 29791
rect 4587 29420 4629 29429
rect 4587 29380 4588 29420
rect 4628 29380 4629 29420
rect 4587 29371 4629 29380
rect 4204 28960 4436 29000
rect 4492 28960 4628 29000
rect 3531 28916 3573 28925
rect 3436 28876 3532 28916
rect 3572 28876 3573 28916
rect 3436 28328 3476 28876
rect 3531 28867 3573 28876
rect 3532 28782 3572 28867
rect 3688 28748 4056 28757
rect 3728 28708 3770 28748
rect 3810 28708 3852 28748
rect 3892 28708 3934 28748
rect 3974 28708 4016 28748
rect 3688 28699 4056 28708
rect 3915 28412 3957 28421
rect 3915 28372 3916 28412
rect 3956 28372 3957 28412
rect 3915 28363 3957 28372
rect 3436 28279 3476 28288
rect 3531 28328 3573 28337
rect 3531 28288 3532 28328
rect 3572 28288 3573 28328
rect 3531 28279 3573 28288
rect 3532 28194 3572 28279
rect 3435 27992 3477 28001
rect 3435 27952 3436 27992
rect 3476 27952 3477 27992
rect 3435 27943 3477 27952
rect 3339 27908 3381 27917
rect 3339 27868 3340 27908
rect 3380 27868 3381 27908
rect 3339 27859 3381 27868
rect 3340 27824 3380 27859
rect 3340 27773 3380 27784
rect 2996 27616 3284 27656
rect 2956 27607 2996 27616
rect 3148 27404 3188 27413
rect 3051 27152 3093 27161
rect 3051 27112 3052 27152
rect 3092 27112 3093 27152
rect 3051 27103 3093 27112
rect 2859 26480 2901 26489
rect 2859 26440 2860 26480
rect 2900 26440 2901 26480
rect 2859 26431 2901 26440
rect 2764 26272 2900 26312
rect 2763 26144 2805 26153
rect 2763 26104 2764 26144
rect 2804 26104 2805 26144
rect 2763 26095 2805 26104
rect 2764 26010 2804 26095
rect 2763 25892 2805 25901
rect 2763 25852 2764 25892
rect 2804 25852 2805 25892
rect 2763 25843 2805 25852
rect 2764 25388 2804 25843
rect 2860 25565 2900 26272
rect 2956 25892 2996 25901
rect 2859 25556 2901 25565
rect 2859 25516 2860 25556
rect 2900 25516 2901 25556
rect 2859 25507 2901 25516
rect 2956 25397 2996 25852
rect 2667 25304 2709 25313
rect 2667 25264 2668 25304
rect 2708 25264 2709 25304
rect 2667 25255 2709 25264
rect 2764 25229 2804 25348
rect 2955 25388 2997 25397
rect 2955 25348 2956 25388
rect 2996 25348 2997 25388
rect 2955 25339 2997 25348
rect 3052 25313 3092 27103
rect 3148 26825 3188 27364
rect 3436 26909 3476 27943
rect 3627 27824 3669 27833
rect 3627 27784 3628 27824
rect 3668 27784 3669 27824
rect 3627 27775 3669 27784
rect 3531 27740 3573 27749
rect 3531 27700 3532 27740
rect 3572 27700 3573 27740
rect 3531 27691 3573 27700
rect 3532 27656 3572 27691
rect 3532 27605 3572 27616
rect 3628 27488 3668 27775
rect 3532 27448 3668 27488
rect 3435 26900 3477 26909
rect 3435 26860 3436 26900
rect 3476 26860 3477 26900
rect 3435 26851 3477 26860
rect 3147 26816 3189 26825
rect 3147 26776 3148 26816
rect 3188 26776 3189 26816
rect 3147 26767 3189 26776
rect 3148 26144 3188 26767
rect 3244 26144 3284 26153
rect 3148 26104 3244 26144
rect 3244 26095 3284 26104
rect 3339 26144 3381 26153
rect 3339 26104 3340 26144
rect 3380 26104 3381 26144
rect 3339 26095 3381 26104
rect 3340 26010 3380 26095
rect 3435 25724 3477 25733
rect 3435 25684 3436 25724
rect 3476 25684 3477 25724
rect 3435 25675 3477 25684
rect 3339 25556 3381 25565
rect 3339 25516 3340 25556
rect 3380 25516 3381 25556
rect 3339 25507 3381 25516
rect 2859 25304 2901 25313
rect 2859 25264 2860 25304
rect 2900 25264 2901 25304
rect 2859 25255 2901 25264
rect 3051 25304 3093 25313
rect 3051 25264 3052 25304
rect 3092 25264 3093 25304
rect 3051 25255 3093 25264
rect 3340 25304 3380 25507
rect 3436 25313 3476 25675
rect 3340 25255 3380 25264
rect 3435 25304 3477 25313
rect 3435 25264 3436 25304
rect 3476 25264 3477 25304
rect 3435 25255 3477 25264
rect 2763 25220 2805 25229
rect 2763 25180 2764 25220
rect 2804 25180 2805 25220
rect 2763 25171 2805 25180
rect 2860 25170 2900 25255
rect 3532 24809 3572 27448
rect 3916 27404 3956 28363
rect 4012 28328 4052 28337
rect 4052 28288 4340 28328
rect 4012 28279 4052 28288
rect 3916 27364 4148 27404
rect 3688 27236 4056 27245
rect 3728 27196 3770 27236
rect 3810 27196 3852 27236
rect 3892 27196 3934 27236
rect 3974 27196 4016 27236
rect 3688 27187 4056 27196
rect 4108 26984 4148 27364
rect 4012 26944 4148 26984
rect 3627 26900 3669 26909
rect 3627 26860 3628 26900
rect 3668 26860 3669 26900
rect 3627 26851 3669 26860
rect 3628 26816 3668 26851
rect 3628 26765 3668 26776
rect 3915 26816 3957 26825
rect 3915 26776 3916 26816
rect 3956 26776 3957 26816
rect 3915 26767 3957 26776
rect 3916 26682 3956 26767
rect 3819 26648 3861 26657
rect 3819 26608 3820 26648
rect 3860 26608 3861 26648
rect 3819 26599 3861 26608
rect 3820 26514 3860 26599
rect 3820 26144 3860 26153
rect 4012 26144 4052 26944
rect 4108 26816 4148 26827
rect 4108 26741 4148 26776
rect 4107 26732 4149 26741
rect 4107 26692 4108 26732
rect 4148 26692 4149 26732
rect 4107 26683 4149 26692
rect 3860 26104 4052 26144
rect 4300 26144 4340 28288
rect 4396 27917 4436 28960
rect 4588 28337 4628 28960
rect 4684 28664 4724 30304
rect 5260 30101 5300 30547
rect 5452 30428 5492 31984
rect 5643 31940 5685 31949
rect 5643 31900 5644 31940
rect 5684 31900 5685 31940
rect 5643 31891 5685 31900
rect 5644 31806 5684 31891
rect 5835 31772 5877 31781
rect 5835 31732 5836 31772
rect 5876 31732 5877 31772
rect 5835 31723 5877 31732
rect 5548 31352 5588 31363
rect 5548 31277 5588 31312
rect 5547 31268 5589 31277
rect 5547 31228 5548 31268
rect 5588 31228 5589 31268
rect 5547 31219 5589 31228
rect 5548 30857 5588 31219
rect 5739 31184 5781 31193
rect 5739 31144 5740 31184
rect 5780 31144 5781 31184
rect 5739 31135 5781 31144
rect 5740 31050 5780 31135
rect 5547 30848 5589 30857
rect 5547 30808 5548 30848
rect 5588 30808 5589 30848
rect 5547 30799 5589 30808
rect 5836 30680 5876 31723
rect 5836 30631 5876 30640
rect 5356 30388 5492 30428
rect 5259 30092 5301 30101
rect 5259 30052 5260 30092
rect 5300 30052 5301 30092
rect 5259 30043 5301 30052
rect 4780 29849 4820 29934
rect 4779 29840 4821 29849
rect 4779 29800 4780 29840
rect 4820 29800 4821 29840
rect 4779 29791 4821 29800
rect 4972 29672 5012 29681
rect 4780 29632 4972 29672
rect 4780 29177 4820 29632
rect 4972 29623 5012 29632
rect 4928 29504 5296 29513
rect 4968 29464 5010 29504
rect 5050 29464 5092 29504
rect 5132 29464 5174 29504
rect 5214 29464 5256 29504
rect 4928 29455 5296 29464
rect 5163 29336 5205 29345
rect 5163 29296 5164 29336
rect 5204 29296 5205 29336
rect 5163 29287 5205 29296
rect 4779 29168 4821 29177
rect 4779 29128 4780 29168
rect 4820 29128 4821 29168
rect 4779 29119 4821 29128
rect 5164 29168 5204 29287
rect 5356 29261 5396 30388
rect 5932 30344 5972 32152
rect 6027 31940 6069 31949
rect 6027 31900 6028 31940
rect 6068 31900 6069 31940
rect 6027 31891 6069 31900
rect 6028 31352 6068 31891
rect 6028 31303 6068 31312
rect 6124 31352 6164 31361
rect 6124 30689 6164 31312
rect 6123 30680 6165 30689
rect 6123 30640 6124 30680
rect 6164 30640 6165 30680
rect 6123 30631 6165 30640
rect 6220 30512 6260 32152
rect 6316 32117 6356 32152
rect 6315 32108 6357 32117
rect 6315 32068 6316 32108
rect 6356 32068 6357 32108
rect 6315 32059 6357 32068
rect 6507 32024 6549 32033
rect 6507 31984 6508 32024
rect 6548 31984 6549 32024
rect 6507 31975 6549 31984
rect 6508 31436 6548 31975
rect 6604 31781 6644 32656
rect 6603 31772 6645 31781
rect 6603 31732 6604 31772
rect 6644 31732 6645 31772
rect 6603 31723 6645 31732
rect 6412 31396 6508 31436
rect 6412 31277 6452 31396
rect 6508 31387 6548 31396
rect 6604 31394 6644 31403
rect 6411 31268 6453 31277
rect 6411 31228 6412 31268
rect 6452 31228 6453 31268
rect 6411 31219 6453 31228
rect 6315 31184 6357 31193
rect 6315 31144 6316 31184
rect 6356 31144 6357 31184
rect 6315 31135 6357 31144
rect 6507 31184 6549 31193
rect 6507 31144 6508 31184
rect 6548 31144 6549 31184
rect 6507 31135 6549 31144
rect 6316 30675 6356 31135
rect 6508 30848 6548 31135
rect 6508 30799 6548 30808
rect 6604 30773 6644 31354
rect 6700 31193 6740 35419
rect 6699 31184 6741 31193
rect 6699 31144 6700 31184
rect 6740 31144 6741 31184
rect 6699 31135 6741 31144
rect 6699 31016 6741 31025
rect 6699 30976 6700 31016
rect 6740 30976 6741 31016
rect 6699 30967 6741 30976
rect 6603 30764 6645 30773
rect 6603 30724 6604 30764
rect 6644 30724 6645 30764
rect 6603 30715 6645 30724
rect 6316 30626 6356 30635
rect 6124 30472 6260 30512
rect 5932 30304 6068 30344
rect 5932 30008 5972 30017
rect 5740 29968 5932 30008
rect 5452 29840 5492 29849
rect 5452 29345 5492 29800
rect 5547 29840 5589 29849
rect 5547 29800 5548 29840
rect 5588 29800 5589 29840
rect 5547 29791 5589 29800
rect 5740 29840 5780 29968
rect 5932 29959 5972 29968
rect 5740 29791 5780 29800
rect 5931 29840 5973 29849
rect 5931 29800 5932 29840
rect 5972 29800 5973 29840
rect 5931 29791 5973 29800
rect 5451 29336 5493 29345
rect 5451 29296 5452 29336
rect 5492 29296 5493 29336
rect 5451 29287 5493 29296
rect 5355 29252 5397 29261
rect 5355 29212 5356 29252
rect 5396 29212 5397 29252
rect 5355 29203 5397 29212
rect 5548 29168 5588 29791
rect 5932 29706 5972 29791
rect 6028 29765 6068 30304
rect 6027 29756 6069 29765
rect 6027 29716 6028 29756
rect 6068 29716 6069 29756
rect 6027 29707 6069 29716
rect 5643 29672 5685 29681
rect 5643 29632 5644 29672
rect 5684 29632 5685 29672
rect 5643 29623 5685 29632
rect 5644 29538 5684 29623
rect 5644 29168 5684 29177
rect 5548 29128 5644 29168
rect 5164 29119 5204 29128
rect 4780 29000 4820 29119
rect 4780 28960 5012 29000
rect 4684 28624 4820 28664
rect 4683 28496 4725 28505
rect 4683 28456 4684 28496
rect 4724 28456 4725 28496
rect 4683 28447 4725 28456
rect 4492 28328 4532 28337
rect 4492 28169 4532 28288
rect 4587 28328 4629 28337
rect 4587 28288 4588 28328
rect 4628 28288 4629 28328
rect 4587 28279 4629 28288
rect 4491 28160 4533 28169
rect 4491 28120 4492 28160
rect 4532 28120 4533 28160
rect 4491 28111 4533 28120
rect 4395 27908 4437 27917
rect 4395 27868 4396 27908
rect 4436 27868 4437 27908
rect 4395 27859 4437 27868
rect 4396 27581 4436 27859
rect 4588 27833 4628 28279
rect 4587 27824 4629 27833
rect 4587 27784 4588 27824
rect 4628 27784 4629 27824
rect 4587 27775 4629 27784
rect 4395 27572 4437 27581
rect 4395 27532 4396 27572
rect 4436 27532 4437 27572
rect 4395 27523 4437 27532
rect 4587 27572 4629 27581
rect 4587 27532 4588 27572
rect 4628 27532 4629 27572
rect 4587 27523 4629 27532
rect 3723 26060 3765 26069
rect 3723 26020 3724 26060
rect 3764 26020 3765 26060
rect 3723 26011 3765 26020
rect 3724 25926 3764 26011
rect 3820 25901 3860 26104
rect 3819 25892 3861 25901
rect 3819 25852 3820 25892
rect 3860 25852 3861 25892
rect 3819 25843 3861 25852
rect 3688 25724 4056 25733
rect 3728 25684 3770 25724
rect 3810 25684 3852 25724
rect 3892 25684 3934 25724
rect 3974 25684 4016 25724
rect 3688 25675 4056 25684
rect 4300 25481 4340 26104
rect 4395 25640 4437 25649
rect 4395 25600 4396 25640
rect 4436 25600 4437 25640
rect 4395 25591 4437 25600
rect 4299 25472 4341 25481
rect 4299 25432 4300 25472
rect 4340 25432 4341 25472
rect 4299 25423 4341 25432
rect 3819 25388 3861 25397
rect 3819 25348 3820 25388
rect 3860 25348 3861 25388
rect 3819 25339 3861 25348
rect 3820 25318 3860 25339
rect 4396 25313 4436 25591
rect 3820 25253 3860 25278
rect 4395 25304 4437 25313
rect 4395 25264 4396 25304
rect 4436 25264 4437 25304
rect 4395 25255 4437 25264
rect 4011 25220 4053 25229
rect 4011 25180 4012 25220
rect 4052 25180 4053 25220
rect 4011 25171 4053 25180
rect 4012 25086 4052 25171
rect 4396 25170 4436 25255
rect 3531 24800 3573 24809
rect 3531 24760 3532 24800
rect 3572 24760 3573 24800
rect 3531 24751 3573 24760
rect 4588 24641 4628 27523
rect 3340 24632 3380 24641
rect 3244 24592 3340 24632
rect 3052 23792 3092 23801
rect 2667 23624 2709 23633
rect 2667 23584 2668 23624
rect 2708 23584 2709 23624
rect 2667 23575 2709 23584
rect 2668 23490 2708 23575
rect 3052 23372 3092 23752
rect 2668 23332 3092 23372
rect 3148 23792 3188 23801
rect 2668 23288 2708 23332
rect 2668 23239 2708 23248
rect 2475 23120 2517 23129
rect 2475 23080 2476 23120
rect 2516 23080 2517 23120
rect 2475 23071 2517 23080
rect 2571 23120 2613 23129
rect 2571 23080 2572 23120
rect 2612 23080 2613 23120
rect 2571 23071 2613 23080
rect 3052 23120 3092 23129
rect 2476 22986 2516 23071
rect 2763 22952 2805 22961
rect 2763 22912 2764 22952
rect 2804 22912 2805 22952
rect 2763 22903 2805 22912
rect 2476 22280 2516 22289
rect 2571 22280 2613 22289
rect 2516 22240 2572 22280
rect 2612 22240 2613 22280
rect 2476 22231 2516 22240
rect 2571 22231 2613 22240
rect 2764 22280 2804 22903
rect 3052 22709 3092 23080
rect 3148 22961 3188 23752
rect 3147 22952 3189 22961
rect 3147 22912 3148 22952
rect 3188 22912 3189 22952
rect 3147 22903 3189 22912
rect 3244 22784 3284 24592
rect 3340 24583 3380 24592
rect 3436 24632 3476 24641
rect 3628 24632 3668 24641
rect 3436 24464 3476 24592
rect 3148 22744 3284 22784
rect 3340 24424 3476 24464
rect 3532 24592 3628 24632
rect 3051 22700 3093 22709
rect 3051 22660 3052 22700
rect 3092 22660 3093 22700
rect 3051 22651 3093 22660
rect 2859 22616 2901 22625
rect 2859 22576 2860 22616
rect 2900 22576 2901 22616
rect 2859 22567 2901 22576
rect 2764 22231 2804 22240
rect 2860 22280 2900 22567
rect 3148 22532 3188 22744
rect 3340 22616 3380 24424
rect 3532 24380 3572 24592
rect 3628 24583 3668 24592
rect 4587 24632 4629 24641
rect 4587 24592 4588 24632
rect 4628 24592 4629 24632
rect 4587 24583 4629 24592
rect 4684 24464 4724 28447
rect 4780 28085 4820 28624
rect 4972 28342 5012 28960
rect 5644 28925 5684 29128
rect 5740 29168 5780 29179
rect 5836 29177 5876 29262
rect 5740 29093 5780 29128
rect 5835 29168 5877 29177
rect 5835 29128 5836 29168
rect 5876 29128 5877 29168
rect 5835 29119 5877 29128
rect 6027 29168 6069 29177
rect 6027 29128 6028 29168
rect 6068 29128 6069 29168
rect 6027 29119 6069 29128
rect 5739 29084 5781 29093
rect 5739 29044 5740 29084
rect 5780 29044 5781 29084
rect 5739 29035 5781 29044
rect 5356 28916 5396 28925
rect 5643 28916 5685 28925
rect 5396 28876 5492 28916
rect 5356 28867 5396 28876
rect 4972 28293 5012 28302
rect 5163 28244 5205 28253
rect 5163 28204 5164 28244
rect 5204 28204 5205 28244
rect 5163 28195 5205 28204
rect 5164 28110 5204 28195
rect 4779 28076 4821 28085
rect 4779 28036 4780 28076
rect 4820 28036 4821 28076
rect 4779 28027 4821 28036
rect 4928 27992 5296 28001
rect 4968 27952 5010 27992
rect 5050 27952 5092 27992
rect 5132 27952 5174 27992
rect 5214 27952 5256 27992
rect 4928 27943 5296 27952
rect 4779 27656 4821 27665
rect 4779 27616 4780 27656
rect 4820 27616 4821 27656
rect 4779 27607 4821 27616
rect 5452 27656 5492 28876
rect 5643 28876 5644 28916
rect 5684 28876 5685 28916
rect 5643 28867 5685 28876
rect 5740 28505 5780 29035
rect 5835 29000 5877 29009
rect 5835 28960 5836 29000
rect 5876 28960 5877 29000
rect 5835 28951 5877 28960
rect 6028 29000 6068 29119
rect 6124 29000 6164 30472
rect 6219 30092 6261 30101
rect 6219 30052 6220 30092
rect 6260 30052 6261 30092
rect 6219 30043 6261 30052
rect 6220 29840 6260 30043
rect 6220 29791 6260 29800
rect 6700 29840 6740 30967
rect 6700 29791 6740 29800
rect 6603 29756 6645 29765
rect 6603 29716 6604 29756
rect 6644 29716 6645 29756
rect 6603 29707 6645 29716
rect 6315 29672 6357 29681
rect 6315 29632 6316 29672
rect 6356 29632 6357 29672
rect 6315 29623 6357 29632
rect 6219 29252 6261 29261
rect 6219 29212 6220 29252
rect 6260 29212 6261 29252
rect 6219 29203 6261 29212
rect 6220 29168 6260 29203
rect 6220 29117 6260 29128
rect 6316 29168 6356 29623
rect 6316 29119 6356 29128
rect 6411 29168 6453 29177
rect 6411 29128 6412 29168
rect 6452 29128 6453 29168
rect 6411 29119 6453 29128
rect 6508 29168 6548 29177
rect 6412 29034 6452 29119
rect 6508 29009 6548 29128
rect 6604 29093 6644 29707
rect 6699 29504 6741 29513
rect 6699 29464 6700 29504
rect 6740 29464 6741 29504
rect 6699 29455 6741 29464
rect 6603 29084 6645 29093
rect 6603 29044 6604 29084
rect 6644 29044 6645 29084
rect 6603 29035 6645 29044
rect 6507 29000 6549 29009
rect 6124 28960 6356 29000
rect 6028 28951 6068 28960
rect 5739 28496 5781 28505
rect 5739 28456 5740 28496
rect 5780 28456 5781 28496
rect 5739 28447 5781 28456
rect 5739 28328 5781 28337
rect 5739 28288 5740 28328
rect 5780 28288 5781 28328
rect 5739 28279 5781 28288
rect 5643 28244 5685 28253
rect 5643 28204 5644 28244
rect 5684 28204 5685 28244
rect 5643 28195 5685 28204
rect 5644 27656 5684 28195
rect 5740 28194 5780 28279
rect 5836 27740 5876 28951
rect 5931 28496 5973 28505
rect 5931 28456 5932 28496
rect 5972 28456 5973 28496
rect 5931 28447 5973 28456
rect 5836 27691 5876 27700
rect 5740 27656 5780 27665
rect 5644 27616 5740 27656
rect 5452 27607 5492 27616
rect 5740 27607 5780 27616
rect 4780 27522 4820 27607
rect 5451 27488 5493 27497
rect 5451 27448 5452 27488
rect 5492 27448 5493 27488
rect 5451 27439 5493 27448
rect 5355 27152 5397 27161
rect 5355 27112 5356 27152
rect 5396 27112 5397 27152
rect 5355 27103 5397 27112
rect 5356 26816 5396 27103
rect 5356 26767 5396 26776
rect 5355 26648 5397 26657
rect 5355 26608 5356 26648
rect 5396 26608 5397 26648
rect 5355 26599 5397 26608
rect 4928 26480 5296 26489
rect 4968 26440 5010 26480
rect 5050 26440 5092 26480
rect 5132 26440 5174 26480
rect 5214 26440 5256 26480
rect 4928 26431 5296 26440
rect 4779 26396 4821 26405
rect 4779 26356 4780 26396
rect 4820 26356 4821 26396
rect 4779 26347 4821 26356
rect 4780 26139 4820 26347
rect 4971 26312 5013 26321
rect 5356 26312 5396 26599
rect 4971 26272 4972 26312
rect 5012 26272 5013 26312
rect 4971 26263 5013 26272
rect 5164 26272 5396 26312
rect 4972 26178 5012 26263
rect 4780 26090 4820 26099
rect 5164 26144 5204 26272
rect 5164 26095 5204 26104
rect 5356 26144 5396 26153
rect 5163 25976 5205 25985
rect 5163 25936 5164 25976
rect 5204 25936 5205 25976
rect 5356 25976 5396 26104
rect 5452 26144 5492 27439
rect 5739 27152 5781 27161
rect 5739 27112 5740 27152
rect 5780 27112 5781 27152
rect 5739 27103 5781 27112
rect 5643 26816 5685 26825
rect 5643 26776 5644 26816
rect 5684 26776 5685 26816
rect 5643 26767 5685 26776
rect 5548 26648 5588 26657
rect 5548 26405 5588 26608
rect 5547 26396 5589 26405
rect 5547 26356 5548 26396
rect 5588 26356 5589 26396
rect 5547 26347 5589 26356
rect 5452 26095 5492 26104
rect 5644 25976 5684 26767
rect 5740 26480 5780 27103
rect 5932 26909 5972 28447
rect 6123 27656 6165 27665
rect 6123 27616 6124 27656
rect 6164 27616 6165 27656
rect 6123 27607 6165 27616
rect 6124 27488 6164 27607
rect 6124 27439 6164 27448
rect 6220 26984 6260 26993
rect 5931 26900 5973 26909
rect 5931 26860 5932 26900
rect 5972 26860 5973 26900
rect 5931 26851 5973 26860
rect 5835 26816 5877 26825
rect 5835 26776 5836 26816
rect 5876 26776 5877 26816
rect 5835 26767 5877 26776
rect 5932 26816 5972 26851
rect 6220 26825 6260 26944
rect 5836 26682 5876 26767
rect 5932 26766 5972 26776
rect 6028 26816 6068 26825
rect 6028 26489 6068 26776
rect 6219 26816 6261 26825
rect 6219 26776 6220 26816
rect 6260 26776 6261 26816
rect 6219 26767 6261 26776
rect 6219 26648 6261 26657
rect 6219 26608 6220 26648
rect 6260 26608 6261 26648
rect 6219 26599 6261 26608
rect 6027 26480 6069 26489
rect 5740 26440 5972 26480
rect 5356 25936 5684 25976
rect 5740 26144 5780 26153
rect 5163 25927 5205 25936
rect 5164 25842 5204 25927
rect 5355 25724 5397 25733
rect 5355 25684 5356 25724
rect 5396 25684 5397 25724
rect 5355 25675 5397 25684
rect 4928 24968 5296 24977
rect 4968 24928 5010 24968
rect 5050 24928 5092 24968
rect 5132 24928 5174 24968
rect 5214 24928 5256 24968
rect 4928 24919 5296 24928
rect 4780 24641 4820 24726
rect 4779 24632 4821 24641
rect 4779 24592 4780 24632
rect 4820 24592 4821 24632
rect 4779 24583 4821 24592
rect 4684 24424 4820 24464
rect 3628 24380 3668 24389
rect 3436 24340 3572 24380
rect 3615 24340 3628 24380
rect 3436 23633 3476 24340
rect 3615 24331 3668 24340
rect 3615 24296 3655 24331
rect 3532 24256 3655 24296
rect 3532 23969 3572 24256
rect 3688 24212 4056 24221
rect 3728 24172 3770 24212
rect 3810 24172 3852 24212
rect 3892 24172 3934 24212
rect 3974 24172 4016 24212
rect 3688 24163 4056 24172
rect 3531 23960 3573 23969
rect 3531 23920 3532 23960
rect 3572 23920 3573 23960
rect 3531 23911 3573 23920
rect 4011 23960 4053 23969
rect 4011 23920 4012 23960
rect 4052 23920 4053 23960
rect 4011 23911 4053 23920
rect 3531 23792 3573 23801
rect 3531 23752 3532 23792
rect 3572 23752 3573 23792
rect 3531 23743 3573 23752
rect 3628 23792 3668 23801
rect 3532 23658 3572 23743
rect 3435 23624 3477 23633
rect 3435 23584 3436 23624
rect 3476 23584 3477 23624
rect 3435 23575 3477 23584
rect 3628 22868 3668 23752
rect 3148 22483 3188 22492
rect 3244 22576 3380 22616
rect 3532 22828 3668 22868
rect 4012 22868 4052 23911
rect 4108 23792 4148 23801
rect 4108 23045 4148 23752
rect 4588 23797 4628 23806
rect 4492 23288 4532 23297
rect 4588 23288 4628 23757
rect 4780 23708 4820 24424
rect 5260 23969 5300 24054
rect 5259 23960 5301 23969
rect 5259 23920 5260 23960
rect 5300 23920 5301 23960
rect 5259 23911 5301 23920
rect 4971 23792 5013 23801
rect 4971 23752 4972 23792
rect 5012 23752 5013 23792
rect 4971 23743 5013 23752
rect 5259 23792 5301 23801
rect 5259 23752 5260 23792
rect 5300 23752 5301 23792
rect 5259 23743 5301 23752
rect 4780 23659 4820 23668
rect 4972 23658 5012 23743
rect 5260 23658 5300 23743
rect 4683 23624 4725 23633
rect 4683 23584 4684 23624
rect 4724 23584 4725 23624
rect 4683 23575 4725 23584
rect 4532 23248 4628 23288
rect 4492 23239 4532 23248
rect 4299 23120 4341 23129
rect 4299 23080 4300 23120
rect 4340 23080 4341 23120
rect 4299 23071 4341 23080
rect 4684 23120 4724 23575
rect 4928 23456 5296 23465
rect 4968 23416 5010 23456
rect 5050 23416 5092 23456
rect 5132 23416 5174 23456
rect 5214 23416 5256 23456
rect 4928 23407 5296 23416
rect 4684 23071 4724 23080
rect 4971 23120 5013 23129
rect 4971 23080 4972 23120
rect 5012 23080 5013 23120
rect 4971 23071 5013 23080
rect 4107 23036 4149 23045
rect 4107 22996 4108 23036
rect 4148 22996 4149 23036
rect 4107 22987 4149 22996
rect 4300 22986 4340 23071
rect 4972 22986 5012 23071
rect 4780 22868 4820 22877
rect 4012 22828 4148 22868
rect 3244 22280 3284 22576
rect 2860 22231 2900 22240
rect 3052 22240 3284 22280
rect 3340 22448 3380 22457
rect 2476 21608 2516 21617
rect 2380 21568 2476 21608
rect 2476 20768 2516 21568
rect 2572 21533 2612 22231
rect 3052 21776 3092 22240
rect 3244 21869 3284 21929
rect 3243 21860 3285 21869
rect 3243 21811 3244 21860
rect 3284 21811 3285 21860
rect 3244 21785 3284 21794
rect 3052 21727 3092 21736
rect 2668 21692 2708 21703
rect 3340 21692 3380 22408
rect 3532 22196 3572 22828
rect 3688 22700 4056 22709
rect 3728 22660 3770 22700
rect 3810 22660 3852 22700
rect 3892 22660 3934 22700
rect 3974 22660 4016 22700
rect 3688 22651 4056 22660
rect 4012 22289 4052 22374
rect 3724 22280 3764 22289
rect 3627 22196 3669 22205
rect 3532 22156 3628 22196
rect 3668 22156 3669 22196
rect 3627 22147 3669 22156
rect 3628 22062 3668 22147
rect 3724 21953 3764 22240
rect 4011 22280 4053 22289
rect 4011 22240 4012 22280
rect 4052 22240 4053 22280
rect 4011 22231 4053 22240
rect 4108 22112 4148 22828
rect 4396 22828 4780 22868
rect 4203 22700 4245 22709
rect 4203 22660 4204 22700
rect 4244 22660 4245 22700
rect 4203 22651 4245 22660
rect 4012 22072 4148 22112
rect 3723 21944 3765 21953
rect 3723 21904 3724 21944
rect 3764 21904 3765 21944
rect 3723 21895 3765 21904
rect 2668 21617 2708 21652
rect 3244 21652 3380 21692
rect 2667 21608 2709 21617
rect 2667 21568 2668 21608
rect 2708 21568 2709 21608
rect 2667 21559 2709 21568
rect 2955 21608 2997 21617
rect 2955 21568 2956 21608
rect 2996 21568 2997 21608
rect 2955 21559 2997 21568
rect 3147 21608 3189 21617
rect 3147 21568 3148 21608
rect 3188 21568 3189 21608
rect 3147 21559 3189 21568
rect 2571 21524 2613 21533
rect 2571 21484 2572 21524
rect 2612 21484 2613 21524
rect 2571 21475 2613 21484
rect 2572 21020 2612 21475
rect 2956 21474 2996 21559
rect 2763 21440 2805 21449
rect 2763 21400 2764 21440
rect 2804 21400 2805 21440
rect 2763 21391 2805 21400
rect 2668 21020 2708 21029
rect 2572 20980 2668 21020
rect 2668 20777 2708 20980
rect 2764 20945 2804 21391
rect 3052 21356 3092 21365
rect 3052 20945 3092 21316
rect 2763 20936 2805 20945
rect 2763 20896 2764 20936
rect 2804 20896 2805 20936
rect 2763 20887 2805 20896
rect 3051 20936 3093 20945
rect 3051 20896 3052 20936
rect 3092 20896 3093 20936
rect 3051 20887 3093 20896
rect 2955 20852 2997 20861
rect 2955 20812 2956 20852
rect 2996 20812 2997 20852
rect 2955 20803 2997 20812
rect 2380 20728 2476 20768
rect 2283 20264 2325 20273
rect 2188 20224 2284 20264
rect 2324 20224 2325 20264
rect 2283 20215 2325 20224
rect 2036 19384 2132 19424
rect 1996 19375 2036 19384
rect 1803 19256 1845 19265
rect 1803 19216 1804 19256
rect 1844 19216 1845 19256
rect 1803 19207 1845 19216
rect 1996 19256 2036 19265
rect 1707 19004 1749 19013
rect 1707 18964 1708 19004
rect 1748 18964 1749 19004
rect 1707 18955 1749 18964
rect 1996 18752 2036 19216
rect 1708 18712 2036 18752
rect 1708 18584 1748 18712
rect 1708 17753 1748 18544
rect 1804 18584 1844 18593
rect 1707 17744 1749 17753
rect 1707 17704 1708 17744
rect 1748 17704 1749 17744
rect 1707 17695 1749 17704
rect 1804 17585 1844 18544
rect 1803 17576 1845 17585
rect 1803 17536 1804 17576
rect 1844 17536 1845 17576
rect 1803 17527 1845 17536
rect 1899 15896 1941 15905
rect 1899 15856 1900 15896
rect 1940 15856 1941 15896
rect 1899 15847 1941 15856
rect 1611 15644 1653 15653
rect 1611 15604 1612 15644
rect 1652 15604 1653 15644
rect 1611 15595 1653 15604
rect 1268 15520 1460 15560
rect 1228 15511 1268 15520
rect 1323 14216 1365 14225
rect 1323 14176 1324 14216
rect 1364 14176 1365 14216
rect 1323 14167 1365 14176
rect 1324 13460 1364 14167
rect 1324 13411 1364 13420
rect 1228 11024 1268 11033
rect 1420 11024 1460 15520
rect 1515 15560 1557 15569
rect 1515 15520 1516 15560
rect 1556 15520 1557 15560
rect 1515 15511 1557 15520
rect 1516 14972 1556 15511
rect 1516 14923 1556 14932
rect 1900 14972 1940 15847
rect 2092 15821 2132 19384
rect 2187 19088 2229 19097
rect 2187 19048 2188 19088
rect 2228 19048 2229 19088
rect 2187 19039 2229 19048
rect 2188 18954 2228 19039
rect 2187 18836 2229 18845
rect 2284 18836 2324 20215
rect 2187 18796 2188 18836
rect 2228 18796 2324 18836
rect 2187 18787 2229 18796
rect 2188 18584 2228 18787
rect 2283 18668 2325 18677
rect 2283 18628 2284 18668
rect 2324 18628 2325 18668
rect 2283 18619 2325 18628
rect 2188 18535 2228 18544
rect 2284 18584 2324 18619
rect 2284 18533 2324 18544
rect 2380 18005 2420 20728
rect 2476 20719 2516 20728
rect 2667 20768 2709 20777
rect 2667 20728 2668 20768
rect 2708 20728 2709 20768
rect 2667 20719 2709 20728
rect 2956 20768 2996 20803
rect 2667 20264 2709 20273
rect 2667 20224 2668 20264
rect 2708 20224 2709 20264
rect 2667 20215 2709 20224
rect 2668 20130 2708 20215
rect 2956 20180 2996 20728
rect 3051 20768 3093 20777
rect 3051 20728 3052 20768
rect 3092 20728 3093 20768
rect 3051 20719 3093 20728
rect 3148 20768 3188 21559
rect 3244 20945 3284 21652
rect 3436 21608 3476 21617
rect 3340 21566 3380 21575
rect 3339 21526 3340 21533
rect 3380 21526 3381 21533
rect 3339 21524 3381 21526
rect 3339 21484 3340 21524
rect 3380 21484 3381 21524
rect 3339 21475 3381 21484
rect 3340 21431 3380 21475
rect 3243 20936 3285 20945
rect 3243 20896 3244 20936
rect 3284 20896 3285 20936
rect 3243 20887 3285 20896
rect 3148 20719 3188 20728
rect 3244 20768 3284 20777
rect 3436 20768 3476 21568
rect 3916 21608 3956 21617
rect 3723 21440 3765 21449
rect 3723 21400 3724 21440
rect 3764 21400 3765 21440
rect 3723 21391 3765 21400
rect 3531 21356 3573 21365
rect 3531 21316 3532 21356
rect 3572 21316 3573 21356
rect 3531 21307 3573 21316
rect 3532 21020 3572 21307
rect 3724 21306 3764 21391
rect 3916 21365 3956 21568
rect 4012 21524 4052 22072
rect 4204 22028 4244 22651
rect 4012 21475 4052 21484
rect 4108 21988 4244 22028
rect 4300 22448 4340 22457
rect 4108 21440 4148 21988
rect 4300 21608 4340 22408
rect 4300 21559 4340 21568
rect 4204 21524 4244 21535
rect 4204 21449 4244 21484
rect 4108 21391 4148 21400
rect 4203 21440 4245 21449
rect 4203 21400 4204 21440
rect 4244 21400 4245 21440
rect 4203 21391 4245 21400
rect 3915 21356 3957 21365
rect 3915 21316 3916 21356
rect 3956 21316 3957 21356
rect 3915 21307 3957 21316
rect 4203 21272 4245 21281
rect 4108 21232 4204 21272
rect 4244 21232 4245 21272
rect 3688 21188 4056 21197
rect 3728 21148 3770 21188
rect 3810 21148 3852 21188
rect 3892 21148 3934 21188
rect 3974 21148 4016 21188
rect 3688 21139 4056 21148
rect 3532 20980 3764 21020
rect 3531 20852 3573 20861
rect 3531 20812 3532 20852
rect 3572 20812 3573 20852
rect 3531 20803 3573 20812
rect 3284 20728 3476 20768
rect 3532 20768 3572 20803
rect 3244 20719 3284 20728
rect 3052 20634 3092 20719
rect 3532 20717 3572 20728
rect 3627 20768 3669 20777
rect 3627 20728 3628 20768
rect 3668 20728 3669 20768
rect 3627 20719 3669 20728
rect 3628 20634 3668 20719
rect 3724 20684 3764 20980
rect 4108 20936 4148 21232
rect 4203 21223 4245 21232
rect 4396 21104 4436 22828
rect 4780 22819 4820 22828
rect 4491 22448 4533 22457
rect 4491 22408 4492 22448
rect 4532 22408 4533 22448
rect 4491 22399 4533 22408
rect 4492 22121 4532 22399
rect 5067 22364 5109 22373
rect 5067 22324 5068 22364
rect 5108 22324 5109 22364
rect 5067 22315 5109 22324
rect 4588 22280 4628 22289
rect 4491 22112 4533 22121
rect 4491 22072 4492 22112
rect 4532 22072 4533 22112
rect 4491 22063 4533 22072
rect 4492 21776 4532 21785
rect 4588 21776 4628 22240
rect 4683 22280 4725 22289
rect 4683 22240 4684 22280
rect 4724 22240 4725 22280
rect 4683 22231 4725 22240
rect 5068 22280 5108 22315
rect 4532 21736 4628 21776
rect 4492 21727 4532 21736
rect 4684 21692 4724 22231
rect 5068 22229 5108 22240
rect 4780 22054 4820 22063
rect 4780 21776 4820 22014
rect 4928 21944 5296 21953
rect 4968 21904 5010 21944
rect 5050 21904 5092 21944
rect 5132 21904 5174 21944
rect 5214 21904 5256 21944
rect 4928 21895 5296 21904
rect 4780 21736 5012 21776
rect 4684 21652 4820 21692
rect 4587 21608 4629 21617
rect 4587 21568 4588 21608
rect 4628 21568 4629 21608
rect 4780 21608 4820 21652
rect 4587 21559 4629 21568
rect 4684 21566 4724 21575
rect 4588 21474 4628 21559
rect 4780 21559 4820 21568
rect 4108 20887 4148 20896
rect 4204 21064 4436 21104
rect 4204 20777 4244 21064
rect 4684 20945 4724 21526
rect 4972 21020 5012 21736
rect 5067 21608 5109 21617
rect 5067 21568 5068 21608
rect 5108 21568 5109 21608
rect 5067 21559 5109 21568
rect 5068 21474 5108 21559
rect 4972 20971 5012 20980
rect 4300 20936 4340 20945
rect 4683 20936 4725 20945
rect 4340 20896 4628 20936
rect 4300 20887 4340 20896
rect 3819 20768 3861 20777
rect 3819 20728 3820 20768
rect 3860 20728 3861 20768
rect 3819 20719 3861 20728
rect 4108 20768 4148 20777
rect 3724 20635 3764 20644
rect 3820 20634 3860 20719
rect 3339 20600 3381 20609
rect 3339 20560 3340 20600
rect 3380 20560 3381 20600
rect 3339 20551 3381 20560
rect 3915 20600 3957 20609
rect 3915 20560 3916 20600
rect 3956 20560 3957 20600
rect 3915 20551 3957 20560
rect 2956 20140 3092 20180
rect 2476 20096 2516 20107
rect 2476 20021 2516 20056
rect 2859 20096 2901 20105
rect 2859 20056 2860 20096
rect 2900 20056 2901 20096
rect 2859 20047 2901 20056
rect 2475 20012 2517 20021
rect 2475 19972 2476 20012
rect 2516 19972 2517 20012
rect 2475 19963 2517 19972
rect 2860 19962 2900 20047
rect 2668 19844 2708 19853
rect 2476 19804 2668 19844
rect 2476 19256 2516 19804
rect 2668 19795 2708 19804
rect 2476 19207 2516 19216
rect 2571 19256 2613 19265
rect 2571 19216 2572 19256
rect 2612 19216 2613 19256
rect 2571 19207 2613 19216
rect 2763 19256 2805 19265
rect 2763 19216 2764 19256
rect 2804 19216 2805 19256
rect 2763 19207 2805 19216
rect 2956 19256 2996 19265
rect 2572 19088 2612 19207
rect 2476 19048 2612 19088
rect 2379 17996 2421 18005
rect 2379 17956 2380 17996
rect 2420 17956 2421 17996
rect 2379 17947 2421 17956
rect 2476 17912 2516 19048
rect 2764 18929 2804 19207
rect 2763 18920 2805 18929
rect 2763 18880 2764 18920
rect 2804 18880 2805 18920
rect 2763 18871 2805 18880
rect 2764 18584 2804 18871
rect 2956 18845 2996 19216
rect 3052 19256 3092 20140
rect 2955 18836 2997 18845
rect 2955 18796 2956 18836
rect 2996 18796 2997 18836
rect 2955 18787 2997 18796
rect 2764 18535 2804 18544
rect 2956 18509 2996 18787
rect 3052 18677 3092 19216
rect 3147 19088 3189 19097
rect 3147 19048 3148 19088
rect 3188 19048 3189 19088
rect 3147 19039 3189 19048
rect 3051 18668 3093 18677
rect 3051 18628 3052 18668
rect 3092 18628 3093 18668
rect 3051 18619 3093 18628
rect 2955 18500 2997 18509
rect 2955 18460 2956 18500
rect 2996 18460 2997 18500
rect 2955 18451 2997 18460
rect 2763 18416 2805 18425
rect 2763 18376 2764 18416
rect 2804 18376 2805 18416
rect 2763 18367 2805 18376
rect 2476 17872 2612 17912
rect 2476 17744 2516 17753
rect 2379 17072 2421 17081
rect 2379 17032 2380 17072
rect 2420 17032 2421 17072
rect 2379 17023 2421 17032
rect 2476 17067 2516 17704
rect 2572 17585 2612 17872
rect 2667 17744 2709 17753
rect 2667 17704 2668 17744
rect 2708 17704 2709 17744
rect 2667 17695 2709 17704
rect 2668 17660 2708 17695
rect 2668 17609 2708 17620
rect 2571 17576 2613 17585
rect 2571 17536 2572 17576
rect 2612 17536 2613 17576
rect 2571 17527 2613 17536
rect 2764 17240 2804 18367
rect 2859 18332 2901 18341
rect 2859 18292 2860 18332
rect 2900 18292 2901 18332
rect 2859 18283 2901 18292
rect 2764 17191 2804 17200
rect 2476 17051 2612 17067
rect 2476 17027 2572 17051
rect 2091 15812 2133 15821
rect 2091 15772 2092 15812
rect 2132 15772 2133 15812
rect 2091 15763 2133 15772
rect 2380 15485 2420 17023
rect 2476 15560 2516 17027
rect 2572 17002 2612 17011
rect 2764 16820 2804 16829
rect 2668 16780 2764 16820
rect 2668 15989 2708 16780
rect 2764 16771 2804 16780
rect 2764 16232 2804 16241
rect 2667 15980 2709 15989
rect 2667 15940 2668 15980
rect 2708 15940 2709 15980
rect 2667 15931 2709 15940
rect 2764 15560 2804 16192
rect 2860 15653 2900 18283
rect 3148 17744 3188 19039
rect 3244 18570 3284 18579
rect 3244 18425 3284 18530
rect 3243 18416 3285 18425
rect 3243 18376 3244 18416
rect 3284 18376 3285 18416
rect 3243 18367 3285 18376
rect 3340 18080 3380 20551
rect 3916 20189 3956 20551
rect 4108 20273 4148 20728
rect 4203 20768 4245 20777
rect 4203 20728 4204 20768
rect 4244 20728 4245 20768
rect 4203 20719 4245 20728
rect 4588 20768 4628 20896
rect 4683 20896 4684 20936
rect 4724 20896 4725 20936
rect 4683 20887 4725 20896
rect 5067 20852 5109 20861
rect 5067 20812 5068 20852
rect 5108 20812 5109 20852
rect 5067 20803 5109 20812
rect 4588 20719 4628 20728
rect 4684 20768 4724 20777
rect 4492 20600 4532 20609
rect 4300 20560 4492 20600
rect 4107 20264 4149 20273
rect 4107 20224 4108 20264
rect 4148 20224 4149 20264
rect 4107 20215 4149 20224
rect 3915 20180 3957 20189
rect 3915 20140 3916 20180
rect 3956 20140 3957 20180
rect 3915 20131 3957 20140
rect 4108 20096 4148 20105
rect 4012 20021 4052 20040
rect 4011 20012 4053 20021
rect 4108 20012 4148 20056
rect 4203 20096 4245 20105
rect 4203 20056 4204 20096
rect 4244 20056 4245 20096
rect 4203 20047 4245 20056
rect 4011 19972 4012 20012
rect 4052 19972 4148 20012
rect 4011 19963 4053 19972
rect 4108 19853 4148 19972
rect 4107 19844 4149 19853
rect 4107 19804 4108 19844
rect 4148 19804 4149 19844
rect 4107 19795 4149 19804
rect 3688 19676 4056 19685
rect 3728 19636 3770 19676
rect 3810 19636 3852 19676
rect 3892 19636 3934 19676
rect 3974 19636 4016 19676
rect 3688 19627 4056 19636
rect 4060 19265 4100 19274
rect 3531 19256 3573 19265
rect 3531 19216 3532 19256
rect 3572 19216 3573 19256
rect 4100 19225 4148 19256
rect 4060 19216 4148 19225
rect 3531 19207 3573 19216
rect 3532 19122 3572 19207
rect 4108 19004 4148 19216
rect 4204 19172 4244 20047
rect 4300 20021 4340 20560
rect 4492 20551 4532 20560
rect 4395 20180 4437 20189
rect 4684 20180 4724 20728
rect 4395 20140 4396 20180
rect 4436 20140 4437 20180
rect 4395 20131 4437 20140
rect 4588 20140 4724 20180
rect 4780 20768 4820 20777
rect 4299 20012 4341 20021
rect 4299 19972 4300 20012
rect 4340 19972 4341 20012
rect 4396 20012 4436 20131
rect 4588 20096 4628 20140
rect 4492 20012 4532 20021
rect 4396 19972 4492 20012
rect 4299 19963 4341 19972
rect 4492 19963 4532 19972
rect 4204 19123 4244 19132
rect 4300 19844 4340 19853
rect 4300 19004 4340 19804
rect 4396 19601 4436 19603
rect 4395 19592 4437 19601
rect 4395 19552 4396 19592
rect 4436 19552 4437 19592
rect 4395 19543 4437 19552
rect 4396 19508 4436 19543
rect 4396 19459 4436 19468
rect 4588 19424 4628 20056
rect 4683 20012 4725 20021
rect 4683 19972 4684 20012
rect 4724 19972 4725 20012
rect 4683 19963 4725 19972
rect 4492 19384 4628 19424
rect 4395 19340 4437 19349
rect 4395 19300 4396 19340
rect 4436 19300 4437 19340
rect 4395 19291 4437 19300
rect 4108 18964 4340 19004
rect 4300 18761 4340 18964
rect 4299 18752 4341 18761
rect 4299 18712 4300 18752
rect 4340 18712 4341 18752
rect 4299 18703 4341 18712
rect 3435 18668 3477 18677
rect 3435 18628 3436 18668
rect 3476 18628 3477 18668
rect 3435 18619 3477 18628
rect 3436 18534 3476 18619
rect 3628 18584 3668 18593
rect 3532 18544 3628 18584
rect 3148 17695 3188 17704
rect 3244 18040 3380 18080
rect 3244 17744 3284 18040
rect 3532 17996 3572 18544
rect 3628 18535 3668 18544
rect 3820 18584 3860 18593
rect 3628 18341 3668 18426
rect 3820 18425 3860 18544
rect 3916 18584 3956 18593
rect 4107 18584 4149 18593
rect 3956 18544 4108 18584
rect 4148 18544 4149 18584
rect 3916 18535 3956 18544
rect 4107 18535 4149 18544
rect 4204 18584 4244 18593
rect 4300 18584 4340 18703
rect 4244 18544 4340 18584
rect 4396 18584 4436 19291
rect 4204 18535 4244 18544
rect 4396 18535 4436 18544
rect 3819 18416 3861 18425
rect 3819 18376 3820 18416
rect 3860 18376 3861 18416
rect 3819 18367 3861 18376
rect 3627 18332 3669 18341
rect 3627 18292 3628 18332
rect 3668 18292 3669 18332
rect 3627 18283 3669 18292
rect 3688 18164 4056 18173
rect 3728 18124 3770 18164
rect 3810 18124 3852 18164
rect 3892 18124 3934 18164
rect 3974 18124 4016 18164
rect 3688 18115 4056 18124
rect 3628 17996 3668 18005
rect 3532 17956 3628 17996
rect 3628 17837 3668 17956
rect 3819 17996 3861 18005
rect 3819 17956 3820 17996
rect 3860 17956 3861 17996
rect 3819 17947 3861 17956
rect 3339 17828 3381 17837
rect 3339 17788 3340 17828
rect 3380 17788 3381 17828
rect 3339 17779 3381 17788
rect 3627 17828 3669 17837
rect 3627 17788 3628 17828
rect 3668 17788 3669 17828
rect 3627 17779 3669 17788
rect 3244 17669 3284 17704
rect 3340 17744 3380 17779
rect 3340 17693 3380 17704
rect 3531 17744 3573 17753
rect 3531 17704 3532 17744
rect 3572 17704 3573 17744
rect 3531 17695 3573 17704
rect 3820 17744 3860 17947
rect 4108 17837 4148 18535
rect 4204 18341 4244 18426
rect 4203 18332 4245 18341
rect 4203 18292 4204 18332
rect 4244 18292 4245 18332
rect 4203 18283 4245 18292
rect 4492 18173 4532 19384
rect 4587 19256 4629 19265
rect 4587 19216 4588 19256
rect 4628 19216 4629 19256
rect 4587 19207 4629 19216
rect 4588 19122 4628 19207
rect 4587 18752 4629 18761
rect 4587 18712 4588 18752
rect 4628 18712 4629 18752
rect 4587 18703 4629 18712
rect 4588 18584 4628 18703
rect 4588 18535 4628 18544
rect 4684 18584 4724 19963
rect 4780 19853 4820 20728
rect 5068 20768 5108 20803
rect 5068 20717 5108 20728
rect 4928 20432 5296 20441
rect 4968 20392 5010 20432
rect 5050 20392 5092 20432
rect 5132 20392 5174 20432
rect 5214 20392 5256 20432
rect 5356 20432 5396 25675
rect 5740 25556 5780 26104
rect 5836 25556 5876 25565
rect 5740 25516 5836 25556
rect 5836 25507 5876 25516
rect 5644 25304 5684 25313
rect 5644 25220 5684 25264
rect 5932 25220 5972 26440
rect 6027 26440 6028 26480
rect 6068 26440 6069 26480
rect 6027 26431 6069 26440
rect 6027 26312 6069 26321
rect 6027 26272 6028 26312
rect 6068 26272 6069 26312
rect 6027 26263 6069 26272
rect 6028 26144 6068 26263
rect 6123 26228 6165 26237
rect 6123 26188 6124 26228
rect 6164 26188 6165 26228
rect 6123 26179 6165 26188
rect 6028 26095 6068 26104
rect 6124 26094 6164 26179
rect 5644 25180 5972 25220
rect 5835 24968 5877 24977
rect 5835 24928 5836 24968
rect 5876 24928 5877 24968
rect 5835 24919 5877 24928
rect 5836 24221 5876 24919
rect 5835 24212 5877 24221
rect 5835 24172 5836 24212
rect 5876 24172 5877 24212
rect 5835 24163 5877 24172
rect 5451 23960 5493 23969
rect 5451 23920 5452 23960
rect 5492 23920 5493 23960
rect 5451 23911 5493 23920
rect 5452 23792 5492 23911
rect 5452 23743 5492 23752
rect 5643 23792 5685 23801
rect 5643 23752 5644 23792
rect 5684 23752 5685 23792
rect 5643 23743 5685 23752
rect 5740 23792 5780 23801
rect 5547 23708 5589 23717
rect 5547 23668 5548 23708
rect 5588 23668 5589 23708
rect 5547 23659 5589 23668
rect 5548 23574 5588 23659
rect 5644 23658 5684 23743
rect 5643 23456 5685 23465
rect 5643 23416 5644 23456
rect 5684 23416 5685 23456
rect 5643 23407 5685 23416
rect 5547 23372 5589 23381
rect 5547 23332 5548 23372
rect 5588 23332 5589 23372
rect 5547 23323 5589 23332
rect 5548 22877 5588 23323
rect 5547 22868 5589 22877
rect 5547 22828 5548 22868
rect 5588 22828 5589 22868
rect 5547 22819 5589 22828
rect 5547 21524 5589 21533
rect 5547 21484 5548 21524
rect 5588 21484 5589 21524
rect 5547 21475 5589 21484
rect 5548 20768 5588 21475
rect 5644 20945 5684 23407
rect 5740 22625 5780 23752
rect 5836 23465 5876 24163
rect 5835 23456 5877 23465
rect 5835 23416 5836 23456
rect 5876 23416 5877 23456
rect 5835 23407 5877 23416
rect 5835 23036 5877 23045
rect 5835 22996 5836 23036
rect 5876 22996 5877 23036
rect 5835 22987 5877 22996
rect 5739 22616 5781 22625
rect 5739 22576 5740 22616
rect 5780 22576 5781 22616
rect 5739 22567 5781 22576
rect 5740 21029 5780 22567
rect 5739 21020 5781 21029
rect 5739 20980 5740 21020
rect 5780 20980 5781 21020
rect 5739 20971 5781 20980
rect 5643 20936 5685 20945
rect 5643 20896 5644 20936
rect 5684 20896 5685 20936
rect 5643 20887 5685 20896
rect 5739 20852 5781 20861
rect 5739 20812 5740 20852
rect 5780 20812 5781 20852
rect 5739 20803 5781 20812
rect 5548 20719 5588 20728
rect 5643 20768 5685 20777
rect 5643 20728 5644 20768
rect 5684 20728 5685 20768
rect 5643 20719 5685 20728
rect 5740 20768 5780 20803
rect 5644 20634 5684 20719
rect 5740 20717 5780 20728
rect 5452 20600 5492 20609
rect 5836 20600 5876 22987
rect 5932 22952 5972 25180
rect 6028 25304 6068 25313
rect 6220 25304 6260 26599
rect 6068 25264 6260 25304
rect 6028 24977 6068 25264
rect 6027 24968 6069 24977
rect 6027 24928 6028 24968
rect 6068 24928 6069 24968
rect 6027 24919 6069 24928
rect 6028 24632 6068 24641
rect 6123 24632 6165 24641
rect 6068 24592 6124 24632
rect 6164 24592 6165 24632
rect 6028 24583 6068 24592
rect 6123 24583 6165 24592
rect 6027 24464 6069 24473
rect 6027 24424 6028 24464
rect 6068 24424 6069 24464
rect 6027 24415 6069 24424
rect 6028 23792 6068 24415
rect 6124 24212 6164 24583
rect 6219 24464 6261 24473
rect 6219 24424 6220 24464
rect 6260 24424 6261 24464
rect 6219 24415 6261 24424
rect 6220 24330 6260 24415
rect 6124 24172 6260 24212
rect 6028 23743 6068 23752
rect 6124 23792 6164 23801
rect 6124 23549 6164 23752
rect 6123 23540 6165 23549
rect 6123 23500 6124 23540
rect 6164 23500 6165 23540
rect 6123 23491 6165 23500
rect 6220 23120 6260 24172
rect 6220 23071 6260 23080
rect 5932 22912 6260 22952
rect 5931 22616 5973 22625
rect 5931 22576 5932 22616
rect 5972 22576 5973 22616
rect 5931 22567 5973 22576
rect 5932 21617 5972 22567
rect 6027 21776 6069 21785
rect 6027 21736 6028 21776
rect 6068 21736 6069 21776
rect 6027 21727 6069 21736
rect 5931 21608 5973 21617
rect 5931 21568 5932 21608
rect 5972 21568 5973 21608
rect 5931 21559 5973 21568
rect 6028 21020 6068 21727
rect 6123 21440 6165 21449
rect 6123 21400 6124 21440
rect 6164 21400 6165 21440
rect 6123 21391 6165 21400
rect 5492 20560 5588 20600
rect 5452 20551 5492 20560
rect 5356 20392 5492 20432
rect 4928 20383 5296 20392
rect 4972 20096 5012 20105
rect 4779 19844 4821 19853
rect 4779 19804 4780 19844
rect 4820 19804 4821 19844
rect 4779 19795 4821 19804
rect 4780 19349 4820 19795
rect 4875 19760 4917 19769
rect 4875 19720 4876 19760
rect 4916 19720 4917 19760
rect 4875 19711 4917 19720
rect 4779 19340 4821 19349
rect 4779 19300 4780 19340
rect 4820 19300 4821 19340
rect 4779 19291 4821 19300
rect 4876 19265 4916 19711
rect 4972 19601 5012 20056
rect 5259 20096 5301 20105
rect 5259 20056 5260 20096
rect 5300 20056 5301 20096
rect 5259 20047 5301 20056
rect 5356 20096 5396 20105
rect 5260 19962 5300 20047
rect 4971 19592 5013 19601
rect 4971 19552 4972 19592
rect 5012 19552 5013 19592
rect 4971 19543 5013 19552
rect 4875 19256 4917 19265
rect 4875 19216 4876 19256
rect 4916 19216 4917 19256
rect 4875 19207 4917 19216
rect 4928 18920 5296 18929
rect 4968 18880 5010 18920
rect 5050 18880 5092 18920
rect 5132 18880 5174 18920
rect 5214 18880 5256 18920
rect 4928 18871 5296 18880
rect 5356 18761 5396 20056
rect 4875 18752 4917 18761
rect 4875 18712 4876 18752
rect 4916 18712 4917 18752
rect 4875 18703 4917 18712
rect 5355 18752 5397 18761
rect 5355 18712 5356 18752
rect 5396 18712 5397 18752
rect 5355 18703 5397 18712
rect 4876 18618 4916 18703
rect 4684 18535 4724 18544
rect 4780 18584 4820 18593
rect 4780 18416 4820 18544
rect 5067 18584 5109 18593
rect 5067 18544 5068 18584
rect 5108 18544 5109 18584
rect 5067 18535 5109 18544
rect 4684 18376 4820 18416
rect 4587 18332 4629 18341
rect 4684 18332 4724 18376
rect 4587 18292 4588 18332
rect 4628 18292 4724 18332
rect 4587 18283 4629 18292
rect 4203 18164 4245 18173
rect 4203 18124 4204 18164
rect 4244 18124 4245 18164
rect 4203 18115 4245 18124
rect 4491 18164 4533 18173
rect 4491 18124 4492 18164
rect 4532 18124 4533 18164
rect 4491 18115 4533 18124
rect 4779 18164 4821 18173
rect 4779 18124 4780 18164
rect 4820 18124 4821 18164
rect 4779 18115 4821 18124
rect 4107 17828 4149 17837
rect 4107 17788 4108 17828
rect 4148 17788 4149 17828
rect 4107 17779 4149 17788
rect 3820 17695 3860 17704
rect 3243 17660 3285 17669
rect 3243 17620 3244 17660
rect 3284 17620 3285 17660
rect 3243 17611 3285 17620
rect 3435 17660 3477 17669
rect 3435 17620 3436 17660
rect 3476 17620 3477 17660
rect 3435 17611 3477 17620
rect 3052 17576 3092 17585
rect 3244 17580 3284 17611
rect 2956 17536 3052 17576
rect 2956 16661 2996 17536
rect 3052 17527 3092 17536
rect 3148 17072 3188 17081
rect 2955 16652 2997 16661
rect 2955 16612 2956 16652
rect 2996 16612 2997 16652
rect 2955 16603 2997 16612
rect 3148 16493 3188 17032
rect 3339 16652 3381 16661
rect 3339 16612 3340 16652
rect 3380 16612 3381 16652
rect 3339 16603 3381 16612
rect 3147 16484 3189 16493
rect 3147 16444 3148 16484
rect 3188 16444 3189 16484
rect 3147 16435 3189 16444
rect 2955 16400 2997 16409
rect 2955 16360 2956 16400
rect 2996 16360 2997 16400
rect 2955 16351 2997 16360
rect 3243 16400 3285 16409
rect 3243 16360 3244 16400
rect 3284 16360 3285 16400
rect 3243 16351 3285 16360
rect 2956 16266 2996 16351
rect 3244 16232 3284 16351
rect 3244 16183 3284 16192
rect 3340 16064 3380 16603
rect 3436 16232 3476 17611
rect 3532 17610 3572 17695
rect 3688 16652 4056 16661
rect 3728 16612 3770 16652
rect 3810 16612 3852 16652
rect 3892 16612 3934 16652
rect 3974 16612 4016 16652
rect 3688 16603 4056 16612
rect 3723 16484 3765 16493
rect 3723 16444 3724 16484
rect 3764 16444 3765 16484
rect 3723 16435 3765 16444
rect 3532 16232 3572 16241
rect 3436 16192 3532 16232
rect 3532 16183 3572 16192
rect 3244 16024 3380 16064
rect 3628 16148 3668 16157
rect 3147 15980 3189 15989
rect 3147 15940 3148 15980
rect 3188 15940 3189 15980
rect 3147 15931 3189 15940
rect 2859 15644 2901 15653
rect 2859 15604 2860 15644
rect 2900 15604 2901 15644
rect 2859 15595 2901 15604
rect 2516 15520 2804 15560
rect 3148 15560 3188 15931
rect 2476 15511 2516 15520
rect 2379 15476 2421 15485
rect 2379 15436 2380 15476
rect 2420 15436 2421 15476
rect 2379 15427 2421 15436
rect 1900 14923 1940 14932
rect 2283 14888 2325 14897
rect 2283 14848 2284 14888
rect 2324 14848 2325 14888
rect 2283 14839 2325 14848
rect 1708 14804 1748 14813
rect 1612 14764 1708 14804
rect 1515 14552 1557 14561
rect 1515 14512 1516 14552
rect 1556 14512 1557 14552
rect 1515 14503 1557 14512
rect 1516 14216 1556 14503
rect 1516 14167 1556 14176
rect 1515 13292 1557 13301
rect 1515 13252 1516 13292
rect 1556 13252 1557 13292
rect 1515 13243 1557 13252
rect 1516 13158 1556 13243
rect 1515 12872 1557 12881
rect 1515 12832 1516 12872
rect 1556 12832 1557 12872
rect 1515 12823 1557 12832
rect 1516 12368 1556 12823
rect 1612 12377 1652 14764
rect 1708 14755 1748 14764
rect 2091 14804 2133 14813
rect 2091 14764 2092 14804
rect 2132 14764 2133 14804
rect 2091 14755 2133 14764
rect 2092 14670 2132 14755
rect 1995 14468 2037 14477
rect 1995 14428 1996 14468
rect 2036 14428 2037 14468
rect 1995 14419 2037 14428
rect 1707 14048 1749 14057
rect 1707 14008 1708 14048
rect 1748 14008 1749 14048
rect 1707 13999 1749 14008
rect 1708 13964 1748 13999
rect 1708 13913 1748 13924
rect 1899 13880 1941 13889
rect 1899 13840 1900 13880
rect 1940 13840 1941 13880
rect 1899 13831 1941 13840
rect 1900 13746 1940 13831
rect 1803 13544 1845 13553
rect 1803 13504 1804 13544
rect 1844 13504 1845 13544
rect 1803 13495 1845 13504
rect 1708 13040 1748 13049
rect 1708 12629 1748 13000
rect 1707 12620 1749 12629
rect 1707 12580 1708 12620
rect 1748 12580 1749 12620
rect 1707 12571 1749 12580
rect 1708 12452 1748 12461
rect 1516 12319 1556 12328
rect 1611 12368 1653 12377
rect 1611 12328 1612 12368
rect 1652 12328 1653 12368
rect 1611 12319 1653 12328
rect 1708 12293 1748 12412
rect 1707 12284 1749 12293
rect 1707 12244 1708 12284
rect 1748 12244 1749 12284
rect 1707 12235 1749 12244
rect 1515 12200 1557 12209
rect 1515 12160 1516 12200
rect 1556 12160 1557 12200
rect 1515 12151 1557 12160
rect 1516 11948 1556 12151
rect 1804 11948 1844 13495
rect 1900 13292 1940 13301
rect 1996 13292 2036 14419
rect 2284 14216 2324 14839
rect 2284 14167 2324 14176
rect 2572 13973 2612 15520
rect 3148 15511 3188 15520
rect 3244 15560 3284 16024
rect 3436 15728 3476 15737
rect 3628 15728 3668 16108
rect 3476 15688 3668 15728
rect 3436 15679 3476 15688
rect 3339 15644 3381 15653
rect 3339 15604 3340 15644
rect 3380 15604 3381 15644
rect 3339 15595 3381 15604
rect 3244 15511 3284 15520
rect 3340 15560 3380 15595
rect 3340 15509 3380 15520
rect 2668 15308 2708 15317
rect 3724 15308 3764 16435
rect 3916 16400 3956 16409
rect 3956 16360 4148 16400
rect 3916 16351 3956 16360
rect 3819 15980 3861 15989
rect 3819 15940 3820 15980
rect 3860 15940 3861 15980
rect 3819 15931 3861 15940
rect 3820 15560 3860 15931
rect 3820 15511 3860 15520
rect 2668 14720 2708 15268
rect 3532 15268 3764 15308
rect 2668 14671 2708 14680
rect 2764 14720 2804 14729
rect 3148 14720 3188 14729
rect 2804 14680 3092 14720
rect 2764 14671 2804 14680
rect 2667 14132 2709 14141
rect 2667 14092 2668 14132
rect 2708 14092 2709 14132
rect 2667 14083 2709 14092
rect 2668 14048 2708 14083
rect 2668 13997 2708 14008
rect 2091 13964 2133 13973
rect 2091 13924 2092 13964
rect 2132 13924 2133 13964
rect 2091 13915 2133 13924
rect 2476 13964 2516 13973
rect 2092 13830 2132 13915
rect 1940 13252 2036 13292
rect 1900 13243 1940 13252
rect 2092 13208 2132 13219
rect 2092 13133 2132 13168
rect 1899 13124 1941 13133
rect 1899 13084 1900 13124
rect 1940 13084 1941 13124
rect 1899 13075 1941 13084
rect 2091 13124 2133 13133
rect 2091 13084 2092 13124
rect 2132 13084 2133 13124
rect 2091 13075 2133 13084
rect 1900 12368 1940 13075
rect 1995 12956 2037 12965
rect 1995 12916 1996 12956
rect 2036 12916 2037 12956
rect 1995 12907 2037 12916
rect 1900 12319 1940 12328
rect 1900 11948 1940 11957
rect 1804 11908 1900 11948
rect 1516 11899 1556 11908
rect 1900 11899 1940 11908
rect 1707 11780 1749 11789
rect 1707 11740 1708 11780
rect 1748 11740 1749 11780
rect 1707 11731 1749 11740
rect 1708 11646 1748 11731
rect 1803 11528 1845 11537
rect 1803 11488 1804 11528
rect 1844 11488 1845 11528
rect 1803 11479 1845 11488
rect 1515 11360 1557 11369
rect 1515 11320 1516 11360
rect 1556 11320 1557 11360
rect 1515 11311 1557 11320
rect 1268 10984 1460 11024
rect 1228 10975 1268 10984
rect 1323 10856 1365 10865
rect 1323 10816 1324 10856
rect 1364 10816 1365 10856
rect 1323 10807 1365 10816
rect 555 9260 597 9269
rect 555 9220 556 9260
rect 596 9220 597 9260
rect 555 9211 597 9220
rect 556 8513 596 9211
rect 555 8504 597 8513
rect 555 8464 556 8504
rect 596 8464 597 8504
rect 555 8455 597 8464
rect 1324 8168 1364 10807
rect 1420 10361 1460 10984
rect 1419 10352 1461 10361
rect 1419 10312 1420 10352
rect 1460 10312 1461 10352
rect 1419 10303 1461 10312
rect 1419 10184 1461 10193
rect 1419 10144 1420 10184
rect 1460 10144 1461 10184
rect 1419 10135 1461 10144
rect 1516 10184 1556 11311
rect 1707 11276 1749 11285
rect 1707 11236 1708 11276
rect 1748 11236 1749 11276
rect 1707 11227 1749 11236
rect 1516 10135 1556 10144
rect 1420 9680 1460 10135
rect 1611 10016 1653 10025
rect 1611 9976 1612 10016
rect 1652 9976 1653 10016
rect 1611 9967 1653 9976
rect 1516 9680 1556 9689
rect 1420 9640 1516 9680
rect 1516 9631 1556 9640
rect 1515 8840 1557 8849
rect 1515 8800 1516 8840
rect 1556 8800 1557 8840
rect 1515 8791 1557 8800
rect 1516 8706 1556 8791
rect 1612 8756 1652 9967
rect 1708 9428 1748 11227
rect 1708 9379 1748 9388
rect 1804 8840 1844 11479
rect 1899 10100 1941 10109
rect 1899 10060 1900 10100
rect 1940 10060 1941 10100
rect 1899 10051 1941 10060
rect 1900 9512 1940 10051
rect 1900 9463 1940 9472
rect 1996 8933 2036 12907
rect 2476 12713 2516 13924
rect 2571 13964 2613 13973
rect 2571 13924 2572 13964
rect 2612 13924 2613 13964
rect 2571 13915 2613 13924
rect 2475 12704 2517 12713
rect 2475 12664 2476 12704
rect 2516 12664 2517 12704
rect 2475 12655 2517 12664
rect 2955 12620 2997 12629
rect 2955 12580 2956 12620
rect 2996 12580 2997 12620
rect 2955 12571 2997 12580
rect 2475 12536 2517 12545
rect 2475 12496 2476 12536
rect 2516 12496 2517 12536
rect 2475 12487 2517 12496
rect 2091 12452 2133 12461
rect 2091 12412 2092 12452
rect 2132 12412 2133 12452
rect 2091 12403 2133 12412
rect 2092 12318 2132 12403
rect 2092 11780 2132 11789
rect 2092 9773 2132 11740
rect 2476 11369 2516 12487
rect 2668 11696 2708 11705
rect 2475 11360 2517 11369
rect 2475 11320 2476 11360
rect 2516 11320 2517 11360
rect 2475 11311 2517 11320
rect 2187 11192 2229 11201
rect 2187 11152 2188 11192
rect 2228 11152 2229 11192
rect 2187 11143 2229 11152
rect 2668 11192 2708 11656
rect 2668 11143 2708 11152
rect 2764 11696 2804 11705
rect 2091 9764 2133 9773
rect 2091 9724 2092 9764
rect 2132 9724 2133 9764
rect 2091 9715 2133 9724
rect 1995 8924 2037 8933
rect 1995 8884 1996 8924
rect 2036 8884 2037 8924
rect 1995 8875 2037 8884
rect 1900 8840 1940 8849
rect 1804 8800 1900 8840
rect 1900 8791 1940 8800
rect 1708 8756 1748 8765
rect 1612 8716 1708 8756
rect 1708 8707 1748 8716
rect 1995 8756 2037 8765
rect 1995 8716 1996 8756
rect 2036 8716 2037 8756
rect 1995 8707 2037 8716
rect 2092 8756 2132 8765
rect 1803 8672 1845 8681
rect 1803 8632 1804 8672
rect 1844 8632 1845 8672
rect 1803 8623 1845 8632
rect 1804 8336 1844 8623
rect 1708 8296 1844 8336
rect 1420 8168 1460 8177
rect 1324 8128 1420 8168
rect 1420 8119 1460 8128
rect 1611 7916 1653 7925
rect 1611 7876 1612 7916
rect 1652 7876 1653 7916
rect 1611 7867 1653 7876
rect 1323 7832 1365 7841
rect 1323 7792 1324 7832
rect 1364 7792 1365 7832
rect 1323 7783 1365 7792
rect 1324 7412 1364 7783
rect 1612 7782 1652 7867
rect 1420 7412 1460 7421
rect 1324 7372 1420 7412
rect 1420 7363 1460 7372
rect 1611 7244 1653 7253
rect 1611 7204 1612 7244
rect 1652 7204 1653 7244
rect 1611 7195 1653 7204
rect 1612 7110 1652 7195
rect 1708 6992 1748 8296
rect 1803 8168 1845 8177
rect 1803 8128 1804 8168
rect 1844 8128 1845 8168
rect 1803 8119 1845 8128
rect 1804 8034 1844 8119
rect 1996 7916 2036 8707
rect 2092 8597 2132 8716
rect 2091 8588 2133 8597
rect 2091 8548 2092 8588
rect 2132 8548 2133 8588
rect 2091 8539 2133 8548
rect 2188 8168 2228 11143
rect 2475 11024 2517 11033
rect 2475 10984 2476 11024
rect 2516 10984 2517 11024
rect 2475 10975 2517 10984
rect 2476 10890 2516 10975
rect 2764 10445 2804 11656
rect 2860 10772 2900 10781
rect 2860 10529 2900 10732
rect 2859 10520 2901 10529
rect 2859 10480 2860 10520
rect 2900 10480 2901 10520
rect 2859 10471 2901 10480
rect 2763 10436 2805 10445
rect 2763 10396 2764 10436
rect 2804 10396 2805 10436
rect 2763 10387 2805 10396
rect 2956 10268 2996 12571
rect 3052 11612 3092 14680
rect 3148 13217 3188 14680
rect 3243 14720 3285 14729
rect 3243 14680 3244 14720
rect 3284 14680 3285 14720
rect 3243 14671 3285 14680
rect 3244 14586 3284 14671
rect 3339 13964 3381 13973
rect 3339 13924 3340 13964
rect 3380 13924 3381 13964
rect 3339 13915 3381 13924
rect 3147 13208 3189 13217
rect 3147 13168 3148 13208
rect 3188 13168 3189 13208
rect 3147 13159 3189 13168
rect 3340 13208 3380 13915
rect 3532 13301 3572 15268
rect 3688 15140 4056 15149
rect 3728 15100 3770 15140
rect 3810 15100 3852 15140
rect 3892 15100 3934 15140
rect 3974 15100 4016 15140
rect 3688 15091 4056 15100
rect 4108 14897 4148 16360
rect 4204 15728 4244 18115
rect 4395 18080 4437 18089
rect 4395 18040 4396 18080
rect 4436 18040 4437 18080
rect 4395 18031 4437 18040
rect 4396 17753 4436 18031
rect 4491 17828 4533 17837
rect 4491 17788 4492 17828
rect 4532 17788 4533 17828
rect 4491 17779 4533 17788
rect 4395 17744 4437 17753
rect 4395 17704 4396 17744
rect 4436 17704 4437 17744
rect 4395 17695 4437 17704
rect 4396 17072 4436 17695
rect 4396 17023 4436 17032
rect 4492 17030 4532 17779
rect 4780 17240 4820 18115
rect 5068 17753 5108 18535
rect 5355 18080 5397 18089
rect 5355 18040 5356 18080
rect 5396 18040 5397 18080
rect 5355 18031 5397 18040
rect 5067 17744 5109 17753
rect 5067 17704 5068 17744
rect 5108 17704 5109 17744
rect 5067 17695 5109 17704
rect 5068 17610 5108 17695
rect 5259 17660 5301 17669
rect 5259 17620 5260 17660
rect 5300 17620 5301 17660
rect 5259 17611 5301 17620
rect 5260 17526 5300 17611
rect 4928 17408 5296 17417
rect 4968 17368 5010 17408
rect 5050 17368 5092 17408
rect 5132 17368 5174 17408
rect 5214 17368 5256 17408
rect 4928 17359 5296 17368
rect 4780 17200 5012 17240
rect 4588 17156 4628 17165
rect 4628 17116 4916 17156
rect 4588 17107 4628 17116
rect 4876 17072 4916 17116
rect 4492 16990 4628 17030
rect 4876 17023 4916 17032
rect 4972 17072 5012 17200
rect 4299 16232 4341 16241
rect 4299 16192 4300 16232
rect 4340 16192 4341 16232
rect 4299 16183 4341 16192
rect 4300 16098 4340 16183
rect 4204 15688 4340 15728
rect 4107 14888 4149 14897
rect 4107 14848 4108 14888
rect 4148 14848 4149 14888
rect 4107 14839 4149 14848
rect 3724 14720 3764 14731
rect 3724 14645 3764 14680
rect 4204 14725 4244 14734
rect 3723 14636 3765 14645
rect 3723 14596 3724 14636
rect 3764 14596 3765 14636
rect 3723 14587 3765 14596
rect 4108 14216 4148 14225
rect 4204 14216 4244 14685
rect 4148 14176 4244 14216
rect 4108 14167 4148 14176
rect 4300 14141 4340 15688
rect 4395 14804 4437 14813
rect 4395 14764 4396 14804
rect 4436 14764 4437 14804
rect 4395 14755 4437 14764
rect 4396 14636 4436 14755
rect 4396 14587 4436 14596
rect 4299 14132 4341 14141
rect 4299 14092 4300 14132
rect 4340 14092 4341 14132
rect 4299 14083 4341 14092
rect 3916 14048 3956 14059
rect 3916 13973 3956 14008
rect 3915 13964 3957 13973
rect 3915 13924 3916 13964
rect 3956 13924 3957 13964
rect 3915 13915 3957 13924
rect 3688 13628 4056 13637
rect 3728 13588 3770 13628
rect 3810 13588 3852 13628
rect 3892 13588 3934 13628
rect 3974 13588 4016 13628
rect 3688 13579 4056 13588
rect 3531 13292 3573 13301
rect 3531 13252 3532 13292
rect 3572 13252 3573 13292
rect 3531 13243 3573 13252
rect 3340 13159 3380 13168
rect 3820 13208 3860 13217
rect 3148 11780 3188 13159
rect 3532 13124 3572 13133
rect 3820 13124 3860 13168
rect 3572 13084 3860 13124
rect 3916 13208 3956 13217
rect 3532 13075 3572 13084
rect 3916 12545 3956 13168
rect 4300 13208 4340 14083
rect 4107 12620 4149 12629
rect 4107 12580 4108 12620
rect 4148 12580 4149 12620
rect 4107 12571 4149 12580
rect 3724 12536 3764 12545
rect 3148 11731 3188 11740
rect 3532 12496 3724 12536
rect 3532 11705 3572 12496
rect 3724 12487 3764 12496
rect 3915 12536 3957 12545
rect 3915 12496 3916 12536
rect 3956 12496 3957 12536
rect 3915 12487 3957 12496
rect 4108 12536 4148 12571
rect 4108 12485 4148 12496
rect 3916 12284 3956 12293
rect 3956 12244 4244 12284
rect 3916 12235 3956 12244
rect 3688 12116 4056 12125
rect 3728 12076 3770 12116
rect 3810 12076 3852 12116
rect 3892 12076 3934 12116
rect 3974 12076 4016 12116
rect 3688 12067 4056 12076
rect 4204 11710 4244 12244
rect 3244 11696 3284 11705
rect 3244 11612 3284 11656
rect 3531 11696 3573 11705
rect 3531 11656 3532 11696
rect 3572 11656 3573 11696
rect 3531 11647 3573 11656
rect 3724 11696 3764 11705
rect 4204 11661 4244 11670
rect 3052 11572 3284 11612
rect 3147 11444 3189 11453
rect 3052 11404 3148 11444
rect 3188 11404 3189 11444
rect 3052 10940 3092 11404
rect 3147 11395 3189 11404
rect 3244 11360 3284 11572
rect 3244 11320 3380 11360
rect 3052 10891 3092 10900
rect 2860 10228 2996 10268
rect 2379 10184 2421 10193
rect 2379 10144 2380 10184
rect 2420 10144 2421 10184
rect 2379 10135 2421 10144
rect 2764 10184 2804 10193
rect 2283 9512 2325 9521
rect 2283 9472 2284 9512
rect 2324 9472 2325 9512
rect 2283 9463 2325 9472
rect 2284 8840 2324 9463
rect 2284 8791 2324 8800
rect 1996 7867 2036 7876
rect 2092 8128 2228 8168
rect 2092 7748 2132 8128
rect 2188 8000 2228 8009
rect 2188 7757 2228 7960
rect 1900 7708 2132 7748
rect 2187 7748 2229 7757
rect 2187 7708 2188 7748
rect 2228 7708 2229 7748
rect 1803 7496 1845 7505
rect 1803 7456 1804 7496
rect 1844 7456 1845 7496
rect 1803 7447 1845 7456
rect 1804 7412 1844 7447
rect 1804 7361 1844 7372
rect 1612 6952 1748 6992
rect 1515 6824 1557 6833
rect 1515 6784 1516 6824
rect 1556 6784 1557 6824
rect 1515 6775 1557 6784
rect 1516 6656 1556 6775
rect 1516 6607 1556 6616
rect 1419 5732 1461 5741
rect 1419 5692 1420 5732
rect 1460 5692 1461 5732
rect 1419 5683 1461 5692
rect 1228 5648 1268 5657
rect 1323 5648 1365 5657
rect 1268 5608 1324 5648
rect 1364 5608 1365 5648
rect 1228 5599 1268 5608
rect 1323 5599 1365 5608
rect 1323 4976 1365 4985
rect 1323 4936 1324 4976
rect 1364 4936 1365 4976
rect 1323 4927 1365 4936
rect 1324 4808 1364 4927
rect 1324 4759 1364 4768
rect 1323 4640 1365 4649
rect 1323 4600 1324 4640
rect 1364 4600 1365 4640
rect 1323 4591 1365 4600
rect 1228 4136 1268 4145
rect 1324 4136 1364 4591
rect 1268 4096 1364 4136
rect 1228 4087 1268 4096
rect 363 3884 405 3893
rect 363 3844 364 3884
rect 404 3844 405 3884
rect 363 3835 405 3844
rect 364 1121 404 3835
rect 1420 2381 1460 5683
rect 1516 4892 1556 4901
rect 1516 3977 1556 4852
rect 1515 3968 1557 3977
rect 1515 3928 1516 3968
rect 1556 3928 1557 3968
rect 1515 3919 1557 3928
rect 1612 3380 1652 6952
rect 1900 6656 1940 7708
rect 2187 7699 2229 7708
rect 1995 7412 2037 7421
rect 1995 7372 1996 7412
rect 2036 7372 2037 7412
rect 1995 7363 2037 7372
rect 1996 7244 2036 7363
rect 2380 7328 2420 10135
rect 2571 10100 2613 10109
rect 2571 10060 2572 10100
rect 2612 10060 2613 10100
rect 2571 10051 2613 10060
rect 2475 9932 2517 9941
rect 2475 9892 2476 9932
rect 2516 9892 2517 9932
rect 2475 9883 2517 9892
rect 2476 8756 2516 9883
rect 2476 8707 2516 8716
rect 2475 7580 2517 7589
rect 2475 7540 2476 7580
rect 2516 7540 2517 7580
rect 2475 7531 2517 7540
rect 1996 7195 2036 7204
rect 2284 7288 2420 7328
rect 2187 6992 2229 7001
rect 2187 6952 2188 6992
rect 2228 6952 2229 6992
rect 2187 6943 2229 6952
rect 1995 6908 2037 6917
rect 1995 6868 1996 6908
rect 2036 6868 2037 6908
rect 1995 6859 2037 6868
rect 1900 6607 1940 6616
rect 1803 6572 1845 6581
rect 1803 6532 1804 6572
rect 1844 6532 1845 6572
rect 1803 6523 1845 6532
rect 1708 6413 1748 6498
rect 1707 6404 1749 6413
rect 1707 6364 1708 6404
rect 1748 6364 1749 6404
rect 1707 6355 1749 6364
rect 1707 5480 1749 5489
rect 1707 5440 1708 5480
rect 1748 5440 1749 5480
rect 1707 5431 1749 5440
rect 1708 4808 1748 5431
rect 1708 4759 1748 4768
rect 1708 3380 1748 3389
rect 1612 3340 1708 3380
rect 1708 3331 1748 3340
rect 1515 3212 1557 3221
rect 1515 3172 1516 3212
rect 1556 3172 1557 3212
rect 1515 3163 1557 3172
rect 1516 3078 1556 3163
rect 1708 2708 1748 2717
rect 1804 2708 1844 6523
rect 1996 6320 2036 6859
rect 2188 6858 2228 6943
rect 2091 6656 2133 6665
rect 2091 6616 2092 6656
rect 2132 6616 2133 6656
rect 2091 6607 2133 6616
rect 2092 6404 2132 6607
rect 2284 6413 2324 7288
rect 2380 7160 2420 7169
rect 2476 7160 2516 7531
rect 2420 7120 2516 7160
rect 2092 6355 2132 6364
rect 2283 6404 2325 6413
rect 2283 6364 2284 6404
rect 2324 6364 2325 6404
rect 2283 6355 2325 6364
rect 1900 6280 2036 6320
rect 1900 4892 1940 6280
rect 2284 6236 2324 6245
rect 2187 5900 2229 5909
rect 2187 5860 2188 5900
rect 2228 5860 2229 5900
rect 2187 5851 2229 5860
rect 1995 5396 2037 5405
rect 1995 5356 1996 5396
rect 2036 5356 2037 5396
rect 1995 5347 2037 5356
rect 1900 4843 1940 4852
rect 1899 4136 1941 4145
rect 1899 4096 1900 4136
rect 1940 4096 1941 4136
rect 1899 4087 1941 4096
rect 1900 3632 1940 4087
rect 1900 3583 1940 3592
rect 1899 2792 1941 2801
rect 1899 2752 1900 2792
rect 1940 2752 1941 2792
rect 1899 2743 1941 2752
rect 1748 2668 1844 2708
rect 1708 2659 1748 2668
rect 1900 2658 1940 2743
rect 1996 2708 2036 5347
rect 2092 4985 2132 5070
rect 2091 4976 2133 4985
rect 2091 4936 2092 4976
rect 2132 4936 2133 4976
rect 2091 4927 2133 4936
rect 2188 4808 2228 5851
rect 2284 5153 2324 6196
rect 2380 5648 2420 7120
rect 2476 6393 2516 6415
rect 2476 6329 2516 6353
rect 2475 6320 2517 6329
rect 2475 6280 2476 6320
rect 2516 6280 2517 6320
rect 2475 6271 2517 6280
rect 2476 5648 2516 5657
rect 2380 5608 2476 5648
rect 2283 5144 2325 5153
rect 2283 5104 2284 5144
rect 2324 5104 2325 5144
rect 2283 5095 2325 5104
rect 2476 5069 2516 5608
rect 2475 5060 2517 5069
rect 2475 5020 2476 5060
rect 2516 5020 2517 5060
rect 2475 5011 2517 5020
rect 2092 4768 2228 4808
rect 2092 3380 2132 4768
rect 2475 4136 2517 4145
rect 2475 4096 2476 4136
rect 2516 4096 2517 4136
rect 2475 4087 2517 4096
rect 2476 4002 2516 4087
rect 2187 3800 2229 3809
rect 2187 3760 2188 3800
rect 2228 3760 2229 3800
rect 2187 3751 2229 3760
rect 2092 3331 2132 3340
rect 2188 2876 2228 3751
rect 2475 3632 2517 3641
rect 2475 3592 2476 3632
rect 2516 3592 2517 3632
rect 2475 3583 2517 3592
rect 2283 3464 2325 3473
rect 2283 3424 2284 3464
rect 2324 3424 2325 3464
rect 2283 3415 2325 3424
rect 2284 3296 2324 3415
rect 2476 3380 2516 3583
rect 2476 3331 2516 3340
rect 2284 3247 2324 3256
rect 2379 3128 2421 3137
rect 2379 3088 2380 3128
rect 2420 3088 2421 3128
rect 2379 3079 2421 3088
rect 2284 2876 2324 2885
rect 2188 2836 2284 2876
rect 2284 2827 2324 2836
rect 2092 2708 2132 2717
rect 1996 2668 2092 2708
rect 2092 2659 2132 2668
rect 2380 2549 2420 3079
rect 2475 2708 2517 2717
rect 2475 2668 2476 2708
rect 2516 2668 2517 2708
rect 2475 2659 2517 2668
rect 2476 2574 2516 2659
rect 1995 2540 2037 2549
rect 1995 2500 1996 2540
rect 2036 2500 2037 2540
rect 1995 2491 2037 2500
rect 2379 2540 2421 2549
rect 2379 2500 2380 2540
rect 2420 2500 2421 2540
rect 2572 2540 2612 10051
rect 2667 9176 2709 9185
rect 2667 9136 2668 9176
rect 2708 9136 2709 9176
rect 2667 9127 2709 9136
rect 2668 8840 2708 9127
rect 2668 8791 2708 8800
rect 2764 8597 2804 10144
rect 2860 10109 2900 10228
rect 3244 10184 3284 10193
rect 2859 10100 2901 10109
rect 2859 10060 2860 10100
rect 2900 10060 2901 10100
rect 2859 10051 2901 10060
rect 2956 10100 2996 10109
rect 3244 10100 3284 10144
rect 2996 10060 3284 10100
rect 3340 10184 3380 11320
rect 3532 11033 3572 11647
rect 3531 11024 3573 11033
rect 3531 10984 3532 11024
rect 3572 10984 3573 11024
rect 3531 10975 3573 10984
rect 3724 10781 3764 11656
rect 3915 11612 3957 11621
rect 3915 11572 3916 11612
rect 3956 11572 3957 11612
rect 3915 11563 3957 11572
rect 3916 11024 3956 11563
rect 3916 10975 3956 10984
rect 3723 10772 3765 10781
rect 3723 10732 3724 10772
rect 3764 10732 3765 10772
rect 3723 10723 3765 10732
rect 4203 10772 4245 10781
rect 4203 10732 4204 10772
rect 4244 10732 4245 10772
rect 4203 10723 4245 10732
rect 3688 10604 4056 10613
rect 3728 10564 3770 10604
rect 3810 10564 3852 10604
rect 3892 10564 3934 10604
rect 3974 10564 4016 10604
rect 3688 10555 4056 10564
rect 4204 10445 4244 10723
rect 3915 10436 3957 10445
rect 3915 10396 3916 10436
rect 3956 10396 3957 10436
rect 3915 10387 3957 10396
rect 4203 10436 4245 10445
rect 4203 10396 4204 10436
rect 4244 10396 4245 10436
rect 4203 10387 4245 10396
rect 3531 10352 3573 10361
rect 3531 10312 3532 10352
rect 3572 10312 3573 10352
rect 3531 10303 3573 10312
rect 2956 10051 2996 10060
rect 3340 9848 3380 10144
rect 3244 9808 3380 9848
rect 2859 9596 2901 9605
rect 2859 9556 2860 9596
rect 2900 9556 2901 9596
rect 2859 9547 2901 9556
rect 2860 8756 2900 9547
rect 3051 9512 3093 9521
rect 3148 9512 3188 9521
rect 3051 9472 3052 9512
rect 3092 9472 3148 9512
rect 3051 9463 3093 9472
rect 3148 9463 3188 9472
rect 2860 8707 2900 8716
rect 2763 8588 2805 8597
rect 2763 8548 2764 8588
rect 2804 8548 2805 8588
rect 2763 8539 2805 8548
rect 2764 7589 2804 8539
rect 3052 7841 3092 9463
rect 3147 9344 3189 9353
rect 3147 9304 3148 9344
rect 3188 9304 3189 9344
rect 3147 9295 3189 9304
rect 3051 7832 3093 7841
rect 3051 7792 3052 7832
rect 3092 7792 3093 7832
rect 3051 7783 3093 7792
rect 2763 7580 2805 7589
rect 2763 7540 2764 7580
rect 2804 7540 2805 7580
rect 2763 7531 2805 7540
rect 2859 6992 2901 7001
rect 2859 6952 2860 6992
rect 2900 6952 2901 6992
rect 2859 6943 2901 6952
rect 2667 6572 2709 6581
rect 2667 6532 2668 6572
rect 2708 6532 2709 6572
rect 2667 6523 2709 6532
rect 2668 6438 2708 6523
rect 2763 6488 2805 6497
rect 2763 6448 2764 6488
rect 2804 6448 2805 6488
rect 2763 6439 2805 6448
rect 2860 6483 2900 6943
rect 2955 6740 2997 6749
rect 2955 6700 2956 6740
rect 2996 6700 2997 6740
rect 2955 6691 2997 6700
rect 2668 5900 2708 5909
rect 2764 5900 2804 6439
rect 2860 6434 2900 6443
rect 2708 5860 2804 5900
rect 2860 5900 2900 5909
rect 2956 5900 2996 6691
rect 2900 5860 2996 5900
rect 2668 5851 2708 5860
rect 2860 5851 2900 5860
rect 3052 5732 3092 5741
rect 3052 4985 3092 5692
rect 3051 4976 3093 4985
rect 3051 4936 3052 4976
rect 3092 4936 3093 4976
rect 3051 4927 3093 4936
rect 3051 4808 3093 4817
rect 3051 4768 3052 4808
rect 3092 4768 3093 4808
rect 3051 4759 3093 4768
rect 3052 4313 3092 4759
rect 3051 4304 3093 4313
rect 3051 4264 3052 4304
rect 3092 4264 3093 4304
rect 3051 4255 3093 4264
rect 3148 4229 3188 9295
rect 3244 8261 3284 9808
rect 3340 9680 3380 9689
rect 3380 9640 3476 9680
rect 3340 9631 3380 9640
rect 3436 9521 3476 9640
rect 3435 9512 3477 9521
rect 3435 9472 3436 9512
rect 3476 9472 3477 9512
rect 3435 9463 3477 9472
rect 3532 8672 3572 10303
rect 3819 10268 3861 10277
rect 3819 10228 3820 10268
rect 3860 10228 3861 10268
rect 3819 10219 3861 10228
rect 3724 10184 3764 10195
rect 3724 10109 3764 10144
rect 3820 10134 3860 10219
rect 3723 10100 3765 10109
rect 3723 10060 3724 10100
rect 3764 10060 3765 10100
rect 3723 10051 3765 10060
rect 3723 9512 3765 9521
rect 3723 9472 3724 9512
rect 3764 9472 3765 9512
rect 3723 9463 3765 9472
rect 3820 9512 3860 9521
rect 3916 9512 3956 10387
rect 4204 10268 4244 10387
rect 4300 10352 4340 13168
rect 4395 13208 4437 13217
rect 4395 13168 4396 13208
rect 4436 13168 4437 13208
rect 4395 13159 4437 13168
rect 4396 13074 4436 13159
rect 4491 12536 4533 12545
rect 4491 12496 4492 12536
rect 4532 12496 4533 12536
rect 4491 12487 4533 12496
rect 4395 11528 4437 11537
rect 4395 11488 4396 11528
rect 4436 11488 4437 11528
rect 4395 11479 4437 11488
rect 4396 11394 4436 11479
rect 4492 10697 4532 12487
rect 4491 10688 4533 10697
rect 4491 10648 4492 10688
rect 4532 10648 4533 10688
rect 4491 10639 4533 10648
rect 4588 10352 4628 16990
rect 4972 16409 5012 17032
rect 5356 17072 5396 18031
rect 5452 17744 5492 20392
rect 5548 20105 5588 20560
rect 5740 20560 5876 20600
rect 5932 20980 6068 21020
rect 5932 20596 5972 20980
rect 6027 20852 6069 20861
rect 6027 20812 6028 20852
rect 6068 20812 6069 20852
rect 6027 20803 6069 20812
rect 6028 20768 6068 20803
rect 6028 20717 6068 20728
rect 6124 20768 6164 21391
rect 6124 20719 6164 20728
rect 6220 20600 6260 22912
rect 6316 22709 6356 28960
rect 6507 28960 6508 29000
rect 6548 28960 6549 29000
rect 6507 28951 6549 28960
rect 6603 28916 6645 28925
rect 6603 28876 6604 28916
rect 6644 28876 6645 28916
rect 6603 28867 6645 28876
rect 6604 27161 6644 28867
rect 6700 27656 6740 29455
rect 6700 27329 6740 27616
rect 6699 27320 6741 27329
rect 6699 27280 6700 27320
rect 6740 27280 6741 27320
rect 6699 27271 6741 27280
rect 6603 27152 6645 27161
rect 6603 27112 6604 27152
rect 6644 27112 6645 27152
rect 6796 27152 6836 35596
rect 6892 34880 6932 36436
rect 6988 35057 7028 36604
rect 6987 35048 7029 35057
rect 6987 35008 6988 35048
rect 7028 35008 7029 35048
rect 6987 34999 7029 35008
rect 6892 34840 7028 34880
rect 6988 33125 7028 34840
rect 6987 33116 7029 33125
rect 6987 33076 6988 33116
rect 7028 33076 7029 33116
rect 6987 33067 7029 33076
rect 6988 32864 7028 32873
rect 7084 32864 7124 36856
rect 7180 36737 7220 37444
rect 7179 36728 7221 36737
rect 7179 36688 7180 36728
rect 7220 36688 7221 36728
rect 7179 36679 7221 36688
rect 7276 35384 7316 39787
rect 7372 39752 7412 40879
rect 7660 40433 7700 40464
rect 7659 40424 7701 40433
rect 7659 40384 7660 40424
rect 7700 40384 7701 40424
rect 7659 40375 7701 40384
rect 7467 40340 7509 40349
rect 7467 40300 7468 40340
rect 7508 40300 7509 40340
rect 7467 40291 7509 40300
rect 7660 40340 7700 40375
rect 7468 40206 7508 40291
rect 7467 40088 7509 40097
rect 7467 40048 7468 40088
rect 7508 40048 7509 40088
rect 7467 40039 7509 40048
rect 7372 39703 7412 39712
rect 7468 38921 7508 40039
rect 7467 38912 7509 38921
rect 7467 38872 7468 38912
rect 7508 38872 7509 38912
rect 7467 38863 7509 38872
rect 7660 38408 7700 40300
rect 7468 38368 7700 38408
rect 7468 38165 7508 38368
rect 7563 38240 7605 38249
rect 7563 38200 7564 38240
rect 7604 38200 7605 38240
rect 7563 38191 7605 38200
rect 7660 38240 7700 38249
rect 7467 38156 7509 38165
rect 7467 38116 7468 38156
rect 7508 38116 7509 38156
rect 7467 38107 7509 38116
rect 7372 37400 7412 37409
rect 7372 36905 7412 37360
rect 7467 37232 7509 37241
rect 7467 37192 7468 37232
rect 7508 37192 7509 37232
rect 7467 37183 7509 37192
rect 7468 37098 7508 37183
rect 7371 36896 7413 36905
rect 7371 36856 7372 36896
rect 7412 36856 7413 36896
rect 7371 36847 7413 36856
rect 7372 35468 7412 36847
rect 7468 36728 7508 36737
rect 7468 36569 7508 36688
rect 7467 36560 7509 36569
rect 7467 36520 7468 36560
rect 7508 36520 7509 36560
rect 7467 36511 7509 36520
rect 7564 36401 7604 38191
rect 7660 37829 7700 38200
rect 7659 37820 7701 37829
rect 7659 37780 7660 37820
rect 7700 37780 7701 37820
rect 7659 37771 7701 37780
rect 7756 37661 7796 40972
rect 7948 40963 7988 40972
rect 8044 40853 8084 41215
rect 8140 41213 8180 41224
rect 8332 41105 8372 42928
rect 8524 41525 8564 42928
rect 8523 41516 8565 41525
rect 8523 41476 8524 41516
rect 8564 41476 8565 41516
rect 8523 41467 8565 41476
rect 8331 41096 8373 41105
rect 8331 41056 8332 41096
rect 8372 41056 8373 41096
rect 8331 41047 8373 41056
rect 8043 40844 8085 40853
rect 8043 40804 8044 40844
rect 8084 40804 8085 40844
rect 8043 40795 8085 40804
rect 7947 40676 7989 40685
rect 7947 40636 7948 40676
rect 7988 40636 7989 40676
rect 7947 40627 7989 40636
rect 7948 40542 7988 40627
rect 8332 40552 8564 40592
rect 8139 40508 8181 40517
rect 8139 40468 8140 40508
rect 8180 40468 8181 40508
rect 8139 40459 8181 40468
rect 8140 40374 8180 40459
rect 7851 40340 7893 40349
rect 7851 40300 7852 40340
rect 7892 40300 7893 40340
rect 7851 40291 7893 40300
rect 7852 39747 7892 40291
rect 8235 40004 8277 40013
rect 8235 39964 8236 40004
rect 8276 39964 8277 40004
rect 8235 39955 8277 39964
rect 8236 39920 8276 39955
rect 8236 39869 8276 39880
rect 8044 39836 8084 39847
rect 8044 39761 8084 39796
rect 7852 39698 7892 39707
rect 8043 39752 8085 39761
rect 8043 39712 8044 39752
rect 8084 39712 8085 39752
rect 8043 39703 8085 39712
rect 8332 38837 8372 40552
rect 8428 40424 8468 40433
rect 8428 39080 8468 40384
rect 8524 40424 8564 40552
rect 8524 40375 8564 40384
rect 8523 40172 8565 40181
rect 8523 40132 8524 40172
rect 8564 40132 8565 40172
rect 8523 40123 8565 40132
rect 8524 39752 8564 40123
rect 8524 39425 8564 39712
rect 8523 39416 8565 39425
rect 8523 39376 8524 39416
rect 8564 39376 8565 39416
rect 8523 39367 8565 39376
rect 8620 39080 8660 39089
rect 8428 39040 8620 39080
rect 8620 39031 8660 39040
rect 8427 38912 8469 38921
rect 8427 38872 8428 38912
rect 8468 38872 8469 38912
rect 8427 38863 8469 38872
rect 8331 38828 8373 38837
rect 8331 38788 8332 38828
rect 8372 38788 8373 38828
rect 8331 38779 8373 38788
rect 8043 38408 8085 38417
rect 8043 38368 8044 38408
rect 8084 38368 8085 38408
rect 8043 38359 8085 38368
rect 8044 38274 8084 38359
rect 8332 38072 8372 38081
rect 7852 37988 7892 37997
rect 7755 37652 7797 37661
rect 7755 37612 7756 37652
rect 7796 37612 7797 37652
rect 7755 37603 7797 37612
rect 7852 37409 7892 37948
rect 8043 37736 8085 37745
rect 8043 37696 8044 37736
rect 8084 37696 8085 37736
rect 8043 37687 8085 37696
rect 8044 37493 8084 37687
rect 8332 37493 8372 38032
rect 8428 37829 8468 38863
rect 8523 38408 8565 38417
rect 8523 38368 8524 38408
rect 8564 38368 8565 38408
rect 8523 38359 8565 38368
rect 8427 37820 8469 37829
rect 8427 37780 8428 37820
rect 8468 37780 8469 37820
rect 8427 37771 8469 37780
rect 8043 37484 8085 37493
rect 8043 37444 8044 37484
rect 8084 37444 8085 37484
rect 8043 37435 8085 37444
rect 8331 37484 8373 37493
rect 8331 37444 8332 37484
rect 8372 37444 8373 37484
rect 8331 37435 8373 37444
rect 7660 37400 7700 37409
rect 7660 36737 7700 37360
rect 7851 37400 7893 37409
rect 7851 37360 7852 37400
rect 7892 37360 7893 37400
rect 7851 37351 7893 37360
rect 7948 37400 7988 37409
rect 7852 37232 7892 37241
rect 7756 37192 7852 37232
rect 7659 36728 7701 36737
rect 7659 36688 7660 36728
rect 7700 36688 7701 36728
rect 7659 36679 7701 36688
rect 7563 36392 7605 36401
rect 7563 36352 7564 36392
rect 7604 36352 7605 36392
rect 7563 36343 7605 36352
rect 7372 35428 7508 35468
rect 7468 35384 7508 35428
rect 7276 35344 7412 35384
rect 7276 35216 7316 35225
rect 7180 35176 7276 35216
rect 7180 34637 7220 35176
rect 7276 35167 7316 35176
rect 7179 34628 7221 34637
rect 7179 34588 7180 34628
rect 7220 34588 7221 34628
rect 7179 34579 7221 34588
rect 7180 34049 7220 34579
rect 7179 34040 7221 34049
rect 7179 34000 7180 34040
rect 7220 34000 7221 34040
rect 7179 33991 7221 34000
rect 7028 32824 7124 32864
rect 7180 33704 7220 33991
rect 6988 28505 7028 32824
rect 7083 31772 7125 31781
rect 7083 31732 7084 31772
rect 7124 31732 7125 31772
rect 7083 31723 7125 31732
rect 7084 31520 7124 31723
rect 7083 31480 7124 31520
rect 7083 31361 7123 31480
rect 7083 31352 7124 31361
rect 7083 31321 7084 31352
rect 7084 31303 7124 31312
rect 7083 29420 7125 29429
rect 7083 29380 7084 29420
rect 7124 29380 7125 29420
rect 7083 29371 7125 29380
rect 7084 28580 7124 29371
rect 7180 28925 7220 33664
rect 7372 33620 7412 35344
rect 7468 35309 7508 35344
rect 7467 35300 7509 35309
rect 7467 35260 7468 35300
rect 7508 35260 7604 35300
rect 7467 35251 7509 35260
rect 7468 35220 7508 35251
rect 7564 34469 7604 35260
rect 7660 35225 7700 36679
rect 7756 35981 7796 37192
rect 7852 37183 7892 37192
rect 7948 36989 7988 37360
rect 8140 37232 8180 37241
rect 8044 37192 8140 37232
rect 7947 36980 7989 36989
rect 7947 36940 7948 36980
rect 7988 36940 7989 36980
rect 7947 36931 7989 36940
rect 8044 36812 8084 37192
rect 8140 37183 8180 37192
rect 8332 36896 8372 37435
rect 8427 37400 8469 37409
rect 8427 37360 8428 37400
rect 8468 37360 8469 37400
rect 8427 37351 8469 37360
rect 8524 37400 8564 38359
rect 8619 38240 8661 38249
rect 8619 38200 8620 38240
rect 8660 38200 8661 38240
rect 8619 38191 8661 38200
rect 8620 38106 8660 38191
rect 8524 37351 8564 37360
rect 8428 37266 8468 37351
rect 8332 36847 8372 36856
rect 8619 36896 8661 36905
rect 8619 36856 8620 36896
rect 8660 36856 8661 36896
rect 8619 36847 8661 36856
rect 7852 36772 8084 36812
rect 8140 36812 8180 36821
rect 7755 35972 7797 35981
rect 7755 35932 7756 35972
rect 7796 35932 7797 35972
rect 7755 35923 7797 35932
rect 7659 35216 7701 35225
rect 7659 35176 7660 35216
rect 7700 35176 7701 35216
rect 7659 35167 7701 35176
rect 7756 35141 7796 35923
rect 7755 35132 7797 35141
rect 7755 35092 7756 35132
rect 7796 35092 7797 35132
rect 7755 35083 7797 35092
rect 7659 34964 7701 34973
rect 7659 34924 7660 34964
rect 7700 34924 7701 34964
rect 7659 34915 7701 34924
rect 7660 34721 7700 34915
rect 7659 34712 7701 34721
rect 7659 34672 7660 34712
rect 7700 34672 7701 34712
rect 7659 34663 7701 34672
rect 7755 34628 7797 34637
rect 7755 34588 7756 34628
rect 7796 34588 7797 34628
rect 7755 34579 7797 34588
rect 7563 34460 7605 34469
rect 7563 34420 7564 34460
rect 7604 34420 7605 34460
rect 7563 34411 7605 34420
rect 7564 33713 7604 34411
rect 7756 34376 7796 34579
rect 7756 34327 7796 34336
rect 7852 33965 7892 36772
rect 8140 36728 8180 36772
rect 8620 36728 8660 36847
rect 7996 36686 8036 36695
rect 8140 36688 8564 36728
rect 7996 36644 8036 36646
rect 7996 36604 8084 36644
rect 8044 36140 8084 36604
rect 8428 36560 8468 36569
rect 8236 36140 8276 36149
rect 8044 36100 8236 36140
rect 8236 36091 8276 36100
rect 8428 36056 8468 36520
rect 8428 36007 8468 36016
rect 8044 35888 8084 35897
rect 8524 35888 8564 36688
rect 8620 36679 8660 36688
rect 8044 35729 8084 35848
rect 8428 35848 8564 35888
rect 8043 35720 8085 35729
rect 8043 35680 8044 35720
rect 8084 35680 8085 35720
rect 8043 35671 8085 35680
rect 8428 35393 8468 35848
rect 8524 35720 8564 35729
rect 8427 35384 8469 35393
rect 8427 35344 8428 35384
rect 8468 35344 8469 35384
rect 8427 35335 8469 35344
rect 8043 35300 8085 35309
rect 8043 35260 8044 35300
rect 8084 35260 8085 35300
rect 8043 35251 8085 35260
rect 7947 35216 7989 35225
rect 7947 35176 7948 35216
rect 7988 35176 7989 35216
rect 7947 35167 7989 35176
rect 7948 34301 7988 35167
rect 8044 35166 8084 35251
rect 8140 35216 8180 35225
rect 8043 35048 8085 35057
rect 8043 35008 8044 35048
rect 8084 35008 8085 35048
rect 8043 34999 8085 35008
rect 7947 34292 7989 34301
rect 7947 34252 7948 34292
rect 7988 34252 7989 34292
rect 7947 34243 7989 34252
rect 8044 34124 8084 34999
rect 8140 34637 8180 35176
rect 8236 35216 8276 35225
rect 8236 35048 8276 35176
rect 8428 35048 8468 35057
rect 8236 35008 8428 35048
rect 8428 34999 8468 35008
rect 8524 34973 8564 35680
rect 8716 35468 8756 42928
rect 8908 42197 8948 42928
rect 8907 42188 8949 42197
rect 8907 42148 8908 42188
rect 8948 42148 8949 42188
rect 8907 42139 8949 42148
rect 8908 40433 8948 40518
rect 9003 40508 9045 40517
rect 9003 40468 9004 40508
rect 9044 40468 9045 40508
rect 9003 40459 9045 40468
rect 8907 40424 8949 40433
rect 8907 40384 8908 40424
rect 8948 40384 8949 40424
rect 8907 40375 8949 40384
rect 9004 40374 9044 40459
rect 8907 40256 8949 40265
rect 8907 40216 8908 40256
rect 8948 40216 8949 40256
rect 8907 40207 8949 40216
rect 8811 38996 8853 39005
rect 8811 38956 8812 38996
rect 8852 38956 8853 38996
rect 8811 38947 8853 38956
rect 8812 38912 8852 38947
rect 8812 38669 8852 38872
rect 8811 38660 8853 38669
rect 8811 38620 8812 38660
rect 8852 38620 8853 38660
rect 8811 38611 8853 38620
rect 8908 37400 8948 40207
rect 9100 38165 9140 42928
rect 9292 42281 9332 42928
rect 9291 42272 9333 42281
rect 9291 42232 9292 42272
rect 9332 42232 9333 42272
rect 9291 42223 9333 42232
rect 9291 42104 9333 42113
rect 9291 42064 9292 42104
rect 9332 42064 9333 42104
rect 9291 42055 9333 42064
rect 9195 42020 9237 42029
rect 9195 41980 9196 42020
rect 9236 41980 9237 42020
rect 9195 41971 9237 41980
rect 9196 40013 9236 41971
rect 9292 41189 9332 42055
rect 9484 41609 9524 42928
rect 9579 42608 9621 42617
rect 9579 42568 9580 42608
rect 9620 42568 9621 42608
rect 9579 42559 9621 42568
rect 9483 41600 9525 41609
rect 9483 41560 9484 41600
rect 9524 41560 9525 41600
rect 9483 41551 9525 41560
rect 9387 41432 9429 41441
rect 9580 41432 9620 42559
rect 9387 41392 9388 41432
rect 9428 41392 9429 41432
rect 9387 41383 9429 41392
rect 9484 41392 9620 41432
rect 9388 41273 9428 41383
rect 9387 41264 9429 41273
rect 9387 41224 9388 41264
rect 9428 41224 9429 41264
rect 9387 41215 9429 41224
rect 9291 41180 9333 41189
rect 9291 41140 9292 41180
rect 9332 41140 9333 41180
rect 9291 41131 9333 41140
rect 9388 41130 9428 41215
rect 9484 40424 9524 41392
rect 9579 41180 9621 41189
rect 9579 41140 9580 41180
rect 9620 41140 9621 41180
rect 9579 41131 9621 41140
rect 9580 41096 9620 41131
rect 9580 41045 9620 41056
rect 9484 40375 9524 40384
rect 9676 40256 9716 42928
rect 9388 40216 9716 40256
rect 9772 41180 9812 41189
rect 9195 40004 9237 40013
rect 9195 39964 9196 40004
rect 9236 39964 9237 40004
rect 9195 39955 9237 39964
rect 9099 38156 9141 38165
rect 9099 38116 9100 38156
rect 9140 38116 9141 38156
rect 9099 38107 9141 38116
rect 9388 37820 9428 40216
rect 9483 40004 9525 40013
rect 9483 39964 9484 40004
rect 9524 39964 9525 40004
rect 9483 39955 9525 39964
rect 9196 37780 9428 37820
rect 9003 37484 9045 37493
rect 9003 37444 9004 37484
rect 9044 37444 9045 37484
rect 9003 37435 9045 37444
rect 8620 35428 8756 35468
rect 8812 37360 8908 37400
rect 8523 34964 8565 34973
rect 8523 34924 8524 34964
rect 8564 34924 8565 34964
rect 8523 34915 8565 34924
rect 8139 34628 8181 34637
rect 8139 34588 8140 34628
rect 8180 34588 8181 34628
rect 8139 34579 8181 34588
rect 8331 34376 8373 34385
rect 8331 34336 8332 34376
rect 8372 34336 8373 34376
rect 8331 34327 8373 34336
rect 7948 34084 8084 34124
rect 8139 34124 8181 34133
rect 8139 34084 8140 34124
rect 8180 34084 8181 34124
rect 7851 33956 7893 33965
rect 7851 33916 7852 33956
rect 7892 33916 7893 33956
rect 7851 33907 7893 33916
rect 7852 33713 7892 33798
rect 7563 33704 7605 33713
rect 7563 33664 7564 33704
rect 7604 33664 7605 33704
rect 7851 33704 7893 33713
rect 7563 33655 7605 33664
rect 7660 33691 7700 33700
rect 7851 33664 7852 33704
rect 7892 33664 7893 33704
rect 7851 33655 7893 33664
rect 7660 33629 7700 33651
rect 7659 33620 7701 33629
rect 7372 33580 7508 33620
rect 7371 33452 7413 33461
rect 7371 33412 7372 33452
rect 7412 33412 7413 33452
rect 7371 33403 7413 33412
rect 7372 33318 7412 33403
rect 7371 33116 7413 33125
rect 7371 33076 7372 33116
rect 7412 33076 7413 33116
rect 7371 33067 7413 33076
rect 7372 31025 7412 33067
rect 7371 31016 7413 31025
rect 7371 30976 7372 31016
rect 7412 30976 7413 31016
rect 7371 30967 7413 30976
rect 7468 30269 7508 33580
rect 7659 33580 7660 33620
rect 7700 33580 7701 33620
rect 7659 33571 7701 33580
rect 7948 33620 7988 34084
rect 8139 34075 8181 34084
rect 7948 33571 7988 33580
rect 8140 33620 8180 34075
rect 8236 33713 8276 33798
rect 8235 33704 8277 33713
rect 8235 33664 8236 33704
rect 8276 33664 8277 33704
rect 8235 33655 8277 33664
rect 7660 33556 7700 33571
rect 8043 33536 8085 33545
rect 8043 33496 8044 33536
rect 8084 33496 8085 33536
rect 8043 33487 8085 33496
rect 7564 33452 7604 33461
rect 7564 32873 7604 33412
rect 7947 33452 7989 33461
rect 7947 33412 7948 33452
rect 7988 33412 7989 33452
rect 7947 33403 7989 33412
rect 7948 32957 7988 33403
rect 8044 33402 8084 33487
rect 8140 33452 8180 33580
rect 8140 33412 8276 33452
rect 8139 33284 8181 33293
rect 8139 33244 8140 33284
rect 8180 33244 8181 33284
rect 8139 33235 8181 33244
rect 7947 32948 7989 32957
rect 7947 32908 7948 32948
rect 7988 32908 8084 32948
rect 7947 32899 7989 32908
rect 7563 32864 7605 32873
rect 7563 32824 7564 32864
rect 7604 32824 7605 32864
rect 7563 32815 7605 32824
rect 7563 32444 7605 32453
rect 7563 32404 7564 32444
rect 7604 32404 7605 32444
rect 7563 32395 7605 32404
rect 7564 32192 7604 32395
rect 7564 31529 7604 32152
rect 7948 32192 7988 32201
rect 7756 31940 7796 31949
rect 7660 31900 7756 31940
rect 7563 31520 7605 31529
rect 7563 31480 7564 31520
rect 7604 31480 7605 31520
rect 7563 31471 7605 31480
rect 7564 31357 7604 31366
rect 7660 31352 7700 31900
rect 7756 31891 7796 31900
rect 7948 31613 7988 32152
rect 8044 32192 8084 32908
rect 8140 32360 8180 33235
rect 8236 33032 8276 33412
rect 8332 33293 8372 34327
rect 8524 34217 8564 34915
rect 8620 34544 8660 35428
rect 8812 35393 8852 37360
rect 8908 37351 8948 37360
rect 9004 37350 9044 37435
rect 9099 37232 9141 37241
rect 9099 37192 9100 37232
rect 9140 37192 9141 37232
rect 9099 37183 9141 37192
rect 8908 36737 8948 36822
rect 8907 36728 8949 36737
rect 8907 36688 8908 36728
rect 8948 36688 8949 36728
rect 8907 36679 8949 36688
rect 8908 36476 8948 36485
rect 8811 35384 8853 35393
rect 8811 35344 8812 35384
rect 8852 35344 8853 35384
rect 8811 35335 8853 35344
rect 8811 35216 8853 35225
rect 8716 35174 8756 35183
rect 8811 35176 8812 35216
rect 8852 35176 8853 35216
rect 8811 35167 8853 35176
rect 8716 34973 8756 35134
rect 8812 35082 8852 35167
rect 8715 34964 8757 34973
rect 8715 34924 8716 34964
rect 8756 34924 8757 34964
rect 8715 34915 8757 34924
rect 8908 34880 8948 36436
rect 9003 36476 9045 36485
rect 9003 36436 9004 36476
rect 9044 36436 9045 36476
rect 9003 36427 9045 36436
rect 9004 35888 9044 36427
rect 9100 35972 9140 37183
rect 9196 36233 9236 37780
rect 9484 37400 9524 39955
rect 9772 39929 9812 41140
rect 9868 40265 9908 42928
rect 9963 41936 10005 41945
rect 9963 41896 9964 41936
rect 10004 41896 10005 41936
rect 9963 41887 10005 41896
rect 9964 41432 10004 41887
rect 9964 41383 10004 41392
rect 9964 40429 10004 40438
rect 10060 40433 10100 42928
rect 10155 41180 10197 41189
rect 10155 41140 10156 41180
rect 10196 41140 10197 41180
rect 10155 41131 10197 41140
rect 10156 41046 10196 41131
rect 9867 40256 9909 40265
rect 9867 40216 9868 40256
rect 9908 40216 9909 40256
rect 9867 40207 9909 40216
rect 9771 39920 9813 39929
rect 9771 39880 9772 39920
rect 9812 39880 9813 39920
rect 9771 39871 9813 39880
rect 9964 39920 10004 40389
rect 10059 40424 10101 40433
rect 10059 40384 10060 40424
rect 10100 40384 10101 40424
rect 10059 40375 10101 40384
rect 9964 39871 10004 39880
rect 10156 40256 10196 40265
rect 10252 40256 10292 42928
rect 10347 41852 10389 41861
rect 10347 41812 10348 41852
rect 10388 41812 10389 41852
rect 10347 41803 10389 41812
rect 10348 41432 10388 41803
rect 10444 41609 10484 42928
rect 10443 41600 10485 41609
rect 10443 41560 10444 41600
rect 10484 41560 10485 41600
rect 10443 41551 10485 41560
rect 10348 41383 10388 41392
rect 10540 41180 10580 41189
rect 10444 41140 10540 41180
rect 10347 40592 10389 40601
rect 10347 40552 10348 40592
rect 10388 40552 10389 40592
rect 10347 40543 10389 40552
rect 10348 40424 10388 40543
rect 10348 40375 10388 40384
rect 10252 40216 10388 40256
rect 9772 39752 9812 39761
rect 9812 39712 9908 39752
rect 9772 39703 9812 39712
rect 9868 38921 9908 39712
rect 9867 38912 9909 38921
rect 9867 38872 9868 38912
rect 9908 38872 9909 38912
rect 9867 38863 9909 38872
rect 10060 38912 10100 38921
rect 9868 38585 9908 38863
rect 10060 38585 10100 38872
rect 9867 38576 9909 38585
rect 9867 38536 9868 38576
rect 9908 38536 9909 38576
rect 9867 38527 9909 38536
rect 10059 38576 10101 38585
rect 10059 38536 10060 38576
rect 10100 38536 10101 38576
rect 10059 38527 10101 38536
rect 9868 38240 9908 38527
rect 9868 38191 9908 38200
rect 10060 37988 10100 37997
rect 9964 37948 10060 37988
rect 9964 37414 10004 37948
rect 10060 37939 10100 37948
rect 10156 37820 10196 40216
rect 10251 40088 10293 40097
rect 10251 40048 10252 40088
rect 10292 40048 10293 40088
rect 10251 40039 10293 40048
rect 10252 39752 10292 40039
rect 10252 39703 10292 39712
rect 10251 38828 10293 38837
rect 10251 38788 10252 38828
rect 10292 38788 10293 38828
rect 10251 38779 10293 38788
rect 10252 38694 10292 38779
rect 10156 37780 10292 37820
rect 9964 37365 10004 37374
rect 9484 37064 9524 37360
rect 10156 37232 10196 37241
rect 9292 37024 9524 37064
rect 10060 37192 10156 37232
rect 9195 36224 9237 36233
rect 9195 36184 9196 36224
rect 9236 36184 9237 36224
rect 9195 36175 9237 36184
rect 9100 35923 9140 35932
rect 9196 36056 9236 36065
rect 9004 35729 9044 35848
rect 9003 35720 9045 35729
rect 9003 35680 9004 35720
rect 9044 35680 9045 35720
rect 9003 35671 9045 35680
rect 9100 35216 9140 35225
rect 9100 35141 9140 35176
rect 9099 35132 9141 35141
rect 9099 35092 9100 35132
rect 9140 35092 9141 35132
rect 9099 35083 9141 35092
rect 8812 34840 8948 34880
rect 8620 34504 8756 34544
rect 8619 34376 8661 34385
rect 8619 34336 8620 34376
rect 8660 34336 8661 34376
rect 8619 34327 8661 34336
rect 8523 34208 8565 34217
rect 8523 34168 8524 34208
rect 8564 34168 8565 34208
rect 8523 34159 8565 34168
rect 8524 34074 8564 34159
rect 8524 33704 8564 33713
rect 8620 33704 8660 34327
rect 8564 33664 8660 33704
rect 8524 33461 8564 33664
rect 8523 33452 8565 33461
rect 8523 33412 8524 33452
rect 8564 33412 8565 33452
rect 8523 33403 8565 33412
rect 8331 33284 8373 33293
rect 8331 33244 8332 33284
rect 8372 33244 8373 33284
rect 8331 33235 8373 33244
rect 8716 33032 8756 34504
rect 8812 34124 8852 34840
rect 9100 34796 9140 35083
rect 8908 34756 9140 34796
rect 8908 34385 8948 34756
rect 9196 34628 9236 36016
rect 9292 35972 9332 37024
rect 9483 36896 9525 36905
rect 9483 36856 9484 36896
rect 9524 36856 9525 36896
rect 9483 36847 9525 36856
rect 9484 36728 9524 36847
rect 9484 36653 9524 36688
rect 9483 36644 9525 36653
rect 9483 36604 9484 36644
rect 9524 36604 9525 36644
rect 9483 36595 9525 36604
rect 9387 36476 9429 36485
rect 9387 36436 9388 36476
rect 9428 36436 9429 36476
rect 9387 36427 9429 36436
rect 9388 36065 9428 36427
rect 10060 36233 10100 37192
rect 10156 37183 10196 37192
rect 10155 36728 10197 36737
rect 10155 36688 10156 36728
rect 10196 36688 10197 36728
rect 10155 36679 10197 36688
rect 10059 36224 10101 36233
rect 10059 36184 10060 36224
rect 10100 36184 10101 36224
rect 10059 36175 10101 36184
rect 9387 36056 9429 36065
rect 9387 36016 9388 36056
rect 9428 36016 9429 36056
rect 9387 36007 9429 36016
rect 9292 35923 9332 35932
rect 9388 35888 9428 35897
rect 9291 35804 9333 35813
rect 9291 35764 9292 35804
rect 9332 35764 9333 35804
rect 9291 35755 9333 35764
rect 9292 35645 9332 35755
rect 9291 35636 9333 35645
rect 9291 35596 9292 35636
rect 9332 35596 9333 35636
rect 9291 35587 9333 35596
rect 9004 34588 9236 34628
rect 9292 34628 9332 35587
rect 9388 35057 9428 35848
rect 9579 35888 9621 35897
rect 9579 35848 9580 35888
rect 9620 35848 9621 35888
rect 9579 35839 9621 35848
rect 9580 35561 9620 35839
rect 10156 35813 10196 36679
rect 10155 35804 10197 35813
rect 10155 35764 10156 35804
rect 10196 35764 10197 35804
rect 10155 35755 10197 35764
rect 10252 35729 10292 37780
rect 10348 36653 10388 40216
rect 10444 39089 10484 41140
rect 10540 41131 10580 41140
rect 10636 39089 10676 42928
rect 10731 40508 10773 40517
rect 10828 40508 10868 42928
rect 10731 40468 10732 40508
rect 10772 40468 10868 40508
rect 10731 40459 10773 40468
rect 10443 39080 10485 39089
rect 10443 39040 10444 39080
rect 10484 39040 10485 39080
rect 10443 39031 10485 39040
rect 10635 39080 10677 39089
rect 10635 39040 10636 39080
rect 10676 39040 10677 39080
rect 10635 39031 10677 39040
rect 10540 38912 10580 38923
rect 10540 38837 10580 38872
rect 10635 38912 10677 38921
rect 10635 38872 10636 38912
rect 10676 38872 10677 38912
rect 10635 38863 10677 38872
rect 10539 38828 10581 38837
rect 10539 38788 10540 38828
rect 10580 38788 10581 38828
rect 10539 38779 10581 38788
rect 10636 38778 10676 38863
rect 10635 38408 10677 38417
rect 10635 38368 10636 38408
rect 10676 38368 10677 38408
rect 10635 38359 10677 38368
rect 10636 38240 10676 38359
rect 10732 38249 10772 40459
rect 10923 40424 10965 40433
rect 10923 40384 10924 40424
rect 10964 40384 10965 40424
rect 10923 40375 10965 40384
rect 10539 37988 10581 37997
rect 10636 37988 10676 38200
rect 10731 38240 10773 38249
rect 10731 38200 10732 38240
rect 10772 38200 10773 38240
rect 10731 38191 10773 38200
rect 10539 37948 10540 37988
rect 10580 37948 10676 37988
rect 10539 37939 10581 37948
rect 10347 36644 10389 36653
rect 10347 36604 10348 36644
rect 10388 36604 10389 36644
rect 10347 36595 10389 36604
rect 10347 36224 10389 36233
rect 10347 36184 10348 36224
rect 10388 36184 10389 36224
rect 10347 36175 10389 36184
rect 10251 35720 10293 35729
rect 10251 35680 10252 35720
rect 10292 35680 10293 35720
rect 10251 35671 10293 35680
rect 10059 35636 10101 35645
rect 10059 35596 10060 35636
rect 10100 35596 10101 35636
rect 10348 35636 10388 36175
rect 10348 35596 10484 35636
rect 10059 35587 10101 35596
rect 9579 35552 9621 35561
rect 9579 35512 9580 35552
rect 9620 35512 9621 35552
rect 9579 35503 9621 35512
rect 10060 35393 10100 35587
rect 10059 35384 10101 35393
rect 10059 35344 10060 35384
rect 10100 35344 10101 35384
rect 10059 35335 10101 35344
rect 10156 35388 10196 35397
rect 9867 35300 9909 35309
rect 9867 35260 9868 35300
rect 9908 35260 9909 35300
rect 9867 35251 9909 35260
rect 9479 35216 9519 35225
rect 9580 35216 9620 35225
rect 9519 35176 9524 35216
rect 9479 35167 9524 35176
rect 9387 35048 9429 35057
rect 9387 35008 9388 35048
rect 9428 35008 9429 35048
rect 9387 34999 9429 35008
rect 9292 34588 9439 34628
rect 9004 34385 9044 34588
rect 8907 34376 8949 34385
rect 8907 34336 8908 34376
rect 8948 34336 8949 34376
rect 9004 34376 9050 34385
rect 9004 34336 9009 34376
rect 9049 34336 9050 34376
rect 8907 34327 8949 34336
rect 9008 34327 9050 34336
rect 9196 34376 9236 34387
rect 8908 34242 8948 34327
rect 9196 34301 9236 34336
rect 9292 34376 9332 34385
rect 9399 34365 9439 34588
rect 9332 34336 9439 34365
rect 9292 34325 9439 34336
rect 9195 34292 9237 34301
rect 9195 34252 9196 34292
rect 9236 34252 9237 34292
rect 9195 34243 9237 34252
rect 9484 34217 9524 35167
rect 9580 34721 9620 35176
rect 9676 35216 9716 35225
rect 9676 34805 9716 35176
rect 9868 35216 9908 35251
rect 9868 35165 9908 35176
rect 9964 35216 10004 35225
rect 10059 35216 10101 35225
rect 10004 35176 10060 35216
rect 10100 35176 10101 35216
rect 9964 35167 10004 35176
rect 10059 35167 10101 35176
rect 9963 34964 10005 34973
rect 9963 34924 9964 34964
rect 10004 34924 10005 34964
rect 9963 34915 10005 34924
rect 9964 34830 10004 34915
rect 9675 34796 9717 34805
rect 9675 34756 9676 34796
rect 9716 34756 9717 34796
rect 9675 34747 9717 34756
rect 9579 34712 9621 34721
rect 9579 34672 9580 34712
rect 9620 34672 9621 34712
rect 9579 34663 9621 34672
rect 9963 34712 10005 34721
rect 9963 34672 9964 34712
rect 10004 34672 10005 34712
rect 9963 34663 10005 34672
rect 9771 34628 9813 34637
rect 9771 34588 9772 34628
rect 9812 34588 9813 34628
rect 9771 34579 9813 34588
rect 9580 34544 9620 34553
rect 9620 34504 9716 34544
rect 9580 34495 9620 34504
rect 9579 34376 9621 34385
rect 9579 34336 9580 34376
rect 9620 34336 9621 34376
rect 9579 34327 9621 34336
rect 9099 34208 9141 34217
rect 9099 34168 9100 34208
rect 9140 34168 9141 34208
rect 9099 34159 9141 34168
rect 9483 34208 9525 34217
rect 9483 34168 9484 34208
rect 9524 34168 9525 34208
rect 9483 34159 9525 34168
rect 8812 34084 9044 34124
rect 8811 33704 8853 33713
rect 8811 33664 8812 33704
rect 8852 33664 8853 33704
rect 8811 33655 8853 33664
rect 8908 33704 8948 33715
rect 8812 33570 8852 33655
rect 8908 33629 8948 33664
rect 8907 33620 8949 33629
rect 8907 33580 8908 33620
rect 8948 33580 8949 33620
rect 8907 33571 8949 33580
rect 8236 32992 8372 33032
rect 8236 32864 8276 32873
rect 8332 32864 8372 32992
rect 8620 32992 8756 33032
rect 8332 32824 8564 32864
rect 8236 32537 8276 32824
rect 8428 32696 8468 32705
rect 8332 32656 8428 32696
rect 8235 32528 8277 32537
rect 8235 32488 8236 32528
rect 8276 32488 8277 32528
rect 8235 32479 8277 32488
rect 8236 32360 8276 32369
rect 8140 32320 8236 32360
rect 8236 32311 8276 32320
rect 8044 32143 8084 32152
rect 7947 31604 7989 31613
rect 7947 31564 7948 31604
rect 7988 31564 7989 31604
rect 7947 31555 7989 31564
rect 7755 31520 7797 31529
rect 7755 31480 7756 31520
rect 7796 31480 7797 31520
rect 7755 31471 7797 31480
rect 7604 31317 7700 31352
rect 7564 31312 7700 31317
rect 7756 31352 7796 31471
rect 8332 31352 8372 32656
rect 8428 32647 8468 32656
rect 8524 31529 8564 32824
rect 8523 31520 8565 31529
rect 8523 31480 8524 31520
rect 8564 31480 8565 31520
rect 8523 31471 8565 31480
rect 7756 31312 7988 31352
rect 7564 31308 7604 31312
rect 7755 31184 7797 31193
rect 7755 31144 7756 31184
rect 7796 31144 7797 31184
rect 7755 31135 7797 31144
rect 7563 31100 7605 31109
rect 7563 31060 7564 31100
rect 7604 31060 7605 31100
rect 7563 31051 7605 31060
rect 7467 30260 7509 30269
rect 7467 30220 7468 30260
rect 7508 30220 7509 30260
rect 7467 30211 7509 30220
rect 7371 29756 7413 29765
rect 7371 29716 7372 29756
rect 7412 29716 7413 29756
rect 7371 29707 7413 29716
rect 7372 29168 7412 29707
rect 7467 29336 7509 29345
rect 7467 29296 7468 29336
rect 7508 29296 7509 29336
rect 7467 29287 7509 29296
rect 7179 28916 7221 28925
rect 7179 28876 7180 28916
rect 7220 28876 7221 28916
rect 7179 28867 7221 28876
rect 7372 28757 7412 29128
rect 7468 29168 7508 29287
rect 7179 28748 7221 28757
rect 7179 28708 7180 28748
rect 7220 28708 7221 28748
rect 7179 28699 7221 28708
rect 7371 28748 7413 28757
rect 7371 28708 7372 28748
rect 7412 28708 7413 28748
rect 7371 28699 7413 28708
rect 7180 28580 7220 28699
rect 7084 28540 7135 28580
rect 6987 28496 7029 28505
rect 6987 28456 6988 28496
rect 7028 28456 7029 28496
rect 6987 28447 7029 28456
rect 7095 28412 7135 28540
rect 7180 28531 7220 28540
rect 6988 28370 7028 28379
rect 7095 28372 7220 28412
rect 6988 28001 7028 28330
rect 7083 28244 7125 28253
rect 7083 28204 7084 28244
rect 7124 28204 7125 28244
rect 7083 28195 7125 28204
rect 6987 27992 7029 28001
rect 6987 27952 6988 27992
rect 7028 27952 7029 27992
rect 6987 27943 7029 27952
rect 6796 27112 6932 27152
rect 6603 27103 6645 27112
rect 6892 26900 6932 27112
rect 6987 26984 7029 26993
rect 6987 26944 6988 26984
rect 7028 26944 7029 26984
rect 7084 26984 7124 28195
rect 7180 27068 7220 28372
rect 7372 28347 7412 28699
rect 7468 28505 7508 29128
rect 7467 28496 7509 28505
rect 7467 28456 7468 28496
rect 7508 28456 7509 28496
rect 7564 28496 7604 31051
rect 7756 31050 7796 31135
rect 7755 30932 7797 30941
rect 7755 30892 7756 30932
rect 7796 30892 7797 30932
rect 7755 30883 7797 30892
rect 7659 29336 7701 29345
rect 7659 29296 7660 29336
rect 7700 29296 7701 29336
rect 7659 29287 7701 29296
rect 7660 29202 7700 29287
rect 7564 28456 7700 28496
rect 7467 28447 7509 28456
rect 7468 28347 7508 28356
rect 7372 28307 7468 28347
rect 7468 28298 7508 28307
rect 7564 28328 7604 28337
rect 7564 28244 7604 28288
rect 7468 28204 7604 28244
rect 7468 28085 7508 28204
rect 7660 28160 7700 28456
rect 7564 28120 7700 28160
rect 7467 28076 7509 28085
rect 7467 28036 7468 28076
rect 7508 28036 7509 28076
rect 7467 28027 7509 28036
rect 7180 27028 7316 27068
rect 7084 26944 7220 26984
rect 6987 26935 7029 26944
rect 6796 26860 6932 26900
rect 6412 26816 6452 26825
rect 6412 26489 6452 26776
rect 6508 26816 6548 26825
rect 6411 26480 6453 26489
rect 6411 26440 6412 26480
rect 6452 26440 6453 26480
rect 6411 26431 6453 26440
rect 6508 25985 6548 26776
rect 6603 26816 6645 26825
rect 6603 26776 6604 26816
rect 6644 26776 6645 26816
rect 6603 26767 6645 26776
rect 6604 26682 6644 26767
rect 6700 26648 6740 26657
rect 6700 26237 6740 26608
rect 6699 26228 6741 26237
rect 6699 26188 6700 26228
rect 6740 26188 6741 26228
rect 6699 26179 6741 26188
rect 6507 25976 6549 25985
rect 6507 25936 6508 25976
rect 6548 25936 6549 25976
rect 6507 25927 6549 25936
rect 6412 25892 6452 25901
rect 6412 24893 6452 25852
rect 6796 25052 6836 26860
rect 6891 26732 6933 26741
rect 6891 26692 6892 26732
rect 6932 26692 6933 26732
rect 6891 26683 6933 26692
rect 6700 25012 6836 25052
rect 6411 24884 6453 24893
rect 6411 24844 6412 24884
rect 6452 24844 6453 24884
rect 6411 24835 6453 24844
rect 6604 24632 6644 24641
rect 6412 24592 6604 24632
rect 6412 23801 6452 24592
rect 6604 24583 6644 24592
rect 6700 24632 6740 25012
rect 6507 24296 6549 24305
rect 6507 24256 6508 24296
rect 6548 24256 6549 24296
rect 6507 24247 6549 24256
rect 6508 23876 6548 24247
rect 6700 24137 6740 24592
rect 6796 24632 6836 24641
rect 6796 24473 6836 24592
rect 6795 24464 6837 24473
rect 6795 24424 6796 24464
rect 6836 24424 6837 24464
rect 6795 24415 6837 24424
rect 6699 24128 6741 24137
rect 6699 24088 6700 24128
rect 6740 24088 6741 24128
rect 6699 24079 6741 24088
rect 6603 23960 6645 23969
rect 6603 23920 6604 23960
rect 6644 23920 6645 23960
rect 6603 23911 6645 23920
rect 6508 23827 6548 23836
rect 6411 23792 6453 23801
rect 6411 23752 6412 23792
rect 6452 23752 6453 23792
rect 6411 23743 6453 23752
rect 6604 23792 6644 23911
rect 6892 23885 6932 26683
rect 6988 24548 7028 26935
rect 7083 26816 7125 26825
rect 7083 26776 7084 26816
rect 7124 26776 7125 26816
rect 7083 26767 7125 26776
rect 7084 26682 7124 26767
rect 7180 26657 7220 26944
rect 7179 26648 7221 26657
rect 7179 26608 7180 26648
rect 7220 26608 7221 26648
rect 7179 26599 7221 26608
rect 7083 26480 7125 26489
rect 7083 26440 7084 26480
rect 7124 26440 7125 26480
rect 7083 26431 7125 26440
rect 7084 24632 7124 26431
rect 7276 25397 7316 27028
rect 7468 26312 7508 28027
rect 7372 26272 7508 26312
rect 7372 26069 7412 26272
rect 7371 26060 7413 26069
rect 7371 26020 7372 26060
rect 7412 26020 7413 26060
rect 7371 26011 7413 26020
rect 7275 25388 7317 25397
rect 7275 25348 7276 25388
rect 7316 25348 7317 25388
rect 7275 25339 7317 25348
rect 7179 25304 7221 25313
rect 7179 25264 7180 25304
rect 7220 25264 7221 25304
rect 7179 25255 7221 25264
rect 7276 25304 7316 25339
rect 7180 25136 7220 25255
rect 7276 25254 7316 25264
rect 7180 25096 7316 25136
rect 7084 24592 7220 24632
rect 6988 24508 7124 24548
rect 6988 24380 7028 24389
rect 6891 23876 6933 23885
rect 6891 23836 6892 23876
rect 6932 23836 6933 23876
rect 6891 23827 6933 23836
rect 6988 23801 7028 24340
rect 6412 23381 6452 23743
rect 6507 23624 6549 23633
rect 6507 23584 6508 23624
rect 6548 23584 6549 23624
rect 6507 23575 6549 23584
rect 6411 23372 6453 23381
rect 6411 23332 6412 23372
rect 6452 23332 6453 23372
rect 6411 23323 6453 23332
rect 6412 23288 6452 23323
rect 6412 23237 6452 23248
rect 6508 22709 6548 23575
rect 6604 23549 6644 23752
rect 6987 23792 7029 23801
rect 6987 23752 6988 23792
rect 7028 23752 7029 23792
rect 6987 23743 7029 23752
rect 7084 23792 7124 24508
rect 6603 23540 6645 23549
rect 6603 23500 6604 23540
rect 6644 23500 6645 23540
rect 6603 23491 6645 23500
rect 6987 23456 7029 23465
rect 6987 23416 6988 23456
rect 7028 23416 7029 23456
rect 6987 23407 7029 23416
rect 6604 23120 6644 23129
rect 6315 22700 6357 22709
rect 6315 22660 6316 22700
rect 6356 22660 6357 22700
rect 6315 22651 6357 22660
rect 6507 22700 6549 22709
rect 6507 22660 6508 22700
rect 6548 22660 6549 22700
rect 6507 22651 6549 22660
rect 6507 22448 6549 22457
rect 6412 22408 6508 22448
rect 6548 22408 6549 22448
rect 5547 20096 5589 20105
rect 5547 20056 5548 20096
rect 5588 20056 5589 20096
rect 5547 20047 5589 20056
rect 5644 19844 5684 19853
rect 5644 19013 5684 19804
rect 5643 19004 5685 19013
rect 5643 18964 5644 19004
rect 5684 18964 5685 19004
rect 5643 18955 5685 18964
rect 5643 18836 5685 18845
rect 5643 18796 5644 18836
rect 5684 18796 5685 18836
rect 5643 18787 5685 18796
rect 5644 18584 5684 18787
rect 5644 18535 5684 18544
rect 5452 17695 5492 17704
rect 5740 17072 5780 20560
rect 5835 20264 5877 20273
rect 5835 20224 5836 20264
rect 5876 20224 5877 20264
rect 5835 20215 5877 20224
rect 5836 20096 5876 20215
rect 5932 20189 5972 20556
rect 6028 20560 6260 20600
rect 6316 22280 6356 22289
rect 6316 21608 6356 22240
rect 5931 20180 5973 20189
rect 5931 20140 5932 20180
rect 5972 20140 5973 20180
rect 5931 20131 5973 20140
rect 5836 20047 5876 20056
rect 5931 19844 5973 19853
rect 5931 19804 5932 19844
rect 5972 19804 5973 19844
rect 5931 19795 5973 19804
rect 5932 19710 5972 19795
rect 5835 19256 5877 19265
rect 5835 19216 5836 19256
rect 5876 19216 5877 19256
rect 5835 19207 5877 19216
rect 5836 19122 5876 19207
rect 5932 17072 5972 17081
rect 5356 17023 5396 17032
rect 5548 17032 5932 17072
rect 5452 16988 5492 16997
rect 5452 16745 5492 16948
rect 5451 16736 5493 16745
rect 5451 16696 5452 16736
rect 5492 16696 5493 16736
rect 5451 16687 5493 16696
rect 4971 16400 5013 16409
rect 4971 16360 4972 16400
rect 5012 16360 5013 16400
rect 4971 16351 5013 16360
rect 5355 16400 5397 16409
rect 5548 16400 5588 17032
rect 5932 17023 5972 17032
rect 6028 16493 6068 20560
rect 6123 20432 6165 20441
rect 6123 20392 6124 20432
rect 6164 20392 6165 20432
rect 6123 20383 6165 20392
rect 6027 16484 6069 16493
rect 6027 16444 6028 16484
rect 6068 16444 6069 16484
rect 6027 16435 6069 16444
rect 5355 16360 5356 16400
rect 5396 16360 5397 16400
rect 5355 16351 5397 16360
rect 5452 16360 5588 16400
rect 4928 15896 5296 15905
rect 4968 15856 5010 15896
rect 5050 15856 5092 15896
rect 5132 15856 5174 15896
rect 5214 15856 5256 15896
rect 4928 15847 5296 15856
rect 5259 15728 5301 15737
rect 5259 15688 5260 15728
rect 5300 15688 5301 15728
rect 5259 15679 5301 15688
rect 5067 15644 5109 15653
rect 5067 15604 5068 15644
rect 5108 15604 5109 15644
rect 5067 15595 5109 15604
rect 5068 15560 5108 15595
rect 5260 15594 5300 15679
rect 5068 15509 5108 15520
rect 5356 15476 5396 16351
rect 5452 15905 5492 16360
rect 5548 16232 5588 16241
rect 5451 15896 5493 15905
rect 5451 15856 5452 15896
rect 5492 15856 5493 15896
rect 5451 15847 5493 15856
rect 5548 15653 5588 16192
rect 5932 16232 5972 16241
rect 5740 16148 5780 16157
rect 5644 16108 5740 16148
rect 5547 15644 5589 15653
rect 5547 15604 5548 15644
rect 5588 15604 5589 15644
rect 5547 15595 5589 15604
rect 5451 15560 5493 15569
rect 5451 15520 5452 15560
rect 5492 15520 5493 15560
rect 5451 15511 5493 15520
rect 5164 15436 5396 15476
rect 5164 15392 5204 15436
rect 5452 15426 5492 15511
rect 5068 15352 5204 15392
rect 5068 14888 5108 15352
rect 5260 15308 5300 15317
rect 4780 14848 5108 14888
rect 5164 15268 5260 15308
rect 4780 14216 4820 14848
rect 5067 14720 5109 14729
rect 5067 14680 5068 14720
rect 5108 14680 5109 14720
rect 5067 14671 5109 14680
rect 5068 14586 5108 14671
rect 5164 14552 5204 15268
rect 5260 15259 5300 15268
rect 5644 15056 5684 16108
rect 5740 16099 5780 16108
rect 5835 16064 5877 16073
rect 5835 16024 5836 16064
rect 5876 16024 5877 16064
rect 5835 16015 5877 16024
rect 5739 15896 5781 15905
rect 5739 15856 5740 15896
rect 5780 15856 5781 15896
rect 5739 15847 5781 15856
rect 5260 15016 5684 15056
rect 5260 14720 5300 15016
rect 5356 14888 5396 14897
rect 5396 14848 5588 14888
rect 5356 14839 5396 14848
rect 5260 14671 5300 14680
rect 5356 14720 5396 14729
rect 5356 14552 5396 14680
rect 5451 14720 5493 14729
rect 5451 14680 5452 14720
rect 5492 14680 5493 14720
rect 5451 14671 5493 14680
rect 5548 14720 5588 14848
rect 5548 14671 5588 14680
rect 5644 14720 5684 15016
rect 5644 14671 5684 14680
rect 5164 14512 5396 14552
rect 4928 14384 5296 14393
rect 4968 14344 5010 14384
rect 5050 14344 5092 14384
rect 5132 14344 5174 14384
rect 5214 14344 5256 14384
rect 4928 14335 5296 14344
rect 5452 14216 5492 14671
rect 5740 14552 5780 15847
rect 5836 14720 5876 16015
rect 5932 15737 5972 16192
rect 6028 16232 6068 16241
rect 6028 15905 6068 16192
rect 6027 15896 6069 15905
rect 6027 15856 6028 15896
rect 6068 15856 6069 15896
rect 6027 15847 6069 15856
rect 6124 15812 6164 20383
rect 6316 20264 6356 21568
rect 6412 21197 6452 22408
rect 6507 22399 6549 22408
rect 6508 22314 6548 22399
rect 6507 21524 6549 21533
rect 6507 21484 6508 21524
rect 6548 21484 6549 21524
rect 6507 21475 6549 21484
rect 6508 21440 6548 21475
rect 6604 21449 6644 23080
rect 6700 23120 6740 23129
rect 6700 21785 6740 23080
rect 6796 23120 6836 23129
rect 6796 22457 6836 23080
rect 6892 23120 6932 23129
rect 6892 23045 6932 23080
rect 6891 23036 6933 23045
rect 6891 22996 6892 23036
rect 6932 22996 6933 23036
rect 6891 22987 6933 22996
rect 6892 22985 6932 22987
rect 6988 22457 7028 23407
rect 7084 23288 7124 23752
rect 7180 23465 7220 24592
rect 7179 23456 7221 23465
rect 7179 23416 7180 23456
rect 7220 23416 7221 23456
rect 7179 23407 7221 23416
rect 7084 23248 7220 23288
rect 7180 23120 7220 23248
rect 7180 23045 7220 23080
rect 7179 23036 7221 23045
rect 7179 22996 7180 23036
rect 7220 22996 7221 23036
rect 7179 22987 7221 22996
rect 7180 22956 7220 22987
rect 7083 22700 7125 22709
rect 7083 22660 7084 22700
rect 7124 22660 7125 22700
rect 7083 22651 7125 22660
rect 6795 22448 6837 22457
rect 6795 22408 6796 22448
rect 6836 22408 6837 22448
rect 6795 22399 6837 22408
rect 6987 22448 7029 22457
rect 6987 22408 6988 22448
rect 7028 22408 7029 22448
rect 6987 22399 7029 22408
rect 6796 22280 6836 22399
rect 6796 22231 6836 22240
rect 7084 22280 7124 22651
rect 7084 22231 7124 22240
rect 7180 22205 7220 22290
rect 7179 22196 7221 22205
rect 7179 22156 7180 22196
rect 7220 22156 7221 22196
rect 7179 22147 7221 22156
rect 7276 21785 7316 25096
rect 6699 21776 6741 21785
rect 6699 21736 6700 21776
rect 6740 21736 6741 21776
rect 6699 21727 6741 21736
rect 7275 21776 7317 21785
rect 7275 21736 7276 21776
rect 7316 21736 7317 21776
rect 7275 21727 7317 21736
rect 7372 21701 7412 26011
rect 7467 25136 7509 25145
rect 7467 25096 7468 25136
rect 7508 25096 7509 25136
rect 7467 25087 7509 25096
rect 7468 25002 7508 25087
rect 7564 23969 7604 28120
rect 7659 26144 7701 26153
rect 7659 26104 7660 26144
rect 7700 26104 7701 26144
rect 7659 26095 7701 26104
rect 7660 25304 7700 26095
rect 7660 25255 7700 25264
rect 7659 25136 7701 25145
rect 7659 25096 7660 25136
rect 7700 25096 7701 25136
rect 7659 25087 7701 25096
rect 7660 24632 7700 25087
rect 7660 24583 7700 24592
rect 7756 24464 7796 30883
rect 7851 30260 7893 30269
rect 7851 30220 7852 30260
rect 7892 30220 7893 30260
rect 7851 30211 7893 30220
rect 7852 29000 7892 30211
rect 7852 28951 7892 28960
rect 7948 29840 7988 31312
rect 8332 31303 8372 31312
rect 8427 31352 8469 31361
rect 8427 31312 8428 31352
rect 8468 31312 8469 31352
rect 8427 31303 8469 31312
rect 8428 31218 8468 31303
rect 8524 31109 8564 31471
rect 8523 31100 8565 31109
rect 8523 31060 8524 31100
rect 8564 31060 8565 31100
rect 8523 31051 8565 31060
rect 8620 30941 8660 32992
rect 8716 32864 8756 32873
rect 8716 32621 8756 32824
rect 8811 32864 8853 32873
rect 8811 32824 8812 32864
rect 8852 32824 8853 32864
rect 8811 32815 8853 32824
rect 9004 32864 9044 34084
rect 9100 33041 9140 34159
rect 9387 33956 9429 33965
rect 9387 33916 9388 33956
rect 9428 33916 9524 33956
rect 9387 33907 9429 33916
rect 9484 33872 9524 33916
rect 9484 33832 9528 33872
rect 9388 33704 9428 33713
rect 9488 33704 9528 33832
rect 9580 33788 9620 34327
rect 9676 33872 9716 34504
rect 9772 34494 9812 34579
rect 9868 34365 9908 34374
rect 9868 34217 9908 34325
rect 9867 34208 9909 34217
rect 9867 34168 9868 34208
rect 9908 34168 9909 34208
rect 9867 34159 9909 34168
rect 9964 34040 10004 34663
rect 10060 34628 10100 35167
rect 10060 34579 10100 34588
rect 9964 34000 10100 34040
rect 9676 33832 9908 33872
rect 9580 33748 9812 33788
rect 9383 33664 9388 33704
rect 9383 33655 9428 33664
rect 9484 33664 9528 33704
rect 9772 33704 9812 33748
rect 9383 33536 9423 33655
rect 9484 33620 9524 33664
rect 9772 33655 9812 33664
rect 9484 33571 9524 33580
rect 9676 33620 9716 33631
rect 9676 33545 9716 33580
rect 9580 33536 9620 33545
rect 9383 33496 9428 33536
rect 9196 33452 9236 33461
rect 9291 33452 9333 33461
rect 9236 33412 9292 33452
rect 9332 33412 9333 33452
rect 9196 33403 9236 33412
rect 9291 33403 9333 33412
rect 9195 33116 9237 33125
rect 9195 33076 9196 33116
rect 9236 33076 9237 33116
rect 9195 33067 9237 33076
rect 9292 33116 9332 33125
rect 9388 33116 9428 33496
rect 9580 33293 9620 33496
rect 9675 33536 9717 33545
rect 9675 33496 9676 33536
rect 9716 33496 9717 33536
rect 9675 33487 9717 33496
rect 9579 33284 9621 33293
rect 9579 33244 9580 33284
rect 9620 33244 9621 33284
rect 9579 33235 9621 33244
rect 9332 33076 9428 33116
rect 9292 33067 9332 33076
rect 9099 33032 9141 33041
rect 9099 32992 9100 33032
rect 9140 32992 9141 33032
rect 9099 32983 9141 32992
rect 9004 32815 9044 32824
rect 9100 32864 9140 32873
rect 9196 32864 9236 33067
rect 9484 33041 9524 33126
rect 9483 33032 9525 33041
rect 9483 32992 9484 33032
rect 9524 32992 9525 33032
rect 9483 32983 9525 32992
rect 9387 32948 9429 32957
rect 9140 32824 9236 32864
rect 9292 32908 9388 32948
rect 9428 32908 9429 32948
rect 9292 32864 9332 32908
rect 9387 32899 9429 32908
rect 9676 32873 9716 32958
rect 9100 32815 9140 32824
rect 9292 32815 9332 32824
rect 9483 32864 9525 32873
rect 9483 32824 9484 32864
rect 9524 32824 9525 32864
rect 9483 32815 9525 32824
rect 9675 32864 9717 32873
rect 9675 32824 9676 32864
rect 9716 32824 9717 32864
rect 9675 32815 9717 32824
rect 9772 32864 9812 32873
rect 9868 32864 9908 33832
rect 9963 33788 10005 33797
rect 9963 33748 9964 33788
rect 10004 33748 10005 33788
rect 9963 33739 10005 33748
rect 9964 33704 10004 33739
rect 9964 33653 10004 33664
rect 9963 33452 10005 33461
rect 9963 33412 9964 33452
rect 10004 33412 10005 33452
rect 9963 33403 10005 33412
rect 9812 32824 9908 32864
rect 9964 32864 10004 33403
rect 9772 32815 9812 32824
rect 9964 32815 10004 32824
rect 8812 32730 8852 32815
rect 9387 32780 9429 32789
rect 9387 32740 9388 32780
rect 9428 32740 9429 32780
rect 9387 32731 9429 32740
rect 8715 32612 8757 32621
rect 8715 32572 8716 32612
rect 8756 32572 8757 32612
rect 8715 32563 8757 32572
rect 8715 32192 8757 32201
rect 8715 32152 8716 32192
rect 8756 32152 8757 32192
rect 8715 32143 8757 32152
rect 8716 32058 8756 32143
rect 8907 31520 8949 31529
rect 8907 31480 8908 31520
rect 8948 31480 8949 31520
rect 8907 31471 8949 31480
rect 8908 31436 8948 31471
rect 8908 31385 8948 31396
rect 8812 31352 8852 31363
rect 8812 31277 8852 31312
rect 9388 31352 9428 32731
rect 9484 32730 9524 32815
rect 10060 32780 10100 34000
rect 10156 33293 10196 35348
rect 10251 35216 10293 35225
rect 10251 35176 10252 35216
rect 10292 35176 10293 35216
rect 10251 35167 10293 35176
rect 10348 35216 10388 35225
rect 10252 35082 10292 35167
rect 10348 34973 10388 35176
rect 10347 34964 10389 34973
rect 10347 34924 10348 34964
rect 10388 34924 10389 34964
rect 10347 34915 10389 34924
rect 10251 34376 10293 34385
rect 10251 34336 10252 34376
rect 10292 34336 10293 34376
rect 10251 34327 10293 34336
rect 10252 34133 10292 34327
rect 10347 34208 10389 34217
rect 10347 34168 10348 34208
rect 10388 34168 10389 34208
rect 10347 34159 10389 34168
rect 10251 34124 10293 34133
rect 10251 34084 10252 34124
rect 10292 34084 10293 34124
rect 10251 34075 10293 34084
rect 10251 33788 10293 33797
rect 10251 33748 10252 33788
rect 10292 33748 10293 33788
rect 10251 33739 10293 33748
rect 10252 33461 10292 33739
rect 10251 33452 10293 33461
rect 10251 33412 10252 33452
rect 10292 33412 10293 33452
rect 10251 33403 10293 33412
rect 10155 33284 10197 33293
rect 10155 33244 10156 33284
rect 10196 33244 10197 33284
rect 10155 33235 10197 33244
rect 10156 32864 10196 32873
rect 10348 32864 10388 34159
rect 10444 33209 10484 35596
rect 10443 33200 10485 33209
rect 10443 33160 10444 33200
rect 10484 33160 10485 33200
rect 10443 33151 10485 33160
rect 10540 33032 10580 37939
rect 10924 37325 10964 40375
rect 11020 40349 11060 42928
rect 11019 40340 11061 40349
rect 11019 40300 11020 40340
rect 11060 40300 11061 40340
rect 11019 40291 11061 40300
rect 11115 39080 11157 39089
rect 11115 39040 11116 39080
rect 11156 39040 11157 39080
rect 11115 39031 11157 39040
rect 11116 38996 11156 39031
rect 11116 38945 11156 38956
rect 11019 38912 11061 38921
rect 11019 38872 11020 38912
rect 11060 38872 11061 38912
rect 11019 38863 11061 38872
rect 11020 38778 11060 38863
rect 10923 37316 10965 37325
rect 10923 37276 10924 37316
rect 10964 37276 10965 37316
rect 10923 37267 10965 37276
rect 11212 37148 11252 42928
rect 11404 42113 11444 42928
rect 11403 42104 11445 42113
rect 11403 42064 11404 42104
rect 11444 42064 11445 42104
rect 11403 42055 11445 42064
rect 11307 41684 11349 41693
rect 11596 41684 11636 42928
rect 11307 41644 11308 41684
rect 11348 41644 11349 41684
rect 11307 41635 11349 41644
rect 11404 41644 11636 41684
rect 11308 41357 11348 41635
rect 11307 41348 11349 41357
rect 11307 41308 11308 41348
rect 11348 41308 11349 41348
rect 11307 41299 11349 41308
rect 10636 37108 11252 37148
rect 10636 36317 10676 37108
rect 10731 36728 10773 36737
rect 11212 36728 11252 36737
rect 10731 36688 10732 36728
rect 10772 36688 10773 36728
rect 10731 36679 10773 36688
rect 11020 36688 11212 36728
rect 10732 36594 10772 36679
rect 10924 36476 10964 36485
rect 10635 36308 10677 36317
rect 10635 36268 10636 36308
rect 10676 36268 10677 36308
rect 10635 36259 10677 36268
rect 10924 36149 10964 36436
rect 10923 36140 10965 36149
rect 10923 36100 10924 36140
rect 10964 36100 10965 36140
rect 10923 36091 10965 36100
rect 11020 36140 11060 36688
rect 11212 36679 11252 36688
rect 11308 36728 11348 36737
rect 11115 36560 11157 36569
rect 11115 36520 11116 36560
rect 11156 36520 11157 36560
rect 11115 36511 11157 36520
rect 11020 36091 11060 36100
rect 10828 35909 10868 35918
rect 11116 35888 11156 36511
rect 11308 36392 11348 36688
rect 11404 36569 11444 41644
rect 11788 41525 11828 42928
rect 11883 42104 11925 42113
rect 11883 42064 11884 42104
rect 11924 42064 11925 42104
rect 11883 42055 11925 42064
rect 11787 41516 11829 41525
rect 11787 41476 11788 41516
rect 11828 41476 11829 41516
rect 11787 41467 11829 41476
rect 11884 41348 11924 42055
rect 11980 41936 12020 42928
rect 11980 41896 12116 41936
rect 11881 41308 11924 41348
rect 11881 41264 11921 41308
rect 11788 41224 11921 41264
rect 11980 41264 12020 41273
rect 11595 41180 11637 41189
rect 11595 41140 11596 41180
rect 11636 41140 11637 41180
rect 11595 41131 11637 41140
rect 11596 41046 11636 41131
rect 11788 41096 11828 41224
rect 11788 41047 11828 41056
rect 11980 40760 12020 41224
rect 12076 40937 12116 41896
rect 12075 40928 12117 40937
rect 12075 40888 12076 40928
rect 12116 40888 12117 40928
rect 12075 40879 12117 40888
rect 11692 40720 12020 40760
rect 11596 40445 11636 40454
rect 11500 40405 11596 40429
rect 11692 40433 11732 40720
rect 11980 40592 12020 40601
rect 11884 40552 11980 40592
rect 11500 40389 11636 40405
rect 11691 40424 11733 40433
rect 11500 40181 11540 40389
rect 11691 40384 11692 40424
rect 11732 40384 11733 40424
rect 11691 40375 11733 40384
rect 11787 40340 11829 40349
rect 11787 40300 11788 40340
rect 11828 40300 11829 40340
rect 11787 40291 11829 40300
rect 11788 40206 11828 40291
rect 11499 40172 11541 40181
rect 11499 40132 11500 40172
rect 11540 40132 11541 40172
rect 11499 40123 11541 40132
rect 11500 39752 11540 40123
rect 11787 40004 11829 40013
rect 11787 39964 11788 40004
rect 11828 39964 11829 40004
rect 11787 39955 11829 39964
rect 11692 39836 11732 39847
rect 11692 39761 11732 39796
rect 11500 38585 11540 39712
rect 11691 39752 11733 39761
rect 11691 39712 11692 39752
rect 11732 39712 11733 39752
rect 11691 39703 11733 39712
rect 11596 38912 11636 38921
rect 11788 38912 11828 39955
rect 11884 39752 11924 40552
rect 11980 40543 12020 40552
rect 11980 40424 12020 40435
rect 11980 40349 12020 40384
rect 12076 40424 12116 40433
rect 11979 40340 12021 40349
rect 11979 40300 11980 40340
rect 12020 40300 12021 40340
rect 11979 40291 12021 40300
rect 12076 40088 12116 40384
rect 12172 40097 12212 42928
rect 12364 42617 12404 42928
rect 12363 42608 12405 42617
rect 12363 42568 12364 42608
rect 12404 42568 12405 42608
rect 12363 42559 12405 42568
rect 12556 41609 12596 42928
rect 12555 41600 12597 41609
rect 12555 41560 12556 41600
rect 12596 41560 12597 41600
rect 12555 41551 12597 41560
rect 12267 40424 12309 40433
rect 12267 40384 12268 40424
rect 12308 40384 12309 40424
rect 12267 40375 12309 40384
rect 12556 40424 12596 40433
rect 12748 40424 12788 42928
rect 12748 40384 12884 40424
rect 12268 40290 12308 40375
rect 12363 40340 12405 40349
rect 12363 40300 12364 40340
rect 12404 40300 12405 40340
rect 12363 40291 12405 40300
rect 11980 40048 12116 40088
rect 12171 40088 12213 40097
rect 12171 40048 12172 40088
rect 12212 40048 12213 40088
rect 11980 39761 12020 40048
rect 12171 40039 12213 40048
rect 12076 39920 12116 39929
rect 11884 39703 11924 39712
rect 11979 39752 12021 39761
rect 11979 39712 11980 39752
rect 12020 39712 12021 39752
rect 11979 39703 12021 39712
rect 11980 39618 12020 39703
rect 11979 39332 12021 39341
rect 11979 39292 11980 39332
rect 12020 39292 12021 39332
rect 11979 39283 12021 39292
rect 11636 38872 11828 38912
rect 11596 38863 11636 38872
rect 11499 38576 11541 38585
rect 11499 38536 11500 38576
rect 11540 38536 11541 38576
rect 11499 38527 11541 38536
rect 11883 38576 11925 38585
rect 11883 38536 11884 38576
rect 11924 38536 11925 38576
rect 11883 38527 11925 38536
rect 11884 38240 11924 38527
rect 11884 38191 11924 38200
rect 11595 37736 11637 37745
rect 11595 37696 11596 37736
rect 11636 37696 11637 37736
rect 11595 37687 11637 37696
rect 11500 37400 11540 37409
rect 11596 37400 11636 37687
rect 11540 37360 11636 37400
rect 11500 37351 11540 37360
rect 11403 36560 11445 36569
rect 11403 36520 11404 36560
rect 11444 36520 11445 36560
rect 11403 36511 11445 36520
rect 11308 36352 11444 36392
rect 11307 36140 11349 36149
rect 11307 36100 11308 36140
rect 11348 36100 11349 36140
rect 11307 36091 11349 36100
rect 10731 35720 10773 35729
rect 10731 35680 10732 35720
rect 10772 35680 10773 35720
rect 10731 35671 10773 35680
rect 10636 34922 10676 34931
rect 10636 34049 10676 34882
rect 10635 34040 10677 34049
rect 10635 34000 10636 34040
rect 10676 34000 10677 34040
rect 10635 33991 10677 34000
rect 10540 32992 10676 33032
rect 10196 32824 10388 32864
rect 10156 32815 10196 32824
rect 10060 32731 10100 32740
rect 9675 32696 9717 32705
rect 9675 32656 9676 32696
rect 9716 32656 9717 32696
rect 9675 32647 9717 32656
rect 9579 32360 9621 32369
rect 9579 32320 9580 32360
rect 9620 32320 9621 32360
rect 9579 32311 9621 32320
rect 9428 31312 9524 31352
rect 9388 31303 9428 31312
rect 8811 31268 8853 31277
rect 8811 31228 8812 31268
rect 8852 31228 8853 31268
rect 8811 31219 8853 31228
rect 8619 30932 8661 30941
rect 8619 30892 8620 30932
rect 8660 30892 8661 30932
rect 8619 30883 8661 30892
rect 9099 30932 9141 30941
rect 9099 30892 9100 30932
rect 9140 30892 9141 30932
rect 9099 30883 9141 30892
rect 8812 30848 8852 30857
rect 8716 30808 8812 30848
rect 8619 30764 8661 30773
rect 8619 30724 8620 30764
rect 8660 30724 8661 30764
rect 8619 30715 8661 30724
rect 8524 30680 8564 30689
rect 8524 30269 8564 30640
rect 8620 30680 8660 30715
rect 8620 30629 8660 30640
rect 8716 30512 8756 30808
rect 8812 30799 8852 30808
rect 9003 30680 9045 30689
rect 9003 30640 9004 30680
rect 9044 30640 9045 30680
rect 9003 30631 9045 30640
rect 9004 30546 9044 30631
rect 9100 30521 9140 30883
rect 8620 30472 8756 30512
rect 9099 30512 9141 30521
rect 9099 30472 9100 30512
rect 9140 30472 9141 30512
rect 8523 30260 8565 30269
rect 8523 30220 8524 30260
rect 8564 30220 8565 30260
rect 8523 30211 8565 30220
rect 7948 28496 7988 29800
rect 8332 29840 8372 29849
rect 8140 29756 8180 29765
rect 8332 29756 8372 29800
rect 8180 29716 8372 29756
rect 8140 29707 8180 29716
rect 8428 29672 8468 29681
rect 8620 29672 8660 30472
rect 9099 30463 9141 30472
rect 8811 30260 8853 30269
rect 8811 30220 8812 30260
rect 8852 30220 8853 30260
rect 8811 30211 8853 30220
rect 8812 30017 8852 30211
rect 8811 30008 8853 30017
rect 8811 29968 8812 30008
rect 8852 29968 8853 30008
rect 8811 29959 8853 29968
rect 9387 30008 9429 30017
rect 9387 29968 9388 30008
rect 9428 29968 9429 30008
rect 9387 29959 9429 29968
rect 8716 29849 8756 29934
rect 8715 29840 8757 29849
rect 8715 29800 8716 29840
rect 8756 29800 8757 29840
rect 8715 29791 8757 29800
rect 8812 29840 8852 29959
rect 9004 29849 9044 29934
rect 8812 29765 8852 29800
rect 9003 29840 9045 29849
rect 9196 29840 9236 29849
rect 9003 29800 9004 29840
rect 9044 29800 9045 29840
rect 9003 29791 9045 29800
rect 9100 29800 9196 29840
rect 8811 29756 8853 29765
rect 8811 29716 8812 29756
rect 8852 29716 8853 29756
rect 8811 29707 8853 29716
rect 8908 29672 8948 29681
rect 8236 29632 8428 29672
rect 8468 29632 8564 29672
rect 8620 29632 8756 29672
rect 8139 29336 8181 29345
rect 8139 29296 8140 29336
rect 8180 29296 8181 29336
rect 8139 29287 8181 29296
rect 8140 29168 8180 29287
rect 8140 29119 8180 29128
rect 8236 29168 8276 29632
rect 8428 29623 8468 29632
rect 8236 29119 8276 29128
rect 8332 29340 8372 29349
rect 8235 28832 8277 28841
rect 8235 28792 8236 28832
rect 8276 28792 8277 28832
rect 8235 28783 8277 28792
rect 7852 28456 7988 28496
rect 7852 28001 7892 28456
rect 7948 28328 7988 28337
rect 7851 27992 7893 28001
rect 7851 27952 7852 27992
rect 7892 27952 7893 27992
rect 7851 27943 7893 27952
rect 7852 27656 7892 27943
rect 7948 27824 7988 28288
rect 8044 28328 8084 28337
rect 8044 28001 8084 28288
rect 8043 27992 8085 28001
rect 8043 27952 8044 27992
rect 8084 27952 8085 27992
rect 8043 27943 8085 27952
rect 7948 27784 8084 27824
rect 7948 27656 7988 27665
rect 7852 27616 7948 27656
rect 7948 27607 7988 27616
rect 8044 25229 8084 27784
rect 8139 27572 8181 27581
rect 8139 27532 8140 27572
rect 8180 27532 8181 27572
rect 8139 27523 8181 27532
rect 8140 27488 8180 27523
rect 8140 27437 8180 27448
rect 8236 26909 8276 28783
rect 8332 28253 8372 29300
rect 8524 29168 8564 29632
rect 8524 29119 8564 29128
rect 8619 29168 8661 29177
rect 8619 29128 8620 29168
rect 8660 29128 8661 29168
rect 8716 29168 8756 29632
rect 8948 29632 9044 29672
rect 8908 29623 8948 29632
rect 8812 29345 8852 29430
rect 8811 29336 8853 29345
rect 8811 29296 8812 29336
rect 8852 29296 8853 29336
rect 8811 29287 8853 29296
rect 8907 29252 8949 29261
rect 8907 29212 8908 29252
rect 8948 29212 8949 29252
rect 8907 29203 8949 29212
rect 8812 29168 8852 29177
rect 8716 29128 8812 29168
rect 8619 29119 8661 29128
rect 8812 29119 8852 29128
rect 8908 29168 8948 29203
rect 9004 29177 9044 29632
rect 9004 29168 9049 29177
rect 9004 29128 9009 29168
rect 8620 29034 8660 29119
rect 8908 29117 8948 29128
rect 9009 29119 9049 29128
rect 8427 29000 8469 29009
rect 8427 28960 8428 29000
rect 8468 28960 8469 29000
rect 8427 28951 8469 28960
rect 8715 29000 8757 29009
rect 8715 28960 8716 29000
rect 8756 28960 8757 29000
rect 8715 28951 8757 28960
rect 8331 28244 8373 28253
rect 8331 28204 8332 28244
rect 8372 28204 8373 28244
rect 8331 28195 8373 28204
rect 8331 26984 8373 26993
rect 8331 26944 8332 26984
rect 8372 26944 8373 26984
rect 8331 26935 8373 26944
rect 8235 26900 8277 26909
rect 8235 26860 8236 26900
rect 8276 26860 8277 26900
rect 8235 26851 8277 26860
rect 8043 25220 8085 25229
rect 8043 25180 8044 25220
rect 8084 25180 8085 25220
rect 8043 25171 8085 25180
rect 7948 24632 7988 24641
rect 7660 24424 7796 24464
rect 7852 24592 7948 24632
rect 7563 23960 7605 23969
rect 7563 23920 7564 23960
rect 7604 23920 7605 23960
rect 7563 23911 7605 23920
rect 7564 23797 7604 23806
rect 7564 23381 7604 23757
rect 7660 23540 7700 24424
rect 7756 23708 7796 23717
rect 7852 23708 7892 24592
rect 7948 24583 7988 24592
rect 8044 24632 8084 24641
rect 7947 24464 7989 24473
rect 7947 24424 7948 24464
rect 7988 24424 7989 24464
rect 7947 24415 7989 24424
rect 7948 23792 7988 24415
rect 8044 24044 8084 24592
rect 8236 24128 8276 26851
rect 8332 26816 8372 26935
rect 8332 24641 8372 26776
rect 8428 25976 8468 28951
rect 8523 28328 8565 28337
rect 8523 28288 8524 28328
rect 8564 28288 8565 28328
rect 8523 28279 8565 28288
rect 8524 28194 8564 28279
rect 8524 27656 8564 27665
rect 8716 27656 8756 28951
rect 8907 28916 8949 28925
rect 8907 28876 8908 28916
rect 8948 28876 8949 28916
rect 8907 28867 8949 28876
rect 8811 27740 8853 27749
rect 8811 27700 8812 27740
rect 8852 27700 8853 27740
rect 8811 27691 8853 27700
rect 8564 27616 8756 27656
rect 8812 27656 8852 27691
rect 8524 27607 8564 27616
rect 8812 27605 8852 27616
rect 8811 27488 8853 27497
rect 8811 27448 8812 27488
rect 8852 27448 8853 27488
rect 8811 27439 8853 27448
rect 8715 27404 8757 27413
rect 8715 27364 8716 27404
rect 8756 27364 8757 27404
rect 8715 27355 8757 27364
rect 8523 26816 8565 26825
rect 8523 26776 8524 26816
rect 8564 26776 8565 26816
rect 8523 26767 8565 26776
rect 8524 26732 8564 26767
rect 8524 26681 8564 26692
rect 8428 25936 8564 25976
rect 8427 25808 8469 25817
rect 8427 25768 8428 25808
rect 8468 25768 8469 25808
rect 8427 25759 8469 25768
rect 8331 24632 8373 24641
rect 8331 24592 8332 24632
rect 8372 24592 8373 24632
rect 8331 24583 8373 24592
rect 8331 24380 8373 24389
rect 8331 24340 8332 24380
rect 8372 24340 8373 24380
rect 8331 24331 8373 24340
rect 8332 24246 8372 24331
rect 8236 24088 8372 24128
rect 8044 24004 8276 24044
rect 7948 23743 7988 23752
rect 8044 23792 8084 23803
rect 8044 23717 8084 23752
rect 8139 23792 8181 23801
rect 8139 23752 8140 23792
rect 8180 23752 8181 23792
rect 8139 23743 8181 23752
rect 8236 23792 8276 24004
rect 8236 23743 8276 23752
rect 7796 23668 7892 23708
rect 8043 23708 8085 23717
rect 8043 23668 8044 23708
rect 8084 23668 8085 23708
rect 7756 23659 7796 23668
rect 8043 23659 8085 23668
rect 8140 23658 8180 23743
rect 7660 23500 8276 23540
rect 7563 23372 7605 23381
rect 7563 23332 7564 23372
rect 7604 23332 7605 23372
rect 7563 23323 7605 23332
rect 8139 23288 8181 23297
rect 8139 23248 8140 23288
rect 8180 23248 8181 23288
rect 8139 23239 8181 23248
rect 7468 23129 7508 23214
rect 7755 23204 7797 23213
rect 7755 23164 7756 23204
rect 7796 23164 7797 23204
rect 7755 23155 7797 23164
rect 7467 23120 7509 23129
rect 7660 23120 7700 23129
rect 7467 23080 7468 23120
rect 7508 23080 7509 23120
rect 7467 23071 7509 23080
rect 7564 23080 7660 23120
rect 7468 22952 7508 22961
rect 7564 22952 7604 23080
rect 7660 23071 7700 23080
rect 7508 22912 7604 22952
rect 7468 22903 7508 22912
rect 7660 22868 7700 22877
rect 7563 22700 7605 22709
rect 7563 22660 7564 22700
rect 7604 22660 7605 22700
rect 7563 22651 7605 22660
rect 7468 22448 7508 22457
rect 7371 21692 7413 21701
rect 7371 21652 7372 21692
rect 7412 21652 7413 21692
rect 7371 21643 7413 21652
rect 6700 21608 6740 21617
rect 6508 21389 6548 21400
rect 6603 21440 6645 21449
rect 6603 21400 6604 21440
rect 6644 21400 6645 21440
rect 6603 21391 6645 21400
rect 6700 21197 6740 21568
rect 7083 21608 7125 21617
rect 7083 21568 7084 21608
rect 7124 21568 7125 21608
rect 7083 21559 7125 21568
rect 7276 21608 7316 21619
rect 6796 21524 6836 21533
rect 6411 21188 6453 21197
rect 6411 21148 6412 21188
rect 6452 21148 6453 21188
rect 6411 21139 6453 21148
rect 6699 21188 6741 21197
rect 6699 21148 6700 21188
rect 6740 21148 6741 21188
rect 6699 21139 6741 21148
rect 6412 21020 6452 21029
rect 6796 21020 6836 21484
rect 6988 21524 7028 21533
rect 6891 21440 6933 21449
rect 6891 21400 6892 21440
rect 6932 21400 6933 21440
rect 6891 21391 6933 21400
rect 6892 21306 6932 21391
rect 6891 21188 6933 21197
rect 6891 21148 6892 21188
rect 6932 21148 6933 21188
rect 6891 21139 6933 21148
rect 6452 20980 6836 21020
rect 6412 20971 6452 20980
rect 6699 20852 6741 20861
rect 6801 20852 6843 20861
rect 6699 20812 6700 20852
rect 6740 20812 6741 20852
rect 6699 20803 6741 20812
rect 6796 20812 6802 20852
rect 6842 20812 6843 20852
rect 6796 20803 6843 20812
rect 6700 20768 6740 20803
rect 6220 20224 6356 20264
rect 6604 20268 6644 20277
rect 6220 20021 6260 20224
rect 6412 20180 6452 20189
rect 6604 20180 6644 20228
rect 6452 20140 6644 20180
rect 6412 20131 6452 20140
rect 6316 20096 6356 20105
rect 6219 20012 6261 20021
rect 6219 19972 6220 20012
rect 6260 19972 6261 20012
rect 6219 19963 6261 19972
rect 6219 19844 6261 19853
rect 6219 19804 6220 19844
rect 6260 19804 6261 19844
rect 6219 19795 6261 19804
rect 6220 17165 6260 19795
rect 6316 19685 6356 20056
rect 6700 20096 6740 20728
rect 6796 20432 6836 20803
rect 6892 20516 6932 21139
rect 6988 20936 7028 21484
rect 7084 21474 7124 21559
rect 7276 21533 7316 21568
rect 7275 21524 7317 21533
rect 7275 21484 7276 21524
rect 7316 21484 7317 21524
rect 7275 21475 7317 21484
rect 7083 21356 7125 21365
rect 7371 21356 7413 21365
rect 7083 21316 7084 21356
rect 7124 21316 7125 21356
rect 7083 21307 7125 21316
rect 7276 21316 7372 21356
rect 7412 21316 7413 21356
rect 7084 21197 7124 21307
rect 7083 21188 7125 21197
rect 7083 21148 7084 21188
rect 7124 21148 7125 21188
rect 7083 21139 7125 21148
rect 6988 20896 7220 20936
rect 6988 20768 7028 20779
rect 6988 20693 7028 20728
rect 7083 20768 7125 20777
rect 7083 20728 7084 20768
rect 7124 20728 7125 20768
rect 7083 20719 7125 20728
rect 6987 20684 7029 20693
rect 6987 20644 6988 20684
rect 7028 20644 7029 20684
rect 6987 20635 7029 20644
rect 7084 20634 7124 20719
rect 6892 20476 7124 20516
rect 6796 20392 7028 20432
rect 6700 20047 6740 20056
rect 6795 20096 6837 20105
rect 6795 20056 6796 20096
rect 6836 20056 6837 20096
rect 6795 20047 6837 20056
rect 6796 19962 6836 20047
rect 6891 20012 6933 20021
rect 6891 19972 6892 20012
rect 6932 19972 6933 20012
rect 6891 19963 6933 19972
rect 6795 19844 6837 19853
rect 6795 19804 6796 19844
rect 6836 19804 6837 19844
rect 6795 19795 6837 19804
rect 6315 19676 6357 19685
rect 6315 19636 6316 19676
rect 6356 19636 6357 19676
rect 6315 19627 6357 19636
rect 6315 19256 6357 19265
rect 6315 19216 6316 19256
rect 6356 19216 6357 19256
rect 6315 19207 6357 19216
rect 6508 19256 6548 19265
rect 6316 19097 6356 19207
rect 6508 19097 6548 19216
rect 6315 19088 6357 19097
rect 6315 19048 6316 19088
rect 6356 19048 6357 19088
rect 6315 19039 6357 19048
rect 6507 19088 6549 19097
rect 6507 19048 6508 19088
rect 6548 19048 6549 19088
rect 6507 19039 6549 19048
rect 6603 18920 6645 18929
rect 6603 18880 6604 18920
rect 6644 18880 6645 18920
rect 6603 18871 6645 18880
rect 6507 18752 6549 18761
rect 6507 18712 6508 18752
rect 6548 18712 6549 18752
rect 6507 18703 6549 18712
rect 6411 17660 6453 17669
rect 6411 17620 6412 17660
rect 6452 17620 6453 17660
rect 6411 17611 6453 17620
rect 6219 17156 6261 17165
rect 6219 17116 6220 17156
rect 6260 17116 6261 17156
rect 6219 17107 6261 17116
rect 6220 16409 6260 17107
rect 6412 17067 6452 17611
rect 6412 17018 6452 17027
rect 6219 16400 6261 16409
rect 6508 16400 6548 18703
rect 6604 17501 6644 18871
rect 6796 18341 6836 19795
rect 6892 18584 6932 19963
rect 6795 18332 6837 18341
rect 6795 18292 6796 18332
rect 6836 18292 6837 18332
rect 6795 18283 6837 18292
rect 6700 17744 6740 17753
rect 6700 17669 6740 17704
rect 6699 17660 6741 17669
rect 6699 17620 6700 17660
rect 6740 17620 6741 17660
rect 6699 17611 6741 17620
rect 6603 17492 6645 17501
rect 6603 17452 6604 17492
rect 6644 17452 6645 17492
rect 6603 17443 6645 17452
rect 6219 16360 6220 16400
rect 6260 16360 6261 16400
rect 6219 16351 6261 16360
rect 6316 16360 6548 16400
rect 6219 16064 6261 16073
rect 6219 16024 6220 16064
rect 6260 16024 6261 16064
rect 6219 16015 6261 16024
rect 6220 15930 6260 16015
rect 6124 15772 6260 15812
rect 5931 15728 5973 15737
rect 5931 15688 5932 15728
rect 5972 15688 6068 15728
rect 5931 15679 5973 15688
rect 6028 14729 6068 15688
rect 5836 14671 5876 14680
rect 5931 14720 5973 14729
rect 5931 14680 5932 14720
rect 5972 14680 5973 14720
rect 6028 14720 6073 14729
rect 6028 14680 6033 14720
rect 5931 14671 5973 14680
rect 6033 14671 6073 14680
rect 5932 14586 5972 14671
rect 6220 14552 6260 15772
rect 5740 14503 5780 14512
rect 6124 14512 6260 14552
rect 5835 14468 5877 14477
rect 5835 14428 5836 14468
rect 5876 14428 5877 14468
rect 5835 14419 5877 14428
rect 4780 14176 5108 14216
rect 5452 14176 5780 14216
rect 5068 14048 5108 14176
rect 5068 13805 5108 14008
rect 5547 14048 5589 14057
rect 5547 14008 5548 14048
rect 5588 14008 5589 14048
rect 5547 13999 5589 14008
rect 5259 13964 5301 13973
rect 5259 13924 5260 13964
rect 5300 13924 5301 13964
rect 5259 13915 5301 13924
rect 5067 13796 5109 13805
rect 5067 13756 5068 13796
rect 5108 13756 5109 13796
rect 5067 13747 5109 13756
rect 4876 13208 4916 13217
rect 4300 10312 4436 10352
rect 4204 10228 4340 10268
rect 4300 10184 4340 10228
rect 4300 10135 4340 10144
rect 4203 10100 4245 10109
rect 4203 10060 4204 10100
rect 4244 10060 4245 10100
rect 4203 10051 4245 10060
rect 3860 9472 4148 9512
rect 3820 9463 3860 9472
rect 3724 9378 3764 9463
rect 3688 9092 4056 9101
rect 3728 9052 3770 9092
rect 3810 9052 3852 9092
rect 3892 9052 3934 9092
rect 3974 9052 4016 9092
rect 3688 9043 4056 9052
rect 3532 8623 3572 8632
rect 3243 8252 3285 8261
rect 3243 8212 3244 8252
rect 3284 8212 3285 8252
rect 3243 8203 3285 8212
rect 3436 8000 3476 8009
rect 3436 7841 3476 7960
rect 4108 7916 4148 9472
rect 4204 9428 4244 10051
rect 4204 9185 4244 9388
rect 4299 9428 4341 9437
rect 4396 9428 4436 10312
rect 4492 10312 4628 10352
rect 4684 13168 4876 13208
rect 4492 9521 4532 10312
rect 4684 10277 4724 13168
rect 4876 13159 4916 13168
rect 5260 13124 5300 13915
rect 5404 13217 5444 13226
rect 5444 13177 5492 13208
rect 5404 13168 5492 13177
rect 5260 13084 5396 13124
rect 4928 12872 5296 12881
rect 4968 12832 5010 12872
rect 5050 12832 5092 12872
rect 5132 12832 5174 12872
rect 5214 12832 5256 12872
rect 4928 12823 5296 12832
rect 5356 12536 5396 13084
rect 5452 12704 5492 13168
rect 5548 13124 5588 13999
rect 5643 13796 5685 13805
rect 5643 13756 5644 13796
rect 5684 13756 5685 13796
rect 5643 13747 5685 13756
rect 5548 13075 5588 13084
rect 5548 12704 5588 12713
rect 5452 12664 5548 12704
rect 5548 12655 5588 12664
rect 5356 12487 5396 12496
rect 5067 11864 5109 11873
rect 5067 11824 5068 11864
rect 5108 11824 5109 11864
rect 5067 11815 5109 11824
rect 5068 11696 5108 11815
rect 5068 11647 5108 11656
rect 4928 11360 5296 11369
rect 5644 11360 5684 13747
rect 4968 11320 5010 11360
rect 5050 11320 5092 11360
rect 5132 11320 5174 11360
rect 5214 11320 5256 11360
rect 4928 11311 5296 11320
rect 5452 11320 5684 11360
rect 5355 11108 5397 11117
rect 5355 11068 5356 11108
rect 5396 11068 5397 11108
rect 5355 11059 5397 11068
rect 5164 11024 5204 11033
rect 5164 10277 5204 10984
rect 5356 10974 5396 11059
rect 4683 10268 4725 10277
rect 4588 10228 4684 10268
rect 4724 10228 4725 10268
rect 4491 9512 4533 9521
rect 4491 9472 4492 9512
rect 4532 9472 4533 9512
rect 4491 9463 4533 9472
rect 4299 9388 4300 9428
rect 4340 9388 4436 9428
rect 4299 9379 4341 9388
rect 4300 9294 4340 9379
rect 4203 9176 4245 9185
rect 4203 9136 4204 9176
rect 4244 9136 4245 9176
rect 4203 9127 4245 9136
rect 4299 8252 4341 8261
rect 4299 8212 4300 8252
rect 4340 8212 4341 8252
rect 4299 8203 4341 8212
rect 4203 8168 4245 8177
rect 4203 8128 4204 8168
rect 4244 8128 4245 8168
rect 4203 8119 4245 8128
rect 4204 8042 4244 8119
rect 4204 7993 4244 8002
rect 4108 7876 4244 7916
rect 3435 7832 3477 7841
rect 3435 7792 3436 7832
rect 3476 7792 3477 7832
rect 3435 7783 3477 7792
rect 3339 6992 3381 7001
rect 3339 6952 3340 6992
rect 3380 6952 3381 6992
rect 3339 6943 3381 6952
rect 3340 6488 3380 6943
rect 3340 6439 3380 6448
rect 3436 5900 3476 7783
rect 3628 7748 3668 7757
rect 3532 7708 3628 7748
rect 3532 7169 3572 7708
rect 3628 7699 3668 7708
rect 4107 7748 4149 7757
rect 4107 7708 4108 7748
rect 4148 7708 4149 7748
rect 4107 7699 4149 7708
rect 3688 7580 4056 7589
rect 3728 7540 3770 7580
rect 3810 7540 3852 7580
rect 3892 7540 3934 7580
rect 3974 7540 4016 7580
rect 3688 7531 4056 7540
rect 4108 7412 4148 7699
rect 3628 7372 4148 7412
rect 3531 7160 3573 7169
rect 3531 7120 3532 7160
rect 3572 7120 3573 7160
rect 3531 7111 3573 7120
rect 3628 7160 3668 7372
rect 3628 7111 3668 7120
rect 3915 7160 3957 7169
rect 3915 7120 3916 7160
rect 3956 7120 3957 7160
rect 3915 7111 3957 7120
rect 4012 7160 4052 7169
rect 3916 7026 3956 7111
rect 3819 6740 3861 6749
rect 3819 6700 3820 6740
rect 3860 6700 3861 6740
rect 3819 6691 3861 6700
rect 3820 6488 3860 6691
rect 3915 6572 3957 6581
rect 3915 6532 3916 6572
rect 3956 6532 3957 6572
rect 3915 6523 3957 6532
rect 3820 6439 3860 6448
rect 3916 6488 3956 6523
rect 3916 6437 3956 6448
rect 4012 6413 4052 7120
rect 4011 6404 4053 6413
rect 4011 6364 4012 6404
rect 4052 6364 4053 6404
rect 4011 6355 4053 6364
rect 3688 6068 4056 6077
rect 3728 6028 3770 6068
rect 3810 6028 3852 6068
rect 3892 6028 3934 6068
rect 3974 6028 4016 6068
rect 3688 6019 4056 6028
rect 3436 5860 3668 5900
rect 3436 5732 3476 5741
rect 3244 5480 3284 5489
rect 3147 4220 3189 4229
rect 3147 4180 3148 4220
rect 3188 4180 3189 4220
rect 3147 4171 3189 4180
rect 3004 4145 3044 4154
rect 2764 4105 3004 4136
rect 2764 4096 3044 4105
rect 2667 4052 2709 4061
rect 2667 4012 2668 4052
rect 2708 4012 2709 4052
rect 2667 4003 2709 4012
rect 2668 3918 2708 4003
rect 2668 3632 2708 3641
rect 2764 3632 2804 4096
rect 2859 3968 2901 3977
rect 2859 3928 2860 3968
rect 2900 3928 2901 3968
rect 2859 3919 2901 3928
rect 2860 3834 2900 3919
rect 2955 3800 2997 3809
rect 2955 3760 2956 3800
rect 2996 3760 2997 3800
rect 2955 3751 2997 3760
rect 2708 3592 2804 3632
rect 2668 3583 2708 3592
rect 2860 3464 2900 3473
rect 2956 3464 2996 3751
rect 2900 3424 2996 3464
rect 2860 3415 2900 3424
rect 3147 2792 3189 2801
rect 3147 2752 3148 2792
rect 3188 2752 3189 2792
rect 3147 2743 3189 2752
rect 3052 2624 3092 2633
rect 2572 2500 2996 2540
rect 2379 2491 2421 2500
rect 1515 2456 1557 2465
rect 1515 2416 1516 2456
rect 1556 2416 1557 2456
rect 1515 2407 1557 2416
rect 1803 2456 1845 2465
rect 1803 2416 1804 2456
rect 1844 2416 1845 2456
rect 1803 2407 1845 2416
rect 1419 2372 1461 2381
rect 1419 2332 1420 2372
rect 1460 2332 1461 2372
rect 1419 2323 1461 2332
rect 1516 2322 1556 2407
rect 1420 1952 1460 1961
rect 1420 1625 1460 1912
rect 1515 1784 1557 1793
rect 1515 1744 1516 1784
rect 1556 1744 1557 1784
rect 1515 1735 1557 1744
rect 1419 1616 1461 1625
rect 1419 1576 1420 1616
rect 1460 1576 1461 1616
rect 1419 1567 1461 1576
rect 1516 1280 1556 1735
rect 1516 1231 1556 1240
rect 1708 1196 1748 1205
rect 363 1112 405 1121
rect 363 1072 364 1112
rect 404 1072 405 1112
rect 363 1063 405 1072
rect 1708 1037 1748 1156
rect 1707 1028 1749 1037
rect 1707 988 1708 1028
rect 1748 988 1749 1028
rect 1707 979 1749 988
rect 1804 80 1844 2407
rect 1899 2120 1941 2129
rect 1899 2080 1900 2120
rect 1940 2080 1941 2120
rect 1899 2071 1941 2080
rect 1900 1280 1940 2071
rect 1900 1231 1940 1240
rect 1996 80 2036 2491
rect 2956 2381 2996 2500
rect 2091 2372 2133 2381
rect 2091 2332 2092 2372
rect 2132 2332 2133 2372
rect 2091 2323 2133 2332
rect 2955 2372 2997 2381
rect 2955 2332 2956 2372
rect 2996 2332 2997 2372
rect 2955 2323 2997 2332
rect 2092 1196 2132 2323
rect 2571 2204 2613 2213
rect 2571 2164 2572 2204
rect 2612 2164 2613 2204
rect 2571 2155 2613 2164
rect 2475 2120 2517 2129
rect 2475 2080 2476 2120
rect 2516 2080 2517 2120
rect 2475 2071 2517 2080
rect 2283 1448 2325 1457
rect 2283 1408 2284 1448
rect 2324 1408 2325 1448
rect 2283 1399 2325 1408
rect 2187 1364 2229 1373
rect 2187 1324 2188 1364
rect 2228 1324 2229 1364
rect 2187 1315 2229 1324
rect 2092 1147 2132 1156
rect 2188 80 2228 1315
rect 2284 1280 2324 1399
rect 2284 1231 2324 1240
rect 2476 1196 2516 2071
rect 2476 1147 2516 1156
rect 2379 692 2421 701
rect 2379 652 2380 692
rect 2420 652 2421 692
rect 2379 643 2421 652
rect 2380 80 2420 643
rect 2572 80 2612 2155
rect 2860 2120 2900 2129
rect 3052 2120 3092 2584
rect 3148 2624 3188 2743
rect 3148 2575 3188 2584
rect 3244 2540 3284 5440
rect 3339 5060 3381 5069
rect 3339 5020 3340 5060
rect 3380 5020 3381 5060
rect 3339 5011 3381 5020
rect 3340 4976 3380 5011
rect 3340 3809 3380 4936
rect 3339 3800 3381 3809
rect 3339 3760 3340 3800
rect 3380 3760 3381 3800
rect 3339 3751 3381 3760
rect 3436 2549 3476 5692
rect 3531 5060 3573 5069
rect 3531 5020 3532 5060
rect 3572 5020 3573 5060
rect 3531 5011 3573 5020
rect 3532 4926 3572 5011
rect 3628 4817 3668 5860
rect 3915 5060 3957 5069
rect 4107 5060 4149 5069
rect 3915 5020 3916 5060
rect 3956 5020 3957 5060
rect 3915 5011 3957 5020
rect 4012 5020 4108 5060
rect 4148 5020 4149 5060
rect 3916 4976 3956 5011
rect 3916 4925 3956 4936
rect 4012 4976 4052 5020
rect 4107 5011 4149 5020
rect 4012 4927 4052 4936
rect 3627 4808 3669 4817
rect 3627 4768 3628 4808
rect 3668 4768 3669 4808
rect 3627 4759 3669 4768
rect 3531 4724 3573 4733
rect 3531 4684 3532 4724
rect 3572 4684 3573 4724
rect 3531 4675 3573 4684
rect 3532 4136 3572 4675
rect 3688 4556 4056 4565
rect 3728 4516 3770 4556
rect 3810 4516 3852 4556
rect 3892 4516 3934 4556
rect 3974 4516 4016 4556
rect 3688 4507 4056 4516
rect 4108 4397 4148 5011
rect 4204 4817 4244 7876
rect 4300 6749 4340 8203
rect 4492 7505 4532 9463
rect 4491 7496 4533 7505
rect 4491 7456 4492 7496
rect 4532 7456 4533 7496
rect 4491 7447 4533 7456
rect 4491 7328 4533 7337
rect 4491 7288 4492 7328
rect 4532 7288 4533 7328
rect 4491 7279 4533 7288
rect 4395 7244 4437 7253
rect 4395 7204 4396 7244
rect 4436 7204 4437 7244
rect 4395 7195 4437 7204
rect 4492 7244 4532 7279
rect 4299 6740 4341 6749
rect 4299 6700 4300 6740
rect 4340 6700 4341 6740
rect 4396 6740 4436 7195
rect 4492 7193 4532 7204
rect 4396 6700 4532 6740
rect 4299 6691 4341 6700
rect 4396 6497 4436 6582
rect 4300 6488 4340 6497
rect 4300 6413 4340 6448
rect 4395 6488 4437 6497
rect 4395 6448 4396 6488
rect 4436 6448 4437 6488
rect 4395 6439 4437 6448
rect 4299 6404 4341 6413
rect 4299 6364 4300 6404
rect 4340 6364 4341 6404
rect 4492 6393 4532 6700
rect 4588 6581 4628 10228
rect 4683 10219 4725 10228
rect 5163 10268 5205 10277
rect 5163 10228 5164 10268
rect 5204 10228 5205 10268
rect 5163 10219 5205 10228
rect 4780 10189 4820 10198
rect 4683 9848 4725 9857
rect 4683 9808 4684 9848
rect 4724 9808 4725 9848
rect 4683 9799 4725 9808
rect 4684 9017 4724 9799
rect 4780 9680 4820 10149
rect 4971 10100 5013 10109
rect 4971 10060 4972 10100
rect 5012 10060 5013 10100
rect 4971 10051 5013 10060
rect 4972 9966 5012 10051
rect 4928 9848 5296 9857
rect 4968 9808 5010 9848
rect 5050 9808 5092 9848
rect 5132 9808 5174 9848
rect 5214 9808 5256 9848
rect 4928 9799 5296 9808
rect 5452 9764 5492 11320
rect 5643 11108 5685 11117
rect 5643 11068 5644 11108
rect 5684 11068 5685 11108
rect 5643 11059 5685 11068
rect 5644 11024 5684 11059
rect 5644 10973 5684 10984
rect 5740 11024 5780 14176
rect 5836 11276 5876 14419
rect 5931 14048 5973 14057
rect 5931 14008 5932 14048
rect 5972 14008 5973 14048
rect 5931 13999 5973 14008
rect 5932 11360 5972 13999
rect 5932 11320 6068 11360
rect 5836 11236 5972 11276
rect 5835 11108 5877 11117
rect 5835 11068 5836 11108
rect 5876 11068 5877 11108
rect 5835 11059 5877 11068
rect 5547 10352 5589 10361
rect 5547 10312 5548 10352
rect 5588 10312 5589 10352
rect 5547 10303 5589 10312
rect 5548 10184 5588 10303
rect 5548 10135 5588 10144
rect 5452 9724 5588 9764
rect 4780 9640 4916 9680
rect 4779 9512 4821 9521
rect 4779 9472 4780 9512
rect 4820 9472 4821 9512
rect 4779 9463 4821 9472
rect 4780 9378 4820 9463
rect 4683 9008 4725 9017
rect 4683 8968 4684 9008
rect 4724 8968 4725 9008
rect 4683 8959 4725 8968
rect 4683 8840 4725 8849
rect 4683 8800 4684 8840
rect 4724 8800 4725 8840
rect 4876 8840 4916 9640
rect 5451 9596 5493 9605
rect 5451 9556 5452 9596
rect 5492 9556 5493 9596
rect 5451 9547 5493 9556
rect 5308 9470 5348 9479
rect 5452 9462 5492 9547
rect 5308 9428 5348 9430
rect 5308 9388 5396 9428
rect 4972 8840 5012 8849
rect 4876 8800 4972 8840
rect 4683 8791 4725 8800
rect 4972 8791 5012 8800
rect 4684 7757 4724 8791
rect 4780 8672 4820 8683
rect 5356 8672 5396 9388
rect 5548 8849 5588 9724
rect 5740 8849 5780 10984
rect 5547 8840 5589 8849
rect 5547 8800 5548 8840
rect 5588 8800 5589 8840
rect 5547 8791 5589 8800
rect 5739 8840 5781 8849
rect 5739 8800 5740 8840
rect 5780 8800 5781 8840
rect 5739 8791 5781 8800
rect 5644 8672 5684 8681
rect 5356 8632 5588 8672
rect 4780 8597 4820 8632
rect 4779 8588 4821 8597
rect 4779 8548 4780 8588
rect 4820 8548 4821 8588
rect 4779 8539 4821 8548
rect 4780 8009 4820 8539
rect 4928 8336 5296 8345
rect 4968 8296 5010 8336
rect 5050 8296 5092 8336
rect 5132 8296 5174 8336
rect 5214 8296 5256 8336
rect 4928 8287 5296 8296
rect 5548 8168 5588 8632
rect 5684 8632 5780 8672
rect 5644 8623 5684 8632
rect 5740 8177 5780 8632
rect 5644 8168 5684 8177
rect 5548 8128 5644 8168
rect 5644 8119 5684 8128
rect 5739 8168 5781 8177
rect 5739 8128 5740 8168
rect 5780 8128 5781 8168
rect 5739 8119 5781 8128
rect 4779 8000 4821 8009
rect 4779 7960 4780 8000
rect 4820 7960 4821 8000
rect 4779 7951 4821 7960
rect 5452 8000 5492 8009
rect 5452 7841 5492 7960
rect 5451 7832 5493 7841
rect 5451 7792 5452 7832
rect 5492 7792 5493 7832
rect 5451 7783 5493 7792
rect 4683 7748 4725 7757
rect 4683 7708 4684 7748
rect 4724 7708 4725 7748
rect 4683 7699 4725 7708
rect 4587 6572 4629 6581
rect 4587 6532 4588 6572
rect 4628 6532 4629 6572
rect 4587 6523 4629 6532
rect 4684 6488 4724 7699
rect 4779 7496 4821 7505
rect 4779 7456 4780 7496
rect 4820 7456 4821 7496
rect 4779 7447 4821 7456
rect 4684 6439 4724 6448
rect 4299 6355 4341 6364
rect 4203 4808 4245 4817
rect 4203 4768 4204 4808
rect 4244 4768 4245 4808
rect 4203 4759 4245 4768
rect 4203 4640 4245 4649
rect 4203 4600 4204 4640
rect 4244 4600 4245 4640
rect 4203 4591 4245 4600
rect 4107 4388 4149 4397
rect 4012 4348 4108 4388
rect 4148 4348 4149 4388
rect 4012 4220 4052 4348
rect 4107 4339 4149 4348
rect 4204 4304 4244 4591
rect 4300 4565 4340 6355
rect 4396 6353 4532 6393
rect 4396 4976 4436 6353
rect 4491 6236 4533 6245
rect 4491 6196 4492 6236
rect 4532 6196 4533 6236
rect 4491 6187 4533 6196
rect 4492 5657 4532 6187
rect 4491 5648 4533 5657
rect 4491 5608 4492 5648
rect 4532 5608 4533 5648
rect 4491 5599 4533 5608
rect 4492 5514 4532 5599
rect 4780 5396 4820 7447
rect 5836 7328 5876 11059
rect 5356 7288 5876 7328
rect 4971 7244 5013 7253
rect 4971 7204 4972 7244
rect 5012 7204 5013 7244
rect 4971 7195 5013 7204
rect 4972 7160 5012 7195
rect 4972 7001 5012 7120
rect 4971 6992 5013 7001
rect 4971 6952 4972 6992
rect 5012 6952 5013 6992
rect 4971 6943 5013 6952
rect 4928 6824 5296 6833
rect 4968 6784 5010 6824
rect 5050 6784 5092 6824
rect 5132 6784 5174 6824
rect 5214 6784 5256 6824
rect 4928 6775 5296 6784
rect 4396 4927 4436 4936
rect 4492 5356 4820 5396
rect 4492 4976 4532 5356
rect 4928 5312 5296 5321
rect 4968 5272 5010 5312
rect 5050 5272 5092 5312
rect 5132 5272 5174 5312
rect 5214 5272 5256 5312
rect 4928 5263 5296 5272
rect 4972 4976 5012 4985
rect 4395 4808 4437 4817
rect 4395 4768 4396 4808
rect 4436 4768 4437 4808
rect 4395 4759 4437 4768
rect 4299 4556 4341 4565
rect 4299 4516 4300 4556
rect 4340 4516 4341 4556
rect 4299 4507 4341 4516
rect 4299 4304 4341 4313
rect 4204 4264 4300 4304
rect 4340 4264 4341 4304
rect 4299 4255 4341 4264
rect 4012 4171 4052 4180
rect 4107 4220 4149 4229
rect 4107 4180 4108 4220
rect 4148 4180 4149 4220
rect 4107 4171 4149 4180
rect 3532 2624 3572 4096
rect 4108 4086 4148 4171
rect 4107 3968 4149 3977
rect 4107 3928 4108 3968
rect 4148 3928 4149 3968
rect 4107 3919 4149 3928
rect 4108 3464 4148 3919
rect 4108 3415 4148 3424
rect 4300 3464 4340 4255
rect 4396 3968 4436 4759
rect 4492 4733 4532 4936
rect 4780 4936 4972 4976
rect 4491 4724 4533 4733
rect 4491 4684 4492 4724
rect 4532 4684 4533 4724
rect 4491 4675 4533 4684
rect 4491 4556 4533 4565
rect 4491 4516 4492 4556
rect 4532 4516 4533 4556
rect 4491 4507 4533 4516
rect 4492 4136 4532 4507
rect 4492 4087 4532 4096
rect 4588 4136 4628 4147
rect 4588 4061 4628 4096
rect 4587 4052 4629 4061
rect 4587 4012 4588 4052
rect 4628 4012 4629 4052
rect 4587 4003 4629 4012
rect 4683 3968 4725 3977
rect 4396 3928 4532 3968
rect 4395 3800 4437 3809
rect 4395 3760 4396 3800
rect 4436 3760 4437 3800
rect 4395 3751 4437 3760
rect 4396 3473 4436 3751
rect 4300 3415 4340 3424
rect 4395 3464 4437 3473
rect 4395 3424 4396 3464
rect 4436 3424 4437 3464
rect 4395 3415 4437 3424
rect 3688 3044 4056 3053
rect 3728 3004 3770 3044
rect 3810 3004 3852 3044
rect 3892 3004 3934 3044
rect 3974 3004 4016 3044
rect 3688 2995 4056 3004
rect 4107 2876 4149 2885
rect 4107 2836 4108 2876
rect 4148 2836 4149 2876
rect 4107 2827 4149 2836
rect 3628 2633 3668 2718
rect 3532 2575 3572 2584
rect 3627 2624 3669 2633
rect 3627 2584 3628 2624
rect 3668 2584 3669 2624
rect 3627 2575 3669 2584
rect 4108 2624 4148 2827
rect 4108 2575 4148 2584
rect 3435 2540 3477 2549
rect 3244 2500 3380 2540
rect 3147 2372 3189 2381
rect 3147 2332 3148 2372
rect 3188 2332 3189 2372
rect 3147 2323 3189 2332
rect 2900 2080 3092 2120
rect 2860 2071 2900 2080
rect 3148 2036 3188 2323
rect 3052 1996 3284 2036
rect 3052 1994 3092 1996
rect 2667 1952 2709 1961
rect 2667 1912 2668 1952
rect 2708 1912 2709 1952
rect 3052 1945 3092 1954
rect 2667 1903 2709 1912
rect 2668 1818 2708 1903
rect 2859 1700 2901 1709
rect 2859 1660 2860 1700
rect 2900 1660 2901 1700
rect 2859 1651 2901 1660
rect 2763 1280 2805 1289
rect 2763 1240 2764 1280
rect 2804 1240 2805 1280
rect 2763 1231 2805 1240
rect 2668 944 2708 953
rect 2668 197 2708 904
rect 2667 188 2709 197
rect 2667 148 2668 188
rect 2708 148 2709 188
rect 2667 139 2709 148
rect 2764 80 2804 1231
rect 2860 1196 2900 1651
rect 2955 1280 2997 1289
rect 2955 1240 2956 1280
rect 2996 1240 2997 1280
rect 2955 1231 2997 1240
rect 3147 1280 3189 1289
rect 3147 1240 3148 1280
rect 3188 1240 3189 1280
rect 3147 1231 3189 1240
rect 2860 1147 2900 1156
rect 2956 80 2996 1231
rect 3148 80 3188 1231
rect 3244 1112 3284 1996
rect 3244 1063 3284 1072
rect 3340 785 3380 2500
rect 3435 2500 3436 2540
rect 3476 2500 3477 2540
rect 3435 2491 3477 2500
rect 3723 2540 3765 2549
rect 3723 2500 3724 2540
rect 3764 2500 3765 2540
rect 3723 2491 3765 2500
rect 4203 2540 4245 2549
rect 4203 2500 4204 2540
rect 4244 2500 4245 2540
rect 4203 2491 4245 2500
rect 3724 1793 3764 2491
rect 3723 1784 3765 1793
rect 3723 1744 3724 1784
rect 3764 1744 3765 1784
rect 3723 1735 3765 1744
rect 3688 1532 4056 1541
rect 3728 1492 3770 1532
rect 3810 1492 3852 1532
rect 3892 1492 3934 1532
rect 3974 1492 4016 1532
rect 3688 1483 4056 1492
rect 3531 1280 3573 1289
rect 3531 1240 3532 1280
rect 3572 1240 3573 1280
rect 3531 1231 3573 1240
rect 3339 776 3381 785
rect 3339 736 3340 776
rect 3380 736 3381 776
rect 3339 727 3381 736
rect 3339 608 3381 617
rect 3339 568 3340 608
rect 3380 568 3381 608
rect 3339 559 3381 568
rect 3340 80 3380 559
rect 3532 80 3572 1231
rect 3915 1196 3957 1205
rect 3915 1156 3916 1196
rect 3956 1156 3957 1196
rect 3915 1147 3957 1156
rect 3723 356 3765 365
rect 3723 316 3724 356
rect 3764 316 3765 356
rect 3723 307 3765 316
rect 3724 80 3764 307
rect 3916 80 3956 1147
rect 4107 860 4149 869
rect 4107 820 4108 860
rect 4148 820 4149 860
rect 4107 811 4149 820
rect 4108 80 4148 811
rect 4204 449 4244 2491
rect 4396 1961 4436 3415
rect 4492 2801 4532 3928
rect 4683 3928 4684 3968
rect 4724 3928 4725 3968
rect 4683 3919 4725 3928
rect 4491 2792 4533 2801
rect 4491 2752 4492 2792
rect 4532 2752 4533 2792
rect 4491 2743 4533 2752
rect 4491 2624 4533 2633
rect 4491 2584 4492 2624
rect 4532 2584 4533 2624
rect 4491 2575 4533 2584
rect 4588 2629 4628 2638
rect 4492 2120 4532 2575
rect 4492 2071 4532 2080
rect 4300 1952 4340 1961
rect 4300 1457 4340 1912
rect 4395 1952 4437 1961
rect 4395 1912 4396 1952
rect 4436 1912 4437 1952
rect 4395 1903 4437 1912
rect 4299 1448 4341 1457
rect 4299 1408 4300 1448
rect 4340 1408 4341 1448
rect 4299 1399 4341 1408
rect 4299 1112 4341 1121
rect 4299 1072 4300 1112
rect 4340 1072 4341 1112
rect 4396 1112 4436 1903
rect 4588 1280 4628 2589
rect 4684 1952 4724 3919
rect 4780 2969 4820 4936
rect 4972 4927 5012 4936
rect 5067 4220 5109 4229
rect 5067 4180 5068 4220
rect 5108 4180 5109 4220
rect 5067 4171 5109 4180
rect 5068 4086 5108 4171
rect 4876 3977 4916 4062
rect 4875 3968 4917 3977
rect 4875 3928 4876 3968
rect 4916 3928 4917 3968
rect 4875 3919 4917 3928
rect 4928 3800 5296 3809
rect 4968 3760 5010 3800
rect 5050 3760 5092 3800
rect 5132 3760 5174 3800
rect 5214 3760 5256 3800
rect 4928 3751 5296 3760
rect 4779 2960 4821 2969
rect 4779 2920 4780 2960
rect 4820 2920 4821 2960
rect 4779 2911 4821 2920
rect 4779 2708 4821 2717
rect 4779 2668 4780 2708
rect 4820 2668 4821 2708
rect 4779 2659 4821 2668
rect 5163 2708 5205 2717
rect 5163 2668 5164 2708
rect 5204 2668 5205 2708
rect 5163 2659 5205 2668
rect 4780 2540 4820 2659
rect 5164 2574 5204 2659
rect 4780 2491 4820 2500
rect 4875 2540 4917 2549
rect 4875 2500 4876 2540
rect 4916 2500 5012 2540
rect 4875 2491 4917 2500
rect 4972 2456 5012 2500
rect 4972 2407 5012 2416
rect 4928 2288 5296 2297
rect 4968 2248 5010 2288
rect 5050 2248 5092 2288
rect 5132 2248 5174 2288
rect 5214 2248 5256 2288
rect 4928 2239 5296 2248
rect 4875 2036 4917 2045
rect 4875 1996 4876 2036
rect 4916 1996 4917 2036
rect 4875 1987 4917 1996
rect 4684 1903 4724 1912
rect 4684 1280 4724 1289
rect 4588 1240 4684 1280
rect 4684 1231 4724 1240
rect 4876 1196 4916 1987
rect 5356 1280 5396 7288
rect 5932 7244 5972 11236
rect 5740 7204 5972 7244
rect 5500 7169 5540 7178
rect 5540 7129 5588 7160
rect 5500 7120 5588 7129
rect 5548 5909 5588 7120
rect 5643 6992 5685 7001
rect 5643 6952 5644 6992
rect 5684 6952 5685 6992
rect 5643 6943 5685 6952
rect 5644 6858 5684 6943
rect 5643 6740 5685 6749
rect 5643 6700 5644 6740
rect 5684 6700 5685 6740
rect 5643 6691 5685 6700
rect 5547 5900 5589 5909
rect 5547 5860 5548 5900
rect 5588 5860 5589 5900
rect 5547 5851 5589 5860
rect 5644 5228 5684 6691
rect 5740 5816 5780 7204
rect 5835 6740 5877 6749
rect 5835 6700 5836 6740
rect 5876 6700 5877 6740
rect 5835 6691 5877 6700
rect 5836 6068 5876 6691
rect 5931 6488 5973 6497
rect 5931 6448 5932 6488
rect 5972 6448 5973 6488
rect 5931 6439 5973 6448
rect 5932 6354 5972 6439
rect 6028 6152 6068 11320
rect 6124 11117 6164 14512
rect 6316 14216 6356 16360
rect 6508 16232 6548 16360
rect 6508 16183 6548 16192
rect 6604 17156 6644 17165
rect 6412 16064 6452 16073
rect 6412 14729 6452 16024
rect 6507 14804 6549 14813
rect 6507 14764 6508 14804
rect 6548 14764 6549 14804
rect 6507 14755 6549 14764
rect 6411 14720 6453 14729
rect 6411 14680 6412 14720
rect 6452 14680 6453 14720
rect 6411 14671 6453 14680
rect 6508 14720 6548 14755
rect 6508 14669 6548 14680
rect 6604 14393 6644 17116
rect 6700 16493 6740 17611
rect 6699 16484 6741 16493
rect 6699 16444 6700 16484
rect 6740 16444 6741 16484
rect 6699 16435 6741 16444
rect 6699 15560 6741 15569
rect 6699 15520 6700 15560
rect 6740 15520 6741 15560
rect 6699 15511 6741 15520
rect 6700 15317 6740 15511
rect 6796 15392 6836 18283
rect 6892 17837 6932 18544
rect 6988 18416 7028 20392
rect 7084 19928 7124 20476
rect 7180 19928 7220 20896
rect 7276 20516 7316 21316
rect 7371 21307 7413 21316
rect 7372 21222 7412 21307
rect 7468 21188 7508 22408
rect 7564 21776 7604 22651
rect 7564 21727 7604 21736
rect 7660 21533 7700 22828
rect 7756 21608 7796 23155
rect 7851 23120 7893 23129
rect 7851 23080 7852 23120
rect 7892 23080 7893 23120
rect 7851 23071 7893 23080
rect 7948 23120 7988 23129
rect 7852 22986 7892 23071
rect 7851 22616 7893 22625
rect 7851 22576 7852 22616
rect 7892 22576 7893 22616
rect 7851 22567 7893 22576
rect 7852 21944 7892 22567
rect 7948 22121 7988 23080
rect 8043 23120 8085 23129
rect 8043 23080 8044 23120
rect 8084 23080 8085 23120
rect 8043 23071 8085 23080
rect 8140 23120 8180 23239
rect 8140 23071 8180 23080
rect 8044 22709 8084 23071
rect 8139 22952 8181 22961
rect 8139 22912 8140 22952
rect 8180 22912 8181 22952
rect 8139 22903 8181 22912
rect 8043 22700 8085 22709
rect 8043 22660 8044 22700
rect 8084 22660 8085 22700
rect 8043 22651 8085 22660
rect 8044 22280 8084 22651
rect 8044 22231 8084 22240
rect 8140 22280 8180 22903
rect 7947 22112 7989 22121
rect 7947 22072 7948 22112
rect 7988 22072 7989 22112
rect 7947 22063 7989 22072
rect 7852 21904 8084 21944
rect 7659 21524 7701 21533
rect 7659 21484 7660 21524
rect 7700 21484 7701 21524
rect 7659 21475 7701 21484
rect 7659 21356 7701 21365
rect 7659 21316 7660 21356
rect 7700 21316 7701 21356
rect 7659 21307 7701 21316
rect 7468 21148 7604 21188
rect 7372 20936 7412 20945
rect 7372 20600 7412 20896
rect 7564 20768 7604 21148
rect 7564 20719 7604 20728
rect 7660 20768 7700 21307
rect 7660 20719 7700 20728
rect 7372 20560 7604 20600
rect 7276 20476 7508 20516
rect 7276 20096 7316 20105
rect 7371 20096 7413 20105
rect 7316 20056 7372 20096
rect 7412 20056 7413 20096
rect 7276 20047 7316 20056
rect 7371 20047 7413 20056
rect 7468 20096 7508 20476
rect 7468 20047 7508 20056
rect 7564 20096 7604 20560
rect 7756 20348 7796 21568
rect 7851 21608 7893 21617
rect 7851 21568 7852 21608
rect 7892 21568 7893 21608
rect 7851 21559 7893 21568
rect 7852 21020 7892 21559
rect 7852 20971 7892 20980
rect 7564 20047 7604 20056
rect 7660 20308 7796 20348
rect 7852 20768 7892 20777
rect 7276 19928 7316 19937
rect 7180 19888 7276 19928
rect 7084 19879 7124 19888
rect 7276 19879 7316 19888
rect 7084 18752 7124 18761
rect 7372 18752 7412 20047
rect 7660 19769 7700 20308
rect 7852 20264 7892 20728
rect 7852 20215 7892 20224
rect 7755 20096 7797 20105
rect 7755 20056 7756 20096
rect 7796 20056 7797 20096
rect 7755 20047 7797 20056
rect 7756 19962 7796 20047
rect 7659 19760 7701 19769
rect 7659 19720 7660 19760
rect 7700 19720 7701 19760
rect 7659 19711 7701 19720
rect 8044 19340 8084 21904
rect 8140 20693 8180 22240
rect 8139 20684 8181 20693
rect 8139 20644 8140 20684
rect 8180 20644 8181 20684
rect 8139 20635 8181 20644
rect 8236 19424 8276 23500
rect 8332 20180 8372 24088
rect 8428 23717 8468 25759
rect 8427 23708 8469 23717
rect 8427 23668 8428 23708
rect 8468 23668 8469 23708
rect 8427 23659 8469 23668
rect 8524 22616 8564 25936
rect 8428 22576 8564 22616
rect 8428 20441 8468 22576
rect 8716 22457 8756 27355
rect 8812 27354 8852 27439
rect 8908 27404 8948 28867
rect 9003 28412 9045 28421
rect 9003 28372 9004 28412
rect 9044 28372 9045 28412
rect 9003 28363 9045 28372
rect 9004 28342 9044 28363
rect 9004 27656 9044 28302
rect 9100 27740 9140 29800
rect 9196 29791 9236 29800
rect 9388 29840 9428 29959
rect 9484 29849 9524 31312
rect 9388 29791 9428 29800
rect 9483 29840 9525 29849
rect 9483 29800 9484 29840
rect 9524 29800 9525 29840
rect 9483 29791 9525 29800
rect 9484 29706 9524 29791
rect 9580 29765 9620 32311
rect 9579 29756 9621 29765
rect 9579 29716 9580 29756
rect 9620 29716 9621 29756
rect 9579 29707 9621 29716
rect 9195 29672 9237 29681
rect 9195 29632 9196 29672
rect 9236 29632 9237 29672
rect 9195 29623 9237 29632
rect 9292 29672 9332 29681
rect 9196 28421 9236 29623
rect 9292 29177 9332 29632
rect 9676 29588 9716 32647
rect 9963 32444 10005 32453
rect 9963 32404 9964 32444
rect 10004 32404 10005 32444
rect 9963 32395 10005 32404
rect 9964 32192 10004 32395
rect 10004 32152 10292 32192
rect 9964 32143 10004 32152
rect 10156 31940 10196 31949
rect 9964 31900 10156 31940
rect 9964 31436 10004 31900
rect 10156 31891 10196 31900
rect 9916 31396 10004 31436
rect 9916 31394 9956 31396
rect 9916 31345 9956 31354
rect 10060 31184 10100 31193
rect 9771 30764 9813 30773
rect 9771 30724 9772 30764
rect 9812 30724 9813 30764
rect 9771 30715 9813 30724
rect 9580 29548 9716 29588
rect 9291 29168 9333 29177
rect 9291 29128 9292 29168
rect 9332 29128 9333 29168
rect 9291 29119 9333 29128
rect 9291 29000 9333 29009
rect 9291 28960 9292 29000
rect 9332 28960 9333 29000
rect 9291 28951 9333 28960
rect 9195 28412 9237 28421
rect 9195 28372 9196 28412
rect 9236 28372 9237 28412
rect 9195 28363 9237 28372
rect 9195 28244 9237 28253
rect 9195 28204 9196 28244
rect 9236 28204 9237 28244
rect 9195 28195 9237 28204
rect 9196 28110 9236 28195
rect 9195 27992 9237 28001
rect 9195 27952 9196 27992
rect 9236 27952 9237 27992
rect 9195 27943 9237 27952
rect 9100 27691 9140 27700
rect 9004 27581 9044 27616
rect 9003 27572 9045 27581
rect 9003 27532 9004 27572
rect 9044 27532 9045 27572
rect 9003 27523 9045 27532
rect 9004 27492 9044 27523
rect 8908 27364 9044 27404
rect 8811 27236 8853 27245
rect 8811 27196 8812 27236
rect 8852 27196 8853 27236
rect 8811 27187 8853 27196
rect 8812 25565 8852 27187
rect 8907 26816 8949 26825
rect 8907 26776 8908 26816
rect 8948 26776 8949 26816
rect 8907 26767 8949 26776
rect 9004 26816 9044 27364
rect 8908 26144 8948 26767
rect 9004 26321 9044 26776
rect 9099 26396 9141 26405
rect 9099 26356 9100 26396
rect 9140 26356 9141 26396
rect 9099 26347 9141 26356
rect 9003 26312 9045 26321
rect 9003 26272 9004 26312
rect 9044 26272 9045 26312
rect 9003 26263 9045 26272
rect 8908 26095 8948 26104
rect 9004 26144 9044 26153
rect 9100 26144 9140 26347
rect 9196 26228 9236 27943
rect 9292 26405 9332 28951
rect 9484 28916 9524 28925
rect 9387 28580 9429 28589
rect 9387 28540 9388 28580
rect 9428 28540 9429 28580
rect 9387 28531 9429 28540
rect 9388 28076 9428 28531
rect 9484 28328 9524 28876
rect 9580 28589 9620 29548
rect 9676 29177 9716 29262
rect 9675 29168 9717 29177
rect 9675 29128 9676 29168
rect 9716 29128 9717 29168
rect 9675 29119 9717 29128
rect 9772 29093 9812 30715
rect 10060 30008 10100 31144
rect 10252 30773 10292 32152
rect 10636 32117 10676 32992
rect 10635 32108 10677 32117
rect 10635 32068 10636 32108
rect 10676 32068 10677 32108
rect 10635 32059 10677 32068
rect 10444 31352 10484 31361
rect 10444 30848 10484 31312
rect 10540 31352 10580 31361
rect 10540 31025 10580 31312
rect 10539 31016 10581 31025
rect 10539 30976 10540 31016
rect 10580 30976 10581 31016
rect 10539 30967 10581 30976
rect 10444 30799 10484 30808
rect 10251 30764 10293 30773
rect 10251 30724 10252 30764
rect 10292 30724 10293 30764
rect 10251 30715 10293 30724
rect 10252 30680 10292 30715
rect 10252 30630 10292 30640
rect 10443 30344 10485 30353
rect 10443 30304 10444 30344
rect 10484 30304 10485 30344
rect 10443 30295 10485 30304
rect 10347 30176 10389 30185
rect 10347 30136 10348 30176
rect 10388 30136 10389 30176
rect 10347 30127 10389 30136
rect 9964 29968 10100 30008
rect 9867 29840 9909 29849
rect 9867 29800 9868 29840
rect 9908 29800 9909 29840
rect 9867 29791 9909 29800
rect 9771 29084 9813 29093
rect 9771 29044 9772 29084
rect 9812 29044 9813 29084
rect 9771 29035 9813 29044
rect 9579 28580 9621 28589
rect 9579 28540 9580 28580
rect 9620 28540 9621 28580
rect 9579 28531 9621 28540
rect 9484 28253 9524 28288
rect 9580 28328 9620 28337
rect 9483 28244 9525 28253
rect 9483 28204 9484 28244
rect 9524 28204 9525 28244
rect 9483 28195 9525 28204
rect 9580 28085 9620 28288
rect 9675 28328 9717 28337
rect 9675 28288 9676 28328
rect 9716 28288 9717 28328
rect 9675 28279 9717 28288
rect 9579 28076 9621 28085
rect 9388 28036 9524 28076
rect 9388 27645 9428 27654
rect 9388 27581 9428 27605
rect 9387 27572 9429 27581
rect 9387 27532 9388 27572
rect 9428 27532 9429 27572
rect 9387 27523 9429 27532
rect 9388 27510 9428 27523
rect 9387 27404 9429 27413
rect 9387 27364 9388 27404
rect 9428 27364 9429 27404
rect 9387 27355 9429 27364
rect 9388 27270 9428 27355
rect 9291 26396 9333 26405
rect 9291 26356 9292 26396
rect 9332 26356 9333 26396
rect 9291 26347 9333 26356
rect 9484 26228 9524 28036
rect 9579 28036 9580 28076
rect 9620 28036 9621 28076
rect 9579 28027 9621 28036
rect 9580 27749 9620 27780
rect 9579 27740 9621 27749
rect 9579 27700 9580 27740
rect 9620 27700 9621 27740
rect 9579 27691 9621 27700
rect 9580 27656 9620 27691
rect 9580 26825 9620 27616
rect 9676 27656 9716 28279
rect 9771 27740 9813 27749
rect 9771 27700 9772 27740
rect 9812 27700 9813 27740
rect 9771 27691 9813 27700
rect 9676 27581 9716 27616
rect 9675 27572 9717 27581
rect 9675 27532 9676 27572
rect 9716 27532 9717 27572
rect 9675 27523 9717 27532
rect 9579 26816 9621 26825
rect 9579 26776 9580 26816
rect 9620 26776 9621 26816
rect 9579 26767 9621 26776
rect 9196 26188 9332 26228
rect 9044 26104 9236 26144
rect 9004 26095 9044 26104
rect 8811 25556 8853 25565
rect 8811 25516 8812 25556
rect 8852 25516 8853 25556
rect 8811 25507 8853 25516
rect 8907 25388 8949 25397
rect 8907 25348 8908 25388
rect 8948 25348 8949 25388
rect 8907 25339 8949 25348
rect 8908 25304 8948 25339
rect 8811 24548 8853 24557
rect 8811 24508 8812 24548
rect 8852 24508 8853 24548
rect 8811 24499 8853 24508
rect 8520 22448 8562 22457
rect 8715 22448 8757 22457
rect 8520 22408 8521 22448
rect 8561 22408 8564 22448
rect 8520 22399 8564 22408
rect 8715 22408 8716 22448
rect 8756 22408 8757 22448
rect 8715 22399 8757 22408
rect 8524 22364 8564 22399
rect 8524 22315 8564 22324
rect 8620 22289 8660 22374
rect 8619 22280 8661 22289
rect 8619 22240 8620 22280
rect 8660 22240 8661 22280
rect 8619 22231 8661 22240
rect 8619 22112 8661 22121
rect 8619 22072 8620 22112
rect 8660 22072 8661 22112
rect 8619 22063 8661 22072
rect 8427 20432 8469 20441
rect 8427 20392 8428 20432
rect 8468 20392 8469 20432
rect 8427 20383 8469 20392
rect 8332 20140 8564 20180
rect 8236 19384 8468 19424
rect 7852 19300 8084 19340
rect 7467 19256 7509 19265
rect 7467 19216 7468 19256
rect 7508 19216 7509 19256
rect 7467 19207 7509 19216
rect 7756 19256 7796 19265
rect 7124 18712 7412 18752
rect 7084 18703 7124 18712
rect 6988 18376 7316 18416
rect 6891 17828 6933 17837
rect 6891 17788 6892 17828
rect 6932 17788 6933 17828
rect 6891 17779 6933 17788
rect 7180 17744 7220 17753
rect 6892 17660 6932 17669
rect 7180 17660 7220 17704
rect 6932 17620 7220 17660
rect 7276 17744 7316 18376
rect 6892 17611 6932 17620
rect 6987 17492 7029 17501
rect 6987 17452 6988 17492
rect 7028 17452 7029 17492
rect 6987 17443 7029 17452
rect 6891 15644 6933 15653
rect 6891 15604 6892 15644
rect 6932 15604 6933 15644
rect 6891 15595 6933 15604
rect 6892 15510 6932 15595
rect 6988 15476 7028 17443
rect 7276 17249 7316 17704
rect 7468 17669 7508 19207
rect 7756 18593 7796 19216
rect 7755 18584 7797 18593
rect 7755 18544 7756 18584
rect 7796 18544 7797 18584
rect 7755 18535 7797 18544
rect 7659 18500 7701 18509
rect 7659 18460 7660 18500
rect 7700 18460 7701 18500
rect 7659 18451 7701 18460
rect 7660 17828 7700 18451
rect 7660 17779 7700 17788
rect 7756 17744 7796 17753
rect 7467 17660 7509 17669
rect 7467 17620 7468 17660
rect 7508 17620 7509 17660
rect 7467 17611 7509 17620
rect 7756 17585 7796 17704
rect 7755 17576 7797 17585
rect 7755 17536 7756 17576
rect 7796 17536 7797 17576
rect 7755 17527 7797 17536
rect 7275 17240 7317 17249
rect 7275 17200 7276 17240
rect 7316 17200 7317 17240
rect 7275 17191 7317 17200
rect 7467 16652 7509 16661
rect 7467 16612 7468 16652
rect 7508 16612 7509 16652
rect 7467 16603 7509 16612
rect 7371 16400 7413 16409
rect 7371 16360 7372 16400
rect 7412 16360 7413 16400
rect 7371 16351 7413 16360
rect 7372 16232 7412 16351
rect 7180 15653 7220 15675
rect 7179 15644 7221 15653
rect 7179 15604 7180 15644
rect 7220 15604 7221 15644
rect 7179 15595 7221 15604
rect 7180 15580 7220 15595
rect 7180 15531 7220 15540
rect 7275 15560 7317 15569
rect 7275 15520 7276 15560
rect 7316 15520 7317 15560
rect 7275 15511 7317 15520
rect 6988 15436 7220 15476
rect 6796 15352 7124 15392
rect 6699 15308 6741 15317
rect 6699 15268 6700 15308
rect 6740 15268 6741 15308
rect 6699 15259 6741 15268
rect 6891 15140 6933 15149
rect 6891 15100 6892 15140
rect 6932 15100 6933 15140
rect 6891 15091 6933 15100
rect 6603 14384 6645 14393
rect 6603 14344 6604 14384
rect 6644 14344 6645 14384
rect 6603 14335 6645 14344
rect 6220 14176 6356 14216
rect 6220 13880 6260 14176
rect 6508 14132 6548 14141
rect 6548 14092 6644 14132
rect 6508 14083 6548 14092
rect 6316 14048 6356 14057
rect 6316 13964 6356 14008
rect 6604 14043 6644 14092
rect 6892 14057 6932 15091
rect 6796 14048 6836 14057
rect 6604 14008 6796 14043
rect 6604 14003 6836 14008
rect 6796 13999 6836 14003
rect 6891 14048 6933 14057
rect 6891 14008 6892 14048
rect 6932 14008 6933 14048
rect 6891 13999 6933 14008
rect 6411 13964 6453 13973
rect 6316 13924 6412 13964
rect 6452 13924 6453 13964
rect 6411 13915 6453 13924
rect 6892 13914 6932 13999
rect 6220 13840 6356 13880
rect 6316 11864 6356 13840
rect 7084 13796 7124 15352
rect 6892 13756 7124 13796
rect 6892 13124 6932 13756
rect 6988 13208 7028 13217
rect 6988 13124 7028 13168
rect 6892 13084 7028 13124
rect 6411 12956 6453 12965
rect 6411 12916 6412 12956
rect 6452 12916 6453 12956
rect 6411 12907 6453 12916
rect 6220 11824 6356 11864
rect 6123 11108 6165 11117
rect 6123 11068 6124 11108
rect 6164 11068 6165 11108
rect 6123 11059 6165 11068
rect 6220 11033 6260 11824
rect 6315 11696 6357 11705
rect 6315 11656 6316 11696
rect 6356 11656 6357 11696
rect 6315 11647 6357 11656
rect 6316 11562 6356 11647
rect 6219 11024 6261 11033
rect 6219 10984 6220 11024
rect 6260 10984 6261 11024
rect 6219 10975 6261 10984
rect 6123 10940 6165 10949
rect 6123 10900 6124 10940
rect 6164 10900 6165 10940
rect 6123 10891 6165 10900
rect 6124 10806 6164 10891
rect 6220 10890 6260 10975
rect 6219 8840 6261 8849
rect 6219 8800 6220 8840
rect 6260 8800 6261 8840
rect 6219 8791 6261 8800
rect 6123 8168 6165 8177
rect 6123 8128 6124 8168
rect 6164 8128 6165 8168
rect 6123 8119 6165 8128
rect 6124 8000 6164 8119
rect 6124 7951 6164 7960
rect 6220 7328 6260 8791
rect 6220 7288 6356 7328
rect 6220 7160 6260 7169
rect 6124 6656 6164 6665
rect 6220 6656 6260 7120
rect 6316 7160 6356 7288
rect 6316 6749 6356 7120
rect 6315 6740 6357 6749
rect 6315 6700 6316 6740
rect 6356 6700 6357 6740
rect 6315 6691 6357 6700
rect 6164 6616 6260 6656
rect 6124 6607 6164 6616
rect 6316 6446 6356 6455
rect 6316 6245 6356 6406
rect 6315 6236 6357 6245
rect 6315 6196 6316 6236
rect 6356 6196 6357 6236
rect 6315 6187 6357 6196
rect 6028 6112 6260 6152
rect 5836 6028 6068 6068
rect 6028 5984 6068 6028
rect 6028 5944 6164 5984
rect 5931 5900 5973 5909
rect 5931 5860 5932 5900
rect 5972 5860 5973 5900
rect 5931 5851 5973 5860
rect 5740 5776 5876 5816
rect 5548 5188 5684 5228
rect 5740 5648 5780 5657
rect 5452 4962 5492 4971
rect 5452 3725 5492 4922
rect 5451 3716 5493 3725
rect 5451 3676 5452 3716
rect 5492 3676 5493 3716
rect 5451 3667 5493 3676
rect 5548 3632 5588 5188
rect 5644 5060 5684 5071
rect 5644 4985 5684 5020
rect 5643 4976 5685 4985
rect 5643 4936 5644 4976
rect 5684 4936 5685 4976
rect 5643 4927 5685 4936
rect 5643 4640 5685 4649
rect 5643 4600 5644 4640
rect 5684 4600 5685 4640
rect 5643 4591 5685 4600
rect 5644 4313 5684 4591
rect 5740 4397 5780 5608
rect 5836 5228 5876 5776
rect 5932 5766 5972 5851
rect 5836 5188 5972 5228
rect 5835 5060 5877 5069
rect 5835 5020 5836 5060
rect 5876 5020 5877 5060
rect 5835 5011 5877 5020
rect 5739 4388 5781 4397
rect 5739 4348 5740 4388
rect 5780 4348 5781 4388
rect 5739 4339 5781 4348
rect 5643 4304 5685 4313
rect 5643 4264 5644 4304
rect 5684 4264 5685 4304
rect 5643 4255 5685 4264
rect 5644 4136 5684 4255
rect 5644 4087 5684 4096
rect 5739 3716 5781 3725
rect 5739 3676 5740 3716
rect 5780 3676 5781 3716
rect 5739 3667 5781 3676
rect 5740 3632 5780 3667
rect 5548 3592 5684 3632
rect 5547 3464 5589 3473
rect 5547 3424 5548 3464
rect 5588 3424 5589 3464
rect 5547 3415 5589 3424
rect 5548 3330 5588 3415
rect 5644 2960 5684 3592
rect 5740 3581 5780 3592
rect 5644 2920 5780 2960
rect 5452 2633 5492 2718
rect 5547 2708 5589 2717
rect 5547 2668 5548 2708
rect 5588 2668 5589 2708
rect 5547 2659 5589 2668
rect 5451 2624 5493 2633
rect 5451 2584 5452 2624
rect 5492 2584 5493 2624
rect 5451 2575 5493 2584
rect 5548 2624 5588 2659
rect 5548 2465 5588 2584
rect 5643 2624 5685 2633
rect 5643 2584 5644 2624
rect 5684 2584 5685 2624
rect 5643 2575 5685 2584
rect 5547 2456 5589 2465
rect 5547 2416 5548 2456
rect 5588 2416 5589 2456
rect 5547 2407 5589 2416
rect 4876 1147 4916 1156
rect 5260 1240 5396 1280
rect 4492 1112 4532 1121
rect 4396 1072 4492 1112
rect 4299 1063 4341 1072
rect 4492 1063 4532 1072
rect 5067 1112 5109 1121
rect 5067 1072 5068 1112
rect 5108 1072 5109 1112
rect 5067 1063 5109 1072
rect 4203 440 4245 449
rect 4203 400 4204 440
rect 4244 400 4245 440
rect 4203 391 4245 400
rect 4300 80 4340 1063
rect 4491 944 4533 953
rect 4491 904 4492 944
rect 4532 904 4533 944
rect 4491 895 4533 904
rect 5068 944 5108 1063
rect 5260 953 5300 1240
rect 5356 1112 5396 1121
rect 5068 895 5108 904
rect 5259 944 5301 953
rect 5259 904 5260 944
rect 5300 904 5301 944
rect 5259 895 5301 904
rect 4492 80 4532 895
rect 5356 785 5396 1072
rect 4928 776 5296 785
rect 4968 736 5010 776
rect 5050 736 5092 776
rect 5132 736 5174 776
rect 5214 736 5256 776
rect 4928 727 5296 736
rect 5355 776 5397 785
rect 5355 736 5356 776
rect 5396 736 5397 776
rect 5355 727 5397 736
rect 5451 692 5493 701
rect 5451 652 5452 692
rect 5492 652 5493 692
rect 5451 643 5493 652
rect 5067 608 5109 617
rect 5067 568 5068 608
rect 5108 568 5109 608
rect 5067 559 5109 568
rect 4683 440 4725 449
rect 4683 400 4684 440
rect 4724 400 4725 440
rect 4683 391 4725 400
rect 4684 80 4724 391
rect 4875 272 4917 281
rect 4875 232 4876 272
rect 4916 232 4917 272
rect 4875 223 4917 232
rect 4876 80 4916 223
rect 5068 80 5108 559
rect 5259 272 5301 281
rect 5259 232 5260 272
rect 5300 232 5301 272
rect 5259 223 5301 232
rect 5260 80 5300 223
rect 5452 80 5492 643
rect 5644 80 5684 2575
rect 5740 2540 5780 2920
rect 5836 2717 5876 5011
rect 5932 4649 5972 5188
rect 6124 5069 6164 5944
rect 6123 5060 6165 5069
rect 6123 5020 6124 5060
rect 6164 5020 6165 5060
rect 6123 5011 6165 5020
rect 6028 4976 6068 4985
rect 5931 4640 5973 4649
rect 5931 4600 5932 4640
rect 5972 4600 5973 4640
rect 5931 4591 5973 4600
rect 5931 4304 5973 4313
rect 5931 4264 5932 4304
rect 5972 4264 5973 4304
rect 5931 4255 5973 4264
rect 5932 3296 5972 4255
rect 6028 3716 6068 4936
rect 6124 4976 6164 5011
rect 6124 4926 6164 4936
rect 6028 3676 6164 3716
rect 6027 3548 6069 3557
rect 6027 3508 6028 3548
rect 6068 3508 6069 3548
rect 6027 3499 6069 3508
rect 6028 3464 6068 3499
rect 6028 3413 6068 3424
rect 5932 3256 6068 3296
rect 5931 2876 5973 2885
rect 5931 2836 5932 2876
rect 5972 2836 5973 2876
rect 5931 2827 5973 2836
rect 5835 2708 5877 2717
rect 5835 2668 5836 2708
rect 5876 2668 5877 2708
rect 5835 2659 5877 2668
rect 5932 2708 5972 2827
rect 5932 2633 5972 2668
rect 6028 2708 6068 3256
rect 6028 2659 6068 2668
rect 5931 2624 5973 2633
rect 5931 2584 5932 2624
rect 5972 2584 5973 2624
rect 5931 2575 5973 2584
rect 5932 2544 5972 2575
rect 5740 2500 5876 2540
rect 5836 80 5876 2500
rect 6124 2120 6164 3676
rect 6124 2071 6164 2080
rect 5932 1952 5972 1961
rect 5932 1457 5972 1912
rect 5931 1448 5973 1457
rect 5931 1408 5932 1448
rect 5972 1408 5973 1448
rect 5931 1399 5973 1408
rect 6027 272 6069 281
rect 6027 232 6028 272
rect 6068 232 6069 272
rect 6027 223 6069 232
rect 6028 80 6068 223
rect 6220 80 6260 6112
rect 6412 3473 6452 12907
rect 6796 11696 6836 11705
rect 6508 11612 6548 11621
rect 6796 11612 6836 11656
rect 6548 11572 6836 11612
rect 6892 11696 6932 11705
rect 6508 11563 6548 11572
rect 6892 11528 6932 11656
rect 6796 11488 6932 11528
rect 6699 11360 6741 11369
rect 6699 11320 6700 11360
rect 6740 11320 6741 11360
rect 6699 11311 6741 11320
rect 6700 11024 6740 11311
rect 6700 10975 6740 10984
rect 6796 10949 6836 11488
rect 6891 11024 6933 11033
rect 6891 10984 6892 11024
rect 6932 10984 6933 11024
rect 6891 10975 6933 10984
rect 6795 10940 6837 10949
rect 6795 10900 6796 10940
rect 6836 10900 6837 10940
rect 6795 10891 6837 10900
rect 6603 10604 6645 10613
rect 6603 10564 6604 10604
rect 6644 10564 6645 10604
rect 6603 10555 6645 10564
rect 6604 7505 6644 10555
rect 6796 10352 6836 10891
rect 6700 10312 6836 10352
rect 6603 7496 6645 7505
rect 6603 7456 6604 7496
rect 6644 7456 6645 7496
rect 6603 7447 6645 7456
rect 6700 7244 6740 10312
rect 6795 10184 6837 10193
rect 6795 10144 6796 10184
rect 6836 10144 6837 10184
rect 6795 10135 6837 10144
rect 6796 10050 6836 10135
rect 6892 8840 6932 10975
rect 6988 10613 7028 13084
rect 7180 11108 7220 15436
rect 7276 15426 7316 15511
rect 7372 15485 7412 16192
rect 7371 15476 7413 15485
rect 7371 15436 7372 15476
rect 7412 15436 7413 15476
rect 7371 15427 7413 15436
rect 7275 14720 7317 14729
rect 7275 14680 7276 14720
rect 7316 14680 7317 14720
rect 7275 14671 7317 14680
rect 7276 14048 7316 14671
rect 7371 14132 7413 14141
rect 7371 14092 7372 14132
rect 7412 14092 7413 14132
rect 7371 14083 7413 14092
rect 7276 13999 7316 14008
rect 7372 14048 7412 14083
rect 7372 13997 7412 14008
rect 7468 12704 7508 16603
rect 7755 15560 7797 15569
rect 7755 15520 7756 15560
rect 7796 15520 7797 15560
rect 7755 15511 7797 15520
rect 7660 15476 7700 15485
rect 7660 15149 7700 15436
rect 7756 15426 7796 15511
rect 7755 15308 7797 15317
rect 7755 15268 7756 15308
rect 7796 15268 7797 15308
rect 7755 15259 7797 15268
rect 7659 15140 7701 15149
rect 7659 15100 7660 15140
rect 7700 15100 7701 15140
rect 7659 15091 7701 15100
rect 7756 14720 7796 15259
rect 7756 14671 7796 14680
rect 7852 14216 7892 19300
rect 8236 19256 8276 19264
rect 8140 19255 8276 19256
rect 8140 19216 8236 19255
rect 7948 19172 7988 19181
rect 8140 19172 8180 19216
rect 8236 19206 8276 19215
rect 8332 19256 8372 19267
rect 8332 19181 8372 19216
rect 7988 19132 8180 19172
rect 8331 19172 8373 19181
rect 8331 19132 8332 19172
rect 8372 19132 8373 19172
rect 7948 19123 7988 19132
rect 8331 19123 8373 19132
rect 8428 18761 8468 19384
rect 8427 18752 8469 18761
rect 8427 18712 8428 18752
rect 8468 18712 8469 18752
rect 8427 18703 8469 18712
rect 8428 18584 8468 18593
rect 8428 18425 8468 18544
rect 8139 18416 8181 18425
rect 8139 18376 8140 18416
rect 8180 18376 8181 18416
rect 8139 18367 8181 18376
rect 8427 18416 8469 18425
rect 8427 18376 8428 18416
rect 8468 18376 8469 18416
rect 8427 18367 8469 18376
rect 7947 14972 7989 14981
rect 7947 14932 7948 14972
rect 7988 14932 7989 14972
rect 7947 14923 7989 14932
rect 7948 14838 7988 14923
rect 8140 14720 8180 18367
rect 8524 18248 8564 20140
rect 8332 18208 8564 18248
rect 8236 17744 8276 17753
rect 8332 17744 8372 18208
rect 8276 17704 8372 17744
rect 8523 17744 8565 17753
rect 8523 17704 8524 17744
rect 8564 17704 8565 17744
rect 8236 15980 8276 17704
rect 8523 17695 8565 17704
rect 8331 17156 8373 17165
rect 8331 17116 8332 17156
rect 8372 17116 8373 17156
rect 8331 17107 8373 17116
rect 8332 17072 8372 17107
rect 8332 17021 8372 17032
rect 8236 15940 8372 15980
rect 8236 15560 8276 15569
rect 8236 14729 8276 15520
rect 8044 14680 8140 14720
rect 7852 14176 7988 14216
rect 7851 14048 7893 14057
rect 7851 14008 7852 14048
rect 7892 14008 7893 14048
rect 7851 13999 7893 14008
rect 7755 13796 7797 13805
rect 7755 13756 7756 13796
rect 7796 13756 7797 13796
rect 7755 13747 7797 13756
rect 7659 13712 7701 13721
rect 7659 13672 7660 13712
rect 7700 13672 7701 13712
rect 7659 13663 7701 13672
rect 7276 12664 7508 12704
rect 7276 11780 7316 12664
rect 7468 12494 7508 12503
rect 7508 12454 7604 12494
rect 7468 12445 7508 12454
rect 7564 12209 7604 12454
rect 7563 12200 7605 12209
rect 7563 12160 7564 12200
rect 7604 12160 7605 12200
rect 7563 12151 7605 12160
rect 7276 11369 7316 11740
rect 7372 11696 7412 11705
rect 7372 11537 7412 11656
rect 7371 11528 7413 11537
rect 7371 11488 7372 11528
rect 7412 11488 7413 11528
rect 7371 11479 7413 11488
rect 7275 11360 7317 11369
rect 7275 11320 7276 11360
rect 7316 11320 7317 11360
rect 7275 11311 7317 11320
rect 7467 11360 7509 11369
rect 7467 11320 7468 11360
rect 7508 11320 7509 11360
rect 7467 11311 7509 11320
rect 7371 11192 7413 11201
rect 7371 11152 7372 11192
rect 7412 11152 7413 11192
rect 7371 11143 7413 11152
rect 7180 11068 7316 11108
rect 7180 11010 7220 11019
rect 6987 10604 7029 10613
rect 6987 10564 6988 10604
rect 7028 10564 7029 10604
rect 6987 10555 7029 10564
rect 6988 10361 7028 10446
rect 7180 10361 7220 10970
rect 6987 10352 7029 10361
rect 6987 10312 6988 10352
rect 7028 10312 7029 10352
rect 6987 10303 7029 10312
rect 7179 10352 7221 10361
rect 7179 10312 7180 10352
rect 7220 10312 7221 10352
rect 7179 10303 7221 10312
rect 6987 10184 7029 10193
rect 6987 10144 6988 10184
rect 7028 10144 7029 10184
rect 6987 10135 7029 10144
rect 7179 10184 7221 10193
rect 7179 10144 7180 10184
rect 7220 10144 7221 10184
rect 7179 10135 7221 10144
rect 6508 7204 6700 7244
rect 6508 4976 6548 7204
rect 6700 7195 6740 7204
rect 6796 8800 6932 8840
rect 6796 7244 6836 8800
rect 6892 8672 6932 8681
rect 6892 8513 6932 8632
rect 6891 8504 6933 8513
rect 6891 8464 6892 8504
rect 6932 8464 6933 8504
rect 6891 8455 6933 8464
rect 6891 7496 6933 7505
rect 6891 7456 6892 7496
rect 6932 7456 6933 7496
rect 6891 7447 6933 7456
rect 6796 6824 6836 7204
rect 6411 3464 6453 3473
rect 6411 3424 6412 3464
rect 6452 3424 6453 3464
rect 6411 3415 6453 3424
rect 6508 2885 6548 4936
rect 6604 6784 6836 6824
rect 6604 4976 6644 6784
rect 6892 6245 6932 7447
rect 6891 6236 6933 6245
rect 6891 6196 6892 6236
rect 6932 6196 6933 6236
rect 6891 6187 6933 6196
rect 6699 6068 6741 6077
rect 6699 6028 6700 6068
rect 6740 6028 6741 6068
rect 6699 6019 6741 6028
rect 6700 5648 6740 6019
rect 6740 5608 6836 5648
rect 6700 5599 6740 5608
rect 6604 4313 6644 4936
rect 6699 4976 6741 4985
rect 6699 4936 6700 4976
rect 6740 4936 6741 4976
rect 6699 4927 6741 4936
rect 6603 4304 6645 4313
rect 6603 4264 6604 4304
rect 6644 4264 6645 4304
rect 6603 4255 6645 4264
rect 6507 2876 6549 2885
rect 6507 2836 6508 2876
rect 6548 2836 6549 2876
rect 6507 2827 6549 2836
rect 6508 2624 6548 2633
rect 6700 2624 6740 4927
rect 6796 3557 6836 5608
rect 6892 4136 6932 4145
rect 6988 4136 7028 10135
rect 7180 10050 7220 10135
rect 7179 9764 7221 9773
rect 7179 9724 7180 9764
rect 7220 9724 7221 9764
rect 7179 9715 7221 9724
rect 7180 9680 7220 9715
rect 7180 9629 7220 9640
rect 7276 9092 7316 11068
rect 7372 11058 7412 11143
rect 7180 9052 7316 9092
rect 7372 9498 7412 9507
rect 7083 8840 7125 8849
rect 7083 8800 7084 8840
rect 7124 8800 7125 8840
rect 7083 8791 7125 8800
rect 7084 8706 7124 8791
rect 7083 4976 7125 4985
rect 7083 4936 7084 4976
rect 7124 4936 7125 4976
rect 7083 4927 7125 4936
rect 7084 4842 7124 4927
rect 7083 4388 7125 4397
rect 7083 4348 7084 4388
rect 7124 4348 7125 4388
rect 7083 4339 7125 4348
rect 7084 4254 7124 4339
rect 7180 4150 7220 9052
rect 7276 8924 7316 8933
rect 7372 8924 7412 9458
rect 7316 8884 7412 8924
rect 7276 8875 7316 8884
rect 7468 8840 7508 11311
rect 7372 8800 7508 8840
rect 7564 11024 7604 11033
rect 7660 11024 7700 13663
rect 7604 10984 7700 11024
rect 7372 8168 7412 8800
rect 7468 8672 7508 8681
rect 7468 8513 7508 8632
rect 7467 8504 7509 8513
rect 7467 8464 7468 8504
rect 7508 8464 7509 8504
rect 7467 8455 7509 8464
rect 7276 8128 7412 8168
rect 7276 7160 7316 8128
rect 7371 8000 7413 8009
rect 7371 7960 7372 8000
rect 7412 7960 7413 8000
rect 7371 7951 7413 7960
rect 7276 4985 7316 7120
rect 7372 5909 7412 7951
rect 7564 7916 7604 10984
rect 7756 8168 7796 13747
rect 7852 12032 7892 13999
rect 7948 12209 7988 14176
rect 8044 13805 8084 14680
rect 8140 14671 8180 14680
rect 8235 14720 8277 14729
rect 8235 14680 8236 14720
rect 8276 14680 8277 14720
rect 8235 14671 8277 14680
rect 8332 14645 8372 15940
rect 8331 14636 8373 14645
rect 8331 14596 8332 14636
rect 8372 14596 8373 14636
rect 8331 14587 8373 14596
rect 8139 14468 8181 14477
rect 8139 14428 8140 14468
rect 8180 14428 8181 14468
rect 8139 14419 8181 14428
rect 8043 13796 8085 13805
rect 8043 13756 8044 13796
rect 8084 13756 8085 13796
rect 8043 13747 8085 13756
rect 7947 12200 7989 12209
rect 7947 12160 7948 12200
rect 7988 12160 7989 12200
rect 7947 12151 7989 12160
rect 7852 11992 7988 12032
rect 7851 11696 7893 11705
rect 7851 11656 7852 11696
rect 7892 11656 7893 11696
rect 7851 11647 7893 11656
rect 7852 11562 7892 11647
rect 7851 9680 7893 9689
rect 7851 9640 7852 9680
rect 7892 9640 7893 9680
rect 7851 9631 7893 9640
rect 7852 9521 7892 9631
rect 7851 9512 7893 9521
rect 7851 9472 7852 9512
rect 7892 9472 7893 9512
rect 7851 9463 7893 9472
rect 7852 9378 7892 9463
rect 7851 8756 7893 8765
rect 7851 8716 7852 8756
rect 7892 8716 7893 8756
rect 7851 8707 7893 8716
rect 7468 7876 7604 7916
rect 7660 8128 7796 8168
rect 7468 6245 7508 7876
rect 7563 7748 7605 7757
rect 7563 7708 7564 7748
rect 7604 7708 7605 7748
rect 7563 7699 7605 7708
rect 7564 7614 7604 7699
rect 7563 7496 7605 7505
rect 7563 7456 7564 7496
rect 7604 7456 7605 7496
rect 7563 7447 7605 7456
rect 7564 6497 7604 7447
rect 7563 6488 7605 6497
rect 7563 6448 7564 6488
rect 7604 6448 7605 6488
rect 7563 6439 7605 6448
rect 7467 6236 7509 6245
rect 7467 6196 7468 6236
rect 7508 6196 7509 6236
rect 7467 6187 7509 6196
rect 7371 5900 7413 5909
rect 7371 5860 7372 5900
rect 7412 5860 7413 5900
rect 7371 5851 7413 5860
rect 7564 5657 7604 6439
rect 7563 5648 7605 5657
rect 7563 5608 7564 5648
rect 7604 5608 7605 5648
rect 7563 5599 7605 5608
rect 7467 5060 7509 5069
rect 7467 5020 7468 5060
rect 7508 5020 7509 5060
rect 7467 5011 7509 5020
rect 7275 4976 7317 4985
rect 7275 4936 7276 4976
rect 7316 4936 7317 4976
rect 7275 4927 7317 4936
rect 6932 4096 7028 4136
rect 7084 4110 7220 4150
rect 7372 4136 7412 4145
rect 6795 3548 6837 3557
rect 6795 3508 6796 3548
rect 6836 3508 6837 3548
rect 6795 3499 6837 3508
rect 6548 2584 6740 2624
rect 6508 2575 6548 2584
rect 6892 2540 6932 4096
rect 6604 2500 6932 2540
rect 6988 2629 7028 2638
rect 6411 2372 6453 2381
rect 6411 2332 6412 2372
rect 6452 2332 6453 2372
rect 6411 2323 6453 2332
rect 6412 1952 6452 2323
rect 6412 1903 6452 1912
rect 6604 1457 6644 2500
rect 6988 1700 7028 2589
rect 6796 1660 7028 1700
rect 6603 1448 6645 1457
rect 6603 1408 6604 1448
rect 6644 1408 6645 1448
rect 6603 1399 6645 1408
rect 6411 1280 6453 1289
rect 6411 1240 6412 1280
rect 6452 1240 6453 1280
rect 6411 1231 6453 1240
rect 6412 80 6452 1231
rect 6604 1112 6644 1399
rect 6796 1280 6836 1660
rect 6796 1231 6836 1240
rect 6987 1280 7029 1289
rect 6987 1240 6988 1280
rect 7028 1240 7029 1280
rect 7084 1280 7124 4110
rect 7179 4052 7221 4061
rect 7179 4012 7180 4052
rect 7220 4012 7221 4052
rect 7179 4003 7221 4012
rect 7180 2540 7220 4003
rect 7372 3632 7412 4096
rect 7468 4136 7508 5011
rect 7564 4962 7604 4971
rect 7564 4397 7604 4922
rect 7563 4388 7605 4397
rect 7563 4348 7564 4388
rect 7604 4348 7605 4388
rect 7563 4339 7605 4348
rect 7660 4220 7700 8128
rect 7756 8000 7796 8009
rect 7852 8000 7892 8707
rect 7796 7960 7892 8000
rect 7756 7951 7796 7960
rect 7948 7337 7988 11992
rect 8043 9428 8085 9437
rect 8043 9388 8044 9428
rect 8084 9388 8085 9428
rect 8043 9379 8085 9388
rect 7947 7328 7989 7337
rect 7947 7288 7948 7328
rect 7988 7288 7989 7328
rect 7947 7279 7989 7288
rect 7851 7244 7893 7253
rect 7851 7204 7852 7244
rect 7892 7204 7893 7244
rect 7851 7195 7893 7204
rect 7756 7165 7796 7174
rect 7756 6656 7796 7125
rect 7756 6607 7796 6616
rect 7756 5144 7796 5153
rect 7852 5144 7892 7195
rect 7948 7076 7988 7279
rect 8044 7253 8084 9379
rect 8043 7244 8085 7253
rect 8043 7204 8044 7244
rect 8084 7204 8085 7244
rect 8043 7195 8085 7204
rect 7948 7027 7988 7036
rect 8043 6992 8085 7001
rect 8043 6952 8044 6992
rect 8084 6952 8085 6992
rect 8043 6943 8085 6952
rect 7947 5900 7989 5909
rect 7947 5860 7948 5900
rect 7988 5860 7989 5900
rect 7947 5851 7989 5860
rect 7948 5648 7988 5851
rect 7948 5573 7988 5608
rect 7947 5564 7989 5573
rect 7947 5524 7948 5564
rect 7988 5524 7989 5564
rect 7947 5515 7989 5524
rect 7948 5484 7988 5515
rect 8044 5405 8084 6943
rect 8140 6824 8180 14419
rect 8524 14300 8564 17695
rect 8620 16745 8660 22063
rect 8715 21272 8757 21281
rect 8812 21272 8852 24499
rect 8908 23885 8948 25264
rect 9099 25304 9141 25313
rect 9099 25264 9100 25304
rect 9140 25264 9141 25304
rect 9099 25255 9141 25264
rect 9100 25136 9140 25255
rect 9004 25096 9100 25136
rect 9004 24632 9044 25096
rect 9100 25087 9140 25096
rect 9004 24583 9044 24592
rect 9100 24632 9140 24641
rect 9196 24632 9236 26104
rect 9292 25304 9332 26188
rect 9388 26188 9716 26228
rect 9388 26144 9428 26188
rect 9388 26095 9428 26104
rect 9292 25255 9332 25264
rect 9484 26060 9524 26069
rect 9484 25229 9524 26020
rect 9580 25481 9620 25566
rect 9579 25472 9621 25481
rect 9579 25432 9580 25472
rect 9620 25432 9621 25472
rect 9579 25423 9621 25432
rect 9579 25304 9621 25313
rect 9579 25264 9580 25304
rect 9620 25264 9621 25304
rect 9579 25255 9621 25264
rect 9483 25220 9525 25229
rect 9483 25180 9484 25220
rect 9524 25180 9525 25220
rect 9483 25171 9525 25180
rect 9484 25052 9524 25171
rect 9580 25170 9620 25255
rect 9484 25012 9620 25052
rect 9140 24592 9236 24632
rect 9100 24583 9140 24592
rect 9099 24296 9141 24305
rect 9099 24256 9100 24296
rect 9140 24256 9141 24296
rect 9099 24247 9141 24256
rect 8907 23876 8949 23885
rect 8907 23836 8908 23876
rect 8948 23836 8949 23876
rect 8907 23827 8949 23836
rect 8908 23213 8948 23827
rect 8907 23204 8949 23213
rect 8907 23164 8908 23204
rect 8948 23164 8949 23204
rect 8907 23155 8949 23164
rect 8907 23036 8949 23045
rect 8907 22996 8908 23036
rect 8948 22996 8949 23036
rect 8907 22987 8949 22996
rect 8715 21232 8716 21272
rect 8756 21232 8852 21272
rect 8715 21223 8757 21232
rect 8716 19340 8756 21223
rect 8908 20180 8948 22987
rect 9100 22280 9140 24247
rect 9100 22231 9140 22240
rect 9003 21860 9045 21869
rect 9003 21820 9004 21860
rect 9044 21820 9045 21860
rect 9003 21811 9045 21820
rect 9004 21608 9044 21811
rect 9004 21559 9044 21568
rect 9196 21440 9236 24592
rect 9484 24557 9524 24642
rect 9483 24548 9525 24557
rect 9483 24508 9484 24548
rect 9524 24508 9525 24548
rect 9483 24499 9525 24508
rect 9580 24548 9620 25012
rect 9676 24557 9716 26188
rect 9772 25136 9812 27691
rect 9868 26909 9908 29791
rect 9964 29588 10004 29968
rect 10059 29840 10101 29849
rect 10059 29800 10060 29840
rect 10100 29800 10101 29840
rect 10059 29791 10101 29800
rect 10252 29840 10292 29849
rect 10060 29706 10100 29791
rect 10156 29672 10196 29681
rect 9964 29548 10100 29588
rect 10060 28580 10100 29548
rect 10156 28664 10196 29632
rect 10252 29000 10292 29800
rect 10348 29681 10388 30127
rect 10444 29840 10484 30295
rect 10539 29924 10581 29933
rect 10539 29884 10540 29924
rect 10580 29884 10581 29924
rect 10539 29875 10581 29884
rect 10347 29672 10389 29681
rect 10347 29632 10348 29672
rect 10388 29632 10389 29672
rect 10347 29623 10389 29632
rect 10444 29429 10484 29800
rect 10443 29420 10485 29429
rect 10443 29380 10444 29420
rect 10484 29380 10485 29420
rect 10443 29371 10485 29380
rect 10252 28960 10388 29000
rect 10156 28624 10292 28664
rect 10060 28540 10196 28580
rect 9964 28328 10004 28337
rect 9964 28169 10004 28288
rect 10059 28328 10101 28337
rect 10059 28288 10060 28328
rect 10100 28288 10101 28328
rect 10059 28279 10101 28288
rect 10060 28194 10100 28279
rect 9963 28160 10005 28169
rect 9963 28120 9964 28160
rect 10004 28120 10005 28160
rect 9963 28111 10005 28120
rect 10059 28076 10101 28085
rect 10059 28036 10060 28076
rect 10100 28036 10101 28076
rect 10059 28027 10101 28036
rect 9867 26900 9909 26909
rect 9867 26860 9868 26900
rect 9908 26860 9909 26900
rect 9867 26851 9909 26860
rect 10060 26564 10100 28027
rect 10156 26648 10196 28540
rect 10252 28253 10292 28624
rect 10348 28505 10388 28960
rect 10347 28496 10389 28505
rect 10347 28456 10348 28496
rect 10388 28456 10389 28496
rect 10347 28447 10389 28456
rect 10347 28328 10389 28337
rect 10347 28288 10348 28328
rect 10388 28288 10389 28328
rect 10347 28279 10389 28288
rect 10540 28328 10580 29875
rect 10251 28244 10293 28253
rect 10251 28204 10252 28244
rect 10292 28204 10293 28244
rect 10251 28195 10293 28204
rect 10348 27749 10388 28279
rect 10443 28160 10485 28169
rect 10443 28120 10444 28160
rect 10484 28120 10485 28160
rect 10443 28111 10485 28120
rect 10444 27917 10484 28111
rect 10540 28085 10580 28288
rect 10539 28076 10581 28085
rect 10539 28036 10540 28076
rect 10580 28036 10581 28076
rect 10539 28027 10581 28036
rect 10443 27908 10485 27917
rect 10443 27868 10444 27908
rect 10484 27868 10485 27908
rect 10443 27859 10485 27868
rect 10347 27740 10389 27749
rect 10347 27700 10348 27740
rect 10388 27700 10389 27740
rect 10347 27691 10389 27700
rect 10444 27656 10484 27859
rect 10444 27607 10484 27616
rect 10251 26984 10293 26993
rect 10251 26944 10252 26984
rect 10292 26944 10293 26984
rect 10251 26935 10293 26944
rect 10252 26816 10292 26935
rect 10636 26816 10676 32059
rect 10732 28841 10772 35671
rect 10828 35645 10868 35869
rect 11020 35848 11156 35888
rect 11308 35888 11348 36091
rect 10827 35636 10869 35645
rect 10827 35596 10828 35636
rect 10868 35596 10869 35636
rect 10827 35587 10869 35596
rect 10828 35309 10868 35394
rect 10827 35300 10869 35309
rect 10827 35260 10828 35300
rect 10868 35260 10869 35300
rect 10827 35251 10869 35260
rect 11020 35216 11060 35848
rect 11308 35839 11348 35848
rect 11404 35888 11444 36352
rect 11404 35813 11444 35848
rect 11403 35804 11445 35813
rect 11403 35764 11404 35804
rect 11444 35764 11445 35804
rect 11403 35755 11445 35764
rect 11307 35720 11349 35729
rect 11307 35680 11308 35720
rect 11348 35680 11349 35720
rect 11307 35671 11349 35680
rect 11211 35636 11253 35645
rect 11211 35596 11212 35636
rect 11252 35596 11253 35636
rect 11211 35587 11253 35596
rect 10924 35174 10964 35183
rect 11020 35167 11060 35176
rect 11115 35216 11157 35225
rect 11115 35176 11116 35216
rect 11156 35176 11157 35216
rect 11115 35167 11157 35176
rect 10924 34973 10964 35134
rect 10923 34964 10965 34973
rect 10923 34924 10924 34964
rect 10964 34924 10965 34964
rect 10923 34915 10965 34924
rect 11116 34217 11156 35167
rect 11115 34208 11157 34217
rect 11115 34168 11116 34208
rect 11156 34168 11157 34208
rect 11115 34159 11157 34168
rect 11212 33704 11252 35587
rect 11308 35216 11348 35671
rect 11308 34973 11348 35176
rect 11499 35216 11541 35225
rect 11499 35176 11500 35216
rect 11540 35176 11541 35216
rect 11499 35167 11541 35176
rect 11403 35132 11445 35141
rect 11403 35092 11404 35132
rect 11444 35092 11445 35132
rect 11403 35083 11445 35092
rect 11404 34998 11444 35083
rect 11500 35082 11540 35167
rect 11307 34964 11349 34973
rect 11307 34924 11308 34964
rect 11348 34924 11349 34964
rect 11307 34915 11349 34924
rect 11500 34376 11540 34385
rect 11403 33788 11445 33797
rect 11403 33748 11404 33788
rect 11444 33748 11445 33788
rect 11403 33739 11445 33748
rect 11019 33116 11061 33125
rect 11019 33076 11020 33116
rect 11060 33076 11061 33116
rect 11019 33067 11061 33076
rect 10923 31688 10965 31697
rect 10923 31648 10924 31688
rect 10964 31648 10965 31688
rect 10923 31639 10965 31648
rect 10924 31436 10964 31639
rect 10924 31387 10964 31396
rect 11020 31436 11060 33067
rect 10827 31352 10869 31361
rect 10827 31312 10828 31352
rect 10868 31312 10869 31352
rect 10827 31303 10869 31312
rect 10828 30680 10868 31303
rect 10731 28832 10773 28841
rect 10731 28792 10732 28832
rect 10772 28792 10773 28832
rect 10731 28783 10773 28792
rect 10732 28589 10772 28783
rect 10731 28580 10773 28589
rect 10731 28540 10732 28580
rect 10772 28540 10773 28580
rect 10731 28531 10773 28540
rect 10828 27068 10868 30640
rect 10923 30260 10965 30269
rect 10923 30220 10924 30260
rect 10964 30220 10965 30260
rect 10923 30211 10965 30220
rect 10924 29168 10964 30211
rect 10924 27245 10964 29128
rect 11020 29009 11060 31396
rect 11212 31277 11252 33664
rect 11404 33654 11444 33739
rect 11500 33410 11540 34336
rect 11404 33377 11540 33410
rect 11403 33370 11540 33377
rect 11403 33368 11445 33370
rect 11403 33328 11404 33368
rect 11444 33328 11445 33368
rect 11403 33319 11445 33328
rect 11499 33284 11541 33293
rect 11499 33244 11500 33284
rect 11540 33244 11541 33284
rect 11499 33235 11541 33244
rect 11500 31352 11540 33235
rect 11500 31303 11540 31312
rect 11211 31268 11253 31277
rect 11211 31228 11212 31268
rect 11252 31228 11253 31268
rect 11211 31219 11253 31228
rect 11212 30857 11252 31219
rect 11211 30848 11253 30857
rect 11211 30808 11212 30848
rect 11252 30808 11253 30848
rect 11211 30799 11253 30808
rect 11596 30269 11636 37360
rect 11692 36644 11732 36653
rect 11692 35477 11732 36604
rect 11787 36644 11829 36653
rect 11787 36604 11788 36644
rect 11828 36604 11924 36644
rect 11787 36595 11829 36604
rect 11788 36510 11828 36595
rect 11884 36140 11924 36604
rect 11884 36100 11929 36140
rect 11889 35939 11929 36100
rect 11884 35930 11929 35939
rect 11787 35888 11829 35897
rect 11787 35848 11788 35888
rect 11828 35848 11829 35888
rect 11924 35890 11929 35930
rect 11884 35857 11929 35890
rect 11787 35839 11829 35848
rect 11691 35468 11733 35477
rect 11691 35428 11692 35468
rect 11732 35428 11733 35468
rect 11691 35419 11733 35428
rect 11788 34460 11828 35839
rect 11980 35300 12020 39283
rect 12076 39080 12116 39880
rect 12171 39920 12213 39929
rect 12171 39880 12172 39920
rect 12212 39880 12213 39920
rect 12171 39871 12213 39880
rect 12172 39752 12212 39871
rect 12364 39761 12404 40291
rect 12172 39703 12212 39712
rect 12268 39752 12308 39761
rect 12364 39752 12409 39761
rect 12364 39712 12369 39752
rect 12268 39173 12308 39712
rect 12369 39703 12409 39712
rect 12556 39500 12596 40384
rect 12651 40340 12693 40349
rect 12651 40300 12652 40340
rect 12692 40300 12693 40340
rect 12651 40291 12693 40300
rect 12652 39752 12692 40291
rect 12748 39761 12788 39846
rect 12652 39703 12692 39712
rect 12747 39752 12789 39761
rect 12747 39712 12748 39752
rect 12788 39712 12789 39752
rect 12747 39703 12789 39712
rect 12844 39584 12884 40384
rect 12940 40097 12980 42928
rect 13132 42701 13172 42928
rect 13131 42692 13173 42701
rect 13131 42652 13132 42692
rect 13172 42652 13173 42692
rect 13131 42643 13173 42652
rect 13131 42524 13173 42533
rect 13131 42484 13132 42524
rect 13172 42484 13173 42524
rect 13131 42475 13173 42484
rect 12939 40088 12981 40097
rect 12939 40048 12940 40088
rect 12980 40048 12981 40088
rect 12939 40039 12981 40048
rect 12939 39920 12981 39929
rect 12939 39880 12940 39920
rect 12980 39880 12981 39920
rect 12939 39871 12981 39880
rect 12940 39786 12980 39871
rect 13035 39752 13077 39761
rect 13035 39712 13036 39752
rect 13076 39712 13077 39752
rect 13035 39703 13077 39712
rect 12425 39460 12596 39500
rect 12652 39544 12884 39584
rect 12425 39416 12465 39460
rect 12369 39376 12465 39416
rect 12369 39332 12409 39376
rect 12364 39292 12409 39332
rect 12267 39164 12309 39173
rect 12267 39124 12268 39164
rect 12308 39124 12309 39164
rect 12267 39115 12309 39124
rect 12076 39040 12212 39080
rect 12076 38917 12116 38926
rect 12076 38408 12116 38877
rect 12076 38359 12116 38368
rect 12075 36980 12117 36989
rect 12075 36940 12076 36980
rect 12116 36940 12117 36980
rect 12075 36931 12117 36940
rect 12076 36737 12116 36931
rect 12075 36728 12117 36737
rect 12075 36688 12076 36728
rect 12116 36688 12117 36728
rect 12172 36728 12212 39040
rect 12364 39005 12404 39292
rect 12459 39164 12501 39173
rect 12459 39124 12460 39164
rect 12500 39124 12501 39164
rect 12459 39115 12501 39124
rect 12460 39030 12500 39115
rect 12555 39080 12597 39089
rect 12555 39040 12556 39080
rect 12596 39040 12597 39080
rect 12555 39031 12597 39040
rect 12363 38996 12405 39005
rect 12363 38956 12364 38996
rect 12404 38956 12405 38996
rect 12363 38947 12405 38956
rect 12268 38744 12308 38753
rect 12268 37820 12308 38704
rect 12364 38081 12404 38947
rect 12556 38912 12596 39031
rect 12556 38165 12596 38872
rect 12555 38156 12597 38165
rect 12555 38116 12556 38156
rect 12596 38116 12597 38156
rect 12555 38107 12597 38116
rect 12363 38072 12405 38081
rect 12363 38032 12364 38072
rect 12404 38032 12405 38072
rect 12363 38023 12405 38032
rect 12268 37780 12596 37820
rect 12268 36728 12308 36737
rect 12172 36688 12268 36728
rect 12075 36679 12117 36688
rect 12268 35888 12308 36688
rect 12459 36728 12501 36737
rect 12459 36688 12460 36728
rect 12500 36688 12501 36728
rect 12459 36679 12501 36688
rect 12364 35888 12404 35897
rect 12268 35848 12364 35888
rect 12364 35839 12404 35848
rect 12363 35720 12405 35729
rect 12363 35680 12364 35720
rect 12404 35680 12405 35720
rect 12363 35671 12405 35680
rect 12171 35636 12213 35645
rect 12171 35596 12172 35636
rect 12212 35596 12213 35636
rect 12171 35587 12213 35596
rect 11884 35260 12020 35300
rect 11884 35216 11924 35260
rect 11884 35167 11924 35176
rect 12172 35132 12212 35587
rect 12076 35092 12212 35132
rect 11788 34420 12020 34460
rect 11692 34376 11732 34385
rect 11692 33965 11732 34336
rect 11691 33956 11733 33965
rect 11691 33916 11692 33956
rect 11732 33916 11733 33956
rect 11691 33907 11733 33916
rect 11691 33788 11733 33797
rect 11691 33748 11692 33788
rect 11732 33748 11733 33788
rect 11691 33739 11733 33748
rect 11692 33704 11732 33739
rect 11692 33653 11732 33664
rect 11788 33704 11828 33713
rect 11595 30260 11637 30269
rect 11595 30220 11596 30260
rect 11636 30220 11637 30260
rect 11595 30211 11637 30220
rect 11403 30008 11445 30017
rect 11403 29968 11404 30008
rect 11444 29968 11445 30008
rect 11403 29959 11445 29968
rect 11691 30008 11733 30017
rect 11691 29968 11692 30008
rect 11732 29968 11733 30008
rect 11691 29959 11733 29968
rect 11404 29177 11444 29959
rect 11692 29840 11732 29959
rect 11692 29791 11732 29800
rect 11308 29168 11348 29177
rect 11019 29000 11061 29009
rect 11019 28960 11020 29000
rect 11060 28960 11061 29000
rect 11019 28951 11061 28960
rect 11115 28496 11157 28505
rect 11115 28456 11116 28496
rect 11156 28456 11157 28496
rect 11115 28447 11157 28456
rect 11020 28337 11060 28342
rect 11019 28333 11061 28337
rect 11019 28288 11020 28333
rect 11060 28288 11061 28333
rect 11019 28279 11061 28288
rect 11020 28198 11060 28279
rect 11116 28244 11156 28447
rect 11308 28421 11348 29128
rect 11403 29168 11445 29177
rect 11403 29128 11404 29168
rect 11444 29128 11445 29168
rect 11403 29119 11445 29128
rect 11596 29168 11636 29177
rect 11596 29009 11636 29128
rect 11692 29168 11732 29179
rect 11692 29093 11732 29128
rect 11691 29084 11733 29093
rect 11691 29044 11692 29084
rect 11732 29044 11733 29084
rect 11691 29035 11733 29044
rect 11595 29000 11637 29009
rect 11595 28960 11596 29000
rect 11636 28960 11637 29000
rect 11595 28951 11637 28960
rect 11692 28505 11732 29035
rect 11788 28589 11828 33664
rect 11884 32864 11924 32873
rect 11884 32453 11924 32824
rect 11883 32444 11925 32453
rect 11883 32404 11884 32444
rect 11924 32404 11925 32444
rect 11883 32395 11925 32404
rect 11884 31268 11924 32395
rect 11980 31697 12020 34420
rect 12076 31865 12116 35092
rect 12364 33797 12404 35671
rect 12363 33788 12405 33797
rect 12363 33748 12364 33788
rect 12404 33748 12405 33788
rect 12363 33739 12405 33748
rect 12172 33620 12212 33629
rect 12075 31856 12117 31865
rect 12075 31816 12076 31856
rect 12116 31816 12117 31856
rect 12075 31807 12117 31816
rect 11979 31688 12021 31697
rect 11979 31648 11980 31688
rect 12020 31648 12021 31688
rect 11979 31639 12021 31648
rect 12172 31529 12212 33580
rect 12267 33620 12309 33629
rect 12267 33580 12268 33620
rect 12308 33580 12309 33620
rect 12267 33571 12309 33580
rect 12268 32789 12308 33571
rect 12267 32780 12309 32789
rect 12267 32740 12268 32780
rect 12308 32740 12309 32780
rect 12267 32731 12309 32740
rect 12171 31520 12213 31529
rect 12171 31480 12172 31520
rect 12212 31480 12213 31520
rect 12171 31471 12213 31480
rect 12028 31361 12068 31370
rect 12068 31321 12308 31352
rect 12028 31312 12308 31321
rect 11884 31228 12020 31268
rect 11883 30092 11925 30101
rect 11883 30052 11884 30092
rect 11924 30052 11925 30092
rect 11883 30043 11925 30052
rect 11884 29849 11924 30043
rect 11883 29840 11925 29849
rect 11883 29800 11884 29840
rect 11924 29800 11925 29840
rect 11883 29791 11925 29800
rect 11980 29093 12020 31228
rect 12171 31184 12213 31193
rect 12171 31144 12172 31184
rect 12212 31144 12213 31184
rect 12171 31135 12213 31144
rect 12172 31050 12212 31135
rect 12268 30848 12308 31312
rect 12460 30848 12500 36679
rect 12556 35729 12596 37780
rect 12555 35720 12597 35729
rect 12555 35680 12556 35720
rect 12596 35680 12597 35720
rect 12555 35671 12597 35680
rect 12555 35468 12597 35477
rect 12555 35428 12556 35468
rect 12596 35428 12597 35468
rect 12555 35419 12597 35428
rect 12556 33881 12596 35419
rect 12555 33872 12597 33881
rect 12555 33832 12556 33872
rect 12596 33832 12597 33872
rect 12555 33823 12597 33832
rect 12652 33377 12692 39544
rect 12939 39500 12981 39509
rect 12939 39460 12940 39500
rect 12980 39460 12981 39500
rect 12939 39451 12981 39460
rect 12940 39341 12980 39451
rect 12939 39332 12981 39341
rect 12939 39292 12940 39332
rect 12980 39292 12981 39332
rect 12939 39283 12981 39292
rect 13036 39257 13076 39703
rect 13035 39248 13077 39257
rect 13035 39208 13036 39248
rect 13076 39208 13077 39248
rect 13035 39199 13077 39208
rect 13132 39173 13172 42475
rect 13324 41609 13364 42928
rect 13516 41693 13556 42928
rect 13515 41684 13557 41693
rect 13515 41644 13516 41684
rect 13556 41644 13557 41684
rect 13515 41635 13557 41644
rect 13708 41609 13748 42928
rect 13900 41777 13940 42928
rect 13899 41768 13941 41777
rect 13899 41728 13900 41768
rect 13940 41728 13941 41768
rect 13899 41719 13941 41728
rect 14092 41609 14132 42928
rect 14284 41693 14324 42928
rect 14283 41684 14325 41693
rect 14283 41644 14284 41684
rect 14324 41644 14325 41684
rect 14283 41635 14325 41644
rect 14476 41609 14516 42928
rect 14668 41609 14708 42928
rect 13323 41600 13365 41609
rect 13323 41560 13324 41600
rect 13364 41560 13365 41600
rect 13323 41551 13365 41560
rect 13707 41600 13749 41609
rect 13707 41560 13708 41600
rect 13748 41560 13749 41600
rect 13707 41551 13749 41560
rect 14091 41600 14133 41609
rect 14091 41560 14092 41600
rect 14132 41560 14133 41600
rect 14091 41551 14133 41560
rect 14475 41600 14517 41609
rect 14475 41560 14476 41600
rect 14516 41560 14517 41600
rect 14475 41551 14517 41560
rect 14667 41600 14709 41609
rect 14667 41560 14668 41600
rect 14708 41560 14709 41600
rect 14667 41551 14709 41560
rect 13803 41432 13845 41441
rect 13803 41392 13804 41432
rect 13844 41392 13845 41432
rect 13803 41383 13845 41392
rect 13804 41298 13844 41383
rect 13228 41264 13268 41273
rect 13228 40685 13268 41224
rect 13611 41180 13653 41189
rect 13611 41140 13612 41180
rect 13652 41140 13653 41180
rect 13611 41131 13653 41140
rect 13996 41180 14036 41189
rect 14572 41180 14612 41189
rect 14860 41180 14900 42928
rect 14036 41140 14132 41180
rect 13996 41131 14036 41140
rect 13420 41012 13460 41021
rect 13324 40972 13420 41012
rect 13227 40676 13269 40685
rect 13227 40636 13228 40676
rect 13268 40636 13269 40676
rect 13227 40627 13269 40636
rect 13324 39752 13364 40972
rect 13420 40963 13460 40972
rect 13612 40937 13652 41131
rect 13611 40928 13653 40937
rect 13611 40888 13612 40928
rect 13652 40888 13653 40928
rect 13611 40879 13653 40888
rect 13419 40424 13461 40433
rect 13419 40384 13420 40424
rect 13460 40384 13461 40424
rect 13419 40375 13461 40384
rect 13324 39703 13364 39712
rect 13420 39752 13460 40375
rect 13515 40172 13557 40181
rect 13515 40132 13516 40172
rect 13556 40132 13557 40172
rect 13515 40123 13557 40132
rect 13420 39257 13460 39712
rect 13419 39248 13461 39257
rect 13419 39208 13420 39248
rect 13460 39208 13461 39248
rect 13419 39199 13461 39208
rect 12843 39164 12885 39173
rect 12843 39124 12844 39164
rect 12884 39124 12885 39164
rect 12843 39115 12885 39124
rect 13131 39164 13173 39173
rect 13131 39124 13132 39164
rect 13172 39124 13173 39164
rect 13131 39115 13173 39124
rect 12844 39080 12884 39115
rect 12844 39029 12884 39040
rect 13036 38996 13076 39005
rect 12844 38240 12884 38249
rect 12747 37820 12789 37829
rect 12747 37780 12748 37820
rect 12788 37780 12789 37820
rect 12844 37820 12884 38200
rect 13036 38165 13076 38956
rect 13035 38156 13077 38165
rect 13035 38116 13036 38156
rect 13076 38116 13077 38156
rect 13035 38107 13077 38116
rect 13419 37820 13461 37829
rect 12844 37780 13076 37820
rect 12747 37771 12789 37780
rect 12748 37400 12788 37771
rect 12748 37351 12788 37360
rect 12940 37232 12980 37241
rect 12844 37192 12940 37232
rect 12844 36728 12884 37192
rect 12940 37183 12980 37192
rect 12796 36718 12884 36728
rect 12836 36688 12884 36718
rect 12940 36812 12980 36821
rect 12796 36669 12836 36678
rect 12940 36056 12980 36772
rect 13036 36401 13076 37780
rect 13419 37780 13420 37820
rect 13460 37780 13461 37820
rect 13419 37771 13461 37780
rect 13035 36392 13077 36401
rect 13035 36352 13036 36392
rect 13076 36352 13077 36392
rect 13035 36343 13077 36352
rect 12748 36016 12980 36056
rect 12748 34889 12788 36016
rect 12892 35897 12932 35906
rect 12932 35857 13364 35888
rect 12892 35848 13364 35857
rect 13035 35720 13077 35729
rect 13035 35680 13036 35720
rect 13076 35680 13077 35720
rect 13035 35671 13077 35680
rect 13036 35586 13076 35671
rect 12843 35552 12885 35561
rect 12843 35512 12844 35552
rect 12884 35512 12885 35552
rect 12843 35503 12885 35512
rect 12747 34880 12789 34889
rect 12747 34840 12748 34880
rect 12788 34840 12789 34880
rect 12747 34831 12789 34840
rect 12747 33788 12789 33797
rect 12747 33748 12748 33788
rect 12788 33748 12789 33788
rect 12747 33739 12789 33748
rect 12748 33704 12788 33739
rect 12844 33713 12884 35503
rect 13324 35384 13364 35848
rect 13324 35335 13364 35344
rect 13035 35216 13077 35225
rect 13035 35176 13036 35216
rect 13076 35176 13077 35216
rect 13035 35167 13077 35176
rect 13132 35216 13172 35227
rect 12939 34544 12981 34553
rect 12939 34504 12940 34544
rect 12980 34504 12981 34544
rect 12939 34495 12981 34504
rect 12940 34376 12980 34495
rect 12940 34327 12980 34336
rect 13036 34208 13076 35167
rect 13132 35141 13172 35176
rect 13131 35132 13173 35141
rect 13131 35092 13132 35132
rect 13172 35092 13268 35132
rect 13131 35083 13173 35092
rect 13132 34301 13172 34386
rect 13131 34292 13173 34301
rect 13131 34252 13132 34292
rect 13172 34252 13173 34292
rect 13131 34243 13173 34252
rect 12940 34168 13076 34208
rect 12748 33653 12788 33664
rect 12843 33704 12885 33713
rect 12843 33664 12844 33704
rect 12884 33664 12885 33704
rect 12843 33655 12885 33664
rect 12844 33536 12884 33655
rect 12748 33496 12884 33536
rect 12651 33368 12693 33377
rect 12651 33328 12652 33368
rect 12692 33328 12693 33368
rect 12651 33319 12693 33328
rect 12748 32192 12788 33496
rect 12843 33368 12885 33377
rect 12843 33328 12844 33368
rect 12884 33328 12885 33368
rect 12843 33319 12885 33328
rect 12268 30799 12308 30808
rect 12364 30808 12500 30848
rect 12652 32152 12788 32192
rect 12075 30764 12117 30773
rect 12075 30724 12076 30764
rect 12116 30724 12117 30764
rect 12075 30715 12117 30724
rect 12076 30680 12116 30715
rect 12076 30629 12116 30640
rect 12364 30353 12404 30808
rect 12460 30680 12500 30689
rect 12363 30344 12405 30353
rect 12363 30304 12364 30344
rect 12404 30304 12405 30344
rect 12363 30295 12405 30304
rect 12075 29840 12117 29849
rect 12075 29800 12076 29840
rect 12116 29800 12117 29840
rect 12075 29791 12117 29800
rect 12076 29513 12116 29791
rect 12075 29504 12117 29513
rect 12075 29464 12076 29504
rect 12116 29464 12117 29504
rect 12075 29455 12117 29464
rect 12364 29147 12404 30295
rect 12460 30101 12500 30640
rect 12555 30428 12597 30437
rect 12555 30388 12556 30428
rect 12596 30388 12597 30428
rect 12555 30379 12597 30388
rect 12556 30294 12596 30379
rect 12459 30092 12501 30101
rect 12459 30052 12460 30092
rect 12500 30052 12501 30092
rect 12459 30043 12501 30052
rect 12268 29126 12404 29147
rect 11979 29084 12021 29093
rect 11979 29044 11980 29084
rect 12020 29044 12021 29084
rect 12308 29107 12404 29126
rect 12268 29077 12308 29086
rect 11979 29035 12021 29044
rect 12652 29000 12692 32152
rect 12747 31352 12789 31361
rect 12747 31312 12748 31352
rect 12788 31312 12789 31352
rect 12747 31303 12789 31312
rect 12748 31218 12788 31303
rect 12652 28960 12788 29000
rect 11979 28916 12021 28925
rect 11979 28876 11980 28916
rect 12020 28876 12021 28916
rect 11979 28867 12021 28876
rect 11980 28782 12020 28867
rect 11787 28580 11829 28589
rect 11787 28540 11788 28580
rect 11828 28540 11829 28580
rect 11787 28531 11829 28540
rect 11403 28496 11445 28505
rect 11403 28456 11404 28496
rect 11444 28456 11445 28496
rect 11403 28447 11445 28456
rect 11691 28496 11733 28505
rect 11691 28456 11692 28496
rect 11732 28456 11733 28496
rect 11691 28447 11733 28456
rect 12172 28496 12212 28505
rect 12212 28456 12596 28496
rect 12172 28447 12212 28456
rect 11307 28412 11349 28421
rect 11307 28372 11308 28412
rect 11348 28372 11349 28412
rect 11307 28363 11349 28372
rect 11404 28328 11444 28447
rect 11787 28412 11829 28421
rect 11787 28372 11788 28412
rect 11828 28372 11829 28412
rect 11787 28363 11829 28372
rect 11404 28279 11444 28288
rect 11788 28328 11828 28363
rect 11212 28244 11252 28253
rect 11116 28204 11212 28244
rect 11212 28195 11252 28204
rect 11499 28160 11541 28169
rect 11499 28120 11500 28160
rect 11540 28120 11541 28160
rect 11499 28111 11541 28120
rect 11691 28160 11733 28169
rect 11691 28116 11692 28160
rect 11732 28116 11733 28160
rect 11691 28111 11733 28116
rect 11211 28076 11253 28085
rect 11211 28036 11212 28076
rect 11252 28036 11253 28076
rect 11211 28027 11253 28036
rect 10923 27236 10965 27245
rect 10923 27196 10924 27236
rect 10964 27196 10965 27236
rect 10923 27187 10965 27196
rect 10828 27028 11060 27068
rect 10732 26825 10772 26910
rect 10828 26909 10868 26940
rect 10827 26900 10869 26909
rect 10827 26860 10828 26900
rect 10868 26860 10869 26900
rect 10827 26851 10869 26860
rect 10252 26767 10292 26776
rect 10348 26776 10676 26816
rect 10731 26816 10773 26825
rect 10731 26776 10732 26816
rect 10772 26776 10773 26816
rect 10156 26608 10292 26648
rect 10060 26524 10196 26564
rect 9963 26396 10005 26405
rect 9963 26356 9964 26396
rect 10004 26356 10005 26396
rect 9963 26347 10005 26356
rect 9964 26144 10004 26347
rect 9964 26095 10004 26104
rect 9867 25472 9909 25481
rect 9867 25432 9868 25472
rect 9908 25432 9909 25472
rect 9867 25423 9909 25432
rect 9868 25304 9908 25423
rect 10060 25313 10100 25398
rect 9868 25255 9908 25264
rect 10059 25304 10101 25313
rect 10059 25264 10060 25304
rect 10100 25264 10101 25304
rect 10059 25255 10101 25264
rect 10156 25304 10196 26524
rect 10156 25229 10196 25264
rect 10155 25220 10197 25229
rect 10155 25180 10156 25220
rect 10196 25180 10197 25220
rect 10155 25171 10197 25180
rect 9964 25136 10004 25145
rect 9772 25096 9908 25136
rect 9580 24053 9620 24508
rect 9675 24548 9717 24557
rect 9675 24508 9676 24548
rect 9716 24508 9717 24548
rect 9675 24499 9717 24508
rect 9579 24044 9621 24053
rect 9579 24004 9580 24044
rect 9620 24004 9621 24044
rect 9579 23995 9621 24004
rect 9388 23792 9428 23801
rect 9292 23752 9388 23792
rect 9292 23045 9332 23752
rect 9388 23743 9428 23752
rect 9387 23204 9429 23213
rect 9387 23164 9388 23204
rect 9428 23164 9429 23204
rect 9387 23155 9429 23164
rect 9579 23204 9621 23213
rect 9579 23164 9580 23204
rect 9620 23164 9621 23204
rect 9579 23155 9621 23164
rect 9388 23120 9428 23155
rect 9388 23069 9428 23080
rect 9291 23036 9333 23045
rect 9291 22996 9292 23036
rect 9332 22996 9333 23036
rect 9291 22987 9333 22996
rect 9580 22868 9620 23155
rect 9772 22868 9812 22877
rect 9291 22532 9333 22541
rect 9291 22492 9292 22532
rect 9332 22492 9333 22532
rect 9291 22483 9333 22492
rect 9292 22289 9332 22483
rect 9291 22280 9333 22289
rect 9580 22285 9620 22828
rect 9291 22240 9292 22280
rect 9332 22240 9333 22280
rect 9291 22231 9333 22240
rect 9388 22245 9580 22280
rect 9388 22240 9620 22245
rect 9292 21608 9332 22231
rect 9292 21559 9332 21568
rect 9004 21400 9236 21440
rect 9004 20516 9044 21400
rect 9388 20768 9428 22240
rect 9580 22236 9620 22240
rect 9676 22828 9772 22868
rect 9483 21524 9525 21533
rect 9483 21484 9484 21524
rect 9524 21484 9525 21524
rect 9483 21475 9525 21484
rect 9388 20719 9428 20728
rect 9484 20768 9524 21475
rect 9484 20719 9524 20728
rect 9580 20768 9620 20777
rect 9676 20768 9716 22828
rect 9772 22819 9812 22828
rect 9771 22448 9813 22457
rect 9771 22408 9772 22448
rect 9812 22408 9813 22448
rect 9771 22399 9813 22408
rect 9772 22070 9812 22399
rect 9772 22021 9812 22030
rect 9868 21944 9908 25096
rect 9964 24977 10004 25096
rect 9963 24968 10005 24977
rect 9963 24928 9964 24968
rect 10004 24928 10005 24968
rect 9963 24919 10005 24928
rect 10059 24716 10101 24725
rect 10059 24676 10060 24716
rect 10100 24676 10101 24716
rect 10059 24667 10101 24676
rect 10060 24632 10100 24667
rect 10060 24581 10100 24592
rect 10059 24128 10101 24137
rect 10059 24088 10060 24128
rect 10100 24088 10101 24128
rect 10059 24079 10101 24088
rect 9964 23213 10004 23227
rect 9963 23204 10005 23213
rect 9963 23164 9964 23204
rect 10004 23164 10005 23204
rect 9963 23155 10005 23164
rect 9964 23132 10004 23155
rect 9964 23083 10004 23092
rect 10060 23120 10100 24079
rect 10060 23071 10100 23080
rect 10155 23120 10197 23129
rect 10155 23080 10156 23120
rect 10196 23080 10197 23120
rect 10155 23071 10197 23080
rect 10156 22986 10196 23071
rect 9964 22285 10004 22289
rect 10155 22285 10197 22289
rect 9964 22280 10197 22285
rect 10004 22245 10156 22280
rect 10004 22240 10007 22245
rect 10155 22240 10156 22245
rect 10196 22240 10197 22280
rect 9964 22231 10004 22240
rect 10155 22231 10197 22240
rect 9620 20728 9716 20768
rect 9772 21904 9908 21944
rect 9580 20719 9620 20728
rect 9675 20600 9717 20609
rect 9675 20560 9676 20600
rect 9716 20560 9717 20600
rect 9675 20551 9717 20560
rect 9004 20476 9140 20516
rect 8908 20140 9044 20180
rect 8812 19349 8852 19380
rect 8716 19291 8756 19300
rect 8811 19340 8853 19349
rect 8811 19300 8812 19340
rect 8852 19300 8853 19340
rect 8811 19291 8853 19300
rect 8812 19256 8852 19291
rect 8812 18677 8852 19216
rect 8811 18668 8853 18677
rect 8811 18628 8812 18668
rect 8852 18628 8853 18668
rect 8811 18619 8853 18628
rect 8716 17749 8756 17758
rect 8619 16736 8661 16745
rect 8619 16696 8620 16736
rect 8660 16696 8661 16736
rect 8619 16687 8661 16696
rect 8619 16484 8661 16493
rect 8619 16444 8620 16484
rect 8660 16444 8661 16484
rect 8716 16484 8756 17709
rect 8907 17660 8949 17669
rect 8907 17620 8908 17660
rect 8948 17620 8949 17660
rect 8907 17611 8949 17620
rect 8908 17526 8948 17611
rect 8812 16484 8852 16493
rect 8716 16444 8812 16484
rect 8619 16435 8661 16444
rect 8812 16435 8852 16444
rect 8620 16232 8660 16435
rect 9004 16325 9044 20140
rect 9100 19349 9140 20476
rect 9676 20466 9716 20551
rect 9772 20180 9812 21904
rect 10155 21440 10197 21449
rect 10155 21400 10156 21440
rect 10196 21400 10197 21440
rect 10155 21391 10197 21400
rect 9867 21356 9909 21365
rect 9867 21316 9868 21356
rect 9908 21316 9909 21356
rect 9867 21307 9909 21316
rect 9388 20140 9812 20180
rect 9292 20096 9332 20105
rect 9196 20056 9292 20096
rect 9196 19433 9236 20056
rect 9292 20047 9332 20056
rect 9291 19676 9333 19685
rect 9291 19636 9292 19676
rect 9332 19636 9333 19676
rect 9291 19627 9333 19636
rect 9195 19424 9237 19433
rect 9195 19384 9196 19424
rect 9236 19384 9237 19424
rect 9195 19375 9237 19384
rect 9099 19340 9141 19349
rect 9099 19300 9100 19340
rect 9140 19300 9141 19340
rect 9099 19291 9141 19300
rect 9196 19172 9236 19375
rect 9292 19256 9332 19627
rect 9292 19207 9332 19216
rect 9100 19132 9236 19172
rect 9003 16316 9045 16325
rect 9003 16276 9004 16316
rect 9044 16276 9045 16316
rect 9003 16267 9045 16276
rect 8620 16183 8660 16192
rect 9100 16148 9140 19132
rect 9291 19088 9333 19097
rect 9291 19048 9292 19088
rect 9332 19048 9333 19088
rect 9291 19039 9333 19048
rect 9195 17072 9237 17081
rect 9195 17032 9196 17072
rect 9236 17032 9237 17072
rect 9195 17023 9237 17032
rect 9196 16493 9236 17023
rect 9195 16484 9237 16493
rect 9195 16444 9196 16484
rect 9236 16444 9237 16484
rect 9195 16435 9237 16444
rect 9004 16108 9140 16148
rect 8907 15812 8949 15821
rect 8907 15772 8908 15812
rect 8948 15772 8949 15812
rect 8907 15763 8949 15772
rect 8908 15728 8948 15763
rect 8908 15677 8948 15688
rect 8811 15560 8853 15569
rect 8716 15546 8756 15555
rect 8811 15520 8812 15560
rect 8852 15520 8853 15560
rect 8811 15511 8853 15520
rect 8716 14981 8756 15506
rect 8715 14972 8757 14981
rect 8715 14932 8716 14972
rect 8756 14932 8757 14972
rect 8715 14923 8757 14932
rect 8524 14260 8660 14300
rect 8524 14132 8564 14141
rect 8380 14006 8420 14015
rect 8235 13964 8277 13973
rect 8235 13924 8236 13964
rect 8276 13924 8277 13964
rect 8380 13964 8420 13966
rect 8380 13924 8468 13964
rect 8235 13915 8277 13924
rect 8236 13208 8276 13915
rect 8428 13460 8468 13924
rect 8428 13411 8468 13420
rect 8236 12545 8276 13168
rect 8235 12536 8277 12545
rect 8235 12496 8236 12536
rect 8276 12496 8277 12536
rect 8235 12487 8277 12496
rect 8524 12461 8564 14092
rect 8523 12452 8565 12461
rect 8523 12412 8524 12452
rect 8564 12412 8565 12452
rect 8523 12403 8565 12412
rect 8523 11780 8565 11789
rect 8523 11740 8524 11780
rect 8564 11740 8565 11780
rect 8523 11731 8565 11740
rect 8332 11701 8372 11710
rect 8235 11528 8277 11537
rect 8235 11488 8236 11528
rect 8276 11488 8277 11528
rect 8235 11479 8277 11488
rect 8236 9521 8276 11479
rect 8332 11201 8372 11661
rect 8427 11612 8469 11621
rect 8427 11572 8428 11612
rect 8468 11572 8469 11612
rect 8427 11563 8469 11572
rect 8524 11612 8564 11731
rect 8524 11563 8564 11572
rect 8331 11192 8373 11201
rect 8331 11152 8332 11192
rect 8372 11152 8373 11192
rect 8331 11143 8373 11152
rect 8428 10781 8468 11563
rect 8620 11360 8660 14260
rect 8715 13544 8757 13553
rect 8715 13504 8716 13544
rect 8756 13504 8757 13544
rect 8715 13495 8757 13504
rect 8716 13301 8756 13495
rect 8715 13292 8757 13301
rect 8715 13252 8716 13292
rect 8756 13252 8757 13292
rect 8715 13243 8757 13252
rect 8716 13208 8756 13243
rect 8716 13157 8756 13168
rect 8715 12536 8757 12545
rect 8715 12496 8716 12536
rect 8756 12496 8757 12536
rect 8715 12487 8757 12496
rect 8716 12402 8756 12487
rect 8715 12200 8757 12209
rect 8715 12160 8716 12200
rect 8756 12160 8757 12200
rect 8715 12151 8757 12160
rect 8524 11320 8660 11360
rect 8716 11696 8756 12151
rect 8427 10772 8469 10781
rect 8427 10732 8428 10772
rect 8468 10732 8469 10772
rect 8427 10723 8469 10732
rect 8331 10268 8373 10277
rect 8331 10228 8332 10268
rect 8372 10228 8373 10268
rect 8331 10219 8373 10228
rect 8235 9512 8277 9521
rect 8235 9472 8236 9512
rect 8276 9472 8277 9512
rect 8235 9463 8277 9472
rect 8332 9512 8372 10219
rect 8428 10184 8468 10723
rect 8428 10025 8468 10144
rect 8427 10016 8469 10025
rect 8427 9976 8428 10016
rect 8468 9976 8469 10016
rect 8427 9967 8469 9976
rect 8332 9463 8372 9472
rect 8427 9512 8469 9521
rect 8427 9472 8428 9512
rect 8468 9472 8469 9512
rect 8427 9463 8469 9472
rect 8428 9378 8468 9463
rect 8427 7244 8469 7253
rect 8427 7204 8428 7244
rect 8468 7204 8469 7244
rect 8427 7195 8469 7204
rect 8428 7174 8468 7195
rect 8428 7109 8468 7134
rect 8236 7001 8276 7086
rect 8524 7076 8564 11320
rect 8619 10352 8661 10361
rect 8619 10312 8620 10352
rect 8660 10312 8661 10352
rect 8619 10303 8661 10312
rect 8620 10218 8660 10303
rect 8716 9773 8756 11656
rect 8812 11192 8852 15511
rect 8908 12629 8948 12714
rect 8907 12620 8949 12629
rect 8907 12580 8908 12620
rect 8948 12580 8949 12620
rect 8907 12571 8949 12580
rect 8907 12452 8949 12461
rect 8907 12412 8908 12452
rect 8948 12412 8949 12452
rect 8907 12403 8949 12412
rect 8908 11369 8948 12403
rect 9004 11537 9044 16108
rect 9099 14636 9141 14645
rect 9099 14596 9100 14636
rect 9140 14596 9141 14636
rect 9099 14587 9141 14596
rect 9003 11528 9045 11537
rect 9003 11488 9004 11528
rect 9044 11488 9045 11528
rect 9003 11479 9045 11488
rect 8907 11360 8949 11369
rect 8907 11320 8908 11360
rect 8948 11320 8949 11360
rect 8907 11311 8949 11320
rect 9003 11192 9045 11201
rect 8812 11152 8948 11192
rect 8812 11024 8852 11033
rect 8812 10781 8852 10984
rect 8811 10772 8853 10781
rect 8811 10732 8812 10772
rect 8852 10732 8853 10772
rect 8811 10723 8853 10732
rect 8811 10604 8853 10613
rect 8811 10564 8812 10604
rect 8852 10564 8853 10604
rect 8811 10555 8853 10564
rect 8812 10445 8852 10555
rect 8908 10529 8948 11152
rect 9003 11152 9004 11192
rect 9044 11152 9045 11192
rect 9003 11143 9045 11152
rect 9004 11058 9044 11143
rect 9003 10604 9045 10613
rect 9003 10564 9004 10604
rect 9044 10564 9045 10604
rect 9003 10555 9045 10564
rect 8907 10520 8949 10529
rect 8907 10480 8908 10520
rect 8948 10480 8949 10520
rect 8907 10471 8949 10480
rect 8811 10436 8853 10445
rect 8811 10396 8812 10436
rect 8852 10396 8853 10436
rect 8811 10387 8853 10396
rect 8715 9764 8757 9773
rect 8715 9724 8716 9764
rect 8756 9724 8757 9764
rect 8715 9715 8757 9724
rect 8812 9680 8852 10387
rect 8907 10352 8949 10361
rect 8907 10312 8908 10352
rect 8948 10312 8949 10352
rect 8907 10303 8949 10312
rect 8908 10184 8948 10303
rect 8908 10135 8948 10144
rect 9004 10184 9044 10555
rect 9100 10361 9140 14587
rect 9196 14552 9236 16435
rect 9292 16073 9332 19039
rect 9291 16064 9333 16073
rect 9291 16024 9292 16064
rect 9332 16024 9333 16064
rect 9291 16015 9333 16024
rect 9388 15821 9428 20140
rect 9868 20096 9908 21307
rect 9676 20056 9908 20096
rect 9483 19676 9525 19685
rect 9483 19636 9484 19676
rect 9524 19636 9525 19676
rect 9483 19627 9525 19636
rect 9484 16400 9524 19627
rect 9579 19508 9621 19517
rect 9579 19468 9580 19508
rect 9620 19468 9621 19508
rect 9579 19459 9621 19468
rect 9580 18089 9620 19459
rect 9676 18593 9716 20056
rect 9820 19265 9860 19274
rect 9860 19225 9908 19256
rect 9820 19216 9908 19225
rect 9771 18920 9813 18929
rect 9771 18880 9772 18920
rect 9812 18880 9813 18920
rect 9771 18871 9813 18880
rect 9675 18584 9717 18593
rect 9675 18544 9676 18584
rect 9716 18544 9717 18584
rect 9675 18535 9717 18544
rect 9676 18450 9716 18535
rect 9579 18080 9621 18089
rect 9579 18040 9580 18080
rect 9620 18040 9621 18080
rect 9579 18031 9621 18040
rect 9676 17744 9716 17753
rect 9676 17240 9716 17704
rect 9772 17744 9812 18871
rect 9868 18752 9908 19216
rect 10156 19172 10196 21391
rect 10252 20189 10292 26608
rect 10348 23801 10388 26776
rect 10731 26767 10773 26776
rect 10828 26816 10868 26851
rect 10443 26648 10485 26657
rect 10443 26608 10444 26648
rect 10484 26608 10485 26648
rect 10443 26599 10485 26608
rect 10444 26139 10484 26599
rect 10828 26564 10868 26776
rect 10924 26816 10964 26825
rect 10924 26657 10964 26776
rect 10923 26648 10965 26657
rect 10923 26608 10924 26648
rect 10964 26608 10965 26648
rect 10923 26599 10965 26608
rect 10444 26090 10484 26099
rect 10540 26524 10868 26564
rect 10443 25304 10485 25313
rect 10443 25264 10444 25304
rect 10484 25264 10485 25304
rect 10443 25255 10485 25264
rect 10540 25304 10580 26524
rect 10827 26396 10869 26405
rect 10827 26356 10828 26396
rect 10868 26356 10869 26396
rect 10827 26347 10869 26356
rect 10828 26237 10868 26347
rect 10636 26228 10676 26237
rect 10636 25481 10676 26188
rect 10827 26228 10869 26237
rect 10827 26188 10828 26228
rect 10868 26188 10869 26228
rect 10827 26179 10869 26188
rect 10828 26144 10868 26179
rect 10828 26094 10868 26104
rect 10635 25472 10677 25481
rect 10635 25432 10636 25472
rect 10676 25432 10677 25472
rect 10635 25423 10677 25432
rect 10444 25170 10484 25255
rect 10540 25052 10580 25264
rect 10444 25012 10580 25052
rect 10636 25304 10676 25313
rect 10347 23792 10389 23801
rect 10347 23752 10348 23792
rect 10388 23752 10389 23792
rect 10347 23743 10389 23752
rect 10348 23129 10388 23743
rect 10347 23120 10389 23129
rect 10347 23080 10348 23120
rect 10388 23080 10389 23120
rect 10347 23071 10389 23080
rect 10347 22700 10389 22709
rect 10347 22660 10348 22700
rect 10388 22660 10389 22700
rect 10347 22651 10389 22660
rect 10251 20180 10293 20189
rect 10251 20140 10252 20180
rect 10292 20140 10293 20180
rect 10251 20131 10293 20140
rect 10348 19181 10388 22651
rect 10347 19172 10389 19181
rect 10156 19132 10303 19172
rect 9963 19088 10005 19097
rect 9963 19048 9964 19088
rect 10004 19048 10005 19088
rect 9963 19039 10005 19048
rect 9964 18954 10004 19039
rect 10263 18920 10303 19132
rect 10347 19132 10348 19172
rect 10388 19132 10389 19172
rect 10347 19123 10389 19132
rect 10252 18880 10303 18920
rect 9868 18703 9908 18712
rect 9963 18752 10005 18761
rect 9963 18712 9964 18752
rect 10004 18712 10005 18752
rect 9963 18703 10005 18712
rect 9812 17704 9908 17744
rect 9772 17695 9812 17704
rect 9772 17240 9812 17249
rect 9676 17200 9772 17240
rect 9772 17191 9812 17200
rect 9579 17072 9621 17081
rect 9579 17032 9580 17072
rect 9620 17032 9621 17072
rect 9579 17023 9621 17032
rect 9580 16938 9620 17023
rect 9771 16568 9813 16577
rect 9868 16568 9908 17704
rect 9964 16661 10004 18703
rect 10060 18584 10100 18593
rect 10060 18341 10100 18544
rect 10059 18332 10101 18341
rect 10059 18292 10060 18332
rect 10100 18292 10101 18332
rect 10059 18283 10101 18292
rect 10252 17828 10292 18880
rect 10252 17779 10292 17788
rect 10155 17744 10197 17753
rect 10155 17704 10156 17744
rect 10196 17704 10197 17744
rect 10155 17695 10197 17704
rect 10156 17610 10196 17695
rect 10444 17240 10484 25012
rect 10540 24622 10580 24631
rect 10636 24622 10676 25264
rect 11020 25229 11060 27028
rect 11115 26816 11157 26825
rect 11115 26776 11116 26816
rect 11156 26776 11157 26816
rect 11115 26767 11157 26776
rect 11116 26648 11156 26767
rect 11116 26599 11156 26608
rect 11019 25220 11061 25229
rect 11019 25180 11020 25220
rect 11060 25180 11061 25220
rect 11019 25171 11061 25180
rect 10827 25136 10869 25145
rect 10827 25096 10828 25136
rect 10868 25096 10869 25136
rect 10827 25087 10869 25096
rect 11115 25136 11157 25145
rect 11115 25096 11116 25136
rect 11156 25096 11157 25136
rect 11115 25087 11157 25096
rect 10828 25002 10868 25087
rect 10923 24968 10965 24977
rect 10923 24928 10924 24968
rect 10964 24928 10965 24968
rect 10923 24919 10965 24928
rect 10731 24716 10773 24725
rect 10731 24676 10732 24716
rect 10772 24676 10773 24716
rect 10924 24716 10964 24919
rect 10924 24676 11060 24716
rect 10731 24667 10773 24676
rect 10580 24582 10676 24622
rect 10732 24582 10772 24667
rect 11020 24653 11060 24676
rect 11020 24604 11060 24613
rect 11116 24632 11156 25087
rect 11212 24800 11252 28027
rect 11500 28026 11540 28111
rect 11692 28025 11732 28111
rect 11788 27824 11828 28288
rect 11884 28328 11924 28337
rect 12363 28328 12405 28337
rect 11924 28288 12212 28328
rect 11884 28279 11924 28288
rect 11884 27868 12116 27908
rect 11884 27824 11924 27868
rect 11788 27784 11884 27824
rect 11884 27775 11924 27784
rect 11979 27740 12021 27749
rect 11979 27700 11980 27740
rect 12020 27700 12021 27740
rect 11979 27691 12021 27700
rect 11692 27656 11732 27665
rect 11403 27404 11445 27413
rect 11403 27364 11404 27404
rect 11444 27364 11445 27404
rect 11403 27355 11445 27364
rect 11308 26816 11348 26825
rect 11308 26573 11348 26776
rect 11404 26816 11444 27355
rect 11404 26767 11444 26776
rect 11499 26816 11541 26825
rect 11499 26776 11500 26816
rect 11540 26776 11541 26816
rect 11499 26767 11541 26776
rect 11500 26682 11540 26767
rect 11403 26648 11445 26657
rect 11403 26608 11404 26648
rect 11444 26608 11445 26648
rect 11403 26599 11445 26608
rect 11596 26648 11636 26657
rect 11307 26564 11349 26573
rect 11307 26524 11308 26564
rect 11348 26524 11349 26564
rect 11307 26515 11349 26524
rect 11212 24760 11348 24800
rect 10924 24587 10964 24596
rect 10540 24573 10580 24582
rect 10539 24464 10581 24473
rect 10539 24424 10540 24464
rect 10580 24424 10581 24464
rect 10636 24464 10676 24582
rect 11116 24583 11156 24592
rect 11211 24632 11253 24641
rect 11211 24592 11212 24632
rect 11252 24592 11253 24632
rect 11211 24583 11253 24592
rect 10924 24464 10964 24547
rect 11212 24498 11252 24583
rect 10636 24424 10964 24464
rect 10539 24415 10581 24424
rect 10540 22625 10580 24415
rect 10828 24044 10868 24053
rect 10924 24044 10964 24424
rect 10868 24004 10964 24044
rect 10828 23995 10868 24004
rect 10635 23876 10677 23885
rect 10635 23836 10636 23876
rect 10676 23836 10677 23876
rect 10635 23827 10677 23836
rect 10636 23792 10676 23827
rect 10636 23633 10676 23752
rect 10635 23624 10677 23633
rect 10635 23584 10636 23624
rect 10676 23584 10677 23624
rect 10635 23575 10677 23584
rect 11211 23624 11253 23633
rect 11211 23584 11212 23624
rect 11252 23584 11253 23624
rect 11211 23575 11253 23584
rect 11019 23204 11061 23213
rect 11019 23164 11020 23204
rect 11060 23164 11061 23204
rect 11019 23155 11061 23164
rect 10635 23120 10677 23129
rect 10635 23080 10636 23120
rect 10676 23080 10677 23120
rect 10635 23071 10677 23080
rect 10636 22986 10676 23071
rect 10539 22616 10581 22625
rect 10539 22576 10540 22616
rect 10580 22576 10581 22616
rect 10539 22567 10581 22576
rect 11020 21944 11060 23155
rect 11212 22280 11252 23575
rect 11308 22373 11348 24760
rect 11404 23969 11444 26599
rect 11499 26480 11541 26489
rect 11499 26440 11500 26480
rect 11540 26440 11541 26480
rect 11499 26431 11541 26440
rect 11500 24800 11540 26431
rect 11596 25976 11636 26608
rect 11692 26153 11732 27616
rect 11884 26900 11924 26909
rect 11980 26900 12020 27691
rect 12076 27656 12116 27868
rect 12172 27824 12212 28288
rect 12363 28288 12364 28328
rect 12404 28288 12405 28328
rect 12363 28279 12405 28288
rect 12556 28328 12596 28456
rect 12556 28279 12596 28288
rect 12652 28328 12692 28337
rect 12364 28194 12404 28279
rect 12652 28169 12692 28288
rect 12459 28160 12501 28169
rect 12459 28120 12460 28160
rect 12500 28120 12501 28160
rect 12459 28111 12501 28120
rect 12651 28160 12693 28169
rect 12651 28120 12652 28160
rect 12692 28120 12693 28160
rect 12651 28111 12693 28120
rect 12460 28026 12500 28111
rect 12364 27824 12404 27833
rect 12172 27784 12364 27824
rect 12364 27775 12404 27784
rect 12459 27824 12501 27833
rect 12459 27784 12460 27824
rect 12500 27784 12501 27824
rect 12459 27775 12501 27784
rect 12076 27607 12116 27616
rect 12172 27656 12212 27667
rect 12172 27581 12212 27616
rect 12268 27656 12308 27665
rect 12460 27656 12500 27775
rect 12308 27616 12500 27656
rect 12171 27572 12213 27581
rect 12171 27532 12172 27572
rect 12212 27532 12213 27572
rect 12171 27523 12213 27532
rect 12075 27236 12117 27245
rect 12075 27196 12076 27236
rect 12116 27196 12117 27236
rect 12075 27187 12117 27196
rect 12076 26909 12116 27187
rect 11924 26860 12020 26900
rect 12075 26900 12117 26909
rect 12075 26860 12076 26900
rect 12116 26860 12117 26900
rect 11884 26851 11924 26860
rect 12075 26851 12117 26860
rect 11787 26816 11829 26825
rect 11787 26776 11788 26816
rect 11828 26776 11829 26816
rect 11787 26767 11829 26776
rect 11788 26682 11828 26767
rect 11691 26144 11733 26153
rect 11691 26104 11692 26144
rect 11732 26104 11733 26144
rect 11691 26095 11733 26104
rect 12076 26144 12116 26851
rect 12268 26825 12308 27616
rect 12555 27572 12597 27581
rect 12555 27532 12556 27572
rect 12596 27532 12597 27572
rect 12555 27523 12597 27532
rect 12459 27404 12501 27413
rect 12459 27364 12460 27404
rect 12500 27364 12501 27404
rect 12459 27355 12501 27364
rect 12363 26900 12405 26909
rect 12363 26860 12364 26900
rect 12404 26860 12405 26900
rect 12363 26851 12405 26860
rect 12267 26816 12309 26825
rect 12267 26776 12268 26816
rect 12308 26776 12309 26816
rect 12267 26767 12309 26776
rect 12364 26816 12404 26851
rect 11596 25936 12020 25976
rect 11595 25640 11637 25649
rect 11595 25600 11596 25640
rect 11636 25600 11637 25640
rect 11595 25591 11637 25600
rect 11596 25304 11636 25591
rect 11883 25472 11925 25481
rect 11883 25432 11884 25472
rect 11924 25432 11925 25472
rect 11883 25423 11925 25432
rect 11596 25255 11636 25264
rect 11884 25304 11924 25423
rect 11884 25255 11924 25264
rect 11980 25304 12020 25936
rect 11980 25255 12020 25264
rect 11500 24760 11636 24800
rect 11500 24632 11540 24641
rect 11403 23960 11445 23969
rect 11403 23920 11404 23960
rect 11444 23920 11445 23960
rect 11403 23911 11445 23920
rect 11404 23792 11444 23801
rect 11404 22457 11444 23752
rect 11500 23297 11540 24592
rect 11596 24548 11636 24760
rect 12076 24725 12116 26104
rect 12268 25892 12308 25901
rect 12268 25649 12308 25852
rect 12267 25640 12309 25649
rect 12267 25600 12268 25640
rect 12308 25600 12309 25640
rect 12267 25591 12309 25600
rect 12268 25472 12308 25481
rect 11691 24716 11733 24725
rect 12075 24716 12117 24725
rect 11691 24676 11692 24716
rect 11732 24676 11828 24716
rect 11691 24667 11733 24676
rect 11788 24632 11828 24676
rect 12075 24676 12076 24716
rect 12116 24676 12117 24716
rect 12075 24667 12117 24676
rect 11788 24583 11828 24592
rect 11883 24632 11925 24641
rect 11883 24592 11884 24632
rect 11924 24592 11925 24632
rect 11883 24583 11925 24592
rect 11596 24508 11732 24548
rect 11595 23960 11637 23969
rect 11595 23920 11596 23960
rect 11636 23920 11637 23960
rect 11595 23911 11637 23920
rect 11499 23288 11541 23297
rect 11499 23248 11500 23288
rect 11540 23248 11541 23288
rect 11499 23239 11541 23248
rect 11403 22448 11445 22457
rect 11403 22408 11404 22448
rect 11444 22408 11445 22448
rect 11403 22399 11445 22408
rect 11307 22364 11349 22373
rect 11307 22324 11308 22364
rect 11348 22324 11349 22364
rect 11307 22315 11349 22324
rect 11499 22364 11541 22373
rect 11499 22324 11500 22364
rect 11540 22324 11541 22364
rect 11499 22315 11541 22324
rect 11212 22231 11252 22240
rect 11404 22196 11444 22205
rect 11500 22196 11540 22315
rect 11444 22156 11540 22196
rect 11404 22147 11444 22156
rect 11596 22037 11636 23911
rect 11692 22952 11732 24508
rect 11884 24498 11924 24583
rect 12172 24380 12212 24389
rect 11883 23456 11925 23465
rect 11883 23416 11884 23456
rect 11924 23416 11925 23456
rect 11883 23407 11925 23416
rect 11884 23120 11924 23407
rect 12076 23297 12116 23382
rect 12075 23288 12117 23297
rect 12075 23248 12076 23288
rect 12116 23248 12117 23288
rect 12075 23239 12117 23248
rect 11884 23071 11924 23080
rect 11692 22912 11924 22952
rect 11787 22784 11829 22793
rect 11787 22744 11788 22784
rect 11828 22744 11829 22784
rect 11787 22735 11829 22744
rect 11691 22364 11733 22373
rect 11691 22324 11692 22364
rect 11732 22324 11733 22364
rect 11691 22315 11733 22324
rect 11692 22280 11732 22315
rect 11692 22229 11732 22240
rect 11595 22028 11637 22037
rect 11500 21988 11596 22028
rect 11636 21988 11637 22028
rect 11020 21904 11156 21944
rect 10732 21692 10772 21701
rect 10772 21652 11060 21692
rect 10732 21643 10772 21652
rect 10540 21608 10580 21617
rect 10540 21449 10580 21568
rect 11020 21608 11060 21652
rect 11020 21559 11060 21568
rect 11116 21608 11156 21904
rect 10539 21440 10581 21449
rect 10539 21400 10540 21440
rect 10580 21400 10581 21440
rect 10539 21391 10581 21400
rect 11116 20693 11156 21568
rect 11500 21608 11540 21988
rect 11595 21979 11637 21988
rect 11500 21559 11540 21568
rect 11595 21608 11637 21617
rect 11595 21568 11596 21608
rect 11636 21568 11637 21608
rect 11595 21559 11637 21568
rect 11596 21474 11636 21559
rect 11595 21188 11637 21197
rect 11595 21148 11596 21188
rect 11636 21148 11637 21188
rect 11595 21139 11637 21148
rect 11307 20768 11349 20777
rect 11307 20728 11308 20768
rect 11348 20728 11349 20768
rect 11307 20719 11349 20728
rect 11115 20684 11157 20693
rect 11115 20644 11116 20684
rect 11156 20644 11157 20684
rect 11115 20635 11157 20644
rect 11308 20634 11348 20719
rect 11596 20441 11636 21139
rect 11595 20432 11637 20441
rect 11595 20392 11596 20432
rect 11636 20392 11637 20432
rect 11595 20383 11637 20392
rect 10635 20264 10677 20273
rect 10635 20224 10636 20264
rect 10676 20224 10677 20264
rect 10635 20215 10677 20224
rect 10540 20096 10580 20105
rect 10540 19349 10580 20056
rect 10539 19340 10581 19349
rect 10539 19300 10540 19340
rect 10580 19300 10581 19340
rect 10539 19291 10581 19300
rect 10539 19088 10581 19097
rect 10539 19048 10540 19088
rect 10580 19048 10581 19088
rect 10539 19039 10581 19048
rect 10540 18341 10580 19039
rect 10539 18332 10581 18341
rect 10539 18292 10540 18332
rect 10580 18292 10581 18332
rect 10539 18283 10581 18292
rect 10444 17200 10580 17240
rect 10444 17072 10484 17083
rect 10444 16997 10484 17032
rect 10443 16988 10485 16997
rect 10443 16948 10444 16988
rect 10484 16948 10485 16988
rect 10443 16939 10485 16948
rect 9963 16652 10005 16661
rect 9963 16612 9964 16652
rect 10004 16612 10005 16652
rect 9963 16603 10005 16612
rect 9771 16528 9772 16568
rect 9812 16528 9908 16568
rect 9771 16519 9813 16528
rect 9484 16360 9908 16400
rect 9580 16232 9620 16241
rect 9387 15812 9429 15821
rect 9387 15772 9388 15812
rect 9428 15772 9524 15812
rect 9387 15763 9429 15772
rect 9387 15308 9429 15317
rect 9387 15268 9388 15308
rect 9428 15268 9429 15308
rect 9387 15259 9429 15268
rect 9388 14720 9428 15259
rect 9484 14804 9524 15772
rect 9580 14972 9620 16192
rect 9676 16232 9716 16243
rect 9676 16157 9716 16192
rect 9675 16148 9717 16157
rect 9675 16108 9676 16148
rect 9716 16108 9717 16148
rect 9675 16099 9717 16108
rect 9771 16064 9813 16073
rect 9771 16024 9772 16064
rect 9812 16024 9813 16064
rect 9771 16015 9813 16024
rect 9580 14923 9620 14932
rect 9772 15560 9812 16015
rect 9484 14764 9716 14804
rect 9388 14671 9428 14680
rect 9196 14512 9620 14552
rect 9195 12620 9237 12629
rect 9195 12580 9196 12620
rect 9236 12580 9237 12620
rect 9195 12571 9237 12580
rect 9196 12536 9236 12571
rect 9196 12485 9236 12496
rect 9292 12536 9332 12545
rect 9332 12496 9524 12536
rect 9292 12487 9332 12496
rect 9195 11024 9237 11033
rect 9195 10984 9196 11024
rect 9236 10984 9237 11024
rect 9195 10975 9237 10984
rect 9099 10352 9141 10361
rect 9099 10312 9100 10352
rect 9140 10312 9141 10352
rect 9099 10303 9141 10312
rect 9004 10135 9044 10144
rect 8812 9640 9044 9680
rect 8812 9512 8852 9521
rect 8715 8756 8757 8765
rect 8715 8716 8716 8756
rect 8756 8716 8757 8756
rect 8715 8707 8757 8716
rect 8716 8672 8756 8707
rect 8716 8621 8756 8632
rect 8812 7589 8852 9472
rect 8908 9512 8948 9521
rect 8908 8849 8948 9472
rect 8907 8840 8949 8849
rect 8907 8800 8908 8840
rect 8948 8800 8949 8840
rect 8907 8791 8949 8800
rect 9004 8168 9044 9640
rect 9196 9512 9236 10975
rect 9387 10268 9429 10277
rect 9387 10228 9388 10268
rect 9428 10228 9429 10268
rect 9387 10219 9429 10228
rect 9291 10184 9333 10193
rect 9291 10144 9292 10184
rect 9332 10144 9333 10184
rect 9291 10135 9333 10144
rect 9196 9463 9236 9472
rect 8908 8128 9044 8168
rect 8811 7580 8853 7589
rect 8811 7540 8812 7580
rect 8852 7540 8853 7580
rect 8811 7531 8853 7540
rect 8908 7202 8948 8128
rect 9003 8000 9045 8009
rect 9003 7960 9004 8000
rect 9044 7960 9045 8000
rect 9003 7951 9045 7960
rect 9004 7866 9044 7951
rect 9196 7748 9236 7757
rect 9196 7253 9236 7708
rect 8811 7165 8853 7169
rect 8811 7162 8908 7165
rect 9195 7244 9237 7253
rect 9195 7204 9196 7244
rect 9236 7204 9237 7244
rect 9195 7195 9237 7204
rect 8948 7162 9140 7165
rect 8811 7160 9140 7162
rect 8811 7120 8812 7160
rect 8852 7125 9140 7160
rect 8852 7120 8853 7125
rect 8811 7111 8853 7120
rect 8524 7036 8756 7076
rect 8235 6992 8277 7001
rect 8235 6952 8236 6992
rect 8276 6952 8277 6992
rect 8235 6943 8277 6952
rect 8427 6908 8469 6917
rect 8427 6868 8428 6908
rect 8468 6868 8469 6908
rect 8427 6859 8469 6868
rect 8140 6784 8276 6824
rect 8139 5900 8181 5909
rect 8139 5860 8140 5900
rect 8180 5860 8181 5900
rect 8139 5851 8181 5860
rect 8140 5766 8180 5851
rect 8139 5648 8181 5657
rect 8139 5608 8140 5648
rect 8180 5608 8181 5648
rect 8139 5599 8181 5608
rect 8043 5396 8085 5405
rect 8043 5356 8044 5396
rect 8084 5356 8085 5396
rect 8043 5347 8085 5356
rect 7796 5104 7892 5144
rect 7756 5095 7796 5104
rect 7755 4892 7797 4901
rect 7755 4852 7756 4892
rect 7796 4852 7797 4892
rect 7755 4843 7797 4852
rect 7468 4087 7508 4096
rect 7564 4180 7700 4220
rect 7468 3632 7508 3641
rect 7372 3592 7468 3632
rect 7468 3583 7508 3592
rect 7276 3464 7316 3475
rect 7276 3389 7316 3424
rect 7467 3464 7509 3473
rect 7467 3424 7468 3464
rect 7508 3424 7509 3464
rect 7467 3415 7509 3424
rect 7275 3380 7317 3389
rect 7275 3340 7276 3380
rect 7316 3340 7317 3380
rect 7275 3331 7317 3340
rect 7180 2491 7220 2500
rect 7084 1240 7220 1280
rect 6987 1231 7029 1240
rect 6604 1063 6644 1072
rect 6603 944 6645 953
rect 6603 904 6604 944
rect 6644 904 6645 944
rect 6603 895 6645 904
rect 6604 80 6644 895
rect 6795 776 6837 785
rect 6795 736 6796 776
rect 6836 736 6837 776
rect 6795 727 6837 736
rect 6796 80 6836 727
rect 6988 80 7028 1231
rect 7180 80 7220 1240
rect 7371 1196 7413 1205
rect 7371 1156 7372 1196
rect 7412 1156 7413 1196
rect 7371 1147 7413 1156
rect 7468 1196 7508 3415
rect 7468 1147 7508 1156
rect 7372 80 7412 1147
rect 7564 80 7604 4180
rect 7756 3464 7796 4843
rect 7947 4724 7989 4733
rect 7947 4684 7948 4724
rect 7988 4684 7989 4724
rect 7947 4675 7989 4684
rect 7851 4304 7893 4313
rect 7851 4264 7852 4304
rect 7892 4264 7893 4304
rect 7851 4255 7893 4264
rect 7852 4220 7892 4255
rect 7852 4169 7892 4180
rect 7948 4220 7988 4675
rect 7948 4171 7988 4180
rect 7756 3415 7796 3424
rect 7659 2876 7701 2885
rect 7659 2836 7660 2876
rect 7700 2836 7701 2876
rect 7659 2827 7701 2836
rect 8043 2876 8085 2885
rect 8043 2836 8044 2876
rect 8084 2836 8085 2876
rect 8043 2827 8085 2836
rect 7660 2742 7700 2827
rect 8044 2742 8084 2827
rect 7852 2708 7892 2717
rect 7852 2540 7892 2668
rect 7756 2500 7892 2540
rect 7659 2204 7701 2213
rect 7659 2164 7660 2204
rect 7700 2164 7701 2204
rect 7659 2155 7701 2164
rect 7660 1952 7700 2155
rect 7660 1373 7700 1912
rect 7756 1448 7796 2500
rect 8140 2213 8180 5599
rect 8236 4808 8276 6784
rect 8428 6656 8468 6859
rect 8428 6607 8468 6616
rect 8572 6446 8612 6455
rect 8572 6404 8612 6406
rect 8332 6364 8612 6404
rect 8332 5900 8372 6364
rect 8332 5851 8372 5860
rect 8524 5648 8564 5659
rect 8524 5573 8564 5608
rect 8523 5564 8565 5573
rect 8523 5524 8524 5564
rect 8564 5524 8565 5564
rect 8523 5515 8565 5524
rect 8332 4985 8372 5070
rect 8331 4976 8373 4985
rect 8331 4936 8332 4976
rect 8372 4936 8373 4976
rect 8331 4927 8373 4936
rect 8427 4808 8469 4817
rect 8236 4768 8372 4808
rect 8236 2708 8276 2717
rect 8236 2540 8276 2668
rect 8332 2624 8372 4768
rect 8427 4768 8428 4808
rect 8468 4768 8469 4808
rect 8427 4759 8469 4768
rect 8428 4136 8468 4759
rect 8428 3977 8468 4096
rect 8427 3968 8469 3977
rect 8427 3928 8428 3968
rect 8468 3928 8469 3968
rect 8427 3919 8469 3928
rect 8716 3800 8756 7036
rect 8811 6992 8853 7001
rect 8811 6952 8812 6992
rect 8852 6952 8853 6992
rect 8811 6943 8853 6952
rect 8812 5825 8852 6943
rect 8907 6908 8949 6917
rect 8907 6868 8908 6908
rect 8948 6868 8949 6908
rect 8907 6859 8949 6868
rect 8811 5816 8853 5825
rect 8811 5776 8812 5816
rect 8852 5776 8853 5816
rect 8811 5767 8853 5776
rect 8908 5648 8948 6859
rect 9100 6488 9140 7125
rect 9100 6439 9140 6448
rect 8428 3760 8756 3800
rect 8812 5608 8948 5648
rect 8428 2719 8468 3760
rect 8428 2670 8468 2679
rect 8332 2584 8468 2624
rect 8428 2540 8468 2584
rect 8715 2540 8757 2549
rect 8236 2500 8372 2540
rect 8428 2500 8564 2540
rect 8235 2288 8277 2297
rect 8235 2248 8236 2288
rect 8276 2248 8277 2288
rect 8235 2239 8277 2248
rect 8139 2204 8181 2213
rect 8139 2164 8140 2204
rect 8180 2164 8181 2204
rect 8139 2155 8181 2164
rect 7852 2036 7892 2045
rect 7892 1996 8180 2036
rect 7852 1987 7892 1996
rect 8140 1952 8180 1996
rect 8140 1903 8180 1912
rect 8236 1952 8276 2239
rect 8236 1903 8276 1912
rect 7756 1408 8180 1448
rect 7659 1364 7701 1373
rect 7659 1324 7660 1364
rect 7700 1324 7701 1364
rect 7659 1315 7701 1324
rect 7851 1280 7893 1289
rect 7851 1240 7852 1280
rect 7892 1240 7893 1280
rect 7851 1231 7893 1240
rect 7852 1146 7892 1231
rect 7947 1196 7989 1205
rect 7947 1156 7948 1196
rect 7988 1156 7989 1196
rect 7947 1147 7989 1156
rect 8044 1196 8084 1205
rect 7659 944 7701 953
rect 7659 904 7660 944
rect 7700 904 7701 944
rect 7659 895 7701 904
rect 7660 810 7700 895
rect 7755 692 7797 701
rect 7755 652 7756 692
rect 7796 652 7797 692
rect 7755 643 7797 652
rect 7756 80 7796 643
rect 7948 80 7988 1147
rect 8044 617 8084 1156
rect 8043 608 8085 617
rect 8043 568 8044 608
rect 8084 568 8085 608
rect 8043 559 8085 568
rect 8140 80 8180 1408
rect 8236 1112 8276 1121
rect 8236 785 8276 1072
rect 8332 1028 8372 2500
rect 8524 1373 8564 2500
rect 8715 2500 8716 2540
rect 8756 2500 8757 2540
rect 8715 2491 8757 2500
rect 8619 2456 8661 2465
rect 8619 2416 8620 2456
rect 8660 2416 8661 2456
rect 8619 2407 8661 2416
rect 8620 2322 8660 2407
rect 8716 2381 8756 2491
rect 8715 2372 8757 2381
rect 8715 2332 8716 2372
rect 8756 2332 8757 2372
rect 8715 2323 8757 2332
rect 8716 1952 8756 2323
rect 8716 1903 8756 1912
rect 8620 1868 8660 1877
rect 8523 1364 8565 1373
rect 8523 1324 8524 1364
rect 8564 1324 8565 1364
rect 8523 1315 8565 1324
rect 8332 988 8564 1028
rect 8235 776 8277 785
rect 8235 736 8236 776
rect 8276 736 8277 776
rect 8235 727 8277 736
rect 8331 608 8373 617
rect 8331 568 8332 608
rect 8372 568 8373 608
rect 8331 559 8373 568
rect 8332 80 8372 559
rect 8524 80 8564 988
rect 8620 869 8660 1828
rect 8715 944 8757 953
rect 8715 904 8716 944
rect 8756 904 8757 944
rect 8715 895 8757 904
rect 8619 860 8661 869
rect 8619 820 8620 860
rect 8660 820 8661 860
rect 8619 811 8661 820
rect 8716 80 8756 895
rect 8812 701 8852 5608
rect 8956 4145 8996 4154
rect 8996 4105 9236 4136
rect 8956 4096 9236 4105
rect 9100 3968 9140 3977
rect 9003 3464 9045 3473
rect 9003 3424 9004 3464
rect 9044 3424 9045 3464
rect 9003 3415 9045 3424
rect 9004 3330 9044 3415
rect 9100 1709 9140 3928
rect 9196 3632 9236 4096
rect 9196 3583 9236 3592
rect 9292 2708 9332 10135
rect 9388 10134 9428 10219
rect 9484 10193 9524 12496
rect 9580 11201 9620 14512
rect 9676 12536 9716 14764
rect 9772 12629 9812 15520
rect 9771 12620 9813 12629
rect 9771 12580 9772 12620
rect 9812 12580 9813 12620
rect 9771 12571 9813 12580
rect 9868 12545 9908 16360
rect 10060 16232 10100 16241
rect 9963 15308 10005 15317
rect 9963 15268 9964 15308
rect 10004 15268 10005 15308
rect 9963 15259 10005 15268
rect 9964 13208 10004 15259
rect 10060 15149 10100 16192
rect 10155 16232 10197 16241
rect 10155 16192 10156 16232
rect 10196 16192 10197 16232
rect 10155 16183 10197 16192
rect 10156 15401 10196 16183
rect 10251 16148 10293 16157
rect 10251 16108 10252 16148
rect 10292 16108 10293 16148
rect 10251 16099 10293 16108
rect 10155 15392 10197 15401
rect 10155 15352 10156 15392
rect 10196 15352 10197 15392
rect 10155 15343 10197 15352
rect 10059 15140 10101 15149
rect 10059 15100 10060 15140
rect 10100 15100 10101 15140
rect 10059 15091 10101 15100
rect 10156 14720 10196 14729
rect 10060 14680 10156 14720
rect 10060 13880 10100 14680
rect 10156 14671 10196 14680
rect 10252 14720 10292 16099
rect 10540 15905 10580 17200
rect 10636 16232 10676 20215
rect 10732 20180 10772 20189
rect 11115 20180 11157 20189
rect 10772 20140 11060 20180
rect 10732 20131 10772 20140
rect 11020 20096 11060 20140
rect 11115 20140 11116 20180
rect 11156 20140 11157 20180
rect 11115 20131 11157 20140
rect 11020 20047 11060 20056
rect 11116 20096 11156 20131
rect 11116 19928 11156 20056
rect 11596 20096 11636 20383
rect 11596 20047 11636 20056
rect 11500 20012 11540 20023
rect 11500 19937 11540 19972
rect 11020 19888 11156 19928
rect 11499 19928 11541 19937
rect 11499 19888 11500 19928
rect 11540 19888 11541 19928
rect 10923 18836 10965 18845
rect 10923 18796 10924 18836
rect 10964 18796 10965 18836
rect 10923 18787 10965 18796
rect 10731 18164 10773 18173
rect 10731 18124 10732 18164
rect 10772 18124 10773 18164
rect 10731 18115 10773 18124
rect 10732 17744 10772 18115
rect 10827 18080 10869 18089
rect 10827 18040 10828 18080
rect 10868 18040 10869 18080
rect 10827 18031 10869 18040
rect 10732 17695 10772 17704
rect 10828 16316 10868 18031
rect 10539 15896 10581 15905
rect 10539 15856 10540 15896
rect 10580 15856 10581 15896
rect 10539 15847 10581 15856
rect 10636 15821 10676 16192
rect 10732 16276 10868 16316
rect 10635 15812 10677 15821
rect 10635 15772 10636 15812
rect 10676 15772 10677 15812
rect 10635 15763 10677 15772
rect 10732 15560 10772 16276
rect 10827 15812 10869 15821
rect 10827 15772 10828 15812
rect 10868 15772 10869 15812
rect 10827 15763 10869 15772
rect 10636 15520 10772 15560
rect 10636 15485 10676 15520
rect 10347 15476 10389 15485
rect 10347 15436 10348 15476
rect 10388 15436 10389 15476
rect 10347 15427 10389 15436
rect 10634 15476 10676 15485
rect 10634 15436 10635 15476
rect 10675 15436 10676 15476
rect 10634 15427 10676 15436
rect 10156 14057 10196 14142
rect 10155 14048 10197 14057
rect 10155 14008 10156 14048
rect 10196 14008 10197 14048
rect 10155 13999 10197 14008
rect 10252 14048 10292 14680
rect 10060 13840 10196 13880
rect 10059 13628 10101 13637
rect 10059 13588 10060 13628
rect 10100 13588 10101 13628
rect 10059 13579 10101 13588
rect 9964 13159 10004 13168
rect 9579 11192 9621 11201
rect 9579 11152 9580 11192
rect 9620 11152 9621 11192
rect 9579 11143 9621 11152
rect 9579 11024 9621 11033
rect 9579 10984 9580 11024
rect 9620 10984 9621 11024
rect 9579 10975 9621 10984
rect 9580 10890 9620 10975
rect 9579 10520 9621 10529
rect 9579 10480 9580 10520
rect 9620 10480 9621 10520
rect 9579 10471 9621 10480
rect 9483 10184 9525 10193
rect 9483 10144 9484 10184
rect 9524 10144 9525 10184
rect 9483 10135 9525 10144
rect 9484 10050 9524 10135
rect 9483 9848 9525 9857
rect 9483 9808 9484 9848
rect 9524 9808 9525 9848
rect 9483 9799 9525 9808
rect 9388 8000 9428 8009
rect 9388 7841 9428 7960
rect 9387 7832 9429 7841
rect 9387 7792 9388 7832
rect 9428 7792 9429 7832
rect 9387 7783 9429 7792
rect 9387 7580 9429 7589
rect 9387 7540 9388 7580
rect 9428 7540 9429 7580
rect 9387 7531 9429 7540
rect 9388 7244 9428 7531
rect 9484 7328 9524 9799
rect 9580 7841 9620 10471
rect 9676 10277 9716 12496
rect 9867 12536 9909 12545
rect 9867 12496 9868 12536
rect 9908 12496 9909 12536
rect 9867 12487 9909 12496
rect 9771 12452 9813 12461
rect 9771 12412 9772 12452
rect 9812 12412 9813 12452
rect 9771 12403 9813 12412
rect 9772 12318 9812 12403
rect 10060 11948 10100 13579
rect 10156 13460 10196 13840
rect 10156 13411 10196 13420
rect 10252 13208 10292 14008
rect 10156 13168 10292 13208
rect 10156 12368 10196 13168
rect 10252 12545 10292 12630
rect 10251 12536 10293 12545
rect 10251 12496 10252 12536
rect 10292 12496 10293 12536
rect 10251 12487 10293 12496
rect 10156 12328 10292 12368
rect 10156 11948 10196 11957
rect 10060 11908 10156 11948
rect 10156 11899 10196 11908
rect 9964 11789 10004 11833
rect 9771 11780 9813 11789
rect 9771 11740 9772 11780
rect 9812 11740 9813 11780
rect 9771 11731 9813 11740
rect 9963 11780 10005 11789
rect 9963 11740 9964 11780
rect 10004 11740 10005 11780
rect 9963 11738 10005 11740
rect 9963 11731 9964 11738
rect 9675 10268 9717 10277
rect 9675 10228 9676 10268
rect 9716 10228 9717 10268
rect 9675 10219 9717 10228
rect 9772 8840 9812 11731
rect 10004 11731 10005 11738
rect 9964 11689 10004 11698
rect 9867 11528 9909 11537
rect 9867 11488 9868 11528
rect 9908 11488 9909 11528
rect 9867 11479 9909 11488
rect 9676 8800 9812 8840
rect 9676 8084 9716 8800
rect 9868 8765 9908 11479
rect 10059 11108 10101 11117
rect 10059 11068 10060 11108
rect 10100 11068 10101 11108
rect 10059 11059 10101 11068
rect 10060 10445 10100 11059
rect 10155 10604 10197 10613
rect 10155 10564 10156 10604
rect 10196 10564 10197 10604
rect 10155 10555 10197 10564
rect 10059 10436 10101 10445
rect 10059 10396 10060 10436
rect 10100 10396 10101 10436
rect 10059 10387 10101 10396
rect 9963 10352 10005 10361
rect 9963 10312 9964 10352
rect 10004 10312 10005 10352
rect 9963 10303 10005 10312
rect 9964 10184 10004 10303
rect 9964 10135 10004 10144
rect 9867 8756 9909 8765
rect 9867 8716 9868 8756
rect 9908 8716 9909 8756
rect 9867 8707 9909 8716
rect 9772 8672 9812 8681
rect 9772 8588 9812 8632
rect 9868 8588 9908 8707
rect 9772 8548 9908 8588
rect 9676 8044 9908 8084
rect 9579 7832 9621 7841
rect 9579 7792 9580 7832
rect 9620 7792 9621 7832
rect 9579 7783 9621 7792
rect 9771 7832 9813 7841
rect 9771 7792 9772 7832
rect 9812 7792 9813 7832
rect 9771 7783 9813 7792
rect 9484 7288 9620 7328
rect 9388 7195 9428 7204
rect 9484 7160 9524 7169
rect 9387 7076 9429 7085
rect 9484 7076 9524 7120
rect 9387 7036 9388 7076
rect 9428 7036 9524 7076
rect 9387 7027 9429 7036
rect 9484 6908 9524 7036
rect 9388 6868 9524 6908
rect 9388 6581 9428 6868
rect 9580 6656 9620 7288
rect 9484 6616 9620 6656
rect 9387 6572 9429 6581
rect 9387 6532 9388 6572
rect 9428 6532 9429 6572
rect 9387 6523 9429 6532
rect 9484 4976 9524 6616
rect 9675 6572 9717 6581
rect 9675 6532 9676 6572
rect 9716 6532 9717 6572
rect 9675 6523 9717 6532
rect 9579 6488 9621 6497
rect 9579 6448 9580 6488
rect 9620 6448 9621 6488
rect 9579 6439 9621 6448
rect 9676 6488 9716 6523
rect 9580 6404 9620 6439
rect 9676 6437 9716 6448
rect 9580 6353 9620 6364
rect 9675 6236 9717 6245
rect 9675 6196 9676 6236
rect 9716 6196 9717 6236
rect 9675 6187 9717 6196
rect 9676 5573 9716 6187
rect 9772 5648 9812 7783
rect 9868 7505 9908 8044
rect 9963 7748 10005 7757
rect 9963 7708 9964 7748
rect 10004 7708 10005 7748
rect 9963 7699 10005 7708
rect 9867 7496 9909 7505
rect 9867 7456 9868 7496
rect 9908 7456 9909 7496
rect 9867 7447 9909 7456
rect 9867 7160 9909 7169
rect 9867 7120 9868 7160
rect 9908 7120 9909 7160
rect 9867 7111 9909 7120
rect 9964 7160 10004 7699
rect 10059 7580 10101 7589
rect 10059 7540 10060 7580
rect 10100 7540 10101 7580
rect 10059 7531 10101 7540
rect 9964 7111 10004 7120
rect 9868 7026 9908 7111
rect 10060 6488 10100 7531
rect 10156 7169 10196 10555
rect 10155 7160 10197 7169
rect 10155 7120 10156 7160
rect 10196 7120 10197 7160
rect 10155 7111 10197 7120
rect 10060 6439 10100 6448
rect 10156 6488 10196 6497
rect 10156 5909 10196 6448
rect 10155 5900 10197 5909
rect 10155 5860 10156 5900
rect 10196 5860 10197 5900
rect 10155 5851 10197 5860
rect 9675 5564 9717 5573
rect 9675 5524 9676 5564
rect 9716 5524 9717 5564
rect 9675 5515 9717 5524
rect 9579 4976 9621 4985
rect 9484 4936 9580 4976
rect 9620 4936 9621 4976
rect 9579 4927 9621 4936
rect 9580 4842 9620 4927
rect 9580 3464 9620 3473
rect 9676 3464 9716 5515
rect 9772 4901 9812 5608
rect 9963 5648 10005 5657
rect 9963 5608 9964 5648
rect 10004 5608 10005 5648
rect 9963 5599 10005 5608
rect 9964 5514 10004 5599
rect 9964 4976 10004 4985
rect 9771 4892 9813 4901
rect 9771 4852 9772 4892
rect 9812 4852 9813 4892
rect 9771 4843 9813 4852
rect 9772 4724 9812 4733
rect 9772 4145 9812 4684
rect 9964 4649 10004 4936
rect 9963 4640 10005 4649
rect 9963 4600 9964 4640
rect 10004 4600 10005 4640
rect 9963 4591 10005 4600
rect 9771 4136 9813 4145
rect 9771 4096 9772 4136
rect 9812 4096 9813 4136
rect 9771 4087 9813 4096
rect 10155 4136 10197 4145
rect 10155 4096 10156 4136
rect 10196 4096 10197 4136
rect 10155 4087 10197 4096
rect 10252 4136 10292 12328
rect 10348 11696 10388 15427
rect 10731 15392 10773 15401
rect 10731 15352 10732 15392
rect 10772 15352 10773 15392
rect 10731 15343 10773 15352
rect 10635 15140 10677 15149
rect 10635 15100 10636 15140
rect 10676 15100 10677 15140
rect 10635 15091 10677 15100
rect 10636 14720 10676 15091
rect 10636 14048 10676 14680
rect 10636 13999 10676 14008
rect 10732 14804 10772 15343
rect 10732 14048 10772 14764
rect 10828 14729 10868 15763
rect 10827 14720 10869 14729
rect 10827 14680 10828 14720
rect 10868 14680 10869 14720
rect 10827 14671 10869 14680
rect 10732 13208 10772 14008
rect 10924 13217 10964 18787
rect 11020 16913 11060 19888
rect 11499 19879 11541 19888
rect 11595 19844 11637 19853
rect 11595 19804 11596 19844
rect 11636 19804 11637 19844
rect 11595 19795 11637 19804
rect 11307 19340 11349 19349
rect 11307 19300 11308 19340
rect 11348 19300 11349 19340
rect 11307 19291 11349 19300
rect 11116 19256 11156 19267
rect 11116 19181 11156 19216
rect 11115 19172 11157 19181
rect 11115 19132 11116 19172
rect 11156 19132 11157 19172
rect 11115 19123 11157 19132
rect 11308 18584 11348 19291
rect 11116 18544 11308 18584
rect 11116 17081 11156 18544
rect 11308 18535 11348 18544
rect 11500 18332 11540 18341
rect 11308 18292 11500 18332
rect 11308 17828 11348 18292
rect 11500 18283 11540 18292
rect 11260 17788 11348 17828
rect 11260 17786 11300 17788
rect 11260 17737 11300 17746
rect 11403 17660 11445 17669
rect 11403 17620 11404 17660
rect 11444 17620 11445 17660
rect 11403 17611 11445 17620
rect 11404 17526 11444 17611
rect 11115 17072 11157 17081
rect 11115 17032 11116 17072
rect 11156 17032 11157 17072
rect 11115 17023 11157 17032
rect 11019 16904 11061 16913
rect 11019 16864 11020 16904
rect 11060 16864 11061 16904
rect 11019 16855 11061 16864
rect 11164 16241 11204 16250
rect 11596 16232 11636 19795
rect 11788 19088 11828 22735
rect 11884 20021 11924 22912
rect 11979 22280 12021 22289
rect 11979 22240 11980 22280
rect 12020 22240 12021 22280
rect 11979 22231 12021 22240
rect 11980 22146 12020 22231
rect 12076 22196 12116 22205
rect 12076 21776 12116 22156
rect 11980 21736 12116 21776
rect 11980 20609 12020 21736
rect 12076 21608 12116 21619
rect 12076 21533 12116 21568
rect 12075 21524 12117 21533
rect 12075 21484 12076 21524
rect 12116 21484 12117 21524
rect 12075 21475 12117 21484
rect 11979 20600 12021 20609
rect 11979 20560 11980 20600
rect 12020 20560 12021 20600
rect 11979 20551 12021 20560
rect 12172 20525 12212 24340
rect 12268 22121 12308 25432
rect 12364 25229 12404 26776
rect 12363 25220 12405 25229
rect 12363 25180 12364 25220
rect 12404 25180 12405 25220
rect 12363 25171 12405 25180
rect 12364 22448 12404 22457
rect 12267 22112 12309 22121
rect 12267 22072 12268 22112
rect 12308 22072 12309 22112
rect 12267 22063 12309 22072
rect 12267 21104 12309 21113
rect 12267 21064 12268 21104
rect 12308 21064 12309 21104
rect 12267 21055 12309 21064
rect 12268 20777 12308 21055
rect 12364 20945 12404 22408
rect 12363 20936 12405 20945
rect 12363 20896 12364 20936
rect 12404 20896 12405 20936
rect 12363 20887 12405 20896
rect 12267 20768 12309 20777
rect 12267 20728 12268 20768
rect 12308 20728 12309 20768
rect 12267 20719 12309 20728
rect 12171 20516 12213 20525
rect 12171 20476 12172 20516
rect 12212 20476 12213 20516
rect 12171 20467 12213 20476
rect 12076 20096 12116 20105
rect 11883 20012 11925 20021
rect 11883 19972 11884 20012
rect 11924 19972 11925 20012
rect 11883 19963 11925 19972
rect 11692 19048 11828 19088
rect 11692 17165 11732 19048
rect 11787 18920 11829 18929
rect 11787 18880 11788 18920
rect 11828 18880 11829 18920
rect 11787 18871 11829 18880
rect 11691 17156 11733 17165
rect 11691 17116 11692 17156
rect 11732 17116 11733 17156
rect 11691 17107 11733 17116
rect 11788 17072 11828 18871
rect 11884 18005 11924 19963
rect 12076 19853 12116 20056
rect 12171 19928 12213 19937
rect 12171 19888 12172 19928
rect 12212 19888 12213 19928
rect 12171 19879 12213 19888
rect 12075 19844 12117 19853
rect 12075 19804 12076 19844
rect 12116 19804 12117 19844
rect 12075 19795 12117 19804
rect 12075 19508 12117 19517
rect 12075 19468 12076 19508
rect 12116 19468 12117 19508
rect 12075 19459 12117 19468
rect 11979 18584 12021 18593
rect 11979 18544 11980 18584
rect 12020 18544 12021 18584
rect 11979 18535 12021 18544
rect 12076 18584 12116 19459
rect 12076 18535 12116 18544
rect 11883 17996 11925 18005
rect 11883 17956 11884 17996
rect 11924 17956 11925 17996
rect 11883 17947 11925 17956
rect 11884 17669 11924 17947
rect 11883 17660 11925 17669
rect 11883 17620 11884 17660
rect 11924 17620 11925 17660
rect 11883 17611 11925 17620
rect 11980 17501 12020 18535
rect 12172 18416 12212 19879
rect 12076 18376 12212 18416
rect 12076 17921 12116 18376
rect 12075 17912 12117 17921
rect 12075 17872 12076 17912
rect 12116 17872 12117 17912
rect 12075 17863 12117 17872
rect 12171 17828 12213 17837
rect 12171 17788 12172 17828
rect 12212 17788 12213 17828
rect 12171 17779 12213 17788
rect 12076 17744 12116 17753
rect 11979 17492 12021 17501
rect 11979 17452 11980 17492
rect 12020 17452 12021 17492
rect 11979 17443 12021 17452
rect 12076 17324 12116 17704
rect 12172 17744 12212 17779
rect 12172 17693 12212 17704
rect 11884 17284 12116 17324
rect 11884 17240 11924 17284
rect 11884 17191 11924 17200
rect 12076 17072 12116 17081
rect 11692 17030 11732 17039
rect 11788 17032 12076 17072
rect 11692 16988 11732 16990
rect 11692 16948 11828 16988
rect 11691 16820 11733 16829
rect 11691 16780 11692 16820
rect 11732 16780 11733 16820
rect 11691 16771 11733 16780
rect 11204 16201 11252 16232
rect 11164 16192 11252 16201
rect 11115 15896 11157 15905
rect 11115 15856 11116 15896
rect 11156 15856 11157 15896
rect 11115 15847 11157 15856
rect 11020 15653 11060 15684
rect 11019 15644 11061 15653
rect 11019 15604 11020 15644
rect 11060 15604 11061 15644
rect 11019 15595 11061 15604
rect 11020 15560 11060 15595
rect 11020 15317 11060 15520
rect 11019 15308 11061 15317
rect 11019 15268 11020 15308
rect 11060 15268 11061 15308
rect 11019 15259 11061 15268
rect 10348 11033 10388 11656
rect 10636 13168 10772 13208
rect 10923 13208 10965 13217
rect 10923 13168 10924 13208
rect 10964 13168 10965 13208
rect 10636 11360 10676 13168
rect 10923 13159 10965 13168
rect 10924 13074 10964 13159
rect 10923 12704 10965 12713
rect 10923 12664 10924 12704
rect 10964 12664 10965 12704
rect 10923 12655 10965 12664
rect 10924 12570 10964 12655
rect 10780 12526 10820 12535
rect 10820 12486 11060 12526
rect 10780 12477 10820 12486
rect 10923 11612 10965 11621
rect 10923 11572 10924 11612
rect 10964 11572 10965 11612
rect 10923 11563 10965 11572
rect 10636 11320 10772 11360
rect 10347 11024 10389 11033
rect 10347 10984 10348 11024
rect 10388 10984 10389 11024
rect 10347 10975 10389 10984
rect 10539 10688 10581 10697
rect 10539 10648 10540 10688
rect 10580 10648 10581 10688
rect 10539 10639 10581 10648
rect 10540 10361 10580 10639
rect 10539 10352 10581 10361
rect 10539 10312 10540 10352
rect 10580 10312 10581 10352
rect 10539 10303 10581 10312
rect 10492 10193 10532 10202
rect 10532 10153 10580 10184
rect 10492 10144 10580 10153
rect 10443 10016 10485 10025
rect 10443 9976 10444 10016
rect 10484 9976 10485 10016
rect 10443 9967 10485 9976
rect 10444 9512 10484 9967
rect 10540 9680 10580 10144
rect 10635 10016 10677 10025
rect 10635 9976 10636 10016
rect 10676 9976 10677 10016
rect 10635 9967 10677 9976
rect 10636 9882 10676 9967
rect 10636 9680 10676 9689
rect 10540 9640 10636 9680
rect 10636 9631 10676 9640
rect 10484 9472 10676 9512
rect 10444 9463 10484 9472
rect 10539 9344 10581 9353
rect 10539 9304 10540 9344
rect 10580 9304 10581 9344
rect 10539 9295 10581 9304
rect 10443 7160 10485 7169
rect 10443 7120 10444 7160
rect 10484 7120 10485 7160
rect 10443 7111 10485 7120
rect 10444 4313 10484 7111
rect 10443 4304 10485 4313
rect 10443 4264 10444 4304
rect 10484 4264 10485 4304
rect 10443 4255 10485 4264
rect 10156 4002 10196 4087
rect 9620 3424 9716 3464
rect 9580 3415 9620 3424
rect 9867 3380 9909 3389
rect 9867 3340 9868 3380
rect 9908 3340 9909 3380
rect 9867 3331 9909 3340
rect 9388 2708 9428 2717
rect 9292 2668 9388 2708
rect 9388 2659 9428 2668
rect 9771 2708 9813 2717
rect 9771 2668 9772 2708
rect 9812 2668 9813 2708
rect 9771 2659 9813 2668
rect 9772 2574 9812 2659
rect 9291 2456 9333 2465
rect 9291 2416 9292 2456
rect 9332 2416 9333 2456
rect 9291 2407 9333 2416
rect 9580 2456 9620 2465
rect 9195 1952 9237 1961
rect 9195 1912 9196 1952
rect 9236 1912 9237 1952
rect 9195 1903 9237 1912
rect 9196 1818 9236 1903
rect 9099 1700 9141 1709
rect 9099 1660 9100 1700
rect 9140 1660 9141 1700
rect 9099 1651 9141 1660
rect 8907 776 8949 785
rect 8907 736 8908 776
rect 8948 736 8949 776
rect 8907 727 8949 736
rect 8811 692 8853 701
rect 8811 652 8812 692
rect 8852 652 8853 692
rect 8811 643 8853 652
rect 8908 80 8948 727
rect 9099 608 9141 617
rect 9099 568 9100 608
rect 9140 568 9141 608
rect 9099 559 9141 568
rect 9100 80 9140 559
rect 9292 80 9332 2407
rect 9580 2297 9620 2416
rect 9579 2288 9621 2297
rect 9579 2248 9580 2288
rect 9620 2248 9621 2288
rect 9579 2239 9621 2248
rect 9868 2120 9908 3331
rect 10156 2708 10196 2717
rect 10156 2549 10196 2668
rect 10155 2540 10197 2549
rect 10155 2500 10156 2540
rect 10196 2500 10197 2540
rect 10155 2491 10197 2500
rect 9868 2071 9908 2080
rect 9964 2456 10004 2465
rect 9676 1938 9716 1947
rect 9676 1364 9716 1898
rect 9867 1700 9909 1709
rect 9867 1660 9868 1700
rect 9908 1660 9909 1700
rect 9867 1651 9909 1660
rect 9676 1315 9716 1324
rect 9483 1280 9525 1289
rect 9483 1240 9484 1280
rect 9524 1240 9525 1280
rect 9483 1231 9525 1240
rect 9387 1112 9429 1121
rect 9387 1072 9388 1112
rect 9428 1072 9429 1112
rect 9387 1063 9429 1072
rect 9484 1112 9524 1231
rect 9388 524 9428 1063
rect 9484 701 9524 1072
rect 9483 692 9525 701
rect 9483 652 9484 692
rect 9524 652 9525 692
rect 9483 643 9525 652
rect 9388 484 9524 524
rect 9484 80 9524 484
rect 9675 440 9717 449
rect 9675 400 9676 440
rect 9716 400 9717 440
rect 9675 391 9717 400
rect 9676 80 9716 391
rect 9868 80 9908 1651
rect 9964 1028 10004 2416
rect 10155 2288 10197 2297
rect 10155 2248 10156 2288
rect 10196 2248 10197 2288
rect 10155 2239 10197 2248
rect 10059 1868 10101 1877
rect 10059 1828 10060 1868
rect 10100 1828 10101 1868
rect 10059 1819 10101 1828
rect 10060 1734 10100 1819
rect 10059 1616 10101 1625
rect 10059 1576 10060 1616
rect 10100 1576 10101 1616
rect 10059 1567 10101 1576
rect 10060 1196 10100 1567
rect 10060 1147 10100 1156
rect 9964 988 10100 1028
rect 10060 80 10100 988
rect 10156 533 10196 2239
rect 10252 1961 10292 4096
rect 10348 2456 10388 2465
rect 10251 1952 10293 1961
rect 10251 1912 10252 1952
rect 10292 1912 10293 1952
rect 10251 1903 10293 1912
rect 10252 1700 10292 1709
rect 10252 1121 10292 1660
rect 10251 1112 10293 1121
rect 10251 1072 10252 1112
rect 10292 1072 10293 1112
rect 10251 1063 10293 1072
rect 10252 944 10292 953
rect 10155 524 10197 533
rect 10155 484 10156 524
rect 10196 484 10197 524
rect 10155 475 10197 484
rect 10252 80 10292 904
rect 10348 365 10388 2416
rect 10443 1868 10485 1877
rect 10443 1828 10444 1868
rect 10484 1828 10485 1868
rect 10443 1819 10485 1828
rect 10444 1734 10484 1819
rect 10444 1196 10484 1205
rect 10540 1196 10580 9295
rect 10636 8597 10676 9472
rect 10635 8588 10677 8597
rect 10635 8548 10636 8588
rect 10676 8548 10677 8588
rect 10635 8539 10677 8548
rect 10636 8000 10676 8539
rect 10636 7951 10676 7960
rect 10732 7748 10772 11320
rect 10828 11024 10868 11035
rect 10828 10949 10868 10984
rect 10827 10940 10869 10949
rect 10827 10900 10828 10940
rect 10868 10900 10869 10940
rect 10827 10891 10869 10900
rect 10828 8513 10868 10891
rect 10827 8504 10869 8513
rect 10827 8464 10828 8504
rect 10868 8464 10869 8504
rect 10827 8455 10869 8464
rect 10827 8084 10869 8093
rect 10827 8044 10828 8084
rect 10868 8044 10869 8084
rect 10827 8035 10869 8044
rect 10828 7950 10868 8035
rect 10636 7708 10772 7748
rect 10636 4220 10676 7708
rect 10731 5144 10773 5153
rect 10731 5104 10732 5144
rect 10772 5104 10773 5144
rect 10731 5095 10773 5104
rect 10636 4171 10676 4180
rect 10732 4220 10772 5095
rect 10732 4171 10772 4180
rect 10924 3968 10964 11563
rect 11020 11192 11060 12486
rect 11020 11143 11060 11152
rect 11019 10604 11061 10613
rect 11019 10564 11020 10604
rect 11060 10564 11061 10604
rect 11019 10555 11061 10564
rect 11020 9680 11060 10555
rect 11116 10016 11156 15847
rect 11212 15728 11252 16192
rect 11500 16192 11636 16232
rect 11308 16148 11348 16157
rect 11500 16148 11540 16192
rect 11348 16108 11540 16148
rect 11308 16099 11348 16108
rect 11212 15679 11252 15688
rect 11404 15476 11444 16108
rect 11595 15644 11637 15653
rect 11595 15604 11596 15644
rect 11636 15604 11637 15644
rect 11595 15595 11637 15604
rect 11596 15560 11636 15595
rect 11596 15509 11636 15520
rect 11308 15436 11444 15476
rect 11308 15140 11348 15436
rect 11692 15392 11732 16771
rect 11788 15653 11828 16948
rect 11883 16232 11925 16241
rect 11883 16192 11884 16232
rect 11924 16192 11925 16232
rect 11883 16183 11925 16192
rect 11884 16098 11924 16183
rect 11787 15644 11829 15653
rect 11787 15604 11788 15644
rect 11828 15604 11829 15644
rect 11787 15595 11829 15604
rect 11692 15352 11924 15392
rect 11404 15308 11444 15317
rect 11444 15268 11732 15308
rect 11404 15259 11444 15268
rect 11308 15100 11540 15140
rect 11211 14720 11253 14729
rect 11211 14680 11212 14720
rect 11252 14680 11253 14720
rect 11211 14671 11253 14680
rect 11212 14048 11252 14671
rect 11212 13999 11252 14008
rect 11403 12452 11445 12461
rect 11403 12412 11404 12452
rect 11444 12412 11445 12452
rect 11403 12403 11445 12412
rect 11211 10856 11253 10865
rect 11211 10816 11212 10856
rect 11252 10816 11253 10856
rect 11211 10807 11253 10816
rect 11212 10184 11252 10807
rect 11212 10135 11252 10144
rect 11307 10184 11349 10193
rect 11307 10144 11308 10184
rect 11348 10144 11349 10184
rect 11307 10135 11349 10144
rect 11308 10050 11348 10135
rect 11116 9976 11252 10016
rect 11020 9640 11156 9680
rect 11020 9512 11060 9521
rect 11020 8924 11060 9472
rect 11116 9512 11156 9640
rect 11116 9463 11156 9472
rect 11212 9437 11252 9976
rect 11211 9428 11253 9437
rect 11211 9388 11212 9428
rect 11252 9388 11253 9428
rect 11211 9379 11253 9388
rect 11212 8924 11252 8933
rect 11020 8884 11212 8924
rect 11212 8875 11252 8884
rect 11020 8672 11060 8683
rect 11020 8597 11060 8632
rect 11019 8588 11061 8597
rect 11019 8548 11020 8588
rect 11060 8548 11061 8588
rect 11019 8539 11061 8548
rect 11115 8084 11157 8093
rect 11115 8044 11116 8084
rect 11156 8044 11157 8084
rect 11115 8035 11157 8044
rect 11116 8000 11156 8035
rect 11116 7949 11156 7960
rect 11212 8000 11252 8009
rect 11404 8000 11444 12403
rect 11500 10100 11540 15100
rect 11692 14734 11732 15268
rect 11692 14685 11732 14694
rect 11884 14636 11924 15352
rect 11596 14596 11884 14636
rect 11596 12704 11636 14596
rect 11884 14587 11924 14596
rect 11980 14384 12020 17032
rect 12076 17023 12116 17032
rect 12171 16652 12213 16661
rect 12171 16612 12172 16652
rect 12212 16612 12213 16652
rect 12171 16603 12213 16612
rect 12075 16484 12117 16493
rect 12075 16444 12076 16484
rect 12116 16444 12117 16484
rect 12075 16435 12117 16444
rect 12076 15737 12116 16435
rect 12075 15728 12117 15737
rect 12075 15688 12076 15728
rect 12116 15688 12117 15728
rect 12075 15679 12117 15688
rect 11788 14344 12020 14384
rect 11692 14057 11732 14138
rect 11691 14048 11733 14057
rect 11691 14003 11692 14048
rect 11732 14003 11733 14048
rect 11691 13999 11733 14003
rect 11692 13994 11732 13999
rect 11691 13796 11733 13805
rect 11691 13756 11692 13796
rect 11732 13756 11733 13796
rect 11691 13747 11733 13756
rect 11692 13460 11732 13747
rect 11788 13721 11828 14344
rect 11883 14216 11925 14225
rect 11883 14176 11884 14216
rect 11924 14176 11925 14216
rect 11883 14167 11925 14176
rect 11787 13712 11829 13721
rect 11787 13672 11788 13712
rect 11828 13672 11829 13712
rect 11787 13663 11829 13672
rect 11692 13420 11828 13460
rect 11596 12664 11732 12704
rect 11596 12536 11636 12545
rect 11596 12284 11636 12496
rect 11692 12461 11732 12664
rect 11788 12629 11828 13420
rect 11787 12620 11829 12629
rect 11787 12580 11788 12620
rect 11828 12580 11829 12620
rect 11787 12571 11829 12580
rect 11691 12452 11733 12461
rect 11691 12412 11692 12452
rect 11732 12412 11733 12452
rect 11691 12403 11733 12412
rect 11788 12284 11828 12571
rect 11596 12244 11828 12284
rect 11595 11696 11637 11705
rect 11595 11656 11596 11696
rect 11636 11656 11637 11696
rect 11595 11647 11637 11656
rect 11596 11562 11636 11647
rect 11884 11621 11924 14167
rect 12076 13208 12116 15679
rect 12172 14048 12212 16603
rect 12268 15821 12308 20719
rect 12363 19340 12405 19349
rect 12363 19300 12364 19340
rect 12404 19300 12405 19340
rect 12363 19291 12405 19300
rect 12364 19256 12404 19291
rect 12364 19205 12404 19216
rect 12363 18248 12405 18257
rect 12363 18208 12364 18248
rect 12404 18208 12405 18248
rect 12363 18199 12405 18208
rect 12364 16232 12404 18199
rect 12460 17921 12500 27355
rect 12556 26396 12596 27523
rect 12556 26356 12692 26396
rect 12556 26153 12596 26238
rect 12555 26144 12597 26153
rect 12555 26104 12556 26144
rect 12596 26104 12597 26144
rect 12555 26095 12597 26104
rect 12652 25976 12692 26356
rect 12556 25936 12692 25976
rect 12556 22793 12596 25936
rect 12652 24632 12692 24641
rect 12652 23969 12692 24592
rect 12651 23960 12693 23969
rect 12651 23920 12652 23960
rect 12692 23920 12693 23960
rect 12651 23911 12693 23920
rect 12652 23792 12692 23801
rect 12652 23549 12692 23752
rect 12748 23624 12788 28960
rect 12844 28673 12884 33319
rect 12940 32696 12980 34168
rect 13131 34124 13173 34133
rect 13131 34084 13132 34124
rect 13172 34084 13173 34124
rect 13131 34075 13173 34084
rect 13035 33956 13077 33965
rect 13035 33916 13036 33956
rect 13076 33916 13077 33956
rect 13035 33907 13077 33916
rect 13036 32864 13076 33907
rect 13132 33536 13172 34075
rect 13228 33788 13268 35092
rect 13420 34544 13460 37771
rect 13516 34553 13556 40123
rect 13612 38912 13652 40879
rect 13803 40676 13845 40685
rect 13803 40636 13804 40676
rect 13844 40636 13845 40676
rect 13803 40627 13845 40636
rect 13804 40433 13844 40627
rect 13803 40424 13845 40433
rect 13803 40384 13804 40424
rect 13844 40384 13845 40424
rect 13803 40375 13845 40384
rect 13804 40290 13844 40375
rect 13996 40256 14036 40265
rect 13803 39668 13845 39677
rect 13803 39628 13804 39668
rect 13844 39628 13845 39668
rect 13803 39619 13845 39628
rect 13900 39668 13940 39677
rect 13804 39534 13844 39619
rect 13900 39416 13940 39628
rect 13804 39376 13940 39416
rect 13804 39089 13844 39376
rect 13899 39248 13941 39257
rect 13899 39208 13900 39248
rect 13940 39208 13941 39248
rect 13899 39199 13941 39208
rect 13803 39080 13845 39089
rect 13803 39040 13804 39080
rect 13844 39040 13845 39080
rect 13803 39031 13845 39040
rect 13612 38872 13844 38912
rect 13611 38156 13653 38165
rect 13611 38116 13612 38156
rect 13652 38116 13653 38156
rect 13611 38107 13653 38116
rect 13324 34504 13460 34544
rect 13515 34544 13557 34553
rect 13515 34504 13516 34544
rect 13556 34504 13557 34544
rect 13324 33965 13364 34504
rect 13515 34495 13557 34504
rect 13420 34376 13460 34385
rect 13420 34217 13460 34336
rect 13516 34376 13556 34387
rect 13516 34301 13556 34336
rect 13515 34292 13557 34301
rect 13515 34252 13516 34292
rect 13556 34252 13557 34292
rect 13515 34243 13557 34252
rect 13419 34208 13461 34217
rect 13419 34168 13420 34208
rect 13460 34168 13461 34208
rect 13419 34159 13461 34168
rect 13612 34040 13652 38107
rect 13707 35216 13749 35225
rect 13707 35176 13708 35216
rect 13748 35176 13749 35216
rect 13707 35167 13749 35176
rect 13708 35082 13748 35167
rect 13804 34796 13844 38872
rect 13900 37409 13940 39199
rect 13996 38912 14036 40216
rect 14092 39341 14132 41140
rect 14612 41140 14900 41180
rect 14956 41180 14996 41189
rect 15052 41180 15092 42928
rect 14996 41140 15092 41180
rect 14572 41131 14612 41140
rect 14956 41131 14996 41140
rect 14380 41012 14420 41021
rect 14380 40685 14420 40972
rect 14763 41012 14805 41021
rect 14763 40972 14764 41012
rect 14804 40972 14805 41012
rect 14763 40963 14805 40972
rect 15147 41012 15189 41021
rect 15147 40972 15148 41012
rect 15188 40972 15189 41012
rect 15147 40963 15189 40972
rect 14764 40878 14804 40963
rect 15148 40878 15188 40963
rect 14379 40676 14421 40685
rect 14379 40636 14380 40676
rect 14420 40636 14421 40676
rect 14379 40627 14421 40636
rect 14380 40433 14420 40518
rect 15244 40517 15284 42928
rect 15340 41180 15380 41189
rect 15436 41180 15476 42928
rect 15628 41432 15668 42928
rect 15820 41684 15860 42928
rect 16012 41768 16052 42928
rect 16012 41728 16148 41768
rect 15820 41644 16052 41684
rect 15724 41432 15764 41441
rect 15628 41392 15724 41432
rect 15724 41383 15764 41392
rect 15380 41140 15476 41180
rect 15916 41180 15956 41189
rect 15340 41131 15380 41140
rect 15819 40592 15861 40601
rect 15819 40552 15820 40592
rect 15860 40552 15861 40592
rect 15819 40543 15861 40552
rect 15243 40508 15285 40517
rect 15243 40468 15244 40508
rect 15284 40468 15285 40508
rect 15243 40459 15285 40468
rect 15820 40458 15860 40543
rect 14379 40424 14421 40433
rect 14284 40384 14380 40424
rect 14420 40384 14421 40424
rect 14187 40256 14229 40265
rect 14187 40216 14188 40256
rect 14228 40216 14229 40256
rect 14187 40207 14229 40216
rect 14188 40122 14228 40207
rect 14091 39332 14133 39341
rect 14091 39292 14092 39332
rect 14132 39292 14133 39332
rect 14091 39283 14133 39292
rect 14187 39248 14229 39257
rect 14187 39208 14188 39248
rect 14228 39208 14229 39248
rect 14187 39199 14229 39208
rect 14092 38912 14132 38921
rect 13996 38872 14092 38912
rect 14092 38863 14132 38872
rect 14188 38912 14228 39199
rect 14188 38863 14228 38872
rect 14092 38240 14132 38249
rect 14284 38240 14324 40384
rect 14379 40375 14421 40384
rect 15627 40424 15669 40433
rect 15627 40384 15628 40424
rect 15668 40384 15669 40424
rect 15627 40375 15669 40384
rect 15435 40340 15477 40349
rect 15435 40300 15436 40340
rect 15476 40300 15477 40340
rect 15435 40291 15477 40300
rect 14859 40256 14901 40265
rect 14859 40216 14860 40256
rect 14900 40216 14901 40256
rect 14859 40207 14901 40216
rect 14379 40088 14421 40097
rect 14379 40048 14380 40088
rect 14420 40048 14421 40088
rect 14379 40039 14421 40048
rect 14380 39752 14420 40039
rect 14420 39712 14516 39752
rect 14380 39703 14420 39712
rect 14379 39332 14421 39341
rect 14379 39292 14380 39332
rect 14420 39292 14421 39332
rect 14379 39283 14421 39292
rect 14132 38200 14324 38240
rect 14092 38072 14132 38200
rect 13996 38032 14132 38072
rect 13899 37400 13941 37409
rect 13899 37360 13900 37400
rect 13940 37360 13941 37400
rect 13899 37351 13941 37360
rect 13420 34000 13652 34040
rect 13708 34756 13844 34796
rect 13323 33956 13365 33965
rect 13323 33916 13324 33956
rect 13364 33916 13365 33956
rect 13323 33907 13365 33916
rect 13420 33914 13460 34000
rect 13420 33865 13460 33874
rect 13228 33748 13364 33788
rect 13324 33704 13364 33748
rect 13612 33704 13652 33713
rect 13228 33690 13268 33699
rect 13324 33664 13460 33704
rect 13228 33620 13268 33650
rect 13228 33580 13364 33620
rect 13132 33496 13268 33536
rect 13132 32873 13172 32958
rect 13131 32864 13173 32873
rect 13036 32824 13132 32864
rect 13172 32824 13173 32864
rect 13131 32815 13173 32824
rect 12940 32656 13172 32696
rect 13035 32528 13077 32537
rect 13035 32488 13036 32528
rect 13076 32488 13077 32528
rect 13035 32479 13077 32488
rect 12939 32192 12981 32201
rect 12939 32152 12940 32192
rect 12980 32152 12981 32192
rect 12939 32143 12981 32152
rect 12940 30605 12980 32143
rect 12939 30596 12981 30605
rect 12939 30556 12940 30596
rect 12980 30556 12981 30596
rect 12939 30547 12981 30556
rect 12939 30428 12981 30437
rect 12939 30388 12940 30428
rect 12980 30388 12981 30428
rect 12939 30379 12981 30388
rect 12843 28664 12885 28673
rect 12843 28624 12844 28664
rect 12884 28624 12885 28664
rect 12843 28615 12885 28624
rect 12844 28328 12884 28337
rect 12940 28328 12980 30379
rect 13036 29420 13076 32479
rect 13132 29681 13172 32656
rect 13131 29672 13173 29681
rect 13131 29632 13132 29672
rect 13172 29632 13173 29672
rect 13131 29623 13173 29632
rect 13228 29504 13268 33496
rect 13324 33116 13364 33580
rect 13324 33067 13364 33076
rect 13323 32864 13365 32873
rect 13323 32824 13324 32864
rect 13364 32824 13365 32864
rect 13323 32815 13365 32824
rect 13324 31277 13364 32815
rect 13323 31268 13365 31277
rect 13323 31228 13324 31268
rect 13364 31228 13365 31268
rect 13323 31219 13365 31228
rect 13324 30941 13364 31219
rect 13323 30932 13365 30941
rect 13323 30892 13324 30932
rect 13364 30892 13365 30932
rect 13323 30883 13365 30892
rect 13324 29840 13364 30883
rect 13420 30773 13460 33664
rect 13515 31688 13557 31697
rect 13515 31648 13516 31688
rect 13556 31648 13557 31688
rect 13515 31639 13557 31648
rect 13419 30764 13461 30773
rect 13419 30724 13420 30764
rect 13460 30724 13461 30764
rect 13419 30715 13461 30724
rect 13324 29791 13364 29800
rect 13420 29588 13460 30715
rect 13516 30269 13556 31639
rect 13515 30260 13557 30269
rect 13515 30220 13516 30260
rect 13556 30220 13557 30260
rect 13515 30211 13557 30220
rect 13612 30101 13652 33664
rect 13708 32201 13748 34756
rect 13996 34712 14036 38032
rect 14284 37988 14324 37997
rect 14092 37948 14284 37988
rect 14092 37400 14132 37948
rect 14284 37939 14324 37948
rect 14283 37736 14325 37745
rect 14283 37696 14284 37736
rect 14324 37696 14325 37736
rect 14283 37687 14325 37696
rect 14092 37351 14132 37360
rect 14187 37400 14229 37409
rect 14187 37360 14188 37400
rect 14228 37360 14229 37400
rect 14187 37351 14229 37360
rect 13804 34672 14036 34712
rect 13804 34385 13844 34672
rect 13900 34469 13940 34500
rect 13899 34460 13941 34469
rect 13899 34420 13900 34460
rect 13940 34420 13941 34460
rect 13899 34411 13941 34420
rect 13803 34376 13845 34385
rect 13803 34336 13804 34376
rect 13844 34336 13845 34376
rect 13803 34327 13845 34336
rect 13900 34376 13940 34411
rect 13803 33788 13845 33797
rect 13803 33748 13804 33788
rect 13844 33748 13845 33788
rect 13803 33739 13845 33748
rect 13804 32789 13844 33739
rect 13803 32780 13845 32789
rect 13803 32740 13804 32780
rect 13844 32740 13845 32780
rect 13803 32731 13845 32740
rect 13707 32192 13749 32201
rect 13707 32152 13708 32192
rect 13748 32152 13749 32192
rect 13707 32143 13749 32152
rect 13900 32024 13940 34336
rect 13995 34376 14037 34385
rect 13995 34336 13996 34376
rect 14036 34336 14037 34376
rect 13995 34327 14037 34336
rect 13996 34242 14036 34327
rect 14188 34301 14228 37351
rect 14187 34292 14229 34301
rect 14187 34252 14188 34292
rect 14228 34252 14229 34292
rect 14187 34243 14229 34252
rect 14284 34049 14324 37687
rect 14380 34805 14420 39283
rect 14476 38921 14516 39712
rect 14860 39747 14900 40207
rect 14860 39698 14900 39707
rect 15052 39836 15092 39845
rect 14571 39668 14613 39677
rect 14571 39628 14572 39668
rect 14612 39628 14613 39668
rect 14571 39619 14613 39628
rect 14572 38996 14612 39619
rect 14667 39080 14709 39089
rect 14667 39040 14668 39080
rect 14708 39040 14709 39080
rect 14667 39031 14709 39040
rect 14475 38912 14517 38921
rect 14475 38872 14476 38912
rect 14516 38872 14517 38912
rect 14475 38863 14517 38872
rect 14476 38240 14516 38249
rect 14476 37997 14516 38200
rect 14475 37988 14517 37997
rect 14475 37948 14476 37988
rect 14516 37948 14517 37988
rect 14475 37939 14517 37948
rect 14475 37820 14517 37829
rect 14475 37780 14476 37820
rect 14516 37780 14517 37820
rect 14475 37771 14517 37780
rect 14379 34796 14421 34805
rect 14379 34756 14380 34796
rect 14420 34756 14421 34796
rect 14379 34747 14421 34756
rect 14476 34376 14516 37771
rect 14572 37400 14612 38956
rect 14572 34469 14612 37360
rect 14668 38996 14708 39031
rect 14668 37400 14708 38956
rect 15052 37829 15092 39796
rect 15436 39752 15476 40291
rect 15628 40290 15668 40375
rect 15476 39712 15764 39752
rect 15436 39703 15476 39712
rect 15244 39500 15284 39509
rect 15284 39460 15668 39500
rect 15244 39451 15284 39460
rect 15339 39332 15381 39341
rect 15339 39292 15340 39332
rect 15380 39292 15381 39332
rect 15339 39283 15381 39292
rect 15147 38912 15189 38921
rect 15147 38872 15148 38912
rect 15188 38872 15189 38912
rect 15147 38863 15189 38872
rect 15148 37913 15188 38863
rect 15147 37904 15189 37913
rect 15147 37864 15148 37904
rect 15188 37864 15189 37904
rect 15147 37855 15189 37864
rect 15051 37820 15093 37829
rect 15051 37780 15052 37820
rect 15092 37780 15093 37820
rect 15051 37771 15093 37780
rect 14571 34460 14613 34469
rect 14571 34420 14572 34460
rect 14612 34420 14613 34460
rect 14571 34411 14613 34420
rect 14668 34385 14708 37360
rect 15148 37400 15188 37855
rect 15148 37351 15188 37360
rect 14955 36980 14997 36989
rect 14955 36940 14956 36980
rect 14996 36940 14997 36980
rect 14955 36931 14997 36940
rect 14956 35561 14996 36931
rect 15147 36812 15189 36821
rect 15147 36772 15148 36812
rect 15188 36772 15189 36812
rect 15147 36763 15189 36772
rect 15148 36728 15188 36763
rect 15148 36677 15188 36688
rect 15340 36065 15380 39283
rect 15628 38926 15668 39460
rect 15628 38877 15668 38886
rect 15627 38492 15669 38501
rect 15627 38452 15628 38492
rect 15668 38452 15669 38492
rect 15627 38443 15669 38452
rect 15531 38240 15573 38249
rect 15531 38200 15532 38240
rect 15572 38200 15573 38240
rect 15531 38191 15573 38200
rect 15339 36056 15381 36065
rect 15339 36016 15340 36056
rect 15380 36016 15381 36056
rect 15339 36007 15381 36016
rect 15340 35888 15380 35897
rect 14955 35552 14997 35561
rect 14955 35512 14956 35552
rect 14996 35512 14997 35552
rect 14955 35503 14997 35512
rect 14956 35216 14996 35503
rect 15148 35384 15188 35393
rect 15340 35384 15380 35848
rect 15436 35888 15476 35897
rect 15436 35813 15476 35848
rect 15435 35804 15477 35813
rect 15435 35764 15436 35804
rect 15476 35764 15477 35804
rect 15435 35755 15477 35764
rect 15436 35477 15476 35755
rect 15435 35468 15477 35477
rect 15435 35428 15436 35468
rect 15476 35428 15477 35468
rect 15435 35419 15477 35428
rect 15188 35344 15380 35384
rect 15148 35335 15188 35344
rect 15340 35216 15380 35344
rect 15436 35216 15476 35225
rect 15340 35176 15436 35216
rect 14956 35141 14996 35176
rect 15436 35167 15476 35176
rect 15532 35216 15572 38191
rect 15628 37913 15668 38443
rect 15724 38240 15764 39712
rect 15820 38744 15860 38753
rect 15916 38744 15956 41140
rect 16012 40676 16052 41644
rect 16108 41609 16148 41728
rect 16107 41600 16149 41609
rect 16107 41560 16108 41600
rect 16148 41560 16149 41600
rect 16107 41551 16149 41560
rect 16108 41432 16148 41441
rect 16204 41432 16244 42928
rect 16148 41392 16244 41432
rect 16108 41383 16148 41392
rect 16300 41180 16340 41189
rect 16204 40676 16244 40685
rect 16012 40636 16204 40676
rect 16204 40627 16244 40636
rect 16011 40508 16053 40517
rect 16011 40468 16012 40508
rect 16052 40468 16053 40508
rect 16011 40459 16053 40468
rect 16012 40374 16052 40459
rect 16107 40424 16149 40433
rect 16107 40384 16108 40424
rect 16148 40384 16149 40424
rect 16107 40375 16149 40384
rect 16011 39752 16053 39761
rect 16011 39712 16012 39752
rect 16052 39712 16053 39752
rect 16011 39703 16053 39712
rect 16012 38912 16052 39703
rect 16012 38863 16052 38872
rect 15916 38704 16052 38744
rect 15820 38249 15860 38704
rect 15724 38191 15764 38200
rect 15819 38240 15861 38249
rect 15819 38200 15820 38240
rect 15860 38200 15861 38240
rect 15819 38191 15861 38200
rect 15916 37988 15956 37997
rect 15627 37904 15669 37913
rect 15627 37864 15628 37904
rect 15668 37864 15669 37904
rect 15627 37855 15669 37864
rect 15916 37820 15956 37948
rect 15724 37780 15956 37820
rect 15724 37484 15764 37780
rect 16012 37661 16052 38704
rect 16108 38156 16148 40375
rect 16300 39920 16340 41140
rect 16396 40685 16436 42928
rect 16588 41609 16628 42928
rect 16587 41600 16629 41609
rect 16587 41560 16588 41600
rect 16628 41560 16629 41600
rect 16587 41551 16629 41560
rect 16491 41516 16533 41525
rect 16491 41476 16492 41516
rect 16532 41476 16533 41516
rect 16491 41467 16533 41476
rect 16395 40676 16437 40685
rect 16395 40636 16396 40676
rect 16436 40636 16437 40676
rect 16492 40676 16532 41467
rect 16780 41264 16820 42928
rect 16972 41432 17012 42928
rect 17164 41693 17204 42928
rect 17163 41684 17205 41693
rect 17163 41644 17164 41684
rect 17204 41644 17205 41684
rect 17163 41635 17205 41644
rect 17356 41609 17396 42928
rect 17355 41600 17397 41609
rect 17355 41560 17356 41600
rect 17396 41560 17397 41600
rect 17355 41551 17397 41560
rect 17260 41432 17300 41441
rect 16972 41392 17260 41432
rect 17260 41383 17300 41392
rect 16684 41224 16820 41264
rect 16587 41180 16629 41189
rect 16587 41140 16588 41180
rect 16628 41140 16629 41180
rect 16587 41131 16629 41140
rect 16588 41046 16628 41131
rect 16588 40676 16628 40685
rect 16492 40636 16588 40676
rect 16395 40627 16437 40636
rect 16588 40627 16628 40636
rect 16396 40508 16436 40517
rect 16396 40181 16436 40468
rect 16684 40349 16724 41224
rect 16972 41180 17012 41189
rect 17452 41180 17492 41189
rect 16876 41140 16972 41180
rect 16779 41096 16821 41105
rect 16779 41056 16780 41096
rect 16820 41056 16821 41096
rect 16779 41047 16821 41056
rect 16780 40962 16820 41047
rect 16780 40508 16820 40519
rect 16780 40433 16820 40468
rect 16779 40424 16821 40433
rect 16779 40384 16780 40424
rect 16820 40384 16821 40424
rect 16779 40375 16821 40384
rect 16683 40340 16725 40349
rect 16683 40300 16684 40340
rect 16724 40300 16725 40340
rect 16683 40291 16725 40300
rect 16395 40172 16437 40181
rect 16395 40132 16396 40172
rect 16436 40132 16437 40172
rect 16395 40123 16437 40132
rect 16204 39880 16340 39920
rect 16204 39341 16244 39880
rect 16299 39752 16341 39761
rect 16299 39712 16300 39752
rect 16340 39712 16341 39752
rect 16299 39703 16341 39712
rect 16684 39752 16724 39761
rect 16203 39332 16245 39341
rect 16203 39292 16204 39332
rect 16244 39292 16245 39332
rect 16203 39283 16245 39292
rect 16203 39164 16245 39173
rect 16203 39124 16204 39164
rect 16244 39124 16245 39164
rect 16203 39115 16245 39124
rect 16204 38408 16244 39115
rect 16300 39080 16340 39703
rect 16300 39031 16340 39040
rect 16395 39080 16437 39089
rect 16395 39040 16396 39080
rect 16436 39040 16437 39080
rect 16395 39031 16437 39040
rect 16300 38912 16340 38921
rect 16396 38912 16436 39031
rect 16340 38872 16436 38912
rect 16492 38912 16532 38921
rect 16300 38863 16340 38872
rect 16300 38408 16340 38417
rect 16204 38368 16300 38408
rect 16300 38359 16340 38368
rect 16108 38107 16148 38116
rect 16203 37904 16245 37913
rect 16203 37864 16204 37904
rect 16244 37864 16245 37904
rect 16203 37855 16245 37864
rect 16011 37652 16053 37661
rect 16011 37612 16012 37652
rect 16052 37612 16053 37652
rect 16011 37603 16053 37612
rect 15676 37444 15764 37484
rect 15676 37442 15716 37444
rect 15676 37393 15716 37402
rect 16204 37400 16244 37855
rect 16395 37568 16437 37577
rect 16395 37528 16396 37568
rect 16436 37528 16437 37568
rect 16395 37519 16437 37528
rect 16107 37316 16149 37325
rect 16107 37276 16108 37316
rect 16148 37276 16149 37316
rect 16107 37267 16149 37276
rect 15819 37232 15861 37241
rect 15819 37192 15820 37232
rect 15860 37192 15861 37232
rect 15819 37183 15861 37192
rect 15820 36569 15860 37183
rect 16011 36644 16053 36653
rect 16011 36604 16012 36644
rect 16052 36604 16053 36644
rect 16011 36595 16053 36604
rect 15819 36560 15861 36569
rect 15819 36520 15820 36560
rect 15860 36520 15861 36560
rect 15819 36511 15861 36520
rect 15820 35888 15860 35897
rect 15820 35645 15860 35848
rect 15915 35888 15957 35897
rect 15915 35848 15916 35888
rect 15956 35848 15957 35888
rect 15915 35839 15957 35848
rect 15916 35754 15956 35839
rect 15819 35636 15861 35645
rect 15819 35596 15820 35636
rect 15860 35596 15861 35636
rect 15819 35587 15861 35596
rect 15819 35468 15861 35477
rect 15819 35428 15820 35468
rect 15860 35428 15861 35468
rect 15819 35419 15861 35428
rect 15572 35176 15668 35216
rect 15532 35167 15572 35176
rect 14955 35132 14997 35141
rect 14955 35092 14956 35132
rect 14996 35092 14997 35132
rect 14955 35083 14997 35092
rect 14956 35052 14996 35083
rect 14859 34796 14901 34805
rect 14859 34756 14860 34796
rect 14900 34756 14901 34796
rect 14859 34747 14901 34756
rect 14763 34544 14805 34553
rect 14763 34504 14764 34544
rect 14804 34504 14805 34544
rect 14763 34495 14805 34504
rect 14476 34133 14516 34336
rect 14667 34376 14709 34385
rect 14667 34336 14668 34376
rect 14708 34336 14709 34376
rect 14667 34327 14709 34336
rect 14475 34124 14517 34133
rect 14475 34084 14476 34124
rect 14516 34084 14517 34124
rect 14475 34075 14517 34084
rect 14283 34040 14325 34049
rect 14283 34000 14284 34040
rect 14324 34000 14325 34040
rect 14283 33991 14325 34000
rect 14091 33368 14133 33377
rect 14091 33328 14092 33368
rect 14132 33328 14133 33368
rect 14091 33319 14133 33328
rect 14092 32957 14132 33319
rect 14091 32948 14133 32957
rect 14091 32908 14092 32948
rect 14132 32908 14133 32948
rect 14091 32899 14133 32908
rect 14092 32864 14132 32899
rect 14092 32814 14132 32824
rect 13708 31984 13940 32024
rect 14188 32192 14228 32201
rect 13611 30092 13653 30101
rect 13611 30052 13612 30092
rect 13652 30052 13653 30092
rect 13611 30043 13653 30052
rect 13515 30008 13557 30017
rect 13515 29968 13516 30008
rect 13556 29968 13557 30008
rect 13515 29959 13557 29968
rect 13516 29874 13556 29959
rect 13708 29924 13748 31984
rect 14188 31949 14228 32152
rect 13995 31940 14037 31949
rect 13995 31900 13996 31940
rect 14036 31900 14037 31940
rect 13995 31891 14037 31900
rect 14187 31940 14229 31949
rect 14187 31900 14188 31940
rect 14228 31900 14229 31940
rect 14187 31891 14229 31900
rect 13996 31352 14036 31891
rect 14284 31781 14324 33991
rect 14571 32192 14613 32201
rect 14571 32152 14572 32192
rect 14612 32152 14613 32192
rect 14571 32143 14613 32152
rect 14572 32058 14612 32143
rect 14668 32117 14708 34327
rect 14764 33704 14804 34495
rect 14860 34292 14900 34747
rect 15243 34712 15285 34721
rect 15243 34672 15244 34712
rect 15284 34672 15285 34712
rect 15243 34663 15285 34672
rect 15004 34385 15044 34394
rect 15044 34345 15092 34376
rect 15004 34336 15092 34345
rect 14860 34252 14996 34292
rect 14860 33704 14900 33713
rect 14764 33664 14860 33704
rect 14667 32108 14709 32117
rect 14667 32068 14668 32108
rect 14708 32068 14709 32108
rect 14667 32059 14709 32068
rect 14860 31949 14900 33664
rect 14380 31940 14420 31949
rect 14668 31940 14708 31949
rect 14859 31940 14901 31949
rect 14420 31900 14612 31940
rect 14380 31891 14420 31900
rect 14283 31772 14325 31781
rect 14283 31732 14284 31772
rect 14324 31732 14325 31772
rect 14283 31723 14325 31732
rect 13996 30857 14036 31312
rect 14188 31520 14228 31529
rect 14228 31480 14516 31520
rect 13995 30848 14037 30857
rect 13995 30808 13996 30848
rect 14036 30808 14037 30848
rect 13995 30799 14037 30808
rect 13995 30680 14037 30689
rect 13995 30640 13996 30680
rect 14036 30640 14037 30680
rect 13995 30631 14037 30640
rect 14188 30680 14228 31480
rect 14476 31361 14516 31480
rect 14572 31361 14612 31900
rect 14708 31900 14804 31940
rect 14668 31891 14708 31900
rect 14667 31520 14709 31529
rect 14667 31480 14668 31520
rect 14708 31480 14709 31520
rect 14667 31471 14709 31480
rect 14283 31352 14325 31361
rect 14283 31312 14284 31352
rect 14324 31312 14325 31352
rect 14283 31303 14325 31312
rect 14380 31352 14420 31361
rect 14188 30631 14228 30640
rect 14284 30680 14324 31303
rect 14284 30631 14324 30640
rect 13996 30546 14036 30631
rect 14187 30512 14229 30521
rect 14187 30472 14188 30512
rect 14228 30472 14229 30512
rect 14187 30463 14229 30472
rect 14284 30512 14324 30521
rect 14380 30512 14420 31312
rect 14476 31352 14518 31361
rect 14516 31312 14518 31352
rect 14476 31308 14518 31312
rect 14571 31352 14613 31361
rect 14571 31312 14572 31352
rect 14612 31312 14613 31352
rect 14476 31303 14516 31308
rect 14571 31303 14613 31312
rect 14668 31352 14708 31471
rect 14668 31303 14708 31312
rect 14764 31352 14804 31900
rect 14859 31900 14860 31940
rect 14900 31900 14901 31940
rect 14859 31891 14901 31900
rect 14865 31361 14905 31446
rect 14764 31303 14804 31312
rect 14864 31352 14906 31361
rect 14864 31312 14865 31352
rect 14905 31312 14906 31352
rect 14864 31303 14906 31312
rect 14763 31184 14805 31193
rect 14763 31144 14764 31184
rect 14804 31144 14805 31184
rect 14763 31135 14805 31144
rect 14860 31184 14900 31193
rect 14667 31100 14709 31109
rect 14667 31060 14668 31100
rect 14708 31060 14709 31100
rect 14667 31051 14709 31060
rect 14475 30680 14517 30689
rect 14475 30640 14476 30680
rect 14516 30640 14517 30680
rect 14475 30631 14517 30640
rect 14324 30472 14420 30512
rect 14284 30463 14324 30472
rect 13803 30008 13845 30017
rect 13803 29968 13804 30008
rect 13844 29968 13845 30008
rect 13803 29959 13845 29968
rect 13612 29884 13748 29924
rect 13420 29548 13556 29588
rect 13228 29464 13460 29504
rect 13036 29380 13364 29420
rect 13131 28916 13173 28925
rect 13131 28876 13132 28916
rect 13172 28876 13173 28916
rect 13131 28867 13173 28876
rect 12884 28288 12980 28328
rect 13036 28328 13076 28337
rect 12844 28279 12884 28288
rect 12939 28160 12981 28169
rect 12939 28120 12940 28160
rect 12980 28120 12981 28160
rect 12939 28111 12981 28120
rect 12940 28026 12980 28111
rect 12843 27824 12885 27833
rect 12843 27784 12844 27824
rect 12884 27784 12885 27824
rect 12843 27775 12885 27784
rect 12844 26153 12884 27775
rect 13036 27749 13076 28288
rect 13132 28328 13172 28867
rect 13227 28664 13269 28673
rect 13227 28624 13228 28664
rect 13268 28624 13269 28664
rect 13227 28615 13269 28624
rect 13132 28279 13172 28288
rect 13035 27740 13077 27749
rect 13035 27700 13036 27740
rect 13076 27700 13077 27740
rect 13035 27691 13077 27700
rect 13035 26228 13077 26237
rect 13035 26188 13036 26228
rect 13076 26188 13077 26228
rect 13035 26179 13077 26188
rect 12843 26144 12885 26153
rect 12843 26104 12844 26144
rect 12884 26104 12885 26144
rect 12843 26095 12885 26104
rect 12844 25733 12884 26095
rect 12843 25724 12885 25733
rect 12843 25684 12844 25724
rect 12884 25684 12885 25724
rect 12843 25675 12885 25684
rect 12844 23960 12884 23971
rect 12844 23885 12884 23920
rect 12843 23876 12885 23885
rect 12843 23836 12844 23876
rect 12884 23836 12885 23876
rect 12843 23827 12885 23836
rect 12748 23584 12980 23624
rect 12651 23540 12693 23549
rect 12651 23500 12652 23540
rect 12692 23500 12693 23540
rect 12651 23491 12693 23500
rect 12555 22784 12597 22793
rect 12555 22744 12556 22784
rect 12596 22744 12597 22784
rect 12555 22735 12597 22744
rect 12555 22448 12597 22457
rect 12555 22408 12556 22448
rect 12596 22408 12597 22448
rect 12555 22399 12597 22408
rect 12556 21869 12596 22399
rect 12555 21860 12597 21869
rect 12555 21820 12556 21860
rect 12596 21820 12597 21860
rect 12555 21811 12597 21820
rect 12747 21692 12789 21701
rect 12747 21652 12748 21692
rect 12788 21652 12789 21692
rect 12747 21643 12789 21652
rect 12604 21566 12644 21575
rect 12748 21558 12788 21643
rect 12940 21608 12980 23584
rect 12844 21568 12940 21608
rect 12604 21524 12644 21526
rect 12604 21484 12692 21524
rect 12652 21020 12692 21484
rect 12748 21020 12788 21029
rect 12652 20980 12748 21020
rect 12748 20971 12788 20980
rect 12555 20768 12597 20777
rect 12555 20728 12556 20768
rect 12596 20728 12597 20768
rect 12555 20719 12597 20728
rect 12556 20634 12596 20719
rect 12748 20180 12788 20220
rect 12748 20105 12788 20140
rect 12747 20096 12789 20105
rect 12556 20082 12596 20091
rect 12747 20056 12748 20096
rect 12788 20056 12789 20096
rect 12747 20047 12789 20056
rect 12748 20045 12788 20047
rect 12556 19508 12596 20042
rect 12556 19459 12596 19468
rect 12844 18752 12884 21568
rect 12940 21559 12980 21568
rect 12939 20684 12981 20693
rect 12939 20644 12940 20684
rect 12980 20644 12981 20684
rect 12939 20635 12981 20644
rect 12748 18712 12884 18752
rect 12940 20096 12980 20635
rect 12651 18500 12693 18509
rect 12651 18460 12652 18500
rect 12692 18460 12693 18500
rect 12651 18451 12693 18460
rect 12652 18089 12692 18451
rect 12651 18080 12693 18089
rect 12651 18040 12652 18080
rect 12692 18040 12693 18080
rect 12651 18031 12693 18040
rect 12748 17921 12788 18712
rect 12843 18584 12885 18593
rect 12843 18544 12844 18584
rect 12884 18544 12885 18584
rect 12843 18535 12885 18544
rect 12844 18089 12884 18535
rect 12940 18509 12980 20056
rect 12939 18500 12981 18509
rect 12939 18460 12940 18500
rect 12980 18460 12981 18500
rect 12939 18451 12981 18460
rect 12843 18080 12885 18089
rect 12843 18040 12844 18080
rect 12884 18040 12885 18080
rect 12843 18031 12885 18040
rect 12459 17912 12501 17921
rect 12459 17872 12460 17912
rect 12500 17872 12501 17912
rect 12459 17863 12501 17872
rect 12747 17912 12789 17921
rect 12747 17872 12748 17912
rect 12788 17872 12789 17912
rect 12747 17863 12789 17872
rect 12459 17744 12501 17753
rect 12459 17704 12460 17744
rect 12500 17704 12501 17744
rect 12459 17695 12501 17704
rect 12556 17744 12596 17755
rect 12844 17753 12884 18031
rect 12939 17912 12981 17921
rect 12939 17872 12940 17912
rect 12980 17872 12981 17912
rect 12939 17863 12981 17872
rect 12460 16493 12500 17695
rect 12556 17669 12596 17704
rect 12652 17744 12692 17753
rect 12843 17744 12885 17753
rect 12692 17704 12788 17744
rect 12652 17695 12692 17704
rect 12555 17660 12597 17669
rect 12555 17620 12556 17660
rect 12596 17620 12597 17660
rect 12555 17611 12597 17620
rect 12748 17417 12788 17704
rect 12843 17704 12844 17744
rect 12884 17704 12885 17744
rect 12843 17695 12885 17704
rect 12843 17576 12885 17585
rect 12843 17536 12844 17576
rect 12884 17536 12885 17576
rect 12843 17527 12885 17536
rect 12747 17408 12789 17417
rect 12747 17368 12748 17408
rect 12788 17368 12789 17408
rect 12747 17359 12789 17368
rect 12459 16484 12501 16493
rect 12459 16444 12460 16484
rect 12500 16444 12501 16484
rect 12459 16435 12501 16444
rect 12459 16232 12501 16241
rect 12364 16192 12460 16232
rect 12500 16192 12501 16232
rect 12459 16183 12501 16192
rect 12267 15812 12309 15821
rect 12267 15772 12268 15812
rect 12308 15772 12309 15812
rect 12267 15763 12309 15772
rect 12363 14048 12405 14057
rect 12212 14008 12308 14048
rect 12172 13999 12212 14008
rect 12172 13208 12212 13217
rect 12076 13168 12172 13208
rect 12076 11789 12116 13168
rect 12172 13159 12212 13168
rect 12075 11780 12117 11789
rect 12075 11740 12076 11780
rect 12116 11740 12117 11780
rect 12075 11731 12117 11740
rect 11883 11612 11925 11621
rect 11883 11572 11884 11612
rect 11924 11572 11925 11612
rect 11883 11563 11925 11572
rect 11788 11528 11828 11537
rect 11596 11024 11636 11033
rect 11596 10445 11636 10984
rect 11788 10865 11828 11488
rect 11787 10856 11829 10865
rect 11787 10816 11788 10856
rect 11828 10816 11829 10856
rect 11787 10807 11829 10816
rect 11691 10772 11733 10781
rect 11691 10732 11692 10772
rect 11732 10732 11733 10772
rect 11691 10723 11733 10732
rect 11595 10436 11637 10445
rect 11595 10396 11596 10436
rect 11636 10396 11637 10436
rect 11595 10387 11637 10396
rect 11692 10268 11732 10723
rect 11500 10060 11636 10100
rect 11596 9521 11636 10060
rect 11595 9512 11637 9521
rect 11595 9472 11596 9512
rect 11636 9472 11637 9512
rect 11595 9463 11637 9472
rect 11500 9428 11540 9437
rect 11500 9260 11540 9388
rect 11596 9378 11636 9463
rect 11692 9260 11732 10228
rect 11788 10184 11828 10193
rect 11788 9689 11828 10144
rect 11787 9680 11829 9689
rect 11787 9640 11788 9680
rect 11828 9640 11829 9680
rect 11787 9631 11829 9640
rect 11787 9428 11829 9437
rect 11787 9388 11788 9428
rect 11828 9388 11829 9428
rect 11787 9379 11829 9388
rect 11500 9220 11732 9260
rect 11691 8924 11733 8933
rect 11691 8884 11692 8924
rect 11732 8884 11733 8924
rect 11691 8875 11733 8884
rect 11595 8756 11637 8765
rect 11595 8716 11596 8756
rect 11636 8716 11637 8756
rect 11595 8707 11637 8716
rect 11596 8672 11636 8707
rect 11596 8177 11636 8632
rect 11595 8168 11637 8177
rect 11595 8128 11596 8168
rect 11636 8128 11637 8168
rect 11595 8119 11637 8128
rect 11596 8000 11636 8009
rect 11404 7960 11596 8000
rect 11212 7916 11252 7960
rect 11596 7951 11636 7960
rect 11692 8000 11732 8875
rect 11212 7876 11444 7916
rect 11308 6488 11348 6497
rect 11308 5900 11348 6448
rect 11404 6488 11444 7876
rect 11692 7589 11732 7960
rect 11691 7580 11733 7589
rect 11691 7540 11692 7580
rect 11732 7540 11733 7580
rect 11691 7531 11733 7540
rect 11788 7253 11828 9379
rect 11787 7244 11829 7253
rect 11787 7204 11788 7244
rect 11828 7204 11829 7244
rect 11787 7195 11829 7204
rect 11595 7160 11637 7169
rect 11595 7120 11596 7160
rect 11636 7120 11637 7160
rect 11595 7111 11637 7120
rect 11444 6448 11540 6488
rect 11404 6439 11444 6448
rect 11404 5900 11444 5928
rect 11308 5860 11404 5900
rect 11500 5900 11540 6448
rect 11596 6077 11636 7111
rect 11787 6572 11829 6581
rect 11787 6532 11788 6572
rect 11828 6532 11829 6572
rect 11787 6523 11829 6532
rect 11788 6404 11828 6523
rect 11884 6488 11924 11563
rect 12268 10865 12308 14008
rect 12363 14008 12364 14048
rect 12404 14008 12405 14048
rect 12363 13999 12405 14008
rect 12364 13460 12404 13999
rect 12364 13411 12404 13420
rect 12267 10856 12309 10865
rect 12267 10816 12268 10856
rect 12308 10816 12309 10856
rect 12267 10807 12309 10816
rect 12267 10520 12309 10529
rect 12267 10480 12268 10520
rect 12308 10480 12309 10520
rect 12267 10471 12309 10480
rect 12171 10268 12213 10277
rect 12171 10228 12172 10268
rect 12212 10228 12213 10268
rect 12171 10219 12213 10228
rect 12172 9848 12212 10219
rect 12268 10184 12308 10471
rect 12308 10144 12404 10184
rect 12268 10135 12308 10144
rect 12172 9808 12308 9848
rect 12171 9680 12213 9689
rect 12171 9640 12172 9680
rect 12212 9640 12213 9680
rect 12171 9631 12213 9640
rect 12076 9512 12116 9523
rect 12076 9437 12116 9472
rect 12075 9428 12117 9437
rect 12075 9388 12076 9428
rect 12116 9388 12117 9428
rect 12075 9379 12117 9388
rect 11979 8840 12021 8849
rect 11979 8800 11980 8840
rect 12020 8800 12021 8840
rect 11979 8791 12021 8800
rect 11884 6439 11924 6448
rect 11788 6320 11828 6364
rect 11980 6320 12020 8791
rect 12075 8756 12117 8765
rect 12075 8716 12076 8756
rect 12116 8716 12117 8756
rect 12075 8707 12117 8716
rect 12076 8597 12116 8707
rect 12075 8588 12117 8597
rect 12075 8548 12076 8588
rect 12116 8548 12117 8588
rect 12075 8539 12117 8548
rect 12172 8168 12212 9631
rect 11788 6280 12020 6320
rect 12076 8128 12212 8168
rect 12076 6236 12116 8128
rect 12172 8000 12212 8009
rect 12172 7253 12212 7960
rect 12268 7757 12308 9808
rect 12267 7748 12309 7757
rect 12267 7708 12268 7748
rect 12308 7708 12309 7748
rect 12267 7699 12309 7708
rect 12267 7580 12309 7589
rect 12267 7540 12268 7580
rect 12308 7540 12309 7580
rect 12267 7531 12309 7540
rect 12171 7244 12213 7253
rect 12171 7204 12172 7244
rect 12212 7204 12213 7244
rect 12171 7195 12213 7204
rect 12171 7076 12213 7085
rect 12171 7036 12172 7076
rect 12212 7036 12213 7076
rect 12171 7027 12213 7036
rect 12172 6917 12212 7027
rect 12171 6908 12213 6917
rect 12171 6868 12172 6908
rect 12212 6868 12213 6908
rect 12171 6859 12213 6868
rect 11788 6196 12116 6236
rect 11595 6068 11637 6077
rect 11595 6028 11596 6068
rect 11636 6028 11637 6068
rect 11595 6019 11637 6028
rect 11500 5860 11636 5900
rect 11404 5851 11444 5860
rect 11212 5648 11252 5657
rect 11212 5489 11252 5608
rect 11403 5648 11445 5657
rect 11403 5608 11404 5648
rect 11444 5608 11445 5648
rect 11403 5599 11445 5608
rect 11211 5480 11253 5489
rect 11211 5440 11212 5480
rect 11252 5440 11253 5480
rect 11211 5431 11253 5440
rect 11404 5321 11444 5599
rect 11403 5312 11445 5321
rect 11596 5312 11636 5860
rect 11691 5648 11733 5657
rect 11691 5608 11692 5648
rect 11732 5608 11733 5648
rect 11691 5599 11733 5608
rect 11692 5514 11732 5599
rect 11403 5272 11404 5312
rect 11444 5272 11445 5312
rect 11403 5263 11445 5272
rect 11500 5272 11636 5312
rect 11691 5312 11733 5321
rect 11691 5272 11692 5312
rect 11732 5272 11733 5312
rect 11019 4976 11061 4985
rect 11019 4936 11020 4976
rect 11060 4936 11061 4976
rect 11019 4927 11061 4936
rect 11211 4976 11253 4985
rect 11211 4936 11212 4976
rect 11252 4936 11253 4976
rect 11211 4927 11253 4936
rect 10732 3928 10964 3968
rect 10636 1700 10676 1709
rect 10636 1289 10676 1660
rect 10732 1625 10772 3928
rect 11020 3884 11060 4927
rect 11212 4842 11252 4927
rect 11404 4724 11444 4733
rect 11404 4397 11444 4684
rect 11403 4388 11445 4397
rect 11403 4348 11404 4388
rect 11444 4348 11445 4388
rect 11403 4339 11445 4348
rect 11211 4304 11253 4313
rect 11211 4264 11212 4304
rect 11252 4264 11253 4304
rect 11211 4255 11253 4264
rect 11212 4136 11252 4255
rect 11212 4087 11252 4096
rect 10828 3844 11060 3884
rect 10828 3473 10868 3844
rect 11020 3548 11060 3557
rect 11060 3508 11348 3548
rect 11020 3499 11060 3508
rect 10827 3464 10869 3473
rect 10827 3424 10828 3464
rect 10868 3424 10869 3464
rect 10827 3415 10869 3424
rect 11308 3464 11348 3508
rect 11308 3415 11348 3424
rect 11404 3464 11444 3473
rect 11500 3464 11540 5272
rect 11691 5263 11733 5272
rect 11595 5060 11637 5069
rect 11595 5020 11596 5060
rect 11636 5020 11637 5060
rect 11595 5011 11637 5020
rect 11596 4976 11636 5011
rect 11596 4925 11636 4936
rect 11692 4808 11732 5263
rect 11444 3424 11540 3464
rect 11596 4768 11732 4808
rect 10828 3330 10868 3415
rect 11404 3137 11444 3424
rect 11403 3128 11445 3137
rect 11403 3088 11404 3128
rect 11444 3088 11445 3128
rect 11403 3079 11445 3088
rect 11115 2708 11157 2717
rect 11115 2668 11116 2708
rect 11156 2668 11157 2708
rect 11115 2659 11157 2668
rect 11116 2574 11156 2659
rect 11596 2624 11636 4768
rect 11691 4388 11733 4397
rect 11691 4348 11692 4388
rect 11732 4348 11733 4388
rect 11691 4339 11733 4348
rect 11692 4150 11732 4339
rect 11692 4101 11732 4110
rect 11788 3464 11828 6196
rect 11883 4220 11925 4229
rect 11883 4180 11884 4220
rect 11924 4180 11925 4220
rect 11883 4171 11925 4180
rect 11884 4052 11924 4171
rect 11884 4003 11924 4012
rect 11788 3389 11828 3424
rect 11884 3464 11924 3473
rect 12172 3464 12212 6859
rect 11924 3424 12212 3464
rect 11884 3415 11924 3424
rect 11787 3380 11829 3389
rect 11787 3340 11788 3380
rect 11828 3340 11829 3380
rect 11787 3331 11829 3340
rect 11788 3300 11828 3331
rect 11884 2624 11924 2633
rect 11596 2584 11884 2624
rect 11884 2575 11924 2584
rect 10924 2456 10964 2465
rect 10827 1700 10869 1709
rect 10827 1660 10828 1700
rect 10868 1660 10869 1700
rect 10827 1651 10869 1660
rect 10731 1616 10773 1625
rect 10731 1576 10732 1616
rect 10772 1576 10773 1616
rect 10731 1567 10773 1576
rect 10828 1566 10868 1651
rect 10731 1364 10773 1373
rect 10731 1324 10732 1364
rect 10772 1324 10773 1364
rect 10731 1315 10773 1324
rect 10635 1280 10677 1289
rect 10635 1240 10636 1280
rect 10676 1240 10677 1280
rect 10635 1231 10677 1240
rect 10484 1156 10580 1196
rect 10444 1147 10484 1156
rect 10635 944 10677 953
rect 10635 904 10636 944
rect 10676 904 10677 944
rect 10635 895 10677 904
rect 10443 860 10485 869
rect 10443 820 10444 860
rect 10484 820 10485 860
rect 10443 811 10485 820
rect 10347 356 10389 365
rect 10347 316 10348 356
rect 10388 316 10389 356
rect 10347 307 10389 316
rect 10444 80 10484 811
rect 10636 810 10676 895
rect 10732 608 10772 1315
rect 10827 1196 10869 1205
rect 10827 1156 10828 1196
rect 10868 1156 10869 1196
rect 10827 1147 10869 1156
rect 10828 1062 10868 1147
rect 10924 869 10964 2416
rect 11019 2456 11061 2465
rect 11019 2416 11020 2456
rect 11060 2416 11061 2456
rect 11019 2407 11061 2416
rect 11020 1868 11060 2407
rect 11020 1819 11060 1828
rect 11211 1868 11253 1877
rect 11211 1828 11212 1868
rect 11252 1828 11253 1868
rect 11211 1819 11253 1828
rect 11595 1868 11637 1877
rect 11595 1828 11596 1868
rect 11636 1828 11637 1868
rect 11595 1819 11637 1828
rect 12268 1868 12308 7531
rect 12364 6488 12404 10144
rect 12460 7169 12500 16183
rect 12651 16064 12693 16073
rect 12651 16024 12652 16064
rect 12692 16024 12693 16064
rect 12651 16015 12693 16024
rect 12556 9498 12596 9507
rect 12556 8849 12596 9458
rect 12555 8840 12597 8849
rect 12555 8800 12556 8840
rect 12596 8800 12597 8840
rect 12555 8791 12597 8800
rect 12652 8084 12692 16015
rect 12844 15560 12884 17527
rect 12844 15149 12884 15520
rect 12843 15140 12885 15149
rect 12843 15100 12844 15140
rect 12884 15100 12885 15140
rect 12843 15091 12885 15100
rect 12843 14972 12885 14981
rect 12843 14932 12844 14972
rect 12884 14932 12885 14972
rect 12843 14923 12885 14932
rect 12844 13553 12884 14923
rect 12843 13544 12885 13553
rect 12843 13504 12844 13544
rect 12884 13504 12885 13544
rect 12843 13495 12885 13504
rect 12844 12788 12884 13495
rect 12940 13301 12980 17863
rect 13036 14057 13076 26179
rect 13131 25136 13173 25145
rect 13131 25096 13132 25136
rect 13172 25096 13173 25136
rect 13131 25087 13173 25096
rect 13132 24044 13172 25087
rect 13228 24473 13268 28615
rect 13227 24464 13269 24473
rect 13227 24424 13228 24464
rect 13268 24424 13269 24464
rect 13227 24415 13269 24424
rect 13132 24004 13268 24044
rect 13131 23876 13173 23885
rect 13131 23836 13132 23876
rect 13172 23836 13173 23876
rect 13131 23827 13173 23836
rect 13132 23792 13172 23827
rect 13132 23741 13172 23752
rect 13228 23792 13268 24004
rect 13324 23969 13364 29380
rect 13323 23960 13365 23969
rect 13323 23920 13324 23960
rect 13364 23920 13365 23960
rect 13323 23911 13365 23920
rect 13268 23752 13364 23792
rect 13228 23743 13268 23752
rect 13227 22280 13269 22289
rect 13227 22240 13228 22280
rect 13268 22240 13269 22280
rect 13227 22231 13269 22240
rect 13324 22280 13364 23752
rect 13228 22146 13268 22231
rect 13324 22028 13364 22240
rect 13228 21988 13364 22028
rect 13228 19937 13268 21988
rect 13420 21029 13460 29464
rect 13516 29168 13556 29548
rect 13516 27824 13556 29128
rect 13612 29154 13652 29884
rect 13804 29840 13844 29959
rect 13804 29791 13844 29800
rect 13900 29840 13940 29849
rect 13940 29800 14132 29840
rect 13900 29791 13940 29800
rect 14092 29261 14132 29800
rect 13708 29252 13748 29261
rect 14091 29252 14133 29261
rect 13748 29212 14036 29252
rect 13708 29203 13748 29212
rect 13996 29188 14036 29212
rect 14091 29212 14092 29252
rect 14132 29212 14133 29252
rect 14091 29203 14133 29212
rect 13612 29114 13748 29154
rect 13996 29139 14036 29148
rect 14092 29188 14132 29203
rect 14092 29139 14132 29148
rect 13516 27784 13652 27824
rect 13516 27656 13556 27665
rect 13516 27161 13556 27616
rect 13515 27152 13557 27161
rect 13515 27112 13516 27152
rect 13556 27112 13557 27152
rect 13515 27103 13557 27112
rect 13612 26816 13652 27784
rect 13612 26405 13652 26776
rect 13611 26396 13653 26405
rect 13611 26356 13612 26396
rect 13652 26356 13653 26396
rect 13611 26347 13653 26356
rect 13515 25304 13557 25313
rect 13515 25264 13516 25304
rect 13556 25264 13557 25304
rect 13515 25255 13557 25264
rect 13516 25170 13556 25255
rect 13611 25220 13653 25229
rect 13611 25180 13612 25220
rect 13652 25180 13653 25220
rect 13611 25171 13653 25180
rect 13612 25086 13652 25171
rect 13708 24557 13748 29114
rect 14188 29084 14228 30463
rect 14284 29840 14324 29849
rect 14284 29513 14324 29800
rect 14379 29840 14421 29849
rect 14379 29800 14380 29840
rect 14420 29800 14421 29840
rect 14379 29791 14421 29800
rect 14380 29706 14420 29791
rect 14476 29588 14516 30631
rect 14571 29840 14613 29849
rect 14571 29800 14572 29840
rect 14612 29800 14613 29840
rect 14571 29791 14613 29800
rect 14380 29548 14516 29588
rect 14283 29504 14325 29513
rect 14283 29464 14284 29504
rect 14324 29464 14325 29504
rect 14283 29455 14325 29464
rect 14380 29336 14420 29548
rect 13900 29044 14228 29084
rect 14284 29296 14420 29336
rect 13803 28832 13845 28841
rect 13803 28792 13804 28832
rect 13844 28792 13845 28832
rect 13803 28783 13845 28792
rect 13804 27833 13844 28783
rect 13803 27824 13845 27833
rect 13803 27784 13804 27824
rect 13844 27784 13845 27824
rect 13803 27775 13845 27784
rect 13803 26816 13845 26825
rect 13803 26776 13804 26816
rect 13844 26776 13845 26816
rect 13803 26767 13845 26776
rect 13804 26732 13844 26767
rect 13804 26681 13844 26692
rect 13803 26396 13845 26405
rect 13803 26356 13804 26396
rect 13844 26356 13845 26396
rect 13803 26347 13845 26356
rect 13804 26144 13844 26347
rect 13804 26095 13844 26104
rect 13803 25724 13845 25733
rect 13803 25684 13804 25724
rect 13844 25684 13845 25724
rect 13803 25675 13845 25684
rect 13804 25304 13844 25675
rect 13900 25388 13940 29044
rect 13995 27740 14037 27749
rect 13995 27700 13996 27740
rect 14036 27700 14037 27740
rect 13995 27691 14037 27700
rect 13996 26312 14036 27691
rect 14187 27656 14229 27665
rect 14187 27616 14188 27656
rect 14228 27616 14229 27656
rect 14187 27607 14229 27616
rect 14188 27068 14228 27607
rect 14188 27019 14228 27028
rect 14091 26816 14133 26825
rect 14091 26776 14092 26816
rect 14132 26776 14133 26816
rect 14091 26767 14133 26776
rect 14092 26682 14132 26767
rect 13996 26263 14036 26272
rect 14188 26648 14228 26657
rect 14188 26144 14228 26608
rect 14284 26321 14324 29296
rect 14475 29252 14517 29261
rect 14475 29212 14476 29252
rect 14516 29212 14517 29252
rect 14475 29203 14517 29212
rect 14476 29168 14516 29203
rect 14476 29117 14516 29128
rect 14572 29168 14612 29791
rect 14476 28328 14516 28337
rect 14380 28160 14420 28169
rect 14380 26405 14420 28120
rect 14476 27749 14516 28288
rect 14475 27740 14517 27749
rect 14475 27700 14476 27740
rect 14516 27700 14517 27740
rect 14475 27691 14517 27700
rect 14572 27077 14612 29128
rect 14668 28328 14708 31051
rect 14764 29261 14804 31135
rect 14860 29840 14900 31144
rect 14956 30269 14996 34252
rect 15052 33872 15092 34336
rect 15147 34208 15189 34217
rect 15147 34168 15148 34208
rect 15188 34168 15189 34208
rect 15147 34159 15189 34168
rect 15148 34074 15188 34159
rect 15052 33823 15092 33832
rect 15244 32696 15284 34663
rect 15532 34376 15572 34385
rect 15435 33704 15477 33713
rect 15435 33664 15436 33704
rect 15476 33664 15477 33704
rect 15435 33655 15477 33664
rect 15339 33620 15381 33629
rect 15339 33580 15340 33620
rect 15380 33580 15381 33620
rect 15339 33571 15381 33580
rect 15340 32873 15380 33571
rect 15436 33125 15476 33655
rect 15435 33116 15477 33125
rect 15435 33076 15436 33116
rect 15476 33076 15477 33116
rect 15435 33067 15477 33076
rect 15532 32948 15572 34336
rect 15628 33041 15668 35176
rect 15627 33032 15669 33041
rect 15627 32992 15628 33032
rect 15668 32992 15669 33032
rect 15820 33032 15860 35419
rect 15915 35132 15957 35141
rect 15915 35092 15916 35132
rect 15956 35092 15957 35132
rect 15915 35083 15957 35092
rect 16012 35132 16052 36595
rect 15916 34998 15956 35083
rect 16012 34217 16052 35092
rect 16011 34208 16053 34217
rect 16011 34168 16012 34208
rect 16052 34168 16053 34208
rect 16011 34159 16053 34168
rect 16011 33032 16053 33041
rect 15820 32992 15956 33032
rect 15627 32983 15669 32992
rect 15436 32908 15572 32948
rect 15339 32864 15381 32873
rect 15339 32824 15340 32864
rect 15380 32824 15381 32864
rect 15339 32815 15381 32824
rect 15244 32656 15380 32696
rect 15051 32024 15093 32033
rect 15051 31984 15052 32024
rect 15092 31984 15093 32024
rect 15051 31975 15093 31984
rect 15052 31109 15092 31975
rect 15243 31436 15285 31445
rect 15243 31396 15244 31436
rect 15284 31396 15285 31436
rect 15243 31387 15285 31396
rect 15147 31352 15189 31361
rect 15147 31312 15148 31352
rect 15188 31312 15189 31352
rect 15147 31303 15189 31312
rect 15244 31352 15284 31387
rect 15148 31218 15188 31303
rect 15244 31301 15284 31312
rect 15340 31184 15380 32656
rect 15436 32612 15476 32908
rect 15916 32873 15956 32992
rect 16011 32992 16012 33032
rect 16052 32992 16053 33032
rect 16011 32983 16053 32992
rect 15820 32864 15860 32873
rect 15532 32780 15572 32789
rect 15820 32780 15860 32824
rect 15915 32864 15957 32873
rect 15915 32824 15916 32864
rect 15956 32824 15957 32864
rect 15915 32815 15957 32824
rect 15572 32740 15860 32780
rect 15532 32731 15572 32740
rect 15436 32572 15572 32612
rect 15435 31520 15477 31529
rect 15435 31480 15436 31520
rect 15476 31480 15477 31520
rect 15435 31471 15477 31480
rect 15244 31144 15380 31184
rect 15436 31184 15476 31471
rect 15051 31100 15093 31109
rect 15051 31060 15052 31100
rect 15092 31060 15093 31100
rect 15051 31051 15093 31060
rect 15147 31016 15189 31025
rect 15147 30976 15148 31016
rect 15188 30976 15189 31016
rect 15147 30967 15189 30976
rect 14955 30260 14997 30269
rect 14955 30220 14956 30260
rect 14996 30220 14997 30260
rect 14955 30211 14997 30220
rect 14900 29800 15092 29840
rect 14860 29791 14900 29800
rect 14763 29252 14805 29261
rect 14763 29212 14764 29252
rect 14804 29212 14805 29252
rect 14763 29203 14805 29212
rect 14764 29084 14804 29203
rect 15052 29168 15092 29800
rect 15052 29119 15092 29128
rect 14764 29044 14900 29084
rect 14668 28253 14708 28288
rect 14667 28244 14709 28253
rect 14667 28204 14668 28244
rect 14708 28204 14709 28244
rect 14667 28195 14709 28204
rect 14764 27656 14804 27665
rect 14668 27616 14764 27656
rect 14668 27413 14708 27616
rect 14764 27607 14804 27616
rect 14667 27404 14709 27413
rect 14667 27364 14668 27404
rect 14708 27364 14709 27404
rect 14667 27355 14709 27364
rect 14571 27068 14613 27077
rect 14571 27028 14572 27068
rect 14612 27028 14613 27068
rect 14571 27019 14613 27028
rect 14475 26816 14517 26825
rect 14475 26776 14476 26816
rect 14516 26776 14612 26816
rect 14475 26767 14517 26776
rect 14476 26682 14516 26767
rect 14379 26396 14421 26405
rect 14379 26356 14380 26396
rect 14420 26356 14421 26396
rect 14379 26347 14421 26356
rect 14283 26312 14325 26321
rect 14283 26272 14284 26312
rect 14324 26272 14325 26312
rect 14283 26263 14325 26272
rect 14475 26312 14517 26321
rect 14475 26272 14476 26312
rect 14516 26272 14517 26312
rect 14475 26263 14517 26272
rect 14476 26178 14516 26263
rect 14188 25733 14228 26104
rect 14284 26144 14324 26153
rect 14284 25901 14324 26104
rect 14380 26144 14420 26153
rect 14572 26144 14612 26776
rect 14668 26489 14708 27355
rect 14860 27320 14900 29044
rect 15148 27824 15188 30967
rect 15052 27784 15188 27824
rect 14764 27280 14900 27320
rect 14956 27404 14996 27413
rect 14764 26816 14804 27280
rect 14859 27068 14901 27077
rect 14859 27028 14860 27068
rect 14900 27028 14901 27068
rect 14859 27019 14901 27028
rect 14667 26480 14709 26489
rect 14667 26440 14668 26480
rect 14708 26440 14709 26480
rect 14667 26431 14709 26440
rect 14764 26312 14804 26776
rect 14860 26816 14900 27019
rect 14860 26767 14900 26776
rect 14956 26489 14996 27364
rect 15052 27245 15092 27784
rect 15147 27656 15189 27665
rect 15147 27616 15148 27656
rect 15188 27616 15189 27656
rect 15147 27607 15189 27616
rect 15244 27656 15284 31144
rect 15436 31135 15476 31144
rect 15532 30605 15572 32572
rect 15724 32192 15764 32740
rect 15916 32730 15956 32815
rect 15916 32192 15956 32201
rect 15724 32152 15916 32192
rect 15916 32143 15956 32152
rect 16012 32192 16052 32983
rect 16012 31109 16052 32152
rect 16011 31100 16053 31109
rect 16011 31060 16012 31100
rect 16052 31060 16053 31100
rect 16011 31051 16053 31060
rect 16108 31025 16148 37267
rect 16107 31016 16149 31025
rect 16107 30976 16108 31016
rect 16148 30976 16149 31016
rect 16107 30967 16149 30976
rect 15723 30932 15765 30941
rect 15723 30892 15724 30932
rect 15764 30892 15765 30932
rect 15723 30883 15765 30892
rect 15724 30680 15764 30883
rect 15724 30605 15764 30640
rect 15531 30596 15573 30605
rect 15531 30556 15532 30596
rect 15572 30556 15573 30596
rect 15531 30547 15573 30556
rect 15723 30596 15765 30605
rect 15723 30556 15724 30596
rect 15764 30556 15765 30596
rect 15723 30547 15765 30556
rect 15724 30516 15764 30547
rect 15916 30428 15956 30437
rect 15627 30260 15669 30269
rect 15627 30220 15628 30260
rect 15668 30220 15669 30260
rect 15627 30211 15669 30220
rect 15339 29924 15381 29933
rect 15339 29884 15340 29924
rect 15380 29884 15381 29924
rect 15339 29875 15381 29884
rect 15340 29854 15380 29875
rect 15340 29789 15380 29814
rect 15531 29756 15573 29765
rect 15531 29716 15532 29756
rect 15572 29716 15573 29756
rect 15531 29707 15573 29716
rect 15532 29622 15572 29707
rect 15532 29154 15572 29163
rect 15532 28589 15572 29114
rect 15531 28580 15573 28589
rect 15531 28540 15532 28580
rect 15572 28540 15573 28580
rect 15531 28531 15573 28540
rect 15628 27992 15668 30211
rect 15916 29933 15956 30388
rect 16011 30428 16053 30437
rect 16011 30388 16012 30428
rect 16052 30388 16053 30428
rect 16011 30379 16053 30388
rect 15915 29924 15957 29933
rect 15915 29884 15916 29924
rect 15956 29884 15957 29924
rect 15915 29875 15957 29884
rect 15724 29840 15764 29849
rect 15764 29800 15860 29840
rect 15724 29791 15764 29800
rect 15820 29345 15860 29800
rect 15819 29336 15861 29345
rect 15819 29296 15820 29336
rect 15860 29296 15861 29336
rect 15819 29287 15861 29296
rect 15723 29252 15765 29261
rect 15723 29212 15724 29252
rect 15764 29212 15765 29252
rect 15723 29203 15765 29212
rect 15724 29118 15764 29203
rect 15532 27952 15668 27992
rect 15916 28328 15956 28337
rect 15339 27740 15381 27749
rect 15339 27700 15340 27740
rect 15380 27700 15381 27740
rect 15339 27691 15381 27700
rect 15148 27522 15188 27607
rect 15244 27245 15284 27616
rect 15340 27656 15380 27691
rect 15340 27605 15380 27616
rect 15435 27656 15477 27665
rect 15435 27616 15436 27656
rect 15476 27616 15477 27656
rect 15435 27607 15477 27616
rect 15436 27522 15476 27607
rect 15051 27236 15093 27245
rect 15051 27196 15052 27236
rect 15092 27196 15093 27236
rect 15051 27187 15093 27196
rect 15243 27236 15285 27245
rect 15243 27196 15244 27236
rect 15284 27196 15285 27236
rect 15243 27187 15285 27196
rect 15051 26984 15093 26993
rect 15051 26944 15052 26984
rect 15092 26944 15093 26984
rect 15051 26935 15093 26944
rect 15148 26984 15188 26993
rect 15532 26984 15572 27952
rect 15724 27656 15764 27665
rect 15724 27245 15764 27616
rect 15819 27488 15861 27497
rect 15819 27448 15820 27488
rect 15860 27448 15861 27488
rect 15819 27439 15861 27448
rect 15723 27236 15765 27245
rect 15723 27196 15724 27236
rect 15764 27196 15765 27236
rect 15820 27236 15860 27439
rect 15916 27413 15956 28288
rect 15915 27404 15957 27413
rect 15915 27364 15916 27404
rect 15956 27364 15957 27404
rect 15915 27355 15957 27364
rect 15820 27196 15956 27236
rect 15723 27187 15765 27196
rect 15916 27068 15956 27196
rect 15916 27019 15956 27028
rect 14955 26480 14997 26489
rect 14955 26440 14956 26480
rect 14996 26440 14997 26480
rect 14955 26431 14997 26440
rect 14764 26272 14900 26312
rect 14764 26144 14804 26153
rect 14572 26104 14764 26144
rect 14283 25892 14325 25901
rect 14283 25852 14284 25892
rect 14324 25852 14325 25892
rect 14283 25843 14325 25852
rect 14187 25724 14229 25733
rect 14187 25684 14188 25724
rect 14228 25684 14229 25724
rect 14187 25675 14229 25684
rect 14092 25556 14132 25565
rect 14380 25556 14420 26104
rect 14132 25516 14420 25556
rect 14092 25507 14132 25516
rect 14091 25388 14133 25397
rect 13900 25348 14036 25388
rect 13804 25255 13844 25264
rect 13900 25262 13940 25271
rect 13899 25222 13900 25229
rect 13940 25222 13941 25229
rect 13899 25220 13941 25222
rect 13899 25180 13900 25220
rect 13940 25180 13941 25220
rect 13899 25171 13941 25180
rect 13900 25127 13940 25171
rect 13900 24641 13940 24726
rect 13899 24632 13941 24641
rect 13899 24592 13900 24632
rect 13940 24592 13941 24632
rect 13899 24583 13941 24592
rect 13707 24548 13749 24557
rect 13707 24508 13708 24548
rect 13748 24508 13749 24548
rect 13707 24499 13749 24508
rect 13899 24464 13941 24473
rect 13899 24424 13900 24464
rect 13940 24424 13941 24464
rect 13899 24415 13941 24424
rect 13707 23960 13749 23969
rect 13707 23920 13708 23960
rect 13748 23920 13749 23960
rect 13707 23911 13749 23920
rect 13708 23876 13748 23911
rect 13612 23792 13652 23801
rect 13612 23381 13652 23752
rect 13611 23372 13653 23381
rect 13611 23332 13612 23372
rect 13652 23332 13653 23372
rect 13611 23323 13653 23332
rect 13708 23204 13748 23836
rect 13803 23792 13845 23801
rect 13803 23752 13804 23792
rect 13844 23752 13845 23792
rect 13803 23743 13845 23752
rect 13804 23633 13844 23743
rect 13803 23624 13845 23633
rect 13803 23584 13804 23624
rect 13844 23584 13845 23624
rect 13803 23575 13845 23584
rect 13900 23288 13940 24415
rect 13612 23164 13748 23204
rect 13804 23248 13940 23288
rect 13612 22196 13652 23164
rect 13804 22868 13844 23248
rect 13899 23120 13941 23129
rect 13899 23080 13900 23120
rect 13940 23080 13941 23120
rect 13899 23071 13941 23080
rect 13900 22986 13940 23071
rect 13804 22828 13940 22868
rect 13708 22373 13748 22458
rect 13707 22364 13749 22373
rect 13707 22324 13708 22364
rect 13748 22324 13749 22364
rect 13707 22315 13749 22324
rect 13804 22280 13844 22289
rect 13804 22196 13844 22240
rect 13612 22156 13844 22196
rect 13612 21197 13652 22156
rect 13611 21188 13653 21197
rect 13611 21148 13612 21188
rect 13652 21148 13653 21188
rect 13611 21139 13653 21148
rect 13419 21020 13461 21029
rect 13419 20980 13420 21020
rect 13460 20980 13461 21020
rect 13419 20971 13461 20980
rect 13611 21020 13653 21029
rect 13611 20980 13612 21020
rect 13652 20980 13653 21020
rect 13611 20971 13653 20980
rect 13324 20777 13364 20862
rect 13323 20768 13365 20777
rect 13323 20728 13324 20768
rect 13364 20728 13365 20768
rect 13323 20719 13365 20728
rect 13612 20180 13652 20971
rect 13516 20140 13652 20180
rect 13900 20180 13940 22828
rect 13996 22037 14036 25348
rect 14091 25348 14092 25388
rect 14132 25348 14133 25388
rect 14091 25339 14133 25348
rect 14092 25304 14132 25339
rect 14092 25253 14132 25264
rect 14284 25304 14324 25313
rect 14284 24800 14324 25264
rect 14476 25304 14516 25313
rect 14379 25220 14421 25229
rect 14379 25180 14380 25220
rect 14420 25180 14421 25220
rect 14379 25171 14421 25180
rect 14380 25086 14420 25171
rect 14380 24800 14420 24809
rect 14284 24760 14380 24800
rect 14380 24751 14420 24760
rect 14284 24632 14324 24641
rect 14476 24632 14516 25264
rect 14572 25304 14612 25313
rect 14572 24809 14612 25264
rect 14571 24800 14613 24809
rect 14571 24760 14572 24800
rect 14612 24760 14613 24800
rect 14571 24751 14613 24760
rect 14324 24592 14516 24632
rect 14571 24632 14613 24641
rect 14571 24592 14572 24632
rect 14612 24592 14613 24632
rect 14668 24632 14708 26104
rect 14764 26095 14804 26104
rect 14860 25649 14900 26272
rect 15052 26153 15092 26935
rect 15148 26825 15188 26944
rect 15244 26944 15476 26984
rect 15147 26816 15189 26825
rect 15147 26776 15148 26816
rect 15188 26776 15189 26816
rect 15147 26767 15189 26776
rect 15244 26321 15284 26944
rect 15436 26919 15476 26944
rect 15532 26935 15572 26944
rect 15723 26984 15765 26993
rect 15723 26944 15724 26984
rect 15764 26944 15765 26984
rect 15723 26935 15765 26944
rect 15436 26910 15477 26919
rect 15436 26870 15437 26910
rect 15436 26860 15477 26870
rect 15628 26900 15668 26909
rect 15340 26816 15380 26827
rect 15340 26741 15380 26776
rect 15339 26732 15381 26741
rect 15339 26692 15340 26732
rect 15380 26692 15381 26732
rect 15339 26683 15381 26692
rect 15628 26564 15668 26860
rect 15724 26858 15764 26935
rect 15724 26809 15764 26818
rect 15532 26524 15668 26564
rect 15243 26312 15285 26321
rect 15243 26272 15244 26312
rect 15284 26272 15285 26312
rect 15243 26263 15285 26272
rect 15051 26144 15093 26153
rect 15051 26104 15052 26144
rect 15092 26104 15093 26144
rect 15051 26095 15093 26104
rect 15148 26144 15188 26153
rect 15148 25976 15188 26104
rect 15052 25936 15188 25976
rect 14859 25640 14901 25649
rect 14859 25600 14860 25640
rect 14900 25600 14901 25640
rect 14859 25591 14901 25600
rect 15052 25481 15092 25936
rect 15436 25892 15476 25901
rect 15244 25852 15436 25892
rect 15051 25472 15093 25481
rect 15051 25432 15052 25472
rect 15092 25432 15093 25472
rect 15051 25423 15093 25432
rect 14764 25304 14804 25313
rect 14764 24809 14804 25264
rect 14860 25304 14900 25315
rect 14860 25229 14900 25264
rect 14956 25304 14996 25313
rect 14859 25220 14901 25229
rect 14859 25180 14860 25220
rect 14900 25180 14901 25220
rect 14859 25171 14901 25180
rect 14763 24800 14805 24809
rect 14763 24760 14764 24800
rect 14804 24760 14805 24800
rect 14956 24800 14996 25264
rect 15244 25304 15284 25852
rect 15436 25843 15476 25852
rect 15435 25724 15477 25733
rect 15435 25684 15436 25724
rect 15476 25684 15477 25724
rect 15435 25675 15477 25684
rect 15339 25388 15381 25397
rect 15339 25348 15340 25388
rect 15380 25348 15381 25388
rect 15339 25339 15381 25348
rect 15244 25255 15284 25264
rect 15340 25304 15380 25339
rect 15340 25253 15380 25264
rect 15051 25220 15093 25229
rect 15051 25180 15052 25220
rect 15092 25180 15093 25220
rect 15051 25171 15093 25180
rect 15052 25086 15092 25171
rect 15339 24800 15381 24809
rect 14956 24760 15092 24800
rect 14763 24751 14805 24760
rect 14668 24619 14804 24632
rect 14668 24592 14764 24619
rect 14092 24380 14132 24389
rect 14284 24380 14324 24592
rect 14571 24583 14613 24592
rect 14572 24498 14612 24583
rect 14764 24570 14804 24579
rect 14860 24557 14900 24642
rect 14955 24632 14997 24641
rect 14955 24592 14956 24632
rect 14996 24592 14997 24632
rect 14955 24583 14997 24592
rect 14859 24548 14901 24557
rect 14859 24508 14860 24548
rect 14900 24508 14901 24548
rect 14859 24499 14901 24508
rect 14956 24498 14996 24583
rect 14379 24464 14421 24473
rect 14379 24424 14380 24464
rect 14420 24424 14421 24464
rect 14379 24415 14421 24424
rect 14132 24340 14324 24380
rect 14092 23801 14132 24340
rect 14091 23792 14133 23801
rect 14091 23752 14092 23792
rect 14132 23752 14133 23792
rect 14091 23743 14133 23752
rect 14188 23792 14228 23803
rect 14188 23717 14228 23752
rect 14187 23708 14229 23717
rect 14187 23668 14188 23708
rect 14228 23668 14229 23708
rect 14187 23659 14229 23668
rect 14091 23624 14133 23633
rect 14091 23584 14092 23624
rect 14132 23584 14133 23624
rect 14091 23575 14133 23584
rect 13995 22028 14037 22037
rect 13995 21988 13996 22028
rect 14036 21988 14037 22028
rect 13995 21979 14037 21988
rect 14092 20189 14132 23575
rect 14188 22280 14228 23659
rect 14380 23549 14420 24415
rect 14955 24380 14997 24389
rect 14955 24340 14956 24380
rect 14996 24340 14997 24380
rect 14955 24331 14997 24340
rect 14571 24296 14613 24305
rect 14571 24256 14572 24296
rect 14612 24256 14613 24296
rect 14571 24247 14613 24256
rect 14379 23540 14421 23549
rect 14379 23500 14380 23540
rect 14420 23500 14421 23540
rect 14379 23491 14421 23500
rect 14380 23129 14420 23491
rect 14379 23120 14421 23129
rect 14379 23080 14380 23120
rect 14420 23080 14421 23120
rect 14379 23071 14421 23080
rect 14475 22700 14517 22709
rect 14475 22660 14476 22700
rect 14516 22660 14517 22700
rect 14475 22651 14517 22660
rect 14284 22280 14324 22289
rect 14188 22240 14284 22280
rect 14284 22231 14324 22240
rect 14379 22280 14421 22289
rect 14379 22240 14380 22280
rect 14420 22240 14421 22280
rect 14379 22231 14421 22240
rect 14283 22028 14325 22037
rect 14283 21988 14284 22028
rect 14324 21988 14325 22028
rect 14283 21979 14325 21988
rect 14188 21608 14228 21617
rect 14188 21029 14228 21568
rect 14187 21020 14229 21029
rect 14187 20980 14188 21020
rect 14228 20980 14229 21020
rect 14187 20971 14229 20980
rect 14091 20180 14133 20189
rect 13900 20140 14036 20180
rect 13227 19928 13269 19937
rect 13227 19888 13228 19928
rect 13268 19888 13269 19928
rect 13227 19879 13269 19888
rect 13227 19760 13269 19769
rect 13227 19720 13228 19760
rect 13268 19720 13269 19760
rect 13227 19711 13269 19720
rect 13131 17744 13173 17753
rect 13131 17704 13132 17744
rect 13172 17704 13173 17744
rect 13131 17695 13173 17704
rect 13132 17610 13172 17695
rect 13131 16400 13173 16409
rect 13131 16360 13132 16400
rect 13172 16360 13173 16400
rect 13131 16351 13173 16360
rect 13132 16232 13172 16351
rect 13132 15653 13172 16192
rect 13131 15644 13173 15653
rect 13131 15604 13132 15644
rect 13172 15604 13173 15644
rect 13131 15595 13173 15604
rect 13035 14048 13077 14057
rect 13035 14008 13036 14048
rect 13076 14008 13077 14048
rect 13035 13999 13077 14008
rect 12939 13292 12981 13301
rect 12939 13252 12940 13292
rect 12980 13252 12981 13292
rect 12939 13243 12981 13252
rect 13036 13208 13076 13217
rect 12844 12748 12980 12788
rect 12844 12536 12884 12545
rect 12844 12125 12884 12496
rect 12940 12461 12980 12748
rect 13036 12704 13076 13168
rect 13036 12655 13076 12664
rect 13132 13208 13172 13217
rect 13228 13208 13268 19711
rect 13516 18836 13556 20140
rect 13899 20012 13941 20021
rect 13899 19972 13900 20012
rect 13940 19972 13941 20012
rect 13899 19963 13941 19972
rect 13420 18796 13556 18836
rect 13323 18584 13365 18593
rect 13323 18544 13324 18584
rect 13364 18544 13365 18584
rect 13323 18535 13365 18544
rect 13324 18450 13364 18535
rect 13324 17072 13364 17081
rect 13324 16409 13364 17032
rect 13323 16400 13365 16409
rect 13323 16360 13324 16400
rect 13364 16360 13365 16400
rect 13323 16351 13365 16360
rect 13420 16316 13460 18796
rect 13900 18752 13940 19963
rect 13996 19928 14036 20140
rect 14091 20140 14092 20180
rect 14132 20140 14133 20180
rect 14091 20131 14133 20140
rect 14188 20096 14228 20105
rect 14284 20096 14324 21979
rect 14380 21776 14420 22231
rect 14380 21727 14420 21736
rect 14379 20096 14421 20105
rect 14284 20056 14380 20096
rect 14420 20056 14421 20096
rect 14188 20012 14228 20056
rect 14379 20047 14421 20056
rect 14188 19972 14324 20012
rect 13996 19888 14228 19928
rect 13995 19760 14037 19769
rect 13995 19720 13996 19760
rect 14036 19720 14037 19760
rect 13995 19711 14037 19720
rect 13996 19256 14036 19711
rect 14091 19676 14133 19685
rect 14091 19636 14092 19676
rect 14132 19636 14133 19676
rect 14091 19627 14133 19636
rect 13996 19207 14036 19216
rect 14092 19256 14132 19627
rect 13900 18712 14036 18752
rect 13516 18668 13556 18677
rect 13556 18628 13844 18668
rect 13516 18619 13556 18628
rect 13804 18584 13844 18628
rect 13804 18535 13844 18544
rect 13899 18584 13941 18593
rect 13899 18544 13900 18584
rect 13940 18544 13941 18584
rect 13899 18535 13941 18544
rect 13803 17912 13845 17921
rect 13803 17872 13804 17912
rect 13844 17872 13845 17912
rect 13803 17863 13845 17872
rect 13612 17749 13652 17758
rect 13516 17240 13556 17249
rect 13612 17240 13652 17709
rect 13804 17660 13844 17863
rect 13900 17837 13940 18535
rect 13899 17828 13941 17837
rect 13899 17788 13900 17828
rect 13940 17788 13941 17828
rect 13899 17779 13941 17788
rect 13804 17611 13844 17620
rect 13900 17324 13940 17779
rect 13556 17200 13652 17240
rect 13708 17284 13940 17324
rect 13516 17191 13556 17200
rect 13611 16316 13653 16325
rect 13420 16276 13556 16316
rect 13323 16241 13365 16250
rect 13323 16201 13324 16241
rect 13364 16201 13365 16241
rect 13323 16192 13365 16201
rect 13324 16148 13364 16192
rect 13324 16099 13364 16108
rect 13323 15980 13365 15989
rect 13323 15940 13324 15980
rect 13364 15940 13365 15980
rect 13323 15931 13365 15940
rect 13172 13168 13268 13208
rect 12939 12452 12981 12461
rect 12939 12412 12940 12452
rect 12980 12412 12981 12452
rect 12939 12403 12981 12412
rect 13132 12368 13172 13168
rect 13228 12545 13268 12630
rect 13227 12536 13269 12545
rect 13227 12496 13228 12536
rect 13268 12496 13269 12536
rect 13227 12487 13269 12496
rect 13132 12328 13268 12368
rect 13131 12200 13173 12209
rect 13131 12160 13132 12200
rect 13172 12160 13173 12200
rect 13131 12151 13173 12160
rect 12843 12116 12885 12125
rect 12843 12076 12844 12116
rect 12884 12076 12885 12116
rect 12843 12067 12885 12076
rect 12843 11696 12885 11705
rect 12843 11656 12844 11696
rect 12884 11656 12885 11696
rect 12843 11647 12885 11656
rect 12844 11024 12884 11647
rect 12844 10975 12884 10984
rect 13036 10772 13076 10781
rect 12844 10732 13036 10772
rect 12844 10268 12884 10732
rect 13036 10723 13076 10732
rect 13132 10352 13172 12151
rect 13228 10436 13268 12328
rect 13324 10613 13364 15931
rect 13420 14048 13460 14059
rect 13420 13973 13460 14008
rect 13419 13964 13461 13973
rect 13419 13924 13420 13964
rect 13460 13924 13461 13964
rect 13419 13915 13461 13924
rect 13516 13292 13556 16276
rect 13611 16276 13612 16316
rect 13652 16276 13653 16316
rect 13611 16267 13653 16276
rect 13612 16232 13652 16267
rect 13612 16181 13652 16192
rect 13708 16232 13748 17284
rect 13708 15989 13748 16192
rect 13803 16232 13845 16241
rect 13803 16192 13804 16232
rect 13844 16192 13845 16232
rect 13803 16183 13845 16192
rect 13707 15980 13749 15989
rect 13707 15940 13708 15980
rect 13748 15940 13749 15980
rect 13707 15931 13749 15940
rect 13612 14720 13652 14729
rect 13612 14216 13652 14680
rect 13612 14167 13652 14176
rect 13708 14720 13748 14729
rect 13804 14720 13844 16183
rect 13899 15560 13941 15569
rect 13899 15520 13900 15560
rect 13940 15520 13941 15560
rect 13899 15511 13941 15520
rect 13900 15426 13940 15511
rect 13748 14680 13844 14720
rect 13516 13243 13556 13252
rect 13419 13208 13461 13217
rect 13419 13168 13420 13208
rect 13460 13168 13461 13208
rect 13419 13159 13461 13168
rect 13611 13208 13653 13217
rect 13611 13168 13612 13208
rect 13652 13168 13653 13208
rect 13611 13159 13653 13168
rect 13323 10604 13365 10613
rect 13323 10564 13324 10604
rect 13364 10564 13365 10604
rect 13323 10555 13365 10564
rect 13228 10396 13364 10436
rect 13132 10312 13268 10352
rect 12796 10228 12884 10268
rect 12939 10268 12981 10277
rect 12939 10228 12940 10268
rect 12980 10228 12981 10268
rect 12796 10226 12836 10228
rect 12939 10219 12981 10228
rect 12796 10177 12836 10186
rect 12940 10100 12980 10219
rect 13131 10184 13173 10193
rect 13131 10144 13132 10184
rect 13172 10144 13173 10184
rect 13131 10135 13173 10144
rect 12940 10051 12980 10060
rect 13132 10050 13172 10135
rect 12747 9596 12789 9605
rect 12747 9556 12748 9596
rect 12788 9556 12789 9596
rect 12747 9547 12789 9556
rect 12748 9462 12788 9547
rect 13035 8840 13077 8849
rect 13035 8800 13036 8840
rect 13076 8800 13077 8840
rect 13035 8791 13077 8800
rect 12844 8765 12884 8767
rect 12843 8756 12885 8765
rect 12843 8716 12844 8756
rect 12884 8716 12885 8756
rect 12843 8707 12885 8716
rect 12844 8672 12884 8707
rect 13036 8706 13076 8791
rect 12844 8623 12884 8632
rect 12844 8093 12884 8178
rect 12604 8044 12692 8084
rect 12843 8084 12885 8093
rect 12843 8044 12844 8084
rect 12884 8044 12885 8084
rect 12604 7832 12644 8044
rect 12843 8035 12885 8044
rect 12700 7958 12740 7967
rect 12700 7916 12740 7918
rect 12700 7876 13076 7916
rect 12604 7792 12692 7832
rect 12459 7160 12501 7169
rect 12459 7120 12460 7160
rect 12500 7120 12501 7160
rect 12459 7111 12501 7120
rect 12555 6656 12597 6665
rect 12555 6616 12556 6656
rect 12596 6616 12597 6656
rect 12555 6607 12597 6616
rect 12364 3464 12404 6448
rect 12556 3977 12596 6607
rect 12555 3968 12597 3977
rect 12555 3928 12556 3968
rect 12596 3928 12597 3968
rect 12555 3919 12597 3928
rect 12364 2969 12404 3424
rect 12363 2960 12405 2969
rect 12363 2920 12364 2960
rect 12404 2920 12405 2960
rect 12363 2911 12405 2920
rect 12459 2288 12501 2297
rect 12459 2248 12460 2288
rect 12500 2248 12501 2288
rect 12459 2239 12501 2248
rect 12460 1952 12500 2239
rect 12460 1903 12500 1912
rect 12268 1819 12308 1828
rect 11212 1734 11252 1819
rect 11596 1734 11636 1819
rect 12652 1709 12692 7792
rect 13036 7412 13076 7876
rect 13036 7363 13076 7372
rect 12843 7160 12885 7169
rect 12843 7120 12844 7160
rect 12884 7120 12885 7160
rect 12843 7111 12885 7120
rect 12844 7026 12884 7111
rect 13228 6833 13268 10312
rect 13324 7673 13364 10396
rect 13420 8672 13460 13159
rect 13612 13074 13652 13159
rect 13515 12536 13557 12545
rect 13515 12496 13516 12536
rect 13556 12496 13557 12536
rect 13515 12487 13557 12496
rect 13516 11360 13556 12487
rect 13708 12209 13748 14680
rect 13803 14048 13845 14057
rect 13803 14008 13804 14048
rect 13844 14008 13845 14048
rect 13803 13999 13845 14008
rect 13707 12200 13749 12209
rect 13707 12160 13708 12200
rect 13748 12160 13749 12200
rect 13707 12151 13749 12160
rect 13516 11320 13748 11360
rect 13515 10520 13557 10529
rect 13515 10480 13516 10520
rect 13556 10480 13557 10520
rect 13515 10471 13557 10480
rect 13420 8345 13460 8632
rect 13419 8336 13461 8345
rect 13419 8296 13420 8336
rect 13460 8296 13461 8336
rect 13419 8287 13461 8296
rect 13323 7664 13365 7673
rect 13323 7624 13324 7664
rect 13364 7624 13365 7664
rect 13323 7615 13365 7624
rect 13227 6824 13269 6833
rect 13227 6784 13228 6824
rect 13268 6784 13269 6824
rect 13227 6775 13269 6784
rect 13036 6581 13076 6666
rect 13035 6572 13077 6581
rect 13035 6532 13036 6572
rect 13076 6532 13077 6572
rect 13035 6523 13077 6532
rect 13228 6488 13268 6497
rect 12892 6446 12932 6455
rect 12892 6404 12932 6406
rect 12892 6364 13172 6404
rect 13132 5900 13172 6364
rect 13132 5851 13172 5860
rect 12940 5657 12980 5742
rect 12939 5648 12981 5657
rect 12939 5608 12940 5648
rect 12980 5608 12981 5648
rect 12939 5599 12981 5608
rect 13228 5480 13268 6448
rect 13420 5657 13460 8287
rect 13419 5648 13461 5657
rect 13419 5608 13420 5648
rect 13460 5608 13461 5648
rect 13419 5599 13461 5608
rect 13516 5480 13556 10471
rect 13611 9092 13653 9101
rect 13611 9052 13612 9092
rect 13652 9052 13653 9092
rect 13611 9043 13653 9052
rect 12940 5440 13268 5480
rect 13438 5440 13556 5480
rect 13612 8000 13652 9043
rect 12940 4985 12980 5440
rect 13438 5396 13478 5440
rect 13420 5356 13478 5396
rect 13036 5060 13076 5069
rect 13076 5020 13172 5060
rect 13036 5011 13076 5020
rect 12747 4976 12789 4985
rect 12844 4976 12884 4985
rect 12747 4936 12748 4976
rect 12788 4936 12844 4976
rect 12747 4927 12789 4936
rect 12844 4927 12884 4936
rect 12939 4976 12981 4985
rect 12939 4936 12940 4976
rect 12980 4936 12981 4976
rect 13132 4976 13172 5020
rect 13420 4976 13460 5356
rect 13515 5312 13557 5321
rect 13515 5272 13516 5312
rect 13556 5272 13557 5312
rect 13515 5263 13557 5272
rect 13132 4957 13364 4976
rect 13132 4936 13324 4957
rect 12939 4927 12981 4936
rect 12748 4145 12788 4927
rect 13324 4908 13364 4917
rect 12747 4136 12789 4145
rect 12747 4096 12748 4136
rect 12788 4096 12789 4136
rect 12747 4087 12789 4096
rect 13228 4136 13268 4145
rect 12748 2717 12788 4087
rect 13228 3977 13268 4096
rect 13227 3968 13269 3977
rect 13227 3928 13228 3968
rect 13268 3928 13269 3968
rect 13227 3919 13269 3928
rect 12940 3676 13364 3716
rect 12940 3464 12980 3676
rect 12892 3454 12980 3464
rect 12932 3424 12980 3454
rect 13036 3548 13076 3557
rect 12892 3405 12932 3414
rect 12747 2708 12789 2717
rect 12747 2668 12748 2708
rect 12788 2668 12789 2708
rect 12747 2659 12789 2668
rect 13036 2540 13076 3508
rect 13324 2876 13364 3676
rect 13420 3221 13460 4936
rect 13516 3464 13556 5263
rect 13516 3415 13556 3424
rect 13419 3212 13461 3221
rect 13419 3172 13420 3212
rect 13460 3172 13461 3212
rect 13419 3163 13461 3172
rect 13324 2827 13364 2836
rect 13131 2708 13173 2717
rect 13131 2668 13132 2708
rect 13172 2668 13173 2708
rect 13131 2659 13173 2668
rect 13132 2624 13172 2659
rect 13132 2573 13172 2584
rect 12748 2500 13076 2540
rect 12748 2129 12788 2500
rect 13516 2456 13556 2465
rect 12940 2416 13516 2456
rect 12747 2120 12789 2129
rect 12747 2080 12748 2120
rect 12788 2080 12789 2120
rect 12747 2071 12789 2080
rect 11404 1700 11444 1709
rect 11788 1700 11828 1709
rect 12076 1700 12116 1709
rect 11444 1660 11540 1700
rect 11404 1651 11444 1660
rect 11211 1196 11253 1205
rect 11211 1156 11212 1196
rect 11252 1156 11253 1196
rect 11211 1147 11253 1156
rect 11212 1062 11252 1147
rect 11307 1112 11349 1121
rect 11307 1072 11308 1112
rect 11348 1072 11349 1112
rect 11307 1063 11349 1072
rect 11020 944 11060 953
rect 10923 860 10965 869
rect 10923 820 10924 860
rect 10964 820 10965 860
rect 10923 811 10965 820
rect 10636 568 10772 608
rect 10636 80 10676 568
rect 11020 533 11060 904
rect 11211 944 11253 953
rect 11211 904 11212 944
rect 11252 904 11253 944
rect 11211 895 11253 904
rect 10827 524 10869 533
rect 10827 484 10828 524
rect 10868 484 10869 524
rect 10827 475 10869 484
rect 11019 524 11061 533
rect 11019 484 11020 524
rect 11060 484 11061 524
rect 11019 475 11061 484
rect 10828 80 10868 475
rect 11019 356 11061 365
rect 11019 316 11020 356
rect 11060 316 11061 356
rect 11019 307 11061 316
rect 11020 80 11060 307
rect 11212 80 11252 895
rect 11308 692 11348 1063
rect 11403 944 11445 953
rect 11403 904 11404 944
rect 11444 904 11445 944
rect 11403 895 11445 904
rect 11404 810 11444 895
rect 11500 869 11540 1660
rect 11828 1660 12020 1700
rect 11788 1651 11828 1660
rect 11787 1280 11829 1289
rect 11787 1240 11788 1280
rect 11828 1240 11829 1280
rect 11787 1231 11829 1240
rect 11499 860 11541 869
rect 11499 820 11500 860
rect 11540 820 11541 860
rect 11499 811 11541 820
rect 11308 652 11444 692
rect 11404 80 11444 652
rect 11595 524 11637 533
rect 11595 484 11596 524
rect 11636 484 11637 524
rect 11595 475 11637 484
rect 11596 80 11636 475
rect 11788 80 11828 1231
rect 11980 1112 12020 1660
rect 12076 1373 12116 1660
rect 12651 1700 12693 1709
rect 12651 1660 12652 1700
rect 12692 1660 12693 1700
rect 12651 1651 12693 1660
rect 12075 1364 12117 1373
rect 12075 1324 12076 1364
rect 12116 1324 12117 1364
rect 12075 1315 12117 1324
rect 12651 1196 12693 1205
rect 12651 1156 12652 1196
rect 12692 1156 12693 1196
rect 12651 1147 12693 1156
rect 11980 1072 12404 1112
rect 11979 944 12021 953
rect 11979 904 11980 944
rect 12020 904 12021 944
rect 11979 895 12021 904
rect 11980 80 12020 895
rect 12171 860 12213 869
rect 12171 820 12172 860
rect 12212 820 12213 860
rect 12171 811 12213 820
rect 12172 80 12212 811
rect 12364 80 12404 1072
rect 12652 1062 12692 1147
rect 12460 944 12500 953
rect 12460 449 12500 904
rect 12555 944 12597 953
rect 12555 904 12556 944
rect 12596 904 12597 944
rect 12555 895 12597 904
rect 12844 944 12884 953
rect 12459 440 12501 449
rect 12459 400 12460 440
rect 12500 400 12501 440
rect 12459 391 12501 400
rect 12556 80 12596 895
rect 12844 617 12884 904
rect 12843 608 12885 617
rect 12843 568 12844 608
rect 12884 568 12885 608
rect 12843 559 12885 568
rect 12747 524 12789 533
rect 12747 484 12748 524
rect 12788 484 12789 524
rect 12747 475 12789 484
rect 12748 80 12788 475
rect 12940 80 12980 2416
rect 13516 2407 13556 2416
rect 13323 2204 13365 2213
rect 13323 2164 13324 2204
rect 13364 2164 13365 2204
rect 13323 2155 13365 2164
rect 13035 1196 13077 1205
rect 13035 1156 13036 1196
rect 13076 1156 13077 1196
rect 13035 1147 13077 1156
rect 13036 1062 13076 1147
rect 13227 944 13269 953
rect 13227 904 13228 944
rect 13268 904 13269 944
rect 13227 895 13269 904
rect 13228 810 13268 895
rect 13131 440 13173 449
rect 13131 400 13132 440
rect 13172 400 13173 440
rect 13131 391 13173 400
rect 13132 80 13172 391
rect 13324 80 13364 2155
rect 13612 1961 13652 7960
rect 13708 4985 13748 11320
rect 13804 10613 13844 13999
rect 13899 11696 13941 11705
rect 13899 11656 13900 11696
rect 13940 11656 13941 11696
rect 13899 11647 13941 11656
rect 13900 11033 13940 11647
rect 13899 11024 13941 11033
rect 13899 10984 13900 11024
rect 13940 10984 13941 11024
rect 13899 10975 13941 10984
rect 13803 10604 13845 10613
rect 13803 10564 13804 10604
rect 13844 10564 13845 10604
rect 13803 10555 13845 10564
rect 13803 10436 13845 10445
rect 13803 10396 13804 10436
rect 13844 10396 13845 10436
rect 13803 10387 13845 10396
rect 13707 4976 13749 4985
rect 13707 4936 13708 4976
rect 13748 4936 13749 4976
rect 13707 4927 13749 4936
rect 13804 4976 13844 10387
rect 13900 10193 13940 10975
rect 13899 10184 13941 10193
rect 13899 10144 13900 10184
rect 13940 10144 13941 10184
rect 13899 10135 13941 10144
rect 13900 6992 13940 7001
rect 13900 5741 13940 6952
rect 13899 5732 13941 5741
rect 13899 5692 13900 5732
rect 13940 5692 13941 5732
rect 13899 5683 13941 5692
rect 13804 4927 13844 4936
rect 13996 5648 14036 18712
rect 14092 18593 14132 19216
rect 14188 18929 14228 19888
rect 14284 19349 14324 19972
rect 14380 19844 14420 19853
rect 14380 19685 14420 19804
rect 14379 19676 14421 19685
rect 14379 19636 14380 19676
rect 14420 19636 14421 19676
rect 14379 19627 14421 19636
rect 14476 19424 14516 22651
rect 14572 21617 14612 24247
rect 14668 23801 14708 23887
rect 14667 23797 14709 23801
rect 14667 23752 14668 23797
rect 14708 23752 14709 23797
rect 14956 23792 14996 24331
rect 15052 23960 15092 24760
rect 15339 24760 15340 24800
rect 15380 24760 15381 24800
rect 15339 24751 15381 24760
rect 15244 24632 15284 24641
rect 15052 23911 15092 23920
rect 15148 24592 15244 24632
rect 14956 23752 15092 23792
rect 14667 23743 14709 23752
rect 14859 23708 14901 23717
rect 14859 23668 14860 23708
rect 14900 23668 14901 23708
rect 14859 23659 14901 23668
rect 14860 23574 14900 23659
rect 14764 22289 14804 22294
rect 14763 22285 14805 22289
rect 14763 22240 14764 22285
rect 14804 22240 14805 22285
rect 14763 22231 14805 22240
rect 14571 21608 14613 21617
rect 14571 21568 14572 21608
rect 14612 21568 14613 21608
rect 14571 21559 14613 21568
rect 14764 21608 14804 22231
rect 14956 22112 14996 22121
rect 14956 21617 14996 22072
rect 14860 21608 14900 21617
rect 14764 21568 14860 21608
rect 14572 21474 14612 21559
rect 14667 21440 14709 21449
rect 14667 21400 14668 21440
rect 14708 21400 14709 21440
rect 14667 21391 14709 21400
rect 14571 21020 14613 21029
rect 14571 20980 14572 21020
rect 14612 20980 14613 21020
rect 14571 20971 14613 20980
rect 14572 20768 14612 20971
rect 14572 20719 14612 20728
rect 14380 19384 14516 19424
rect 14283 19340 14325 19349
rect 14283 19300 14284 19340
rect 14324 19300 14325 19340
rect 14283 19291 14325 19300
rect 14187 18920 14229 18929
rect 14187 18880 14188 18920
rect 14228 18880 14229 18920
rect 14187 18871 14229 18880
rect 14283 18836 14325 18845
rect 14283 18796 14284 18836
rect 14324 18796 14325 18836
rect 14283 18787 14325 18796
rect 14091 18584 14133 18593
rect 14091 18544 14092 18584
rect 14132 18544 14133 18584
rect 14091 18535 14133 18544
rect 14187 18500 14229 18509
rect 14187 18460 14188 18500
rect 14228 18460 14229 18500
rect 14187 18451 14229 18460
rect 14284 18500 14324 18787
rect 14380 18668 14420 19384
rect 14572 19265 14612 19350
rect 14476 19256 14516 19265
rect 14476 18845 14516 19216
rect 14571 19256 14613 19265
rect 14571 19216 14572 19256
rect 14612 19216 14613 19256
rect 14571 19207 14613 19216
rect 14668 19088 14708 21391
rect 14764 21020 14804 21568
rect 14860 21559 14900 21568
rect 14955 21608 14997 21617
rect 14955 21568 14956 21608
rect 14996 21568 14997 21608
rect 14955 21559 14997 21568
rect 14764 20971 14804 20980
rect 14860 21356 14900 21365
rect 14763 20600 14805 20609
rect 14763 20560 14764 20600
rect 14804 20560 14805 20600
rect 14763 20551 14805 20560
rect 14764 20466 14804 20551
rect 14763 20348 14805 20357
rect 14763 20308 14764 20348
rect 14804 20308 14805 20348
rect 14860 20348 14900 21316
rect 14955 21188 14997 21197
rect 14955 21148 14956 21188
rect 14996 21148 14997 21188
rect 14955 21139 14997 21148
rect 14956 21020 14996 21139
rect 14956 20971 14996 20980
rect 15052 20357 15092 23752
rect 15148 23372 15188 24592
rect 15244 24583 15284 24592
rect 15340 24128 15380 24751
rect 15244 24088 15380 24128
rect 15244 23885 15284 24088
rect 15436 24044 15476 25675
rect 15532 25556 15572 26524
rect 15819 26480 15861 26489
rect 15819 26440 15820 26480
rect 15860 26440 15861 26480
rect 15819 26431 15861 26440
rect 15723 26312 15765 26321
rect 15723 26272 15724 26312
rect 15764 26272 15765 26312
rect 15723 26263 15765 26272
rect 15724 26178 15764 26263
rect 15532 25507 15572 25516
rect 15628 26144 15668 26153
rect 15628 26060 15668 26104
rect 15820 26060 15860 26431
rect 15916 26144 15956 26153
rect 16012 26144 16052 30379
rect 16204 28925 16244 37360
rect 16396 36989 16436 37519
rect 16395 36980 16437 36989
rect 16395 36940 16396 36980
rect 16436 36940 16437 36980
rect 16395 36931 16437 36940
rect 16396 36728 16436 36931
rect 16396 36679 16436 36688
rect 16395 36560 16437 36569
rect 16395 36520 16396 36560
rect 16436 36520 16437 36560
rect 16395 36511 16437 36520
rect 16396 35888 16436 36511
rect 16492 36485 16532 38872
rect 16684 38417 16724 39712
rect 16876 39257 16916 41140
rect 16972 41131 17012 41140
rect 17356 41140 17452 41180
rect 16971 40676 17013 40685
rect 16971 40636 16972 40676
rect 17012 40636 17013 40676
rect 16971 40627 17013 40636
rect 16972 40542 17012 40627
rect 17164 40508 17204 40517
rect 17068 40468 17164 40508
rect 16971 39752 17013 39761
rect 16971 39712 16972 39752
rect 17012 39712 17013 39752
rect 16971 39703 17013 39712
rect 16972 39618 17012 39703
rect 16972 39500 17012 39509
rect 16875 39248 16917 39257
rect 16875 39208 16876 39248
rect 16916 39208 16917 39248
rect 16875 39199 16917 39208
rect 16972 39005 17012 39460
rect 16971 38996 17013 39005
rect 16971 38956 16972 38996
rect 17012 38956 17013 38996
rect 16971 38947 17013 38956
rect 17068 38921 17108 40468
rect 17164 40459 17204 40468
rect 17356 39836 17396 41140
rect 17452 41131 17492 41140
rect 17548 40685 17588 42928
rect 17740 41432 17780 42928
rect 17836 41432 17876 41441
rect 17740 41392 17836 41432
rect 17836 41383 17876 41392
rect 17643 41180 17685 41189
rect 17643 41140 17644 41180
rect 17684 41140 17685 41180
rect 17643 41131 17685 41140
rect 17547 40676 17589 40685
rect 17547 40636 17548 40676
rect 17588 40636 17589 40676
rect 17547 40627 17589 40636
rect 17547 40340 17589 40349
rect 17547 40300 17548 40340
rect 17588 40300 17589 40340
rect 17547 40291 17589 40300
rect 17548 40206 17588 40291
rect 17644 39929 17684 41131
rect 17739 40844 17781 40853
rect 17739 40804 17740 40844
rect 17780 40804 17781 40844
rect 17739 40795 17781 40804
rect 17740 40508 17780 40795
rect 17932 40769 17972 42928
rect 18124 41432 18164 42928
rect 18316 41525 18356 42928
rect 18315 41516 18357 41525
rect 18315 41476 18316 41516
rect 18356 41476 18357 41516
rect 18315 41467 18357 41476
rect 18124 41383 18164 41392
rect 18508 41348 18548 42928
rect 18700 41600 18740 42928
rect 18892 41693 18932 42928
rect 18891 41684 18933 41693
rect 18891 41644 18892 41684
rect 18932 41644 18933 41684
rect 18891 41635 18933 41644
rect 18412 41308 18548 41348
rect 18604 41560 18740 41600
rect 18795 41600 18837 41609
rect 18795 41560 18796 41600
rect 18836 41560 18837 41600
rect 18027 41180 18069 41189
rect 18316 41180 18356 41189
rect 18027 41140 18028 41180
rect 18068 41140 18069 41180
rect 18027 41131 18069 41140
rect 18220 41140 18316 41180
rect 17931 40760 17973 40769
rect 17931 40720 17932 40760
rect 17972 40720 17973 40760
rect 17931 40711 17973 40720
rect 17740 40459 17780 40468
rect 17932 40592 17972 40601
rect 17932 40433 17972 40552
rect 17931 40424 17973 40433
rect 17931 40384 17932 40424
rect 17972 40384 17973 40424
rect 17931 40375 17973 40384
rect 17643 39920 17685 39929
rect 17643 39880 17644 39920
rect 17684 39880 17685 39920
rect 17643 39871 17685 39880
rect 17356 39796 17492 39836
rect 17164 39752 17204 39761
rect 17164 39089 17204 39712
rect 17260 39752 17300 39761
rect 17300 39712 17396 39752
rect 17260 39703 17300 39712
rect 17163 39080 17205 39089
rect 17163 39040 17164 39080
rect 17204 39040 17205 39080
rect 17163 39031 17205 39040
rect 17067 38912 17109 38921
rect 17067 38872 17068 38912
rect 17108 38872 17109 38912
rect 17067 38863 17109 38872
rect 16683 38408 16725 38417
rect 16683 38368 16684 38408
rect 16724 38368 16725 38408
rect 16683 38359 16725 38368
rect 16588 38240 16628 38249
rect 16588 38081 16628 38200
rect 16683 38240 16725 38249
rect 16683 38200 16684 38240
rect 16724 38200 16725 38240
rect 16683 38191 16725 38200
rect 17259 38240 17301 38249
rect 17259 38200 17260 38240
rect 17300 38200 17301 38240
rect 17259 38191 17301 38200
rect 16684 38106 16724 38191
rect 17068 38156 17108 38165
rect 16780 38116 17068 38156
rect 16587 38072 16629 38081
rect 16587 38032 16588 38072
rect 16628 38032 16629 38072
rect 16587 38023 16629 38032
rect 16683 37736 16725 37745
rect 16683 37696 16684 37736
rect 16724 37696 16725 37736
rect 16683 37687 16725 37696
rect 16587 37400 16629 37409
rect 16587 37360 16588 37400
rect 16628 37360 16629 37400
rect 16587 37351 16629 37360
rect 16588 36896 16628 37351
rect 16588 36847 16628 36856
rect 16587 36644 16629 36653
rect 16684 36644 16724 37687
rect 16587 36604 16588 36644
rect 16628 36604 16724 36644
rect 16587 36595 16629 36604
rect 16491 36476 16533 36485
rect 16491 36436 16492 36476
rect 16532 36436 16533 36476
rect 16491 36427 16533 36436
rect 16396 34544 16436 35848
rect 16491 35300 16533 35309
rect 16491 35260 16492 35300
rect 16532 35260 16533 35300
rect 16491 35251 16533 35260
rect 16492 35216 16532 35251
rect 16492 35165 16532 35176
rect 16588 35141 16628 36595
rect 16780 35813 16820 38116
rect 17068 38107 17108 38116
rect 17163 38156 17205 38165
rect 17163 38116 17164 38156
rect 17204 38116 17205 38156
rect 17163 38107 17205 38116
rect 17164 38022 17204 38107
rect 16875 37988 16917 37997
rect 16875 37948 16876 37988
rect 16916 37948 16917 37988
rect 16875 37939 16917 37948
rect 16876 36149 16916 37939
rect 17163 37736 17205 37745
rect 17163 37696 17164 37736
rect 17204 37696 17205 37736
rect 17163 37687 17205 37696
rect 17164 37325 17204 37687
rect 17163 37316 17205 37325
rect 17163 37276 17164 37316
rect 17204 37276 17205 37316
rect 17163 37267 17205 37276
rect 16972 36644 17012 36653
rect 16972 36485 17012 36604
rect 17163 36560 17205 36569
rect 17163 36520 17164 36560
rect 17204 36520 17205 36560
rect 17163 36511 17205 36520
rect 16971 36476 17013 36485
rect 16971 36436 16972 36476
rect 17012 36436 17013 36476
rect 16971 36427 17013 36436
rect 17164 36426 17204 36511
rect 17067 36392 17109 36401
rect 17067 36352 17068 36392
rect 17108 36352 17109 36392
rect 17067 36343 17109 36352
rect 16875 36140 16917 36149
rect 16875 36100 16876 36140
rect 16916 36100 16917 36140
rect 16875 36091 16917 36100
rect 16924 35897 16964 35906
rect 16964 35857 17012 35888
rect 16924 35848 17012 35857
rect 16779 35804 16821 35813
rect 16779 35764 16780 35804
rect 16820 35764 16821 35804
rect 16779 35755 16821 35764
rect 16875 35720 16917 35729
rect 16875 35680 16876 35720
rect 16916 35680 16917 35720
rect 16875 35671 16917 35680
rect 16683 35552 16725 35561
rect 16683 35512 16684 35552
rect 16724 35512 16725 35552
rect 16683 35503 16725 35512
rect 16587 35132 16629 35141
rect 16587 35092 16588 35132
rect 16628 35092 16629 35132
rect 16587 35083 16629 35092
rect 16396 34504 16532 34544
rect 16395 33872 16437 33881
rect 16395 33832 16396 33872
rect 16436 33832 16437 33872
rect 16395 33823 16437 33832
rect 16299 32864 16341 32873
rect 16299 32824 16300 32864
rect 16340 32824 16341 32864
rect 16299 32815 16341 32824
rect 16396 32864 16436 33823
rect 16300 32730 16340 32815
rect 16396 32612 16436 32824
rect 16492 32705 16532 34504
rect 16491 32696 16533 32705
rect 16491 32656 16492 32696
rect 16532 32656 16533 32696
rect 16491 32647 16533 32656
rect 16300 32572 16436 32612
rect 16300 30680 16340 32572
rect 16588 32528 16628 35083
rect 16684 34376 16724 35503
rect 16780 34376 16820 34385
rect 16684 34336 16780 34376
rect 16780 34327 16820 34336
rect 16876 33965 16916 35671
rect 16972 35202 17012 35848
rect 17068 35804 17108 36343
rect 17260 36308 17300 38191
rect 17356 37241 17396 39712
rect 17452 37997 17492 39796
rect 17548 39752 17588 39761
rect 17548 39089 17588 39712
rect 17644 39752 17684 39761
rect 17547 39080 17589 39089
rect 17547 39040 17548 39080
rect 17588 39040 17589 39080
rect 17644 39080 17684 39712
rect 17740 39752 17780 39761
rect 17780 39712 17876 39752
rect 17740 39703 17780 39712
rect 17739 39080 17781 39089
rect 17644 39040 17740 39080
rect 17780 39040 17781 39080
rect 17547 39031 17589 39040
rect 17739 39031 17781 39040
rect 17548 38585 17588 39031
rect 17739 38912 17781 38921
rect 17644 38872 17740 38912
rect 17780 38872 17781 38912
rect 17547 38576 17589 38585
rect 17547 38536 17548 38576
rect 17588 38536 17589 38576
rect 17547 38527 17589 38536
rect 17644 38408 17684 38872
rect 17739 38863 17781 38872
rect 17740 38778 17780 38863
rect 17836 38669 17876 39712
rect 17932 39500 17972 39509
rect 17932 38921 17972 39460
rect 17931 38912 17973 38921
rect 17931 38872 17932 38912
rect 17972 38872 17973 38912
rect 17931 38863 17973 38872
rect 17932 38744 17972 38753
rect 17835 38660 17877 38669
rect 17835 38620 17836 38660
rect 17876 38620 17877 38660
rect 17835 38611 17877 38620
rect 17548 38368 17684 38408
rect 17451 37988 17493 37997
rect 17451 37948 17452 37988
rect 17492 37948 17493 37988
rect 17451 37939 17493 37948
rect 17451 37820 17493 37829
rect 17451 37780 17452 37820
rect 17492 37780 17493 37820
rect 17451 37771 17493 37780
rect 17452 37568 17492 37771
rect 17548 37745 17588 38368
rect 17644 38240 17684 38249
rect 17684 38200 17780 38240
rect 17644 38191 17684 38200
rect 17643 38072 17685 38081
rect 17643 38032 17644 38072
rect 17684 38032 17685 38072
rect 17643 38023 17685 38032
rect 17547 37736 17589 37745
rect 17547 37696 17548 37736
rect 17588 37696 17589 37736
rect 17547 37687 17589 37696
rect 17644 37652 17684 38023
rect 17644 37603 17684 37612
rect 17452 37528 17588 37568
rect 17452 37400 17492 37409
rect 17452 37325 17492 37360
rect 17451 37316 17493 37325
rect 17451 37276 17452 37316
rect 17492 37276 17493 37316
rect 17451 37267 17493 37276
rect 17452 37265 17492 37267
rect 17355 37232 17397 37241
rect 17355 37192 17356 37232
rect 17396 37192 17397 37232
rect 17355 37183 17397 37192
rect 17356 36728 17396 36739
rect 17356 36653 17396 36688
rect 17451 36728 17493 36737
rect 17451 36688 17452 36728
rect 17492 36688 17493 36728
rect 17451 36679 17493 36688
rect 17355 36644 17397 36653
rect 17355 36604 17356 36644
rect 17396 36604 17397 36644
rect 17355 36595 17397 36604
rect 17452 36594 17492 36679
rect 17068 35755 17108 35764
rect 17164 36268 17300 36308
rect 17067 35384 17109 35393
rect 17067 35344 17068 35384
rect 17108 35344 17109 35384
rect 17067 35335 17109 35344
rect 16972 34628 17012 35162
rect 16972 34579 17012 34588
rect 16971 34208 17013 34217
rect 16971 34168 16972 34208
rect 17012 34168 17013 34208
rect 16971 34159 17013 34168
rect 16683 33956 16725 33965
rect 16683 33916 16684 33956
rect 16724 33916 16725 33956
rect 16683 33907 16725 33916
rect 16875 33956 16917 33965
rect 16875 33916 16876 33956
rect 16916 33916 16917 33956
rect 16875 33907 16917 33916
rect 16684 33704 16724 33907
rect 16875 33788 16917 33797
rect 16875 33748 16876 33788
rect 16916 33748 16917 33788
rect 16875 33739 16917 33748
rect 16684 33629 16724 33664
rect 16876 33654 16916 33739
rect 16683 33620 16725 33629
rect 16683 33580 16684 33620
rect 16724 33580 16725 33620
rect 16683 33571 16725 33580
rect 16972 33032 17012 34159
rect 16396 32488 16628 32528
rect 16780 32992 17012 33032
rect 16396 32117 16436 32488
rect 16395 32108 16437 32117
rect 16395 32068 16396 32108
rect 16436 32068 16437 32108
rect 16395 32059 16437 32068
rect 16492 32108 16532 32117
rect 16492 32024 16532 32068
rect 16780 32024 16820 32992
rect 16876 32864 16916 32873
rect 16876 32705 16916 32824
rect 16971 32780 17013 32789
rect 16971 32740 16972 32780
rect 17012 32740 17013 32780
rect 16971 32731 17013 32740
rect 16875 32696 16917 32705
rect 16875 32656 16876 32696
rect 16916 32656 16917 32696
rect 16875 32647 16917 32656
rect 16492 31984 16820 32024
rect 16395 31940 16437 31949
rect 16395 31900 16396 31940
rect 16436 31900 16437 31940
rect 16395 31891 16437 31900
rect 16300 30631 16340 30640
rect 16299 30512 16341 30521
rect 16299 30472 16300 30512
rect 16340 30472 16341 30512
rect 16396 30512 16436 31891
rect 16683 31436 16725 31445
rect 16683 31396 16684 31436
rect 16724 31396 16725 31436
rect 16683 31387 16725 31396
rect 16491 31352 16533 31361
rect 16491 31312 16492 31352
rect 16532 31312 16533 31352
rect 16491 31303 16533 31312
rect 16492 30848 16532 31303
rect 16684 31193 16724 31387
rect 16683 31184 16725 31193
rect 16683 31144 16684 31184
rect 16724 31144 16725 31184
rect 16683 31135 16725 31144
rect 16492 30799 16532 30808
rect 16588 30689 16628 30774
rect 16587 30680 16629 30689
rect 16587 30640 16588 30680
rect 16628 30640 16629 30680
rect 16587 30631 16629 30640
rect 16396 30472 16724 30512
rect 16299 30463 16341 30472
rect 16203 28916 16245 28925
rect 16203 28876 16204 28916
rect 16244 28876 16245 28916
rect 16203 28867 16245 28876
rect 16107 28580 16149 28589
rect 16107 28540 16108 28580
rect 16148 28540 16149 28580
rect 16107 28531 16149 28540
rect 16108 28446 16148 28531
rect 16107 27656 16149 27665
rect 16107 27616 16108 27656
rect 16148 27616 16149 27656
rect 16107 27607 16149 27616
rect 16108 26984 16148 27607
rect 16203 27236 16245 27245
rect 16203 27196 16204 27236
rect 16244 27196 16245 27236
rect 16203 27187 16245 27196
rect 16108 26935 16148 26944
rect 15956 26104 16052 26144
rect 16108 26816 16148 26825
rect 15916 26095 15956 26104
rect 15628 26020 15860 26060
rect 15628 25388 15668 26020
rect 15723 25892 15765 25901
rect 15723 25852 15724 25892
rect 15764 25852 15765 25892
rect 15723 25843 15765 25852
rect 15532 25348 15668 25388
rect 15532 25304 15572 25348
rect 15532 25255 15572 25264
rect 15627 25136 15669 25145
rect 15627 25096 15628 25136
rect 15668 25096 15669 25136
rect 15627 25087 15669 25096
rect 15628 24716 15668 25087
rect 15628 24667 15668 24676
rect 15340 24004 15476 24044
rect 15532 24632 15572 24641
rect 15243 23876 15285 23885
rect 15243 23836 15244 23876
rect 15284 23836 15285 23876
rect 15243 23827 15285 23836
rect 15244 23792 15284 23827
rect 15244 23742 15284 23752
rect 15340 23792 15380 24004
rect 15340 23456 15380 23752
rect 15435 23792 15477 23801
rect 15435 23752 15436 23792
rect 15476 23752 15477 23792
rect 15435 23743 15477 23752
rect 15436 23658 15476 23743
rect 15532 23717 15572 24592
rect 15724 24548 15764 25843
rect 15819 25556 15861 25565
rect 15819 25516 15820 25556
rect 15860 25516 15861 25556
rect 15819 25507 15861 25516
rect 15628 24508 15764 24548
rect 15531 23708 15573 23717
rect 15531 23668 15532 23708
rect 15572 23668 15573 23708
rect 15531 23659 15573 23668
rect 15340 23416 15476 23456
rect 15148 23332 15380 23372
rect 15340 23288 15380 23332
rect 15340 23239 15380 23248
rect 15243 23120 15285 23129
rect 15148 23099 15244 23120
rect 15188 23080 15244 23099
rect 15284 23080 15285 23120
rect 15243 23071 15285 23080
rect 15148 23050 15188 23059
rect 15436 23036 15476 23416
rect 15340 22996 15476 23036
rect 15147 22784 15189 22793
rect 15147 22744 15148 22784
rect 15188 22744 15189 22784
rect 15147 22735 15189 22744
rect 15148 22028 15188 22735
rect 15340 22373 15380 22996
rect 15628 22793 15668 24508
rect 15723 23792 15765 23801
rect 15723 23752 15724 23792
rect 15764 23752 15765 23792
rect 15723 23743 15765 23752
rect 15724 23658 15764 23743
rect 15724 23120 15764 23129
rect 15820 23120 15860 25507
rect 16011 24548 16053 24557
rect 16108 24548 16148 26776
rect 16204 26237 16244 27187
rect 16300 26489 16340 30463
rect 16395 30344 16437 30353
rect 16395 30304 16396 30344
rect 16436 30304 16437 30344
rect 16395 30295 16437 30304
rect 16396 27236 16436 30295
rect 16588 29168 16628 29177
rect 16588 29009 16628 29128
rect 16587 29000 16629 29009
rect 16587 28960 16588 29000
rect 16628 28960 16629 29000
rect 16684 29000 16724 30472
rect 16780 29261 16820 31984
rect 16876 31949 16916 32647
rect 16972 32192 17012 32731
rect 16875 31940 16917 31949
rect 16875 31900 16876 31940
rect 16916 31900 16917 31940
rect 16875 31891 16917 31900
rect 16972 31772 17012 32152
rect 16876 31732 17012 31772
rect 16876 31445 16916 31732
rect 16875 31436 16917 31445
rect 16875 31396 16876 31436
rect 16916 31396 16917 31436
rect 16875 31387 16917 31396
rect 16875 31268 16917 31277
rect 17068 31268 17108 35335
rect 17164 35300 17204 36268
rect 17355 36140 17397 36149
rect 17355 36100 17356 36140
rect 17396 36100 17397 36140
rect 17355 36091 17397 36100
rect 17452 36140 17492 36149
rect 17548 36140 17588 37528
rect 17740 36989 17780 38200
rect 17836 38081 17876 38611
rect 17932 38585 17972 38704
rect 17931 38576 17973 38585
rect 17931 38536 17932 38576
rect 17972 38536 17973 38576
rect 17931 38527 17973 38536
rect 17931 38324 17973 38333
rect 17931 38284 17932 38324
rect 17972 38284 17973 38324
rect 17931 38275 17973 38284
rect 17835 38072 17877 38081
rect 17835 38032 17836 38072
rect 17876 38032 17877 38072
rect 17835 38023 17877 38032
rect 17835 37064 17877 37073
rect 17835 37024 17836 37064
rect 17876 37024 17877 37064
rect 17835 37015 17877 37024
rect 17739 36980 17781 36989
rect 17739 36940 17740 36980
rect 17780 36940 17781 36980
rect 17739 36931 17781 36940
rect 17644 36728 17684 36737
rect 17684 36688 17780 36728
rect 17644 36679 17684 36688
rect 17643 36560 17685 36569
rect 17643 36520 17644 36560
rect 17684 36520 17685 36560
rect 17643 36511 17685 36520
rect 17644 36426 17684 36511
rect 17492 36100 17588 36140
rect 17452 36091 17492 36100
rect 17164 35251 17204 35260
rect 17260 35972 17300 35981
rect 17163 33788 17205 33797
rect 17163 33748 17164 33788
rect 17204 33748 17205 33788
rect 17163 33739 17205 33748
rect 17164 33704 17204 33739
rect 17164 33653 17204 33664
rect 17260 33461 17300 35932
rect 17356 34460 17396 36091
rect 17644 35972 17684 35981
rect 17547 35132 17589 35141
rect 17547 35092 17548 35132
rect 17588 35092 17589 35132
rect 17547 35083 17589 35092
rect 17452 34460 17492 34469
rect 17356 34420 17452 34460
rect 17452 34411 17492 34420
rect 17548 34292 17588 35083
rect 17644 35057 17684 35932
rect 17643 35048 17685 35057
rect 17643 35008 17644 35048
rect 17684 35008 17685 35048
rect 17643 34999 17685 35008
rect 17644 34914 17684 34999
rect 17643 34544 17685 34553
rect 17643 34504 17644 34544
rect 17684 34504 17685 34544
rect 17643 34495 17685 34504
rect 17644 34410 17684 34495
rect 17356 34252 17588 34292
rect 17259 33452 17301 33461
rect 17259 33412 17260 33452
rect 17300 33412 17301 33452
rect 17259 33403 17301 33412
rect 17356 33284 17396 34252
rect 17740 34208 17780 36688
rect 17836 36140 17876 37015
rect 17932 36392 17972 38275
rect 18028 36728 18068 41131
rect 18123 40676 18165 40685
rect 18123 40636 18124 40676
rect 18164 40636 18165 40676
rect 18123 40627 18165 40636
rect 18124 40542 18164 40627
rect 18220 40349 18260 41140
rect 18316 41131 18356 41140
rect 18316 40508 18356 40517
rect 18219 40340 18261 40349
rect 18219 40300 18220 40340
rect 18260 40300 18261 40340
rect 18219 40291 18261 40300
rect 18316 40088 18356 40468
rect 18124 40048 18356 40088
rect 18124 38753 18164 40048
rect 18315 39920 18357 39929
rect 18315 39880 18316 39920
rect 18356 39880 18357 39920
rect 18412 39920 18452 41308
rect 18507 41180 18549 41189
rect 18507 41140 18508 41180
rect 18548 41140 18549 41180
rect 18507 41131 18549 41140
rect 18508 41046 18548 41131
rect 18507 40760 18549 40769
rect 18507 40720 18508 40760
rect 18548 40720 18549 40760
rect 18507 40711 18549 40720
rect 18508 40676 18548 40711
rect 18508 40625 18548 40636
rect 18508 39920 18548 39929
rect 18412 39880 18508 39920
rect 18315 39871 18357 39880
rect 18508 39871 18548 39880
rect 18316 39786 18356 39871
rect 18604 39752 18644 41560
rect 18795 41551 18837 41560
rect 18699 41432 18741 41441
rect 18699 41392 18700 41432
rect 18740 41392 18741 41432
rect 18699 41383 18741 41392
rect 18700 41298 18740 41383
rect 18796 41264 18836 41551
rect 19084 41432 19124 42928
rect 19276 42113 19316 42928
rect 19275 42104 19317 42113
rect 19275 42064 19276 42104
rect 19316 42064 19317 42104
rect 19275 42055 19317 42064
rect 19275 41684 19317 41693
rect 19275 41644 19276 41684
rect 19316 41644 19317 41684
rect 19275 41635 19317 41644
rect 18988 41392 19124 41432
rect 18796 41224 18932 41264
rect 18892 41096 18932 41224
rect 18892 41047 18932 41056
rect 18988 41021 19028 41392
rect 19083 41180 19125 41189
rect 19083 41140 19084 41180
rect 19124 41140 19125 41180
rect 19083 41131 19125 41140
rect 19084 41046 19124 41131
rect 18699 41012 18741 41021
rect 18699 40972 18700 41012
rect 18740 40972 18741 41012
rect 18699 40963 18741 40972
rect 18987 41012 19029 41021
rect 18987 40972 18988 41012
rect 19028 40972 19029 41012
rect 18987 40963 19029 40972
rect 18700 40676 18740 40963
rect 18808 40844 19176 40853
rect 18848 40804 18890 40844
rect 18930 40804 18972 40844
rect 19012 40804 19054 40844
rect 19094 40804 19136 40844
rect 18808 40795 19176 40804
rect 18891 40676 18933 40685
rect 19276 40676 19316 41635
rect 19468 41441 19508 42928
rect 20048 41600 20416 41609
rect 20088 41560 20130 41600
rect 20170 41560 20212 41600
rect 20252 41560 20294 41600
rect 20334 41560 20376 41600
rect 20048 41551 20416 41560
rect 19755 41516 19797 41525
rect 19755 41476 19756 41516
rect 19796 41476 19797 41516
rect 19755 41467 19797 41476
rect 19467 41432 19509 41441
rect 19467 41392 19468 41432
rect 19508 41392 19509 41432
rect 19467 41383 19509 41392
rect 19756 41432 19796 41467
rect 19756 41381 19796 41392
rect 19371 41348 19413 41357
rect 19371 41308 19372 41348
rect 19412 41308 19413 41348
rect 19371 41299 19413 41308
rect 19372 41180 19412 41299
rect 19372 41131 19412 41140
rect 19948 41180 19988 41189
rect 19564 41012 19604 41021
rect 19604 40972 19700 41012
rect 19564 40963 19604 40972
rect 19371 40928 19413 40937
rect 19371 40888 19372 40928
rect 19412 40888 19413 40928
rect 19371 40879 19413 40888
rect 18700 40636 18836 40676
rect 18700 40508 18740 40517
rect 18700 39929 18740 40468
rect 18699 39920 18741 39929
rect 18699 39880 18700 39920
rect 18740 39880 18741 39920
rect 18699 39871 18741 39880
rect 18412 39712 18644 39752
rect 18315 39668 18357 39677
rect 18315 39628 18316 39668
rect 18356 39628 18357 39668
rect 18315 39619 18357 39628
rect 18219 39584 18261 39593
rect 18219 39544 18220 39584
rect 18260 39544 18261 39584
rect 18219 39535 18261 39544
rect 18220 39450 18260 39535
rect 18316 39332 18356 39619
rect 18220 39292 18356 39332
rect 18123 38744 18165 38753
rect 18123 38704 18124 38744
rect 18164 38704 18165 38744
rect 18123 38695 18165 38704
rect 18123 38576 18165 38585
rect 18123 38536 18124 38576
rect 18164 38536 18165 38576
rect 18123 38527 18165 38536
rect 18124 38235 18164 38527
rect 18124 38186 18164 38195
rect 18220 37652 18260 39292
rect 18315 38324 18357 38333
rect 18315 38284 18316 38324
rect 18356 38284 18357 38324
rect 18315 38275 18357 38284
rect 18316 38190 18356 38275
rect 18316 37652 18356 37661
rect 18220 37612 18316 37652
rect 18316 37603 18356 37612
rect 18124 37484 18164 37493
rect 18124 36896 18164 37444
rect 18315 37232 18357 37241
rect 18315 37192 18316 37232
rect 18356 37192 18357 37232
rect 18315 37183 18357 37192
rect 18124 36847 18164 36856
rect 18316 36728 18356 37183
rect 18412 37073 18452 39712
rect 18796 39677 18836 40636
rect 18891 40636 18892 40676
rect 18932 40636 18933 40676
rect 18891 40627 18933 40636
rect 18988 40636 19316 40676
rect 18892 40542 18932 40627
rect 18892 39920 18932 39929
rect 18988 39920 19028 40636
rect 19084 40508 19124 40517
rect 19372 40508 19412 40879
rect 19563 40592 19605 40601
rect 19563 40552 19564 40592
rect 19604 40552 19605 40592
rect 19563 40543 19605 40552
rect 19124 40468 19220 40508
rect 19084 40459 19124 40468
rect 18932 39880 19028 39920
rect 18892 39871 18932 39880
rect 18700 39668 18740 39677
rect 18604 39080 18644 39089
rect 18700 39080 18740 39628
rect 18795 39668 18837 39677
rect 18795 39628 18796 39668
rect 18836 39628 18837 39668
rect 18795 39619 18837 39628
rect 19083 39668 19125 39677
rect 19083 39628 19084 39668
rect 19124 39628 19125 39668
rect 19083 39619 19125 39628
rect 19084 39534 19124 39619
rect 19180 39500 19220 40468
rect 19372 40459 19412 40468
rect 19564 40458 19604 40543
rect 19371 39836 19413 39845
rect 19371 39796 19372 39836
rect 19412 39796 19413 39836
rect 19371 39787 19413 39796
rect 19180 39460 19316 39500
rect 18808 39332 19176 39341
rect 18848 39292 18890 39332
rect 18930 39292 18972 39332
rect 19012 39292 19054 39332
rect 19094 39292 19136 39332
rect 18808 39283 19176 39292
rect 19276 39164 19316 39460
rect 18644 39040 18740 39080
rect 19180 39124 19316 39164
rect 18604 39031 18644 39040
rect 18891 38996 18933 39005
rect 18891 38956 18892 38996
rect 18932 38956 18933 38996
rect 18891 38947 18933 38956
rect 18796 38912 18836 38921
rect 18507 38744 18549 38753
rect 18507 38704 18508 38744
rect 18548 38704 18549 38744
rect 18507 38695 18549 38704
rect 18508 38610 18548 38695
rect 18796 38669 18836 38872
rect 18892 38912 18932 38947
rect 18892 38861 18932 38872
rect 18987 38912 19029 38921
rect 18987 38872 18988 38912
rect 19028 38872 19029 38912
rect 18987 38863 19029 38872
rect 18988 38778 19028 38863
rect 19084 38744 19124 38753
rect 18795 38660 18837 38669
rect 18795 38620 18796 38660
rect 18836 38620 18837 38660
rect 18795 38611 18837 38620
rect 18795 38324 18837 38333
rect 18988 38324 19028 38333
rect 19084 38324 19124 38704
rect 18795 38284 18796 38324
rect 18836 38284 18932 38324
rect 18795 38275 18837 38284
rect 18604 38240 18644 38249
rect 18507 37232 18549 37241
rect 18507 37192 18508 37232
rect 18548 37192 18549 37232
rect 18507 37183 18549 37192
rect 18508 37098 18548 37183
rect 18411 37064 18453 37073
rect 18411 37024 18412 37064
rect 18452 37024 18453 37064
rect 18411 37015 18453 37024
rect 18412 36896 18452 36905
rect 18604 36896 18644 38200
rect 18892 38240 18932 38284
rect 19028 38284 19124 38324
rect 18988 38275 19028 38284
rect 18892 38191 18932 38200
rect 19180 38081 19220 39124
rect 19372 39080 19412 39787
rect 19468 39668 19508 39677
rect 19660 39668 19700 40972
rect 19948 40517 19988 41140
rect 19852 40508 19892 40517
rect 19852 39761 19892 40468
rect 19947 40508 19989 40517
rect 19947 40468 19948 40508
rect 19988 40468 19989 40508
rect 19947 40459 19989 40468
rect 20523 40424 20565 40433
rect 20523 40384 20524 40424
rect 20564 40384 20565 40424
rect 20523 40375 20565 40384
rect 20044 40256 20084 40265
rect 19948 40216 20044 40256
rect 19851 39752 19893 39761
rect 19851 39712 19852 39752
rect 19892 39712 19893 39752
rect 19851 39703 19893 39712
rect 19660 39628 19796 39668
rect 19468 39425 19508 39628
rect 19756 39584 19796 39628
rect 19851 39584 19893 39593
rect 19756 39544 19852 39584
rect 19892 39544 19893 39584
rect 19851 39535 19893 39544
rect 19660 39500 19700 39509
rect 19700 39460 19796 39500
rect 19660 39451 19700 39460
rect 19467 39416 19509 39425
rect 19467 39376 19468 39416
rect 19508 39376 19509 39416
rect 19467 39367 19509 39376
rect 19276 39040 19412 39080
rect 19276 38996 19316 39040
rect 19660 38996 19700 39005
rect 19276 38947 19316 38956
rect 19564 38956 19660 38996
rect 19371 38912 19413 38921
rect 19371 38872 19372 38912
rect 19412 38872 19413 38912
rect 19371 38863 19413 38872
rect 19179 38072 19221 38081
rect 19179 38032 19180 38072
rect 19220 38032 19221 38072
rect 19179 38023 19221 38032
rect 19275 37988 19317 37997
rect 19275 37948 19276 37988
rect 19316 37948 19317 37988
rect 19275 37939 19317 37948
rect 19276 37854 19316 37939
rect 18808 37820 19176 37829
rect 18848 37780 18890 37820
rect 18930 37780 18972 37820
rect 19012 37780 19054 37820
rect 19094 37780 19136 37820
rect 18808 37771 19176 37780
rect 19179 37652 19221 37661
rect 19179 37612 19180 37652
rect 19220 37612 19221 37652
rect 19179 37603 19221 37612
rect 19180 37518 19220 37603
rect 18988 37400 19028 37409
rect 19028 37360 19316 37400
rect 18988 37351 19028 37360
rect 18699 37316 18741 37325
rect 18699 37276 18700 37316
rect 18740 37276 18741 37316
rect 18699 37267 18741 37276
rect 18452 36856 18644 36896
rect 18412 36847 18452 36856
rect 18028 36688 18356 36728
rect 18220 36560 18260 36569
rect 17932 36352 18164 36392
rect 17836 36091 17876 36100
rect 18027 36140 18069 36149
rect 18027 36100 18028 36140
rect 18068 36100 18069 36140
rect 18027 36091 18069 36100
rect 17835 35888 17877 35897
rect 17835 35848 17836 35888
rect 17876 35848 17877 35888
rect 17835 35839 17877 35848
rect 18028 35888 18068 36091
rect 18028 35839 18068 35848
rect 17836 34376 17876 35839
rect 18027 35216 18069 35225
rect 18027 35176 18028 35216
rect 18068 35176 18069 35216
rect 18027 35167 18069 35176
rect 18124 35216 18164 36352
rect 18220 36233 18260 36520
rect 18219 36224 18261 36233
rect 18219 36184 18220 36224
rect 18260 36184 18261 36224
rect 18219 36175 18261 36184
rect 18316 36056 18356 36688
rect 18604 36728 18644 36737
rect 18700 36728 18740 37267
rect 18891 36896 18933 36905
rect 18891 36856 18892 36896
rect 18932 36856 18933 36896
rect 18891 36847 18933 36856
rect 18644 36688 18740 36728
rect 18604 36679 18644 36688
rect 18892 36560 18932 36847
rect 18124 35167 18164 35176
rect 18220 36016 18356 36056
rect 18412 36520 18932 36560
rect 18028 35082 18068 35167
rect 18123 34628 18165 34637
rect 18123 34588 18124 34628
rect 18164 34588 18165 34628
rect 18123 34579 18165 34588
rect 18028 34376 18068 34385
rect 17836 34327 17876 34336
rect 17932 34336 18028 34376
rect 17932 34208 17972 34336
rect 18028 34327 18068 34336
rect 18124 34376 18164 34579
rect 18124 34327 18164 34336
rect 18220 34208 18260 36016
rect 17740 34168 17972 34208
rect 18028 34168 18260 34208
rect 18316 34376 18356 34385
rect 17931 33956 17973 33965
rect 17931 33916 17932 33956
rect 17972 33916 17973 33956
rect 17931 33907 17973 33916
rect 17164 33244 17396 33284
rect 17452 33704 17492 33713
rect 17164 32285 17204 33244
rect 17259 32864 17301 32873
rect 17259 32824 17260 32864
rect 17300 32824 17301 32864
rect 17259 32815 17301 32824
rect 17356 32869 17396 32878
rect 17163 32276 17205 32285
rect 17163 32236 17164 32276
rect 17204 32236 17205 32276
rect 17163 32227 17205 32236
rect 17164 31613 17204 31698
rect 17163 31604 17205 31613
rect 17163 31564 17164 31604
rect 17204 31564 17205 31604
rect 17163 31555 17205 31564
rect 17164 31361 17204 31446
rect 17163 31352 17205 31361
rect 17163 31312 17164 31352
rect 17204 31312 17205 31352
rect 17163 31303 17205 31312
rect 16875 31228 16876 31268
rect 16916 31228 16917 31268
rect 16875 31219 16917 31228
rect 16972 31228 17108 31268
rect 16876 30689 16916 31219
rect 16875 30680 16917 30689
rect 16875 30640 16876 30680
rect 16916 30640 16917 30680
rect 16875 30631 16917 30640
rect 16972 30680 17012 31228
rect 17067 31100 17109 31109
rect 17067 31060 17068 31100
rect 17108 31060 17109 31100
rect 17067 31051 17109 31060
rect 16875 30512 16917 30521
rect 16875 30472 16876 30512
rect 16916 30472 16917 30512
rect 16875 30463 16917 30472
rect 16779 29252 16821 29261
rect 16779 29212 16780 29252
rect 16820 29212 16821 29252
rect 16779 29203 16821 29212
rect 16684 28960 16820 29000
rect 16587 28951 16629 28960
rect 16492 28328 16532 28337
rect 16492 27749 16532 28288
rect 16588 28328 16628 28337
rect 16588 28085 16628 28288
rect 16587 28076 16629 28085
rect 16587 28036 16588 28076
rect 16628 28036 16629 28076
rect 16587 28027 16629 28036
rect 16491 27740 16533 27749
rect 16491 27700 16492 27740
rect 16532 27700 16533 27740
rect 16491 27691 16533 27700
rect 16396 27196 16532 27236
rect 16396 26993 16436 27078
rect 16395 26984 16437 26993
rect 16395 26944 16396 26984
rect 16436 26944 16437 26984
rect 16395 26935 16437 26944
rect 16396 26816 16436 26825
rect 16299 26480 16341 26489
rect 16299 26440 16300 26480
rect 16340 26440 16341 26480
rect 16299 26431 16341 26440
rect 16396 26321 16436 26776
rect 16395 26312 16437 26321
rect 16395 26272 16396 26312
rect 16436 26272 16437 26312
rect 16395 26263 16437 26272
rect 16203 26228 16245 26237
rect 16203 26188 16204 26228
rect 16244 26188 16245 26228
rect 16203 26179 16245 26188
rect 16395 26144 16437 26153
rect 16395 26104 16396 26144
rect 16436 26104 16437 26144
rect 16395 26095 16437 26104
rect 16203 26060 16245 26069
rect 16203 26020 16204 26060
rect 16244 26020 16245 26060
rect 16203 26011 16245 26020
rect 16011 24508 16012 24548
rect 16052 24508 16148 24548
rect 16011 24499 16053 24508
rect 16204 24464 16244 26011
rect 16299 25304 16341 25313
rect 16299 25264 16300 25304
rect 16340 25264 16341 25304
rect 16299 25255 16341 25264
rect 16300 24641 16340 25255
rect 16299 24632 16341 24641
rect 16299 24592 16300 24632
rect 16340 24592 16341 24632
rect 16299 24583 16341 24592
rect 16108 24424 16244 24464
rect 15916 24380 15956 24389
rect 15916 23381 15956 24340
rect 15915 23372 15957 23381
rect 15915 23332 15916 23372
rect 15956 23332 15957 23372
rect 15915 23323 15957 23332
rect 15764 23080 15860 23120
rect 15724 23071 15764 23080
rect 15820 22793 15860 23080
rect 15627 22784 15669 22793
rect 15627 22744 15628 22784
rect 15668 22744 15669 22784
rect 15627 22735 15669 22744
rect 15819 22784 15861 22793
rect 15819 22744 15820 22784
rect 15860 22744 15861 22784
rect 15819 22735 15861 22744
rect 15339 22364 15381 22373
rect 15339 22324 15340 22364
rect 15380 22324 15381 22364
rect 15339 22315 15381 22324
rect 15436 22324 15860 22364
rect 15243 22280 15285 22289
rect 15243 22240 15244 22280
rect 15284 22240 15285 22280
rect 15243 22231 15285 22240
rect 15340 22280 15380 22315
rect 15244 22146 15284 22231
rect 15340 22230 15380 22240
rect 15436 22280 15476 22324
rect 15436 22205 15476 22240
rect 15820 22280 15860 22324
rect 15916 22289 15956 22374
rect 16108 22289 16148 24424
rect 16203 23372 16245 23381
rect 16203 23332 16204 23372
rect 16244 23332 16245 23372
rect 16203 23323 16245 23332
rect 15820 22231 15860 22240
rect 15915 22280 15957 22289
rect 15915 22240 15916 22280
rect 15956 22240 15957 22280
rect 15915 22231 15957 22240
rect 16012 22280 16052 22289
rect 15435 22196 15477 22205
rect 15435 22156 15436 22196
rect 15476 22156 15477 22196
rect 15435 22147 15477 22156
rect 15628 22112 15668 22121
rect 16012 22112 16052 22240
rect 16107 22280 16149 22289
rect 16107 22240 16108 22280
rect 16148 22240 16149 22280
rect 16107 22231 16149 22240
rect 15668 22072 16052 22112
rect 16108 22112 16148 22121
rect 15628 22063 15668 22072
rect 15148 21988 15380 22028
rect 15244 21608 15284 21617
rect 15244 21197 15284 21568
rect 15243 21188 15285 21197
rect 15243 21148 15244 21188
rect 15284 21148 15285 21188
rect 15243 21139 15285 21148
rect 15147 21020 15189 21029
rect 15147 20980 15148 21020
rect 15188 20980 15189 21020
rect 15147 20971 15189 20980
rect 15148 20768 15188 20971
rect 15148 20719 15188 20728
rect 15147 20600 15189 20609
rect 15147 20560 15148 20600
rect 15188 20560 15189 20600
rect 15147 20551 15189 20560
rect 15051 20348 15093 20357
rect 14860 20308 14996 20348
rect 14763 20299 14805 20308
rect 14572 19048 14708 19088
rect 14475 18836 14517 18845
rect 14475 18796 14476 18836
rect 14516 18796 14517 18836
rect 14475 18787 14517 18796
rect 14380 18628 14516 18668
rect 14188 17744 14228 18451
rect 14188 17695 14228 17704
rect 14284 17669 14324 18460
rect 14379 18500 14421 18509
rect 14379 18460 14380 18500
rect 14420 18460 14421 18500
rect 14379 18451 14421 18460
rect 14091 17660 14133 17669
rect 14091 17620 14092 17660
rect 14132 17620 14133 17660
rect 14091 17611 14133 17620
rect 14283 17660 14325 17669
rect 14283 17620 14284 17660
rect 14324 17620 14325 17660
rect 14283 17611 14325 17620
rect 14092 16241 14132 17611
rect 14380 17417 14420 18451
rect 14379 17408 14421 17417
rect 14379 17368 14380 17408
rect 14420 17368 14421 17408
rect 14379 17359 14421 17368
rect 14188 16325 14228 16410
rect 14380 16325 14420 17359
rect 14187 16316 14229 16325
rect 14187 16276 14188 16316
rect 14228 16276 14229 16316
rect 14187 16267 14229 16276
rect 14379 16316 14421 16325
rect 14379 16276 14380 16316
rect 14420 16276 14421 16316
rect 14379 16267 14421 16276
rect 14091 16232 14133 16241
rect 14091 16192 14092 16232
rect 14132 16192 14133 16232
rect 14091 16183 14133 16192
rect 14091 16064 14133 16073
rect 14091 16024 14092 16064
rect 14132 16024 14133 16064
rect 14091 16015 14133 16024
rect 14092 14804 14132 16015
rect 14283 15140 14325 15149
rect 14283 15100 14284 15140
rect 14324 15100 14325 15140
rect 14283 15091 14325 15100
rect 14092 14755 14132 14764
rect 14187 14804 14229 14813
rect 14187 14764 14188 14804
rect 14228 14764 14229 14804
rect 14187 14755 14229 14764
rect 14188 14670 14228 14755
rect 14091 13460 14133 13469
rect 14091 13420 14092 13460
rect 14132 13420 14133 13460
rect 14091 13411 14133 13420
rect 14092 13208 14132 13411
rect 14092 13159 14132 13168
rect 14284 11705 14324 15091
rect 14476 14300 14516 18628
rect 14380 14260 14516 14300
rect 14283 11696 14325 11705
rect 14283 11656 14284 11696
rect 14324 11656 14325 11696
rect 14283 11647 14325 11656
rect 14091 11444 14133 11453
rect 14091 11404 14092 11444
rect 14132 11404 14133 11444
rect 14091 11395 14133 11404
rect 14092 7916 14132 11395
rect 14283 11192 14325 11201
rect 14283 11152 14284 11192
rect 14324 11152 14325 11192
rect 14380 11192 14420 14260
rect 14572 14216 14612 19048
rect 14667 18752 14709 18761
rect 14667 18712 14668 18752
rect 14708 18712 14709 18752
rect 14667 18703 14709 18712
rect 14668 18089 14708 18703
rect 14667 18080 14709 18089
rect 14667 18040 14668 18080
rect 14708 18040 14709 18080
rect 14667 18031 14709 18040
rect 14667 17744 14709 17753
rect 14667 17704 14668 17744
rect 14708 17704 14709 17744
rect 14667 17695 14709 17704
rect 14668 16232 14708 17695
rect 14668 16073 14708 16192
rect 14667 16064 14709 16073
rect 14667 16024 14668 16064
rect 14708 16024 14709 16064
rect 14667 16015 14709 16024
rect 14764 15812 14804 20299
rect 14859 20096 14901 20105
rect 14859 20056 14860 20096
rect 14900 20056 14901 20096
rect 14859 20047 14901 20056
rect 14956 20096 14996 20308
rect 15051 20308 15052 20348
rect 15092 20308 15093 20348
rect 15051 20299 15093 20308
rect 15051 20180 15093 20189
rect 15051 20140 15052 20180
rect 15092 20140 15093 20180
rect 15051 20131 15093 20140
rect 14956 20047 14996 20056
rect 14860 18761 14900 20047
rect 15052 20046 15092 20131
rect 15148 20096 15188 20551
rect 15340 20180 15380 21988
rect 16108 21860 16148 22072
rect 15628 21820 16148 21860
rect 15628 21692 15668 21820
rect 15628 21643 15668 21652
rect 15531 21608 15573 21617
rect 15531 21568 15532 21608
rect 15572 21568 15573 21608
rect 15531 21559 15573 21568
rect 16107 21608 16149 21617
rect 16107 21568 16108 21608
rect 16148 21568 16149 21608
rect 16107 21559 16149 21568
rect 15532 21474 15572 21559
rect 15627 21524 15669 21533
rect 15627 21484 15628 21524
rect 15668 21484 15669 21524
rect 15627 21475 15669 21484
rect 15148 20047 15188 20056
rect 15244 20140 15380 20180
rect 15244 20096 15284 20140
rect 15147 19340 15189 19349
rect 15147 19300 15148 19340
rect 15188 19300 15189 19340
rect 15147 19291 15189 19300
rect 15052 19256 15092 19265
rect 15052 18929 15092 19216
rect 15051 18920 15093 18929
rect 15051 18880 15052 18920
rect 15092 18880 15093 18920
rect 15051 18871 15093 18880
rect 14859 18752 14901 18761
rect 14859 18712 14860 18752
rect 14900 18712 14901 18752
rect 14859 18703 14901 18712
rect 14860 18584 14900 18593
rect 15052 18584 15092 18871
rect 14900 18544 15092 18584
rect 14860 17753 14900 18544
rect 14859 17744 14901 17753
rect 14859 17704 14860 17744
rect 14900 17704 14901 17744
rect 14859 17695 14901 17704
rect 15148 16409 15188 19291
rect 15244 17921 15284 20056
rect 15532 19265 15572 19351
rect 15531 19261 15573 19265
rect 15531 19216 15532 19261
rect 15572 19216 15573 19261
rect 15531 19207 15573 19216
rect 15628 18920 15668 21475
rect 15915 21440 15957 21449
rect 15915 21400 15916 21440
rect 15956 21400 15957 21440
rect 15915 21391 15957 21400
rect 15916 21306 15956 21391
rect 16108 21113 16148 21559
rect 16107 21104 16149 21113
rect 16107 21064 16108 21104
rect 16148 21064 16149 21104
rect 16107 21055 16149 21064
rect 15724 19552 15956 19592
rect 15724 19265 15764 19552
rect 15916 19508 15956 19552
rect 15916 19459 15956 19468
rect 15819 19424 15861 19433
rect 15819 19384 15820 19424
rect 15860 19384 15861 19424
rect 15819 19375 15861 19384
rect 15723 19256 15765 19265
rect 15723 19216 15724 19256
rect 15764 19216 15765 19256
rect 15723 19207 15765 19216
rect 15820 19088 15860 19375
rect 16107 19340 16149 19349
rect 16107 19300 16108 19340
rect 16148 19300 16149 19340
rect 16107 19298 16149 19300
rect 16107 19291 16108 19298
rect 16148 19291 16149 19298
rect 16108 19205 16148 19258
rect 15724 19048 15860 19088
rect 15724 19046 15764 19048
rect 15724 18997 15764 19006
rect 15820 19004 15860 19048
rect 15820 18964 16052 19004
rect 15628 18880 15860 18920
rect 15532 18677 15572 18762
rect 15531 18668 15573 18677
rect 15531 18628 15532 18668
rect 15572 18628 15573 18668
rect 15531 18619 15573 18628
rect 15388 18542 15428 18551
rect 15388 18416 15428 18502
rect 15388 18376 15668 18416
rect 15531 18248 15573 18257
rect 15531 18208 15532 18248
rect 15572 18208 15573 18248
rect 15531 18199 15573 18208
rect 15435 18080 15477 18089
rect 15435 18040 15436 18080
rect 15476 18040 15477 18080
rect 15435 18031 15477 18040
rect 15243 17912 15285 17921
rect 15243 17872 15244 17912
rect 15284 17872 15285 17912
rect 15243 17863 15285 17872
rect 15436 17744 15476 18031
rect 15532 18005 15572 18199
rect 15531 17996 15573 18005
rect 15531 17956 15532 17996
rect 15572 17956 15573 17996
rect 15531 17947 15573 17956
rect 15628 17996 15668 18376
rect 15628 17947 15668 17956
rect 15436 17695 15476 17704
rect 15532 17072 15572 17947
rect 15627 17660 15669 17669
rect 15627 17620 15628 17660
rect 15668 17620 15669 17660
rect 15627 17611 15669 17620
rect 15339 16484 15381 16493
rect 15339 16444 15340 16484
rect 15380 16444 15381 16484
rect 15339 16435 15381 16444
rect 15147 16400 15189 16409
rect 15052 16360 15148 16400
rect 15188 16360 15189 16400
rect 15052 16148 15092 16360
rect 15147 16351 15189 16360
rect 15196 16241 15236 16250
rect 15236 16232 15275 16241
rect 15236 16201 15284 16232
rect 15196 16192 15284 16201
rect 15052 16108 15188 16148
rect 14764 15772 14900 15812
rect 14667 14972 14709 14981
rect 14667 14932 14668 14972
rect 14708 14932 14709 14972
rect 14667 14923 14709 14932
rect 14668 14720 14708 14923
rect 14668 14671 14708 14680
rect 14476 14176 14612 14216
rect 14476 13124 14516 14176
rect 14620 13217 14660 13226
rect 14660 13177 14708 13208
rect 14620 13168 14708 13177
rect 14476 13084 14612 13124
rect 14475 12536 14517 12545
rect 14475 12496 14476 12536
rect 14516 12496 14517 12536
rect 14475 12487 14517 12496
rect 14476 12402 14516 12487
rect 14380 11152 14516 11192
rect 14283 11143 14325 11152
rect 14284 11024 14324 11143
rect 14284 10975 14324 10984
rect 14380 11024 14420 11033
rect 14380 10697 14420 10984
rect 14379 10688 14421 10697
rect 14379 10648 14380 10688
rect 14420 10648 14421 10688
rect 14379 10639 14421 10648
rect 14476 10445 14516 11152
rect 14475 10436 14517 10445
rect 14475 10396 14476 10436
rect 14516 10396 14517 10436
rect 14475 10387 14517 10396
rect 14283 10268 14325 10277
rect 14283 10228 14284 10268
rect 14324 10228 14325 10268
rect 14283 10219 14325 10228
rect 14379 10268 14421 10277
rect 14572 10268 14612 13084
rect 14668 12704 14708 13168
rect 14668 12655 14708 12664
rect 14764 13040 14804 13049
rect 14764 12293 14804 13000
rect 14763 12284 14805 12293
rect 14763 12244 14764 12284
rect 14804 12244 14805 12284
rect 14763 12235 14805 12244
rect 14860 11360 14900 15772
rect 15148 15560 15188 16108
rect 15244 15728 15284 16192
rect 15340 16148 15380 16435
rect 15532 16232 15572 17032
rect 15532 16183 15572 16192
rect 15380 16108 15476 16148
rect 15340 16099 15380 16108
rect 15340 15728 15380 15737
rect 15244 15688 15340 15728
rect 15340 15679 15380 15688
rect 15148 15511 15188 15520
rect 15196 14729 15236 14738
rect 15236 14689 15284 14720
rect 15196 14680 15284 14689
rect 15244 14216 15284 14680
rect 15339 14552 15381 14561
rect 15339 14512 15340 14552
rect 15380 14512 15381 14552
rect 15339 14503 15381 14512
rect 15340 14418 15380 14503
rect 15244 14167 15284 14176
rect 15052 14048 15092 14059
rect 15052 13973 15092 14008
rect 15051 13964 15093 13973
rect 15051 13924 15052 13964
rect 15092 13924 15093 13964
rect 15051 13915 15093 13924
rect 14955 13292 14997 13301
rect 14955 13252 14956 13292
rect 14996 13252 14997 13292
rect 14955 13243 14997 13252
rect 14956 13208 14996 13243
rect 14956 13157 14996 13168
rect 15243 13208 15285 13217
rect 15243 13168 15244 13208
rect 15284 13168 15285 13208
rect 15243 13159 15285 13168
rect 15051 12452 15093 12461
rect 15051 12412 15052 12452
rect 15092 12412 15093 12452
rect 15051 12403 15093 12412
rect 15052 11789 15092 12403
rect 15051 11780 15093 11789
rect 15051 11740 15052 11780
rect 15092 11740 15093 11780
rect 15051 11731 15093 11740
rect 14860 11320 14996 11360
rect 14667 11192 14709 11201
rect 14667 11152 14668 11192
rect 14708 11152 14709 11192
rect 14667 11143 14709 11152
rect 14859 11192 14901 11201
rect 14859 11152 14860 11192
rect 14900 11152 14901 11192
rect 14859 11143 14901 11152
rect 14379 10228 14380 10268
rect 14420 10228 14421 10268
rect 14379 10226 14421 10228
rect 14379 10219 14380 10226
rect 14187 10184 14229 10193
rect 14187 10144 14188 10184
rect 14228 10144 14229 10184
rect 14187 10135 14229 10144
rect 14188 9017 14228 10135
rect 14284 10016 14324 10219
rect 14420 10219 14421 10226
rect 14486 10228 14612 10268
rect 14380 10133 14420 10186
rect 14486 10100 14526 10228
rect 14476 10060 14526 10100
rect 14572 10100 14612 10109
rect 14668 10100 14708 11143
rect 14860 11024 14900 11143
rect 14860 10975 14900 10984
rect 14763 10940 14805 10949
rect 14763 10900 14764 10940
rect 14804 10900 14805 10940
rect 14763 10891 14805 10900
rect 14764 10806 14804 10891
rect 14763 10436 14805 10445
rect 14763 10396 14764 10436
rect 14804 10396 14805 10436
rect 14763 10387 14805 10396
rect 14612 10060 14708 10100
rect 14284 9976 14420 10016
rect 14283 9512 14325 9521
rect 14283 9472 14284 9512
rect 14324 9472 14325 9512
rect 14283 9463 14325 9472
rect 14284 9378 14324 9463
rect 14283 9092 14325 9101
rect 14283 9052 14284 9092
rect 14324 9052 14325 9092
rect 14283 9043 14325 9052
rect 14187 9008 14229 9017
rect 14187 8968 14188 9008
rect 14228 8968 14229 9008
rect 14187 8959 14229 8968
rect 14092 7876 14228 7916
rect 14091 7748 14133 7757
rect 14091 7708 14092 7748
rect 14132 7708 14133 7748
rect 14091 7699 14133 7708
rect 14092 7174 14132 7699
rect 14092 7125 14132 7134
rect 13899 4892 13941 4901
rect 13899 4852 13900 4892
rect 13940 4852 13941 4892
rect 13899 4843 13941 4852
rect 13900 4565 13940 4843
rect 13899 4556 13941 4565
rect 13899 4516 13900 4556
rect 13940 4516 13941 4556
rect 13899 4507 13941 4516
rect 13996 3977 14036 5608
rect 13995 3968 14037 3977
rect 13995 3928 13996 3968
rect 14036 3928 14037 3968
rect 13995 3919 14037 3928
rect 14188 3305 14228 7876
rect 14187 3296 14229 3305
rect 14187 3256 14188 3296
rect 14228 3256 14229 3296
rect 14187 3247 14229 3256
rect 14284 3128 14324 9043
rect 14380 8765 14420 9976
rect 14379 8756 14421 8765
rect 14379 8716 14380 8756
rect 14420 8716 14421 8756
rect 14379 8707 14421 8716
rect 14380 7925 14420 8707
rect 14379 7916 14421 7925
rect 14379 7876 14380 7916
rect 14420 7876 14421 7916
rect 14379 7867 14421 7876
rect 14380 7169 14420 7867
rect 14379 7160 14421 7169
rect 14379 7120 14380 7160
rect 14420 7120 14421 7160
rect 14379 7111 14421 7120
rect 14476 6908 14516 10060
rect 14572 10051 14612 10060
rect 14668 8672 14708 8681
rect 14668 8513 14708 8632
rect 14667 8504 14709 8513
rect 14667 8464 14668 8504
rect 14708 8464 14709 8504
rect 14667 8455 14709 8464
rect 14571 8420 14613 8429
rect 14571 8380 14572 8420
rect 14612 8380 14613 8420
rect 14571 8371 14613 8380
rect 14572 7160 14612 8371
rect 14668 8177 14708 8455
rect 14667 8168 14709 8177
rect 14667 8128 14668 8168
rect 14708 8128 14709 8168
rect 14667 8119 14709 8128
rect 14572 7111 14612 7120
rect 14476 6868 14612 6908
rect 14475 6488 14517 6497
rect 14475 6448 14476 6488
rect 14516 6448 14517 6488
rect 14475 6439 14517 6448
rect 14379 5816 14421 5825
rect 14379 5776 14380 5816
rect 14420 5776 14421 5816
rect 14379 5767 14421 5776
rect 14380 4976 14420 5767
rect 14380 4565 14420 4936
rect 14379 4556 14421 4565
rect 14379 4516 14380 4556
rect 14420 4516 14421 4556
rect 14379 4507 14421 4516
rect 14379 4388 14421 4397
rect 14379 4348 14380 4388
rect 14420 4348 14421 4388
rect 14379 4339 14421 4348
rect 14188 3088 14324 3128
rect 13707 2708 13749 2717
rect 13707 2668 13708 2708
rect 13748 2668 13749 2708
rect 13707 2659 13749 2668
rect 14091 2708 14133 2717
rect 14091 2668 14092 2708
rect 14132 2668 14133 2708
rect 14091 2659 14133 2668
rect 13708 2574 13748 2659
rect 14092 2574 14132 2659
rect 13803 2456 13845 2465
rect 13803 2416 13804 2456
rect 13844 2416 13845 2456
rect 13803 2407 13845 2416
rect 13900 2456 13940 2465
rect 13707 2372 13749 2381
rect 13707 2332 13708 2372
rect 13748 2332 13749 2372
rect 13707 2323 13749 2332
rect 13611 1952 13653 1961
rect 13611 1912 13612 1952
rect 13652 1912 13653 1952
rect 13611 1903 13653 1912
rect 13708 1952 13748 2323
rect 13708 1903 13748 1912
rect 13804 1364 13844 2407
rect 13900 2213 13940 2416
rect 13995 2372 14037 2381
rect 13995 2332 13996 2372
rect 14036 2332 14037 2372
rect 13995 2323 14037 2332
rect 13899 2204 13941 2213
rect 13899 2164 13900 2204
rect 13940 2164 13941 2204
rect 13899 2155 13941 2164
rect 13899 1784 13941 1793
rect 13899 1744 13900 1784
rect 13940 1744 13941 1784
rect 13899 1735 13941 1744
rect 13900 1650 13940 1735
rect 13708 1324 13844 1364
rect 13419 1196 13461 1205
rect 13419 1156 13420 1196
rect 13460 1156 13461 1196
rect 13419 1147 13461 1156
rect 13420 1062 13460 1147
rect 13515 944 13557 953
rect 13515 904 13516 944
rect 13556 904 13557 944
rect 13515 895 13557 904
rect 13612 944 13652 953
rect 13516 80 13556 895
rect 13612 533 13652 904
rect 13611 524 13653 533
rect 13611 484 13612 524
rect 13652 484 13653 524
rect 13611 475 13653 484
rect 13708 80 13748 1324
rect 13996 1280 14036 2323
rect 14091 1868 14133 1877
rect 14091 1828 14092 1868
rect 14132 1828 14133 1868
rect 14091 1819 14133 1828
rect 14092 1734 14132 1819
rect 13900 1240 14036 1280
rect 13803 1196 13845 1205
rect 13803 1156 13804 1196
rect 13844 1156 13845 1196
rect 13803 1147 13845 1156
rect 13804 1062 13844 1147
rect 13900 80 13940 1240
rect 14091 944 14133 953
rect 14091 904 14092 944
rect 14132 904 14133 944
rect 14091 895 14133 904
rect 14092 810 14132 895
rect 14091 692 14133 701
rect 14091 652 14092 692
rect 14132 652 14133 692
rect 14091 643 14133 652
rect 14092 80 14132 643
rect 14188 524 14228 3088
rect 14380 2801 14420 4339
rect 14476 4145 14516 6439
rect 14475 4136 14517 4145
rect 14475 4096 14476 4136
rect 14516 4096 14517 4136
rect 14475 4087 14517 4096
rect 14476 4002 14516 4087
rect 14379 2792 14421 2801
rect 14379 2752 14380 2792
rect 14420 2752 14421 2792
rect 14379 2743 14421 2752
rect 14475 2708 14517 2717
rect 14475 2668 14476 2708
rect 14516 2668 14517 2708
rect 14475 2659 14517 2668
rect 14476 2574 14516 2659
rect 14283 2456 14325 2465
rect 14283 2416 14284 2456
rect 14324 2416 14325 2456
rect 14283 2407 14325 2416
rect 14284 2322 14324 2407
rect 14572 2288 14612 6868
rect 14667 6656 14709 6665
rect 14667 6616 14668 6656
rect 14708 6616 14709 6656
rect 14667 6607 14709 6616
rect 14668 6522 14708 6607
rect 14764 4817 14804 10387
rect 14956 9428 14996 11320
rect 15052 9521 15092 11731
rect 15147 11696 15189 11705
rect 15147 11656 15148 11696
rect 15188 11656 15189 11696
rect 15147 11647 15189 11656
rect 15148 11562 15188 11647
rect 15147 10604 15189 10613
rect 15147 10564 15148 10604
rect 15188 10564 15189 10604
rect 15147 10555 15189 10564
rect 15051 9512 15093 9521
rect 15051 9472 15052 9512
rect 15092 9472 15093 9512
rect 15051 9463 15093 9472
rect 15148 9437 15188 10555
rect 15244 10277 15284 13159
rect 15436 12713 15476 16108
rect 15628 14300 15668 17611
rect 15820 16913 15860 18880
rect 15915 18668 15957 18677
rect 15915 18628 15916 18668
rect 15956 18628 15957 18668
rect 15915 18619 15957 18628
rect 15916 17669 15956 18619
rect 15915 17660 15957 17669
rect 15915 17620 15916 17660
rect 15956 17620 15957 17660
rect 15915 17611 15957 17620
rect 15819 16904 15861 16913
rect 15819 16864 15820 16904
rect 15860 16864 15861 16904
rect 15819 16855 15861 16864
rect 15820 15065 15860 16855
rect 15819 15056 15861 15065
rect 15532 14260 15668 14300
rect 15724 15016 15820 15056
rect 15860 15016 15861 15056
rect 15532 13469 15572 14260
rect 15628 14132 15668 14141
rect 15628 13889 15668 14092
rect 15627 13880 15669 13889
rect 15627 13840 15628 13880
rect 15668 13840 15669 13880
rect 15627 13831 15669 13840
rect 15531 13460 15573 13469
rect 15531 13420 15532 13460
rect 15572 13420 15668 13460
rect 15531 13411 15573 13420
rect 15435 12704 15477 12713
rect 15435 12664 15436 12704
rect 15476 12664 15572 12704
rect 15435 12655 15477 12664
rect 15340 12536 15380 12545
rect 15340 11948 15380 12496
rect 15340 11899 15380 11908
rect 15436 12536 15476 12545
rect 15436 11201 15476 12496
rect 15435 11192 15477 11201
rect 15435 11152 15436 11192
rect 15476 11152 15477 11192
rect 15435 11143 15477 11152
rect 15340 11024 15380 11033
rect 15243 10268 15285 10277
rect 15243 10228 15244 10268
rect 15284 10228 15285 10268
rect 15243 10219 15285 10228
rect 14860 9388 14996 9428
rect 15147 9428 15189 9437
rect 15147 9388 15148 9428
rect 15188 9388 15189 9428
rect 14860 9008 14900 9388
rect 15147 9379 15189 9388
rect 14860 8968 14996 9008
rect 14859 8840 14901 8849
rect 14859 8800 14860 8840
rect 14900 8800 14901 8840
rect 14859 8791 14901 8800
rect 14860 8706 14900 8791
rect 14860 8000 14900 8011
rect 14860 7925 14900 7960
rect 14859 7916 14901 7925
rect 14859 7876 14860 7916
rect 14900 7876 14901 7916
rect 14859 7867 14901 7876
rect 14859 7664 14901 7673
rect 14859 7624 14860 7664
rect 14900 7624 14901 7664
rect 14859 7615 14901 7624
rect 14860 6497 14900 7615
rect 14859 6488 14901 6497
rect 14859 6448 14860 6488
rect 14900 6448 14901 6488
rect 14859 6439 14901 6448
rect 14860 4962 14900 4971
rect 14763 4808 14805 4817
rect 14763 4768 14764 4808
rect 14804 4768 14805 4808
rect 14763 4759 14805 4768
rect 14860 4640 14900 4922
rect 14668 4600 14900 4640
rect 14668 4388 14708 4600
rect 14956 4556 14996 8968
rect 15148 8672 15188 8681
rect 15052 8168 15092 8177
rect 15148 8168 15188 8632
rect 15092 8128 15188 8168
rect 15244 8672 15284 8681
rect 15052 8119 15092 8128
rect 15244 8009 15284 8632
rect 15340 8429 15380 10984
rect 15532 10949 15572 12664
rect 15628 11360 15668 13420
rect 15724 11537 15764 15016
rect 15819 15007 15861 15016
rect 15916 14552 15956 14561
rect 15820 14512 15916 14552
rect 15820 14043 15860 14512
rect 15916 14503 15956 14512
rect 15820 13994 15860 14003
rect 15819 12704 15861 12713
rect 15819 12664 15820 12704
rect 15860 12664 15861 12704
rect 15819 12655 15861 12664
rect 15820 12536 15860 12655
rect 15820 12487 15860 12496
rect 15916 12536 15956 12545
rect 16012 12536 16052 18964
rect 16108 18509 16148 18594
rect 16107 18500 16149 18509
rect 16107 18460 16108 18500
rect 16148 18460 16149 18500
rect 16107 18451 16149 18460
rect 16107 18332 16149 18341
rect 16107 18292 16108 18332
rect 16148 18292 16149 18332
rect 16107 18283 16149 18292
rect 16108 15224 16148 18283
rect 16204 15401 16244 23323
rect 16300 19433 16340 24583
rect 16396 22289 16436 26095
rect 16492 24221 16532 27196
rect 16588 26816 16628 26825
rect 16588 26405 16628 26776
rect 16683 26816 16725 26825
rect 16683 26776 16684 26816
rect 16724 26776 16725 26816
rect 16683 26767 16725 26776
rect 16684 26682 16724 26767
rect 16587 26396 16629 26405
rect 16587 26356 16588 26396
rect 16628 26356 16629 26396
rect 16587 26347 16629 26356
rect 16587 24632 16629 24641
rect 16587 24592 16588 24632
rect 16628 24592 16629 24632
rect 16587 24583 16629 24592
rect 16588 24498 16628 24583
rect 16780 24380 16820 28960
rect 16876 27329 16916 30463
rect 16972 30017 17012 30640
rect 17068 30353 17108 31051
rect 17260 30689 17300 32815
rect 17356 32789 17396 32829
rect 17355 32780 17397 32789
rect 17355 32740 17356 32780
rect 17396 32740 17397 32780
rect 17452 32780 17492 33664
rect 17548 33704 17588 33713
rect 17548 32864 17588 33664
rect 17836 33452 17876 33461
rect 17548 32824 17684 32864
rect 17452 32740 17588 32780
rect 17355 32731 17397 32740
rect 17356 32612 17396 32731
rect 17548 32696 17588 32740
rect 17548 32647 17588 32656
rect 17356 32572 17492 32612
rect 17452 32187 17492 32572
rect 17644 32360 17684 32824
rect 17739 32780 17781 32789
rect 17739 32740 17740 32780
rect 17780 32740 17781 32780
rect 17739 32731 17781 32740
rect 17740 32646 17780 32731
rect 17644 32311 17684 32320
rect 17452 32138 17492 32147
rect 17836 31445 17876 33412
rect 17932 32864 17972 33907
rect 17932 32815 17972 32824
rect 17644 31436 17684 31445
rect 17548 31396 17644 31436
rect 17355 31352 17397 31361
rect 17355 31312 17356 31352
rect 17396 31312 17397 31352
rect 17355 31303 17397 31312
rect 17452 31352 17492 31361
rect 17356 31218 17396 31303
rect 17452 31109 17492 31312
rect 17451 31100 17493 31109
rect 17451 31060 17452 31100
rect 17492 31060 17493 31100
rect 17451 31051 17493 31060
rect 17259 30680 17301 30689
rect 17259 30640 17260 30680
rect 17300 30640 17301 30680
rect 17259 30631 17301 30640
rect 17163 30596 17205 30605
rect 17163 30556 17164 30596
rect 17204 30556 17205 30596
rect 17163 30547 17205 30556
rect 17356 30596 17396 30605
rect 17067 30344 17109 30353
rect 17067 30304 17068 30344
rect 17108 30304 17109 30344
rect 17067 30295 17109 30304
rect 17164 30092 17204 30547
rect 17259 30344 17301 30353
rect 17259 30304 17260 30344
rect 17300 30304 17301 30344
rect 17259 30295 17301 30304
rect 17164 30043 17204 30052
rect 16971 30008 17013 30017
rect 16971 29968 16972 30008
rect 17012 29968 17013 30008
rect 16971 29959 17013 29968
rect 16971 29840 17013 29849
rect 16971 29800 16972 29840
rect 17012 29800 17013 29840
rect 16971 29791 17013 29800
rect 17163 29840 17205 29849
rect 17163 29800 17164 29840
rect 17204 29800 17205 29840
rect 17163 29791 17205 29800
rect 16972 29706 17012 29791
rect 17067 29756 17109 29765
rect 17067 29716 17068 29756
rect 17108 29716 17109 29756
rect 17067 29707 17109 29716
rect 17068 28505 17108 29707
rect 17164 29177 17204 29791
rect 17163 29168 17205 29177
rect 17163 29128 17164 29168
rect 17204 29128 17205 29168
rect 17163 29119 17205 29128
rect 17067 28496 17109 28505
rect 17067 28456 17068 28496
rect 17108 28456 17109 28496
rect 17067 28447 17109 28456
rect 16971 28412 17013 28421
rect 16971 28372 16972 28412
rect 17012 28372 17013 28412
rect 16971 28363 17013 28372
rect 17068 28412 17108 28447
rect 16972 28278 17012 28363
rect 17068 28362 17108 28372
rect 17164 28244 17204 29119
rect 17068 28204 17204 28244
rect 16972 27656 17012 27665
rect 17068 27656 17108 28204
rect 17163 27740 17205 27749
rect 17163 27700 17164 27740
rect 17204 27700 17205 27740
rect 17163 27691 17205 27700
rect 17012 27616 17108 27656
rect 16875 27320 16917 27329
rect 16875 27280 16876 27320
rect 16916 27280 16917 27320
rect 16875 27271 16917 27280
rect 16972 26321 17012 27616
rect 17164 27606 17204 27691
rect 17067 26480 17109 26489
rect 17067 26440 17068 26480
rect 17108 26440 17109 26480
rect 17067 26431 17109 26440
rect 16971 26312 17013 26321
rect 16971 26272 16972 26312
rect 17012 26272 17013 26312
rect 16971 26263 17013 26272
rect 16971 26144 17013 26153
rect 16971 26104 16972 26144
rect 17012 26104 17013 26144
rect 16971 26095 17013 26104
rect 16875 25892 16917 25901
rect 16875 25852 16876 25892
rect 16916 25852 16917 25892
rect 16875 25843 16917 25852
rect 16876 25304 16916 25843
rect 16876 25255 16916 25264
rect 16972 25304 17012 26095
rect 16972 25255 17012 25264
rect 16875 24548 16917 24557
rect 16875 24508 16876 24548
rect 16916 24508 16917 24548
rect 16875 24499 16917 24508
rect 16694 24340 16820 24380
rect 16694 24296 16734 24340
rect 16684 24256 16734 24296
rect 16491 24212 16533 24221
rect 16684 24212 16724 24256
rect 16491 24172 16492 24212
rect 16532 24172 16533 24212
rect 16491 24163 16533 24172
rect 16588 24172 16724 24212
rect 16779 24212 16821 24221
rect 16779 24172 16780 24212
rect 16820 24172 16821 24212
rect 16491 23120 16533 23129
rect 16491 23080 16492 23120
rect 16532 23080 16533 23120
rect 16491 23071 16533 23080
rect 16395 22280 16437 22289
rect 16395 22240 16396 22280
rect 16436 22240 16437 22280
rect 16395 22231 16437 22240
rect 16396 20768 16436 20777
rect 16396 19937 16436 20728
rect 16492 20273 16532 23071
rect 16491 20264 16533 20273
rect 16491 20224 16492 20264
rect 16532 20224 16533 20264
rect 16491 20215 16533 20224
rect 16492 20096 16532 20105
rect 16395 19928 16437 19937
rect 16395 19888 16396 19928
rect 16436 19888 16437 19928
rect 16395 19879 16437 19888
rect 16395 19760 16437 19769
rect 16395 19720 16396 19760
rect 16436 19720 16437 19760
rect 16395 19711 16437 19720
rect 16299 19424 16341 19433
rect 16299 19384 16300 19424
rect 16340 19384 16341 19424
rect 16299 19375 16341 19384
rect 16299 18752 16341 18761
rect 16299 18712 16300 18752
rect 16340 18712 16341 18752
rect 16299 18703 16341 18712
rect 16300 18618 16340 18703
rect 16396 18509 16436 19711
rect 16492 19685 16532 20056
rect 16491 19676 16533 19685
rect 16491 19636 16492 19676
rect 16532 19636 16533 19676
rect 16491 19627 16533 19636
rect 16492 19517 16532 19627
rect 16491 19508 16533 19517
rect 16491 19468 16492 19508
rect 16532 19468 16533 19508
rect 16491 19459 16533 19468
rect 16491 18752 16533 18761
rect 16491 18712 16492 18752
rect 16532 18712 16533 18752
rect 16491 18703 16533 18712
rect 16492 18618 16532 18703
rect 16395 18500 16437 18509
rect 16395 18460 16396 18500
rect 16436 18460 16437 18500
rect 16395 18451 16437 18460
rect 16299 18416 16341 18425
rect 16299 18376 16300 18416
rect 16340 18376 16341 18416
rect 16299 18367 16341 18376
rect 16300 17837 16340 18367
rect 16299 17828 16341 17837
rect 16299 17788 16300 17828
rect 16340 17788 16341 17828
rect 16299 17779 16341 17788
rect 16396 17081 16436 18451
rect 16588 17753 16628 24172
rect 16779 24163 16821 24172
rect 16683 24044 16725 24053
rect 16683 24004 16684 24044
rect 16724 24004 16725 24044
rect 16683 23995 16725 24004
rect 16684 20189 16724 23995
rect 16683 20180 16725 20189
rect 16683 20140 16684 20180
rect 16724 20140 16725 20180
rect 16683 20131 16725 20140
rect 16684 18500 16724 18509
rect 16587 17744 16629 17753
rect 16587 17704 16588 17744
rect 16628 17704 16629 17744
rect 16587 17695 16629 17704
rect 16684 17324 16724 18460
rect 16588 17284 16724 17324
rect 16395 17072 16437 17081
rect 16395 17032 16396 17072
rect 16436 17032 16437 17072
rect 16395 17023 16437 17032
rect 16588 16241 16628 17284
rect 16780 17240 16820 24163
rect 16876 17996 16916 24499
rect 16972 23792 17012 23801
rect 16972 23120 17012 23752
rect 16972 19349 17012 23080
rect 16971 19340 17013 19349
rect 16971 19300 16972 19340
rect 17012 19300 17013 19340
rect 16971 19291 17013 19300
rect 16876 17956 17012 17996
rect 16972 17828 17012 17956
rect 17068 17912 17108 26431
rect 17164 26144 17204 26153
rect 17164 25985 17204 26104
rect 17163 25976 17205 25985
rect 17163 25936 17164 25976
rect 17204 25936 17205 25976
rect 17163 25927 17205 25936
rect 17260 24557 17300 30295
rect 17356 29681 17396 30556
rect 17451 30596 17493 30605
rect 17451 30556 17452 30596
rect 17492 30556 17493 30596
rect 17451 30547 17493 30556
rect 17452 30462 17492 30547
rect 17452 29840 17492 29849
rect 17355 29672 17397 29681
rect 17355 29632 17356 29672
rect 17396 29632 17397 29672
rect 17355 29623 17397 29632
rect 17355 29504 17397 29513
rect 17355 29464 17356 29504
rect 17396 29464 17397 29504
rect 17355 29455 17397 29464
rect 17356 26060 17396 29455
rect 17452 28841 17492 29800
rect 17451 28832 17493 28841
rect 17451 28792 17452 28832
rect 17492 28792 17493 28832
rect 17451 28783 17493 28792
rect 17452 28673 17492 28783
rect 17451 28664 17493 28673
rect 17451 28624 17452 28664
rect 17492 28624 17493 28664
rect 17451 28615 17493 28624
rect 17548 28496 17588 31396
rect 17644 31387 17684 31396
rect 17835 31436 17877 31445
rect 17835 31396 17836 31436
rect 17876 31396 17877 31436
rect 17835 31387 17877 31396
rect 17836 31184 17876 31193
rect 17836 30017 17876 31144
rect 17931 30680 17973 30689
rect 17931 30640 17932 30680
rect 17972 30640 17973 30680
rect 17931 30631 17973 30640
rect 17932 30546 17972 30631
rect 17835 30008 17877 30017
rect 17835 29968 17836 30008
rect 17876 29968 17877 30008
rect 17835 29959 17877 29968
rect 18028 29840 18068 34168
rect 18316 33872 18356 34336
rect 18220 33832 18356 33872
rect 18123 32192 18165 32201
rect 18123 32152 18124 32192
rect 18164 32152 18165 32192
rect 18123 32143 18165 32152
rect 18124 32058 18164 32143
rect 18220 32033 18260 33832
rect 18316 33704 18356 33713
rect 18412 33704 18452 36520
rect 18808 36308 19176 36317
rect 18848 36268 18890 36308
rect 18930 36268 18972 36308
rect 19012 36268 19054 36308
rect 19094 36268 19136 36308
rect 18808 36259 19176 36268
rect 19179 36056 19221 36065
rect 19179 36016 19180 36056
rect 19220 36016 19221 36056
rect 19276 36056 19316 37360
rect 19372 36317 19412 38863
rect 19564 38837 19604 38956
rect 19660 38947 19700 38956
rect 19756 38921 19796 39460
rect 19755 38912 19797 38921
rect 19755 38872 19756 38912
rect 19796 38872 19797 38912
rect 19755 38863 19797 38872
rect 19563 38828 19605 38837
rect 19563 38788 19564 38828
rect 19604 38788 19605 38828
rect 19563 38779 19605 38788
rect 19467 38744 19509 38753
rect 19852 38744 19892 38753
rect 19467 38704 19468 38744
rect 19508 38704 19509 38744
rect 19467 38695 19509 38704
rect 19660 38704 19852 38744
rect 19468 38610 19508 38695
rect 19467 38492 19509 38501
rect 19467 38452 19468 38492
rect 19508 38452 19509 38492
rect 19467 38443 19509 38452
rect 19468 38072 19508 38443
rect 19468 38023 19508 38032
rect 19563 37484 19605 37493
rect 19563 37444 19564 37484
rect 19604 37444 19605 37484
rect 19563 37435 19605 37444
rect 19564 36905 19604 37435
rect 19660 37241 19700 38704
rect 19852 38695 19892 38704
rect 19755 38240 19797 38249
rect 19755 38200 19756 38240
rect 19796 38200 19797 38240
rect 19755 38191 19797 38200
rect 19852 38240 19892 38249
rect 19756 38106 19796 38191
rect 19659 37232 19701 37241
rect 19659 37192 19660 37232
rect 19700 37192 19701 37232
rect 19659 37183 19701 37192
rect 19563 36896 19605 36905
rect 19563 36856 19564 36896
rect 19604 36856 19605 36896
rect 19852 36896 19892 38200
rect 19948 37157 19988 40216
rect 20044 40207 20084 40216
rect 20048 40088 20416 40097
rect 20088 40048 20130 40088
rect 20170 40048 20212 40088
rect 20252 40048 20294 40088
rect 20334 40048 20376 40088
rect 20048 40039 20416 40048
rect 20044 39668 20084 39677
rect 20044 39509 20084 39628
rect 20043 39500 20085 39509
rect 20043 39460 20044 39500
rect 20084 39460 20085 39500
rect 20043 39451 20085 39460
rect 20236 39500 20276 39509
rect 20044 38996 20084 39005
rect 20044 38837 20084 38956
rect 20236 38921 20276 39460
rect 20331 38996 20373 39005
rect 20331 38956 20332 38996
rect 20372 38956 20373 38996
rect 20331 38947 20373 38956
rect 20235 38912 20277 38921
rect 20235 38872 20236 38912
rect 20276 38872 20277 38912
rect 20235 38863 20277 38872
rect 20043 38828 20085 38837
rect 20043 38788 20044 38828
rect 20084 38788 20085 38828
rect 20043 38779 20085 38788
rect 20236 38744 20276 38753
rect 20332 38744 20372 38947
rect 20276 38704 20372 38744
rect 20236 38695 20276 38704
rect 20048 38576 20416 38585
rect 20088 38536 20130 38576
rect 20170 38536 20212 38576
rect 20252 38536 20294 38576
rect 20334 38536 20376 38576
rect 20048 38527 20416 38536
rect 20140 38240 20180 38249
rect 20180 38200 20276 38240
rect 20140 38172 20180 38200
rect 20043 37484 20085 37493
rect 20043 37444 20044 37484
rect 20084 37444 20085 37484
rect 20043 37435 20085 37444
rect 20044 37350 20084 37435
rect 20236 37409 20276 38200
rect 20524 37577 20564 40375
rect 21291 38996 21333 39005
rect 21291 38956 21292 38996
rect 21332 38956 21333 38996
rect 21291 38947 21333 38956
rect 20811 38828 20853 38837
rect 20811 38788 20812 38828
rect 20852 38788 20853 38828
rect 20811 38779 20853 38788
rect 20523 37568 20565 37577
rect 20523 37528 20524 37568
rect 20564 37528 20565 37568
rect 20523 37519 20565 37528
rect 20235 37400 20277 37409
rect 20235 37360 20236 37400
rect 20276 37360 20277 37400
rect 20235 37351 20277 37360
rect 20236 37232 20276 37241
rect 20276 37192 20660 37232
rect 20236 37183 20276 37192
rect 19947 37148 19989 37157
rect 19947 37108 19948 37148
rect 19988 37108 19989 37148
rect 19947 37099 19989 37108
rect 20048 37064 20416 37073
rect 20088 37024 20130 37064
rect 20170 37024 20212 37064
rect 20252 37024 20294 37064
rect 20334 37024 20376 37064
rect 20048 37015 20416 37024
rect 19852 36856 19988 36896
rect 19563 36847 19605 36856
rect 19467 36812 19509 36821
rect 19467 36772 19468 36812
rect 19508 36772 19509 36812
rect 19467 36763 19509 36772
rect 19755 36812 19797 36821
rect 19755 36772 19756 36812
rect 19796 36772 19797 36812
rect 19755 36763 19797 36772
rect 19371 36308 19413 36317
rect 19371 36268 19372 36308
rect 19412 36268 19413 36308
rect 19371 36259 19413 36268
rect 19468 36140 19508 36763
rect 19659 36644 19701 36653
rect 19659 36604 19660 36644
rect 19700 36604 19701 36644
rect 19659 36595 19701 36604
rect 19468 36091 19508 36100
rect 19276 36016 19412 36056
rect 19179 36007 19221 36016
rect 19180 35888 19220 36007
rect 19276 35888 19316 35897
rect 19180 35848 19276 35888
rect 18507 35636 18549 35645
rect 18507 35596 18508 35636
rect 18548 35596 18549 35636
rect 18507 35587 18549 35596
rect 18508 35216 18548 35587
rect 18508 35167 18548 35176
rect 19084 35216 19124 35227
rect 19084 35141 19124 35176
rect 18604 35132 18644 35141
rect 18604 34889 18644 35092
rect 19083 35132 19125 35141
rect 19083 35092 19084 35132
rect 19124 35092 19125 35132
rect 19083 35083 19125 35092
rect 18603 34880 18645 34889
rect 18603 34840 18604 34880
rect 18644 34840 18645 34880
rect 18603 34831 18645 34840
rect 18808 34796 19176 34805
rect 18848 34756 18890 34796
rect 18930 34756 18972 34796
rect 19012 34756 19054 34796
rect 19094 34756 19136 34796
rect 18808 34747 19176 34756
rect 19276 34721 19316 35848
rect 19275 34712 19317 34721
rect 19275 34672 19276 34712
rect 19316 34672 19317 34712
rect 19275 34663 19317 34672
rect 19275 34460 19317 34469
rect 19275 34420 19276 34460
rect 19316 34420 19317 34460
rect 19275 34411 19317 34420
rect 19276 34049 19316 34411
rect 19275 34040 19317 34049
rect 19275 34000 19276 34040
rect 19316 34000 19317 34040
rect 19275 33991 19317 34000
rect 18356 33664 18452 33704
rect 18316 33655 18356 33664
rect 18808 33284 19176 33293
rect 18848 33244 18890 33284
rect 18930 33244 18972 33284
rect 19012 33244 19054 33284
rect 19094 33244 19136 33284
rect 18808 33235 19176 33244
rect 19180 32864 19220 32873
rect 19276 32864 19316 33991
rect 19220 32824 19316 32864
rect 19180 32815 19220 32824
rect 19372 32276 19412 36016
rect 19468 35720 19508 35729
rect 19508 35680 19604 35720
rect 19468 35671 19508 35680
rect 19564 35211 19604 35680
rect 19660 35309 19700 36595
rect 19756 35888 19796 36763
rect 19851 36728 19893 36737
rect 19851 36688 19852 36728
rect 19892 36688 19893 36728
rect 19851 36679 19893 36688
rect 19852 36594 19892 36679
rect 19948 36401 19988 36856
rect 20044 36644 20084 36653
rect 19947 36392 19989 36401
rect 19947 36352 19948 36392
rect 19988 36352 19989 36392
rect 19947 36343 19989 36352
rect 20044 36149 20084 36604
rect 20236 36476 20276 36485
rect 20276 36436 20564 36476
rect 20236 36427 20276 36436
rect 20043 36140 20085 36149
rect 20043 36100 20044 36140
rect 20084 36100 20085 36140
rect 20043 36091 20085 36100
rect 19756 35839 19796 35848
rect 19851 35888 19893 35897
rect 19851 35848 19852 35888
rect 19892 35848 19893 35888
rect 19851 35839 19893 35848
rect 19948 35888 19988 35897
rect 19852 35754 19892 35839
rect 19659 35300 19701 35309
rect 19659 35260 19660 35300
rect 19700 35260 19701 35300
rect 19659 35251 19701 35260
rect 19756 35300 19796 35309
rect 19796 35260 19892 35300
rect 19756 35251 19796 35260
rect 19467 34712 19509 34721
rect 19467 34672 19468 34712
rect 19508 34672 19509 34712
rect 19467 34663 19509 34672
rect 19468 34376 19508 34663
rect 19564 34637 19604 35171
rect 19755 35132 19797 35141
rect 19755 35092 19756 35132
rect 19796 35092 19797 35132
rect 19755 35083 19797 35092
rect 19563 34628 19605 34637
rect 19563 34588 19564 34628
rect 19604 34588 19605 34628
rect 19563 34579 19605 34588
rect 19756 34628 19796 35083
rect 19756 34579 19796 34588
rect 19564 34376 19604 34385
rect 19468 34336 19564 34376
rect 19564 33713 19604 34336
rect 19563 33704 19605 33713
rect 19563 33664 19564 33704
rect 19604 33664 19605 33704
rect 19563 33655 19605 33664
rect 19564 33570 19604 33655
rect 19756 33452 19796 33461
rect 19564 33412 19756 33452
rect 19468 32864 19508 32873
rect 19564 32864 19604 33412
rect 19756 33403 19796 33412
rect 19852 33284 19892 35260
rect 19948 35225 19988 35848
rect 20140 35729 20180 35814
rect 20139 35720 20181 35729
rect 20139 35680 20140 35720
rect 20180 35680 20181 35720
rect 20139 35671 20181 35680
rect 20048 35552 20416 35561
rect 20088 35512 20130 35552
rect 20170 35512 20212 35552
rect 20252 35512 20294 35552
rect 20334 35512 20376 35552
rect 20048 35503 20416 35512
rect 20139 35384 20181 35393
rect 20139 35344 20140 35384
rect 20180 35344 20181 35384
rect 20139 35335 20181 35344
rect 20043 35300 20085 35309
rect 20043 35260 20044 35300
rect 20084 35260 20085 35300
rect 20043 35251 20085 35260
rect 19947 35216 19989 35225
rect 19947 35176 19948 35216
rect 19988 35176 19989 35216
rect 19947 35167 19989 35176
rect 20044 35216 20084 35251
rect 20140 35237 20180 35335
rect 20140 35188 20180 35197
rect 20236 35216 20276 35225
rect 19948 35082 19988 35167
rect 20044 35165 20084 35176
rect 20236 35057 20276 35176
rect 20043 35048 20085 35057
rect 20043 35008 20044 35048
rect 20084 35008 20085 35048
rect 20043 34999 20085 35008
rect 20235 35048 20277 35057
rect 20235 35008 20236 35048
rect 20276 35008 20277 35048
rect 20235 34999 20277 35008
rect 19947 34460 19989 34469
rect 19947 34420 19948 34460
rect 19988 34420 19989 34460
rect 19947 34411 19989 34420
rect 19948 34326 19988 34411
rect 20044 34208 20084 34999
rect 20140 34217 20180 34302
rect 19948 34168 20084 34208
rect 20139 34208 20181 34217
rect 20139 34168 20140 34208
rect 20180 34168 20181 34208
rect 19948 33788 19988 34168
rect 20139 34159 20181 34168
rect 20048 34040 20416 34049
rect 20088 34000 20130 34040
rect 20170 34000 20212 34040
rect 20252 34000 20294 34040
rect 20334 34000 20376 34040
rect 20048 33991 20416 34000
rect 19948 33748 20084 33788
rect 19948 33620 19988 33629
rect 19948 33377 19988 33580
rect 19947 33368 19989 33377
rect 19947 33328 19948 33368
rect 19988 33328 19989 33368
rect 19947 33319 19989 33328
rect 19756 33244 19892 33284
rect 19659 33032 19701 33041
rect 19659 32992 19660 33032
rect 19700 32992 19701 33032
rect 19659 32983 19701 32992
rect 19508 32824 19604 32864
rect 19468 32815 19508 32824
rect 19084 32236 19412 32276
rect 19084 32192 19124 32236
rect 19084 32143 19124 32152
rect 19276 32108 19316 32119
rect 19276 32033 19316 32068
rect 18219 32024 18261 32033
rect 18219 31984 18220 32024
rect 18260 31984 18261 32024
rect 18219 31975 18261 31984
rect 19275 32024 19317 32033
rect 19275 31984 19276 32024
rect 19316 31984 19317 32024
rect 19275 31975 19317 31984
rect 18808 31772 19176 31781
rect 18848 31732 18890 31772
rect 18930 31732 18972 31772
rect 19012 31732 19054 31772
rect 19094 31732 19136 31772
rect 18808 31723 19176 31732
rect 19372 31604 19412 32236
rect 19660 32192 19700 32983
rect 19756 32864 19796 33244
rect 20044 33200 20084 33748
rect 20140 33452 20180 33461
rect 20140 33209 20180 33412
rect 19756 32815 19796 32824
rect 19852 33160 20084 33200
rect 20139 33200 20181 33209
rect 20139 33160 20140 33200
rect 20180 33160 20181 33200
rect 19852 32864 19892 33160
rect 20139 33151 20181 33160
rect 19947 32948 19989 32957
rect 19947 32908 19948 32948
rect 19988 32908 19989 32948
rect 19947 32899 19989 32908
rect 19852 32815 19892 32824
rect 19948 32612 19988 32899
rect 20140 32705 20180 32749
rect 20139 32696 20181 32705
rect 20139 32656 20140 32696
rect 20180 32656 20181 32696
rect 20139 32654 20181 32656
rect 20139 32647 20140 32654
rect 19852 32572 19988 32612
rect 20180 32647 20181 32654
rect 20140 32605 20180 32614
rect 19852 32201 19892 32572
rect 20524 32537 20564 36436
rect 20620 33545 20660 37192
rect 20715 36224 20757 36233
rect 20715 36184 20716 36224
rect 20756 36184 20757 36224
rect 20715 36175 20757 36184
rect 20716 35888 20756 36175
rect 20812 36065 20852 38779
rect 20811 36056 20853 36065
rect 20811 36016 20812 36056
rect 20852 36016 20853 36056
rect 20811 36007 20853 36016
rect 20716 35848 20852 35888
rect 20715 34208 20757 34217
rect 20715 34168 20716 34208
rect 20756 34168 20757 34208
rect 20715 34159 20757 34168
rect 20619 33536 20661 33545
rect 20619 33496 20620 33536
rect 20660 33496 20661 33536
rect 20619 33487 20661 33496
rect 20619 33200 20661 33209
rect 20619 33160 20620 33200
rect 20660 33160 20661 33200
rect 20619 33151 20661 33160
rect 20048 32528 20416 32537
rect 20088 32488 20130 32528
rect 20170 32488 20212 32528
rect 20252 32488 20294 32528
rect 20334 32488 20376 32528
rect 20048 32479 20416 32488
rect 20523 32528 20565 32537
rect 20523 32488 20524 32528
rect 20564 32488 20565 32528
rect 20523 32479 20565 32488
rect 19468 32152 19700 32192
rect 19851 32192 19893 32201
rect 19851 32152 19852 32192
rect 19892 32152 19893 32192
rect 19468 32024 19508 32152
rect 19851 32143 19893 32152
rect 20043 32192 20085 32201
rect 20043 32152 20044 32192
rect 20084 32152 20085 32192
rect 20043 32143 20085 32152
rect 20044 32108 20084 32143
rect 19468 31975 19508 31984
rect 19660 32097 19700 32106
rect 20044 32057 20084 32068
rect 19660 31697 19700 32057
rect 19851 32024 19893 32033
rect 19851 31984 19852 32024
rect 19892 31984 19893 32024
rect 19851 31975 19893 31984
rect 19852 31890 19892 31975
rect 20236 31940 20276 31949
rect 19659 31688 19701 31697
rect 19659 31648 19660 31688
rect 19700 31648 19701 31688
rect 19659 31639 19701 31648
rect 19372 31564 19604 31604
rect 19275 31520 19317 31529
rect 19275 31480 19276 31520
rect 19316 31480 19317 31520
rect 18316 31445 18356 31476
rect 19275 31471 19317 31480
rect 18315 31436 18357 31445
rect 18315 31396 18316 31436
rect 18356 31396 18357 31436
rect 18315 31387 18357 31396
rect 19179 31436 19221 31445
rect 19179 31396 19180 31436
rect 19220 31396 19221 31436
rect 19179 31387 19221 31396
rect 18123 31352 18165 31361
rect 18123 31312 18124 31352
rect 18164 31312 18165 31352
rect 18123 31303 18165 31312
rect 18220 31352 18260 31363
rect 18124 31218 18164 31303
rect 18220 31277 18260 31312
rect 18316 31352 18356 31387
rect 18219 31268 18261 31277
rect 18219 31228 18220 31268
rect 18260 31228 18261 31268
rect 18219 31219 18261 31228
rect 18316 31016 18356 31312
rect 18507 31352 18549 31361
rect 18700 31352 18740 31361
rect 18507 31312 18508 31352
rect 18548 31312 18549 31352
rect 18507 31303 18549 31312
rect 18604 31312 18700 31352
rect 18508 31184 18548 31303
rect 18508 31135 18548 31144
rect 18316 30976 18452 31016
rect 18315 30848 18357 30857
rect 18315 30808 18316 30848
rect 18356 30808 18357 30848
rect 18315 30799 18357 30808
rect 17452 28456 17588 28496
rect 17740 29800 18068 29840
rect 17452 26144 17492 28456
rect 17547 28328 17589 28337
rect 17547 28288 17548 28328
rect 17588 28288 17589 28328
rect 17547 28279 17589 28288
rect 17548 28194 17588 28279
rect 17548 27656 17588 27665
rect 17548 27329 17588 27616
rect 17547 27320 17589 27329
rect 17547 27280 17548 27320
rect 17588 27280 17589 27320
rect 17547 27271 17589 27280
rect 17548 26144 17588 26153
rect 17452 26104 17548 26144
rect 17356 26020 17492 26060
rect 17355 25892 17397 25901
rect 17355 25852 17356 25892
rect 17396 25852 17397 25892
rect 17355 25843 17397 25852
rect 17356 25758 17396 25843
rect 17355 25640 17397 25649
rect 17355 25600 17356 25640
rect 17396 25600 17397 25640
rect 17355 25591 17397 25600
rect 17356 25388 17396 25591
rect 17259 24548 17301 24557
rect 17259 24508 17260 24548
rect 17300 24508 17301 24548
rect 17259 24499 17301 24508
rect 17356 24221 17396 25348
rect 17452 25304 17492 26020
rect 17355 24212 17397 24221
rect 17355 24172 17356 24212
rect 17396 24172 17397 24212
rect 17355 24163 17397 24172
rect 17452 24053 17492 25264
rect 17451 24044 17493 24053
rect 17451 24004 17452 24044
rect 17492 24004 17493 24044
rect 17451 23995 17493 24004
rect 17548 23969 17588 26104
rect 17547 23960 17589 23969
rect 17547 23920 17548 23960
rect 17588 23920 17589 23960
rect 17547 23911 17589 23920
rect 17356 23792 17396 23801
rect 17260 23752 17356 23792
rect 17164 23624 17204 23633
rect 17164 23129 17204 23584
rect 17260 23213 17300 23752
rect 17356 23743 17396 23752
rect 17452 23792 17492 23801
rect 17356 23288 17396 23297
rect 17452 23288 17492 23752
rect 17548 23792 17588 23801
rect 17548 23297 17588 23752
rect 17643 23624 17685 23633
rect 17643 23584 17644 23624
rect 17684 23584 17685 23624
rect 17643 23575 17685 23584
rect 17644 23490 17684 23575
rect 17396 23248 17492 23288
rect 17547 23288 17589 23297
rect 17547 23248 17548 23288
rect 17588 23248 17589 23288
rect 17356 23239 17396 23248
rect 17547 23239 17589 23248
rect 17259 23204 17301 23213
rect 17259 23164 17260 23204
rect 17300 23164 17301 23204
rect 17259 23155 17301 23164
rect 17163 23120 17205 23129
rect 17163 23080 17164 23120
rect 17204 23080 17205 23120
rect 17163 23071 17205 23080
rect 17164 22952 17204 22961
rect 17260 22952 17300 23155
rect 17548 23120 17588 23129
rect 17204 22912 17300 22952
rect 17355 22952 17397 22961
rect 17355 22912 17356 22952
rect 17396 22912 17397 22952
rect 17164 22903 17204 22912
rect 17355 22903 17397 22912
rect 17164 22280 17204 22289
rect 17164 21701 17204 22240
rect 17259 22280 17301 22289
rect 17259 22240 17260 22280
rect 17300 22240 17301 22280
rect 17259 22231 17301 22240
rect 17163 21692 17205 21701
rect 17163 21652 17164 21692
rect 17204 21652 17205 21692
rect 17163 21643 17205 21652
rect 17163 19592 17205 19601
rect 17163 19552 17164 19592
rect 17204 19552 17205 19592
rect 17163 19543 17205 19552
rect 17164 18593 17204 19543
rect 17260 18845 17300 22231
rect 17356 21608 17396 22903
rect 17548 22877 17588 23080
rect 17643 23120 17685 23129
rect 17643 23080 17644 23120
rect 17684 23080 17685 23120
rect 17643 23071 17685 23080
rect 17547 22868 17589 22877
rect 17547 22828 17548 22868
rect 17588 22828 17589 22868
rect 17547 22819 17589 22828
rect 17644 22793 17684 23071
rect 17643 22784 17685 22793
rect 17643 22744 17644 22784
rect 17684 22744 17685 22784
rect 17643 22735 17685 22744
rect 17740 22532 17780 29800
rect 17835 29672 17877 29681
rect 17835 29632 17836 29672
rect 17876 29632 17877 29672
rect 17835 29623 17877 29632
rect 17836 29177 17876 29623
rect 18027 29588 18069 29597
rect 18027 29548 18028 29588
rect 18068 29548 18069 29588
rect 18027 29539 18069 29548
rect 18028 29336 18068 29539
rect 18028 29287 18068 29296
rect 18316 29336 18356 30799
rect 18412 30666 18452 30976
rect 18604 30932 18644 31312
rect 18700 31303 18740 31312
rect 18796 31352 18836 31361
rect 18412 30101 18452 30626
rect 18508 30892 18644 30932
rect 18411 30092 18453 30101
rect 18411 30052 18412 30092
rect 18452 30052 18453 30092
rect 18411 30043 18453 30052
rect 18411 29588 18453 29597
rect 18411 29548 18412 29588
rect 18452 29548 18453 29588
rect 18411 29539 18453 29548
rect 18316 29287 18356 29296
rect 17835 29168 17877 29177
rect 18220 29168 18260 29177
rect 17835 29128 17836 29168
rect 17876 29128 17877 29168
rect 17835 29119 17877 29128
rect 17932 29128 18220 29168
rect 17836 29034 17876 29119
rect 17836 27665 17876 27750
rect 17835 27656 17877 27665
rect 17835 27616 17836 27656
rect 17876 27616 17877 27656
rect 17835 27607 17877 27616
rect 17836 27488 17876 27497
rect 17932 27488 17972 29128
rect 18220 29119 18260 29128
rect 18412 29168 18452 29539
rect 18508 29345 18548 30892
rect 18796 30857 18836 31312
rect 18892 31352 18932 31361
rect 18795 30848 18837 30857
rect 18795 30808 18796 30848
rect 18836 30808 18837 30848
rect 18795 30799 18837 30808
rect 18604 30764 18644 30773
rect 18507 29336 18549 29345
rect 18507 29296 18508 29336
rect 18548 29296 18549 29336
rect 18507 29287 18549 29296
rect 18604 29177 18644 30724
rect 18796 30680 18836 30689
rect 18700 30640 18796 30680
rect 18700 30008 18740 30640
rect 18796 30631 18836 30640
rect 18892 30521 18932 31312
rect 19180 31352 19220 31387
rect 19180 31301 19220 31312
rect 19276 31352 19316 31471
rect 19372 31361 19412 31446
rect 19276 31303 19316 31312
rect 19371 31352 19413 31361
rect 19371 31312 19372 31352
rect 19412 31312 19413 31352
rect 19371 31303 19413 31312
rect 18987 31184 19029 31193
rect 18987 31144 18988 31184
rect 19028 31144 19029 31184
rect 18987 31135 19029 31144
rect 19468 31184 19508 31193
rect 18988 31050 19028 31135
rect 18891 30512 18933 30521
rect 18891 30472 18892 30512
rect 18932 30472 18933 30512
rect 18891 30463 18933 30472
rect 18808 30260 19176 30269
rect 18848 30220 18890 30260
rect 18930 30220 18972 30260
rect 19012 30220 19054 30260
rect 19094 30220 19136 30260
rect 18808 30211 19176 30220
rect 19468 30101 19508 31144
rect 18891 30092 18933 30101
rect 18891 30052 18892 30092
rect 18932 30052 18933 30092
rect 18891 30043 18933 30052
rect 19467 30092 19509 30101
rect 19467 30052 19468 30092
rect 19508 30052 19509 30092
rect 19467 30043 19509 30052
rect 18700 29968 18836 30008
rect 18699 29840 18741 29849
rect 18699 29800 18700 29840
rect 18740 29800 18741 29840
rect 18699 29791 18741 29800
rect 18700 29706 18740 29791
rect 18699 29420 18741 29429
rect 18699 29380 18700 29420
rect 18740 29380 18741 29420
rect 18699 29371 18741 29380
rect 18412 29119 18452 29128
rect 18498 29168 18548 29177
rect 18498 29128 18499 29168
rect 18498 29119 18548 29128
rect 18603 29168 18645 29177
rect 18603 29128 18604 29168
rect 18644 29128 18645 29168
rect 18603 29119 18645 29128
rect 18508 29000 18548 29119
rect 18700 29084 18740 29371
rect 18700 29035 18740 29044
rect 18412 28960 18548 29000
rect 18603 29000 18645 29009
rect 18603 28960 18604 29000
rect 18644 28960 18645 29000
rect 18028 28916 18068 28925
rect 18028 28342 18068 28876
rect 18068 28302 18164 28342
rect 18028 28293 18068 28302
rect 18124 27665 18164 28302
rect 18219 28160 18261 28169
rect 18219 28120 18220 28160
rect 18260 28120 18261 28160
rect 18219 28111 18261 28120
rect 18220 28026 18260 28111
rect 18219 27908 18261 27917
rect 18219 27868 18220 27908
rect 18260 27868 18261 27908
rect 18219 27859 18261 27868
rect 18123 27656 18165 27665
rect 18123 27616 18124 27656
rect 18164 27616 18165 27656
rect 18123 27607 18165 27616
rect 18220 27656 18260 27859
rect 18124 27522 18164 27607
rect 17876 27448 17972 27488
rect 17836 27439 17876 27448
rect 18027 27068 18069 27077
rect 18027 27028 18028 27068
rect 18068 27028 18069 27068
rect 18027 27019 18069 27028
rect 18028 26489 18068 27019
rect 18123 26984 18165 26993
rect 18123 26944 18124 26984
rect 18164 26944 18165 26984
rect 18123 26935 18165 26944
rect 18027 26480 18069 26489
rect 18027 26440 18028 26480
rect 18068 26440 18069 26480
rect 18027 26431 18069 26440
rect 17835 25976 17877 25985
rect 17835 25936 17836 25976
rect 17876 25936 17877 25976
rect 17835 25927 17877 25936
rect 17836 24632 17876 25927
rect 17931 25304 17973 25313
rect 17931 25264 17932 25304
rect 17972 25264 17973 25304
rect 17931 25255 17973 25264
rect 17932 25170 17972 25255
rect 18027 25220 18069 25229
rect 18027 25180 18028 25220
rect 18068 25180 18069 25220
rect 18027 25171 18069 25180
rect 18028 24800 18068 25171
rect 18028 24751 18068 24760
rect 17836 24583 17876 24592
rect 18124 23465 18164 26935
rect 18123 23456 18165 23465
rect 18123 23416 18124 23456
rect 18164 23416 18165 23456
rect 18123 23407 18165 23416
rect 17835 23372 17877 23381
rect 17835 23332 17836 23372
rect 17876 23332 17877 23372
rect 17835 23323 17877 23332
rect 17836 23120 17876 23323
rect 18123 23288 18165 23297
rect 18123 23248 18124 23288
rect 18164 23248 18165 23288
rect 18123 23239 18165 23248
rect 17931 23204 17973 23213
rect 17931 23164 17932 23204
rect 17972 23164 17973 23204
rect 17931 23155 17973 23164
rect 17836 23071 17876 23080
rect 17932 23120 17972 23155
rect 18124 23154 18164 23239
rect 17932 23069 17972 23080
rect 18028 23120 18068 23129
rect 18028 22952 18068 23080
rect 18220 23036 18260 27616
rect 18315 27656 18357 27665
rect 18315 27616 18316 27656
rect 18356 27616 18357 27656
rect 18315 27607 18357 27616
rect 18316 27522 18356 27607
rect 18412 26993 18452 28960
rect 18603 28951 18645 28960
rect 18508 28328 18548 28337
rect 18604 28328 18644 28951
rect 18796 28916 18836 29968
rect 18892 29958 18932 30043
rect 19564 29924 19604 31564
rect 20236 31529 20276 31900
rect 20235 31520 20277 31529
rect 20235 31480 20236 31520
rect 20276 31480 20277 31520
rect 20235 31471 20277 31480
rect 19660 31436 19700 31445
rect 19660 31025 19700 31396
rect 19755 31436 19797 31445
rect 19755 31396 19756 31436
rect 19796 31396 19797 31436
rect 19755 31387 19797 31396
rect 20043 31436 20085 31445
rect 20043 31396 20044 31436
rect 20084 31396 20085 31436
rect 20043 31387 20085 31396
rect 19659 31016 19701 31025
rect 19659 30976 19660 31016
rect 19700 30976 19701 31016
rect 19659 30967 19701 30976
rect 19756 30437 19796 31387
rect 20044 31302 20084 31387
rect 19852 31184 19892 31193
rect 19755 30428 19797 30437
rect 19755 30388 19756 30428
rect 19796 30388 19797 30428
rect 19755 30379 19797 30388
rect 19659 30092 19701 30101
rect 19659 30052 19660 30092
rect 19700 30052 19701 30092
rect 19659 30043 19701 30052
rect 19276 29884 19604 29924
rect 19276 29840 19316 29884
rect 19660 29840 19700 30043
rect 19276 29791 19316 29800
rect 19564 29800 19700 29840
rect 19755 29840 19797 29849
rect 19755 29800 19756 29840
rect 19796 29800 19797 29840
rect 19179 29756 19221 29765
rect 19179 29716 19180 29756
rect 19220 29716 19221 29756
rect 19179 29707 19221 29716
rect 18891 29336 18933 29345
rect 18891 29296 18892 29336
rect 18932 29296 18933 29336
rect 18891 29287 18933 29296
rect 18892 29202 18932 29287
rect 18987 29252 19029 29261
rect 18987 29212 18988 29252
rect 19028 29212 19029 29252
rect 18987 29203 19029 29212
rect 18988 29093 19028 29203
rect 19180 29168 19220 29707
rect 19564 29252 19604 29800
rect 19755 29791 19797 29800
rect 19564 29203 19604 29212
rect 19660 29672 19700 29681
rect 19180 29119 19220 29128
rect 19467 29168 19509 29177
rect 19467 29128 19468 29168
rect 19508 29128 19509 29168
rect 19467 29119 19509 29128
rect 18987 29084 19029 29093
rect 18987 29044 18988 29084
rect 19028 29044 19029 29084
rect 18987 29035 19029 29044
rect 19468 29034 19508 29119
rect 19275 29000 19317 29009
rect 19275 28960 19276 29000
rect 19316 28960 19317 29000
rect 19275 28951 19317 28960
rect 18548 28288 18644 28328
rect 18700 28876 18836 28916
rect 18508 28279 18548 28288
rect 18507 27824 18549 27833
rect 18507 27784 18508 27824
rect 18548 27784 18549 27824
rect 18507 27775 18549 27784
rect 18508 27690 18548 27775
rect 18700 27572 18740 28876
rect 18808 28748 19176 28757
rect 18848 28708 18890 28748
rect 18930 28708 18972 28748
rect 19012 28708 19054 28748
rect 19094 28708 19136 28748
rect 18808 28699 19176 28708
rect 19179 27656 19221 27665
rect 19179 27616 19180 27656
rect 19220 27616 19221 27656
rect 19179 27607 19221 27616
rect 18700 27161 18740 27532
rect 19180 27522 19220 27607
rect 18891 27488 18933 27497
rect 18891 27448 18892 27488
rect 18932 27448 18933 27488
rect 18891 27439 18933 27448
rect 18892 27354 18932 27439
rect 18808 27236 19176 27245
rect 18848 27196 18890 27236
rect 18930 27196 18972 27236
rect 19012 27196 19054 27236
rect 19094 27196 19136 27236
rect 18808 27187 19176 27196
rect 18699 27152 18741 27161
rect 18699 27112 18700 27152
rect 18740 27112 18741 27152
rect 18699 27103 18741 27112
rect 18411 26984 18453 26993
rect 18411 26944 18412 26984
rect 18452 26944 18453 26984
rect 18411 26935 18453 26944
rect 19276 26900 19316 28951
rect 19467 28160 19509 28169
rect 19467 28120 19468 28160
rect 19508 28120 19509 28160
rect 19467 28111 19509 28120
rect 19468 27656 19508 28111
rect 19563 27740 19605 27749
rect 19563 27700 19564 27740
rect 19604 27700 19605 27740
rect 19563 27691 19605 27700
rect 19468 27607 19508 27616
rect 19564 27606 19604 27691
rect 19372 26900 19412 26909
rect 19276 26860 19372 26900
rect 19372 26851 19412 26860
rect 18411 26816 18453 26825
rect 18316 26776 18412 26816
rect 18452 26776 18453 26816
rect 18316 24053 18356 26776
rect 18411 26767 18453 26776
rect 18604 26816 18644 26825
rect 18795 26816 18837 26825
rect 18644 26776 18740 26816
rect 18604 26767 18644 26776
rect 18412 26682 18452 26767
rect 18508 26732 18548 26741
rect 18411 26312 18453 26321
rect 18411 26272 18412 26312
rect 18452 26272 18453 26312
rect 18411 26263 18453 26272
rect 18412 25318 18452 26263
rect 18412 25229 18452 25278
rect 18411 25220 18453 25229
rect 18411 25180 18412 25220
rect 18452 25180 18453 25220
rect 18411 25171 18453 25180
rect 18412 24968 18452 25171
rect 18508 25145 18548 26692
rect 18603 26480 18645 26489
rect 18603 26440 18604 26480
rect 18644 26440 18645 26480
rect 18603 26431 18645 26440
rect 18604 25220 18644 26431
rect 18700 25901 18740 26776
rect 18795 26776 18796 26816
rect 18836 26776 18837 26816
rect 18795 26767 18837 26776
rect 18892 26816 18932 26825
rect 18796 26682 18836 26767
rect 18892 26489 18932 26776
rect 18987 26816 19029 26825
rect 18987 26776 18988 26816
rect 19028 26776 19029 26816
rect 18987 26767 19029 26776
rect 18891 26480 18933 26489
rect 18891 26440 18892 26480
rect 18932 26440 18933 26480
rect 18891 26431 18933 26440
rect 18988 26312 19028 26767
rect 18988 26153 19028 26272
rect 19084 26648 19124 26657
rect 18796 26144 18836 26153
rect 18796 25985 18836 26104
rect 18987 26144 19029 26153
rect 18987 26104 18988 26144
rect 19028 26104 19029 26144
rect 18987 26095 19029 26104
rect 18795 25976 18837 25985
rect 18795 25936 18796 25976
rect 18836 25936 18837 25976
rect 18795 25927 18837 25936
rect 18699 25892 18741 25901
rect 18699 25852 18700 25892
rect 18740 25852 18741 25892
rect 19084 25892 19124 26608
rect 19563 26648 19605 26657
rect 19563 26608 19564 26648
rect 19604 26608 19605 26648
rect 19563 26599 19605 26608
rect 19564 26514 19604 26599
rect 19660 26396 19700 29632
rect 19756 28328 19796 29791
rect 19852 29597 19892 31144
rect 20236 31184 20276 31193
rect 20276 31144 20564 31184
rect 20236 31135 20276 31144
rect 20048 31016 20416 31025
rect 20088 30976 20130 31016
rect 20170 30976 20212 31016
rect 20252 30976 20294 31016
rect 20334 30976 20376 31016
rect 20048 30967 20416 30976
rect 20043 30680 20085 30689
rect 20043 30640 20044 30680
rect 20084 30640 20085 30680
rect 20043 30631 20085 30640
rect 20044 30546 20084 30631
rect 20236 30428 20276 30437
rect 20236 29765 20276 30388
rect 20235 29756 20277 29765
rect 20235 29716 20236 29756
rect 20276 29716 20277 29756
rect 20235 29707 20277 29716
rect 19851 29588 19893 29597
rect 19851 29548 19852 29588
rect 19892 29548 19893 29588
rect 19851 29539 19893 29548
rect 19947 29504 19989 29513
rect 19947 29464 19948 29504
rect 19988 29464 19989 29504
rect 19947 29455 19989 29464
rect 20048 29504 20416 29513
rect 20088 29464 20130 29504
rect 20170 29464 20212 29504
rect 20252 29464 20294 29504
rect 20334 29464 20376 29504
rect 20048 29455 20416 29464
rect 19948 29084 19988 29455
rect 20524 29261 20564 31144
rect 20620 30521 20660 33151
rect 20716 31025 20756 34159
rect 20715 31016 20757 31025
rect 20715 30976 20716 31016
rect 20756 30976 20757 31016
rect 20715 30967 20757 30976
rect 20619 30512 20661 30521
rect 20619 30472 20620 30512
rect 20660 30472 20661 30512
rect 20619 30463 20661 30472
rect 20619 29336 20661 29345
rect 20619 29296 20620 29336
rect 20660 29296 20661 29336
rect 20619 29287 20661 29296
rect 20523 29252 20565 29261
rect 20523 29212 20524 29252
rect 20564 29212 20565 29252
rect 20523 29203 20565 29212
rect 20044 29084 20084 29093
rect 19948 29044 20044 29084
rect 20044 29035 20084 29044
rect 20523 29084 20565 29093
rect 20523 29044 20524 29084
rect 20564 29044 20565 29084
rect 20523 29035 20565 29044
rect 19851 29000 19893 29009
rect 19851 28960 19852 29000
rect 19892 28960 19893 29000
rect 19851 28951 19893 28960
rect 19852 28866 19892 28951
rect 20236 28916 20276 28925
rect 20236 28505 20276 28876
rect 20235 28496 20277 28505
rect 20235 28456 20236 28496
rect 20276 28456 20277 28496
rect 20235 28447 20277 28456
rect 19756 28279 19796 28288
rect 19948 28160 19988 28169
rect 19948 27665 19988 28120
rect 20048 27992 20416 28001
rect 20088 27952 20130 27992
rect 20170 27952 20212 27992
rect 20252 27952 20294 27992
rect 20334 27952 20376 27992
rect 20048 27943 20416 27952
rect 19947 27656 19989 27665
rect 19947 27616 19948 27656
rect 19988 27616 19989 27656
rect 19947 27607 19989 27616
rect 19851 27404 19893 27413
rect 19851 27364 19852 27404
rect 19892 27364 19893 27404
rect 19851 27355 19893 27364
rect 19852 27270 19892 27355
rect 19947 26984 19989 26993
rect 19947 26944 19948 26984
rect 19988 26944 19989 26984
rect 19947 26935 19989 26944
rect 19756 26900 19796 26909
rect 19756 26741 19796 26860
rect 19948 26850 19988 26935
rect 19755 26732 19797 26741
rect 19755 26692 19756 26732
rect 19796 26692 19797 26732
rect 19755 26683 19797 26692
rect 20048 26480 20416 26489
rect 20088 26440 20130 26480
rect 20170 26440 20212 26480
rect 20252 26440 20294 26480
rect 20334 26440 20376 26480
rect 20048 26431 20416 26440
rect 19660 26356 19988 26396
rect 19179 26312 19221 26321
rect 19179 26272 19180 26312
rect 19220 26272 19221 26312
rect 19179 26263 19221 26272
rect 19276 26272 19604 26312
rect 19180 26144 19220 26263
rect 19180 26095 19220 26104
rect 19276 26144 19316 26272
rect 19276 26095 19316 26104
rect 19371 26144 19413 26153
rect 19371 26104 19372 26144
rect 19412 26104 19413 26144
rect 19371 26095 19413 26104
rect 19468 26144 19508 26153
rect 19372 26010 19412 26095
rect 19084 25852 19316 25892
rect 18699 25843 18741 25852
rect 18700 25556 18740 25843
rect 18808 25724 19176 25733
rect 18848 25684 18890 25724
rect 18930 25684 18972 25724
rect 19012 25684 19054 25724
rect 19094 25684 19136 25724
rect 18808 25675 19176 25684
rect 19276 25556 19316 25852
rect 19371 25808 19413 25817
rect 19371 25768 19372 25808
rect 19412 25768 19413 25808
rect 19371 25759 19413 25768
rect 18700 25516 18836 25556
rect 18796 25388 18836 25516
rect 19084 25516 19316 25556
rect 18891 25388 18933 25397
rect 18796 25348 18892 25388
rect 18932 25348 18933 25388
rect 18891 25339 18933 25348
rect 18699 25304 18741 25313
rect 18699 25264 18700 25304
rect 18740 25264 18741 25304
rect 18699 25255 18741 25264
rect 18892 25304 18932 25339
rect 18604 25171 18644 25180
rect 18507 25136 18549 25145
rect 18507 25096 18508 25136
rect 18548 25096 18549 25136
rect 18507 25087 18549 25096
rect 18700 24968 18740 25255
rect 18892 25253 18932 25264
rect 18795 25136 18837 25145
rect 18795 25096 18796 25136
rect 18836 25096 18837 25136
rect 18795 25087 18837 25096
rect 18412 24928 18548 24968
rect 18508 24842 18548 24928
rect 18508 24793 18548 24802
rect 18604 24928 18740 24968
rect 18604 24632 18644 24928
rect 18700 24632 18740 24641
rect 18604 24592 18700 24632
rect 18700 24583 18740 24592
rect 18796 24632 18836 25087
rect 19084 25052 19124 25516
rect 19372 25472 19412 25759
rect 19276 25432 19412 25472
rect 19180 25304 19220 25315
rect 19180 25229 19220 25264
rect 19276 25304 19316 25432
rect 19468 25388 19508 26104
rect 19564 25556 19604 26272
rect 19659 26060 19701 26069
rect 19659 26020 19660 26060
rect 19700 26020 19701 26060
rect 19659 26011 19701 26020
rect 19660 25926 19700 26011
rect 19852 25892 19892 25901
rect 19852 25733 19892 25852
rect 19851 25724 19893 25733
rect 19851 25684 19852 25724
rect 19892 25684 19893 25724
rect 19851 25675 19893 25684
rect 19564 25507 19604 25516
rect 19276 25255 19316 25264
rect 19372 25348 19508 25388
rect 19659 25388 19701 25397
rect 19659 25348 19660 25388
rect 19700 25348 19796 25388
rect 19179 25220 19221 25229
rect 19179 25180 19180 25220
rect 19220 25180 19221 25220
rect 19179 25171 19221 25180
rect 19084 25012 19316 25052
rect 19180 24641 19220 24726
rect 18796 24583 18836 24592
rect 19179 24632 19221 24641
rect 19179 24592 19180 24632
rect 19220 24592 19221 24632
rect 19179 24583 19221 24592
rect 19276 24632 19316 25012
rect 19276 24583 19316 24592
rect 19372 24632 19412 25348
rect 19659 25339 19701 25348
rect 19756 25304 19796 25348
rect 19756 25255 19796 25264
rect 19852 25304 19892 25313
rect 19755 25136 19797 25145
rect 19755 25096 19756 25136
rect 19796 25096 19797 25136
rect 19755 25087 19797 25096
rect 19372 24583 19412 24592
rect 19468 24632 19508 24641
rect 18603 24464 18645 24473
rect 18603 24424 18604 24464
rect 18644 24424 18645 24464
rect 18603 24415 18645 24424
rect 18988 24464 19028 24473
rect 19468 24464 19508 24592
rect 19028 24424 19508 24464
rect 19660 24548 19700 24557
rect 18988 24415 19028 24424
rect 18315 24044 18357 24053
rect 18315 24004 18316 24044
rect 18356 24004 18357 24044
rect 18315 23995 18357 24004
rect 17932 22912 18068 22952
rect 18124 22996 18260 23036
rect 18316 23792 18356 23801
rect 17932 22793 17972 22912
rect 17931 22784 17973 22793
rect 17931 22744 17932 22784
rect 17972 22744 17973 22784
rect 17931 22735 17973 22744
rect 18027 22532 18069 22541
rect 17740 22492 17876 22532
rect 17740 22289 17780 22374
rect 17644 22280 17684 22289
rect 17644 22196 17684 22240
rect 17739 22280 17781 22289
rect 17739 22240 17740 22280
rect 17780 22240 17781 22280
rect 17739 22231 17781 22240
rect 17356 21113 17396 21568
rect 17452 22156 17684 22196
rect 17355 21104 17397 21113
rect 17355 21064 17356 21104
rect 17396 21064 17397 21104
rect 17355 21055 17397 21064
rect 17356 20768 17396 20777
rect 17356 20021 17396 20728
rect 17452 20768 17492 22156
rect 17836 22112 17876 22492
rect 18027 22492 18028 22532
rect 18068 22492 18069 22532
rect 18027 22483 18069 22492
rect 17931 22280 17973 22289
rect 17931 22240 17932 22280
rect 17972 22240 17973 22280
rect 17931 22231 17973 22240
rect 17644 22072 17876 22112
rect 17547 21692 17589 21701
rect 17547 21652 17548 21692
rect 17588 21652 17589 21692
rect 17547 21643 17589 21652
rect 17548 21558 17588 21643
rect 17452 20441 17492 20728
rect 17451 20432 17493 20441
rect 17451 20392 17452 20432
rect 17492 20392 17493 20432
rect 17451 20383 17493 20392
rect 17355 20012 17397 20021
rect 17355 19972 17356 20012
rect 17396 19972 17397 20012
rect 17355 19963 17397 19972
rect 17356 19256 17396 19267
rect 17356 19181 17396 19216
rect 17355 19172 17397 19181
rect 17355 19132 17356 19172
rect 17396 19132 17397 19172
rect 17355 19123 17397 19132
rect 17259 18836 17301 18845
rect 17259 18796 17260 18836
rect 17300 18796 17301 18836
rect 17259 18787 17301 18796
rect 17163 18584 17205 18593
rect 17163 18544 17164 18584
rect 17204 18544 17205 18584
rect 17163 18535 17205 18544
rect 17164 18450 17204 18535
rect 17068 17872 17588 17912
rect 16972 17788 17396 17828
rect 16684 17200 16820 17240
rect 16876 17744 16916 17753
rect 16876 17240 16916 17704
rect 16972 17724 17012 17733
rect 16972 17669 17012 17684
rect 16971 17660 17013 17669
rect 16971 17620 16972 17660
rect 17012 17620 17013 17660
rect 16971 17611 17013 17620
rect 16972 17589 17012 17611
rect 16972 17240 17012 17249
rect 16876 17200 16972 17240
rect 16587 16232 16629 16241
rect 16587 16192 16588 16232
rect 16628 16192 16629 16232
rect 16587 16183 16629 16192
rect 16299 15560 16341 15569
rect 16299 15520 16300 15560
rect 16340 15520 16341 15560
rect 16299 15511 16341 15520
rect 16396 15560 16436 15569
rect 16300 15426 16340 15511
rect 16203 15392 16245 15401
rect 16203 15352 16204 15392
rect 16244 15352 16245 15392
rect 16203 15343 16245 15352
rect 16108 15184 16244 15224
rect 16107 14720 16149 14729
rect 16107 14680 16108 14720
rect 16148 14680 16149 14720
rect 16107 14671 16149 14680
rect 16108 13208 16148 14671
rect 16204 13880 16244 15184
rect 16396 15149 16436 15520
rect 16395 15140 16437 15149
rect 16395 15100 16396 15140
rect 16436 15100 16437 15140
rect 16395 15091 16437 15100
rect 16299 15056 16341 15065
rect 16299 15016 16300 15056
rect 16340 15016 16341 15056
rect 16299 15007 16341 15016
rect 16300 14048 16340 15007
rect 16684 14813 16724 17200
rect 16972 17191 17012 17200
rect 16779 17072 16821 17081
rect 16779 17032 16780 17072
rect 16820 17032 16821 17072
rect 16779 17023 16821 17032
rect 16780 16938 16820 17023
rect 16779 16232 16821 16241
rect 17068 16232 17108 17788
rect 17356 17744 17396 17788
rect 17356 17695 17396 17704
rect 17451 17744 17493 17753
rect 17451 17704 17452 17744
rect 17492 17704 17493 17744
rect 17451 17695 17493 17704
rect 17259 17660 17301 17669
rect 17259 17620 17260 17660
rect 17300 17620 17301 17660
rect 17259 17611 17301 17620
rect 16779 16192 16780 16232
rect 16820 16192 16821 16232
rect 16779 16183 16821 16192
rect 16876 16192 17108 16232
rect 16780 16098 16820 16183
rect 16876 15896 16916 16192
rect 17164 16148 17204 16157
rect 16780 15856 16916 15896
rect 16972 16064 17012 16073
rect 16780 15560 16820 15856
rect 16972 15569 17012 16024
rect 17164 15569 17204 16108
rect 16683 14804 16725 14813
rect 16683 14764 16684 14804
rect 16724 14764 16725 14804
rect 16683 14755 16725 14764
rect 16491 14552 16533 14561
rect 16491 14512 16492 14552
rect 16532 14512 16533 14552
rect 16491 14503 16533 14512
rect 16300 13999 16340 14008
rect 16204 13840 16340 13880
rect 16204 13208 16244 13217
rect 16108 13168 16204 13208
rect 15956 12496 16052 12536
rect 15819 11780 15861 11789
rect 15819 11740 15820 11780
rect 15860 11740 15861 11780
rect 15819 11731 15861 11740
rect 15820 11696 15860 11731
rect 15820 11645 15860 11656
rect 15723 11528 15765 11537
rect 15723 11488 15724 11528
rect 15764 11488 15765 11528
rect 15723 11479 15765 11488
rect 15628 11320 15764 11360
rect 15531 10940 15573 10949
rect 15531 10900 15532 10940
rect 15572 10900 15573 10940
rect 15531 10891 15573 10900
rect 15532 10184 15572 10193
rect 15436 10144 15532 10184
rect 15436 8849 15476 10144
rect 15532 10135 15572 10144
rect 15628 10184 15668 10193
rect 15628 9773 15668 10144
rect 15724 9857 15764 11320
rect 15820 11010 15860 11019
rect 15723 9848 15765 9857
rect 15723 9808 15724 9848
rect 15764 9808 15765 9848
rect 15723 9799 15765 9808
rect 15627 9764 15669 9773
rect 15627 9724 15628 9764
rect 15668 9724 15669 9764
rect 15627 9715 15669 9724
rect 15532 9512 15572 9521
rect 15532 9353 15572 9472
rect 15531 9344 15573 9353
rect 15531 9304 15532 9344
rect 15572 9304 15573 9344
rect 15531 9295 15573 9304
rect 15531 9008 15573 9017
rect 15531 8968 15532 9008
rect 15572 8968 15573 9008
rect 15531 8959 15573 8968
rect 15435 8840 15477 8849
rect 15435 8800 15436 8840
rect 15476 8800 15477 8840
rect 15435 8791 15477 8800
rect 15339 8420 15381 8429
rect 15339 8380 15340 8420
rect 15380 8380 15381 8420
rect 15339 8371 15381 8380
rect 15051 8000 15093 8009
rect 15051 7960 15052 8000
rect 15092 7960 15093 8000
rect 15051 7951 15093 7960
rect 15243 8000 15285 8009
rect 15243 7960 15244 8000
rect 15284 7960 15285 8000
rect 15243 7951 15285 7960
rect 15436 8000 15476 8009
rect 15052 7244 15092 7951
rect 15243 7748 15285 7757
rect 15243 7708 15244 7748
rect 15284 7708 15285 7748
rect 15243 7699 15285 7708
rect 15244 7614 15284 7699
rect 15436 7673 15476 7960
rect 15435 7664 15477 7673
rect 15435 7624 15436 7664
rect 15476 7624 15477 7664
rect 15435 7615 15477 7624
rect 15532 7412 15572 8959
rect 15628 8924 15668 9715
rect 15724 9680 15764 9689
rect 15820 9680 15860 10970
rect 15764 9640 15860 9680
rect 15724 9631 15764 9640
rect 15916 9512 15956 12496
rect 16204 11705 16244 13168
rect 16203 11696 16245 11705
rect 16203 11656 16204 11696
rect 16244 11656 16245 11696
rect 16203 11647 16245 11656
rect 16203 11528 16245 11537
rect 16203 11488 16204 11528
rect 16244 11488 16245 11528
rect 16203 11479 16245 11488
rect 16011 11276 16053 11285
rect 16011 11236 16012 11276
rect 16052 11236 16053 11276
rect 16011 11227 16053 11236
rect 16012 11192 16052 11227
rect 16012 11141 16052 11152
rect 16107 10940 16149 10949
rect 16107 10900 16108 10940
rect 16148 10900 16149 10940
rect 16107 10891 16149 10900
rect 16011 10268 16053 10277
rect 16011 10228 16012 10268
rect 16052 10228 16053 10268
rect 16011 10219 16053 10228
rect 16108 10268 16148 10891
rect 16204 10529 16244 11479
rect 16203 10520 16245 10529
rect 16203 10480 16204 10520
rect 16244 10480 16245 10520
rect 16203 10471 16245 10480
rect 16108 10219 16148 10228
rect 16012 10134 16052 10219
rect 16011 9932 16053 9941
rect 16011 9892 16012 9932
rect 16052 9892 16053 9932
rect 16011 9883 16053 9892
rect 16012 9521 16052 9883
rect 15820 9472 15956 9512
rect 16011 9512 16053 9521
rect 16011 9472 16012 9512
rect 16052 9472 16053 9512
rect 15628 8884 15764 8924
rect 15627 8756 15669 8765
rect 15627 8716 15628 8756
rect 15668 8716 15669 8756
rect 15627 8707 15669 8716
rect 15724 8756 15764 8884
rect 15820 8849 15860 9472
rect 16011 9463 16053 9472
rect 15915 9344 15957 9353
rect 15915 9304 15916 9344
rect 15956 9304 15957 9344
rect 15915 9295 15957 9304
rect 15819 8840 15861 8849
rect 15819 8800 15820 8840
rect 15860 8800 15861 8840
rect 15819 8791 15861 8800
rect 15628 8622 15668 8707
rect 15052 7195 15092 7204
rect 15244 7372 15572 7412
rect 15148 7160 15188 7171
rect 15148 7085 15188 7120
rect 15147 7076 15189 7085
rect 15147 7036 15148 7076
rect 15188 7036 15189 7076
rect 15147 7027 15189 7036
rect 15244 5816 15284 7372
rect 15724 7328 15764 8716
rect 15819 8000 15861 8009
rect 15819 7960 15820 8000
rect 15860 7960 15861 8000
rect 15819 7951 15861 7960
rect 15148 5776 15284 5816
rect 15340 7288 15764 7328
rect 14668 4339 14708 4348
rect 14860 4516 14996 4556
rect 15052 5060 15092 5069
rect 14763 3716 14805 3725
rect 14763 3676 14764 3716
rect 14804 3676 14805 3716
rect 14763 3667 14805 3676
rect 14764 3464 14804 3667
rect 14860 3464 14900 4516
rect 15052 4397 15092 5020
rect 15148 4976 15188 5776
rect 15244 5648 15284 5657
rect 15244 5489 15284 5608
rect 15243 5480 15285 5489
rect 15243 5440 15244 5480
rect 15284 5440 15285 5480
rect 15243 5431 15285 5440
rect 15244 4976 15284 4985
rect 15148 4936 15244 4976
rect 15244 4927 15284 4936
rect 15147 4556 15189 4565
rect 15147 4516 15148 4556
rect 15188 4516 15189 4556
rect 15147 4507 15189 4516
rect 15051 4388 15093 4397
rect 15051 4348 15052 4388
rect 15092 4348 15093 4388
rect 15051 4339 15093 4348
rect 15148 4220 15188 4507
rect 15340 4304 15380 7288
rect 15820 7244 15860 7951
rect 15916 7925 15956 9295
rect 16012 9017 16052 9463
rect 16107 9428 16149 9437
rect 16107 9388 16108 9428
rect 16148 9388 16149 9428
rect 16107 9379 16149 9388
rect 16011 9008 16053 9017
rect 16011 8968 16012 9008
rect 16052 8968 16053 9008
rect 16011 8959 16053 8968
rect 16108 8849 16148 9379
rect 16107 8840 16149 8849
rect 16107 8800 16108 8840
rect 16148 8800 16149 8840
rect 16107 8791 16149 8800
rect 16204 8672 16244 10471
rect 15915 7916 15957 7925
rect 15915 7876 15916 7916
rect 15956 7876 15957 7916
rect 15915 7867 15957 7876
rect 15532 7204 15860 7244
rect 15435 7160 15477 7169
rect 15435 7120 15436 7160
rect 15476 7120 15477 7160
rect 15435 7111 15477 7120
rect 15532 7160 15572 7204
rect 16012 7169 16052 7254
rect 16011 7160 16053 7169
rect 15532 7111 15572 7120
rect 15628 7140 15668 7149
rect 15436 5900 15476 7111
rect 16011 7120 16012 7160
rect 16052 7120 16053 7160
rect 16011 7111 16053 7120
rect 16108 7160 16148 7169
rect 15628 6665 15668 7100
rect 16108 6992 16148 7120
rect 16204 7076 16244 8632
rect 16204 7036 16247 7076
rect 16207 6992 16247 7036
rect 16012 6952 16148 6992
rect 16191 6952 16247 6992
rect 15627 6656 15669 6665
rect 15627 6616 15628 6656
rect 15668 6616 15669 6656
rect 15627 6607 15669 6616
rect 15820 6488 15860 6497
rect 15820 6245 15860 6448
rect 15819 6236 15861 6245
rect 15819 6196 15820 6236
rect 15860 6196 15861 6236
rect 15819 6187 15861 6196
rect 15436 5851 15476 5860
rect 16012 5657 16052 6952
rect 16191 6908 16231 6952
rect 16108 6868 16231 6908
rect 16011 5648 16053 5657
rect 16011 5608 16012 5648
rect 16052 5608 16053 5648
rect 16011 5599 16053 5608
rect 15819 5564 15861 5573
rect 15819 5524 15820 5564
rect 15860 5524 15861 5564
rect 15819 5515 15861 5524
rect 15340 4264 15572 4304
rect 15052 4180 15188 4220
rect 15532 4220 15572 4264
rect 14956 4136 14996 4145
rect 14956 3632 14996 4096
rect 15052 4136 15092 4180
rect 15052 4087 15092 4096
rect 15435 4136 15477 4145
rect 15435 4096 15436 4136
rect 15476 4096 15477 4136
rect 15435 4087 15477 4096
rect 15436 4002 15476 4087
rect 15532 4061 15572 4180
rect 15531 4052 15573 4061
rect 15531 4012 15532 4052
rect 15572 4012 15573 4052
rect 15531 4003 15573 4012
rect 14956 3583 14996 3592
rect 14860 3424 15092 3464
rect 14764 3415 14804 3424
rect 14955 3296 14997 3305
rect 14955 3256 14956 3296
rect 14996 3256 14997 3296
rect 14955 3247 14997 3256
rect 14763 3212 14805 3221
rect 14763 3172 14764 3212
rect 14804 3172 14805 3212
rect 14763 3163 14805 3172
rect 14668 2465 14708 2550
rect 14667 2456 14709 2465
rect 14667 2416 14668 2456
rect 14708 2416 14709 2456
rect 14667 2407 14709 2416
rect 14572 2248 14708 2288
rect 14283 1868 14325 1877
rect 14283 1828 14284 1868
rect 14324 1828 14325 1868
rect 14283 1819 14325 1828
rect 14380 1868 14420 1877
rect 14284 1196 14324 1819
rect 14380 1709 14420 1828
rect 14379 1700 14421 1709
rect 14379 1660 14380 1700
rect 14420 1660 14421 1700
rect 14379 1651 14421 1660
rect 14571 1700 14613 1709
rect 14571 1660 14572 1700
rect 14612 1660 14613 1700
rect 14571 1651 14613 1660
rect 14572 1566 14612 1651
rect 14284 1147 14324 1156
rect 14668 1196 14708 2248
rect 14764 1205 14804 3163
rect 14859 2708 14901 2717
rect 14859 2668 14860 2708
rect 14900 2668 14901 2708
rect 14859 2659 14901 2668
rect 14860 2574 14900 2659
rect 14860 1952 14900 1961
rect 14860 1793 14900 1912
rect 14956 1952 14996 3247
rect 14859 1784 14901 1793
rect 14859 1744 14860 1784
rect 14900 1744 14901 1784
rect 14859 1735 14901 1744
rect 14956 1541 14996 1912
rect 14955 1532 14997 1541
rect 14955 1492 14956 1532
rect 14996 1492 14997 1532
rect 14955 1483 14997 1492
rect 15052 1364 15092 3424
rect 15435 3380 15477 3389
rect 15435 3340 15436 3380
rect 15476 3340 15477 3380
rect 15435 3331 15477 3340
rect 15436 3246 15476 3331
rect 15244 3212 15284 3221
rect 15147 1952 15189 1961
rect 15147 1912 15148 1952
rect 15188 1912 15189 1952
rect 15147 1903 15189 1912
rect 14956 1324 15092 1364
rect 14668 1147 14708 1156
rect 14763 1196 14805 1205
rect 14763 1156 14764 1196
rect 14804 1156 14805 1196
rect 14763 1147 14805 1156
rect 14476 944 14516 953
rect 14188 484 14420 524
rect 14283 356 14325 365
rect 14283 316 14284 356
rect 14324 316 14325 356
rect 14283 307 14325 316
rect 14284 80 14324 307
rect 14380 272 14420 484
rect 14476 449 14516 904
rect 14860 944 14900 953
rect 14667 860 14709 869
rect 14667 820 14668 860
rect 14708 820 14709 860
rect 14667 811 14709 820
rect 14475 440 14517 449
rect 14475 400 14476 440
rect 14516 400 14517 440
rect 14475 391 14517 400
rect 14380 232 14516 272
rect 14476 80 14516 232
rect 14668 80 14708 811
rect 14860 80 14900 904
rect 14956 701 14996 1324
rect 15148 1289 15188 1903
rect 15147 1280 15189 1289
rect 15147 1240 15148 1280
rect 15188 1240 15189 1280
rect 15147 1231 15189 1240
rect 15051 1196 15093 1205
rect 15051 1156 15052 1196
rect 15092 1156 15093 1196
rect 15051 1147 15093 1156
rect 15052 1062 15092 1147
rect 15147 944 15189 953
rect 15147 904 15148 944
rect 15188 904 15189 944
rect 15147 895 15189 904
rect 14955 692 14997 701
rect 14955 652 14956 692
rect 14996 652 14997 692
rect 14955 643 14997 652
rect 15148 524 15188 895
rect 15244 785 15284 3172
rect 15435 3128 15477 3137
rect 15435 3088 15436 3128
rect 15476 3088 15477 3128
rect 15435 3079 15477 3088
rect 15436 2801 15476 3079
rect 15435 2792 15477 2801
rect 15435 2752 15436 2792
rect 15476 2752 15477 2792
rect 15435 2743 15477 2752
rect 15339 2708 15381 2717
rect 15339 2668 15340 2708
rect 15380 2668 15381 2708
rect 15339 2659 15381 2668
rect 15340 2624 15380 2659
rect 15340 2573 15380 2584
rect 15339 1952 15381 1961
rect 15339 1912 15340 1952
rect 15380 1912 15381 1952
rect 15339 1903 15381 1912
rect 15436 1952 15476 2743
rect 15820 2540 15860 5515
rect 16012 5153 16052 5599
rect 16011 5144 16053 5153
rect 16011 5104 16012 5144
rect 16052 5104 16053 5144
rect 16011 5095 16053 5104
rect 16108 4397 16148 6868
rect 16300 6740 16340 13840
rect 16395 13460 16437 13469
rect 16395 13420 16396 13460
rect 16436 13420 16437 13460
rect 16395 13411 16437 13420
rect 16396 13326 16436 13411
rect 16395 12536 16437 12545
rect 16395 12496 16396 12536
rect 16436 12496 16437 12536
rect 16395 12487 16437 12496
rect 16396 10445 16436 12487
rect 16395 10436 16437 10445
rect 16395 10396 16396 10436
rect 16436 10396 16437 10436
rect 16395 10387 16437 10396
rect 16395 10016 16437 10025
rect 16395 9976 16396 10016
rect 16436 9976 16437 10016
rect 16395 9967 16437 9976
rect 16396 7085 16436 9967
rect 16492 7244 16532 14503
rect 16684 13880 16724 14755
rect 16780 14048 16820 15520
rect 16971 15560 17013 15569
rect 16971 15520 16972 15560
rect 17012 15520 17013 15560
rect 16971 15511 17013 15520
rect 17163 15560 17205 15569
rect 17163 15520 17164 15560
rect 17204 15520 17205 15560
rect 17163 15511 17205 15520
rect 17260 15485 17300 17611
rect 17355 17576 17397 17585
rect 17355 17536 17356 17576
rect 17396 17536 17397 17576
rect 17355 17527 17397 17536
rect 17356 16409 17396 17527
rect 17355 16400 17397 16409
rect 17355 16360 17356 16400
rect 17396 16360 17397 16400
rect 17355 16351 17397 16360
rect 17355 16232 17397 16241
rect 17355 16192 17356 16232
rect 17396 16192 17397 16232
rect 17355 16183 17397 16192
rect 17356 15989 17396 16183
rect 17355 15980 17397 15989
rect 17355 15940 17356 15980
rect 17396 15940 17397 15980
rect 17355 15931 17397 15940
rect 17355 15812 17397 15821
rect 17355 15772 17356 15812
rect 17396 15772 17397 15812
rect 17355 15763 17397 15772
rect 17356 15560 17396 15763
rect 16875 15476 16917 15485
rect 16875 15436 16876 15476
rect 16916 15436 16917 15476
rect 16875 15427 16917 15436
rect 17259 15476 17301 15485
rect 17259 15436 17260 15476
rect 17300 15436 17301 15476
rect 17259 15427 17301 15436
rect 16876 15342 16916 15427
rect 17356 14888 17396 15520
rect 16780 13999 16820 14008
rect 17164 14848 17396 14888
rect 16876 13964 16916 13973
rect 16876 13880 16916 13924
rect 16684 13840 16916 13880
rect 16683 13208 16725 13217
rect 16683 13168 16684 13208
rect 16724 13168 16725 13208
rect 16683 13159 16725 13168
rect 16684 13074 16724 13159
rect 16779 12620 16821 12629
rect 16779 12580 16780 12620
rect 16820 12580 16821 12620
rect 16779 12571 16821 12580
rect 17068 12620 17108 12629
rect 16587 11948 16629 11957
rect 16587 11908 16588 11948
rect 16628 11908 16629 11948
rect 16587 11899 16629 11908
rect 16588 10184 16628 11899
rect 16683 10436 16725 10445
rect 16683 10396 16684 10436
rect 16724 10396 16725 10436
rect 16683 10387 16725 10396
rect 16588 10025 16628 10144
rect 16587 10016 16629 10025
rect 16587 9976 16588 10016
rect 16628 9976 16629 10016
rect 16587 9967 16629 9976
rect 16684 9017 16724 10387
rect 16683 9008 16725 9017
rect 16683 8968 16684 9008
rect 16724 8968 16725 9008
rect 16683 8959 16725 8968
rect 16780 8840 16820 12571
rect 16876 12522 16916 12531
rect 16876 12041 16916 12482
rect 17068 12377 17108 12580
rect 17164 12545 17204 14848
rect 17356 14720 17396 14731
rect 17356 14645 17396 14680
rect 17355 14636 17397 14645
rect 17355 14596 17356 14636
rect 17396 14596 17397 14636
rect 17355 14587 17397 14596
rect 17452 14561 17492 17695
rect 17451 14552 17493 14561
rect 17451 14512 17452 14552
rect 17492 14512 17493 14552
rect 17451 14503 17493 14512
rect 17259 14048 17301 14057
rect 17259 14008 17260 14048
rect 17300 14008 17301 14048
rect 17259 13999 17301 14008
rect 17356 14048 17396 14057
rect 17260 13914 17300 13999
rect 17356 13469 17396 14008
rect 17355 13460 17397 13469
rect 17355 13420 17356 13460
rect 17396 13420 17397 13460
rect 17355 13411 17397 13420
rect 17355 13292 17397 13301
rect 17355 13252 17356 13292
rect 17396 13252 17397 13292
rect 17355 13243 17397 13252
rect 17163 12536 17205 12545
rect 17163 12496 17164 12536
rect 17204 12496 17205 12536
rect 17163 12487 17205 12496
rect 17067 12368 17109 12377
rect 17067 12328 17068 12368
rect 17108 12328 17109 12368
rect 17067 12319 17109 12328
rect 16875 12032 16917 12041
rect 16875 11992 16876 12032
rect 16916 11992 16917 12032
rect 16875 11983 16917 11992
rect 17259 12032 17301 12041
rect 17259 11992 17260 12032
rect 17300 11992 17301 12032
rect 17259 11983 17301 11992
rect 17260 11948 17300 11983
rect 17260 11897 17300 11908
rect 16971 11780 17013 11789
rect 17356 11780 17396 13243
rect 16971 11740 16972 11780
rect 17012 11740 17013 11780
rect 16971 11731 17013 11740
rect 17260 11740 17396 11780
rect 16972 11360 17012 11731
rect 17067 11696 17109 11705
rect 17067 11656 17068 11696
rect 17108 11656 17109 11696
rect 17067 11647 17109 11656
rect 17068 11562 17108 11647
rect 16972 11320 17108 11360
rect 17068 11024 17108 11320
rect 17068 10975 17108 10984
rect 16971 10856 17013 10865
rect 16971 10816 16972 10856
rect 17012 10816 17013 10856
rect 16971 10807 17013 10816
rect 16972 9008 17012 10807
rect 17116 10193 17156 10202
rect 17156 10153 17204 10184
rect 17116 10144 17204 10153
rect 17164 9689 17204 10144
rect 17260 10100 17300 11740
rect 17355 11612 17397 11621
rect 17355 11572 17356 11612
rect 17396 11572 17397 11612
rect 17355 11563 17397 11572
rect 17260 10051 17300 10060
rect 17163 9680 17205 9689
rect 17163 9640 17164 9680
rect 17204 9640 17205 9680
rect 17163 9631 17205 9640
rect 17260 9512 17300 9521
rect 17356 9512 17396 11563
rect 17452 10352 17492 10361
rect 17452 10193 17492 10312
rect 17451 10184 17493 10193
rect 17451 10144 17452 10184
rect 17492 10144 17493 10184
rect 17451 10135 17493 10144
rect 17451 9680 17493 9689
rect 17451 9640 17452 9680
rect 17492 9640 17493 9680
rect 17451 9631 17493 9640
rect 17452 9546 17492 9631
rect 17300 9472 17396 9512
rect 17260 9463 17300 9472
rect 16972 8968 17204 9008
rect 17068 8840 17108 8849
rect 16588 8800 16820 8840
rect 16876 8800 17068 8840
rect 16588 8000 16628 8800
rect 16876 8756 16916 8800
rect 17068 8791 17108 8800
rect 16684 8716 16916 8756
rect 16684 8686 16724 8716
rect 17164 8714 17204 8968
rect 17071 8674 17204 8714
rect 17071 8672 17111 8674
rect 16684 8637 16724 8646
rect 16972 8632 17111 8672
rect 17259 8672 17301 8681
rect 17259 8632 17260 8672
rect 17300 8632 17301 8672
rect 16779 8588 16821 8597
rect 16779 8548 16780 8588
rect 16820 8548 16821 8588
rect 16779 8539 16821 8548
rect 16684 8000 16724 8009
rect 16588 7960 16684 8000
rect 16492 7195 16532 7204
rect 16587 7244 16629 7253
rect 16587 7204 16588 7244
rect 16628 7204 16629 7244
rect 16587 7195 16629 7204
rect 16588 7110 16628 7195
rect 16684 7169 16724 7960
rect 16683 7160 16725 7169
rect 16683 7120 16684 7160
rect 16724 7120 16725 7160
rect 16683 7111 16725 7120
rect 16395 7076 16437 7085
rect 16395 7036 16396 7076
rect 16436 7036 16437 7076
rect 16395 7027 16437 7036
rect 16395 6824 16437 6833
rect 16395 6784 16396 6824
rect 16436 6784 16437 6824
rect 16395 6775 16437 6784
rect 16204 6700 16340 6740
rect 16107 4388 16149 4397
rect 16107 4348 16108 4388
rect 16148 4348 16149 4388
rect 16107 4339 16149 4348
rect 16108 4229 16148 4339
rect 16107 4220 16149 4229
rect 16107 4180 16108 4220
rect 16148 4180 16149 4220
rect 16107 4171 16149 4180
rect 16011 4136 16053 4145
rect 16011 4096 16012 4136
rect 16052 4096 16053 4136
rect 16011 4087 16053 4096
rect 16012 4002 16052 4087
rect 15820 2500 15956 2540
rect 15436 1903 15476 1912
rect 15916 1952 15956 2500
rect 15916 1903 15956 1912
rect 15340 1818 15380 1903
rect 15339 1700 15381 1709
rect 15339 1660 15340 1700
rect 15380 1660 15381 1700
rect 15339 1651 15381 1660
rect 15243 776 15285 785
rect 15243 736 15244 776
rect 15284 736 15285 776
rect 15243 727 15285 736
rect 15340 692 15380 1651
rect 16011 1448 16053 1457
rect 16011 1408 16012 1448
rect 16052 1408 16053 1448
rect 16011 1399 16053 1408
rect 15435 1280 15477 1289
rect 15435 1240 15436 1280
rect 15476 1240 15477 1280
rect 15435 1231 15477 1240
rect 15436 1112 15476 1231
rect 15436 1063 15476 1072
rect 15627 692 15669 701
rect 15340 652 15476 692
rect 15148 484 15284 524
rect 15051 356 15093 365
rect 15051 316 15052 356
rect 15092 316 15093 356
rect 15051 307 15093 316
rect 15052 80 15092 307
rect 15244 80 15284 484
rect 15436 80 15476 652
rect 15627 652 15628 692
rect 15668 652 15669 692
rect 15627 643 15669 652
rect 15628 80 15668 643
rect 15819 608 15861 617
rect 15819 568 15820 608
rect 15860 568 15861 608
rect 15819 559 15861 568
rect 15820 80 15860 559
rect 16012 80 16052 1399
rect 16204 80 16244 6700
rect 16299 6236 16341 6245
rect 16299 6196 16300 6236
rect 16340 6196 16341 6236
rect 16299 6187 16341 6196
rect 16300 5648 16340 6187
rect 16300 5599 16340 5608
rect 16396 2036 16436 6775
rect 16491 5396 16533 5405
rect 16491 5356 16492 5396
rect 16532 5356 16533 5396
rect 16491 5347 16533 5356
rect 16492 4976 16532 5347
rect 16492 4927 16532 4936
rect 16684 4724 16724 4733
rect 16684 4229 16724 4684
rect 16491 4220 16533 4229
rect 16491 4180 16492 4220
rect 16532 4180 16533 4220
rect 16491 4171 16533 4180
rect 16683 4220 16725 4229
rect 16683 4180 16684 4220
rect 16724 4180 16725 4220
rect 16683 4171 16725 4180
rect 16492 4150 16532 4171
rect 16780 4145 16820 8539
rect 16875 8504 16917 8513
rect 16875 8464 16876 8504
rect 16916 8464 16917 8504
rect 16875 8455 16917 8464
rect 16876 8370 16916 8455
rect 16875 8168 16917 8177
rect 16875 8128 16876 8168
rect 16916 8128 16917 8168
rect 16875 8119 16917 8128
rect 16876 6833 16916 8119
rect 16875 6824 16917 6833
rect 16875 6784 16876 6824
rect 16916 6784 16917 6824
rect 16875 6775 16917 6784
rect 16972 5816 17012 8632
rect 17259 8623 17301 8632
rect 17260 7925 17300 8623
rect 17356 8177 17396 9472
rect 17451 9092 17493 9101
rect 17451 9052 17452 9092
rect 17492 9052 17493 9092
rect 17451 9043 17493 9052
rect 17355 8168 17397 8177
rect 17355 8128 17356 8168
rect 17396 8128 17397 8168
rect 17355 8119 17397 8128
rect 17452 8000 17492 9043
rect 17548 8849 17588 17872
rect 17644 15812 17684 22072
rect 17835 21608 17877 21617
rect 17835 21568 17836 21608
rect 17876 21568 17877 21608
rect 17835 21559 17877 21568
rect 17739 21104 17781 21113
rect 17739 21064 17740 21104
rect 17780 21064 17781 21104
rect 17739 21055 17781 21064
rect 17740 20096 17780 21055
rect 17836 20852 17876 21559
rect 17836 20803 17876 20812
rect 17932 20852 17972 22231
rect 17932 20803 17972 20812
rect 17740 19265 17780 20056
rect 17931 20012 17973 20021
rect 17931 19972 17932 20012
rect 17972 19972 17973 20012
rect 17931 19963 17973 19972
rect 17932 19928 17972 19963
rect 17932 19877 17972 19888
rect 17739 19256 17781 19265
rect 17739 19216 17740 19256
rect 17780 19216 17781 19256
rect 17739 19207 17781 19216
rect 17836 19256 17876 19265
rect 17740 18341 17780 19207
rect 17836 19097 17876 19216
rect 17835 19088 17877 19097
rect 17835 19048 17836 19088
rect 17876 19048 17877 19088
rect 17835 19039 17877 19048
rect 17739 18332 17781 18341
rect 17739 18292 17740 18332
rect 17780 18292 17781 18332
rect 17739 18283 17781 18292
rect 17931 18164 17973 18173
rect 17931 18124 17932 18164
rect 17972 18124 17973 18164
rect 17931 18115 17973 18124
rect 17932 17744 17972 18115
rect 17932 17695 17972 17704
rect 18028 16988 18068 22483
rect 18124 22112 18164 22996
rect 18219 22616 18261 22625
rect 18219 22576 18220 22616
rect 18260 22576 18261 22616
rect 18219 22567 18261 22576
rect 18220 22289 18260 22567
rect 18219 22280 18261 22289
rect 18219 22240 18220 22280
rect 18260 22240 18261 22280
rect 18219 22231 18261 22240
rect 18124 22072 18260 22112
rect 18123 21860 18165 21869
rect 18123 21820 18124 21860
rect 18164 21820 18165 21860
rect 18123 21811 18165 21820
rect 18124 21608 18164 21811
rect 18124 20777 18164 21568
rect 18123 20768 18165 20777
rect 18123 20728 18124 20768
rect 18164 20728 18165 20768
rect 18123 20719 18165 20728
rect 18123 20096 18165 20105
rect 18123 20056 18124 20096
rect 18164 20056 18165 20096
rect 18123 20047 18165 20056
rect 18124 19962 18164 20047
rect 18220 19853 18260 22072
rect 18316 21776 18356 23752
rect 18507 23792 18549 23801
rect 18507 23752 18508 23792
rect 18548 23752 18549 23792
rect 18507 23743 18549 23752
rect 18604 23792 18644 24415
rect 18808 24212 19176 24221
rect 18848 24172 18890 24212
rect 18930 24172 18972 24212
rect 19012 24172 19054 24212
rect 19094 24172 19136 24212
rect 18808 24163 19176 24172
rect 19660 24137 19700 24508
rect 19756 24212 19796 25087
rect 19852 24641 19892 25264
rect 19851 24632 19893 24641
rect 19851 24592 19852 24632
rect 19892 24592 19893 24632
rect 19851 24583 19893 24592
rect 19851 24464 19893 24473
rect 19851 24424 19852 24464
rect 19892 24424 19893 24464
rect 19851 24415 19893 24424
rect 19852 24330 19892 24415
rect 19756 24172 19892 24212
rect 19659 24128 19701 24137
rect 19659 24088 19660 24128
rect 19700 24088 19701 24128
rect 19659 24079 19701 24088
rect 18987 24044 19029 24053
rect 18987 24004 18988 24044
rect 19028 24004 19029 24044
rect 18987 23995 19029 24004
rect 18411 23708 18453 23717
rect 18411 23668 18412 23708
rect 18452 23668 18453 23708
rect 18411 23659 18453 23668
rect 18412 23574 18452 23659
rect 18508 23658 18548 23743
rect 18604 23549 18644 23752
rect 18891 23792 18933 23801
rect 18891 23752 18892 23792
rect 18932 23752 18933 23792
rect 18891 23743 18933 23752
rect 18988 23792 19028 23995
rect 19276 23969 19316 24054
rect 19275 23960 19317 23969
rect 19275 23920 19276 23960
rect 19316 23920 19317 23960
rect 19275 23911 19317 23920
rect 19659 23960 19701 23969
rect 19659 23920 19660 23960
rect 19700 23920 19701 23960
rect 19659 23911 19701 23920
rect 19564 23801 19604 23886
rect 18795 23624 18837 23633
rect 18795 23584 18796 23624
rect 18836 23584 18837 23624
rect 18795 23575 18837 23584
rect 18603 23540 18645 23549
rect 18603 23500 18604 23540
rect 18644 23500 18645 23540
rect 18603 23491 18645 23500
rect 18412 23288 18452 23297
rect 18507 23288 18549 23297
rect 18452 23248 18508 23288
rect 18548 23248 18549 23288
rect 18412 23239 18452 23248
rect 18507 23239 18549 23248
rect 18699 23204 18741 23213
rect 18699 23164 18700 23204
rect 18740 23164 18741 23204
rect 18699 23155 18741 23164
rect 18604 23099 18648 23120
rect 18644 23059 18648 23099
rect 18604 23050 18648 23059
rect 18608 22961 18648 23050
rect 18603 22952 18648 22961
rect 18603 22912 18604 22952
rect 18644 22912 18648 22952
rect 18603 22903 18645 22912
rect 18411 22784 18453 22793
rect 18411 22744 18412 22784
rect 18452 22744 18453 22784
rect 18411 22735 18453 22744
rect 18316 21727 18356 21736
rect 18412 21701 18452 22735
rect 18700 22294 18740 23155
rect 18796 22961 18836 23575
rect 18795 22952 18837 22961
rect 18795 22912 18796 22952
rect 18836 22912 18837 22952
rect 18795 22903 18837 22912
rect 18892 22877 18932 23743
rect 18988 23036 19028 23752
rect 19084 23792 19124 23801
rect 19468 23792 19508 23801
rect 19124 23752 19468 23792
rect 19084 23213 19124 23752
rect 19468 23743 19508 23752
rect 19563 23792 19605 23801
rect 19563 23752 19564 23792
rect 19604 23752 19605 23792
rect 19563 23743 19605 23752
rect 19660 23792 19700 23911
rect 19660 23743 19700 23752
rect 19756 23624 19796 23633
rect 19564 23584 19756 23624
rect 19083 23204 19125 23213
rect 19083 23164 19084 23204
rect 19124 23164 19125 23204
rect 19083 23155 19125 23164
rect 18988 22996 19412 23036
rect 18891 22868 18933 22877
rect 18891 22828 18892 22868
rect 18932 22828 18933 22868
rect 18891 22819 18933 22828
rect 18808 22700 19176 22709
rect 18848 22660 18890 22700
rect 18930 22660 18972 22700
rect 19012 22660 19054 22700
rect 19094 22660 19136 22700
rect 18808 22651 19176 22660
rect 18891 22448 18933 22457
rect 18891 22408 18892 22448
rect 18932 22408 18933 22448
rect 18891 22399 18933 22408
rect 18507 22280 18549 22289
rect 18507 22240 18508 22280
rect 18548 22240 18549 22280
rect 18700 22245 18740 22254
rect 18507 22231 18549 22240
rect 18411 21692 18453 21701
rect 18411 21652 18412 21692
rect 18452 21652 18453 21692
rect 18411 21643 18453 21652
rect 18412 21608 18452 21643
rect 18508 21617 18548 22231
rect 18892 22196 18932 22399
rect 19180 22289 19220 22374
rect 19179 22280 19221 22289
rect 19179 22240 19180 22280
rect 19220 22240 19221 22280
rect 19179 22231 19221 22240
rect 18892 22147 18932 22156
rect 19372 22112 19412 22996
rect 19467 22448 19509 22457
rect 19467 22408 19468 22448
rect 19508 22408 19509 22448
rect 19467 22399 19509 22408
rect 19468 22280 19508 22399
rect 19468 22231 19508 22240
rect 19564 22280 19604 23584
rect 19756 23575 19796 23584
rect 19852 23456 19892 24172
rect 19948 23876 19988 26356
rect 20044 26060 20084 26069
rect 20044 25565 20084 26020
rect 20235 25976 20277 25985
rect 20235 25936 20236 25976
rect 20276 25936 20277 25976
rect 20235 25927 20277 25936
rect 20236 25842 20276 25927
rect 20043 25556 20085 25565
rect 20043 25516 20044 25556
rect 20084 25516 20085 25556
rect 20043 25507 20085 25516
rect 20043 25304 20085 25313
rect 20043 25264 20044 25304
rect 20084 25264 20085 25304
rect 20043 25255 20085 25264
rect 20044 25136 20084 25255
rect 20044 25087 20084 25096
rect 20048 24968 20416 24977
rect 20088 24928 20130 24968
rect 20170 24928 20212 24968
rect 20252 24928 20294 24968
rect 20334 24928 20376 24968
rect 20048 24919 20416 24928
rect 20235 24800 20277 24809
rect 20235 24760 20236 24800
rect 20276 24760 20277 24800
rect 20235 24751 20277 24760
rect 20236 24666 20276 24751
rect 19948 23827 19988 23836
rect 20044 24548 20084 24557
rect 20044 23624 20084 24508
rect 20140 23633 20180 23718
rect 19756 23416 19892 23456
rect 19948 23584 20084 23624
rect 20139 23624 20181 23633
rect 20139 23584 20140 23624
rect 20180 23584 20181 23624
rect 19659 22448 19701 22457
rect 19659 22408 19660 22448
rect 19700 22408 19701 22448
rect 19659 22399 19701 22408
rect 19564 22231 19604 22240
rect 19372 22072 19508 22112
rect 18699 21776 18741 21785
rect 18699 21736 18700 21776
rect 18740 21736 18741 21776
rect 18699 21727 18741 21736
rect 18412 21558 18452 21568
rect 18507 21608 18549 21617
rect 18507 21568 18508 21608
rect 18548 21568 18549 21608
rect 18507 21559 18549 21568
rect 18700 21608 18740 21727
rect 18700 21559 18740 21568
rect 18808 21188 19176 21197
rect 18848 21148 18890 21188
rect 18930 21148 18972 21188
rect 19012 21148 19054 21188
rect 19094 21148 19136 21188
rect 18808 21139 19176 21148
rect 18940 20777 18980 20786
rect 18411 20768 18453 20777
rect 18411 20728 18412 20768
rect 18452 20728 18453 20768
rect 18411 20719 18453 20728
rect 18892 20737 18940 20768
rect 19372 20768 19412 20777
rect 18980 20737 19372 20768
rect 18892 20728 19372 20737
rect 18412 20634 18452 20719
rect 18892 20105 18932 20728
rect 19084 20600 19124 20609
rect 18411 20096 18453 20105
rect 18411 20056 18412 20096
rect 18452 20056 18453 20096
rect 18411 20047 18453 20056
rect 18700 20096 18740 20105
rect 18412 19962 18452 20047
rect 18219 19844 18261 19853
rect 18219 19804 18220 19844
rect 18260 19804 18261 19844
rect 18219 19795 18261 19804
rect 18412 19844 18452 19853
rect 18452 19804 18548 19844
rect 18412 19795 18452 19804
rect 18123 18584 18165 18593
rect 18123 18544 18124 18584
rect 18164 18544 18165 18584
rect 18123 18535 18165 18544
rect 17836 16948 18068 16988
rect 17644 15772 17780 15812
rect 17643 14216 17685 14225
rect 17643 14176 17644 14216
rect 17684 14176 17685 14216
rect 17643 14167 17685 14176
rect 17644 14082 17684 14167
rect 17643 13460 17685 13469
rect 17643 13420 17644 13460
rect 17684 13420 17685 13460
rect 17643 13411 17685 13420
rect 17644 10268 17684 13411
rect 17644 10219 17684 10228
rect 17643 9512 17685 9521
rect 17643 9472 17644 9512
rect 17684 9472 17685 9512
rect 17643 9463 17685 9472
rect 17644 9378 17684 9463
rect 17740 8849 17780 15772
rect 17836 15737 17876 16948
rect 18028 16820 18068 16829
rect 18028 15812 18068 16780
rect 18124 16241 18164 18535
rect 18220 17753 18260 19795
rect 18412 18584 18452 18595
rect 18508 18584 18548 19804
rect 18700 18761 18740 20056
rect 18891 20096 18933 20105
rect 18891 20056 18892 20096
rect 18932 20056 18933 20096
rect 18891 20047 18933 20056
rect 19084 19844 19124 20560
rect 19179 20600 19221 20609
rect 19179 20560 19180 20600
rect 19220 20560 19221 20600
rect 19179 20551 19221 20560
rect 19180 20105 19220 20551
rect 19179 20096 19221 20105
rect 19179 20056 19180 20096
rect 19220 20056 19221 20096
rect 19179 20047 19221 20056
rect 19084 19804 19316 19844
rect 19276 19685 19316 19804
rect 18808 19676 19176 19685
rect 18848 19636 18890 19676
rect 18930 19636 18972 19676
rect 19012 19636 19054 19676
rect 19094 19636 19136 19676
rect 18808 19627 19176 19636
rect 19275 19676 19317 19685
rect 19275 19636 19276 19676
rect 19316 19636 19317 19676
rect 19275 19627 19317 19636
rect 19276 19508 19316 19517
rect 19372 19508 19412 20728
rect 19316 19468 19412 19508
rect 19468 20768 19508 22072
rect 19276 19459 19316 19468
rect 19084 19265 19124 19350
rect 19083 19256 19125 19265
rect 19083 19216 19084 19256
rect 19124 19216 19125 19256
rect 19083 19207 19125 19216
rect 19276 19088 19316 19097
rect 18988 19048 19276 19088
rect 18699 18752 18741 18761
rect 18699 18712 18700 18752
rect 18740 18712 18741 18752
rect 18699 18703 18741 18712
rect 18891 18752 18933 18761
rect 18891 18712 18892 18752
rect 18932 18712 18933 18752
rect 18891 18703 18933 18712
rect 18892 18618 18932 18703
rect 18796 18584 18836 18593
rect 18508 18544 18796 18584
rect 18412 18509 18452 18544
rect 18796 18535 18836 18544
rect 18988 18584 19028 19048
rect 19276 19039 19316 19048
rect 19083 18920 19125 18929
rect 19083 18880 19084 18920
rect 19124 18880 19125 18920
rect 19083 18871 19125 18880
rect 18988 18535 19028 18544
rect 19084 18584 19124 18871
rect 19124 18544 19316 18584
rect 19084 18535 19124 18544
rect 18411 18500 18453 18509
rect 18411 18460 18412 18500
rect 18452 18460 18453 18500
rect 18411 18451 18453 18460
rect 18604 18332 18644 18341
rect 18508 18292 18604 18332
rect 18508 17828 18548 18292
rect 18604 18283 18644 18292
rect 18808 18164 19176 18173
rect 18848 18124 18890 18164
rect 18930 18124 18972 18164
rect 19012 18124 19054 18164
rect 19094 18124 19136 18164
rect 18808 18115 19176 18124
rect 18460 17788 18548 17828
rect 18460 17786 18500 17788
rect 18219 17744 18261 17753
rect 18219 17704 18220 17744
rect 18260 17704 18261 17744
rect 18460 17737 18500 17746
rect 18987 17744 19029 17753
rect 18219 17695 18261 17704
rect 18987 17704 18988 17744
rect 19028 17704 19029 17744
rect 18987 17695 19029 17704
rect 18988 17610 19028 17695
rect 19083 17660 19125 17669
rect 19083 17620 19084 17660
rect 19124 17620 19125 17660
rect 19083 17611 19125 17620
rect 18604 17576 18644 17585
rect 18796 17576 18836 17585
rect 18220 17536 18604 17576
rect 18220 16988 18260 17536
rect 18604 17527 18644 17536
rect 18700 17536 18796 17576
rect 18700 17324 18740 17536
rect 18796 17527 18836 17536
rect 18604 17284 18740 17324
rect 18220 16939 18260 16948
rect 18412 17156 18452 17165
rect 18219 16400 18261 16409
rect 18219 16360 18220 16400
rect 18260 16360 18261 16400
rect 18219 16351 18261 16360
rect 18123 16232 18165 16241
rect 18123 16192 18124 16232
rect 18164 16192 18165 16232
rect 18123 16183 18165 16192
rect 17932 15772 18068 15812
rect 17835 15728 17877 15737
rect 17835 15688 17836 15728
rect 17876 15688 17877 15728
rect 17835 15679 17877 15688
rect 17835 15560 17877 15569
rect 17835 15515 17836 15560
rect 17876 15515 17877 15560
rect 17835 15511 17877 15515
rect 17836 15425 17876 15511
rect 17932 15233 17972 15772
rect 18123 15728 18165 15737
rect 18123 15688 18124 15728
rect 18164 15688 18165 15728
rect 18123 15679 18165 15688
rect 18028 15644 18068 15653
rect 17931 15224 17973 15233
rect 17931 15184 17932 15224
rect 17972 15184 17973 15224
rect 17931 15175 17973 15184
rect 17836 14048 17876 14059
rect 17836 13973 17876 14008
rect 17835 13964 17877 13973
rect 17835 13924 17836 13964
rect 17876 13924 17877 13964
rect 17835 13915 17877 13924
rect 18028 13469 18068 15604
rect 18124 14981 18164 15679
rect 18123 14972 18165 14981
rect 18123 14932 18124 14972
rect 18164 14932 18165 14972
rect 18123 14923 18165 14932
rect 18027 13460 18069 13469
rect 18027 13420 18028 13460
rect 18068 13420 18069 13460
rect 18027 13411 18069 13420
rect 18124 13292 18164 14923
rect 18220 13301 18260 16351
rect 18315 15140 18357 15149
rect 18315 15100 18316 15140
rect 18356 15100 18357 15140
rect 18315 15091 18357 15100
rect 18316 14804 18356 15091
rect 18412 14888 18452 17116
rect 18604 17067 18644 17284
rect 18604 17018 18644 17027
rect 19084 17072 19124 17611
rect 19084 17023 19124 17032
rect 18699 16988 18741 16997
rect 18699 16948 18700 16988
rect 18740 16948 18741 16988
rect 18699 16939 18741 16948
rect 18507 16400 18549 16409
rect 18507 16360 18508 16400
rect 18548 16360 18549 16400
rect 18507 16351 18549 16360
rect 18508 15560 18548 16351
rect 18603 16232 18645 16241
rect 18603 16192 18604 16232
rect 18644 16192 18645 16232
rect 18603 16183 18645 16192
rect 18604 16098 18644 16183
rect 18508 15511 18548 15520
rect 18412 14848 18644 14888
rect 18316 14764 18452 14804
rect 18412 14720 18452 14764
rect 18316 14700 18356 14709
rect 18452 14680 18548 14720
rect 18412 14671 18452 14680
rect 18316 14225 18356 14660
rect 18315 14216 18357 14225
rect 18315 14176 18316 14216
rect 18356 14176 18357 14216
rect 18315 14167 18357 14176
rect 18028 13252 18164 13292
rect 18219 13292 18261 13301
rect 18219 13252 18220 13292
rect 18260 13252 18261 13292
rect 17932 13208 17972 13217
rect 17932 11537 17972 13168
rect 17931 11528 17973 11537
rect 17931 11488 17932 11528
rect 17972 11488 17973 11528
rect 17931 11479 17973 11488
rect 18028 10865 18068 13252
rect 18219 13243 18261 13252
rect 18412 13208 18452 13217
rect 18124 13124 18164 13133
rect 18412 13124 18452 13168
rect 18164 13084 18452 13124
rect 18508 13208 18548 14680
rect 18124 13075 18164 13084
rect 18508 12620 18548 13168
rect 18124 12580 18548 12620
rect 18027 10856 18069 10865
rect 18027 10816 18028 10856
rect 18068 10816 18069 10856
rect 18027 10807 18069 10816
rect 18124 10613 18164 12580
rect 18220 11824 18548 11864
rect 18220 11201 18260 11824
rect 18412 11696 18452 11705
rect 18315 11528 18357 11537
rect 18315 11488 18316 11528
rect 18356 11488 18357 11528
rect 18315 11479 18357 11488
rect 18219 11192 18261 11201
rect 18219 11152 18220 11192
rect 18260 11152 18261 11192
rect 18219 11143 18261 11152
rect 17931 10604 17973 10613
rect 17931 10564 17932 10604
rect 17972 10564 17973 10604
rect 17931 10555 17973 10564
rect 18123 10604 18165 10613
rect 18123 10564 18124 10604
rect 18164 10564 18165 10604
rect 18123 10555 18165 10564
rect 17835 9848 17877 9857
rect 17835 9808 17836 9848
rect 17876 9808 17877 9848
rect 17835 9799 17877 9808
rect 17547 8840 17589 8849
rect 17547 8800 17548 8840
rect 17588 8800 17589 8840
rect 17547 8791 17589 8800
rect 17739 8840 17781 8849
rect 17739 8800 17740 8840
rect 17780 8800 17781 8840
rect 17739 8791 17781 8800
rect 17643 8168 17685 8177
rect 17643 8128 17644 8168
rect 17684 8128 17685 8168
rect 17643 8119 17685 8128
rect 17356 7960 17492 8000
rect 17259 7916 17301 7925
rect 17259 7876 17260 7916
rect 17300 7876 17301 7916
rect 17259 7867 17301 7876
rect 17068 7160 17108 7171
rect 17068 7085 17108 7120
rect 17067 7076 17109 7085
rect 17067 7036 17068 7076
rect 17108 7036 17109 7076
rect 17067 7027 17109 7036
rect 17356 6824 17396 7960
rect 17548 7165 17588 7174
rect 17548 6992 17588 7125
rect 17164 6784 17396 6824
rect 17537 6952 17588 6992
rect 17067 6488 17109 6497
rect 17067 6448 17068 6488
rect 17108 6448 17109 6488
rect 17067 6439 17109 6448
rect 17068 6354 17108 6439
rect 17164 6152 17204 6784
rect 17537 6740 17577 6952
rect 17260 6700 17577 6740
rect 17260 6656 17300 6700
rect 17260 6607 17300 6616
rect 16876 5776 17012 5816
rect 17068 6112 17204 6152
rect 17355 6152 17397 6161
rect 17355 6112 17356 6152
rect 17396 6112 17397 6152
rect 16876 4976 16916 5776
rect 16971 5648 17013 5657
rect 16971 5608 16972 5648
rect 17012 5608 17013 5648
rect 16971 5599 17013 5608
rect 16492 4085 16532 4110
rect 16779 4136 16821 4145
rect 16779 4096 16780 4136
rect 16820 4096 16821 4136
rect 16779 4087 16821 4096
rect 16684 3968 16724 3977
rect 16684 3641 16724 3928
rect 16683 3632 16725 3641
rect 16683 3592 16684 3632
rect 16724 3592 16725 3632
rect 16683 3583 16725 3592
rect 16684 3464 16724 3473
rect 16684 2960 16724 3424
rect 16779 3464 16821 3473
rect 16779 3424 16780 3464
rect 16820 3424 16821 3464
rect 16779 3415 16821 3424
rect 16780 3330 16820 3415
rect 16684 2920 16820 2960
rect 16780 2876 16820 2920
rect 16780 2827 16820 2836
rect 16588 2645 16628 2719
rect 16587 2584 16588 2633
rect 16628 2584 16629 2633
rect 16876 2624 16916 4936
rect 16972 3473 17012 5599
rect 16971 3464 17013 3473
rect 16971 3424 16972 3464
rect 17012 3424 17013 3464
rect 16971 3415 17013 3424
rect 16972 2624 17012 2633
rect 16876 2584 16972 2624
rect 16587 2575 16629 2584
rect 16972 2575 17012 2584
rect 16683 2540 16725 2549
rect 16683 2500 16684 2540
rect 16724 2500 16725 2540
rect 16683 2491 16725 2500
rect 16587 2036 16629 2045
rect 16396 1996 16532 2036
rect 16396 1938 16436 1947
rect 16299 1868 16341 1877
rect 16396 1868 16436 1898
rect 16299 1828 16300 1868
rect 16340 1828 16436 1868
rect 16299 1819 16341 1828
rect 16492 1784 16532 1996
rect 16587 1996 16588 2036
rect 16628 1996 16629 2036
rect 16587 1987 16629 1996
rect 16588 1902 16628 1987
rect 16396 1744 16532 1784
rect 16587 1784 16629 1793
rect 16587 1744 16588 1784
rect 16628 1744 16629 1784
rect 16396 80 16436 1744
rect 16587 1735 16629 1744
rect 16588 80 16628 1735
rect 16684 1121 16724 2491
rect 16779 1952 16821 1961
rect 16779 1912 16780 1952
rect 16820 1912 16821 1952
rect 16779 1903 16821 1912
rect 16780 1818 16820 1903
rect 16875 1868 16917 1877
rect 16875 1828 16876 1868
rect 16916 1828 16917 1868
rect 16875 1819 16917 1828
rect 16779 1700 16821 1709
rect 16779 1660 16780 1700
rect 16820 1660 16821 1700
rect 16779 1651 16821 1660
rect 16683 1112 16725 1121
rect 16683 1072 16684 1112
rect 16724 1072 16725 1112
rect 16683 1063 16725 1072
rect 16684 978 16724 1063
rect 16780 80 16820 1651
rect 16876 1364 16916 1819
rect 16876 1315 16916 1324
rect 16971 1112 17013 1121
rect 16971 1072 16972 1112
rect 17012 1072 17013 1112
rect 16971 1063 17013 1072
rect 16972 80 17012 1063
rect 17068 776 17108 6112
rect 17355 6103 17397 6112
rect 17163 4388 17205 4397
rect 17163 4348 17164 4388
rect 17204 4348 17205 4388
rect 17163 4339 17205 4348
rect 17356 4388 17396 6103
rect 17548 5741 17588 5772
rect 17547 5732 17589 5741
rect 17547 5692 17548 5732
rect 17588 5692 17589 5732
rect 17547 5683 17589 5692
rect 17548 5648 17588 5683
rect 17548 5405 17588 5608
rect 17644 5573 17684 8119
rect 17836 7757 17876 9799
rect 17932 8177 17972 10555
rect 18220 10352 18260 11143
rect 18124 10312 18260 10352
rect 18316 11024 18356 11479
rect 18412 11192 18452 11656
rect 18508 11696 18548 11824
rect 18508 11647 18548 11656
rect 18508 11192 18548 11201
rect 18412 11152 18508 11192
rect 18508 11143 18548 11152
rect 18027 10100 18069 10109
rect 18027 10060 18028 10100
rect 18068 10060 18069 10100
rect 18027 10051 18069 10060
rect 18028 9966 18068 10051
rect 18027 9428 18069 9437
rect 18027 9388 18028 9428
rect 18068 9388 18069 9428
rect 18027 9379 18069 9388
rect 17931 8168 17973 8177
rect 17931 8128 17932 8168
rect 17972 8128 17973 8168
rect 17931 8119 17973 8128
rect 17835 7748 17877 7757
rect 17835 7708 17836 7748
rect 17876 7708 17877 7748
rect 17835 7699 17877 7708
rect 17931 7496 17973 7505
rect 17931 7456 17932 7496
rect 17972 7456 17973 7496
rect 17931 7447 17973 7456
rect 17932 7412 17972 7447
rect 17932 7361 17972 7372
rect 18028 7253 18068 9379
rect 18124 8177 18164 10312
rect 18220 10193 18260 10198
rect 18219 10189 18261 10193
rect 18219 10144 18220 10189
rect 18260 10144 18261 10189
rect 18219 10135 18261 10144
rect 18220 10054 18260 10135
rect 18316 8924 18356 10984
rect 18411 10856 18453 10865
rect 18411 10816 18412 10856
rect 18452 10816 18453 10856
rect 18411 10807 18453 10816
rect 18220 8884 18356 8924
rect 18220 8513 18260 8884
rect 18412 8840 18452 10807
rect 18507 10436 18549 10445
rect 18507 10396 18508 10436
rect 18548 10396 18549 10436
rect 18507 10387 18549 10396
rect 18508 9017 18548 10387
rect 18507 9008 18549 9017
rect 18507 8968 18508 9008
rect 18548 8968 18549 9008
rect 18507 8959 18549 8968
rect 18316 8800 18452 8840
rect 18219 8504 18261 8513
rect 18219 8464 18220 8504
rect 18260 8464 18261 8504
rect 18219 8455 18261 8464
rect 18316 8252 18356 8800
rect 18507 8756 18549 8765
rect 18507 8716 18508 8756
rect 18548 8716 18549 8756
rect 18507 8707 18549 8716
rect 18508 8672 18548 8707
rect 18508 8621 18548 8632
rect 18507 8504 18549 8513
rect 18507 8464 18508 8504
rect 18548 8464 18549 8504
rect 18507 8455 18549 8464
rect 18316 8212 18452 8252
rect 18123 8168 18165 8177
rect 18123 8128 18124 8168
rect 18164 8128 18165 8168
rect 18123 8119 18165 8128
rect 18316 8009 18356 8094
rect 18315 8000 18357 8009
rect 18220 7986 18260 7990
rect 18124 7981 18260 7986
rect 18124 7946 18220 7981
rect 18124 7505 18164 7946
rect 18315 7960 18316 8000
rect 18356 7960 18357 8000
rect 18315 7951 18357 7960
rect 18220 7932 18260 7941
rect 18315 7832 18357 7841
rect 18315 7792 18316 7832
rect 18356 7792 18357 7832
rect 18315 7783 18357 7792
rect 18123 7496 18165 7505
rect 18123 7456 18124 7496
rect 18164 7456 18165 7496
rect 18123 7447 18165 7456
rect 18123 7328 18165 7337
rect 18123 7288 18124 7328
rect 18164 7288 18165 7328
rect 18123 7279 18165 7288
rect 18027 7244 18069 7253
rect 18027 7204 18028 7244
rect 18068 7204 18069 7244
rect 18027 7195 18069 7204
rect 17740 6992 17780 7001
rect 18028 6992 18068 7195
rect 18124 7160 18164 7279
rect 18124 7111 18164 7120
rect 18028 6952 18164 6992
rect 17740 6749 17780 6952
rect 17739 6740 17781 6749
rect 17739 6700 17740 6740
rect 17780 6700 17781 6740
rect 17739 6691 17781 6700
rect 18028 6488 18068 6497
rect 17740 6448 18028 6488
rect 17740 5900 17780 6448
rect 18028 6439 18068 6448
rect 18124 6488 18164 6952
rect 18124 6439 18164 6448
rect 17740 5851 17780 5860
rect 17931 5732 17973 5741
rect 17931 5692 17932 5732
rect 17972 5692 17973 5732
rect 17931 5683 17973 5692
rect 17643 5564 17685 5573
rect 17643 5524 17644 5564
rect 17684 5524 17685 5564
rect 17643 5515 17685 5524
rect 17547 5396 17589 5405
rect 17547 5356 17548 5396
rect 17588 5356 17589 5396
rect 17547 5347 17589 5356
rect 17932 5060 17972 5683
rect 18028 5648 18068 5657
rect 18028 5228 18068 5608
rect 18123 5648 18165 5657
rect 18123 5608 18124 5648
rect 18164 5608 18165 5648
rect 18123 5599 18165 5608
rect 18124 5514 18164 5599
rect 18316 5312 18356 7783
rect 18412 5564 18452 8212
rect 18508 6488 18548 8455
rect 18604 7748 18644 14848
rect 18700 14720 18740 16939
rect 18808 16652 19176 16661
rect 18848 16612 18890 16652
rect 18930 16612 18972 16652
rect 19012 16612 19054 16652
rect 19094 16612 19136 16652
rect 18808 16603 19176 16612
rect 19276 16493 19316 18544
rect 19468 18257 19508 20728
rect 19563 20768 19605 20777
rect 19563 20728 19564 20768
rect 19604 20728 19605 20768
rect 19563 20719 19605 20728
rect 19564 20189 19604 20719
rect 19563 20180 19605 20189
rect 19563 20140 19564 20180
rect 19604 20140 19605 20180
rect 19563 20131 19605 20140
rect 19563 19592 19605 19601
rect 19563 19552 19564 19592
rect 19604 19552 19605 19592
rect 19563 19543 19605 19552
rect 19564 19256 19604 19543
rect 19564 19207 19604 19216
rect 19660 19097 19700 22399
rect 19756 20861 19796 23416
rect 19851 23120 19893 23129
rect 19851 23080 19852 23120
rect 19892 23080 19893 23120
rect 19851 23071 19893 23080
rect 19852 22986 19892 23071
rect 19948 22457 19988 23584
rect 20139 23575 20181 23584
rect 20048 23456 20416 23465
rect 20088 23416 20130 23456
rect 20170 23416 20212 23456
rect 20252 23416 20294 23456
rect 20334 23416 20376 23456
rect 20048 23407 20416 23416
rect 19852 22448 19892 22457
rect 19852 21449 19892 22408
rect 19947 22448 19989 22457
rect 19947 22408 19948 22448
rect 19988 22408 19989 22448
rect 19947 22399 19989 22408
rect 19947 22280 19989 22289
rect 19947 22240 19948 22280
rect 19988 22240 19989 22280
rect 19947 22231 19989 22240
rect 19948 21776 19988 22231
rect 20048 21944 20416 21953
rect 20088 21904 20130 21944
rect 20170 21904 20212 21944
rect 20252 21904 20294 21944
rect 20334 21904 20376 21944
rect 20048 21895 20416 21904
rect 20140 21776 20180 21785
rect 19948 21736 20140 21776
rect 20140 21727 20180 21736
rect 19947 21608 19989 21617
rect 19947 21568 19948 21608
rect 19988 21568 19989 21608
rect 19947 21559 19989 21568
rect 19948 21474 19988 21559
rect 19851 21440 19893 21449
rect 19851 21400 19852 21440
rect 19892 21400 19893 21440
rect 19851 21391 19893 21400
rect 20524 21020 20564 29035
rect 20620 28001 20660 29287
rect 20812 29093 20852 35848
rect 21292 35057 21332 38947
rect 21387 38912 21429 38921
rect 21387 38872 21388 38912
rect 21428 38872 21429 38912
rect 21387 38863 21429 38872
rect 21291 35048 21333 35057
rect 21291 35008 21292 35048
rect 21332 35008 21333 35048
rect 21291 34999 21333 35008
rect 21388 34049 21428 38863
rect 21387 34040 21429 34049
rect 21387 34000 21388 34040
rect 21428 34000 21429 34040
rect 21387 33991 21429 34000
rect 21291 32696 21333 32705
rect 21291 32656 21292 32696
rect 21332 32656 21333 32696
rect 21291 32647 21333 32656
rect 21099 30260 21141 30269
rect 21099 30220 21100 30260
rect 21140 30220 21141 30260
rect 21099 30211 21141 30220
rect 20811 29084 20853 29093
rect 20811 29044 20812 29084
rect 20852 29044 20853 29084
rect 20811 29035 20853 29044
rect 20619 27992 20661 28001
rect 20619 27952 20620 27992
rect 20660 27952 20661 27992
rect 20619 27943 20661 27952
rect 20811 27404 20853 27413
rect 20811 27364 20812 27404
rect 20852 27364 20853 27404
rect 20811 27355 20853 27364
rect 20812 21953 20852 27355
rect 20811 21944 20853 21953
rect 20811 21904 20812 21944
rect 20852 21904 20853 21944
rect 20811 21895 20853 21904
rect 20524 20980 20660 21020
rect 19755 20852 19797 20861
rect 19755 20812 19756 20852
rect 19796 20812 19797 20852
rect 19755 20803 19797 20812
rect 19948 20777 19988 20862
rect 19947 20768 19989 20777
rect 19947 20728 19948 20768
rect 19988 20728 19989 20768
rect 19947 20719 19989 20728
rect 20044 20768 20084 20777
rect 19755 20600 19797 20609
rect 20044 20600 20084 20728
rect 20140 20747 20180 20756
rect 20140 20609 20180 20707
rect 19755 20560 19756 20600
rect 19796 20560 19797 20600
rect 19755 20551 19797 20560
rect 19852 20560 20084 20600
rect 20139 20600 20181 20609
rect 20139 20560 20140 20600
rect 20180 20560 20181 20600
rect 19756 20466 19796 20551
rect 19852 20180 19892 20560
rect 20139 20551 20181 20560
rect 20236 20600 20276 20609
rect 20276 20560 20564 20600
rect 20236 20551 20276 20560
rect 20048 20432 20416 20441
rect 20088 20392 20130 20432
rect 20170 20392 20212 20432
rect 20252 20392 20294 20432
rect 20334 20392 20376 20432
rect 20048 20383 20416 20392
rect 20524 20264 20564 20560
rect 19756 20140 19892 20180
rect 20236 20224 20564 20264
rect 19659 19088 19701 19097
rect 19659 19048 19660 19088
rect 19700 19048 19701 19088
rect 19659 19039 19701 19048
rect 19756 18761 19796 20140
rect 19947 20096 19989 20105
rect 20236 20096 20276 20224
rect 20620 20180 20660 20980
rect 19947 20056 19948 20096
rect 19988 20056 19989 20096
rect 19947 20047 19989 20056
rect 20044 20056 20276 20096
rect 20524 20140 20660 20180
rect 19851 19676 19893 19685
rect 19851 19636 19852 19676
rect 19892 19636 19893 19676
rect 19851 19627 19893 19636
rect 19852 19256 19892 19627
rect 19948 19433 19988 20047
rect 19947 19424 19989 19433
rect 19947 19384 19948 19424
rect 19988 19384 19989 19424
rect 19947 19375 19989 19384
rect 19852 19207 19892 19216
rect 19948 19256 19988 19265
rect 20044 19256 20084 20056
rect 20140 19844 20180 19853
rect 20140 19601 20180 19804
rect 20139 19592 20181 19601
rect 20139 19552 20140 19592
rect 20180 19552 20181 19592
rect 20139 19543 20181 19552
rect 20235 19424 20277 19433
rect 20235 19384 20236 19424
rect 20276 19384 20277 19424
rect 20235 19375 20277 19384
rect 20236 19290 20276 19375
rect 19988 19216 20084 19256
rect 19948 19207 19988 19216
rect 20048 18920 20416 18929
rect 20088 18880 20130 18920
rect 20170 18880 20212 18920
rect 20252 18880 20294 18920
rect 20334 18880 20376 18920
rect 20048 18871 20416 18880
rect 19755 18752 19797 18761
rect 19755 18712 19756 18752
rect 19796 18712 19797 18752
rect 19755 18703 19797 18712
rect 19467 18248 19509 18257
rect 19467 18208 19468 18248
rect 19508 18208 19509 18248
rect 19467 18199 19509 18208
rect 19275 16484 19317 16493
rect 19275 16444 19276 16484
rect 19316 16444 19317 16484
rect 19275 16435 19317 16444
rect 18795 16232 18837 16241
rect 18795 16192 18796 16232
rect 18836 16192 18837 16232
rect 18795 16183 18837 16192
rect 18796 16098 18836 16183
rect 18808 15140 19176 15149
rect 18848 15100 18890 15140
rect 18930 15100 18972 15140
rect 19012 15100 19054 15140
rect 19094 15100 19136 15140
rect 18808 15091 19176 15100
rect 18891 14804 18933 14813
rect 18891 14764 18892 14804
rect 18932 14764 18933 14804
rect 18891 14755 18933 14764
rect 18796 14720 18836 14729
rect 18700 14680 18796 14720
rect 18700 13460 18740 14680
rect 18796 14671 18836 14680
rect 18892 14670 18932 14755
rect 19371 14720 19413 14729
rect 19371 14680 19372 14720
rect 19412 14680 19413 14720
rect 19371 14671 19413 14680
rect 19083 14636 19125 14645
rect 19083 14596 19084 14636
rect 19124 14596 19125 14636
rect 19083 14587 19125 14596
rect 19084 14048 19124 14587
rect 19084 13889 19124 14008
rect 19275 14048 19317 14057
rect 19275 14008 19276 14048
rect 19316 14008 19317 14048
rect 19275 13999 19317 14008
rect 19083 13880 19125 13889
rect 19083 13840 19084 13880
rect 19124 13840 19125 13880
rect 19083 13831 19125 13840
rect 18808 13628 19176 13637
rect 18848 13588 18890 13628
rect 18930 13588 18972 13628
rect 19012 13588 19054 13628
rect 19094 13588 19136 13628
rect 18808 13579 19176 13588
rect 18891 13460 18933 13469
rect 18700 13420 18836 13460
rect 18699 13292 18741 13301
rect 18699 13252 18700 13292
rect 18740 13252 18741 13292
rect 18699 13243 18741 13252
rect 18700 12536 18740 13243
rect 18700 12487 18740 12496
rect 18796 12368 18836 13420
rect 18891 13420 18892 13460
rect 18932 13420 18933 13460
rect 18891 13411 18933 13420
rect 18700 12328 18836 12368
rect 18892 13292 18932 13411
rect 19276 13376 19316 13999
rect 19372 13553 19412 14671
rect 19371 13544 19413 13553
rect 19371 13504 19372 13544
rect 19412 13504 19413 13544
rect 19371 13495 19413 13504
rect 18700 11453 18740 12328
rect 18892 12293 18932 13252
rect 18988 13336 19412 13376
rect 18988 13292 19028 13336
rect 18988 13243 19028 13252
rect 18891 12284 18933 12293
rect 18891 12244 18892 12284
rect 18932 12244 18933 12284
rect 18891 12235 18933 12244
rect 18808 12116 19176 12125
rect 18848 12076 18890 12116
rect 18930 12076 18972 12116
rect 19012 12076 19054 12116
rect 19094 12076 19136 12116
rect 18808 12067 19176 12076
rect 18987 11948 19029 11957
rect 18987 11908 18988 11948
rect 19028 11908 19029 11948
rect 18987 11899 19029 11908
rect 18891 11864 18933 11873
rect 18891 11824 18892 11864
rect 18932 11824 18933 11864
rect 18891 11815 18933 11824
rect 18892 11780 18932 11815
rect 18892 11729 18932 11740
rect 18988 11780 19028 11899
rect 19275 11864 19317 11873
rect 19275 11824 19276 11864
rect 19316 11824 19317 11864
rect 19275 11815 19317 11824
rect 18988 11731 19028 11740
rect 18699 11444 18741 11453
rect 18699 11404 18700 11444
rect 18740 11404 18741 11444
rect 18699 11395 18741 11404
rect 18699 11024 18741 11033
rect 18699 10984 18700 11024
rect 18740 10984 18741 11024
rect 18699 10975 18741 10984
rect 18700 10890 18740 10975
rect 18808 10604 19176 10613
rect 18848 10564 18890 10604
rect 18930 10564 18972 10604
rect 19012 10564 19054 10604
rect 19094 10564 19136 10604
rect 18808 10555 19176 10564
rect 18699 10520 18741 10529
rect 18699 10480 18700 10520
rect 18740 10480 18741 10520
rect 18699 10471 18741 10480
rect 18700 10184 18740 10471
rect 19179 10268 19221 10277
rect 19179 10228 19180 10268
rect 19220 10228 19221 10268
rect 19179 10219 19221 10228
rect 19276 10268 19316 11815
rect 19276 10219 19316 10228
rect 18700 10135 18740 10144
rect 19180 10134 19220 10219
rect 18795 10100 18837 10109
rect 18795 10060 18796 10100
rect 18836 10060 18837 10100
rect 18795 10051 18837 10060
rect 18796 9260 18836 10051
rect 19083 9680 19125 9689
rect 19083 9640 19084 9680
rect 19124 9640 19125 9680
rect 19083 9631 19125 9640
rect 19084 9546 19124 9631
rect 18700 9220 18836 9260
rect 18892 9512 18932 9521
rect 18892 9260 18932 9472
rect 19372 9437 19412 13336
rect 19468 13208 19508 18199
rect 20235 17996 20277 18005
rect 20235 17956 20236 17996
rect 20276 17956 20277 17996
rect 20235 17947 20277 17956
rect 19851 17744 19893 17753
rect 19851 17704 19852 17744
rect 19892 17704 19893 17744
rect 19851 17695 19893 17704
rect 20236 17744 20276 17947
rect 20236 17695 20276 17704
rect 19564 16988 19604 16999
rect 19564 16913 19604 16948
rect 19659 16988 19701 16997
rect 19659 16948 19660 16988
rect 19700 16948 19701 16988
rect 19659 16939 19701 16948
rect 19563 16904 19605 16913
rect 19563 16864 19564 16904
rect 19604 16864 19605 16904
rect 19563 16855 19605 16864
rect 19660 16854 19700 16939
rect 19852 16064 19892 17695
rect 20048 17408 20416 17417
rect 20088 17368 20130 17408
rect 20170 17368 20212 17408
rect 20252 17368 20294 17408
rect 20334 17368 20376 17408
rect 20048 17359 20416 17368
rect 20044 17072 20084 17081
rect 20044 16409 20084 17032
rect 20140 17053 20180 17062
rect 20140 16484 20180 17013
rect 20236 16484 20276 16493
rect 20140 16444 20236 16484
rect 20236 16435 20276 16444
rect 20043 16400 20085 16409
rect 20043 16360 20044 16400
rect 20084 16360 20085 16400
rect 20043 16351 20085 16360
rect 20044 16232 20084 16241
rect 20044 16064 20084 16192
rect 19852 16024 20084 16064
rect 19755 15980 19797 15989
rect 19755 15940 19756 15980
rect 19796 15940 19797 15980
rect 19755 15931 19797 15940
rect 19756 15560 19796 15931
rect 19756 15511 19796 15520
rect 19852 15392 19892 16024
rect 20048 15896 20416 15905
rect 20088 15856 20130 15896
rect 20170 15856 20212 15896
rect 20252 15856 20294 15896
rect 20334 15856 20376 15896
rect 20048 15847 20416 15856
rect 19468 11705 19508 13168
rect 19756 15352 19892 15392
rect 19756 12545 19796 15352
rect 19948 15308 19988 15317
rect 19852 15268 19948 15308
rect 19852 14734 19892 15268
rect 19948 15259 19988 15268
rect 20524 15140 20564 20140
rect 20619 19424 20661 19433
rect 20619 19384 20620 19424
rect 20660 19384 20661 19424
rect 20619 19375 20661 19384
rect 20620 17417 20660 19375
rect 20619 17408 20661 17417
rect 20619 17368 20620 17408
rect 20660 17368 20661 17408
rect 20619 17359 20661 17368
rect 21100 15905 21140 30211
rect 21195 27572 21237 27581
rect 21195 27532 21196 27572
rect 21236 27532 21237 27572
rect 21195 27523 21237 27532
rect 21196 18425 21236 27523
rect 21292 19937 21332 32647
rect 21387 29252 21429 29261
rect 21387 29212 21388 29252
rect 21428 29212 21429 29252
rect 21387 29203 21429 29212
rect 21388 29009 21428 29203
rect 21387 29000 21429 29009
rect 21387 28960 21388 29000
rect 21428 28960 21429 29000
rect 21387 28951 21429 28960
rect 21387 25724 21429 25733
rect 21387 25684 21388 25724
rect 21428 25684 21429 25724
rect 21387 25675 21429 25684
rect 21388 25481 21428 25675
rect 21387 25472 21429 25481
rect 21387 25432 21388 25472
rect 21428 25432 21429 25472
rect 21387 25423 21429 25432
rect 21387 24296 21429 24305
rect 21387 24256 21388 24296
rect 21428 24256 21429 24296
rect 21387 24247 21429 24256
rect 21388 23969 21428 24247
rect 21387 23960 21429 23969
rect 21387 23920 21388 23960
rect 21428 23920 21429 23960
rect 21387 23911 21429 23920
rect 21291 19928 21333 19937
rect 21291 19888 21292 19928
rect 21332 19888 21333 19928
rect 21291 19879 21333 19888
rect 21195 18416 21237 18425
rect 21195 18376 21196 18416
rect 21236 18376 21237 18416
rect 21195 18367 21237 18376
rect 21099 15896 21141 15905
rect 21099 15856 21100 15896
rect 21140 15856 21141 15896
rect 21099 15847 21141 15856
rect 20524 15100 20660 15140
rect 19852 14685 19892 14694
rect 20044 14552 20084 14561
rect 19852 14512 20044 14552
rect 19755 12536 19797 12545
rect 19755 12496 19756 12536
rect 19796 12496 19797 12536
rect 19755 12487 19797 12496
rect 19467 11696 19509 11705
rect 19467 11656 19468 11696
rect 19508 11656 19509 11696
rect 19467 11647 19509 11656
rect 19468 11562 19508 11647
rect 19756 11537 19796 12487
rect 19755 11528 19797 11537
rect 19755 11488 19756 11528
rect 19796 11488 19797 11528
rect 19755 11479 19797 11488
rect 19563 11192 19605 11201
rect 19563 11152 19564 11192
rect 19604 11152 19605 11192
rect 19563 11143 19605 11152
rect 19371 9428 19413 9437
rect 19371 9388 19372 9428
rect 19412 9388 19413 9428
rect 19371 9379 19413 9388
rect 19564 9428 19604 11143
rect 19756 11024 19796 11479
rect 19852 11201 19892 14512
rect 20044 14503 20084 14512
rect 20048 14384 20416 14393
rect 20088 14344 20130 14384
rect 20170 14344 20212 14384
rect 20252 14344 20294 14384
rect 20334 14344 20376 14384
rect 20048 14335 20416 14344
rect 19948 13213 19988 13222
rect 19948 12704 19988 13173
rect 20140 13049 20180 13134
rect 20139 13040 20181 13049
rect 20139 13000 20140 13040
rect 20180 13000 20181 13040
rect 20139 12991 20181 13000
rect 20048 12872 20416 12881
rect 20088 12832 20130 12872
rect 20170 12832 20212 12872
rect 20252 12832 20294 12872
rect 20334 12832 20376 12872
rect 20048 12823 20416 12832
rect 20140 12704 20180 12713
rect 19948 12664 20140 12704
rect 20140 12655 20180 12664
rect 19947 12536 19989 12545
rect 19947 12496 19948 12536
rect 19988 12496 19989 12536
rect 19947 12487 19989 12496
rect 19948 12402 19988 12487
rect 19948 11701 19988 11710
rect 19851 11192 19893 11201
rect 19851 11152 19852 11192
rect 19892 11152 19893 11192
rect 19948 11192 19988 11661
rect 20140 11528 20180 11537
rect 20180 11488 20564 11528
rect 20140 11479 20180 11488
rect 20048 11360 20416 11369
rect 20088 11320 20130 11360
rect 20170 11320 20212 11360
rect 20252 11320 20294 11360
rect 20334 11320 20376 11360
rect 20048 11311 20416 11320
rect 20140 11192 20180 11201
rect 19948 11152 20140 11192
rect 19851 11143 19893 11152
rect 20140 11143 20180 11152
rect 19948 11024 19988 11033
rect 19756 10984 19948 11024
rect 19948 10975 19988 10984
rect 19659 10688 19701 10697
rect 19659 10648 19660 10688
rect 19700 10648 19701 10688
rect 19659 10639 19701 10648
rect 19564 9379 19604 9388
rect 19660 10184 19700 10639
rect 19371 9260 19413 9269
rect 18892 9220 19316 9260
rect 18700 8840 18740 9220
rect 18808 9092 19176 9101
rect 18848 9052 18890 9092
rect 18930 9052 18972 9092
rect 19012 9052 19054 9092
rect 19094 9052 19136 9092
rect 18808 9043 19176 9052
rect 18700 8800 18836 8840
rect 18700 8672 18740 8681
rect 18700 8345 18740 8632
rect 18699 8336 18741 8345
rect 18699 8296 18700 8336
rect 18740 8296 18741 8336
rect 18699 8287 18741 8296
rect 18796 8084 18836 8800
rect 19276 8681 19316 9220
rect 19371 9220 19372 9260
rect 19412 9220 19413 9260
rect 19371 9211 19413 9220
rect 19372 9126 19412 9211
rect 19275 8672 19317 8681
rect 19275 8632 19276 8672
rect 19316 8632 19317 8672
rect 19275 8623 19317 8632
rect 18700 8044 18836 8084
rect 19660 8084 19700 10144
rect 19756 10184 19796 10193
rect 19756 9689 19796 10144
rect 19947 10184 19989 10193
rect 19947 10144 19948 10184
rect 19988 10144 19989 10184
rect 19947 10135 19989 10144
rect 19755 9680 19797 9689
rect 19755 9640 19756 9680
rect 19796 9640 19797 9680
rect 19755 9631 19797 9640
rect 19948 8924 19988 10135
rect 20048 9848 20416 9857
rect 20088 9808 20130 9848
rect 20170 9808 20212 9848
rect 20252 9808 20294 9848
rect 20334 9808 20376 9848
rect 20048 9799 20416 9808
rect 20140 8924 20180 8933
rect 19948 8884 20140 8924
rect 20140 8875 20180 8884
rect 19947 8672 19989 8681
rect 19947 8632 19948 8672
rect 19988 8632 19989 8672
rect 19947 8623 19989 8632
rect 19948 8538 19988 8623
rect 20048 8336 20416 8345
rect 20088 8296 20130 8336
rect 20170 8296 20212 8336
rect 20252 8296 20294 8336
rect 20334 8296 20376 8336
rect 20048 8287 20416 8296
rect 19948 8084 19988 8093
rect 19660 8044 19892 8084
rect 18700 8000 18740 8044
rect 18700 7925 18740 7960
rect 19275 8000 19317 8009
rect 19275 7960 19276 8000
rect 19316 7960 19317 8000
rect 19275 7951 19317 7960
rect 19756 7986 19796 7995
rect 18699 7916 18741 7925
rect 18699 7876 18700 7916
rect 18740 7876 18741 7916
rect 18699 7867 18741 7876
rect 18796 7916 18836 7925
rect 18700 7836 18740 7867
rect 18796 7757 18836 7876
rect 18795 7748 18837 7757
rect 18604 7708 18740 7748
rect 18603 7076 18645 7085
rect 18603 7036 18604 7076
rect 18644 7036 18645 7076
rect 18603 7027 18645 7036
rect 18508 5732 18548 6448
rect 18604 6488 18644 7027
rect 18604 6439 18644 6448
rect 18508 5683 18548 5692
rect 18604 5648 18644 5657
rect 18604 5564 18644 5608
rect 18412 5524 18644 5564
rect 18316 5272 18452 5312
rect 18028 5188 18356 5228
rect 18316 5144 18356 5188
rect 18316 5095 18356 5104
rect 18219 5060 18261 5069
rect 17836 5020 18164 5060
rect 17836 4817 17876 5020
rect 18124 4976 18164 5020
rect 18219 5020 18220 5060
rect 18260 5020 18261 5060
rect 18219 5011 18261 5020
rect 18124 4927 18164 4936
rect 17835 4808 17877 4817
rect 18220 4808 18260 5011
rect 17835 4768 17836 4808
rect 17876 4768 17877 4808
rect 17835 4759 17877 4768
rect 18124 4768 18260 4808
rect 17739 4472 17781 4481
rect 17739 4432 17740 4472
rect 17780 4432 17781 4472
rect 17739 4423 17781 4432
rect 17356 4339 17396 4348
rect 17740 4388 17780 4423
rect 17164 3464 17204 4339
rect 17740 4337 17780 4348
rect 17547 4220 17589 4229
rect 17547 4180 17548 4220
rect 17588 4180 17589 4220
rect 17547 4171 17589 4180
rect 17548 4086 17588 4171
rect 17739 4136 17781 4145
rect 17739 4096 17740 4136
rect 17780 4096 17781 4136
rect 17739 4087 17781 4096
rect 17164 3415 17204 3424
rect 17259 3464 17301 3473
rect 17259 3424 17260 3464
rect 17300 3424 17301 3464
rect 17259 3415 17301 3424
rect 17740 3464 17780 4087
rect 17836 3725 17876 4759
rect 17932 4220 17972 4229
rect 18124 4220 18164 4768
rect 18412 4724 18452 5272
rect 18604 4985 18644 5070
rect 18700 5069 18740 7708
rect 18795 7708 18796 7748
rect 18836 7708 18837 7748
rect 18795 7699 18837 7708
rect 18808 7580 19176 7589
rect 18848 7540 18890 7580
rect 18930 7540 18972 7580
rect 19012 7540 19054 7580
rect 19094 7540 19136 7580
rect 18808 7531 19176 7540
rect 19084 6488 19124 6497
rect 19276 6488 19316 7951
rect 19756 7412 19796 7946
rect 19660 7372 19796 7412
rect 19371 7160 19413 7169
rect 19371 7120 19372 7160
rect 19412 7120 19413 7160
rect 19371 7111 19413 7120
rect 19372 7026 19412 7111
rect 19563 6992 19605 7001
rect 19563 6952 19564 6992
rect 19604 6952 19605 6992
rect 19563 6943 19605 6952
rect 19564 6858 19604 6943
rect 19124 6448 19316 6488
rect 19564 6474 19604 6483
rect 19084 6439 19124 6448
rect 18808 6068 19176 6077
rect 18848 6028 18890 6068
rect 18930 6028 18972 6068
rect 19012 6028 19054 6068
rect 19094 6028 19136 6068
rect 18808 6019 19176 6028
rect 19564 5816 19604 6434
rect 19468 5776 19604 5816
rect 19084 5648 19124 5657
rect 19124 5608 19316 5648
rect 19084 5599 19124 5608
rect 18699 5060 18741 5069
rect 18699 5020 18700 5060
rect 18740 5020 18741 5060
rect 18699 5011 18741 5020
rect 18603 4976 18645 4985
rect 18603 4936 18604 4976
rect 18644 4936 18645 4976
rect 18603 4927 18645 4936
rect 18412 4684 18740 4724
rect 17972 4180 18164 4220
rect 18700 4220 18740 4684
rect 18808 4556 19176 4565
rect 18848 4516 18890 4556
rect 18930 4516 18972 4556
rect 19012 4516 19054 4556
rect 19094 4516 19136 4556
rect 18808 4507 19176 4516
rect 18795 4388 18837 4397
rect 18795 4348 18796 4388
rect 18836 4348 18837 4388
rect 18795 4339 18837 4348
rect 17932 4171 17972 4180
rect 18700 4171 18740 4180
rect 18796 4220 18836 4339
rect 18796 4171 18836 4180
rect 18220 4136 18260 4145
rect 18124 4096 18220 4136
rect 17835 3716 17877 3725
rect 17835 3676 17836 3716
rect 17876 3676 17877 3716
rect 17835 3667 17877 3676
rect 18027 3716 18069 3725
rect 18027 3676 18028 3716
rect 18068 3676 18069 3716
rect 18027 3667 18069 3676
rect 17931 3548 17973 3557
rect 17931 3508 17932 3548
rect 17972 3508 17973 3548
rect 17931 3499 17973 3508
rect 17740 3415 17780 3424
rect 17260 3330 17300 3415
rect 17355 1196 17397 1205
rect 17355 1156 17356 1196
rect 17396 1156 17397 1196
rect 17355 1147 17397 1156
rect 17739 1196 17781 1205
rect 17739 1156 17740 1196
rect 17780 1156 17781 1196
rect 17739 1147 17781 1156
rect 17356 1062 17396 1147
rect 17164 953 17204 1038
rect 17163 944 17205 953
rect 17163 904 17164 944
rect 17204 904 17205 944
rect 17163 895 17205 904
rect 17355 944 17397 953
rect 17355 904 17356 944
rect 17396 904 17397 944
rect 17355 895 17397 904
rect 17068 736 17204 776
rect 17164 80 17204 736
rect 17356 80 17396 895
rect 17547 860 17589 869
rect 17547 820 17548 860
rect 17588 820 17589 860
rect 17547 811 17589 820
rect 17548 80 17588 811
rect 17740 80 17780 1147
rect 17932 1037 17972 3499
rect 18028 1952 18068 3667
rect 18124 2120 18164 4096
rect 18220 4087 18260 4096
rect 18316 4136 18356 4147
rect 19276 4145 19316 5608
rect 18316 4061 18356 4096
rect 19275 4136 19317 4145
rect 19275 4096 19276 4136
rect 19316 4096 19317 4136
rect 19275 4087 19317 4096
rect 18315 4052 18357 4061
rect 18315 4012 18316 4052
rect 18356 4012 18357 4052
rect 18315 4003 18357 4012
rect 18507 4052 18549 4061
rect 18507 4012 18508 4052
rect 18548 4012 18549 4052
rect 18507 4003 18549 4012
rect 18412 3557 18452 3642
rect 18411 3548 18453 3557
rect 18411 3508 18412 3548
rect 18452 3508 18453 3548
rect 18411 3499 18453 3508
rect 18268 3422 18308 3431
rect 18268 3380 18308 3382
rect 18268 3340 18452 3380
rect 18412 2876 18452 3340
rect 18412 2827 18452 2836
rect 18220 2633 18260 2718
rect 18219 2624 18261 2633
rect 18219 2584 18220 2624
rect 18260 2584 18261 2624
rect 18219 2575 18261 2584
rect 18508 2540 18548 4003
rect 19276 4002 19316 4087
rect 18603 3968 18645 3977
rect 18603 3928 18604 3968
rect 18644 3928 18645 3968
rect 18603 3919 18645 3928
rect 18604 3464 18644 3919
rect 19468 3641 19508 5776
rect 19564 5653 19604 5662
rect 19467 3632 19509 3641
rect 19467 3592 19468 3632
rect 19508 3592 19509 3632
rect 19467 3583 19509 3592
rect 18604 3415 18644 3424
rect 18808 3044 19176 3053
rect 18848 3004 18890 3044
rect 18930 3004 18972 3044
rect 19012 3004 19054 3044
rect 19094 3004 19136 3044
rect 18808 2995 19176 3004
rect 19564 2885 19604 5613
rect 19660 5228 19700 7372
rect 19756 7244 19796 7253
rect 19756 6656 19796 7204
rect 19756 6607 19796 6616
rect 19852 6152 19892 8044
rect 19948 7421 19988 8044
rect 19947 7412 19989 7421
rect 19947 7372 19948 7412
rect 19988 7372 19989 7412
rect 19947 7363 19989 7372
rect 20048 6824 20416 6833
rect 20088 6784 20130 6824
rect 20170 6784 20212 6824
rect 20252 6784 20294 6824
rect 20334 6784 20376 6824
rect 20048 6775 20416 6784
rect 20121 6401 20161 6410
rect 19947 6320 19989 6329
rect 20121 6320 20161 6361
rect 20524 6320 20564 11488
rect 19947 6280 19948 6320
rect 19988 6280 19989 6320
rect 19947 6271 19989 6280
rect 20044 6280 20161 6320
rect 20236 6280 20564 6320
rect 19948 6186 19988 6271
rect 19756 6112 19892 6152
rect 19756 5825 19796 6112
rect 20044 6068 20084 6280
rect 20236 6236 20276 6280
rect 19852 6028 20084 6068
rect 20140 6196 20276 6236
rect 19755 5816 19797 5825
rect 19755 5776 19756 5816
rect 19796 5776 19797 5816
rect 19755 5767 19797 5776
rect 19756 5564 19796 5573
rect 19852 5564 19892 6028
rect 20140 5743 20180 6196
rect 20140 5694 20180 5703
rect 19796 5524 19892 5564
rect 19756 5515 19796 5524
rect 19947 5480 19989 5489
rect 19947 5440 19948 5480
rect 19988 5440 19989 5480
rect 19947 5431 19989 5440
rect 19948 5346 19988 5431
rect 20048 5312 20416 5321
rect 20088 5272 20130 5312
rect 20170 5272 20212 5312
rect 20252 5272 20294 5312
rect 20334 5272 20376 5312
rect 20048 5263 20416 5272
rect 19660 5188 19988 5228
rect 19948 5060 19988 5188
rect 20044 5060 20084 5069
rect 19948 5020 20044 5060
rect 20044 5011 20084 5020
rect 19852 4976 19892 4985
rect 19852 4817 19892 4936
rect 20523 4892 20565 4901
rect 20523 4852 20524 4892
rect 20564 4852 20565 4892
rect 20523 4843 20565 4852
rect 19851 4808 19893 4817
rect 19851 4768 19852 4808
rect 19892 4768 19893 4808
rect 19851 4759 19893 4768
rect 19756 4141 19796 4150
rect 19756 3389 19796 4101
rect 19852 3464 19892 4759
rect 20524 4313 20564 4843
rect 20523 4304 20565 4313
rect 20523 4264 20524 4304
rect 20564 4264 20565 4304
rect 20523 4255 20565 4264
rect 19947 4220 19989 4229
rect 19947 4180 19948 4220
rect 19988 4180 19989 4220
rect 19947 4171 19989 4180
rect 19948 4052 19988 4171
rect 19948 4003 19988 4012
rect 20048 3800 20416 3809
rect 20088 3760 20130 3800
rect 20170 3760 20212 3800
rect 20252 3760 20294 3800
rect 20334 3760 20376 3800
rect 20048 3751 20416 3760
rect 20043 3632 20085 3641
rect 20043 3592 20044 3632
rect 20084 3592 20085 3632
rect 20043 3583 20085 3592
rect 20044 3498 20084 3583
rect 19755 3380 19797 3389
rect 19755 3340 19756 3380
rect 19796 3340 19797 3380
rect 19755 3331 19797 3340
rect 19563 2876 19605 2885
rect 19563 2836 19564 2876
rect 19604 2836 19605 2876
rect 19563 2827 19605 2836
rect 18603 2708 18645 2717
rect 18603 2668 18604 2708
rect 18644 2668 18645 2708
rect 18603 2659 18645 2668
rect 18604 2624 18644 2659
rect 18604 2573 18644 2584
rect 19852 2624 19892 3424
rect 19947 3380 19989 3389
rect 19947 3340 19948 3380
rect 19988 3340 19989 3380
rect 19947 3331 19989 3340
rect 18412 2500 18548 2540
rect 18220 2120 18260 2129
rect 18124 2080 18220 2120
rect 18220 2071 18260 2080
rect 18028 1709 18068 1912
rect 18027 1700 18069 1709
rect 18027 1660 18028 1700
rect 18068 1660 18069 1700
rect 18027 1651 18069 1660
rect 18412 1196 18452 2500
rect 18508 1952 18548 1961
rect 18508 1289 18548 1912
rect 19756 1952 19796 1961
rect 19852 1952 19892 2584
rect 19948 2120 19988 3331
rect 20043 2876 20085 2885
rect 20043 2836 20044 2876
rect 20084 2836 20085 2876
rect 20043 2827 20085 2836
rect 20044 2742 20084 2827
rect 20048 2288 20416 2297
rect 20088 2248 20130 2288
rect 20170 2248 20212 2288
rect 20252 2248 20294 2288
rect 20334 2248 20376 2288
rect 20048 2239 20416 2248
rect 19948 2071 19988 2080
rect 19796 1912 19892 1952
rect 19756 1903 19796 1912
rect 18808 1532 19176 1541
rect 18848 1492 18890 1532
rect 18930 1492 18972 1532
rect 19012 1492 19054 1532
rect 19094 1492 19136 1532
rect 18808 1483 19176 1492
rect 18891 1364 18933 1373
rect 18891 1324 18892 1364
rect 18932 1324 18933 1364
rect 18891 1315 18933 1324
rect 18507 1280 18549 1289
rect 18507 1240 18508 1280
rect 18548 1240 18549 1280
rect 18507 1231 18549 1240
rect 18412 1147 18452 1156
rect 17931 1028 17973 1037
rect 17931 988 17932 1028
rect 17972 988 17973 1028
rect 17931 979 17973 988
rect 18220 944 18260 953
rect 17931 692 17973 701
rect 17931 652 17932 692
rect 17972 652 17973 692
rect 17931 643 17973 652
rect 18123 692 18165 701
rect 18123 652 18124 692
rect 18164 652 18165 692
rect 18123 643 18165 652
rect 17932 80 17972 643
rect 18124 80 18164 643
rect 18220 365 18260 904
rect 18315 692 18357 701
rect 18315 652 18316 692
rect 18356 652 18357 692
rect 18315 643 18357 652
rect 18507 692 18549 701
rect 18507 652 18508 692
rect 18548 652 18549 692
rect 18507 643 18549 652
rect 18219 356 18261 365
rect 18219 316 18220 356
rect 18260 316 18261 356
rect 18219 307 18261 316
rect 18316 80 18356 643
rect 18508 80 18548 643
rect 18699 524 18741 533
rect 18699 484 18700 524
rect 18740 484 18741 524
rect 18699 475 18741 484
rect 18700 80 18740 475
rect 18892 80 18932 1315
rect 20620 1289 20660 15100
rect 20715 13376 20757 13385
rect 20715 13336 20716 13376
rect 20756 13336 20757 13376
rect 20715 13327 20757 13336
rect 20716 10445 20756 13327
rect 20715 10436 20757 10445
rect 20715 10396 20716 10436
rect 20756 10396 20757 10436
rect 20715 10387 20757 10396
rect 21387 4808 21429 4817
rect 21387 4768 21388 4808
rect 21428 4768 21429 4808
rect 21387 4759 21429 4768
rect 21388 4481 21428 4759
rect 21387 4472 21429 4481
rect 21387 4432 21388 4472
rect 21428 4432 21429 4472
rect 21387 4423 21429 4432
rect 19083 1280 19125 1289
rect 19083 1240 19084 1280
rect 19124 1240 19125 1280
rect 19083 1231 19125 1240
rect 20619 1280 20661 1289
rect 20619 1240 20620 1280
rect 20660 1240 20661 1280
rect 20619 1231 20661 1240
rect 19084 80 19124 1231
rect 20048 776 20416 785
rect 20088 736 20130 776
rect 20170 736 20212 776
rect 20252 736 20294 776
rect 20334 736 20376 776
rect 20048 727 20416 736
rect 19467 692 19509 701
rect 19467 652 19468 692
rect 19508 652 19509 692
rect 19467 643 19509 652
rect 19275 608 19317 617
rect 19275 568 19276 608
rect 19316 568 19317 608
rect 19275 559 19317 568
rect 19276 80 19316 559
rect 19468 80 19508 643
rect 1784 0 1864 80
rect 1976 0 2056 80
rect 2168 0 2248 80
rect 2360 0 2440 80
rect 2552 0 2632 80
rect 2744 0 2824 80
rect 2936 0 3016 80
rect 3128 0 3208 80
rect 3320 0 3400 80
rect 3512 0 3592 80
rect 3704 0 3784 80
rect 3896 0 3976 80
rect 4088 0 4168 80
rect 4280 0 4360 80
rect 4472 0 4552 80
rect 4664 0 4744 80
rect 4856 0 4936 80
rect 5048 0 5128 80
rect 5240 0 5320 80
rect 5432 0 5512 80
rect 5624 0 5704 80
rect 5816 0 5896 80
rect 6008 0 6088 80
rect 6200 0 6280 80
rect 6392 0 6472 80
rect 6584 0 6664 80
rect 6776 0 6856 80
rect 6968 0 7048 80
rect 7160 0 7240 80
rect 7352 0 7432 80
rect 7544 0 7624 80
rect 7736 0 7816 80
rect 7928 0 8008 80
rect 8120 0 8200 80
rect 8312 0 8392 80
rect 8504 0 8584 80
rect 8696 0 8776 80
rect 8888 0 8968 80
rect 9080 0 9160 80
rect 9272 0 9352 80
rect 9464 0 9544 80
rect 9656 0 9736 80
rect 9848 0 9928 80
rect 10040 0 10120 80
rect 10232 0 10312 80
rect 10424 0 10504 80
rect 10616 0 10696 80
rect 10808 0 10888 80
rect 11000 0 11080 80
rect 11192 0 11272 80
rect 11384 0 11464 80
rect 11576 0 11656 80
rect 11768 0 11848 80
rect 11960 0 12040 80
rect 12152 0 12232 80
rect 12344 0 12424 80
rect 12536 0 12616 80
rect 12728 0 12808 80
rect 12920 0 13000 80
rect 13112 0 13192 80
rect 13304 0 13384 80
rect 13496 0 13576 80
rect 13688 0 13768 80
rect 13880 0 13960 80
rect 14072 0 14152 80
rect 14264 0 14344 80
rect 14456 0 14536 80
rect 14648 0 14728 80
rect 14840 0 14920 80
rect 15032 0 15112 80
rect 15224 0 15304 80
rect 15416 0 15496 80
rect 15608 0 15688 80
rect 15800 0 15880 80
rect 15992 0 16072 80
rect 16184 0 16264 80
rect 16376 0 16456 80
rect 16568 0 16648 80
rect 16760 0 16840 80
rect 16952 0 17032 80
rect 17144 0 17224 80
rect 17336 0 17416 80
rect 17528 0 17608 80
rect 17720 0 17800 80
rect 17912 0 17992 80
rect 18104 0 18184 80
rect 18296 0 18376 80
rect 18488 0 18568 80
rect 18680 0 18760 80
rect 18872 0 18952 80
rect 19064 0 19144 80
rect 19256 0 19336 80
rect 19448 0 19528 80
<< via2 >>
rect 1324 40972 1364 41012
rect 1324 40720 1364 40760
rect 1324 40300 1364 40340
rect 1324 39544 1364 39584
rect 1132 39460 1172 39500
rect 1132 39040 1172 39080
rect 1324 38956 1364 38996
rect 1324 38452 1364 38492
rect 1612 42904 1652 42944
rect 1804 42904 1844 42944
rect 1804 42316 1844 42356
rect 1612 42232 1652 42272
rect 1516 40972 1556 41012
rect 1516 40468 1556 40508
rect 1516 40300 1556 40340
rect 1708 41140 1748 41180
rect 1900 41140 1940 41180
rect 1804 40384 1844 40424
rect 1516 39544 1556 39584
rect 1516 39040 1556 39080
rect 1708 38704 1748 38744
rect 1612 38452 1652 38492
rect 1708 38368 1748 38408
rect 1900 40300 1940 40340
rect 2092 41308 2132 41348
rect 2092 40804 2132 40844
rect 1132 37024 1172 37064
rect 1228 36520 1268 36560
rect 1132 36184 1172 36224
rect 1612 37696 1652 37736
rect 1612 36100 1652 36140
rect 1420 35428 1460 35468
rect 1420 35260 1460 35300
rect 1516 34672 1556 34712
rect 1804 37108 1844 37148
rect 2284 40636 2324 40676
rect 2284 40468 2324 40508
rect 2188 40384 2228 40424
rect 2284 39880 2324 39920
rect 2092 39376 2132 39416
rect 1996 39124 2036 39164
rect 1996 38956 2036 38996
rect 2188 38536 2228 38576
rect 2092 38284 2132 38324
rect 1996 37612 2036 37652
rect 1996 37024 2036 37064
rect 2092 36520 2132 36560
rect 2092 36268 2132 36308
rect 1996 35848 2036 35888
rect 1900 35596 1940 35636
rect 2572 41812 2612 41852
rect 2668 41644 2708 41684
rect 2572 39628 2612 39668
rect 2572 39376 2612 39416
rect 2476 39208 2516 39248
rect 2476 38536 2516 38576
rect 2476 38200 2516 38240
rect 2860 40636 2900 40676
rect 3052 42400 3092 42440
rect 3148 41644 3188 41684
rect 3436 42148 3476 42188
rect 2956 39796 2996 39836
rect 2860 39376 2900 39416
rect 3052 39712 3092 39752
rect 3340 41140 3380 41180
rect 3244 40300 3284 40340
rect 3724 42484 3764 42524
rect 4492 42316 4532 42356
rect 4300 42232 4340 42272
rect 4204 41728 4244 41768
rect 4108 41476 4148 41516
rect 3628 41140 3668 41180
rect 3724 41056 3764 41096
rect 3916 40972 3956 41012
rect 3688 40804 3728 40844
rect 3770 40804 3810 40844
rect 3852 40804 3892 40844
rect 3934 40804 3974 40844
rect 4016 40804 4056 40844
rect 3532 40384 3572 40424
rect 3820 40384 3860 40424
rect 3436 39376 3476 39416
rect 2956 38872 2996 38912
rect 2860 38368 2900 38408
rect 3148 38704 3188 38744
rect 2668 38116 2708 38156
rect 2764 37780 2804 37820
rect 2956 38116 2996 38156
rect 4012 39628 4052 39668
rect 3724 39460 3764 39500
rect 3688 39292 3728 39332
rect 3770 39292 3810 39332
rect 3852 39292 3892 39332
rect 3934 39292 3974 39332
rect 4016 39292 4056 39332
rect 4108 39124 4148 39164
rect 3628 39040 3668 39080
rect 3628 38704 3668 38744
rect 3628 38368 3668 38408
rect 4300 39628 4340 39668
rect 4108 38116 4148 38156
rect 2476 37696 2516 37736
rect 2380 36940 2420 36980
rect 2476 36268 2516 36308
rect 2188 36100 2228 36140
rect 2092 35512 2132 35552
rect 1900 35260 1940 35300
rect 1420 34420 1460 34460
rect 1324 34252 1364 34292
rect 940 32992 980 33032
rect 172 31816 212 31856
rect 76 23584 116 23624
rect 1420 32320 1460 32360
rect 1036 32068 1076 32108
rect 1324 31480 1364 31520
rect 1324 30304 1364 30344
rect 1324 29800 1364 29840
rect 1612 34420 1652 34460
rect 1900 34420 1940 34460
rect 1804 34252 1844 34292
rect 1900 33328 1940 33368
rect 2476 35596 2516 35636
rect 2764 37612 2804 37652
rect 2764 36604 2804 36644
rect 2284 33160 2324 33200
rect 2092 32656 2132 32696
rect 1804 32152 1844 32192
rect 2284 32320 2324 32360
rect 2476 33664 2516 33704
rect 2476 33328 2516 33368
rect 1612 31480 1652 31520
rect 1708 30640 1748 30680
rect 1612 30556 1652 30596
rect 1516 28456 1556 28496
rect 1228 27028 1268 27068
rect 1708 28372 1748 28412
rect 1612 28288 1652 28328
rect 1516 28204 1556 28244
rect 1420 27868 1460 27908
rect 1612 27784 1652 27824
rect 1708 27616 1748 27656
rect 1420 27532 1460 27572
rect 1324 26860 1364 26900
rect 1036 26272 1076 26312
rect 1036 25600 1076 25640
rect 940 21568 980 21608
rect 1324 23752 1364 23792
rect 1132 22912 1172 22952
rect 1228 21568 1268 21608
rect 1228 20980 1268 21020
rect 1132 20812 1172 20852
rect 1228 20728 1268 20768
rect 1132 20140 1172 20180
rect 1228 19636 1268 19676
rect 1132 19552 1172 19592
rect 1036 18880 1076 18920
rect 1324 18208 1364 18248
rect 1324 17032 1364 17072
rect 2380 32152 2420 32192
rect 2668 33160 2708 33200
rect 3244 37780 3284 37820
rect 3436 37780 3476 37820
rect 3052 36688 3092 36728
rect 2956 35176 2996 35216
rect 3148 35680 3188 35720
rect 3148 35260 3188 35300
rect 3340 37360 3380 37400
rect 3628 37948 3668 37988
rect 3820 37948 3860 37988
rect 3688 37780 3728 37820
rect 3770 37780 3810 37820
rect 3852 37780 3892 37820
rect 3934 37780 3974 37820
rect 4016 37780 4056 37820
rect 3532 37696 3572 37736
rect 3820 37612 3860 37652
rect 4876 42064 4916 42104
rect 5356 41980 5396 42020
rect 5260 41728 5300 41768
rect 4684 41644 4724 41684
rect 4588 41560 4628 41600
rect 4492 41476 4532 41516
rect 4928 41560 4968 41600
rect 5010 41560 5050 41600
rect 5092 41560 5132 41600
rect 5174 41560 5214 41600
rect 5256 41560 5296 41600
rect 4780 41308 4820 41348
rect 4492 40384 4532 40424
rect 5356 40972 5396 41012
rect 5644 42400 5684 42440
rect 6028 42148 6068 42188
rect 5548 41140 5588 41180
rect 4396 38872 4436 38912
rect 5260 40300 5300 40340
rect 5068 40216 5108 40256
rect 4928 40048 4968 40088
rect 5010 40048 5050 40088
rect 5092 40048 5132 40088
rect 5174 40048 5214 40088
rect 5256 40048 5296 40088
rect 4588 39544 4628 39584
rect 5260 39544 5300 39584
rect 6508 41560 6548 41600
rect 6124 41476 6164 41516
rect 5836 41140 5876 41180
rect 5452 40636 5492 40676
rect 5452 39460 5492 39500
rect 5644 40300 5684 40340
rect 5644 39544 5684 39584
rect 5644 39376 5684 39416
rect 4972 38956 5012 38996
rect 4588 38788 4628 38828
rect 4396 38200 4436 38240
rect 4300 38032 4340 38072
rect 4492 38032 4532 38072
rect 4108 37108 4148 37148
rect 3688 36268 3728 36308
rect 3770 36268 3810 36308
rect 3852 36268 3892 36308
rect 3934 36268 3974 36308
rect 4016 36268 4056 36308
rect 4012 35680 4052 35720
rect 3052 35008 3092 35048
rect 2860 34504 2900 34544
rect 2764 32824 2804 32864
rect 2380 31480 2420 31520
rect 2668 31312 2708 31352
rect 2476 31228 2516 31268
rect 2284 30220 2324 30260
rect 1996 28372 2036 28412
rect 1900 28288 1940 28328
rect 1900 28036 1940 28076
rect 1516 26104 1556 26144
rect 1516 25768 1556 25808
rect 1996 27784 2036 27824
rect 1708 23500 1748 23540
rect 1612 20728 1652 20768
rect 1516 16192 1556 16232
rect 2188 28540 2228 28580
rect 2188 28036 2228 28076
rect 2668 30976 2708 31016
rect 2572 30052 2612 30092
rect 2476 28540 2516 28580
rect 2380 28204 2420 28244
rect 2092 25600 2132 25640
rect 2572 27700 2612 27740
rect 2956 34084 2996 34124
rect 3436 35260 3476 35300
rect 3628 35260 3668 35300
rect 4012 35260 4052 35300
rect 3532 35092 3572 35132
rect 3436 34924 3476 34964
rect 3340 34756 3380 34796
rect 3244 34504 3284 34544
rect 3340 33664 3380 33704
rect 3148 32908 3188 32948
rect 3148 32656 3188 32696
rect 3052 32572 3092 32612
rect 2956 31312 2996 31352
rect 2860 30556 2900 30596
rect 2764 30220 2804 30260
rect 2764 29632 2804 29672
rect 2956 29632 2996 29672
rect 2860 29464 2900 29504
rect 2668 27112 2708 27152
rect 2572 26440 2612 26480
rect 2476 26104 2516 26144
rect 2380 25936 2420 25976
rect 2380 25432 2420 25472
rect 2284 25264 2324 25304
rect 3148 30136 3188 30176
rect 3820 35008 3860 35048
rect 3688 34756 3728 34796
rect 3770 34756 3810 34796
rect 3852 34756 3892 34796
rect 3934 34756 3974 34796
rect 4016 34756 4056 34796
rect 4396 37528 4436 37568
rect 4300 37108 4340 37148
rect 4204 37024 4244 37064
rect 5548 38788 5588 38828
rect 6028 39964 6068 40004
rect 5932 39796 5972 39836
rect 5932 39628 5972 39668
rect 6028 39292 6068 39332
rect 6508 41308 6548 41348
rect 6988 41896 7028 41936
rect 7084 41644 7124 41684
rect 6988 40972 7028 41012
rect 6508 40636 6548 40676
rect 6316 39880 6356 39920
rect 6412 39628 6452 39668
rect 6316 39040 6356 39080
rect 6988 40552 7028 40592
rect 6796 39628 6836 39668
rect 6892 39544 6932 39584
rect 5644 38704 5684 38744
rect 4928 38536 4968 38576
rect 5010 38536 5050 38576
rect 5092 38536 5132 38576
rect 5174 38536 5214 38576
rect 5256 38536 5296 38576
rect 5644 38536 5684 38576
rect 5644 38116 5684 38156
rect 6412 38956 6452 38996
rect 6796 38872 6836 38912
rect 6604 38704 6644 38744
rect 6796 38704 6836 38744
rect 6028 38032 6068 38072
rect 6508 37864 6548 37904
rect 4780 37444 4820 37484
rect 4684 37192 4724 37232
rect 4588 37108 4628 37148
rect 5932 37780 5972 37820
rect 5548 37360 5588 37400
rect 5164 37192 5204 37232
rect 5644 37108 5684 37148
rect 4928 37024 4968 37064
rect 5010 37024 5050 37064
rect 5092 37024 5132 37064
rect 5174 37024 5214 37064
rect 5256 37024 5296 37064
rect 5548 37024 5588 37064
rect 4204 36520 4244 36560
rect 4300 36016 4340 36056
rect 4492 35680 4532 35720
rect 4492 35512 4532 35552
rect 4396 35260 4436 35300
rect 4108 33832 4148 33872
rect 4012 33664 4052 33704
rect 4300 33748 4340 33788
rect 3820 33496 3860 33536
rect 3688 33244 3728 33284
rect 3770 33244 3810 33284
rect 3852 33244 3892 33284
rect 3934 33244 3974 33284
rect 4016 33244 4056 33284
rect 4492 34336 4532 34376
rect 3532 32656 3572 32696
rect 3340 32404 3380 32444
rect 3724 32824 3764 32864
rect 4108 32824 4148 32864
rect 4204 32152 4244 32192
rect 3340 31900 3380 31940
rect 3628 31900 3668 31940
rect 3688 31732 3728 31772
rect 3770 31732 3810 31772
rect 3852 31732 3892 31772
rect 3934 31732 3974 31772
rect 4016 31732 4056 31772
rect 4396 32740 4436 32780
rect 3340 31060 3380 31100
rect 3244 29968 3284 30008
rect 3340 29380 3380 29420
rect 3052 29296 3092 29336
rect 3148 28540 3188 28580
rect 3916 31228 3956 31268
rect 5452 36268 5492 36308
rect 4972 36100 5012 36140
rect 4876 35848 4916 35888
rect 5548 35680 5588 35720
rect 4928 35512 4968 35552
rect 5010 35512 5050 35552
rect 5092 35512 5132 35552
rect 5174 35512 5214 35552
rect 5256 35512 5296 35552
rect 4684 35260 4724 35300
rect 4108 31144 4148 31184
rect 3688 30220 3728 30260
rect 3770 30220 3810 30260
rect 3852 30220 3892 30260
rect 3934 30220 3974 30260
rect 4016 30220 4056 30260
rect 3532 30136 3572 30176
rect 3916 29128 3956 29168
rect 3436 29044 3476 29084
rect 6124 37528 6164 37568
rect 5932 37024 5972 37064
rect 6700 38620 6740 38660
rect 6796 38368 6836 38408
rect 6700 38284 6740 38324
rect 6796 37276 6836 37316
rect 6508 36856 6548 36896
rect 6508 36688 6548 36728
rect 6604 35932 6644 35972
rect 5356 35092 5396 35132
rect 5356 34168 5396 34208
rect 4928 34000 4968 34040
rect 5010 34000 5050 34040
rect 5092 34000 5132 34040
rect 5174 34000 5214 34040
rect 5256 34000 5296 34040
rect 4928 32488 4968 32528
rect 5010 32488 5050 32528
rect 5092 32488 5132 32528
rect 5174 32488 5214 32528
rect 5256 32488 5296 32528
rect 5740 34168 5780 34208
rect 6124 35176 6164 35216
rect 6028 35092 6068 35132
rect 6028 34756 6068 34796
rect 6124 34504 6164 34544
rect 6220 34336 6260 34376
rect 6412 35260 6452 35300
rect 6796 36856 6836 36896
rect 6988 38956 7028 38996
rect 7756 41728 7796 41768
rect 7564 41644 7604 41684
rect 7372 41560 7412 41600
rect 7756 41224 7796 41264
rect 8140 41560 8180 41600
rect 8140 41308 8180 41348
rect 8044 41224 8084 41264
rect 7948 41140 7988 41180
rect 7372 40888 7412 40928
rect 7180 40636 7220 40676
rect 7276 40048 7316 40088
rect 7276 39796 7316 39836
rect 7180 38704 7220 38744
rect 6892 36604 6932 36644
rect 6796 36184 6836 36224
rect 6796 35848 6836 35888
rect 6700 35428 6740 35468
rect 6508 35008 6548 35048
rect 6508 34252 6548 34292
rect 5740 33832 5780 33872
rect 5932 33832 5972 33872
rect 5836 33664 5876 33704
rect 5836 33076 5876 33116
rect 5740 32908 5780 32948
rect 5452 32404 5492 32444
rect 5932 32572 5972 32612
rect 6220 33076 6260 33116
rect 6124 32824 6164 32864
rect 6609 32908 6649 32948
rect 6508 32824 6548 32864
rect 4780 31144 4820 31184
rect 4928 30976 4968 31016
rect 5010 30976 5050 31016
rect 5092 30976 5132 31016
rect 5174 30976 5214 31016
rect 5256 30976 5296 31016
rect 5356 30724 5396 30764
rect 4876 30640 4916 30680
rect 5260 30556 5300 30596
rect 4588 29800 4628 29840
rect 4588 29380 4628 29420
rect 3532 28876 3572 28916
rect 3688 28708 3728 28748
rect 3770 28708 3810 28748
rect 3852 28708 3892 28748
rect 3934 28708 3974 28748
rect 4016 28708 4056 28748
rect 3916 28372 3956 28412
rect 3532 28288 3572 28328
rect 3436 27952 3476 27992
rect 3340 27868 3380 27908
rect 3052 27112 3092 27152
rect 2860 26440 2900 26480
rect 2764 26104 2804 26144
rect 2764 25852 2804 25892
rect 2860 25516 2900 25556
rect 2668 25264 2708 25304
rect 2956 25348 2996 25388
rect 3628 27784 3668 27824
rect 3532 27700 3572 27740
rect 3436 26860 3476 26900
rect 3148 26776 3188 26816
rect 3340 26104 3380 26144
rect 3436 25684 3476 25724
rect 3340 25516 3380 25556
rect 2860 25264 2900 25304
rect 3052 25264 3092 25304
rect 3436 25264 3476 25304
rect 2764 25180 2804 25220
rect 3688 27196 3728 27236
rect 3770 27196 3810 27236
rect 3852 27196 3892 27236
rect 3934 27196 3974 27236
rect 4016 27196 4056 27236
rect 3628 26860 3668 26900
rect 3916 26776 3956 26816
rect 3820 26608 3860 26648
rect 4108 26692 4148 26732
rect 5644 31900 5684 31940
rect 5836 31732 5876 31772
rect 5548 31228 5588 31268
rect 5740 31144 5780 31184
rect 5548 30808 5588 30848
rect 5260 30052 5300 30092
rect 4780 29800 4820 29840
rect 4928 29464 4968 29504
rect 5010 29464 5050 29504
rect 5092 29464 5132 29504
rect 5174 29464 5214 29504
rect 5256 29464 5296 29504
rect 5164 29296 5204 29336
rect 4780 29128 4820 29168
rect 6028 31900 6068 31940
rect 6124 30640 6164 30680
rect 6316 32068 6356 32108
rect 6508 31984 6548 32024
rect 6604 31732 6644 31772
rect 6412 31228 6452 31268
rect 6316 31144 6356 31184
rect 6508 31144 6548 31184
rect 6700 31144 6740 31184
rect 6700 30976 6740 31016
rect 6604 30724 6644 30764
rect 5548 29800 5588 29840
rect 5932 29800 5972 29840
rect 5452 29296 5492 29336
rect 5356 29212 5396 29252
rect 6028 29716 6068 29756
rect 5644 29632 5684 29672
rect 4684 28456 4724 28496
rect 4588 28288 4628 28328
rect 4492 28120 4532 28160
rect 4396 27868 4436 27908
rect 4588 27784 4628 27824
rect 4396 27532 4436 27572
rect 4588 27532 4628 27572
rect 3724 26020 3764 26060
rect 3820 25852 3860 25892
rect 3688 25684 3728 25724
rect 3770 25684 3810 25724
rect 3852 25684 3892 25724
rect 3934 25684 3974 25724
rect 4016 25684 4056 25724
rect 4396 25600 4436 25640
rect 4300 25432 4340 25472
rect 3820 25348 3860 25388
rect 4396 25264 4436 25304
rect 4012 25180 4052 25220
rect 3532 24760 3572 24800
rect 2668 23584 2708 23624
rect 2476 23080 2516 23120
rect 2572 23080 2612 23120
rect 2764 22912 2804 22952
rect 2572 22240 2612 22280
rect 3148 22912 3188 22952
rect 3052 22660 3092 22700
rect 2860 22576 2900 22616
rect 4588 24592 4628 24632
rect 5836 29128 5876 29168
rect 6028 29128 6068 29168
rect 5740 29044 5780 29084
rect 5164 28204 5204 28244
rect 4780 28036 4820 28076
rect 4928 27952 4968 27992
rect 5010 27952 5050 27992
rect 5092 27952 5132 27992
rect 5174 27952 5214 27992
rect 5256 27952 5296 27992
rect 4780 27616 4820 27656
rect 5644 28876 5684 28916
rect 5836 28960 5876 29000
rect 6220 30052 6260 30092
rect 6604 29716 6644 29756
rect 6316 29632 6356 29672
rect 6220 29212 6260 29252
rect 6412 29128 6452 29168
rect 6700 29464 6740 29504
rect 6604 29044 6644 29084
rect 5740 28456 5780 28496
rect 5740 28288 5780 28328
rect 5644 28204 5684 28244
rect 5932 28456 5972 28496
rect 5452 27448 5492 27488
rect 5356 27112 5396 27152
rect 5356 26608 5396 26648
rect 4928 26440 4968 26480
rect 5010 26440 5050 26480
rect 5092 26440 5132 26480
rect 5174 26440 5214 26480
rect 5256 26440 5296 26480
rect 4780 26356 4820 26396
rect 4972 26272 5012 26312
rect 5164 25936 5204 25976
rect 5740 27112 5780 27152
rect 5644 26776 5684 26816
rect 5548 26356 5588 26396
rect 6124 27616 6164 27656
rect 5932 26860 5972 26900
rect 5836 26776 5876 26816
rect 6220 26776 6260 26816
rect 6220 26608 6260 26648
rect 5356 25684 5396 25724
rect 4928 24928 4968 24968
rect 5010 24928 5050 24968
rect 5092 24928 5132 24968
rect 5174 24928 5214 24968
rect 5256 24928 5296 24968
rect 4780 24592 4820 24632
rect 3688 24172 3728 24212
rect 3770 24172 3810 24212
rect 3852 24172 3892 24212
rect 3934 24172 3974 24212
rect 4016 24172 4056 24212
rect 3532 23920 3572 23960
rect 4012 23920 4052 23960
rect 3532 23752 3572 23792
rect 3436 23584 3476 23624
rect 5260 23920 5300 23960
rect 4972 23752 5012 23792
rect 5260 23752 5300 23792
rect 4684 23584 4724 23624
rect 4300 23080 4340 23120
rect 4928 23416 4968 23456
rect 5010 23416 5050 23456
rect 5092 23416 5132 23456
rect 5174 23416 5214 23456
rect 5256 23416 5296 23456
rect 4972 23080 5012 23120
rect 4108 22996 4148 23036
rect 3244 21834 3284 21860
rect 3244 21820 3284 21834
rect 3688 22660 3728 22700
rect 3770 22660 3810 22700
rect 3852 22660 3892 22700
rect 3934 22660 3974 22700
rect 4016 22660 4056 22700
rect 3628 22156 3668 22196
rect 4012 22240 4052 22280
rect 4204 22660 4244 22700
rect 3724 21904 3764 21944
rect 2668 21568 2708 21608
rect 2956 21568 2996 21608
rect 3148 21568 3188 21608
rect 2572 21484 2612 21524
rect 2764 21400 2804 21440
rect 2764 20896 2804 20936
rect 3052 20896 3092 20936
rect 2956 20812 2996 20852
rect 2284 20224 2324 20264
rect 1804 19216 1844 19256
rect 1708 18964 1748 19004
rect 1708 17704 1748 17744
rect 1804 17536 1844 17576
rect 1900 15856 1940 15896
rect 1612 15604 1652 15644
rect 1324 14176 1364 14216
rect 1516 15520 1556 15560
rect 2188 19048 2228 19088
rect 2188 18796 2228 18836
rect 2284 18628 2324 18668
rect 2668 20728 2708 20768
rect 2668 20224 2708 20264
rect 3052 20728 3092 20768
rect 3340 21484 3380 21524
rect 3244 20896 3284 20936
rect 3724 21400 3764 21440
rect 3532 21316 3572 21356
rect 4204 21400 4244 21440
rect 3916 21316 3956 21356
rect 4204 21232 4244 21272
rect 3688 21148 3728 21188
rect 3770 21148 3810 21188
rect 3852 21148 3892 21188
rect 3934 21148 3974 21188
rect 4016 21148 4056 21188
rect 3532 20812 3572 20852
rect 3628 20728 3668 20768
rect 4492 22408 4532 22448
rect 5068 22324 5108 22364
rect 4492 22072 4532 22112
rect 4684 22240 4724 22280
rect 4928 21904 4968 21944
rect 5010 21904 5050 21944
rect 5092 21904 5132 21944
rect 5174 21904 5214 21944
rect 5256 21904 5296 21944
rect 4588 21568 4628 21608
rect 5068 21568 5108 21608
rect 3820 20728 3860 20768
rect 3340 20560 3380 20600
rect 3916 20560 3956 20600
rect 2860 20056 2900 20096
rect 2476 19972 2516 20012
rect 2572 19216 2612 19256
rect 2764 19216 2804 19256
rect 2380 17956 2420 17996
rect 2764 18880 2804 18920
rect 2956 18796 2996 18836
rect 3148 19048 3188 19088
rect 3052 18628 3092 18668
rect 2956 18460 2996 18500
rect 2764 18376 2804 18416
rect 2380 17032 2420 17072
rect 2668 17704 2708 17744
rect 2572 17536 2612 17576
rect 2860 18292 2900 18332
rect 2092 15772 2132 15812
rect 2668 15940 2708 15980
rect 3244 18376 3284 18416
rect 4204 20728 4244 20768
rect 4684 20896 4724 20936
rect 5068 20812 5108 20852
rect 4108 20224 4148 20264
rect 3916 20140 3956 20180
rect 4204 20056 4244 20096
rect 4012 19972 4052 20012
rect 4108 19804 4148 19844
rect 3688 19636 3728 19676
rect 3770 19636 3810 19676
rect 3852 19636 3892 19676
rect 3934 19636 3974 19676
rect 4016 19636 4056 19676
rect 3532 19216 3572 19256
rect 4396 20140 4436 20180
rect 4300 19972 4340 20012
rect 4396 19552 4436 19592
rect 4684 19972 4724 20012
rect 4396 19300 4436 19340
rect 4300 18712 4340 18752
rect 3436 18628 3476 18668
rect 4108 18544 4148 18584
rect 3820 18376 3860 18416
rect 3628 18292 3668 18332
rect 3688 18124 3728 18164
rect 3770 18124 3810 18164
rect 3852 18124 3892 18164
rect 3934 18124 3974 18164
rect 4016 18124 4056 18164
rect 3820 17956 3860 17996
rect 3340 17788 3380 17828
rect 3628 17788 3668 17828
rect 3532 17704 3572 17744
rect 4204 18292 4244 18332
rect 4588 19216 4628 19256
rect 4588 18712 4628 18752
rect 4928 20392 4968 20432
rect 5010 20392 5050 20432
rect 5092 20392 5132 20432
rect 5174 20392 5214 20432
rect 5256 20392 5296 20432
rect 6028 26440 6068 26480
rect 6028 26272 6068 26312
rect 6124 26188 6164 26228
rect 5836 24928 5876 24968
rect 5836 24172 5876 24212
rect 5452 23920 5492 23960
rect 5644 23752 5684 23792
rect 5548 23668 5588 23708
rect 5644 23416 5684 23456
rect 5548 23332 5588 23372
rect 5548 22828 5588 22868
rect 5548 21484 5588 21524
rect 5836 23416 5876 23456
rect 5836 22996 5876 23036
rect 5740 22576 5780 22616
rect 5740 20980 5780 21020
rect 5644 20896 5684 20936
rect 5740 20812 5780 20852
rect 5644 20728 5684 20768
rect 6028 24928 6068 24968
rect 6124 24592 6164 24632
rect 6028 24424 6068 24464
rect 6220 24424 6260 24464
rect 6124 23500 6164 23540
rect 5932 22576 5972 22616
rect 6028 21736 6068 21776
rect 5932 21568 5972 21608
rect 6124 21400 6164 21440
rect 4780 19804 4820 19844
rect 4876 19720 4916 19760
rect 4780 19300 4820 19340
rect 5260 20056 5300 20096
rect 4972 19552 5012 19592
rect 4876 19216 4916 19256
rect 4928 18880 4968 18920
rect 5010 18880 5050 18920
rect 5092 18880 5132 18920
rect 5174 18880 5214 18920
rect 5256 18880 5296 18920
rect 4876 18712 4916 18752
rect 5356 18712 5396 18752
rect 5068 18544 5108 18584
rect 4588 18292 4628 18332
rect 4204 18124 4244 18164
rect 4492 18124 4532 18164
rect 4780 18124 4820 18164
rect 4108 17788 4148 17828
rect 3244 17620 3284 17660
rect 3436 17620 3476 17660
rect 2956 16612 2996 16652
rect 3340 16612 3380 16652
rect 3148 16444 3188 16484
rect 2956 16360 2996 16400
rect 3244 16360 3284 16400
rect 3688 16612 3728 16652
rect 3770 16612 3810 16652
rect 3852 16612 3892 16652
rect 3934 16612 3974 16652
rect 4016 16612 4056 16652
rect 3724 16444 3764 16484
rect 3148 15940 3188 15980
rect 2860 15604 2900 15644
rect 2380 15436 2420 15476
rect 2284 14848 2324 14888
rect 1516 14512 1556 14552
rect 1516 13252 1556 13292
rect 1516 12832 1556 12872
rect 2092 14764 2132 14804
rect 1996 14428 2036 14468
rect 1708 14008 1748 14048
rect 1900 13840 1940 13880
rect 1804 13504 1844 13544
rect 1708 12580 1748 12620
rect 1612 12328 1652 12368
rect 1708 12244 1748 12284
rect 1516 12160 1556 12200
rect 3340 15604 3380 15644
rect 3820 15940 3860 15980
rect 2668 14092 2708 14132
rect 2092 13924 2132 13964
rect 1900 13084 1940 13124
rect 2092 13084 2132 13124
rect 1996 12916 2036 12956
rect 1708 11740 1748 11780
rect 1804 11488 1844 11528
rect 1516 11320 1556 11360
rect 1324 10816 1364 10856
rect 556 9220 596 9260
rect 556 8464 596 8504
rect 1420 10312 1460 10352
rect 1420 10144 1460 10184
rect 1708 11236 1748 11276
rect 1612 9976 1652 10016
rect 1516 8800 1556 8840
rect 1900 10060 1940 10100
rect 2572 13924 2612 13964
rect 2476 12664 2516 12704
rect 2956 12580 2996 12620
rect 2476 12496 2516 12536
rect 2092 12412 2132 12452
rect 2476 11320 2516 11360
rect 2188 11152 2228 11192
rect 2092 9724 2132 9764
rect 1996 8884 2036 8924
rect 1996 8716 2036 8756
rect 1804 8632 1844 8672
rect 1612 7876 1652 7916
rect 1324 7792 1364 7832
rect 1612 7204 1652 7244
rect 1804 8128 1844 8168
rect 2092 8548 2132 8588
rect 2476 10984 2516 11024
rect 2860 10480 2900 10520
rect 2764 10396 2804 10436
rect 3244 14680 3284 14720
rect 3340 13924 3380 13964
rect 3148 13168 3188 13208
rect 3688 15100 3728 15140
rect 3770 15100 3810 15140
rect 3852 15100 3892 15140
rect 3934 15100 3974 15140
rect 4016 15100 4056 15140
rect 4396 18040 4436 18080
rect 4492 17788 4532 17828
rect 4396 17704 4436 17744
rect 5356 18040 5396 18080
rect 5068 17704 5108 17744
rect 5260 17620 5300 17660
rect 4928 17368 4968 17408
rect 5010 17368 5050 17408
rect 5092 17368 5132 17408
rect 5174 17368 5214 17408
rect 5256 17368 5296 17408
rect 4300 16192 4340 16232
rect 4108 14848 4148 14888
rect 3724 14596 3764 14636
rect 4396 14764 4436 14804
rect 4300 14092 4340 14132
rect 3916 13924 3956 13964
rect 3688 13588 3728 13628
rect 3770 13588 3810 13628
rect 3852 13588 3892 13628
rect 3934 13588 3974 13628
rect 4016 13588 4056 13628
rect 3532 13252 3572 13292
rect 4108 12580 4148 12620
rect 3916 12496 3956 12536
rect 3688 12076 3728 12116
rect 3770 12076 3810 12116
rect 3852 12076 3892 12116
rect 3934 12076 3974 12116
rect 4016 12076 4056 12116
rect 3532 11656 3572 11696
rect 3148 11404 3188 11444
rect 2380 10144 2420 10184
rect 2284 9472 2324 9512
rect 2188 7708 2228 7748
rect 1804 7456 1844 7496
rect 1516 6784 1556 6824
rect 1420 5692 1460 5732
rect 1324 5608 1364 5648
rect 1324 4936 1364 4976
rect 1324 4600 1364 4640
rect 364 3844 404 3884
rect 1516 3928 1556 3968
rect 1996 7372 2036 7412
rect 2572 10060 2612 10100
rect 2476 9892 2516 9932
rect 2476 7540 2516 7580
rect 2188 6952 2228 6992
rect 1996 6868 2036 6908
rect 1804 6532 1844 6572
rect 1708 6364 1748 6404
rect 1708 5440 1748 5480
rect 1516 3172 1556 3212
rect 2092 6616 2132 6656
rect 2284 6364 2324 6404
rect 2188 5860 2228 5900
rect 1996 5356 2036 5396
rect 1900 4096 1940 4136
rect 1900 2752 1940 2792
rect 2092 4936 2132 4976
rect 2476 6280 2516 6320
rect 2284 5104 2324 5144
rect 2476 5020 2516 5060
rect 2476 4096 2516 4136
rect 2188 3760 2228 3800
rect 2476 3592 2516 3632
rect 2284 3424 2324 3464
rect 2380 3088 2420 3128
rect 2476 2668 2516 2708
rect 1996 2500 2036 2540
rect 2380 2500 2420 2540
rect 2668 9136 2708 9176
rect 2860 10060 2900 10100
rect 3532 10984 3572 11024
rect 3916 11572 3956 11612
rect 3724 10732 3764 10772
rect 4204 10732 4244 10772
rect 3688 10564 3728 10604
rect 3770 10564 3810 10604
rect 3852 10564 3892 10604
rect 3934 10564 3974 10604
rect 4016 10564 4056 10604
rect 3916 10396 3956 10436
rect 4204 10396 4244 10436
rect 3532 10312 3572 10352
rect 2860 9556 2900 9596
rect 3052 9472 3092 9512
rect 2764 8548 2804 8588
rect 3148 9304 3188 9344
rect 3052 7792 3092 7832
rect 2764 7540 2804 7580
rect 2860 6952 2900 6992
rect 2668 6532 2708 6572
rect 2764 6448 2804 6488
rect 2956 6700 2996 6740
rect 3052 4936 3092 4976
rect 3052 4768 3092 4808
rect 3052 4264 3092 4304
rect 3436 9472 3476 9512
rect 3820 10228 3860 10268
rect 3724 10060 3764 10100
rect 3724 9472 3764 9512
rect 4396 13168 4436 13208
rect 4492 12496 4532 12536
rect 4396 11488 4436 11528
rect 4492 10648 4532 10688
rect 6028 20812 6068 20852
rect 6508 28960 6548 29000
rect 6604 28876 6644 28916
rect 6700 27280 6740 27320
rect 6604 27112 6644 27152
rect 6988 35008 7028 35048
rect 6988 33076 7028 33116
rect 7180 36688 7220 36728
rect 7660 40384 7700 40424
rect 7468 40300 7508 40340
rect 7468 40048 7508 40088
rect 7468 38872 7508 38912
rect 7564 38200 7604 38240
rect 7468 38116 7508 38156
rect 7468 37192 7508 37232
rect 7372 36856 7412 36896
rect 7468 36520 7508 36560
rect 7660 37780 7700 37820
rect 8524 41476 8564 41516
rect 8332 41056 8372 41096
rect 8044 40804 8084 40844
rect 7948 40636 7988 40676
rect 8140 40468 8180 40508
rect 7852 40300 7892 40340
rect 8236 39964 8276 40004
rect 8044 39712 8084 39752
rect 8524 40132 8564 40172
rect 8524 39376 8564 39416
rect 8428 38872 8468 38912
rect 8332 38788 8372 38828
rect 8044 38368 8084 38408
rect 7756 37612 7796 37652
rect 8044 37696 8084 37736
rect 8524 38368 8564 38408
rect 8428 37780 8468 37820
rect 8044 37444 8084 37484
rect 8332 37444 8372 37484
rect 7852 37360 7892 37400
rect 7660 36688 7700 36728
rect 7564 36352 7604 36392
rect 7180 34588 7220 34628
rect 7180 34000 7220 34040
rect 7084 31732 7124 31772
rect 7084 29380 7124 29420
rect 7468 35260 7508 35300
rect 7948 36940 7988 36980
rect 8428 37360 8468 37400
rect 8620 38200 8660 38240
rect 8620 36856 8660 36896
rect 7756 35932 7796 35972
rect 7660 35176 7700 35216
rect 7756 35092 7796 35132
rect 7660 34924 7700 34964
rect 7660 34672 7700 34712
rect 7756 34588 7796 34628
rect 7564 34420 7604 34460
rect 8044 35680 8084 35720
rect 8428 35344 8468 35384
rect 8044 35260 8084 35300
rect 7948 35176 7988 35216
rect 8044 35008 8084 35048
rect 7948 34252 7988 34292
rect 8908 42148 8948 42188
rect 9004 40468 9044 40508
rect 8908 40384 8948 40424
rect 8908 40216 8948 40256
rect 8812 38956 8852 38996
rect 8812 38620 8852 38660
rect 9292 42232 9332 42272
rect 9292 42064 9332 42104
rect 9196 41980 9236 42020
rect 9580 42568 9620 42608
rect 9484 41560 9524 41600
rect 9388 41392 9428 41432
rect 9388 41224 9428 41264
rect 9292 41140 9332 41180
rect 9580 41140 9620 41180
rect 9196 39964 9236 40004
rect 9100 38116 9140 38156
rect 9484 39964 9524 40004
rect 9004 37444 9044 37484
rect 8524 34924 8564 34964
rect 8140 34588 8180 34628
rect 8332 34336 8372 34376
rect 8140 34084 8180 34124
rect 7852 33916 7892 33956
rect 7564 33664 7604 33704
rect 7852 33664 7892 33704
rect 7372 33412 7412 33452
rect 7372 33076 7412 33116
rect 7372 30976 7412 31016
rect 7660 33580 7700 33620
rect 8236 33664 8276 33704
rect 8044 33496 8084 33536
rect 7948 33412 7988 33452
rect 8140 33244 8180 33284
rect 7948 32908 7988 32948
rect 7564 32824 7604 32864
rect 7564 32404 7604 32444
rect 7564 31480 7604 31520
rect 9100 37192 9140 37232
rect 8908 36688 8948 36728
rect 8812 35344 8852 35384
rect 8812 35176 8852 35216
rect 8716 34924 8756 34964
rect 9004 36436 9044 36476
rect 9964 41896 10004 41936
rect 10156 41140 10196 41180
rect 9868 40216 9908 40256
rect 9772 39880 9812 39920
rect 10060 40384 10100 40424
rect 10348 41812 10388 41852
rect 10444 41560 10484 41600
rect 10348 40552 10388 40592
rect 9868 38872 9908 38912
rect 9868 38536 9908 38576
rect 10060 38536 10100 38576
rect 10252 40048 10292 40088
rect 10252 38788 10292 38828
rect 9196 36184 9236 36224
rect 9004 35680 9044 35720
rect 9100 35092 9140 35132
rect 8620 34336 8660 34376
rect 8524 34168 8564 34208
rect 8524 33412 8564 33452
rect 8332 33244 8372 33284
rect 9484 36856 9524 36896
rect 9484 36604 9524 36644
rect 9388 36436 9428 36476
rect 10156 36688 10196 36728
rect 10060 36184 10100 36224
rect 9388 36016 9428 36056
rect 9292 35764 9332 35804
rect 9292 35596 9332 35636
rect 9580 35848 9620 35888
rect 10156 35764 10196 35804
rect 10732 40468 10772 40508
rect 10444 39040 10484 39080
rect 10636 39040 10676 39080
rect 10636 38872 10676 38912
rect 10540 38788 10580 38828
rect 10636 38368 10676 38408
rect 10924 40384 10964 40424
rect 10732 38200 10772 38240
rect 10540 37948 10580 37988
rect 10348 36604 10388 36644
rect 10348 36184 10388 36224
rect 10252 35680 10292 35720
rect 10060 35596 10100 35636
rect 9580 35512 9620 35552
rect 10060 35344 10100 35384
rect 9868 35260 9908 35300
rect 9388 35008 9428 35048
rect 8908 34336 8948 34376
rect 9009 34336 9049 34376
rect 9196 34252 9236 34292
rect 10060 35176 10100 35216
rect 9964 34924 10004 34964
rect 9676 34756 9716 34796
rect 9580 34672 9620 34712
rect 9964 34672 10004 34712
rect 9772 34588 9812 34628
rect 9580 34336 9620 34376
rect 9100 34168 9140 34208
rect 9484 34168 9524 34208
rect 8812 33664 8852 33704
rect 8908 33580 8948 33620
rect 8236 32488 8276 32528
rect 7948 31564 7988 31604
rect 7756 31480 7796 31520
rect 8524 31480 8564 31520
rect 7756 31144 7796 31184
rect 7564 31060 7604 31100
rect 7468 30220 7508 30260
rect 7372 29716 7412 29756
rect 7468 29296 7508 29336
rect 7180 28876 7220 28916
rect 7180 28708 7220 28748
rect 7372 28708 7412 28748
rect 6988 28456 7028 28496
rect 7084 28204 7124 28244
rect 6988 27952 7028 27992
rect 6988 26944 7028 26984
rect 7468 28456 7508 28496
rect 7756 30892 7796 30932
rect 7660 29296 7700 29336
rect 7468 28036 7508 28076
rect 6412 26440 6452 26480
rect 6604 26776 6644 26816
rect 6700 26188 6740 26228
rect 6508 25936 6548 25976
rect 6892 26692 6932 26732
rect 6412 24844 6452 24884
rect 6508 24256 6548 24296
rect 6796 24424 6836 24464
rect 6700 24088 6740 24128
rect 6604 23920 6644 23960
rect 6412 23752 6452 23792
rect 7084 26776 7124 26816
rect 7180 26608 7220 26648
rect 7084 26440 7124 26480
rect 7372 26020 7412 26060
rect 7276 25348 7316 25388
rect 7180 25264 7220 25304
rect 6892 23836 6932 23876
rect 6508 23584 6548 23624
rect 6412 23332 6452 23372
rect 6988 23752 7028 23792
rect 6604 23500 6644 23540
rect 6988 23416 7028 23456
rect 6316 22660 6356 22700
rect 6508 22660 6548 22700
rect 6508 22408 6548 22448
rect 5548 20056 5588 20096
rect 5644 18964 5684 19004
rect 5644 18796 5684 18836
rect 5836 20224 5876 20264
rect 5932 20140 5972 20180
rect 5932 19804 5972 19844
rect 5836 19216 5876 19256
rect 5452 16696 5492 16736
rect 4972 16360 5012 16400
rect 6124 20392 6164 20432
rect 6028 16444 6068 16484
rect 5356 16360 5396 16400
rect 4928 15856 4968 15896
rect 5010 15856 5050 15896
rect 5092 15856 5132 15896
rect 5174 15856 5214 15896
rect 5256 15856 5296 15896
rect 5260 15688 5300 15728
rect 5068 15604 5108 15644
rect 5452 15856 5492 15896
rect 5548 15604 5588 15644
rect 5452 15520 5492 15560
rect 5068 14680 5108 14720
rect 5836 16024 5876 16064
rect 5740 15856 5780 15896
rect 5452 14680 5492 14720
rect 4928 14344 4968 14384
rect 5010 14344 5050 14384
rect 5092 14344 5132 14384
rect 5174 14344 5214 14384
rect 5256 14344 5296 14384
rect 6028 15856 6068 15896
rect 6508 21484 6548 21524
rect 6892 22996 6932 23036
rect 7180 23416 7220 23456
rect 7180 22996 7220 23036
rect 7084 22660 7124 22700
rect 6796 22408 6836 22448
rect 6988 22408 7028 22448
rect 7180 22156 7220 22196
rect 6700 21736 6740 21776
rect 7276 21736 7316 21776
rect 7468 25096 7508 25136
rect 7660 26104 7700 26144
rect 7660 25096 7700 25136
rect 7852 30220 7892 30260
rect 8428 31312 8468 31352
rect 8524 31060 8564 31100
rect 8812 32824 8852 32864
rect 9388 33916 9428 33956
rect 9868 34168 9908 34208
rect 9292 33412 9332 33452
rect 9196 33076 9236 33116
rect 9676 33496 9716 33536
rect 9580 33244 9620 33284
rect 9100 32992 9140 33032
rect 9484 32992 9524 33032
rect 9388 32908 9428 32948
rect 9484 32824 9524 32864
rect 9676 32824 9716 32864
rect 9964 33748 10004 33788
rect 9964 33412 10004 33452
rect 9388 32740 9428 32780
rect 8716 32572 8756 32612
rect 8716 32152 8756 32192
rect 8908 31480 8948 31520
rect 10252 35176 10292 35216
rect 10348 34924 10388 34964
rect 10252 34336 10292 34376
rect 10348 34168 10388 34208
rect 10252 34084 10292 34124
rect 10252 33748 10292 33788
rect 10252 33412 10292 33452
rect 10156 33244 10196 33284
rect 10444 33160 10484 33200
rect 11020 40300 11060 40340
rect 11116 39040 11156 39080
rect 11020 38872 11060 38912
rect 10924 37276 10964 37316
rect 11404 42064 11444 42104
rect 11308 41644 11348 41684
rect 11308 41308 11348 41348
rect 10732 36688 10772 36728
rect 10636 36268 10676 36308
rect 10924 36100 10964 36140
rect 11116 36520 11156 36560
rect 11884 42064 11924 42104
rect 11788 41476 11828 41516
rect 11596 41140 11636 41180
rect 12076 40888 12116 40928
rect 11692 40384 11732 40424
rect 11788 40300 11828 40340
rect 11500 40132 11540 40172
rect 11788 39964 11828 40004
rect 11692 39712 11732 39752
rect 11980 40300 12020 40340
rect 12364 42568 12404 42608
rect 12556 41560 12596 41600
rect 12268 40384 12308 40424
rect 12364 40300 12404 40340
rect 12172 40048 12212 40088
rect 11980 39712 12020 39752
rect 11980 39292 12020 39332
rect 11500 38536 11540 38576
rect 11884 38536 11924 38576
rect 11596 37696 11636 37736
rect 11404 36520 11444 36560
rect 11308 36100 11348 36140
rect 10732 35680 10772 35720
rect 10636 34000 10676 34040
rect 9676 32656 9716 32696
rect 9580 32320 9620 32360
rect 8812 31228 8852 31268
rect 8620 30892 8660 30932
rect 9100 30892 9140 30932
rect 8620 30724 8660 30764
rect 9004 30640 9044 30680
rect 9100 30472 9140 30512
rect 8524 30220 8564 30260
rect 8812 30220 8852 30260
rect 8812 29968 8852 30008
rect 9388 29968 9428 30008
rect 8716 29800 8756 29840
rect 9004 29800 9044 29840
rect 8812 29716 8852 29756
rect 8140 29296 8180 29336
rect 8236 28792 8276 28832
rect 7852 27952 7892 27992
rect 8044 27952 8084 27992
rect 8140 27532 8180 27572
rect 8620 29128 8660 29168
rect 8812 29296 8852 29336
rect 8908 29212 8948 29252
rect 8428 28960 8468 29000
rect 8716 28960 8756 29000
rect 8332 28204 8372 28244
rect 8332 26944 8372 26984
rect 8236 26860 8276 26900
rect 8044 25180 8084 25220
rect 7564 23920 7604 23960
rect 7948 24424 7988 24464
rect 8524 28288 8564 28328
rect 8908 28876 8948 28916
rect 8812 27700 8852 27740
rect 8812 27448 8852 27488
rect 8716 27364 8756 27404
rect 8524 26776 8564 26816
rect 8428 25768 8468 25808
rect 8332 24592 8372 24632
rect 8332 24340 8372 24380
rect 8140 23752 8180 23792
rect 8044 23668 8084 23708
rect 7564 23332 7604 23372
rect 8140 23248 8180 23288
rect 7756 23164 7796 23204
rect 7468 23080 7508 23120
rect 7564 22660 7604 22700
rect 7372 21652 7412 21692
rect 6604 21400 6644 21440
rect 7084 21568 7124 21608
rect 6412 21148 6452 21188
rect 6700 21148 6740 21188
rect 6892 21400 6932 21440
rect 6892 21148 6932 21188
rect 6700 20812 6740 20852
rect 6802 20812 6842 20852
rect 6220 19972 6260 20012
rect 6220 19804 6260 19844
rect 7276 21484 7316 21524
rect 7084 21316 7124 21356
rect 7372 21316 7412 21356
rect 7084 21148 7124 21188
rect 7084 20728 7124 20768
rect 6988 20644 7028 20684
rect 6796 20056 6836 20096
rect 6892 19972 6932 20012
rect 6796 19804 6836 19844
rect 6316 19636 6356 19676
rect 6316 19216 6356 19256
rect 6316 19048 6356 19088
rect 6508 19048 6548 19088
rect 6604 18880 6644 18920
rect 6508 18712 6548 18752
rect 6412 17620 6452 17660
rect 6220 17116 6260 17156
rect 6796 18292 6836 18332
rect 6700 17620 6740 17660
rect 6604 17452 6644 17492
rect 6220 16360 6260 16400
rect 6220 16024 6260 16064
rect 5932 15688 5972 15728
rect 5932 14680 5972 14720
rect 5836 14428 5876 14468
rect 5548 14008 5588 14048
rect 5260 13924 5300 13964
rect 5068 13756 5108 13796
rect 4204 10060 4244 10100
rect 3688 9052 3728 9092
rect 3770 9052 3810 9092
rect 3852 9052 3892 9092
rect 3934 9052 3974 9092
rect 4016 9052 4056 9092
rect 3244 8212 3284 8252
rect 4928 12832 4968 12872
rect 5010 12832 5050 12872
rect 5092 12832 5132 12872
rect 5174 12832 5214 12872
rect 5256 12832 5296 12872
rect 5644 13756 5684 13796
rect 5068 11824 5108 11864
rect 4928 11320 4968 11360
rect 5010 11320 5050 11360
rect 5092 11320 5132 11360
rect 5174 11320 5214 11360
rect 5256 11320 5296 11360
rect 5356 11068 5396 11108
rect 4684 10228 4724 10268
rect 4492 9472 4532 9512
rect 4300 9388 4340 9428
rect 4204 9136 4244 9176
rect 4300 8212 4340 8252
rect 4204 8128 4244 8168
rect 3436 7792 3476 7832
rect 3340 6952 3380 6992
rect 4108 7708 4148 7748
rect 3688 7540 3728 7580
rect 3770 7540 3810 7580
rect 3852 7540 3892 7580
rect 3934 7540 3974 7580
rect 4016 7540 4056 7580
rect 3532 7120 3572 7160
rect 3916 7120 3956 7160
rect 3820 6700 3860 6740
rect 3916 6532 3956 6572
rect 4012 6364 4052 6404
rect 3688 6028 3728 6068
rect 3770 6028 3810 6068
rect 3852 6028 3892 6068
rect 3934 6028 3974 6068
rect 4016 6028 4056 6068
rect 3148 4180 3188 4220
rect 2668 4012 2708 4052
rect 2860 3928 2900 3968
rect 2956 3760 2996 3800
rect 3148 2752 3188 2792
rect 1516 2416 1556 2456
rect 1804 2416 1844 2456
rect 1420 2332 1460 2372
rect 1516 1744 1556 1784
rect 1420 1576 1460 1616
rect 364 1072 404 1112
rect 1708 988 1748 1028
rect 1900 2080 1940 2120
rect 2092 2332 2132 2372
rect 2956 2332 2996 2372
rect 2572 2164 2612 2204
rect 2476 2080 2516 2120
rect 2284 1408 2324 1448
rect 2188 1324 2228 1364
rect 2380 652 2420 692
rect 3340 5020 3380 5060
rect 3340 3760 3380 3800
rect 3532 5020 3572 5060
rect 3916 5020 3956 5060
rect 4108 5020 4148 5060
rect 3628 4768 3668 4808
rect 3532 4684 3572 4724
rect 3688 4516 3728 4556
rect 3770 4516 3810 4556
rect 3852 4516 3892 4556
rect 3934 4516 3974 4556
rect 4016 4516 4056 4556
rect 4492 7456 4532 7496
rect 4492 7288 4532 7328
rect 4396 7204 4436 7244
rect 4300 6700 4340 6740
rect 4396 6448 4436 6488
rect 4300 6364 4340 6404
rect 5164 10228 5204 10268
rect 4684 9808 4724 9848
rect 4972 10060 5012 10100
rect 4928 9808 4968 9848
rect 5010 9808 5050 9848
rect 5092 9808 5132 9848
rect 5174 9808 5214 9848
rect 5256 9808 5296 9848
rect 5644 11068 5684 11108
rect 5932 14008 5972 14048
rect 5836 11068 5876 11108
rect 5548 10312 5588 10352
rect 4780 9472 4820 9512
rect 4684 8968 4724 9008
rect 4684 8800 4724 8840
rect 5452 9556 5492 9596
rect 5548 8800 5588 8840
rect 5740 8800 5780 8840
rect 4780 8548 4820 8588
rect 4928 8296 4968 8336
rect 5010 8296 5050 8336
rect 5092 8296 5132 8336
rect 5174 8296 5214 8336
rect 5256 8296 5296 8336
rect 5740 8128 5780 8168
rect 4780 7960 4820 8000
rect 5452 7792 5492 7832
rect 4684 7708 4724 7748
rect 4588 6532 4628 6572
rect 4780 7456 4820 7496
rect 4204 4768 4244 4808
rect 4204 4600 4244 4640
rect 4108 4348 4148 4388
rect 4492 6196 4532 6236
rect 4492 5608 4532 5648
rect 4972 7204 5012 7244
rect 4972 6952 5012 6992
rect 4928 6784 4968 6824
rect 5010 6784 5050 6824
rect 5092 6784 5132 6824
rect 5174 6784 5214 6824
rect 5256 6784 5296 6824
rect 4928 5272 4968 5312
rect 5010 5272 5050 5312
rect 5092 5272 5132 5312
rect 5174 5272 5214 5312
rect 5256 5272 5296 5312
rect 4396 4768 4436 4808
rect 4300 4516 4340 4556
rect 4300 4264 4340 4304
rect 4108 4180 4148 4220
rect 4108 3928 4148 3968
rect 4492 4684 4532 4724
rect 4492 4516 4532 4556
rect 4588 4012 4628 4052
rect 4396 3760 4436 3800
rect 4396 3424 4436 3464
rect 3688 3004 3728 3044
rect 3770 3004 3810 3044
rect 3852 3004 3892 3044
rect 3934 3004 3974 3044
rect 4016 3004 4056 3044
rect 4108 2836 4148 2876
rect 3628 2584 3668 2624
rect 3148 2332 3188 2372
rect 2668 1912 2708 1952
rect 2860 1660 2900 1700
rect 2764 1240 2804 1280
rect 2668 148 2708 188
rect 2956 1240 2996 1280
rect 3148 1240 3188 1280
rect 3436 2500 3476 2540
rect 3724 2500 3764 2540
rect 4204 2500 4244 2540
rect 3724 1744 3764 1784
rect 3688 1492 3728 1532
rect 3770 1492 3810 1532
rect 3852 1492 3892 1532
rect 3934 1492 3974 1532
rect 4016 1492 4056 1532
rect 3532 1240 3572 1280
rect 3340 736 3380 776
rect 3340 568 3380 608
rect 3916 1156 3956 1196
rect 3724 316 3764 356
rect 4108 820 4148 860
rect 4684 3928 4724 3968
rect 4492 2752 4532 2792
rect 4492 2584 4532 2624
rect 4396 1912 4436 1952
rect 4300 1408 4340 1448
rect 4300 1072 4340 1112
rect 5068 4180 5108 4220
rect 4876 3928 4916 3968
rect 4928 3760 4968 3800
rect 5010 3760 5050 3800
rect 5092 3760 5132 3800
rect 5174 3760 5214 3800
rect 5256 3760 5296 3800
rect 4780 2920 4820 2960
rect 4780 2668 4820 2708
rect 5164 2668 5204 2708
rect 4876 2500 4916 2540
rect 4928 2248 4968 2288
rect 5010 2248 5050 2288
rect 5092 2248 5132 2288
rect 5174 2248 5214 2288
rect 5256 2248 5296 2288
rect 4876 1996 4916 2036
rect 5644 6952 5684 6992
rect 5644 6700 5684 6740
rect 5548 5860 5588 5900
rect 5836 6700 5876 6740
rect 5932 6448 5972 6488
rect 6508 14764 6548 14804
rect 6412 14680 6452 14720
rect 6700 16444 6740 16484
rect 6700 15520 6740 15560
rect 7852 23080 7892 23120
rect 7852 22576 7892 22616
rect 8044 23080 8084 23120
rect 8140 22912 8180 22952
rect 8044 22660 8084 22700
rect 7948 22072 7988 22112
rect 7660 21484 7700 21524
rect 7660 21316 7700 21356
rect 7372 20056 7412 20096
rect 7852 21568 7892 21608
rect 7756 20056 7796 20096
rect 7660 19720 7700 19760
rect 8140 20644 8180 20684
rect 8428 23668 8468 23708
rect 9004 28372 9044 28412
rect 9484 29800 9524 29840
rect 9580 29716 9620 29756
rect 9196 29632 9236 29672
rect 9964 32404 10004 32444
rect 9772 30724 9812 30764
rect 9292 29128 9332 29168
rect 9292 28960 9332 29000
rect 9196 28372 9236 28412
rect 9196 28204 9236 28244
rect 9196 27952 9236 27992
rect 9004 27532 9044 27572
rect 8812 27196 8852 27236
rect 8908 26776 8948 26816
rect 9100 26356 9140 26396
rect 9004 26272 9044 26312
rect 9388 28540 9428 28580
rect 9676 29128 9716 29168
rect 10636 32068 10676 32108
rect 10540 30976 10580 31016
rect 10252 30724 10292 30764
rect 10444 30304 10484 30344
rect 10348 30136 10388 30176
rect 9868 29800 9908 29840
rect 9772 29044 9812 29084
rect 9580 28540 9620 28580
rect 9484 28204 9524 28244
rect 9676 28288 9716 28328
rect 9388 27532 9428 27572
rect 9388 27364 9428 27404
rect 9292 26356 9332 26396
rect 9580 28036 9620 28076
rect 9580 27700 9620 27740
rect 9772 27700 9812 27740
rect 9676 27532 9716 27572
rect 9580 26776 9620 26816
rect 8812 25516 8852 25556
rect 8908 25348 8948 25388
rect 8812 24508 8852 24548
rect 8521 22408 8561 22448
rect 8716 22408 8756 22448
rect 8620 22240 8660 22280
rect 8620 22072 8660 22112
rect 8428 20392 8468 20432
rect 7468 19216 7508 19256
rect 6892 17788 6932 17828
rect 6988 17452 7028 17492
rect 6892 15604 6932 15644
rect 7756 18544 7796 18584
rect 7660 18460 7700 18500
rect 7468 17620 7508 17660
rect 7756 17536 7796 17576
rect 7276 17200 7316 17240
rect 7468 16612 7508 16652
rect 7372 16360 7412 16400
rect 7180 15604 7220 15644
rect 7276 15520 7316 15560
rect 6700 15268 6740 15308
rect 6892 15100 6932 15140
rect 6604 14344 6644 14384
rect 6892 14008 6932 14048
rect 6412 13924 6452 13964
rect 6412 12916 6452 12956
rect 6124 11068 6164 11108
rect 6316 11656 6356 11696
rect 6220 10984 6260 11024
rect 6124 10900 6164 10940
rect 6220 8800 6260 8840
rect 6124 8128 6164 8168
rect 6316 6700 6356 6740
rect 6316 6196 6356 6236
rect 5932 5860 5972 5900
rect 5452 3676 5492 3716
rect 5644 4936 5684 4976
rect 5644 4600 5684 4640
rect 5836 5020 5876 5060
rect 5740 4348 5780 4388
rect 5644 4264 5684 4304
rect 5740 3676 5780 3716
rect 5548 3424 5588 3464
rect 5548 2668 5588 2708
rect 5452 2584 5492 2624
rect 5644 2584 5684 2624
rect 5548 2416 5588 2456
rect 5068 1072 5108 1112
rect 4204 400 4244 440
rect 4492 904 4532 944
rect 5260 904 5300 944
rect 4928 736 4968 776
rect 5010 736 5050 776
rect 5092 736 5132 776
rect 5174 736 5214 776
rect 5256 736 5296 776
rect 5356 736 5396 776
rect 5452 652 5492 692
rect 5068 568 5108 608
rect 4684 400 4724 440
rect 4876 232 4916 272
rect 5260 232 5300 272
rect 6124 5020 6164 5060
rect 5932 4600 5972 4640
rect 5932 4264 5972 4304
rect 6028 3508 6068 3548
rect 5932 2836 5972 2876
rect 5836 2668 5876 2708
rect 5932 2584 5972 2624
rect 5932 1408 5972 1448
rect 6028 232 6068 272
rect 6700 11320 6740 11360
rect 6892 10984 6932 11024
rect 6796 10900 6836 10940
rect 6604 10564 6644 10604
rect 6604 7456 6644 7496
rect 6796 10144 6836 10184
rect 7372 15436 7412 15476
rect 7276 14680 7316 14720
rect 7372 14092 7412 14132
rect 7756 15520 7796 15560
rect 7756 15268 7796 15308
rect 7660 15100 7700 15140
rect 8332 19132 8372 19172
rect 8428 18712 8468 18752
rect 8140 18376 8180 18416
rect 8428 18376 8468 18416
rect 7948 14932 7988 14972
rect 8524 17704 8564 17744
rect 8332 17116 8372 17156
rect 7852 14008 7892 14048
rect 7756 13756 7796 13796
rect 7660 13672 7700 13712
rect 7564 12160 7604 12200
rect 7372 11488 7412 11528
rect 7276 11320 7316 11360
rect 7468 11320 7508 11360
rect 7372 11152 7412 11192
rect 6988 10564 7028 10604
rect 6988 10312 7028 10352
rect 7180 10312 7220 10352
rect 6988 10144 7028 10184
rect 7180 10144 7220 10184
rect 6892 8464 6932 8504
rect 6892 7456 6932 7496
rect 6412 3424 6452 3464
rect 6892 6196 6932 6236
rect 6700 6028 6740 6068
rect 6700 4936 6740 4976
rect 6604 4264 6644 4304
rect 6508 2836 6548 2876
rect 7180 9724 7220 9764
rect 7084 8800 7124 8840
rect 7084 4936 7124 4976
rect 7084 4348 7124 4388
rect 7468 8464 7508 8504
rect 7372 7960 7412 8000
rect 8236 14680 8276 14720
rect 8332 14596 8372 14636
rect 8140 14428 8180 14468
rect 8044 13756 8084 13796
rect 7948 12160 7988 12200
rect 7852 11656 7892 11696
rect 7852 9640 7892 9680
rect 7852 9472 7892 9512
rect 7852 8716 7892 8756
rect 7564 7708 7604 7748
rect 7564 7456 7604 7496
rect 7564 6448 7604 6488
rect 7468 6196 7508 6236
rect 7372 5860 7412 5900
rect 7564 5608 7604 5648
rect 7468 5020 7508 5060
rect 7276 4936 7316 4976
rect 6796 3508 6836 3548
rect 6412 2332 6452 2372
rect 6604 1408 6644 1448
rect 6412 1240 6452 1280
rect 6988 1240 7028 1280
rect 7180 4012 7220 4052
rect 7564 4348 7604 4388
rect 8044 9388 8084 9428
rect 7948 7288 7988 7328
rect 7852 7204 7892 7244
rect 8044 7204 8084 7244
rect 8044 6952 8084 6992
rect 7948 5860 7988 5900
rect 7948 5524 7988 5564
rect 9100 25264 9140 25304
rect 9580 25432 9620 25472
rect 9580 25264 9620 25304
rect 9484 25180 9524 25220
rect 9100 24256 9140 24296
rect 8908 23836 8948 23876
rect 8908 23164 8948 23204
rect 8908 22996 8948 23036
rect 8716 21232 8756 21272
rect 9004 21820 9044 21860
rect 9484 24508 9524 24548
rect 10060 29800 10100 29840
rect 10540 29884 10580 29924
rect 10348 29632 10388 29672
rect 10444 29380 10484 29420
rect 10060 28288 10100 28328
rect 9964 28120 10004 28160
rect 10060 28036 10100 28076
rect 9868 26860 9908 26900
rect 10348 28456 10388 28496
rect 10348 28288 10388 28328
rect 10252 28204 10292 28244
rect 10444 28120 10484 28160
rect 10540 28036 10580 28076
rect 10444 27868 10484 27908
rect 10348 27700 10388 27740
rect 10252 26944 10292 26984
rect 10828 35596 10868 35636
rect 10828 35260 10868 35300
rect 11404 35764 11444 35804
rect 11308 35680 11348 35720
rect 11212 35596 11252 35636
rect 11116 35176 11156 35216
rect 10924 34924 10964 34964
rect 11116 34168 11156 34208
rect 11500 35176 11540 35216
rect 11404 35092 11444 35132
rect 11308 34924 11348 34964
rect 11404 33748 11444 33788
rect 11020 33076 11060 33116
rect 10924 31648 10964 31688
rect 10828 31312 10868 31352
rect 10732 28792 10772 28832
rect 10732 28540 10772 28580
rect 10924 30220 10964 30260
rect 11404 33328 11444 33368
rect 11500 33244 11540 33284
rect 11212 31228 11252 31268
rect 11212 30808 11252 30848
rect 11788 36604 11828 36644
rect 11788 35848 11828 35888
rect 11692 35428 11732 35468
rect 12172 39880 12212 39920
rect 12652 40300 12692 40340
rect 12748 39712 12788 39752
rect 13132 42652 13172 42692
rect 13132 42484 13172 42524
rect 12940 40048 12980 40088
rect 12940 39880 12980 39920
rect 13036 39712 13076 39752
rect 12268 39124 12308 39164
rect 12076 36940 12116 36980
rect 12076 36688 12116 36728
rect 12460 39124 12500 39164
rect 12556 39040 12596 39080
rect 12364 38956 12404 38996
rect 12556 38116 12596 38156
rect 12364 38032 12404 38072
rect 12460 36688 12500 36728
rect 12364 35680 12404 35720
rect 12172 35596 12212 35636
rect 11692 33916 11732 33956
rect 11692 33748 11732 33788
rect 11596 30220 11636 30260
rect 11404 29968 11444 30008
rect 11692 29968 11732 30008
rect 11020 28960 11060 29000
rect 11116 28456 11156 28496
rect 11020 28293 11060 28328
rect 11020 28288 11060 28293
rect 11404 29128 11444 29168
rect 11692 29044 11732 29084
rect 11596 28960 11636 29000
rect 11884 32404 11924 32444
rect 12364 33748 12404 33788
rect 12076 31816 12116 31856
rect 11980 31648 12020 31688
rect 12268 33580 12308 33620
rect 12268 32740 12308 32780
rect 12172 31480 12212 31520
rect 11884 30052 11924 30092
rect 11884 29800 11924 29840
rect 12172 31144 12212 31184
rect 12556 35680 12596 35720
rect 12556 35428 12596 35468
rect 12556 33832 12596 33872
rect 12940 39460 12980 39500
rect 12940 39292 12980 39332
rect 13036 39208 13076 39248
rect 13516 41644 13556 41684
rect 13900 41728 13940 41768
rect 14284 41644 14324 41684
rect 13324 41560 13364 41600
rect 13708 41560 13748 41600
rect 14092 41560 14132 41600
rect 14476 41560 14516 41600
rect 14668 41560 14708 41600
rect 13804 41392 13844 41432
rect 13612 41140 13652 41180
rect 13228 40636 13268 40676
rect 13612 40888 13652 40928
rect 13420 40384 13460 40424
rect 13516 40132 13556 40172
rect 13420 39208 13460 39248
rect 12844 39124 12884 39164
rect 13132 39124 13172 39164
rect 12748 37780 12788 37820
rect 13036 38116 13076 38156
rect 13420 37780 13460 37820
rect 13036 36352 13076 36392
rect 13036 35680 13076 35720
rect 12844 35512 12884 35552
rect 12748 34840 12788 34880
rect 12748 33748 12788 33788
rect 13036 35176 13076 35216
rect 12940 34504 12980 34544
rect 13132 35092 13172 35132
rect 13132 34252 13172 34292
rect 12844 33664 12884 33704
rect 12652 33328 12692 33368
rect 12844 33328 12884 33368
rect 12076 30724 12116 30764
rect 12364 30304 12404 30344
rect 12076 29800 12116 29840
rect 12076 29464 12116 29504
rect 12556 30388 12596 30428
rect 12460 30052 12500 30092
rect 11980 29044 12020 29084
rect 12748 31312 12788 31352
rect 11980 28876 12020 28916
rect 11788 28540 11828 28580
rect 11404 28456 11444 28496
rect 11692 28456 11732 28496
rect 11308 28372 11348 28412
rect 11788 28372 11828 28412
rect 11500 28120 11540 28160
rect 11692 28156 11732 28160
rect 11692 28120 11732 28156
rect 11212 28036 11252 28076
rect 10924 27196 10964 27236
rect 10828 26860 10868 26900
rect 10732 26776 10772 26816
rect 9964 26356 10004 26396
rect 9868 25432 9908 25472
rect 10060 25264 10100 25304
rect 10156 25180 10196 25220
rect 9676 24508 9716 24548
rect 9580 24004 9620 24044
rect 9388 23164 9428 23204
rect 9580 23164 9620 23204
rect 9292 22996 9332 23036
rect 9292 22492 9332 22532
rect 9292 22240 9332 22280
rect 9484 21484 9524 21524
rect 9772 22408 9812 22448
rect 9964 24928 10004 24968
rect 10060 24676 10100 24716
rect 10060 24088 10100 24128
rect 9964 23164 10004 23204
rect 10156 23080 10196 23120
rect 10156 22240 10196 22280
rect 9676 20560 9716 20600
rect 8812 19300 8852 19340
rect 8812 18628 8852 18668
rect 8620 16696 8660 16736
rect 8620 16444 8660 16484
rect 8908 17620 8948 17660
rect 10156 21400 10196 21440
rect 9868 21316 9908 21356
rect 9292 19636 9332 19676
rect 9196 19384 9236 19424
rect 9100 19300 9140 19340
rect 9004 16276 9044 16316
rect 9292 19048 9332 19088
rect 9196 17032 9236 17072
rect 9196 16444 9236 16484
rect 8908 15772 8948 15812
rect 8812 15520 8852 15560
rect 8716 14932 8756 14972
rect 8236 13924 8276 13964
rect 8236 12496 8276 12536
rect 8524 12412 8564 12452
rect 8524 11740 8564 11780
rect 8236 11488 8276 11528
rect 8428 11572 8468 11612
rect 8332 11152 8372 11192
rect 8716 13504 8756 13544
rect 8716 13252 8756 13292
rect 8716 12496 8756 12536
rect 8716 12160 8756 12200
rect 8428 10732 8468 10772
rect 8332 10228 8372 10268
rect 8236 9472 8276 9512
rect 8428 9976 8468 10016
rect 8428 9472 8468 9512
rect 8428 7204 8468 7244
rect 8620 10312 8660 10352
rect 8908 12580 8948 12620
rect 8908 12412 8948 12452
rect 9100 14596 9140 14636
rect 9004 11488 9044 11528
rect 8908 11320 8948 11360
rect 8812 10732 8852 10772
rect 8812 10564 8852 10604
rect 9004 11152 9044 11192
rect 9004 10564 9044 10604
rect 8908 10480 8948 10520
rect 8812 10396 8852 10436
rect 8716 9724 8756 9764
rect 8908 10312 8948 10352
rect 9292 16024 9332 16064
rect 9484 19636 9524 19676
rect 9580 19468 9620 19508
rect 9772 18880 9812 18920
rect 9676 18544 9716 18584
rect 9580 18040 9620 18080
rect 10444 26608 10484 26648
rect 10924 26608 10964 26648
rect 10444 25264 10484 25304
rect 10828 26356 10868 26396
rect 10828 26188 10868 26228
rect 10636 25432 10676 25472
rect 10348 23752 10388 23792
rect 10348 23080 10388 23120
rect 10348 22660 10388 22700
rect 10252 20140 10292 20180
rect 9964 19048 10004 19088
rect 10348 19132 10388 19172
rect 9964 18712 10004 18752
rect 9580 17032 9620 17072
rect 10060 18292 10100 18332
rect 10156 17704 10196 17744
rect 11116 26776 11156 26816
rect 11020 25180 11060 25220
rect 10828 25096 10868 25136
rect 11116 25096 11156 25136
rect 10924 24928 10964 24968
rect 10732 24676 10772 24716
rect 11980 27700 12020 27740
rect 11404 27364 11444 27404
rect 11500 26776 11540 26816
rect 11404 26608 11444 26648
rect 11308 26524 11348 26564
rect 10540 24424 10580 24464
rect 11212 24592 11252 24632
rect 10636 23836 10676 23876
rect 10636 23584 10676 23624
rect 11212 23584 11252 23624
rect 11020 23164 11060 23204
rect 10636 23080 10676 23120
rect 10540 22576 10580 22616
rect 11500 26440 11540 26480
rect 12364 28288 12404 28328
rect 12460 28120 12500 28160
rect 12652 28120 12692 28160
rect 12460 27784 12500 27824
rect 12172 27532 12212 27572
rect 12076 27196 12116 27236
rect 12076 26860 12116 26900
rect 11788 26776 11828 26816
rect 11692 26104 11732 26144
rect 12556 27532 12596 27572
rect 12460 27364 12500 27404
rect 12364 26860 12404 26900
rect 12268 26776 12308 26816
rect 11596 25600 11636 25640
rect 11884 25432 11924 25472
rect 11404 23920 11444 23960
rect 12268 25600 12308 25640
rect 11692 24676 11732 24716
rect 12076 24676 12116 24716
rect 11884 24592 11924 24632
rect 11596 23920 11636 23960
rect 11500 23248 11540 23288
rect 11404 22408 11444 22448
rect 11308 22324 11348 22364
rect 11500 22324 11540 22364
rect 11884 23416 11924 23456
rect 12076 23248 12116 23288
rect 11788 22744 11828 22784
rect 11692 22324 11732 22364
rect 11596 21988 11636 22028
rect 10540 21400 10580 21440
rect 11596 21568 11636 21608
rect 11596 21148 11636 21188
rect 11308 20728 11348 20768
rect 11116 20644 11156 20684
rect 11596 20392 11636 20432
rect 10636 20224 10676 20264
rect 10540 19300 10580 19340
rect 10540 19048 10580 19088
rect 10540 18292 10580 18332
rect 10444 16948 10484 16988
rect 9964 16612 10004 16652
rect 9772 16528 9812 16568
rect 9388 15772 9428 15812
rect 9388 15268 9428 15308
rect 9676 16108 9716 16148
rect 9772 16024 9812 16064
rect 9196 12580 9236 12620
rect 9196 10984 9236 11024
rect 9100 10312 9140 10352
rect 8716 8716 8756 8756
rect 8908 8800 8948 8840
rect 9388 10228 9428 10268
rect 9292 10144 9332 10184
rect 8812 7540 8852 7580
rect 9004 7960 9044 8000
rect 9196 7204 9236 7244
rect 8812 7120 8852 7160
rect 8236 6952 8276 6992
rect 8428 6868 8468 6908
rect 8140 5860 8180 5900
rect 8140 5608 8180 5648
rect 8044 5356 8084 5396
rect 7756 4852 7796 4892
rect 7468 3424 7508 3464
rect 7276 3340 7316 3380
rect 6604 904 6644 944
rect 6796 736 6836 776
rect 7372 1156 7412 1196
rect 7948 4684 7988 4724
rect 7852 4264 7892 4304
rect 7660 2836 7700 2876
rect 8044 2836 8084 2876
rect 7660 2164 7700 2204
rect 8524 5524 8564 5564
rect 8332 4936 8372 4976
rect 8428 4768 8468 4808
rect 8428 3928 8468 3968
rect 8812 6952 8852 6992
rect 8908 6868 8948 6908
rect 8812 5776 8852 5816
rect 8236 2248 8276 2288
rect 8140 2164 8180 2204
rect 7660 1324 7700 1364
rect 7852 1240 7892 1280
rect 7948 1156 7988 1196
rect 7660 904 7700 944
rect 7756 652 7796 692
rect 8044 568 8084 608
rect 8716 2500 8756 2540
rect 8620 2416 8660 2456
rect 8716 2332 8756 2372
rect 8524 1324 8564 1364
rect 8236 736 8276 776
rect 8332 568 8372 608
rect 8716 904 8756 944
rect 8620 820 8660 860
rect 9004 3424 9044 3464
rect 9772 12580 9812 12620
rect 9964 15268 10004 15308
rect 10156 16192 10196 16232
rect 10252 16108 10292 16148
rect 10156 15352 10196 15392
rect 10060 15100 10100 15140
rect 11116 20140 11156 20180
rect 11500 19888 11540 19928
rect 10924 18796 10964 18836
rect 10732 18124 10772 18164
rect 10828 18040 10868 18080
rect 10540 15856 10580 15896
rect 10636 15772 10676 15812
rect 10828 15772 10868 15812
rect 10348 15436 10388 15476
rect 10635 15436 10675 15476
rect 10156 14008 10196 14048
rect 10060 13588 10100 13628
rect 9580 11152 9620 11192
rect 9580 10984 9620 11024
rect 9580 10480 9620 10520
rect 9484 10144 9524 10184
rect 9484 9808 9524 9848
rect 9388 7792 9428 7832
rect 9388 7540 9428 7580
rect 9868 12496 9908 12536
rect 9772 12412 9812 12452
rect 10252 12496 10292 12536
rect 9772 11740 9812 11780
rect 9964 11740 10004 11780
rect 9676 10228 9716 10268
rect 9868 11488 9908 11528
rect 10060 11068 10100 11108
rect 10156 10564 10196 10604
rect 10060 10396 10100 10436
rect 9964 10312 10004 10352
rect 9868 8716 9908 8756
rect 9580 7792 9620 7832
rect 9772 7792 9812 7832
rect 9388 7036 9428 7076
rect 9388 6532 9428 6572
rect 9676 6532 9716 6572
rect 9580 6448 9620 6488
rect 9676 6196 9716 6236
rect 9964 7708 10004 7748
rect 9868 7456 9908 7496
rect 9868 7120 9908 7160
rect 10060 7540 10100 7580
rect 10156 7120 10196 7160
rect 10156 5860 10196 5900
rect 9676 5524 9716 5564
rect 9580 4936 9620 4976
rect 9964 5608 10004 5648
rect 9772 4852 9812 4892
rect 9964 4600 10004 4640
rect 9772 4096 9812 4136
rect 10156 4096 10196 4136
rect 10732 15352 10772 15392
rect 10636 15100 10676 15140
rect 10828 14680 10868 14720
rect 11596 19804 11636 19844
rect 11308 19300 11348 19340
rect 11116 19132 11156 19172
rect 11404 17620 11444 17660
rect 11116 17032 11156 17072
rect 11020 16864 11060 16904
rect 11980 22240 12020 22280
rect 12076 21484 12116 21524
rect 11980 20560 12020 20600
rect 12364 25180 12404 25220
rect 12268 22072 12308 22112
rect 12268 21064 12308 21104
rect 12364 20896 12404 20936
rect 12268 20728 12308 20768
rect 12172 20476 12212 20516
rect 11884 19972 11924 20012
rect 11788 18880 11828 18920
rect 11692 17116 11732 17156
rect 12172 19888 12212 19928
rect 12076 19804 12116 19844
rect 12076 19468 12116 19508
rect 11980 18544 12020 18584
rect 11884 17956 11924 17996
rect 11884 17620 11924 17660
rect 12076 17872 12116 17912
rect 12172 17788 12212 17828
rect 11980 17452 12020 17492
rect 11692 16780 11732 16820
rect 11116 15856 11156 15896
rect 11020 15604 11060 15644
rect 11020 15268 11060 15308
rect 10924 13168 10964 13208
rect 10924 12664 10964 12704
rect 10924 11572 10964 11612
rect 10348 10984 10388 11024
rect 10540 10648 10580 10688
rect 10540 10312 10580 10352
rect 10444 9976 10484 10016
rect 10636 9976 10676 10016
rect 10540 9304 10580 9344
rect 10444 7120 10484 7160
rect 10444 4264 10484 4304
rect 9868 3340 9908 3380
rect 9772 2668 9812 2708
rect 9292 2416 9332 2456
rect 9196 1912 9236 1952
rect 9100 1660 9140 1700
rect 8908 736 8948 776
rect 8812 652 8852 692
rect 9100 568 9140 608
rect 9580 2248 9620 2288
rect 10156 2500 10196 2540
rect 9868 1660 9908 1700
rect 9484 1240 9524 1280
rect 9388 1072 9428 1112
rect 9484 652 9524 692
rect 9676 400 9716 440
rect 10156 2248 10196 2288
rect 10060 1828 10100 1868
rect 10060 1576 10100 1616
rect 10252 1912 10292 1952
rect 10252 1072 10292 1112
rect 10156 484 10196 524
rect 10444 1828 10484 1868
rect 10636 8548 10676 8588
rect 10828 10900 10868 10940
rect 10828 8464 10868 8504
rect 10828 8044 10868 8084
rect 10732 5104 10772 5144
rect 11020 10564 11060 10604
rect 11596 15604 11636 15644
rect 11884 16192 11924 16232
rect 11788 15604 11828 15644
rect 11212 14680 11252 14720
rect 11404 12412 11444 12452
rect 11212 10816 11252 10856
rect 11308 10144 11348 10184
rect 11212 9388 11252 9428
rect 11020 8548 11060 8588
rect 11116 8044 11156 8084
rect 12172 16612 12212 16652
rect 12076 16444 12116 16484
rect 12076 15688 12116 15728
rect 11692 14043 11732 14048
rect 11692 14008 11732 14043
rect 11692 13756 11732 13796
rect 11884 14176 11924 14216
rect 11788 13672 11828 13712
rect 11788 12580 11828 12620
rect 11692 12412 11732 12452
rect 11596 11656 11636 11696
rect 12364 19300 12404 19340
rect 12364 18208 12404 18248
rect 12556 26104 12596 26144
rect 12652 23920 12692 23960
rect 13132 34084 13172 34124
rect 13036 33916 13076 33956
rect 13804 40636 13844 40676
rect 13804 40384 13844 40424
rect 13804 39628 13844 39668
rect 13900 39208 13940 39248
rect 13804 39040 13844 39080
rect 13612 38116 13652 38156
rect 13516 34504 13556 34544
rect 13516 34252 13556 34292
rect 13420 34168 13460 34208
rect 13708 35176 13748 35216
rect 14764 40972 14804 41012
rect 15148 40972 15188 41012
rect 14380 40636 14420 40676
rect 15820 40552 15860 40592
rect 15244 40468 15284 40508
rect 14380 40384 14420 40424
rect 14188 40216 14228 40256
rect 14092 39292 14132 39332
rect 14188 39208 14228 39248
rect 15628 40384 15668 40424
rect 15436 40300 15476 40340
rect 14860 40216 14900 40256
rect 14380 40048 14420 40088
rect 14380 39292 14420 39332
rect 13900 37360 13940 37400
rect 13324 33916 13364 33956
rect 13132 32824 13172 32864
rect 13036 32488 13076 32528
rect 12940 32152 12980 32192
rect 12940 30556 12980 30596
rect 12940 30388 12980 30428
rect 12844 28624 12884 28664
rect 13132 29632 13172 29672
rect 13324 32824 13364 32864
rect 13324 31228 13364 31268
rect 13324 30892 13364 30932
rect 13516 31648 13556 31688
rect 13420 30724 13460 30764
rect 13516 30220 13556 30260
rect 14284 37696 14324 37736
rect 14188 37360 14228 37400
rect 13900 34420 13940 34460
rect 13804 34336 13844 34376
rect 13804 33748 13844 33788
rect 13804 32740 13844 32780
rect 13708 32152 13748 32192
rect 13996 34336 14036 34376
rect 14188 34252 14228 34292
rect 14572 39628 14612 39668
rect 14668 39040 14708 39080
rect 14476 38872 14516 38912
rect 14476 37948 14516 37988
rect 14476 37780 14516 37820
rect 14380 34756 14420 34796
rect 15340 39292 15380 39332
rect 15148 38872 15188 38912
rect 15148 37864 15188 37904
rect 15052 37780 15092 37820
rect 14572 34420 14612 34460
rect 14956 36940 14996 36980
rect 15148 36772 15188 36812
rect 15628 38452 15668 38492
rect 15532 38200 15572 38240
rect 15340 36016 15380 36056
rect 14956 35512 14996 35552
rect 15436 35764 15476 35804
rect 15436 35428 15476 35468
rect 16108 41560 16148 41600
rect 16012 40468 16052 40508
rect 16108 40384 16148 40424
rect 16012 39712 16052 39752
rect 15820 38200 15860 38240
rect 15628 37864 15668 37904
rect 16588 41560 16628 41600
rect 16492 41476 16532 41516
rect 16396 40636 16436 40676
rect 17164 41644 17204 41684
rect 17356 41560 17396 41600
rect 16588 41140 16628 41180
rect 16780 41056 16820 41096
rect 16780 40384 16820 40424
rect 16684 40300 16724 40340
rect 16396 40132 16436 40172
rect 16300 39712 16340 39752
rect 16204 39292 16244 39332
rect 16204 39124 16244 39164
rect 16396 39040 16436 39080
rect 16204 37864 16244 37904
rect 16012 37612 16052 37652
rect 16396 37528 16436 37568
rect 16108 37276 16148 37316
rect 15820 37192 15860 37232
rect 16012 36604 16052 36644
rect 15820 36520 15860 36560
rect 15916 35848 15956 35888
rect 15820 35596 15860 35636
rect 15820 35428 15860 35468
rect 14956 35092 14996 35132
rect 14860 34756 14900 34796
rect 14764 34504 14804 34544
rect 14668 34336 14708 34376
rect 14476 34084 14516 34124
rect 14284 34000 14324 34040
rect 14092 33328 14132 33368
rect 14092 32908 14132 32948
rect 13612 30052 13652 30092
rect 13516 29968 13556 30008
rect 13996 31900 14036 31940
rect 14188 31900 14228 31940
rect 14572 32152 14612 32192
rect 15244 34672 15284 34712
rect 14668 32068 14708 32108
rect 14284 31732 14324 31772
rect 13996 30808 14036 30848
rect 13996 30640 14036 30680
rect 14668 31480 14708 31520
rect 14284 31312 14324 31352
rect 14188 30472 14228 30512
rect 14572 31312 14612 31352
rect 14860 31900 14900 31940
rect 14865 31312 14905 31352
rect 14764 31144 14804 31184
rect 14668 31060 14708 31100
rect 14476 30640 14516 30680
rect 13804 29968 13844 30008
rect 13132 28876 13172 28916
rect 12940 28120 12980 28160
rect 12844 27784 12884 27824
rect 13228 28624 13268 28664
rect 13036 27700 13076 27740
rect 13036 26188 13076 26228
rect 12844 26104 12884 26144
rect 12844 25684 12884 25724
rect 12844 23836 12884 23876
rect 12652 23500 12692 23540
rect 12556 22744 12596 22784
rect 12556 22408 12596 22448
rect 12556 21820 12596 21860
rect 12748 21652 12788 21692
rect 12556 20728 12596 20768
rect 12748 20056 12788 20096
rect 12940 20644 12980 20684
rect 12652 18460 12692 18500
rect 12652 18040 12692 18080
rect 12844 18544 12884 18584
rect 12940 18460 12980 18500
rect 12844 18040 12884 18080
rect 12460 17872 12500 17912
rect 12748 17872 12788 17912
rect 12460 17704 12500 17744
rect 12940 17872 12980 17912
rect 12556 17620 12596 17660
rect 12844 17704 12884 17744
rect 12844 17536 12884 17576
rect 12748 17368 12788 17408
rect 12460 16444 12500 16484
rect 12460 16192 12500 16232
rect 12268 15772 12308 15812
rect 12076 11740 12116 11780
rect 11884 11572 11924 11612
rect 11788 10816 11828 10856
rect 11692 10732 11732 10772
rect 11596 10396 11636 10436
rect 11596 9472 11636 9512
rect 11788 9640 11828 9680
rect 11788 9388 11828 9428
rect 11692 8884 11732 8924
rect 11596 8716 11636 8756
rect 11596 8128 11636 8168
rect 11692 7540 11732 7580
rect 11788 7204 11828 7244
rect 11596 7120 11636 7160
rect 11788 6532 11828 6572
rect 12364 14008 12404 14048
rect 12268 10816 12308 10856
rect 12268 10480 12308 10520
rect 12172 10228 12212 10268
rect 12172 9640 12212 9680
rect 12076 9388 12116 9428
rect 11980 8800 12020 8840
rect 12076 8716 12116 8756
rect 12076 8548 12116 8588
rect 12268 7708 12308 7748
rect 12268 7540 12308 7580
rect 12172 7204 12212 7244
rect 12172 7036 12212 7076
rect 12172 6868 12212 6908
rect 11596 6028 11636 6068
rect 11404 5608 11444 5648
rect 11212 5440 11252 5480
rect 11692 5608 11732 5648
rect 11404 5272 11444 5312
rect 11692 5272 11732 5312
rect 11020 4936 11060 4976
rect 11212 4936 11252 4976
rect 11404 4348 11444 4388
rect 11212 4264 11252 4304
rect 10828 3424 10868 3464
rect 11596 5020 11636 5060
rect 11404 3088 11444 3128
rect 11116 2668 11156 2708
rect 11692 4348 11732 4388
rect 11884 4180 11924 4220
rect 11788 3340 11828 3380
rect 10828 1660 10868 1700
rect 10732 1576 10772 1616
rect 10732 1324 10772 1364
rect 10636 1240 10676 1280
rect 10636 904 10676 944
rect 10444 820 10484 860
rect 10348 316 10388 356
rect 10828 1156 10868 1196
rect 11020 2416 11060 2456
rect 11212 1828 11252 1868
rect 11596 1828 11636 1868
rect 12652 16024 12692 16064
rect 12556 8800 12596 8840
rect 12844 15100 12884 15140
rect 12844 14932 12884 14972
rect 12844 13504 12884 13544
rect 13132 25096 13172 25136
rect 13228 24424 13268 24464
rect 13132 23836 13172 23876
rect 13324 23920 13364 23960
rect 13228 22240 13268 22280
rect 14092 29212 14132 29252
rect 13516 27112 13556 27152
rect 13612 26356 13652 26396
rect 13516 25264 13556 25304
rect 13612 25180 13652 25220
rect 14380 29800 14420 29840
rect 14572 29800 14612 29840
rect 14284 29464 14324 29504
rect 13804 28792 13844 28832
rect 13804 27784 13844 27824
rect 13804 26776 13844 26816
rect 13804 26356 13844 26396
rect 13804 25684 13844 25724
rect 13996 27700 14036 27740
rect 14188 27616 14228 27656
rect 14092 26776 14132 26816
rect 14476 29212 14516 29252
rect 14476 27700 14516 27740
rect 15148 34168 15188 34208
rect 15436 33664 15476 33704
rect 15340 33580 15380 33620
rect 15436 33076 15476 33116
rect 15628 32992 15668 33032
rect 15916 35092 15956 35132
rect 16012 34168 16052 34208
rect 15340 32824 15380 32864
rect 15052 31984 15092 32024
rect 15244 31396 15284 31436
rect 15148 31312 15188 31352
rect 16012 32992 16052 33032
rect 15916 32824 15956 32864
rect 15436 31480 15476 31520
rect 15052 31060 15092 31100
rect 15148 30976 15188 31016
rect 14956 30220 14996 30260
rect 14764 29212 14804 29252
rect 14668 28204 14708 28244
rect 14668 27364 14708 27404
rect 14572 27028 14612 27068
rect 14476 26776 14516 26816
rect 14380 26356 14420 26396
rect 14284 26272 14324 26312
rect 14476 26272 14516 26312
rect 14860 27028 14900 27068
rect 14668 26440 14708 26480
rect 15148 27616 15188 27656
rect 16012 31060 16052 31100
rect 16108 30976 16148 31016
rect 15724 30892 15764 30932
rect 15532 30556 15572 30596
rect 15724 30556 15764 30596
rect 15628 30220 15668 30260
rect 15340 29884 15380 29924
rect 15532 29716 15572 29756
rect 15532 28540 15572 28580
rect 16012 30388 16052 30428
rect 15916 29884 15956 29924
rect 15820 29296 15860 29336
rect 15724 29212 15764 29252
rect 15340 27700 15380 27740
rect 15436 27616 15476 27656
rect 15052 27196 15092 27236
rect 15244 27196 15284 27236
rect 15052 26944 15092 26984
rect 15820 27448 15860 27488
rect 15724 27196 15764 27236
rect 15916 27364 15956 27404
rect 14956 26440 14996 26480
rect 14284 25852 14324 25892
rect 14188 25684 14228 25724
rect 13900 25180 13940 25220
rect 13900 24592 13940 24632
rect 13708 24508 13748 24548
rect 13900 24424 13940 24464
rect 13708 23920 13748 23960
rect 13612 23332 13652 23372
rect 13804 23752 13844 23792
rect 13804 23584 13844 23624
rect 13900 23080 13940 23120
rect 13708 22324 13748 22364
rect 13612 21148 13652 21188
rect 13420 20980 13460 21020
rect 13612 20980 13652 21020
rect 13324 20728 13364 20768
rect 14092 25348 14132 25388
rect 14380 25180 14420 25220
rect 14572 24760 14612 24800
rect 14572 24592 14612 24632
rect 15148 26776 15188 26816
rect 15724 26944 15764 26984
rect 15340 26692 15380 26732
rect 15244 26272 15284 26312
rect 15052 26104 15092 26144
rect 14860 25600 14900 25640
rect 15052 25432 15092 25472
rect 14860 25180 14900 25220
rect 14764 24760 14804 24800
rect 15436 25684 15476 25724
rect 15340 25348 15380 25388
rect 15052 25180 15092 25220
rect 14956 24592 14996 24632
rect 14860 24508 14900 24548
rect 14380 24424 14420 24464
rect 14092 23752 14132 23792
rect 14188 23668 14228 23708
rect 14092 23584 14132 23624
rect 13996 21988 14036 22028
rect 14956 24340 14996 24380
rect 14572 24256 14612 24296
rect 14380 23500 14420 23540
rect 14380 23080 14420 23120
rect 14476 22660 14516 22700
rect 14380 22240 14420 22280
rect 14284 21988 14324 22028
rect 14188 20980 14228 21020
rect 13228 19888 13268 19928
rect 13228 19720 13268 19760
rect 13132 17704 13172 17744
rect 13132 16360 13172 16400
rect 13132 15604 13172 15644
rect 13036 14008 13076 14048
rect 12940 13252 12980 13292
rect 13900 19972 13940 20012
rect 13324 18544 13364 18584
rect 13324 16360 13364 16400
rect 14092 20140 14132 20180
rect 14380 20056 14420 20096
rect 13996 19720 14036 19760
rect 14092 19636 14132 19676
rect 13900 18544 13940 18584
rect 13804 17872 13844 17912
rect 13900 17788 13940 17828
rect 13324 16201 13364 16241
rect 13324 15940 13364 15980
rect 12940 12412 12980 12452
rect 13228 12496 13268 12536
rect 13132 12160 13172 12200
rect 12844 12076 12884 12116
rect 12844 11656 12884 11696
rect 13420 13924 13460 13964
rect 13612 16276 13652 16316
rect 13804 16192 13844 16232
rect 13708 15940 13748 15980
rect 13900 15520 13940 15560
rect 13420 13168 13460 13208
rect 13612 13168 13652 13208
rect 13324 10564 13364 10604
rect 12940 10228 12980 10268
rect 13132 10144 13172 10184
rect 12748 9556 12788 9596
rect 13036 8800 13076 8840
rect 12844 8716 12884 8756
rect 12844 8044 12884 8084
rect 12460 7120 12500 7160
rect 12556 6616 12596 6656
rect 12556 3928 12596 3968
rect 12364 2920 12404 2960
rect 12460 2248 12500 2288
rect 12844 7120 12884 7160
rect 13516 12496 13556 12536
rect 13804 14008 13844 14048
rect 13708 12160 13748 12200
rect 13516 10480 13556 10520
rect 13420 8296 13460 8336
rect 13324 7624 13364 7664
rect 13228 6784 13268 6824
rect 13036 6532 13076 6572
rect 12940 5608 12980 5648
rect 13420 5608 13460 5648
rect 13612 9052 13652 9092
rect 12748 4936 12788 4976
rect 12940 4936 12980 4976
rect 13516 5272 13556 5312
rect 12748 4096 12788 4136
rect 13228 3928 13268 3968
rect 12748 2668 12788 2708
rect 13420 3172 13460 3212
rect 13132 2668 13172 2708
rect 12748 2080 12788 2120
rect 11212 1156 11252 1196
rect 11308 1072 11348 1112
rect 10924 820 10964 860
rect 11212 904 11252 944
rect 10828 484 10868 524
rect 11020 484 11060 524
rect 11020 316 11060 356
rect 11404 904 11444 944
rect 11788 1240 11828 1280
rect 11500 820 11540 860
rect 11596 484 11636 524
rect 12652 1660 12692 1700
rect 12076 1324 12116 1364
rect 12652 1156 12692 1196
rect 11980 904 12020 944
rect 12172 820 12212 860
rect 12556 904 12596 944
rect 12460 400 12500 440
rect 12844 568 12884 608
rect 12748 484 12788 524
rect 13324 2164 13364 2204
rect 13036 1156 13076 1196
rect 13228 904 13268 944
rect 13132 400 13172 440
rect 13900 11656 13940 11696
rect 13900 10984 13940 11024
rect 13804 10564 13844 10604
rect 13804 10396 13844 10436
rect 13708 4936 13748 4976
rect 13900 10144 13940 10184
rect 13900 5692 13940 5732
rect 14380 19636 14420 19676
rect 14668 23757 14708 23792
rect 14668 23752 14708 23757
rect 15340 24760 15380 24800
rect 14860 23668 14900 23708
rect 14764 22245 14804 22280
rect 14764 22240 14804 22245
rect 14572 21568 14612 21608
rect 14668 21400 14708 21440
rect 14572 20980 14612 21020
rect 14284 19300 14324 19340
rect 14188 18880 14228 18920
rect 14284 18796 14324 18836
rect 14092 18544 14132 18584
rect 14188 18460 14228 18500
rect 14572 19216 14612 19256
rect 14956 21568 14996 21608
rect 14764 20560 14804 20600
rect 14764 20308 14804 20348
rect 14956 21148 14996 21188
rect 15820 26440 15860 26480
rect 15724 26272 15764 26312
rect 16396 36940 16436 36980
rect 16396 36520 16436 36560
rect 16972 40636 17012 40676
rect 16972 39712 17012 39752
rect 16876 39208 16916 39248
rect 16972 38956 17012 38996
rect 17644 41140 17684 41180
rect 17548 40636 17588 40676
rect 17548 40300 17588 40340
rect 17740 40804 17780 40844
rect 18316 41476 18356 41516
rect 18892 41644 18932 41684
rect 18796 41560 18836 41600
rect 18028 41140 18068 41180
rect 17932 40720 17972 40760
rect 17932 40384 17972 40424
rect 17644 39880 17684 39920
rect 17164 39040 17204 39080
rect 17068 38872 17108 38912
rect 16684 38368 16724 38408
rect 16684 38200 16724 38240
rect 17260 38200 17300 38240
rect 16588 38032 16628 38072
rect 16684 37696 16724 37736
rect 16588 37360 16628 37400
rect 16588 36604 16628 36644
rect 16492 36436 16532 36476
rect 16492 35260 16532 35300
rect 17164 38116 17204 38156
rect 16876 37948 16916 37988
rect 17164 37696 17204 37736
rect 17164 37276 17204 37316
rect 17164 36520 17204 36560
rect 16972 36436 17012 36476
rect 17068 36352 17108 36392
rect 16876 36100 16916 36140
rect 16780 35764 16820 35804
rect 16876 35680 16916 35720
rect 16684 35512 16724 35552
rect 16588 35092 16628 35132
rect 16396 33832 16436 33872
rect 16300 32824 16340 32864
rect 16492 32656 16532 32696
rect 17548 39040 17588 39080
rect 17740 39040 17780 39080
rect 17740 38872 17780 38912
rect 17548 38536 17588 38576
rect 17932 38872 17972 38912
rect 17836 38620 17876 38660
rect 17452 37948 17492 37988
rect 17452 37780 17492 37820
rect 17644 38032 17684 38072
rect 17548 37696 17588 37736
rect 17452 37276 17492 37316
rect 17356 37192 17396 37232
rect 17452 36688 17492 36728
rect 17356 36604 17396 36644
rect 17068 35344 17108 35384
rect 16972 34168 17012 34208
rect 16684 33916 16724 33956
rect 16876 33916 16916 33956
rect 16876 33748 16916 33788
rect 16684 33580 16724 33620
rect 16396 32068 16436 32108
rect 16972 32740 17012 32780
rect 16876 32656 16916 32696
rect 16396 31900 16436 31940
rect 16300 30472 16340 30512
rect 16684 31396 16724 31436
rect 16492 31312 16532 31352
rect 16684 31144 16724 31184
rect 16588 30640 16628 30680
rect 16204 28876 16244 28916
rect 16108 28540 16148 28580
rect 16108 27616 16148 27656
rect 16204 27196 16244 27236
rect 15724 25852 15764 25892
rect 15628 25096 15668 25136
rect 15244 23836 15284 23876
rect 15436 23752 15476 23792
rect 15820 25516 15860 25556
rect 15532 23668 15572 23708
rect 15244 23080 15284 23120
rect 15148 22744 15188 22784
rect 15724 23752 15764 23792
rect 16396 30304 16436 30344
rect 16588 28960 16628 29000
rect 16876 31900 16916 31940
rect 16876 31396 16916 31436
rect 17356 36100 17396 36140
rect 17932 38536 17972 38576
rect 17932 38284 17972 38324
rect 17836 38032 17876 38072
rect 17836 37024 17876 37064
rect 17740 36940 17780 36980
rect 17644 36520 17684 36560
rect 17164 33748 17204 33788
rect 17548 35092 17588 35132
rect 17644 35008 17684 35048
rect 17644 34504 17684 34544
rect 17260 33412 17300 33452
rect 18124 40636 18164 40676
rect 18220 40300 18260 40340
rect 18316 39880 18356 39920
rect 18508 41140 18548 41180
rect 18508 40720 18548 40760
rect 18700 41392 18740 41432
rect 19276 42064 19316 42104
rect 19276 41644 19316 41684
rect 19084 41140 19124 41180
rect 18700 40972 18740 41012
rect 18988 40972 19028 41012
rect 18808 40804 18848 40844
rect 18890 40804 18930 40844
rect 18972 40804 19012 40844
rect 19054 40804 19094 40844
rect 19136 40804 19176 40844
rect 20048 41560 20088 41600
rect 20130 41560 20170 41600
rect 20212 41560 20252 41600
rect 20294 41560 20334 41600
rect 20376 41560 20416 41600
rect 19756 41476 19796 41516
rect 19468 41392 19508 41432
rect 19372 41308 19412 41348
rect 19372 40888 19412 40928
rect 18700 39880 18740 39920
rect 18316 39628 18356 39668
rect 18220 39544 18260 39584
rect 18124 38704 18164 38744
rect 18124 38536 18164 38576
rect 18316 38284 18356 38324
rect 18316 37192 18356 37232
rect 18892 40636 18932 40676
rect 19564 40552 19604 40592
rect 18796 39628 18836 39668
rect 19084 39628 19124 39668
rect 19372 39796 19412 39836
rect 18808 39292 18848 39332
rect 18890 39292 18930 39332
rect 18972 39292 19012 39332
rect 19054 39292 19094 39332
rect 19136 39292 19176 39332
rect 18892 38956 18932 38996
rect 18508 38704 18548 38744
rect 18988 38872 19028 38912
rect 18796 38620 18836 38660
rect 18796 38284 18836 38324
rect 18508 37192 18548 37232
rect 18412 37024 18452 37064
rect 19948 40468 19988 40508
rect 20524 40384 20564 40424
rect 19852 39712 19892 39752
rect 19852 39544 19892 39584
rect 19468 39376 19508 39416
rect 19372 38872 19412 38912
rect 19180 38032 19220 38072
rect 19276 37948 19316 37988
rect 18808 37780 18848 37820
rect 18890 37780 18930 37820
rect 18972 37780 19012 37820
rect 19054 37780 19094 37820
rect 19136 37780 19176 37820
rect 19180 37612 19220 37652
rect 18700 37276 18740 37316
rect 18028 36100 18068 36140
rect 17836 35848 17876 35888
rect 18028 35176 18068 35216
rect 18220 36184 18260 36224
rect 18892 36856 18932 36896
rect 18124 34588 18164 34628
rect 17932 33916 17972 33956
rect 17260 32824 17300 32864
rect 17164 32236 17204 32276
rect 17164 31564 17204 31604
rect 17164 31312 17204 31352
rect 16876 31228 16916 31268
rect 16876 30640 16916 30680
rect 17068 31060 17108 31100
rect 16876 30472 16916 30512
rect 16780 29212 16820 29252
rect 16588 28036 16628 28076
rect 16492 27700 16532 27740
rect 16396 26944 16436 26984
rect 16300 26440 16340 26480
rect 16396 26272 16436 26312
rect 16204 26188 16244 26228
rect 16396 26104 16436 26144
rect 16204 26020 16244 26060
rect 16012 24508 16052 24548
rect 16300 25264 16340 25304
rect 16300 24592 16340 24632
rect 15916 23332 15956 23372
rect 15628 22744 15668 22784
rect 15820 22744 15860 22784
rect 15340 22324 15380 22364
rect 15244 22240 15284 22280
rect 16204 23332 16244 23372
rect 15916 22240 15956 22280
rect 15436 22156 15476 22196
rect 16108 22240 16148 22280
rect 15244 21148 15284 21188
rect 15148 20980 15188 21020
rect 15148 20560 15188 20600
rect 14476 18796 14516 18836
rect 14380 18460 14420 18500
rect 14092 17620 14132 17660
rect 14284 17620 14324 17660
rect 14380 17368 14420 17408
rect 14188 16276 14228 16316
rect 14380 16276 14420 16316
rect 14092 16192 14132 16232
rect 14092 16024 14132 16064
rect 14284 15100 14324 15140
rect 14188 14764 14228 14804
rect 14092 13420 14132 13460
rect 14284 11656 14324 11696
rect 14092 11404 14132 11444
rect 14284 11152 14324 11192
rect 14668 18712 14708 18752
rect 14668 18040 14708 18080
rect 14668 17704 14708 17744
rect 14668 16024 14708 16064
rect 14860 20056 14900 20096
rect 15052 20308 15092 20348
rect 15052 20140 15092 20180
rect 15532 21568 15572 21608
rect 16108 21568 16148 21608
rect 15628 21484 15668 21524
rect 15148 19300 15188 19340
rect 15052 18880 15092 18920
rect 14860 18712 14900 18752
rect 14860 17704 14900 17744
rect 15532 19221 15572 19256
rect 15532 19216 15572 19221
rect 15916 21400 15956 21440
rect 16108 21064 16148 21104
rect 15820 19384 15860 19424
rect 15724 19216 15764 19256
rect 16108 19300 16148 19340
rect 15532 18628 15572 18668
rect 15532 18208 15572 18248
rect 15436 18040 15476 18080
rect 15244 17872 15284 17912
rect 15532 17956 15572 17996
rect 15628 17620 15668 17660
rect 15340 16444 15380 16484
rect 15148 16360 15188 16400
rect 14668 14932 14708 14972
rect 14476 12496 14516 12536
rect 14380 10648 14420 10688
rect 14476 10396 14516 10436
rect 14284 10228 14324 10268
rect 14764 12244 14804 12284
rect 15340 14512 15380 14552
rect 15052 13924 15092 13964
rect 14956 13252 14996 13292
rect 15244 13168 15284 13208
rect 15052 12412 15092 12452
rect 15052 11740 15092 11780
rect 14668 11152 14708 11192
rect 14860 11152 14900 11192
rect 14380 10228 14420 10268
rect 14188 10144 14228 10184
rect 14764 10900 14804 10940
rect 14764 10396 14804 10436
rect 14284 9472 14324 9512
rect 14284 9052 14324 9092
rect 14188 8968 14228 9008
rect 14092 7708 14132 7748
rect 13900 4852 13940 4892
rect 13900 4516 13940 4556
rect 13996 3928 14036 3968
rect 14188 3256 14228 3296
rect 14380 8716 14420 8756
rect 14380 7876 14420 7916
rect 14380 7120 14420 7160
rect 14668 8464 14708 8504
rect 14572 8380 14612 8420
rect 14668 8128 14708 8168
rect 14476 6448 14516 6488
rect 14380 5776 14420 5816
rect 14380 4516 14420 4556
rect 14380 4348 14420 4388
rect 13708 2668 13748 2708
rect 14092 2668 14132 2708
rect 13804 2416 13844 2456
rect 13708 2332 13748 2372
rect 13612 1912 13652 1952
rect 13996 2332 14036 2372
rect 13900 2164 13940 2204
rect 13900 1744 13940 1784
rect 13420 1156 13460 1196
rect 13516 904 13556 944
rect 13612 484 13652 524
rect 14092 1828 14132 1868
rect 13804 1156 13844 1196
rect 14092 904 14132 944
rect 14092 652 14132 692
rect 14476 4096 14516 4136
rect 14380 2752 14420 2792
rect 14476 2668 14516 2708
rect 14284 2416 14324 2456
rect 14668 6616 14708 6656
rect 15148 11656 15188 11696
rect 15148 10564 15188 10604
rect 15052 9472 15092 9512
rect 15916 18628 15956 18668
rect 15916 17620 15956 17660
rect 15820 16864 15860 16904
rect 15820 15016 15860 15056
rect 15628 13840 15668 13880
rect 15532 13420 15572 13460
rect 15436 12664 15476 12704
rect 15436 11152 15476 11192
rect 15244 10228 15284 10268
rect 15148 9388 15188 9428
rect 14860 8800 14900 8840
rect 14860 7876 14900 7916
rect 14860 7624 14900 7664
rect 14860 6448 14900 6488
rect 14764 4768 14804 4808
rect 15820 12664 15860 12704
rect 16108 18460 16148 18500
rect 16108 18292 16148 18332
rect 16684 26776 16724 26816
rect 16588 26356 16628 26396
rect 16588 24592 16628 24632
rect 17356 32740 17396 32780
rect 17740 32740 17780 32780
rect 17356 31312 17396 31352
rect 17452 31060 17492 31100
rect 17260 30640 17300 30680
rect 17164 30556 17204 30596
rect 17068 30304 17108 30344
rect 17260 30304 17300 30344
rect 16972 29968 17012 30008
rect 16972 29800 17012 29840
rect 17164 29800 17204 29840
rect 17068 29716 17108 29756
rect 17164 29128 17204 29168
rect 17068 28456 17108 28496
rect 16972 28372 17012 28412
rect 17164 27700 17204 27740
rect 16876 27280 16916 27320
rect 17068 26440 17108 26480
rect 16972 26272 17012 26312
rect 16972 26104 17012 26144
rect 16876 25852 16916 25892
rect 16876 24508 16916 24548
rect 16492 24172 16532 24212
rect 16780 24172 16820 24212
rect 16492 23080 16532 23120
rect 16396 22240 16436 22280
rect 16492 20224 16532 20264
rect 16396 19888 16436 19928
rect 16396 19720 16436 19760
rect 16300 19384 16340 19424
rect 16300 18712 16340 18752
rect 16492 19636 16532 19676
rect 16492 19468 16532 19508
rect 16492 18712 16532 18752
rect 16396 18460 16436 18500
rect 16300 18376 16340 18416
rect 16300 17788 16340 17828
rect 16684 24004 16724 24044
rect 16684 20140 16724 20180
rect 16588 17704 16628 17744
rect 16396 17032 16436 17072
rect 16972 19300 17012 19340
rect 17164 25936 17204 25976
rect 17452 30556 17492 30596
rect 17356 29632 17396 29672
rect 17356 29464 17396 29504
rect 17452 28792 17492 28832
rect 17452 28624 17492 28664
rect 17836 31396 17876 31436
rect 17932 30640 17972 30680
rect 17836 29968 17876 30008
rect 18124 32152 18164 32192
rect 18808 36268 18848 36308
rect 18890 36268 18930 36308
rect 18972 36268 19012 36308
rect 19054 36268 19094 36308
rect 19136 36268 19176 36308
rect 19180 36016 19220 36056
rect 19756 38872 19796 38912
rect 19564 38788 19604 38828
rect 19468 38704 19508 38744
rect 19468 38452 19508 38492
rect 19564 37444 19604 37484
rect 19756 38200 19796 38240
rect 19660 37192 19700 37232
rect 19564 36856 19604 36896
rect 20048 40048 20088 40088
rect 20130 40048 20170 40088
rect 20212 40048 20252 40088
rect 20294 40048 20334 40088
rect 20376 40048 20416 40088
rect 20044 39460 20084 39500
rect 20332 38956 20372 38996
rect 20236 38872 20276 38912
rect 20044 38788 20084 38828
rect 20048 38536 20088 38576
rect 20130 38536 20170 38576
rect 20212 38536 20252 38576
rect 20294 38536 20334 38576
rect 20376 38536 20416 38576
rect 20044 37444 20084 37484
rect 21292 38956 21332 38996
rect 20812 38788 20852 38828
rect 20524 37528 20564 37568
rect 20236 37360 20276 37400
rect 19948 37108 19988 37148
rect 20048 37024 20088 37064
rect 20130 37024 20170 37064
rect 20212 37024 20252 37064
rect 20294 37024 20334 37064
rect 20376 37024 20416 37064
rect 19468 36772 19508 36812
rect 19756 36772 19796 36812
rect 19372 36268 19412 36308
rect 19660 36604 19700 36644
rect 18508 35596 18548 35636
rect 19084 35092 19124 35132
rect 18604 34840 18644 34880
rect 18808 34756 18848 34796
rect 18890 34756 18930 34796
rect 18972 34756 19012 34796
rect 19054 34756 19094 34796
rect 19136 34756 19176 34796
rect 19276 34672 19316 34712
rect 19276 34420 19316 34460
rect 19276 34000 19316 34040
rect 18808 33244 18848 33284
rect 18890 33244 18930 33284
rect 18972 33244 19012 33284
rect 19054 33244 19094 33284
rect 19136 33244 19176 33284
rect 19852 36688 19892 36728
rect 19948 36352 19988 36392
rect 20044 36100 20084 36140
rect 19852 35848 19892 35888
rect 19660 35260 19700 35300
rect 19468 34672 19508 34712
rect 19756 35092 19796 35132
rect 19564 34588 19604 34628
rect 19564 33664 19604 33704
rect 20140 35680 20180 35720
rect 20048 35512 20088 35552
rect 20130 35512 20170 35552
rect 20212 35512 20252 35552
rect 20294 35512 20334 35552
rect 20376 35512 20416 35552
rect 20140 35344 20180 35384
rect 20044 35260 20084 35300
rect 19948 35176 19988 35216
rect 20044 35008 20084 35048
rect 20236 35008 20276 35048
rect 19948 34420 19988 34460
rect 20140 34168 20180 34208
rect 20048 34000 20088 34040
rect 20130 34000 20170 34040
rect 20212 34000 20252 34040
rect 20294 34000 20334 34040
rect 20376 34000 20416 34040
rect 19948 33328 19988 33368
rect 19660 32992 19700 33032
rect 18220 31984 18260 32024
rect 19276 31984 19316 32024
rect 18808 31732 18848 31772
rect 18890 31732 18930 31772
rect 18972 31732 19012 31772
rect 19054 31732 19094 31772
rect 19136 31732 19176 31772
rect 20140 33160 20180 33200
rect 19948 32908 19988 32948
rect 20140 32656 20180 32696
rect 20716 36184 20756 36224
rect 20812 36016 20852 36056
rect 20716 34168 20756 34208
rect 20620 33496 20660 33536
rect 20620 33160 20660 33200
rect 20048 32488 20088 32528
rect 20130 32488 20170 32528
rect 20212 32488 20252 32528
rect 20294 32488 20334 32528
rect 20376 32488 20416 32528
rect 20524 32488 20564 32528
rect 19852 32152 19892 32192
rect 20044 32152 20084 32192
rect 19852 31984 19892 32024
rect 19660 31648 19700 31688
rect 19276 31480 19316 31520
rect 18316 31396 18356 31436
rect 19180 31396 19220 31436
rect 18124 31312 18164 31352
rect 18220 31228 18260 31268
rect 18508 31312 18548 31352
rect 18316 30808 18356 30848
rect 17548 28288 17588 28328
rect 17548 27280 17588 27320
rect 17356 25852 17396 25892
rect 17356 25600 17396 25640
rect 17260 24508 17300 24548
rect 17356 24172 17396 24212
rect 17452 24004 17492 24044
rect 17548 23920 17588 23960
rect 17644 23584 17684 23624
rect 17548 23248 17588 23288
rect 17260 23164 17300 23204
rect 17164 23080 17204 23120
rect 17356 22912 17396 22952
rect 17260 22240 17300 22280
rect 17164 21652 17204 21692
rect 17164 19552 17204 19592
rect 17644 23080 17684 23120
rect 17548 22828 17588 22868
rect 17644 22744 17684 22784
rect 17836 29632 17876 29672
rect 18028 29548 18068 29588
rect 18412 30052 18452 30092
rect 18412 29548 18452 29588
rect 17836 29128 17876 29168
rect 17836 27616 17876 27656
rect 18796 30808 18836 30848
rect 18508 29296 18548 29336
rect 19372 31312 19412 31352
rect 18988 31144 19028 31184
rect 18892 30472 18932 30512
rect 18808 30220 18848 30260
rect 18890 30220 18930 30260
rect 18972 30220 19012 30260
rect 19054 30220 19094 30260
rect 19136 30220 19176 30260
rect 18892 30052 18932 30092
rect 19468 30052 19508 30092
rect 18700 29800 18740 29840
rect 18700 29380 18740 29420
rect 18499 29128 18508 29168
rect 18508 29128 18539 29168
rect 18604 29128 18644 29168
rect 18604 28960 18644 29000
rect 18220 28120 18260 28160
rect 18220 27868 18260 27908
rect 18124 27616 18164 27656
rect 18028 27028 18068 27068
rect 18124 26944 18164 26984
rect 18028 26440 18068 26480
rect 17836 25936 17876 25976
rect 17932 25264 17972 25304
rect 18028 25180 18068 25220
rect 18124 23416 18164 23456
rect 17836 23332 17876 23372
rect 18124 23248 18164 23288
rect 17932 23164 17972 23204
rect 18316 27616 18356 27656
rect 20236 31480 20276 31520
rect 19756 31396 19796 31436
rect 20044 31396 20084 31436
rect 19660 30976 19700 31016
rect 19756 30388 19796 30428
rect 19660 30052 19700 30092
rect 19756 29800 19796 29840
rect 19180 29716 19220 29756
rect 18892 29296 18932 29336
rect 18988 29212 19028 29252
rect 19468 29128 19508 29168
rect 18988 29044 19028 29084
rect 19276 28960 19316 29000
rect 18508 27784 18548 27824
rect 18808 28708 18848 28748
rect 18890 28708 18930 28748
rect 18972 28708 19012 28748
rect 19054 28708 19094 28748
rect 19136 28708 19176 28748
rect 19180 27616 19220 27656
rect 18892 27448 18932 27488
rect 18808 27196 18848 27236
rect 18890 27196 18930 27236
rect 18972 27196 19012 27236
rect 19054 27196 19094 27236
rect 19136 27196 19176 27236
rect 18700 27112 18740 27152
rect 18412 26944 18452 26984
rect 19468 28120 19508 28160
rect 19564 27700 19604 27740
rect 18412 26776 18452 26816
rect 18412 26272 18452 26312
rect 18412 25180 18452 25220
rect 18604 26440 18644 26480
rect 18796 26776 18836 26816
rect 18988 26776 19028 26816
rect 18892 26440 18932 26480
rect 18988 26104 19028 26144
rect 18796 25936 18836 25976
rect 18700 25852 18740 25892
rect 19564 26608 19604 26648
rect 20048 30976 20088 31016
rect 20130 30976 20170 31016
rect 20212 30976 20252 31016
rect 20294 30976 20334 31016
rect 20376 30976 20416 31016
rect 20044 30640 20084 30680
rect 20236 29716 20276 29756
rect 19852 29548 19892 29588
rect 19948 29464 19988 29504
rect 20048 29464 20088 29504
rect 20130 29464 20170 29504
rect 20212 29464 20252 29504
rect 20294 29464 20334 29504
rect 20376 29464 20416 29504
rect 20716 30976 20756 31016
rect 20620 30472 20660 30512
rect 20620 29296 20660 29336
rect 20524 29212 20564 29252
rect 20524 29044 20564 29084
rect 19852 28960 19892 29000
rect 20236 28456 20276 28496
rect 20048 27952 20088 27992
rect 20130 27952 20170 27992
rect 20212 27952 20252 27992
rect 20294 27952 20334 27992
rect 20376 27952 20416 27992
rect 19948 27616 19988 27656
rect 19852 27364 19892 27404
rect 19948 26944 19988 26984
rect 19756 26692 19796 26732
rect 20048 26440 20088 26480
rect 20130 26440 20170 26480
rect 20212 26440 20252 26480
rect 20294 26440 20334 26480
rect 20376 26440 20416 26480
rect 19180 26272 19220 26312
rect 19372 26104 19412 26144
rect 18808 25684 18848 25724
rect 18890 25684 18930 25724
rect 18972 25684 19012 25724
rect 19054 25684 19094 25724
rect 19136 25684 19176 25724
rect 19372 25768 19412 25808
rect 18892 25348 18932 25388
rect 18700 25264 18740 25304
rect 18508 25096 18548 25136
rect 18796 25096 18836 25136
rect 19660 26020 19700 26060
rect 19852 25684 19892 25724
rect 19660 25348 19700 25388
rect 19180 25180 19220 25220
rect 19180 24592 19220 24632
rect 19756 25096 19796 25136
rect 18604 24424 18644 24464
rect 18316 24004 18356 24044
rect 17932 22744 17972 22784
rect 17740 22240 17780 22280
rect 17356 21064 17396 21104
rect 18028 22492 18068 22532
rect 17932 22240 17972 22280
rect 17548 21652 17588 21692
rect 17452 20392 17492 20432
rect 17356 19972 17396 20012
rect 17356 19132 17396 19172
rect 17260 18796 17300 18836
rect 17164 18544 17204 18584
rect 16972 17620 17012 17660
rect 16588 16192 16628 16232
rect 16300 15520 16340 15560
rect 16204 15352 16244 15392
rect 16108 14680 16148 14720
rect 16396 15100 16436 15140
rect 16300 15016 16340 15056
rect 16780 17032 16820 17072
rect 17452 17704 17492 17744
rect 17260 17620 17300 17660
rect 16780 16192 16820 16232
rect 16684 14764 16724 14804
rect 16492 14512 16532 14552
rect 15820 11740 15860 11780
rect 15724 11488 15764 11528
rect 15532 10900 15572 10940
rect 15724 9808 15764 9848
rect 15628 9724 15668 9764
rect 15532 9304 15572 9344
rect 15532 8968 15572 9008
rect 15436 8800 15476 8840
rect 15340 8380 15380 8420
rect 15052 7960 15092 8000
rect 15244 7960 15284 8000
rect 15244 7708 15284 7748
rect 15436 7624 15476 7664
rect 16204 11656 16244 11696
rect 16204 11488 16244 11528
rect 16012 11236 16052 11276
rect 16108 10900 16148 10940
rect 16012 10228 16052 10268
rect 16204 10480 16244 10520
rect 16012 9892 16052 9932
rect 16012 9472 16052 9512
rect 15628 8716 15668 8756
rect 15916 9304 15956 9344
rect 15820 8800 15860 8840
rect 15148 7036 15188 7076
rect 15820 7960 15860 8000
rect 14764 3676 14804 3716
rect 15244 5440 15284 5480
rect 15148 4516 15188 4556
rect 15052 4348 15092 4388
rect 16108 9388 16148 9428
rect 16012 8968 16052 9008
rect 16108 8800 16148 8840
rect 15916 7876 15956 7916
rect 15436 7120 15476 7160
rect 16012 7120 16052 7160
rect 15628 6616 15668 6656
rect 15820 6196 15860 6236
rect 16012 5608 16052 5648
rect 15820 5524 15860 5564
rect 15436 4096 15476 4136
rect 15532 4012 15572 4052
rect 14956 3256 14996 3296
rect 14764 3172 14804 3212
rect 14668 2416 14708 2456
rect 14284 1828 14324 1868
rect 14380 1660 14420 1700
rect 14572 1660 14612 1700
rect 14860 2668 14900 2708
rect 14860 1744 14900 1784
rect 14956 1492 14996 1532
rect 15436 3340 15476 3380
rect 15148 1912 15188 1952
rect 14764 1156 14804 1196
rect 14284 316 14324 356
rect 14668 820 14708 860
rect 14476 400 14516 440
rect 15148 1240 15188 1280
rect 15052 1156 15092 1196
rect 15148 904 15188 944
rect 14956 652 14996 692
rect 15436 3088 15476 3128
rect 15436 2752 15476 2792
rect 15340 2668 15380 2708
rect 15340 1912 15380 1952
rect 16012 5104 16052 5144
rect 16396 13420 16436 13460
rect 16396 12496 16436 12536
rect 16396 10396 16436 10436
rect 16396 9976 16436 10016
rect 16972 15520 17012 15560
rect 17164 15520 17204 15560
rect 17356 17536 17396 17576
rect 17356 16360 17396 16400
rect 17356 16192 17396 16232
rect 17356 15940 17396 15980
rect 17356 15772 17396 15812
rect 16876 15436 16916 15476
rect 17260 15436 17300 15476
rect 16684 13168 16724 13208
rect 16780 12580 16820 12620
rect 16588 11908 16628 11948
rect 16684 10396 16724 10436
rect 16588 9976 16628 10016
rect 16684 8968 16724 9008
rect 17356 14596 17396 14636
rect 17452 14512 17492 14552
rect 17260 14008 17300 14048
rect 17356 13420 17396 13460
rect 17356 13252 17396 13292
rect 17164 12496 17204 12536
rect 17068 12328 17108 12368
rect 16876 11992 16916 12032
rect 17260 11992 17300 12032
rect 16972 11740 17012 11780
rect 17068 11656 17108 11696
rect 16972 10816 17012 10856
rect 17356 11572 17396 11612
rect 17164 9640 17204 9680
rect 17452 10144 17492 10184
rect 17452 9640 17492 9680
rect 17260 8632 17300 8672
rect 16780 8548 16820 8588
rect 16588 7204 16628 7244
rect 16684 7120 16724 7160
rect 16396 7036 16436 7076
rect 16396 6784 16436 6824
rect 16108 4348 16148 4388
rect 16108 4180 16148 4220
rect 16012 4096 16052 4136
rect 15340 1660 15380 1700
rect 15244 736 15284 776
rect 16012 1408 16052 1448
rect 15436 1240 15476 1280
rect 15052 316 15092 356
rect 15628 652 15668 692
rect 15820 568 15860 608
rect 16300 6196 16340 6236
rect 16492 5356 16532 5396
rect 16492 4180 16532 4220
rect 16684 4180 16724 4220
rect 16876 8464 16916 8504
rect 16876 8128 16916 8168
rect 16876 6784 16916 6824
rect 17452 9052 17492 9092
rect 17356 8128 17396 8168
rect 17836 21568 17876 21608
rect 17740 21064 17780 21104
rect 17932 19972 17972 20012
rect 17740 19216 17780 19256
rect 17836 19048 17876 19088
rect 17740 18292 17780 18332
rect 17932 18124 17972 18164
rect 18220 22576 18260 22616
rect 18220 22240 18260 22280
rect 18124 21820 18164 21860
rect 18124 20728 18164 20768
rect 18124 20056 18164 20096
rect 18508 23752 18548 23792
rect 18808 24172 18848 24212
rect 18890 24172 18930 24212
rect 18972 24172 19012 24212
rect 19054 24172 19094 24212
rect 19136 24172 19176 24212
rect 19852 24592 19892 24632
rect 19852 24424 19892 24464
rect 19660 24088 19700 24128
rect 18988 24004 19028 24044
rect 18412 23668 18452 23708
rect 18892 23752 18932 23792
rect 19276 23920 19316 23960
rect 19660 23920 19700 23960
rect 18796 23584 18836 23624
rect 18604 23500 18644 23540
rect 18508 23248 18548 23288
rect 18700 23164 18740 23204
rect 18604 22912 18644 22952
rect 18412 22744 18452 22784
rect 18796 22912 18836 22952
rect 19564 23752 19604 23792
rect 19084 23164 19124 23204
rect 18892 22828 18932 22868
rect 18808 22660 18848 22700
rect 18890 22660 18930 22700
rect 18972 22660 19012 22700
rect 19054 22660 19094 22700
rect 19136 22660 19176 22700
rect 18892 22408 18932 22448
rect 18508 22240 18548 22280
rect 18412 21652 18452 21692
rect 19180 22240 19220 22280
rect 19468 22408 19508 22448
rect 20236 25936 20276 25976
rect 20044 25516 20084 25556
rect 20044 25264 20084 25304
rect 20048 24928 20088 24968
rect 20130 24928 20170 24968
rect 20212 24928 20252 24968
rect 20294 24928 20334 24968
rect 20376 24928 20416 24968
rect 20236 24760 20276 24800
rect 20140 23584 20180 23624
rect 19660 22408 19700 22448
rect 18700 21736 18740 21776
rect 18508 21568 18548 21608
rect 18808 21148 18848 21188
rect 18890 21148 18930 21188
rect 18972 21148 19012 21188
rect 19054 21148 19094 21188
rect 19136 21148 19176 21188
rect 18412 20728 18452 20768
rect 18412 20056 18452 20096
rect 18220 19804 18260 19844
rect 18124 18544 18164 18584
rect 17644 14176 17684 14216
rect 17644 13420 17684 13460
rect 17644 9472 17684 9512
rect 18892 20056 18932 20096
rect 19180 20560 19220 20600
rect 19180 20056 19220 20096
rect 18808 19636 18848 19676
rect 18890 19636 18930 19676
rect 18972 19636 19012 19676
rect 19054 19636 19094 19676
rect 19136 19636 19176 19676
rect 19276 19636 19316 19676
rect 19084 19216 19124 19256
rect 18700 18712 18740 18752
rect 18892 18712 18932 18752
rect 19084 18880 19124 18920
rect 18412 18460 18452 18500
rect 18808 18124 18848 18164
rect 18890 18124 18930 18164
rect 18972 18124 19012 18164
rect 19054 18124 19094 18164
rect 19136 18124 19176 18164
rect 18220 17704 18260 17744
rect 18988 17704 19028 17744
rect 19084 17620 19124 17660
rect 18220 16360 18260 16400
rect 18124 16192 18164 16232
rect 17836 15688 17876 15728
rect 17836 15555 17876 15560
rect 17836 15520 17876 15555
rect 18124 15688 18164 15728
rect 17932 15184 17972 15224
rect 17836 13924 17876 13964
rect 18124 14932 18164 14972
rect 18028 13420 18068 13460
rect 18316 15100 18356 15140
rect 18700 16948 18740 16988
rect 18508 16360 18548 16400
rect 18604 16192 18644 16232
rect 18316 14176 18356 14216
rect 18220 13252 18260 13292
rect 17932 11488 17972 11528
rect 18028 10816 18068 10856
rect 18316 11488 18356 11528
rect 18220 11152 18260 11192
rect 17932 10564 17972 10604
rect 18124 10564 18164 10604
rect 17836 9808 17876 9848
rect 17548 8800 17588 8840
rect 17740 8800 17780 8840
rect 17644 8128 17684 8168
rect 17260 7876 17300 7916
rect 17068 7036 17108 7076
rect 17068 6448 17108 6488
rect 17356 6112 17396 6152
rect 16972 5608 17012 5648
rect 16780 4096 16820 4136
rect 16684 3592 16724 3632
rect 16780 3424 16820 3464
rect 16588 2605 16628 2624
rect 16588 2584 16628 2605
rect 16972 3424 17012 3464
rect 16684 2500 16724 2540
rect 16300 1828 16340 1868
rect 16588 1996 16628 2036
rect 16588 1744 16628 1784
rect 16780 1912 16820 1952
rect 16876 1828 16916 1868
rect 16780 1660 16820 1700
rect 16684 1072 16724 1112
rect 16972 1072 17012 1112
rect 17164 4348 17204 4388
rect 17548 5692 17588 5732
rect 18028 10060 18068 10100
rect 18028 9388 18068 9428
rect 17932 8128 17972 8168
rect 17836 7708 17876 7748
rect 17932 7456 17972 7496
rect 18220 10149 18260 10184
rect 18220 10144 18260 10149
rect 18412 10816 18452 10856
rect 18508 10396 18548 10436
rect 18508 8968 18548 9008
rect 18220 8464 18260 8504
rect 18508 8716 18548 8756
rect 18508 8464 18548 8504
rect 18124 8128 18164 8168
rect 18316 7960 18356 8000
rect 18316 7792 18356 7832
rect 18124 7456 18164 7496
rect 18124 7288 18164 7328
rect 18028 7204 18068 7244
rect 17740 6700 17780 6740
rect 17932 5692 17972 5732
rect 17644 5524 17684 5564
rect 17548 5356 17588 5396
rect 18124 5608 18164 5648
rect 18808 16612 18848 16652
rect 18890 16612 18930 16652
rect 18972 16612 19012 16652
rect 19054 16612 19094 16652
rect 19136 16612 19176 16652
rect 19564 20728 19604 20768
rect 19564 20140 19604 20180
rect 19564 19552 19604 19592
rect 19852 23080 19892 23120
rect 20048 23416 20088 23456
rect 20130 23416 20170 23456
rect 20212 23416 20252 23456
rect 20294 23416 20334 23456
rect 20376 23416 20416 23456
rect 19948 22408 19988 22448
rect 19948 22240 19988 22280
rect 20048 21904 20088 21944
rect 20130 21904 20170 21944
rect 20212 21904 20252 21944
rect 20294 21904 20334 21944
rect 20376 21904 20416 21944
rect 19948 21568 19988 21608
rect 19852 21400 19892 21440
rect 21388 38872 21428 38912
rect 21292 35008 21332 35048
rect 21388 34000 21428 34040
rect 21292 32656 21332 32696
rect 21100 30220 21140 30260
rect 20812 29044 20852 29084
rect 20620 27952 20660 27992
rect 20812 27364 20852 27404
rect 20812 21904 20852 21944
rect 19756 20812 19796 20852
rect 19948 20728 19988 20768
rect 19756 20560 19796 20600
rect 20140 20560 20180 20600
rect 20048 20392 20088 20432
rect 20130 20392 20170 20432
rect 20212 20392 20252 20432
rect 20294 20392 20334 20432
rect 20376 20392 20416 20432
rect 19660 19048 19700 19088
rect 19948 20056 19988 20096
rect 19852 19636 19892 19676
rect 19948 19384 19988 19424
rect 20140 19552 20180 19592
rect 20236 19384 20276 19424
rect 20048 18880 20088 18920
rect 20130 18880 20170 18920
rect 20212 18880 20252 18920
rect 20294 18880 20334 18920
rect 20376 18880 20416 18920
rect 19756 18712 19796 18752
rect 19468 18208 19508 18248
rect 19276 16444 19316 16484
rect 18796 16192 18836 16232
rect 18808 15100 18848 15140
rect 18890 15100 18930 15140
rect 18972 15100 19012 15140
rect 19054 15100 19094 15140
rect 19136 15100 19176 15140
rect 18892 14764 18932 14804
rect 19372 14680 19412 14720
rect 19084 14596 19124 14636
rect 19276 14008 19316 14048
rect 19084 13840 19124 13880
rect 18808 13588 18848 13628
rect 18890 13588 18930 13628
rect 18972 13588 19012 13628
rect 19054 13588 19094 13628
rect 19136 13588 19176 13628
rect 18700 13252 18740 13292
rect 18892 13420 18932 13460
rect 19372 13504 19412 13544
rect 18892 12244 18932 12284
rect 18808 12076 18848 12116
rect 18890 12076 18930 12116
rect 18972 12076 19012 12116
rect 19054 12076 19094 12116
rect 19136 12076 19176 12116
rect 18988 11908 19028 11948
rect 18892 11824 18932 11864
rect 19276 11824 19316 11864
rect 18700 11404 18740 11444
rect 18700 10984 18740 11024
rect 18808 10564 18848 10604
rect 18890 10564 18930 10604
rect 18972 10564 19012 10604
rect 19054 10564 19094 10604
rect 19136 10564 19176 10604
rect 18700 10480 18740 10520
rect 19180 10228 19220 10268
rect 18796 10060 18836 10100
rect 19084 9640 19124 9680
rect 20236 17956 20276 17996
rect 19852 17704 19892 17744
rect 19660 16948 19700 16988
rect 19564 16864 19604 16904
rect 20048 17368 20088 17408
rect 20130 17368 20170 17408
rect 20212 17368 20252 17408
rect 20294 17368 20334 17408
rect 20376 17368 20416 17408
rect 20044 16360 20084 16400
rect 19756 15940 19796 15980
rect 20048 15856 20088 15896
rect 20130 15856 20170 15896
rect 20212 15856 20252 15896
rect 20294 15856 20334 15896
rect 20376 15856 20416 15896
rect 20620 19384 20660 19424
rect 20620 17368 20660 17408
rect 21196 27532 21236 27572
rect 21388 29212 21428 29252
rect 21388 28960 21428 29000
rect 21388 25684 21428 25724
rect 21388 25432 21428 25472
rect 21388 24256 21428 24296
rect 21388 23920 21428 23960
rect 21292 19888 21332 19928
rect 21196 18376 21236 18416
rect 21100 15856 21140 15896
rect 19756 12496 19796 12536
rect 19468 11656 19508 11696
rect 19756 11488 19796 11528
rect 19564 11152 19604 11192
rect 19372 9388 19412 9428
rect 20048 14344 20088 14384
rect 20130 14344 20170 14384
rect 20212 14344 20252 14384
rect 20294 14344 20334 14384
rect 20376 14344 20416 14384
rect 20140 13000 20180 13040
rect 20048 12832 20088 12872
rect 20130 12832 20170 12872
rect 20212 12832 20252 12872
rect 20294 12832 20334 12872
rect 20376 12832 20416 12872
rect 19948 12496 19988 12536
rect 19852 11152 19892 11192
rect 20048 11320 20088 11360
rect 20130 11320 20170 11360
rect 20212 11320 20252 11360
rect 20294 11320 20334 11360
rect 20376 11320 20416 11360
rect 19660 10648 19700 10688
rect 18808 9052 18848 9092
rect 18890 9052 18930 9092
rect 18972 9052 19012 9092
rect 19054 9052 19094 9092
rect 19136 9052 19176 9092
rect 18700 8296 18740 8336
rect 19372 9220 19412 9260
rect 19276 8632 19316 8672
rect 19948 10144 19988 10184
rect 19756 9640 19796 9680
rect 20048 9808 20088 9848
rect 20130 9808 20170 9848
rect 20212 9808 20252 9848
rect 20294 9808 20334 9848
rect 20376 9808 20416 9848
rect 19948 8632 19988 8672
rect 20048 8296 20088 8336
rect 20130 8296 20170 8336
rect 20212 8296 20252 8336
rect 20294 8296 20334 8336
rect 20376 8296 20416 8336
rect 19276 7960 19316 8000
rect 18700 7876 18740 7916
rect 18604 7036 18644 7076
rect 18220 5020 18260 5060
rect 17836 4768 17876 4808
rect 17740 4432 17780 4472
rect 17548 4180 17588 4220
rect 17740 4096 17780 4136
rect 17260 3424 17300 3464
rect 18796 7708 18836 7748
rect 18808 7540 18848 7580
rect 18890 7540 18930 7580
rect 18972 7540 19012 7580
rect 19054 7540 19094 7580
rect 19136 7540 19176 7580
rect 19372 7120 19412 7160
rect 19564 6952 19604 6992
rect 18808 6028 18848 6068
rect 18890 6028 18930 6068
rect 18972 6028 19012 6068
rect 19054 6028 19094 6068
rect 19136 6028 19176 6068
rect 18700 5020 18740 5060
rect 18604 4936 18644 4976
rect 18808 4516 18848 4556
rect 18890 4516 18930 4556
rect 18972 4516 19012 4556
rect 19054 4516 19094 4556
rect 19136 4516 19176 4556
rect 18796 4348 18836 4388
rect 17836 3676 17876 3716
rect 18028 3676 18068 3716
rect 17932 3508 17972 3548
rect 17356 1156 17396 1196
rect 17740 1156 17780 1196
rect 17164 904 17204 944
rect 17356 904 17396 944
rect 17548 820 17588 860
rect 19276 4096 19316 4136
rect 18316 4012 18356 4052
rect 18508 4012 18548 4052
rect 18412 3508 18452 3548
rect 18220 2584 18260 2624
rect 18604 3928 18644 3968
rect 19468 3592 19508 3632
rect 18808 3004 18848 3044
rect 18890 3004 18930 3044
rect 18972 3004 19012 3044
rect 19054 3004 19094 3044
rect 19136 3004 19176 3044
rect 19948 7372 19988 7412
rect 20048 6784 20088 6824
rect 20130 6784 20170 6824
rect 20212 6784 20252 6824
rect 20294 6784 20334 6824
rect 20376 6784 20416 6824
rect 19948 6280 19988 6320
rect 19756 5776 19796 5816
rect 19948 5440 19988 5480
rect 20048 5272 20088 5312
rect 20130 5272 20170 5312
rect 20212 5272 20252 5312
rect 20294 5272 20334 5312
rect 20376 5272 20416 5312
rect 20524 4852 20564 4892
rect 19852 4768 19892 4808
rect 20524 4264 20564 4304
rect 19948 4180 19988 4220
rect 20048 3760 20088 3800
rect 20130 3760 20170 3800
rect 20212 3760 20252 3800
rect 20294 3760 20334 3800
rect 20376 3760 20416 3800
rect 20044 3592 20084 3632
rect 19756 3340 19796 3380
rect 19564 2836 19604 2876
rect 18604 2668 18644 2708
rect 19948 3340 19988 3380
rect 18028 1660 18068 1700
rect 20044 2836 20084 2876
rect 20048 2248 20088 2288
rect 20130 2248 20170 2288
rect 20212 2248 20252 2288
rect 20294 2248 20334 2288
rect 20376 2248 20416 2288
rect 18808 1492 18848 1532
rect 18890 1492 18930 1532
rect 18972 1492 19012 1532
rect 19054 1492 19094 1532
rect 19136 1492 19176 1532
rect 18892 1324 18932 1364
rect 18508 1240 18548 1280
rect 17932 988 17972 1028
rect 17932 652 17972 692
rect 18124 652 18164 692
rect 18316 652 18356 692
rect 18508 652 18548 692
rect 18220 316 18260 356
rect 18700 484 18740 524
rect 20716 13336 20756 13376
rect 20716 10396 20756 10436
rect 21388 4768 21428 4808
rect 21388 4432 21428 4472
rect 19084 1240 19124 1280
rect 20620 1240 20660 1280
rect 20048 736 20088 776
rect 20130 736 20170 776
rect 20212 736 20252 776
rect 20294 736 20334 776
rect 20376 736 20416 776
rect 19468 652 19508 692
rect 19276 568 19316 608
<< metal3 >>
rect 1603 42904 1612 42944
rect 1652 42904 1804 42944
rect 1844 42904 1853 42944
rect 0 42776 80 42796
rect 1603 42776 1661 42777
rect 0 42736 1612 42776
rect 1652 42736 1661 42776
rect 0 42716 80 42736
rect 1603 42735 1661 42736
rect 11395 42692 11453 42693
rect 11395 42652 11404 42692
rect 11444 42652 13132 42692
rect 13172 42652 13181 42692
rect 11395 42651 11453 42652
rect 4771 42608 4829 42609
rect 2500 42568 4780 42608
rect 4820 42568 4829 42608
rect 9571 42568 9580 42608
rect 9620 42568 12364 42608
rect 12404 42568 12413 42608
rect 0 42440 80 42460
rect 2500 42440 2540 42568
rect 4771 42567 4829 42568
rect 3715 42484 3724 42524
rect 3764 42484 13132 42524
rect 13172 42484 13181 42524
rect 0 42400 2540 42440
rect 3043 42400 3052 42440
rect 3092 42400 5644 42440
rect 5684 42400 5693 42440
rect 0 42380 80 42400
rect 1795 42316 1804 42356
rect 1844 42316 4492 42356
rect 4532 42316 4541 42356
rect 7747 42272 7805 42273
rect 1603 42232 1612 42272
rect 1652 42232 4300 42272
rect 4340 42232 4349 42272
rect 7747 42232 7756 42272
rect 7796 42232 9292 42272
rect 9332 42232 9341 42272
rect 7747 42231 7805 42232
rect 14659 42188 14717 42189
rect 3427 42148 3436 42188
rect 3476 42148 6028 42188
rect 6068 42148 6077 42188
rect 8899 42148 8908 42188
rect 8948 42148 14668 42188
rect 14708 42148 14717 42188
rect 14659 42147 14717 42148
rect 0 42104 80 42124
rect 0 42064 2540 42104
rect 4867 42064 4876 42104
rect 4916 42064 9292 42104
rect 9332 42064 9341 42104
rect 9388 42064 11404 42104
rect 11444 42064 11453 42104
rect 11875 42064 11884 42104
rect 11924 42064 19276 42104
rect 19316 42064 19325 42104
rect 0 42044 80 42064
rect 2500 42020 2540 42064
rect 9388 42020 9428 42064
rect 2500 41980 5356 42020
rect 5396 41980 5405 42020
rect 9187 41980 9196 42020
rect 9236 41980 9428 42020
rect 6979 41896 6988 41936
rect 7028 41896 9964 41936
rect 10004 41896 10013 41936
rect 2563 41812 2572 41852
rect 2612 41812 10348 41852
rect 10388 41812 10397 41852
rect 0 41768 80 41788
rect 8035 41768 8093 41769
rect 0 41728 2540 41768
rect 4195 41728 4204 41768
rect 4244 41728 5260 41768
rect 5300 41728 5309 41768
rect 7747 41728 7756 41768
rect 7796 41728 8044 41768
rect 8084 41728 8093 41768
rect 0 41708 80 41728
rect 2500 41600 2540 41728
rect 8035 41727 8093 41728
rect 13603 41768 13661 41769
rect 13603 41728 13612 41768
rect 13652 41728 13900 41768
rect 13940 41728 13949 41768
rect 13603 41727 13661 41728
rect 7843 41684 7901 41685
rect 13795 41684 13853 41685
rect 15043 41684 15101 41685
rect 18691 41684 18749 41685
rect 2659 41644 2668 41684
rect 2708 41644 3148 41684
rect 3188 41644 3197 41684
rect 4675 41644 4684 41684
rect 4724 41644 7084 41684
rect 7124 41644 7133 41684
rect 7555 41644 7564 41684
rect 7604 41644 7852 41684
rect 7892 41644 7901 41684
rect 11299 41644 11308 41684
rect 11348 41644 11357 41684
rect 13507 41644 13516 41684
rect 13556 41644 13804 41684
rect 13844 41644 13853 41684
rect 14275 41644 14284 41684
rect 14324 41644 15052 41684
rect 15092 41644 15101 41684
rect 17155 41644 17164 41684
rect 17204 41644 18700 41684
rect 18740 41644 18749 41684
rect 18883 41644 18892 41684
rect 18932 41644 19276 41684
rect 19316 41644 19325 41684
rect 7843 41643 7901 41644
rect 7459 41600 7517 41601
rect 9475 41600 9533 41601
rect 11203 41600 11261 41601
rect 2500 41560 4588 41600
rect 4628 41560 4637 41600
rect 4919 41560 4928 41600
rect 4968 41560 5010 41600
rect 5050 41560 5092 41600
rect 5132 41560 5174 41600
rect 5214 41560 5256 41600
rect 5296 41560 5305 41600
rect 6028 41560 6508 41600
rect 6548 41560 6557 41600
rect 7363 41560 7372 41600
rect 7412 41560 7468 41600
rect 7508 41560 7517 41600
rect 8131 41560 8140 41600
rect 8180 41560 9332 41600
rect 9390 41560 9484 41600
rect 9524 41560 9533 41600
rect 10435 41560 10444 41600
rect 10484 41560 11212 41600
rect 11252 41560 11261 41600
rect 11308 41600 11348 41644
rect 13795 41643 13853 41644
rect 15043 41643 15101 41644
rect 18691 41643 18749 41644
rect 12547 41600 12605 41601
rect 13411 41600 13469 41601
rect 13699 41600 13757 41601
rect 14083 41600 14141 41601
rect 14467 41600 14525 41601
rect 14851 41600 14909 41601
rect 16675 41600 16733 41601
rect 11308 41560 11924 41600
rect 12462 41560 12556 41600
rect 12596 41560 12605 41600
rect 13315 41560 13324 41600
rect 13364 41560 13420 41600
rect 13460 41560 13469 41600
rect 13614 41560 13708 41600
rect 13748 41560 13757 41600
rect 13998 41560 14092 41600
rect 14132 41560 14141 41600
rect 14382 41560 14476 41600
rect 14516 41560 14525 41600
rect 14659 41560 14668 41600
rect 14708 41560 14860 41600
rect 14900 41560 14909 41600
rect 16099 41560 16108 41600
rect 16148 41560 16157 41600
rect 16579 41560 16588 41600
rect 16628 41560 16684 41600
rect 16724 41560 16733 41600
rect 17347 41560 17356 41600
rect 17396 41560 18796 41600
rect 18836 41560 18845 41600
rect 20039 41560 20048 41600
rect 20088 41560 20130 41600
rect 20170 41560 20212 41600
rect 20252 41560 20294 41600
rect 20334 41560 20376 41600
rect 20416 41560 20425 41600
rect 6028 41516 6068 41560
rect 7459 41559 7517 41560
rect 9292 41516 9332 41560
rect 9475 41559 9533 41560
rect 11203 41559 11261 41560
rect 11779 41516 11837 41517
rect 4099 41476 4108 41516
rect 4148 41476 4492 41516
rect 4532 41476 6068 41516
rect 6115 41476 6124 41516
rect 6164 41476 8524 41516
rect 8564 41476 8573 41516
rect 9292 41476 11360 41516
rect 11694 41476 11788 41516
rect 11828 41476 11837 41516
rect 11884 41516 11924 41560
rect 12547 41559 12605 41560
rect 13411 41559 13469 41560
rect 13699 41559 13757 41560
rect 14083 41559 14141 41560
rect 14467 41559 14525 41560
rect 14851 41559 14909 41560
rect 16108 41516 16148 41560
rect 16675 41559 16733 41560
rect 11884 41476 15380 41516
rect 16108 41476 16492 41516
rect 16532 41476 16541 41516
rect 18307 41476 18316 41516
rect 18356 41476 19756 41516
rect 19796 41476 19805 41516
rect 0 41432 80 41452
rect 11320 41432 11360 41476
rect 11779 41475 11837 41476
rect 0 41392 9388 41432
rect 9428 41392 9437 41432
rect 11320 41392 13804 41432
rect 13844 41392 13853 41432
rect 0 41372 80 41392
rect 15340 41348 15380 41476
rect 18691 41392 18700 41432
rect 18740 41392 19468 41432
rect 19508 41392 19517 41432
rect 2083 41308 2092 41348
rect 2132 41308 4780 41348
rect 4820 41308 4829 41348
rect 6499 41308 6508 41348
rect 6548 41308 8140 41348
rect 8180 41308 8189 41348
rect 8236 41308 11308 41348
rect 11348 41308 11357 41348
rect 15340 41308 19372 41348
rect 19412 41308 19421 41348
rect 2500 41224 7756 41264
rect 7796 41224 8044 41264
rect 8084 41224 8093 41264
rect 1699 41140 1708 41180
rect 1748 41140 1900 41180
rect 1940 41140 1949 41180
rect 0 41096 80 41116
rect 2500 41096 2540 41224
rect 5539 41180 5597 41181
rect 3331 41140 3340 41180
rect 3380 41140 3628 41180
rect 3668 41140 3677 41180
rect 5454 41140 5548 41180
rect 5588 41140 5597 41180
rect 5827 41140 5836 41180
rect 5876 41140 7948 41180
rect 7988 41140 7997 41180
rect 5539 41139 5597 41140
rect 0 41056 2540 41096
rect 3427 41096 3485 41097
rect 4195 41096 4253 41097
rect 4771 41096 4829 41097
rect 8236 41096 8276 41308
rect 13987 41264 14045 41265
rect 9379 41224 9388 41264
rect 9428 41224 13652 41264
rect 10243 41180 10301 41181
rect 11683 41180 11741 41181
rect 13612 41180 13652 41224
rect 13987 41224 13996 41264
rect 14036 41224 19124 41264
rect 13987 41223 14045 41224
rect 19084 41180 19124 41224
rect 9283 41140 9292 41180
rect 9332 41140 9580 41180
rect 9620 41140 9629 41180
rect 10147 41140 10156 41180
rect 10196 41140 10252 41180
rect 10292 41140 10301 41180
rect 11587 41140 11596 41180
rect 11636 41140 11692 41180
rect 11732 41140 11741 41180
rect 13603 41140 13612 41180
rect 13652 41140 13661 41180
rect 16579 41140 16588 41180
rect 16628 41140 17644 41180
rect 17684 41140 17693 41180
rect 18019 41140 18028 41180
rect 18068 41140 18508 41180
rect 18548 41140 18557 41180
rect 19075 41140 19084 41180
rect 19124 41140 19133 41180
rect 10243 41139 10301 41140
rect 11683 41139 11741 41140
rect 3427 41056 3436 41096
rect 3476 41056 3724 41096
rect 3764 41056 3773 41096
rect 4195 41056 4204 41096
rect 4244 41056 4780 41096
rect 4820 41056 8276 41096
rect 8323 41056 8332 41096
rect 8372 41056 16780 41096
rect 16820 41056 16829 41096
rect 0 41036 80 41056
rect 3427 41055 3485 41056
rect 4195 41055 4253 41056
rect 4771 41055 4829 41056
rect 14275 41012 14333 41013
rect 15139 41012 15197 41013
rect 1315 40972 1324 41012
rect 1364 40972 1516 41012
rect 1556 40972 1565 41012
rect 2500 40972 3916 41012
rect 3956 40972 3965 41012
rect 5347 40972 5356 41012
rect 5396 40972 6988 41012
rect 7028 40972 7037 41012
rect 14275 40972 14284 41012
rect 14324 40972 14764 41012
rect 14804 40972 14813 41012
rect 15054 40972 15148 41012
rect 15188 40972 15197 41012
rect 18691 40972 18700 41012
rect 18740 40972 18988 41012
rect 19028 40972 19037 41012
rect 2500 40928 2540 40972
rect 14275 40971 14333 40972
rect 15139 40971 15197 40972
rect 2092 40888 2540 40928
rect 7363 40888 7372 40928
rect 7412 40888 12076 40928
rect 12116 40888 12125 40928
rect 13603 40888 13612 40928
rect 13652 40888 19372 40928
rect 19412 40888 19421 40928
rect 2092 40844 2132 40888
rect 12355 40844 12413 40845
rect 17731 40844 17789 40845
rect 2083 40804 2092 40844
rect 2132 40804 2141 40844
rect 3679 40804 3688 40844
rect 3728 40804 3770 40844
rect 3810 40804 3852 40844
rect 3892 40804 3934 40844
rect 3974 40804 4016 40844
rect 4056 40804 4065 40844
rect 8035 40804 8044 40844
rect 8084 40804 12364 40844
rect 12404 40804 17740 40844
rect 17780 40804 17789 40844
rect 18799 40804 18808 40844
rect 18848 40804 18890 40844
rect 18930 40804 18972 40844
rect 19012 40804 19054 40844
rect 19094 40804 19136 40844
rect 19176 40804 19185 40844
rect 12355 40803 12413 40804
rect 17731 40803 17789 40804
rect 0 40760 80 40780
rect 0 40720 1324 40760
rect 1364 40720 1373 40760
rect 17923 40720 17932 40760
rect 17972 40720 18508 40760
rect 18548 40720 18557 40760
rect 0 40700 80 40720
rect 2275 40676 2333 40677
rect 4771 40676 4829 40677
rect 18691 40676 18749 40677
rect 2190 40636 2284 40676
rect 2324 40636 2333 40676
rect 2851 40636 2860 40676
rect 2900 40636 4780 40676
rect 4820 40636 4829 40676
rect 5443 40636 5452 40676
rect 5492 40636 6508 40676
rect 6548 40636 6557 40676
rect 7171 40636 7180 40676
rect 7220 40636 7948 40676
rect 7988 40636 7997 40676
rect 13219 40636 13228 40676
rect 13268 40636 13804 40676
rect 13844 40636 13853 40676
rect 14371 40636 14380 40676
rect 14420 40636 14429 40676
rect 16387 40636 16396 40676
rect 16436 40636 16972 40676
rect 17012 40636 17021 40676
rect 17539 40636 17548 40676
rect 17588 40636 18124 40676
rect 18164 40636 18173 40676
rect 18691 40636 18700 40676
rect 18740 40636 18892 40676
rect 18932 40636 18941 40676
rect 2275 40635 2333 40636
rect 4771 40635 4829 40636
rect 6307 40592 6365 40593
rect 13507 40592 13565 40593
rect 14380 40592 14420 40636
rect 18691 40635 18749 40636
rect 15811 40592 15869 40593
rect 20515 40592 20573 40593
rect 172 40552 6316 40592
rect 6356 40552 6365 40592
rect 6979 40552 6988 40592
rect 7028 40552 10348 40592
rect 10388 40552 11360 40592
rect 0 40424 80 40444
rect 0 40364 116 40424
rect 76 40340 116 40364
rect 172 40340 212 40552
rect 6307 40551 6365 40552
rect 8611 40508 8669 40509
rect 11320 40508 11360 40552
rect 13507 40552 13516 40592
rect 13556 40552 14420 40592
rect 15726 40552 15820 40592
rect 15860 40552 15869 40592
rect 19555 40552 19564 40592
rect 19604 40552 20524 40592
rect 20564 40552 20573 40592
rect 13507 40551 13565 40552
rect 15811 40551 15869 40552
rect 20515 40551 20573 40552
rect 18307 40508 18365 40509
rect 1507 40468 1516 40508
rect 1556 40468 2284 40508
rect 2324 40468 2996 40508
rect 8131 40468 8140 40508
rect 8180 40468 8620 40508
rect 8660 40468 8669 40508
rect 8995 40468 9004 40508
rect 9044 40468 10732 40508
rect 10772 40468 10781 40508
rect 11320 40468 15188 40508
rect 15235 40468 15244 40508
rect 15284 40468 16012 40508
rect 16052 40468 16061 40508
rect 18307 40468 18316 40508
rect 18356 40468 19948 40508
rect 19988 40468 19997 40508
rect 2956 40425 2996 40468
rect 8611 40467 8669 40468
rect 2947 40424 3005 40425
rect 15148 40424 15188 40468
rect 18307 40467 18365 40468
rect 1795 40384 1804 40424
rect 1844 40384 2188 40424
rect 2228 40384 2237 40424
rect 2947 40384 2956 40424
rect 2996 40384 3005 40424
rect 3523 40384 3532 40424
rect 3572 40384 3820 40424
rect 3860 40384 4492 40424
rect 4532 40384 4541 40424
rect 7651 40384 7660 40424
rect 7700 40384 8908 40424
rect 8948 40384 8957 40424
rect 10051 40384 10060 40424
rect 10100 40384 10924 40424
rect 10964 40384 10973 40424
rect 11683 40384 11692 40424
rect 11732 40384 11741 40424
rect 12259 40384 12268 40424
rect 12308 40384 13420 40424
rect 13460 40384 13469 40424
rect 13795 40384 13804 40424
rect 13844 40384 14380 40424
rect 14420 40384 14429 40424
rect 15148 40384 15628 40424
rect 15668 40384 16108 40424
rect 16148 40384 16157 40424
rect 16204 40384 16780 40424
rect 16820 40384 16829 40424
rect 17923 40384 17932 40424
rect 17972 40384 20524 40424
rect 20564 40384 20573 40424
rect 2947 40383 3005 40384
rect 3235 40340 3293 40341
rect 9187 40340 9245 40341
rect 11692 40340 11732 40384
rect 14380 40340 14420 40384
rect 16204 40340 16244 40384
rect 76 40300 212 40340
rect 1315 40300 1324 40340
rect 1364 40300 1516 40340
rect 1556 40300 1565 40340
rect 1891 40300 1900 40340
rect 1940 40300 2228 40340
rect 3150 40300 3244 40340
rect 3284 40300 3293 40340
rect 5251 40300 5260 40340
rect 5300 40300 5644 40340
rect 5684 40300 5693 40340
rect 7459 40300 7468 40340
rect 7508 40300 7852 40340
rect 7892 40300 7901 40340
rect 9187 40300 9196 40340
rect 9236 40300 11020 40340
rect 11060 40300 11069 40340
rect 11320 40300 11732 40340
rect 11779 40300 11788 40340
rect 11828 40300 11980 40340
rect 12020 40300 12364 40340
rect 12404 40300 12652 40340
rect 12692 40300 12701 40340
rect 14380 40300 15436 40340
rect 15476 40300 16244 40340
rect 16291 40340 16349 40341
rect 18115 40340 18173 40341
rect 16291 40300 16300 40340
rect 16340 40300 16684 40340
rect 16724 40300 16733 40340
rect 17539 40300 17548 40340
rect 17588 40300 18124 40340
rect 18164 40300 18220 40340
rect 18260 40300 18288 40340
rect 2188 40256 2228 40300
rect 3235 40299 3293 40300
rect 9187 40299 9245 40300
rect 3523 40256 3581 40257
rect 2188 40216 3532 40256
rect 3572 40216 3581 40256
rect 5059 40216 5068 40256
rect 5108 40216 8852 40256
rect 8899 40216 8908 40256
rect 8948 40216 9868 40256
rect 9908 40216 9917 40256
rect 3523 40215 3581 40216
rect 2284 40132 8524 40172
rect 8564 40132 8573 40172
rect 0 40088 80 40108
rect 1315 40088 1373 40089
rect 2284 40088 2324 40132
rect 8707 40088 8765 40089
rect 8812 40088 8852 40216
rect 11320 40088 11360 40300
rect 16291 40299 16349 40300
rect 18115 40299 18173 40300
rect 14179 40216 14188 40256
rect 14228 40216 14860 40256
rect 14900 40216 14909 40256
rect 11491 40132 11500 40172
rect 11540 40132 13516 40172
rect 13556 40132 16396 40172
rect 16436 40132 16445 40172
rect 21424 40088 21504 40108
rect 0 40048 1324 40088
rect 1364 40048 2324 40088
rect 4919 40048 4928 40088
rect 4968 40048 5010 40088
rect 5050 40048 5092 40088
rect 5132 40048 5174 40088
rect 5214 40048 5256 40088
rect 5296 40048 5305 40088
rect 7267 40048 7276 40088
rect 7316 40048 7468 40088
rect 7508 40048 7517 40088
rect 8688 40048 8716 40088
rect 8756 40048 10252 40088
rect 10292 40048 11360 40088
rect 12163 40048 12172 40088
rect 12212 40048 12221 40088
rect 12931 40048 12940 40088
rect 12980 40048 14380 40088
rect 14420 40048 14429 40088
rect 20039 40048 20048 40088
rect 20088 40048 20130 40088
rect 20170 40048 20212 40088
rect 20252 40048 20294 40088
rect 20334 40048 20376 40088
rect 20416 40048 20425 40088
rect 20524 40048 21504 40088
rect 0 40028 80 40048
rect 1315 40047 1373 40048
rect 8707 40047 8765 40048
rect 1411 40004 1469 40005
rect 7363 40004 7421 40005
rect 11320 40004 11360 40048
rect 12172 40004 12212 40048
rect 1411 39964 1420 40004
rect 1460 39964 6028 40004
rect 6068 39964 6077 40004
rect 7363 39964 7372 40004
rect 7412 39964 8236 40004
rect 8276 39964 8285 40004
rect 9187 39964 9196 40004
rect 9236 39964 9484 40004
rect 9524 39964 9533 40004
rect 11320 39964 11732 40004
rect 11779 39964 11788 40004
rect 11828 39964 12212 40004
rect 17539 40004 17597 40005
rect 20524 40004 20564 40048
rect 21424 40028 21504 40048
rect 17539 39964 17548 40004
rect 17588 39964 20564 40004
rect 1411 39963 1469 39964
rect 7363 39963 7421 39964
rect 8131 39920 8189 39921
rect 2275 39880 2284 39920
rect 2324 39880 6316 39920
rect 6356 39880 6365 39920
rect 8131 39880 8140 39920
rect 8180 39880 9772 39920
rect 9812 39880 9821 39920
rect 8131 39879 8189 39880
rect 11692 39836 11732 39964
rect 17539 39963 17597 39964
rect 17635 39920 17693 39921
rect 12163 39880 12172 39920
rect 12212 39880 12940 39920
rect 12980 39880 12989 39920
rect 17550 39880 17644 39920
rect 17684 39880 17693 39920
rect 18307 39880 18316 39920
rect 18356 39880 18700 39920
rect 18740 39880 18749 39920
rect 17635 39879 17693 39880
rect 2500 39796 2956 39836
rect 2996 39796 3005 39836
rect 5923 39796 5932 39836
rect 5972 39796 7276 39836
rect 7316 39796 7325 39836
rect 11320 39796 11636 39836
rect 11692 39796 19372 39836
rect 19412 39796 19421 39836
rect 0 39752 80 39772
rect 2500 39752 2540 39796
rect 11320 39752 11360 39796
rect 0 39712 2540 39752
rect 3043 39712 3052 39752
rect 3092 39712 8044 39752
rect 8084 39712 11360 39752
rect 0 39692 80 39712
rect 5059 39668 5117 39669
rect 6787 39668 6845 39669
rect 2563 39628 2572 39668
rect 2612 39628 3956 39668
rect 4003 39628 4012 39668
rect 4052 39628 4300 39668
rect 4340 39628 4349 39668
rect 5059 39628 5068 39668
rect 5108 39628 5932 39668
rect 5972 39628 6412 39668
rect 6452 39628 6461 39668
rect 6702 39628 6796 39668
rect 6836 39628 6845 39668
rect 2755 39584 2813 39585
rect 3811 39584 3869 39585
rect 1315 39544 1324 39584
rect 1364 39544 1516 39584
rect 1556 39544 2764 39584
rect 2804 39544 2813 39584
rect 2755 39543 2813 39544
rect 3628 39544 3820 39584
rect 3860 39544 3869 39584
rect 3628 39500 3668 39544
rect 3811 39543 3869 39544
rect 1123 39460 1132 39500
rect 1172 39460 3668 39500
rect 3715 39460 3724 39500
rect 3764 39460 3773 39500
rect 0 39416 80 39436
rect 2275 39416 2333 39417
rect 3724 39416 3764 39460
rect 0 39376 2092 39416
rect 2132 39376 2284 39416
rect 2324 39376 2333 39416
rect 2563 39376 2572 39416
rect 2612 39376 2860 39416
rect 2900 39376 2909 39416
rect 3427 39376 3436 39416
rect 3476 39376 3764 39416
rect 3916 39416 3956 39628
rect 5059 39627 5117 39628
rect 6787 39627 6845 39628
rect 6595 39584 6653 39585
rect 11203 39584 11261 39585
rect 4579 39544 4588 39584
rect 4628 39544 5260 39584
rect 5300 39544 5309 39584
rect 5635 39544 5644 39584
rect 5684 39544 6604 39584
rect 6644 39544 6653 39584
rect 6883 39544 6892 39584
rect 6932 39544 11212 39584
rect 11252 39544 11261 39584
rect 11596 39584 11636 39796
rect 19843 39752 19901 39753
rect 20611 39752 20669 39753
rect 11683 39712 11692 39752
rect 11732 39712 11980 39752
rect 12020 39712 12029 39752
rect 12739 39712 12748 39752
rect 12788 39712 13036 39752
rect 13076 39712 16012 39752
rect 16052 39712 16061 39752
rect 16291 39712 16300 39752
rect 16340 39712 16972 39752
rect 17012 39712 17021 39752
rect 19758 39712 19852 39752
rect 19892 39712 19901 39752
rect 19843 39711 19901 39712
rect 20140 39712 20620 39752
rect 20660 39712 20669 39752
rect 20140 39668 20180 39712
rect 20611 39711 20669 39712
rect 13795 39628 13804 39668
rect 13844 39628 14572 39668
rect 14612 39628 14621 39668
rect 18307 39628 18316 39668
rect 18356 39628 18796 39668
rect 18836 39628 18845 39668
rect 19075 39628 19084 39668
rect 19124 39628 20180 39668
rect 15715 39584 15773 39585
rect 11596 39544 15724 39584
rect 15764 39544 15773 39584
rect 6595 39543 6653 39544
rect 11203 39543 11261 39544
rect 15715 39543 15773 39544
rect 17923 39584 17981 39585
rect 21424 39584 21504 39604
rect 17923 39544 17932 39584
rect 17972 39544 18220 39584
rect 18260 39544 18269 39584
rect 19843 39544 19852 39584
rect 19892 39544 21504 39584
rect 17923 39543 17981 39544
rect 21424 39524 21504 39544
rect 4003 39500 4061 39501
rect 4387 39500 4445 39501
rect 8899 39500 8957 39501
rect 4003 39460 4012 39500
rect 4052 39460 4396 39500
rect 4436 39460 4445 39500
rect 5443 39460 5452 39500
rect 5492 39460 5684 39500
rect 4003 39459 4061 39460
rect 4387 39459 4445 39460
rect 5644 39416 5684 39460
rect 5932 39460 8908 39500
rect 8948 39460 8957 39500
rect 12931 39460 12940 39500
rect 12980 39460 20044 39500
rect 20084 39460 20093 39500
rect 3916 39376 5588 39416
rect 5635 39376 5644 39416
rect 5684 39376 5693 39416
rect 0 39356 80 39376
rect 2275 39375 2333 39376
rect 5548 39332 5588 39376
rect 5932 39332 5972 39460
rect 8899 39459 8957 39460
rect 8515 39376 8524 39416
rect 8564 39376 19468 39416
rect 19508 39376 19517 39416
rect 3679 39292 3688 39332
rect 3728 39292 3770 39332
rect 3810 39292 3852 39332
rect 3892 39292 3934 39332
rect 3974 39292 4016 39332
rect 4056 39292 4065 39332
rect 5548 39292 5972 39332
rect 6019 39292 6028 39332
rect 6068 39292 11980 39332
rect 12020 39292 12940 39332
rect 12980 39292 12989 39332
rect 14083 39292 14092 39332
rect 14132 39292 14380 39332
rect 14420 39292 14429 39332
rect 15331 39292 15340 39332
rect 15380 39292 16204 39332
rect 16244 39292 16253 39332
rect 18799 39292 18808 39332
rect 18848 39292 18890 39332
rect 18930 39292 18972 39332
rect 19012 39292 19054 39332
rect 19094 39292 19136 39332
rect 19176 39292 19185 39332
rect 67 39248 125 39249
rect 19459 39248 19517 39249
rect 67 39208 76 39248
rect 116 39208 2476 39248
rect 2516 39208 13036 39248
rect 13076 39208 13085 39248
rect 13411 39208 13420 39248
rect 13460 39208 13900 39248
rect 13940 39208 14188 39248
rect 14228 39208 14237 39248
rect 16867 39208 16876 39248
rect 16916 39208 19468 39248
rect 19508 39208 19517 39248
rect 67 39207 125 39208
rect 19459 39207 19517 39208
rect 2179 39164 2237 39165
rect 1987 39124 1996 39164
rect 2036 39124 2188 39164
rect 2228 39124 2237 39164
rect 2179 39123 2237 39124
rect 2500 39124 4108 39164
rect 4148 39124 4157 39164
rect 12259 39124 12268 39164
rect 12308 39124 12460 39164
rect 12500 39124 12509 39164
rect 12835 39124 12844 39164
rect 12884 39124 13132 39164
rect 13172 39124 13181 39164
rect 16195 39124 16204 39164
rect 16244 39124 20180 39164
rect 0 39080 80 39100
rect 2500 39080 2540 39124
rect 8227 39080 8285 39081
rect 11299 39080 11357 39081
rect 20140 39080 20180 39124
rect 21424 39080 21504 39100
rect 0 39040 1132 39080
rect 1172 39040 1181 39080
rect 1507 39040 1516 39080
rect 1556 39040 2540 39080
rect 3619 39040 3628 39080
rect 3668 39040 6316 39080
rect 6356 39040 6365 39080
rect 8227 39040 8236 39080
rect 8276 39040 10444 39080
rect 10484 39040 10493 39080
rect 10627 39040 10636 39080
rect 10676 39040 11116 39080
rect 11156 39040 11308 39080
rect 11348 39040 11357 39080
rect 12547 39040 12556 39080
rect 12596 39040 13804 39080
rect 13844 39040 14668 39080
rect 14708 39040 14717 39080
rect 16387 39040 16396 39080
rect 16436 39040 17164 39080
rect 17204 39040 17548 39080
rect 17588 39040 17597 39080
rect 17731 39040 17740 39080
rect 17780 39040 19412 39080
rect 20140 39040 21504 39080
rect 0 39020 80 39040
rect 8227 39039 8285 39040
rect 11299 39039 11357 39040
rect 4675 38996 4733 38997
rect 4963 38996 5021 38997
rect 6691 38996 6749 38997
rect 1315 38956 1324 38996
rect 1364 38956 1996 38996
rect 2036 38956 2045 38996
rect 2500 38956 4684 38996
rect 4724 38956 4733 38996
rect 4878 38956 4972 38996
rect 5012 38956 5021 38996
rect 6403 38956 6412 38996
rect 6452 38956 6700 38996
rect 6740 38956 6749 38996
rect 0 38744 80 38764
rect 1411 38744 1469 38745
rect 2500 38744 2540 38956
rect 4675 38955 4733 38956
rect 4963 38955 5021 38956
rect 6691 38955 6749 38956
rect 6883 38996 6941 38997
rect 6883 38956 6892 38996
rect 6932 38956 6988 38996
rect 7028 38956 7037 38996
rect 8803 38956 8812 38996
rect 8852 38956 12364 38996
rect 12404 38956 12413 38996
rect 16963 38956 16972 38996
rect 17012 38956 18892 38996
rect 18932 38956 18941 38996
rect 6883 38955 6941 38956
rect 10627 38912 10685 38913
rect 2947 38872 2956 38912
rect 2996 38872 3005 38912
rect 4387 38872 4396 38912
rect 4436 38872 6796 38912
rect 6836 38872 6845 38912
rect 7459 38872 7468 38912
rect 7508 38872 8428 38912
rect 8468 38872 9868 38912
rect 9908 38872 9917 38912
rect 10542 38872 10636 38912
rect 10676 38872 10685 38912
rect 2956 38828 2996 38872
rect 10627 38871 10685 38872
rect 10915 38912 10973 38913
rect 19372 38912 19412 39040
rect 21424 39020 21504 39040
rect 20323 38956 20332 38996
rect 20372 38956 21292 38996
rect 21332 38956 21341 38996
rect 10915 38872 10924 38912
rect 10964 38872 11020 38912
rect 11060 38872 11069 38912
rect 14467 38872 14476 38912
rect 14516 38872 15148 38912
rect 15188 38872 15197 38912
rect 17059 38872 17068 38912
rect 17108 38872 17740 38912
rect 17780 38872 17789 38912
rect 17923 38872 17932 38912
rect 17972 38872 18988 38912
rect 19028 38872 19037 38912
rect 19363 38872 19372 38912
rect 19412 38872 19421 38912
rect 19747 38872 19756 38912
rect 19796 38872 20180 38912
rect 20227 38872 20236 38912
rect 20276 38872 21388 38912
rect 21428 38872 21437 38912
rect 10915 38871 10973 38872
rect 6211 38828 6269 38829
rect 19939 38828 19997 38829
rect 20140 38828 20180 38872
rect 2956 38788 4588 38828
rect 4628 38788 4637 38828
rect 5539 38788 5548 38828
rect 5588 38788 6220 38828
rect 6260 38788 8332 38828
rect 8372 38788 8381 38828
rect 10243 38788 10252 38828
rect 10292 38788 10540 38828
rect 10580 38788 10589 38828
rect 15532 38788 19564 38828
rect 19604 38788 19613 38828
rect 19939 38788 19948 38828
rect 19988 38788 20044 38828
rect 20084 38788 20093 38828
rect 20140 38788 20812 38828
rect 20852 38788 20861 38828
rect 6211 38787 6269 38788
rect 15532 38744 15572 38788
rect 19939 38787 19997 38788
rect 0 38704 1420 38744
rect 1460 38704 1469 38744
rect 1699 38704 1708 38744
rect 1748 38704 2540 38744
rect 3139 38704 3148 38744
rect 3188 38704 3628 38744
rect 3668 38704 3677 38744
rect 5635 38704 5644 38744
rect 5684 38704 6604 38744
rect 6644 38704 6653 38744
rect 6787 38704 6796 38744
rect 6836 38704 7180 38744
rect 7220 38704 15572 38744
rect 17443 38744 17501 38745
rect 18499 38744 18557 38745
rect 17443 38704 17452 38744
rect 17492 38704 18124 38744
rect 18164 38704 18173 38744
rect 18414 38704 18508 38744
rect 18548 38704 18557 38744
rect 19459 38704 19468 38744
rect 19508 38704 20660 38744
rect 0 38684 80 38704
rect 1411 38703 1469 38704
rect 17443 38703 17501 38704
rect 18499 38703 18557 38704
rect 2179 38660 2237 38661
rect 2179 38620 2188 38660
rect 2228 38620 2996 38660
rect 2179 38619 2237 38620
rect 2956 38576 2996 38620
rect 3148 38620 6700 38660
rect 6740 38620 6749 38660
rect 6796 38620 8812 38660
rect 8852 38620 8861 38660
rect 17827 38620 17836 38660
rect 17876 38620 18796 38660
rect 18836 38620 18845 38660
rect 3148 38576 3188 38620
rect 6796 38576 6836 38620
rect 19939 38576 19997 38577
rect 20620 38576 20660 38704
rect 21424 38576 21504 38596
rect 2179 38536 2188 38576
rect 2228 38536 2476 38576
rect 2516 38536 2525 38576
rect 2956 38536 3188 38576
rect 4919 38536 4928 38576
rect 4968 38536 5010 38576
rect 5050 38536 5092 38576
rect 5132 38536 5174 38576
rect 5214 38536 5256 38576
rect 5296 38536 5305 38576
rect 5635 38536 5644 38576
rect 5684 38536 6836 38576
rect 9859 38536 9868 38576
rect 9908 38536 10060 38576
rect 10100 38536 11500 38576
rect 11540 38536 11884 38576
rect 11924 38536 11933 38576
rect 17539 38536 17548 38576
rect 17588 38536 17932 38576
rect 17972 38536 18124 38576
rect 18164 38536 18173 38576
rect 19276 38536 19948 38576
rect 19988 38536 19997 38576
rect 20039 38536 20048 38576
rect 20088 38536 20130 38576
rect 20170 38536 20212 38576
rect 20252 38536 20294 38576
rect 20334 38536 20376 38576
rect 20416 38536 20425 38576
rect 20620 38536 21504 38576
rect 19276 38492 19316 38536
rect 19939 38535 19997 38536
rect 21424 38516 21504 38536
rect 19459 38492 19517 38493
rect 1315 38452 1324 38492
rect 1364 38452 1612 38492
rect 1652 38452 15628 38492
rect 15668 38452 15677 38492
rect 16684 38452 19316 38492
rect 19374 38452 19468 38492
rect 19508 38452 19517 38492
rect 0 38408 80 38428
rect 7939 38408 7997 38409
rect 16684 38408 16724 38452
rect 19459 38451 19517 38452
rect 17635 38408 17693 38409
rect 20419 38408 20477 38409
rect 0 38368 1708 38408
rect 1748 38368 1757 38408
rect 2851 38368 2860 38408
rect 2900 38368 3628 38408
rect 3668 38368 6796 38408
rect 6836 38368 6845 38408
rect 7939 38368 7948 38408
rect 7988 38368 8044 38408
rect 8084 38368 8524 38408
rect 8564 38368 8573 38408
rect 10627 38368 10636 38408
rect 10676 38368 16684 38408
rect 16724 38368 16733 38408
rect 17635 38368 17644 38408
rect 17684 38368 20428 38408
rect 20468 38368 20477 38408
rect 0 38348 80 38368
rect 7939 38367 7997 38368
rect 17635 38367 17693 38368
rect 20419 38367 20477 38368
rect 2083 38284 2092 38324
rect 2132 38284 5876 38324
rect 6691 38284 6700 38324
rect 6740 38284 17932 38324
rect 17972 38284 17981 38324
rect 18307 38284 18316 38324
rect 18356 38284 18796 38324
rect 18836 38284 18845 38324
rect 2467 38200 2476 38240
rect 2516 38200 4396 38240
rect 4436 38200 4445 38240
rect 2659 38156 2717 38157
rect 4387 38156 4445 38157
rect 2574 38116 2668 38156
rect 2708 38116 2717 38156
rect 2947 38116 2956 38156
rect 2996 38116 4108 38156
rect 4148 38116 4157 38156
rect 4387 38116 4396 38156
rect 4436 38116 5644 38156
rect 5684 38116 5693 38156
rect 2659 38115 2717 38116
rect 4387 38115 4445 38116
rect 0 38072 80 38092
rect 0 38032 4300 38072
rect 4340 38032 4492 38072
rect 4532 38032 4541 38072
rect 0 38012 80 38032
rect 3811 37988 3869 37989
rect 3619 37948 3628 37988
rect 3668 37948 3677 37988
rect 3726 37948 3820 37988
rect 3860 37948 3869 37988
rect 5836 37988 5876 38284
rect 11587 38240 11645 38241
rect 16684 38240 16724 38284
rect 7555 38200 7564 38240
rect 7604 38200 8620 38240
rect 8660 38200 8669 38240
rect 10723 38200 10732 38240
rect 10772 38200 11596 38240
rect 11636 38200 11645 38240
rect 15523 38200 15532 38240
rect 15572 38200 15820 38240
rect 15860 38200 15869 38240
rect 16675 38200 16684 38240
rect 16724 38200 16733 38240
rect 17251 38200 17260 38240
rect 17300 38200 19756 38240
rect 19796 38200 19805 38240
rect 11587 38199 11645 38200
rect 5923 38156 5981 38157
rect 17155 38156 17213 38157
rect 5923 38116 5932 38156
rect 5972 38116 7468 38156
rect 7508 38116 7517 38156
rect 9091 38116 9100 38156
rect 9140 38116 12556 38156
rect 12596 38116 12605 38156
rect 13027 38116 13036 38156
rect 13076 38116 13612 38156
rect 13652 38116 13661 38156
rect 17070 38116 17164 38156
rect 17204 38116 17213 38156
rect 5923 38115 5981 38116
rect 17155 38115 17213 38116
rect 17347 38156 17405 38157
rect 19843 38156 19901 38157
rect 17347 38116 17356 38156
rect 17396 38116 19852 38156
rect 19892 38116 19901 38156
rect 17347 38115 17405 38116
rect 19843 38115 19901 38116
rect 6019 38072 6077 38073
rect 18691 38072 18749 38073
rect 20515 38072 20573 38073
rect 21424 38072 21504 38092
rect 5934 38032 6028 38072
rect 6068 38032 6077 38072
rect 12355 38032 12364 38072
rect 12404 38032 14612 38072
rect 16579 38032 16588 38072
rect 16628 38032 17644 38072
rect 17684 38032 17836 38072
rect 17876 38032 17885 38072
rect 18691 38032 18700 38072
rect 18740 38032 19180 38072
rect 19220 38032 19229 38072
rect 20515 38032 20524 38072
rect 20564 38032 21504 38072
rect 6019 38031 6077 38032
rect 14572 37988 14612 38032
rect 18691 38031 18749 38032
rect 20515 38031 20573 38032
rect 21424 38012 21504 38032
rect 17347 37988 17405 37989
rect 19267 37988 19325 37989
rect 5836 37948 10540 37988
rect 10580 37948 10589 37988
rect 14467 37948 14476 37988
rect 14516 37948 14525 37988
rect 14572 37948 16876 37988
rect 16916 37948 16925 37988
rect 17347 37948 17356 37988
rect 17396 37948 17452 37988
rect 17492 37948 17501 37988
rect 19182 37948 19276 37988
rect 19316 37948 19325 37988
rect 3628 37904 3668 37948
rect 3811 37947 3869 37948
rect 14476 37904 14516 37948
rect 17347 37947 17405 37948
rect 19267 37947 19325 37948
rect 17251 37904 17309 37905
rect 17539 37904 17597 37905
rect 3244 37864 3668 37904
rect 6499 37864 6508 37904
rect 6548 37864 14516 37904
rect 14572 37864 15148 37904
rect 15188 37864 15197 37904
rect 15619 37864 15628 37904
rect 15668 37864 16204 37904
rect 16244 37864 17260 37904
rect 17300 37864 17309 37904
rect 2467 37820 2525 37821
rect 2659 37820 2717 37821
rect 3244 37820 3284 37864
rect 3427 37820 3485 37821
rect 13987 37820 14045 37821
rect 2448 37780 2476 37820
rect 2516 37780 2612 37820
rect 2467 37779 2525 37780
rect 0 37736 80 37756
rect 2572 37736 2612 37780
rect 2659 37780 2668 37820
rect 2708 37780 2764 37820
rect 2804 37780 2813 37820
rect 3235 37780 3244 37820
rect 3284 37780 3293 37820
rect 3342 37780 3436 37820
rect 3476 37780 3485 37820
rect 3679 37780 3688 37820
rect 3728 37780 3770 37820
rect 3810 37780 3852 37820
rect 3892 37780 3934 37820
rect 3974 37780 4016 37820
rect 4056 37780 4065 37820
rect 5923 37780 5932 37820
rect 5972 37780 7660 37820
rect 7700 37780 8428 37820
rect 8468 37780 8477 37820
rect 12739 37780 12748 37820
rect 12788 37780 13420 37820
rect 13460 37780 13996 37820
rect 14036 37780 14045 37820
rect 2659 37779 2717 37780
rect 3427 37779 3485 37780
rect 13987 37779 14045 37780
rect 14380 37736 14420 37864
rect 14572 37820 14612 37864
rect 17251 37863 17309 37864
rect 17452 37864 17548 37904
rect 17588 37864 17597 37904
rect 17452 37820 17492 37864
rect 17539 37863 17597 37864
rect 14467 37780 14476 37820
rect 14516 37780 14612 37820
rect 15012 37780 15052 37820
rect 15092 37780 15101 37820
rect 17443 37780 17452 37820
rect 17492 37780 17501 37820
rect 18799 37780 18808 37820
rect 18848 37780 18890 37820
rect 18930 37780 18972 37820
rect 19012 37780 19054 37820
rect 19094 37780 19136 37820
rect 19176 37780 19185 37820
rect 0 37696 1268 37736
rect 1603 37696 1612 37736
rect 1652 37696 2476 37736
rect 2516 37696 2525 37736
rect 2572 37696 3532 37736
rect 3572 37696 3581 37736
rect 8035 37696 8044 37736
rect 8084 37696 11596 37736
rect 11636 37696 11645 37736
rect 14275 37696 14284 37736
rect 14324 37696 14420 37736
rect 15052 37736 15092 37780
rect 15052 37696 16684 37736
rect 16724 37696 16733 37736
rect 17155 37696 17164 37736
rect 17204 37696 17548 37736
rect 17588 37696 17597 37736
rect 0 37676 80 37696
rect 1228 37568 1268 37696
rect 1987 37612 1996 37652
rect 2036 37612 2764 37652
rect 2804 37612 2813 37652
rect 3811 37612 3820 37652
rect 3860 37612 7756 37652
rect 7796 37612 7805 37652
rect 16003 37612 16012 37652
rect 16052 37612 19180 37652
rect 19220 37612 19229 37652
rect 2467 37568 2525 37569
rect 4579 37568 4637 37569
rect 11779 37568 11837 37569
rect 18691 37568 18749 37569
rect 21424 37568 21504 37588
rect 1228 37528 2476 37568
rect 2516 37528 2525 37568
rect 4387 37528 4396 37568
rect 4436 37528 4588 37568
rect 4628 37528 4637 37568
rect 6115 37528 6124 37568
rect 6164 37528 11788 37568
rect 11828 37528 11837 37568
rect 16387 37528 16396 37568
rect 16436 37528 18700 37568
rect 18740 37528 18749 37568
rect 20515 37528 20524 37568
rect 20564 37528 21504 37568
rect 2467 37527 2525 37528
rect 4579 37527 4637 37528
rect 11779 37527 11837 37528
rect 18691 37527 18749 37528
rect 21424 37508 21504 37528
rect 2500 37444 4780 37484
rect 4820 37444 8044 37484
rect 8084 37444 8093 37484
rect 8323 37444 8332 37484
rect 8372 37444 9004 37484
rect 9044 37444 9053 37484
rect 19555 37444 19564 37484
rect 19604 37444 20044 37484
rect 20084 37444 20093 37484
rect 0 37400 80 37420
rect 2500 37400 2540 37444
rect 5539 37400 5597 37401
rect 0 37360 2540 37400
rect 3331 37360 3340 37400
rect 3380 37360 3389 37400
rect 5454 37360 5548 37400
rect 5588 37360 5597 37400
rect 7843 37360 7852 37400
rect 7892 37360 8428 37400
rect 8468 37360 8477 37400
rect 13891 37360 13900 37400
rect 13940 37360 14188 37400
rect 14228 37360 14237 37400
rect 16579 37360 16588 37400
rect 16628 37360 20236 37400
rect 20276 37360 20285 37400
rect 0 37340 80 37360
rect 3340 37316 3380 37360
rect 5539 37359 5597 37360
rect 10819 37316 10877 37317
rect 3340 37276 6796 37316
rect 6836 37276 6845 37316
rect 10819 37276 10828 37316
rect 10868 37276 10924 37316
rect 10964 37276 10973 37316
rect 16099 37276 16108 37316
rect 16148 37276 17164 37316
rect 17204 37276 17452 37316
rect 17492 37276 18700 37316
rect 18740 37276 18749 37316
rect 10819 37275 10877 37276
rect 4771 37232 4829 37233
rect 5635 37232 5693 37233
rect 20899 37232 20957 37233
rect 4675 37192 4684 37232
rect 4724 37192 4780 37232
rect 4820 37192 4829 37232
rect 5155 37192 5164 37232
rect 5204 37192 5644 37232
rect 5684 37192 5693 37232
rect 7459 37192 7468 37232
rect 7508 37192 9100 37232
rect 9140 37192 9149 37232
rect 15811 37192 15820 37232
rect 15860 37192 17356 37232
rect 17396 37192 17405 37232
rect 18307 37192 18316 37232
rect 18356 37192 18508 37232
rect 18548 37192 18557 37232
rect 19651 37192 19660 37232
rect 19700 37192 20908 37232
rect 20948 37192 20957 37232
rect 4771 37191 4829 37192
rect 5635 37191 5693 37192
rect 20899 37191 20957 37192
rect 5827 37148 5885 37149
rect 1795 37108 1804 37148
rect 1844 37108 4108 37148
rect 4148 37108 4157 37148
rect 4291 37108 4300 37148
rect 4340 37108 4588 37148
rect 4628 37108 5588 37148
rect 5635 37108 5644 37148
rect 5684 37108 5836 37148
rect 5876 37108 5885 37148
rect 19939 37108 19948 37148
rect 19988 37108 20852 37148
rect 0 37064 80 37084
rect 5548 37064 5588 37108
rect 5827 37107 5885 37108
rect 8995 37064 9053 37065
rect 20812 37064 20852 37108
rect 21424 37064 21504 37084
rect 0 37024 1132 37064
rect 1172 37024 1181 37064
rect 1987 37024 1996 37064
rect 2036 37024 4204 37064
rect 4244 37024 4253 37064
rect 4919 37024 4928 37064
rect 4968 37024 5010 37064
rect 5050 37024 5092 37064
rect 5132 37024 5174 37064
rect 5214 37024 5256 37064
rect 5296 37024 5305 37064
rect 5453 37024 5548 37064
rect 5588 37024 5932 37064
rect 5972 37024 5981 37064
rect 7852 37024 9004 37064
rect 9044 37024 9053 37064
rect 17827 37024 17836 37064
rect 17876 37024 18412 37064
rect 18452 37024 18461 37064
rect 20039 37024 20048 37064
rect 20088 37024 20130 37064
rect 20170 37024 20212 37064
rect 20252 37024 20294 37064
rect 20334 37024 20376 37064
rect 20416 37024 20425 37064
rect 20812 37024 21504 37064
rect 0 37004 80 37024
rect 7852 36980 7892 37024
rect 8995 37023 9053 37024
rect 21424 37004 21504 37024
rect 10723 36980 10781 36981
rect 17827 36980 17885 36981
rect 2371 36940 2380 36980
rect 2420 36940 7892 36980
rect 7939 36940 7948 36980
rect 7988 36940 10732 36980
rect 10772 36940 10781 36980
rect 12067 36940 12076 36980
rect 12116 36940 14956 36980
rect 14996 36940 16396 36980
rect 16436 36940 16445 36980
rect 17731 36940 17740 36980
rect 17780 36940 17836 36980
rect 17876 36940 17885 36980
rect 10723 36939 10781 36940
rect 17827 36939 17885 36940
rect 2500 36856 6508 36896
rect 6548 36856 6796 36896
rect 6836 36856 6845 36896
rect 7363 36856 7372 36896
rect 7412 36856 8620 36896
rect 8660 36856 8669 36896
rect 9475 36856 9484 36896
rect 9524 36856 18892 36896
rect 18932 36856 19564 36896
rect 19604 36856 19613 36896
rect 0 36728 80 36748
rect 2500 36728 2540 36856
rect 16483 36812 16541 36813
rect 3052 36772 15148 36812
rect 15188 36772 16492 36812
rect 16532 36772 16541 36812
rect 3052 36728 3092 36772
rect 16483 36771 16541 36772
rect 17452 36772 19468 36812
rect 19508 36772 19756 36812
rect 19796 36772 19805 36812
rect 7171 36728 7229 36729
rect 17251 36728 17309 36729
rect 17452 36728 17492 36772
rect 17731 36728 17789 36729
rect 0 36688 2540 36728
rect 3043 36688 3052 36728
rect 3092 36688 3101 36728
rect 6499 36688 6508 36728
rect 6548 36688 7180 36728
rect 7220 36688 7229 36728
rect 7651 36688 7660 36728
rect 7700 36688 8908 36728
rect 8948 36688 10156 36728
rect 10196 36688 10205 36728
rect 10723 36688 10732 36728
rect 10772 36688 12076 36728
rect 12116 36688 12125 36728
rect 12451 36688 12460 36728
rect 12500 36688 17260 36728
rect 17300 36688 17309 36728
rect 17443 36688 17452 36728
rect 17492 36688 17501 36728
rect 17731 36688 17740 36728
rect 17780 36688 19852 36728
rect 19892 36688 19901 36728
rect 0 36668 80 36688
rect 7171 36687 7229 36688
rect 17251 36687 17309 36688
rect 17731 36687 17789 36688
rect 7075 36644 7133 36645
rect 10435 36644 10493 36645
rect 2755 36604 2764 36644
rect 2804 36604 4340 36644
rect 6883 36604 6892 36644
rect 6932 36604 7084 36644
rect 7124 36604 7133 36644
rect 1315 36560 1373 36561
rect 1795 36560 1853 36561
rect 1200 36520 1228 36560
rect 1268 36520 1324 36560
rect 1364 36520 1804 36560
rect 1844 36520 1853 36560
rect 2083 36520 2092 36560
rect 2132 36520 4204 36560
rect 4244 36520 4253 36560
rect 1315 36519 1373 36520
rect 1795 36519 1853 36520
rect 4300 36476 4340 36604
rect 7075 36603 7133 36604
rect 7372 36604 9484 36644
rect 9524 36604 9533 36644
rect 10339 36604 10348 36644
rect 10388 36604 10444 36644
rect 10484 36604 10493 36644
rect 11779 36604 11788 36644
rect 11828 36604 16012 36644
rect 16052 36604 16061 36644
rect 16579 36604 16588 36644
rect 16628 36604 17356 36644
rect 17396 36604 17405 36644
rect 17644 36604 19660 36644
rect 19700 36604 19709 36644
rect 4675 36560 4733 36561
rect 7372 36560 7412 36604
rect 10435 36603 10493 36604
rect 17644 36560 17684 36604
rect 21424 36560 21504 36580
rect 4675 36520 4684 36560
rect 4724 36520 7412 36560
rect 7459 36520 7468 36560
rect 7508 36520 11116 36560
rect 11156 36520 11404 36560
rect 11444 36520 11453 36560
rect 15811 36520 15820 36560
rect 15860 36520 16396 36560
rect 16436 36520 16445 36560
rect 17155 36520 17164 36560
rect 17204 36520 17588 36560
rect 17635 36520 17644 36560
rect 17684 36520 17693 36560
rect 17740 36520 21504 36560
rect 4675 36519 4733 36520
rect 17548 36476 17588 36520
rect 17740 36476 17780 36520
rect 21424 36500 21504 36520
rect 4300 36436 9004 36476
rect 9044 36436 9053 36476
rect 9379 36436 9388 36476
rect 9428 36436 16492 36476
rect 16532 36436 16972 36476
rect 17012 36436 17021 36476
rect 17548 36436 17780 36476
rect 0 36392 80 36412
rect 12643 36392 12701 36393
rect 0 36352 7564 36392
rect 7604 36352 12652 36392
rect 12692 36352 13036 36392
rect 13076 36352 13085 36392
rect 17059 36352 17068 36392
rect 17108 36352 19948 36392
rect 19988 36352 19997 36392
rect 0 36332 80 36352
rect 12643 36351 12701 36352
rect 19363 36308 19421 36309
rect 2083 36268 2092 36308
rect 2132 36268 2476 36308
rect 2516 36268 2525 36308
rect 3679 36268 3688 36308
rect 3728 36268 3770 36308
rect 3810 36268 3852 36308
rect 3892 36268 3934 36308
rect 3974 36268 4016 36308
rect 4056 36268 4065 36308
rect 5443 36268 5452 36308
rect 5492 36268 10636 36308
rect 10676 36268 10685 36308
rect 18799 36268 18808 36308
rect 18848 36268 18890 36308
rect 18930 36268 18972 36308
rect 19012 36268 19054 36308
rect 19094 36268 19136 36308
rect 19176 36268 19185 36308
rect 19278 36268 19372 36308
rect 19412 36268 19421 36308
rect 19363 36267 19421 36268
rect 9379 36224 9437 36225
rect 17251 36224 17309 36225
rect 1123 36184 1132 36224
rect 1172 36184 6796 36224
rect 6836 36184 6845 36224
rect 9187 36184 9196 36224
rect 9236 36184 9388 36224
rect 9428 36184 9437 36224
rect 10051 36184 10060 36224
rect 10100 36184 10348 36224
rect 10388 36184 10397 36224
rect 17251 36184 17260 36224
rect 17300 36184 18068 36224
rect 18211 36184 18220 36224
rect 18260 36184 20716 36224
rect 20756 36184 20765 36224
rect 9196 36140 9236 36184
rect 9379 36183 9437 36184
rect 17251 36183 17309 36184
rect 18028 36140 18068 36184
rect 1603 36100 1612 36140
rect 1652 36100 2188 36140
rect 2228 36100 2237 36140
rect 4963 36100 4972 36140
rect 5012 36100 9236 36140
rect 10915 36100 10924 36140
rect 10964 36100 11308 36140
rect 11348 36100 11357 36140
rect 16867 36100 16876 36140
rect 16916 36100 17356 36140
rect 17396 36100 17405 36140
rect 18019 36100 18028 36140
rect 18068 36100 20044 36140
rect 20084 36100 20093 36140
rect 0 36056 80 36076
rect 6307 36056 6365 36057
rect 21424 36056 21504 36076
rect 0 36016 4300 36056
rect 4340 36016 4349 36056
rect 6307 36016 6316 36056
rect 6356 36016 9388 36056
rect 9428 36016 9437 36056
rect 15331 36016 15340 36056
rect 15380 36016 19180 36056
rect 19220 36016 19229 36056
rect 20803 36016 20812 36056
rect 20852 36016 21504 36056
rect 0 35996 80 36016
rect 6307 36015 6365 36016
rect 21424 35996 21504 36016
rect 6595 35932 6604 35972
rect 6644 35932 7756 35972
rect 7796 35932 7805 35972
rect 4867 35888 4925 35889
rect 19363 35888 19421 35889
rect 1987 35848 1996 35888
rect 2036 35848 2540 35888
rect 4782 35848 4876 35888
rect 4916 35848 4925 35888
rect 6787 35848 6796 35888
rect 6836 35848 9580 35888
rect 9620 35848 9629 35888
rect 11779 35848 11788 35888
rect 11828 35848 15916 35888
rect 15956 35848 17836 35888
rect 17876 35848 17885 35888
rect 19363 35848 19372 35888
rect 19412 35848 19852 35888
rect 19892 35848 19901 35888
rect 2500 35804 2540 35848
rect 4867 35847 4925 35848
rect 19363 35847 19421 35848
rect 2500 35764 9292 35804
rect 9332 35764 9341 35804
rect 10147 35764 10156 35804
rect 10196 35764 11348 35804
rect 11395 35764 11404 35804
rect 11444 35764 15436 35804
rect 15476 35764 15485 35804
rect 16771 35764 16780 35804
rect 16820 35764 16829 35804
rect 0 35720 80 35740
rect 4003 35720 4061 35721
rect 9571 35720 9629 35721
rect 11308 35720 11348 35764
rect 13027 35720 13085 35721
rect 0 35680 3148 35720
rect 3188 35680 3197 35720
rect 3918 35680 4012 35720
rect 4052 35680 4492 35720
rect 4532 35680 4541 35720
rect 5539 35680 5548 35720
rect 5588 35680 8044 35720
rect 8084 35680 8093 35720
rect 8995 35680 9004 35720
rect 9044 35680 9580 35720
rect 9620 35680 9629 35720
rect 10243 35680 10252 35720
rect 10292 35680 10732 35720
rect 10772 35680 10781 35720
rect 11299 35680 11308 35720
rect 11348 35680 11357 35720
rect 12355 35680 12364 35720
rect 12404 35680 12556 35720
rect 12596 35680 12605 35720
rect 12942 35680 13036 35720
rect 13076 35680 13085 35720
rect 0 35660 80 35680
rect 4003 35679 4061 35680
rect 9571 35679 9629 35680
rect 13027 35679 13085 35680
rect 16780 35636 16820 35764
rect 17347 35720 17405 35721
rect 16867 35680 16876 35720
rect 16916 35680 17356 35720
rect 17396 35680 17405 35720
rect 20131 35680 20140 35720
rect 20180 35680 20189 35720
rect 17347 35679 17405 35680
rect 20140 35636 20180 35680
rect 1891 35596 1900 35636
rect 1940 35596 2476 35636
rect 2516 35596 6932 35636
rect 9283 35596 9292 35636
rect 9332 35596 10060 35636
rect 10100 35596 10109 35636
rect 10819 35596 10828 35636
rect 10868 35596 11212 35636
rect 11252 35596 11261 35636
rect 12163 35596 12172 35636
rect 12212 35596 15820 35636
rect 15860 35596 18508 35636
rect 18548 35596 18557 35636
rect 19948 35596 20180 35636
rect 2083 35512 2092 35552
rect 2132 35512 4492 35552
rect 4532 35512 4541 35552
rect 4919 35512 4928 35552
rect 4968 35512 5010 35552
rect 5050 35512 5092 35552
rect 5132 35512 5174 35552
rect 5214 35512 5256 35552
rect 5296 35512 5305 35552
rect 6892 35468 6932 35596
rect 9571 35512 9580 35552
rect 9620 35512 12844 35552
rect 12884 35512 12893 35552
rect 14947 35512 14956 35552
rect 14996 35512 16684 35552
rect 16724 35512 16733 35552
rect 1411 35428 1420 35468
rect 1460 35428 6700 35468
rect 6740 35428 6749 35468
rect 6892 35428 11692 35468
rect 11732 35428 12556 35468
rect 12596 35428 12605 35468
rect 15427 35428 15436 35468
rect 15476 35428 15820 35468
rect 15860 35428 15869 35468
rect 0 35384 80 35404
rect 4099 35384 4157 35385
rect 19363 35384 19421 35385
rect 0 35344 4108 35384
rect 4148 35344 4157 35384
rect 0 35324 80 35344
rect 4099 35343 4157 35344
rect 7564 35344 8428 35384
rect 8468 35344 8477 35384
rect 8803 35344 8812 35384
rect 8852 35344 10004 35384
rect 10051 35344 10060 35384
rect 10100 35344 17068 35384
rect 17108 35344 17117 35384
rect 18988 35344 19372 35384
rect 19412 35344 19421 35384
rect 19948 35384 19988 35596
rect 20899 35552 20957 35553
rect 21424 35552 21504 35572
rect 20039 35512 20048 35552
rect 20088 35512 20130 35552
rect 20170 35512 20212 35552
rect 20252 35512 20294 35552
rect 20334 35512 20376 35552
rect 20416 35512 20425 35552
rect 20899 35512 20908 35552
rect 20948 35512 21504 35552
rect 20899 35511 20957 35512
rect 21424 35492 21504 35512
rect 19948 35344 20140 35384
rect 20180 35344 20189 35384
rect 1411 35260 1420 35300
rect 1460 35260 1900 35300
rect 1940 35260 1949 35300
rect 3139 35260 3148 35300
rect 3188 35260 3436 35300
rect 3476 35260 3485 35300
rect 3619 35260 3628 35300
rect 3668 35260 4012 35300
rect 4052 35260 4061 35300
rect 4387 35260 4396 35300
rect 4436 35260 4684 35300
rect 4724 35260 4733 35300
rect 6403 35260 6412 35300
rect 6452 35260 7468 35300
rect 7508 35260 7517 35300
rect 2947 35176 2956 35216
rect 2996 35176 6124 35216
rect 6164 35176 6173 35216
rect 2500 35092 3532 35132
rect 3572 35092 3581 35132
rect 5347 35092 5356 35132
rect 5396 35092 6028 35132
rect 6068 35092 6077 35132
rect 0 35048 80 35068
rect 2500 35048 2540 35092
rect 7459 35048 7517 35049
rect 0 35008 2540 35048
rect 3043 35008 3052 35048
rect 3092 35008 3820 35048
rect 3860 35008 3869 35048
rect 6499 35008 6508 35048
rect 6548 35008 6988 35048
rect 7028 35008 7468 35048
rect 7508 35008 7517 35048
rect 0 34988 80 35008
rect 7459 35007 7517 35008
rect 7564 34964 7604 35344
rect 9964 35300 10004 35344
rect 10051 35300 10109 35301
rect 8035 35260 8044 35300
rect 8084 35260 9868 35300
rect 9908 35260 9917 35300
rect 9964 35260 10060 35300
rect 10100 35260 10109 35300
rect 10051 35259 10109 35260
rect 10723 35300 10781 35301
rect 18988 35300 19028 35344
rect 19363 35343 19421 35344
rect 10723 35260 10732 35300
rect 10772 35260 10828 35300
rect 10868 35260 10877 35300
rect 16483 35260 16492 35300
rect 16532 35260 19028 35300
rect 19651 35260 19660 35300
rect 19700 35260 20044 35300
rect 20084 35260 20093 35300
rect 10723 35259 10781 35260
rect 8803 35216 8861 35217
rect 9091 35216 9149 35217
rect 7651 35176 7660 35216
rect 7700 35176 7948 35216
rect 7988 35176 7997 35216
rect 8718 35176 8812 35216
rect 8852 35176 9100 35216
rect 9140 35176 9149 35216
rect 10051 35176 10060 35216
rect 10100 35176 10252 35216
rect 10292 35176 10301 35216
rect 11107 35176 11116 35216
rect 11156 35176 11500 35216
rect 11540 35176 11549 35216
rect 13027 35176 13036 35216
rect 13076 35176 13708 35216
rect 13748 35176 13757 35216
rect 18019 35176 18028 35216
rect 18068 35176 19948 35216
rect 19988 35176 19997 35216
rect 8803 35175 8861 35176
rect 9091 35175 9149 35176
rect 17827 35132 17885 35133
rect 19756 35132 19796 35176
rect 7747 35092 7756 35132
rect 7796 35092 9100 35132
rect 9140 35092 9149 35132
rect 11320 35092 11404 35132
rect 11444 35092 11453 35132
rect 13123 35092 13132 35132
rect 13172 35092 14956 35132
rect 14996 35092 15005 35132
rect 15907 35092 15916 35132
rect 15956 35092 16588 35132
rect 16628 35092 16637 35132
rect 17539 35092 17548 35132
rect 17588 35092 17836 35132
rect 17876 35092 19084 35132
rect 19124 35092 19133 35132
rect 19747 35092 19756 35132
rect 19796 35092 19836 35132
rect 11320 35048 11360 35092
rect 17827 35091 17885 35092
rect 18691 35048 18749 35049
rect 21424 35048 21504 35068
rect 8035 35008 8044 35048
rect 8084 35008 9388 35048
rect 9428 35008 11360 35048
rect 17635 35008 17644 35048
rect 17684 35008 18700 35048
rect 18740 35008 18749 35048
rect 20035 35008 20044 35048
rect 20084 35008 20236 35048
rect 20276 35008 20285 35048
rect 21283 35008 21292 35048
rect 21332 35008 21504 35048
rect 18691 35007 18749 35008
rect 21424 34988 21504 35008
rect 8899 34964 8957 34965
rect 9667 34964 9725 34965
rect 3427 34924 3436 34964
rect 3476 34924 7660 34964
rect 7700 34924 7728 34964
rect 8515 34924 8524 34964
rect 8564 34924 8716 34964
rect 8756 34924 8765 34964
rect 8899 34924 8908 34964
rect 8948 34924 9676 34964
rect 9716 34924 9725 34964
rect 9955 34924 9964 34964
rect 10004 34924 10348 34964
rect 10388 34924 10397 34964
rect 10915 34924 10924 34964
rect 10964 34924 11308 34964
rect 11348 34924 11357 34964
rect 8899 34923 8957 34924
rect 9667 34923 9725 34924
rect 17155 34880 17213 34881
rect 2500 34840 12748 34880
rect 12788 34840 12797 34880
rect 14284 34840 17164 34880
rect 17204 34840 18604 34880
rect 18644 34840 18653 34880
rect 0 34712 80 34732
rect 2500 34712 2540 34840
rect 3331 34796 3389 34797
rect 9859 34796 9917 34797
rect 14284 34796 14324 34840
rect 17155 34839 17213 34840
rect 3246 34756 3340 34796
rect 3380 34756 3389 34796
rect 3679 34756 3688 34796
rect 3728 34756 3770 34796
rect 3810 34756 3852 34796
rect 3892 34756 3934 34796
rect 3974 34756 4016 34796
rect 4056 34756 4065 34796
rect 6019 34756 6028 34796
rect 6068 34756 9676 34796
rect 9716 34756 9725 34796
rect 9859 34756 9868 34796
rect 9908 34756 14324 34796
rect 14371 34756 14380 34796
rect 14420 34756 14860 34796
rect 14900 34756 14909 34796
rect 18799 34756 18808 34796
rect 18848 34756 18890 34796
rect 18930 34756 18972 34796
rect 19012 34756 19054 34796
rect 19094 34756 19136 34796
rect 19176 34756 19185 34796
rect 3331 34755 3389 34756
rect 9859 34755 9917 34756
rect 9283 34712 9341 34713
rect 0 34672 212 34712
rect 1507 34672 1516 34712
rect 1556 34672 2540 34712
rect 7651 34672 7660 34712
rect 7700 34672 9292 34712
rect 9332 34672 9341 34712
rect 9571 34672 9580 34712
rect 9620 34672 9964 34712
rect 10004 34672 10013 34712
rect 11320 34672 15244 34712
rect 15284 34672 15293 34712
rect 19267 34672 19276 34712
rect 19316 34672 19468 34712
rect 19508 34672 19517 34712
rect 0 34652 80 34672
rect 172 34628 212 34672
rect 9283 34671 9341 34672
rect 9955 34628 10013 34629
rect 172 34588 1940 34628
rect 7171 34588 7180 34628
rect 7220 34588 7756 34628
rect 7796 34588 7805 34628
rect 8131 34588 8140 34628
rect 8180 34588 9772 34628
rect 9812 34588 9964 34628
rect 10004 34588 10013 34628
rect 1900 34460 1940 34588
rect 9955 34587 10013 34588
rect 11320 34544 11360 34672
rect 18115 34588 18124 34628
rect 18164 34588 19564 34628
rect 19604 34588 19613 34628
rect 21424 34544 21504 34564
rect 2851 34504 2860 34544
rect 2900 34504 3244 34544
rect 3284 34504 3293 34544
rect 6115 34504 6124 34544
rect 6164 34504 11360 34544
rect 12931 34504 12940 34544
rect 12980 34504 13516 34544
rect 13556 34504 14764 34544
rect 14804 34504 14813 34544
rect 17635 34504 17644 34544
rect 17684 34504 21504 34544
rect 21424 34484 21504 34504
rect 1411 34420 1420 34460
rect 1460 34420 1612 34460
rect 1652 34420 1661 34460
rect 1891 34420 1900 34460
rect 1940 34420 1949 34460
rect 7555 34420 7564 34460
rect 7604 34420 9908 34460
rect 13891 34420 13900 34460
rect 13940 34420 14572 34460
rect 14612 34420 14621 34460
rect 19267 34420 19276 34460
rect 19316 34420 19948 34460
rect 19988 34420 19997 34460
rect 0 34376 80 34396
rect 4483 34376 4541 34377
rect 0 34336 4340 34376
rect 4398 34336 4492 34376
rect 4532 34336 4541 34376
rect 6211 34336 6220 34376
rect 6260 34336 8332 34376
rect 8372 34336 8381 34376
rect 8611 34336 8620 34376
rect 8660 34336 8908 34376
rect 8948 34336 8957 34376
rect 9000 34336 9009 34376
rect 9049 34336 9580 34376
rect 9620 34336 9629 34376
rect 0 34316 80 34336
rect 4300 34292 4340 34336
rect 4483 34335 4541 34336
rect 7075 34292 7133 34293
rect 8323 34292 8381 34293
rect 1315 34252 1324 34292
rect 1364 34252 1804 34292
rect 1844 34252 1853 34292
rect 4300 34252 6508 34292
rect 6548 34252 7084 34292
rect 7124 34252 7133 34292
rect 7939 34252 7948 34292
rect 7988 34252 8332 34292
rect 8372 34252 8381 34292
rect 7075 34251 7133 34252
rect 8323 34251 8381 34252
rect 8995 34292 9053 34293
rect 9763 34292 9821 34293
rect 8995 34252 9004 34292
rect 9044 34252 9196 34292
rect 9236 34252 9772 34292
rect 9812 34252 9821 34292
rect 8995 34251 9053 34252
rect 9763 34251 9821 34252
rect 6307 34208 6365 34209
rect 8515 34208 8573 34209
rect 9868 34208 9908 34420
rect 10243 34336 10252 34376
rect 10292 34336 13804 34376
rect 13844 34336 13853 34376
rect 13987 34336 13996 34376
rect 14036 34336 14668 34376
rect 14708 34336 14717 34376
rect 15235 34292 15293 34293
rect 13123 34252 13132 34292
rect 13172 34252 13460 34292
rect 13507 34252 13516 34292
rect 13556 34252 14188 34292
rect 14228 34252 15244 34292
rect 15284 34252 15293 34292
rect 13420 34208 13460 34252
rect 15235 34251 15293 34252
rect 172 34168 5356 34208
rect 5396 34168 5405 34208
rect 5731 34168 5740 34208
rect 5780 34168 6316 34208
rect 6356 34168 6365 34208
rect 8430 34168 8524 34208
rect 8564 34168 8573 34208
rect 9091 34168 9100 34208
rect 9140 34168 9484 34208
rect 9524 34168 9533 34208
rect 9859 34168 9868 34208
rect 9908 34168 10348 34208
rect 10388 34168 11116 34208
rect 11156 34168 11165 34208
rect 13411 34168 13420 34208
rect 13460 34168 13469 34208
rect 15139 34168 15148 34208
rect 15188 34168 16012 34208
rect 16052 34168 16972 34208
rect 17012 34168 17021 34208
rect 20131 34168 20140 34208
rect 20180 34168 20716 34208
rect 20756 34168 20765 34208
rect 0 34040 80 34060
rect 172 34040 212 34168
rect 6307 34167 6365 34168
rect 8515 34167 8573 34168
rect 2947 34084 2956 34124
rect 2996 34084 8140 34124
rect 8180 34084 8189 34124
rect 8236 34084 10252 34124
rect 10292 34084 10301 34124
rect 13123 34084 13132 34124
rect 13172 34084 14476 34124
rect 14516 34084 14525 34124
rect 8236 34040 8276 34084
rect 0 34000 212 34040
rect 4919 34000 4928 34040
rect 4968 34000 5010 34040
rect 5050 34000 5092 34040
rect 5132 34000 5174 34040
rect 5214 34000 5256 34040
rect 5296 34000 5305 34040
rect 7171 34000 7180 34040
rect 7220 34000 8276 34040
rect 8419 34040 8477 34041
rect 9475 34040 9533 34041
rect 12067 34040 12125 34041
rect 21424 34040 21504 34060
rect 8419 34000 8428 34040
rect 8468 34000 9484 34040
rect 9524 34000 9533 34040
rect 10627 34000 10636 34040
rect 10676 34000 12076 34040
rect 12116 34000 12125 34040
rect 14275 34000 14284 34040
rect 14324 34000 19276 34040
rect 19316 34000 19325 34040
rect 20039 34000 20048 34040
rect 20088 34000 20130 34040
rect 20170 34000 20212 34040
rect 20252 34000 20294 34040
rect 20334 34000 20376 34040
rect 20416 34000 20425 34040
rect 21379 34000 21388 34040
rect 21428 34000 21504 34040
rect 0 33980 80 34000
rect 8419 33999 8477 34000
rect 9475 33999 9533 34000
rect 12067 33999 12125 34000
rect 21424 33980 21504 34000
rect 2500 33916 5972 33956
rect 7843 33916 7852 33956
rect 7892 33916 9388 33956
rect 9428 33916 9437 33956
rect 11683 33916 11692 33956
rect 11732 33916 11772 33956
rect 13027 33916 13036 33956
rect 13076 33916 13324 33956
rect 13364 33916 13373 33956
rect 16675 33916 16684 33956
rect 16724 33916 16876 33956
rect 16916 33916 17932 33956
rect 17972 33916 17981 33956
rect 2500 33872 2540 33916
rect 5932 33872 5972 33916
rect 11692 33872 11732 33916
rect 11971 33872 12029 33873
rect 1228 33832 2540 33872
rect 4099 33832 4108 33872
rect 4148 33832 5740 33872
rect 5780 33832 5789 33872
rect 5923 33832 5932 33872
rect 5972 33832 11980 33872
rect 12020 33832 12029 33872
rect 12547 33832 12556 33872
rect 12596 33832 16396 33872
rect 16436 33832 16445 33872
rect 0 33704 80 33724
rect 1228 33704 1268 33832
rect 11971 33831 12029 33832
rect 1603 33788 1661 33789
rect 1603 33748 1612 33788
rect 1652 33748 4300 33788
rect 4340 33748 9964 33788
rect 10004 33748 10252 33788
rect 10292 33748 10301 33788
rect 11395 33748 11404 33788
rect 11444 33748 11692 33788
rect 11732 33748 11741 33788
rect 12355 33748 12364 33788
rect 12404 33748 12748 33788
rect 12788 33748 13804 33788
rect 13844 33748 13853 33788
rect 16867 33748 16876 33788
rect 16916 33748 17164 33788
rect 17204 33748 17213 33788
rect 1603 33747 1661 33748
rect 8419 33704 8477 33705
rect 19555 33704 19613 33705
rect 0 33664 1268 33704
rect 2467 33664 2476 33704
rect 2516 33664 3340 33704
rect 3380 33664 3389 33704
rect 4003 33664 4012 33704
rect 4052 33664 5836 33704
rect 5876 33664 5885 33704
rect 7555 33664 7564 33704
rect 7604 33664 7852 33704
rect 7892 33664 7901 33704
rect 8227 33664 8236 33704
rect 8276 33664 8428 33704
rect 8468 33664 8477 33704
rect 8803 33664 8812 33704
rect 8852 33664 11360 33704
rect 12835 33664 12844 33704
rect 12884 33664 15436 33704
rect 15476 33664 15485 33704
rect 19470 33664 19564 33704
rect 19604 33664 19613 33704
rect 0 33644 80 33664
rect 8419 33663 8477 33664
rect 7747 33620 7805 33621
rect 7939 33620 7997 33621
rect 9667 33620 9725 33621
rect 7651 33580 7660 33620
rect 7700 33580 7756 33620
rect 7796 33580 7948 33620
rect 7988 33580 7997 33620
rect 8899 33580 8908 33620
rect 8948 33580 9676 33620
rect 9716 33580 9725 33620
rect 11320 33620 11360 33664
rect 19555 33663 19613 33664
rect 11320 33580 12268 33620
rect 12308 33580 12317 33620
rect 15331 33580 15340 33620
rect 15380 33580 16684 33620
rect 16724 33580 16733 33620
rect 7747 33579 7805 33580
rect 7939 33579 7997 33580
rect 9667 33579 9725 33580
rect 7267 33536 7325 33537
rect 21424 33536 21504 33556
rect 3811 33496 3820 33536
rect 3860 33496 7276 33536
rect 7316 33496 7325 33536
rect 8035 33496 8044 33536
rect 8084 33496 9676 33536
rect 9716 33496 9725 33536
rect 20611 33496 20620 33536
rect 20660 33496 21504 33536
rect 7267 33495 7325 33496
rect 21424 33476 21504 33496
rect 7363 33412 7372 33452
rect 7412 33412 7948 33452
rect 7988 33412 8524 33452
rect 8564 33412 8573 33452
rect 8620 33412 8840 33452
rect 9283 33412 9292 33452
rect 9332 33412 9964 33452
rect 10004 33412 10013 33452
rect 10243 33412 10252 33452
rect 10292 33412 17260 33452
rect 17300 33412 17309 33452
rect 0 33368 80 33388
rect 1699 33368 1757 33369
rect 8620 33368 8660 33412
rect 0 33328 1708 33368
rect 1748 33328 1757 33368
rect 1891 33328 1900 33368
rect 1940 33328 2476 33368
rect 2516 33328 8660 33368
rect 0 33308 80 33328
rect 1699 33327 1757 33328
rect 8800 33284 8840 33412
rect 12259 33368 12317 33369
rect 9484 33328 11404 33368
rect 11444 33328 12268 33368
rect 12308 33328 12317 33368
rect 12643 33328 12652 33368
rect 12692 33328 12844 33368
rect 12884 33328 12893 33368
rect 14083 33328 14092 33368
rect 14132 33328 19948 33368
rect 19988 33328 19997 33368
rect 9484 33284 9524 33328
rect 12259 33327 12317 33328
rect 3679 33244 3688 33284
rect 3728 33244 3770 33284
rect 3810 33244 3852 33284
rect 3892 33244 3934 33284
rect 3974 33244 4016 33284
rect 4056 33244 4065 33284
rect 8131 33244 8140 33284
rect 8180 33244 8332 33284
rect 8372 33244 8381 33284
rect 8800 33244 9524 33284
rect 9571 33244 9580 33284
rect 9620 33244 10156 33284
rect 10196 33244 10205 33284
rect 11320 33244 11500 33284
rect 11540 33244 18068 33284
rect 18799 33244 18808 33284
rect 18848 33244 18890 33284
rect 18930 33244 18972 33284
rect 19012 33244 19054 33284
rect 19094 33244 19136 33284
rect 19176 33244 19185 33284
rect 1891 33200 1949 33201
rect 11320 33200 11360 33244
rect 1891 33160 1900 33200
rect 1940 33160 2284 33200
rect 2324 33160 2333 33200
rect 2659 33160 2668 33200
rect 2708 33160 10444 33200
rect 10484 33160 11360 33200
rect 18028 33200 18068 33244
rect 19363 33200 19421 33201
rect 18028 33160 19372 33200
rect 19412 33160 19421 33200
rect 20131 33160 20140 33200
rect 20180 33160 20620 33200
rect 20660 33160 20669 33200
rect 1891 33159 1949 33160
rect 19363 33159 19421 33160
rect 5827 33076 5836 33116
rect 5876 33076 6220 33116
rect 6260 33076 6269 33116
rect 6979 33076 6988 33116
rect 7028 33076 7372 33116
rect 7412 33076 7421 33116
rect 9004 33076 9196 33116
rect 9236 33076 11020 33116
rect 11060 33076 11069 33116
rect 15427 33076 15436 33116
rect 15476 33076 15485 33116
rect 0 33032 80 33052
rect 9004 33032 9044 33076
rect 0 32992 940 33032
rect 980 32992 989 33032
rect 3148 32992 9044 33032
rect 9091 32992 9100 33032
rect 9140 32992 9484 33032
rect 9524 32992 9533 33032
rect 0 32972 80 32992
rect 3148 32948 3188 32992
rect 12643 32948 12701 32949
rect 15436 32948 15476 33076
rect 21424 33032 21504 33052
rect 15619 32992 15628 33032
rect 15668 32992 16012 33032
rect 16052 32992 16061 33032
rect 19651 32992 19660 33032
rect 19700 32992 21504 33032
rect 21424 32972 21504 32992
rect 3139 32908 3148 32948
rect 3188 32908 3197 32948
rect 5731 32908 5740 32948
rect 5780 32908 6609 32948
rect 6649 32908 6658 32948
rect 7939 32908 7948 32948
rect 7988 32908 9388 32948
rect 9428 32908 9437 32948
rect 12643 32908 12652 32948
rect 12692 32908 14092 32948
rect 14132 32908 14141 32948
rect 15436 32908 19948 32948
rect 19988 32908 19997 32948
rect 12643 32907 12701 32908
rect 9955 32864 10013 32865
rect 14947 32864 15005 32865
rect 15907 32864 15965 32865
rect 2755 32824 2764 32864
rect 2804 32824 3724 32864
rect 3764 32824 3773 32864
rect 4099 32824 4108 32864
rect 4148 32824 6124 32864
rect 6164 32824 6173 32864
rect 6499 32824 6508 32864
rect 6548 32824 7564 32864
rect 7604 32824 7613 32864
rect 8803 32824 8812 32864
rect 8852 32824 9484 32864
rect 9524 32824 9533 32864
rect 9667 32824 9676 32864
rect 9716 32824 9964 32864
rect 10004 32824 10013 32864
rect 13123 32824 13132 32864
rect 13172 32824 13324 32864
rect 13364 32824 13373 32864
rect 14947 32824 14956 32864
rect 14996 32824 15340 32864
rect 15380 32824 15389 32864
rect 15822 32824 15916 32864
rect 15956 32824 15965 32864
rect 16291 32824 16300 32864
rect 16340 32824 17260 32864
rect 17300 32824 17309 32864
rect 9955 32823 10013 32824
rect 14947 32823 15005 32824
rect 15907 32823 15965 32824
rect 4291 32780 4349 32781
rect 4675 32780 4733 32781
rect 4291 32740 4300 32780
rect 4340 32740 4396 32780
rect 4436 32740 4684 32780
rect 4724 32740 4733 32780
rect 4291 32739 4349 32740
rect 4675 32739 4733 32740
rect 9283 32780 9341 32781
rect 9283 32740 9292 32780
rect 9332 32740 9388 32780
rect 9428 32740 9437 32780
rect 12259 32740 12268 32780
rect 12308 32740 13076 32780
rect 13795 32740 13804 32780
rect 13844 32740 16972 32780
rect 17012 32740 17021 32780
rect 17347 32740 17356 32780
rect 17396 32740 17740 32780
rect 17780 32740 17789 32780
rect 9283 32739 9341 32740
rect 0 32696 80 32716
rect 4684 32696 4724 32739
rect 9571 32696 9629 32697
rect 0 32656 2092 32696
rect 2132 32656 2141 32696
rect 3139 32656 3148 32696
rect 3188 32656 3532 32696
rect 3572 32656 3581 32696
rect 4684 32656 8948 32696
rect 0 32636 80 32656
rect 8323 32612 8381 32613
rect 8908 32612 8948 32656
rect 9571 32656 9580 32696
rect 9620 32656 9676 32696
rect 9716 32656 9725 32696
rect 9571 32655 9629 32656
rect 3043 32572 3052 32612
rect 3092 32572 5932 32612
rect 5972 32572 5981 32612
rect 8323 32572 8332 32612
rect 8372 32572 8716 32612
rect 8756 32572 8765 32612
rect 8908 32572 11360 32612
rect 8323 32571 8381 32572
rect 4919 32488 4928 32528
rect 4968 32488 5010 32528
rect 5050 32488 5092 32528
rect 5132 32488 5174 32528
rect 5214 32488 5256 32528
rect 5296 32488 5305 32528
rect 8227 32488 8236 32528
rect 8276 32488 8285 32528
rect 8236 32444 8276 32488
rect 11320 32444 11360 32572
rect 13036 32528 13076 32740
rect 16483 32656 16492 32696
rect 16532 32656 16876 32696
rect 16916 32656 16925 32696
rect 20131 32656 20140 32696
rect 20180 32656 21292 32696
rect 21332 32656 21341 32696
rect 21424 32528 21504 32548
rect 13027 32488 13036 32528
rect 13076 32488 13085 32528
rect 20039 32488 20048 32528
rect 20088 32488 20130 32528
rect 20170 32488 20212 32528
rect 20252 32488 20294 32528
rect 20334 32488 20376 32528
rect 20416 32488 20425 32528
rect 20515 32488 20524 32528
rect 20564 32488 21504 32528
rect 21424 32468 21504 32488
rect 3331 32404 3340 32444
rect 3380 32404 5452 32444
rect 5492 32404 7564 32444
rect 7604 32404 9964 32444
rect 10004 32404 10013 32444
rect 11320 32404 11884 32444
rect 11924 32404 11933 32444
rect 0 32360 80 32380
rect 0 32320 1420 32360
rect 1460 32320 1469 32360
rect 2275 32320 2284 32360
rect 2324 32320 9580 32360
rect 9620 32320 9629 32360
rect 0 32300 80 32320
rect 2500 32236 17164 32276
rect 17204 32236 17213 32276
rect 1795 32152 1804 32192
rect 1844 32152 2380 32192
rect 2420 32152 2429 32192
rect 2500 32108 2540 32236
rect 4387 32192 4445 32193
rect 8707 32192 8765 32193
rect 14659 32192 14717 32193
rect 4195 32152 4204 32192
rect 4244 32152 4396 32192
rect 4436 32152 4445 32192
rect 8622 32152 8716 32192
rect 8756 32152 8765 32192
rect 12931 32152 12940 32192
rect 12980 32152 13708 32192
rect 13748 32152 13757 32192
rect 14563 32152 14572 32192
rect 14612 32152 14668 32192
rect 14708 32152 14717 32192
rect 4387 32151 4445 32152
rect 8707 32151 8765 32152
rect 14659 32151 14717 32152
rect 16579 32192 16637 32193
rect 16579 32152 16588 32192
rect 16628 32152 18124 32192
rect 18164 32152 18173 32192
rect 19843 32152 19852 32192
rect 19892 32152 20044 32192
rect 20084 32152 20093 32192
rect 16579 32151 16637 32152
rect 15331 32108 15389 32109
rect 16387 32108 16445 32109
rect 1027 32068 1036 32108
rect 1076 32068 2540 32108
rect 6307 32068 6316 32108
rect 6356 32068 10636 32108
rect 10676 32068 10685 32108
rect 14659 32068 14668 32108
rect 14708 32068 15340 32108
rect 15380 32068 15389 32108
rect 16302 32068 16396 32108
rect 16436 32068 16445 32108
rect 15331 32067 15389 32068
rect 16387 32067 16445 32068
rect 0 32024 80 32044
rect 21424 32024 21504 32044
rect 0 31984 6508 32024
rect 6548 31984 6557 32024
rect 15043 31984 15052 32024
rect 15092 31984 18220 32024
rect 18260 31984 19276 32024
rect 19316 31984 19325 32024
rect 19843 31984 19852 32024
rect 19892 31984 21504 32024
rect 0 31964 80 31984
rect 21424 31964 21504 31984
rect 3331 31900 3340 31940
rect 3380 31900 3628 31940
rect 3668 31900 3677 31940
rect 5635 31900 5644 31940
rect 5684 31900 6028 31940
rect 6068 31900 6077 31940
rect 13987 31900 13996 31940
rect 14036 31900 14188 31940
rect 14228 31900 14860 31940
rect 14900 31900 14909 31940
rect 16387 31900 16396 31940
rect 16436 31900 16876 31940
rect 16916 31900 16925 31940
rect 163 31816 172 31856
rect 212 31816 12076 31856
rect 12116 31816 12125 31856
rect 14371 31772 14429 31773
rect 3679 31732 3688 31772
rect 3728 31732 3770 31772
rect 3810 31732 3852 31772
rect 3892 31732 3934 31772
rect 3974 31732 4016 31772
rect 4056 31732 4065 31772
rect 5827 31732 5836 31772
rect 5876 31732 6604 31772
rect 6644 31732 7084 31772
rect 7124 31732 7133 31772
rect 14275 31732 14284 31772
rect 14324 31732 14380 31772
rect 14420 31732 14429 31772
rect 18799 31732 18808 31772
rect 18848 31732 18890 31772
rect 18930 31732 18972 31772
rect 19012 31732 19054 31772
rect 19094 31732 19136 31772
rect 19176 31732 19185 31772
rect 14371 31731 14429 31732
rect 0 31688 80 31708
rect 0 31648 10924 31688
rect 10964 31648 11980 31688
rect 12020 31648 12029 31688
rect 13507 31648 13516 31688
rect 13556 31648 19660 31688
rect 19700 31648 19709 31688
rect 0 31628 80 31648
rect 2380 31564 7948 31604
rect 7988 31564 7997 31604
rect 17155 31564 17164 31604
rect 17204 31564 17213 31604
rect 2380 31520 2420 31564
rect 17164 31520 17204 31564
rect 21424 31520 21504 31540
rect 1315 31480 1324 31520
rect 1364 31480 1612 31520
rect 1652 31480 1661 31520
rect 2371 31480 2380 31520
rect 2420 31480 2429 31520
rect 7555 31480 7564 31520
rect 7604 31480 7756 31520
rect 7796 31480 7805 31520
rect 8515 31480 8524 31520
rect 8564 31480 8908 31520
rect 8948 31480 8957 31520
rect 12163 31480 12172 31520
rect 12212 31480 14612 31520
rect 14659 31480 14668 31520
rect 14708 31480 15436 31520
rect 15476 31480 15485 31520
rect 17164 31480 19276 31520
rect 19316 31480 19325 31520
rect 20227 31480 20236 31520
rect 20276 31480 21504 31520
rect 14572 31437 14612 31480
rect 21424 31460 21504 31480
rect 14563 31436 14621 31437
rect 17251 31436 17309 31437
rect 2500 31396 14228 31436
rect 14478 31396 14572 31436
rect 14612 31396 15244 31436
rect 15284 31396 15293 31436
rect 16675 31396 16684 31436
rect 16724 31396 16876 31436
rect 16916 31396 16925 31436
rect 17251 31396 17260 31436
rect 17300 31396 17836 31436
rect 17876 31396 17885 31436
rect 18307 31396 18316 31436
rect 18356 31396 19180 31436
rect 19220 31396 19229 31436
rect 19747 31396 19756 31436
rect 19796 31396 20044 31436
rect 20084 31396 20093 31436
rect 0 31352 80 31372
rect 2500 31352 2540 31396
rect 5443 31352 5501 31353
rect 6403 31352 6461 31353
rect 8707 31352 8765 31353
rect 12355 31352 12413 31353
rect 0 31312 2540 31352
rect 2659 31312 2668 31352
rect 2708 31312 2956 31352
rect 2996 31312 3005 31352
rect 5443 31312 5452 31352
rect 5492 31312 6412 31352
rect 6452 31312 6461 31352
rect 8419 31312 8428 31352
rect 8468 31312 8716 31352
rect 8756 31312 8765 31352
rect 10819 31312 10828 31352
rect 10868 31312 12364 31352
rect 12404 31312 12748 31352
rect 12788 31312 12797 31352
rect 0 31292 80 31312
rect 5443 31311 5501 31312
rect 6403 31311 6461 31312
rect 8707 31311 8765 31312
rect 12355 31311 12413 31312
rect 4483 31268 4541 31269
rect 9283 31268 9341 31269
rect 2467 31228 2476 31268
rect 2516 31228 3916 31268
rect 3956 31228 4492 31268
rect 4532 31228 5548 31268
rect 5588 31228 5597 31268
rect 6403 31228 6412 31268
rect 6452 31228 8812 31268
rect 8852 31228 9292 31268
rect 9332 31228 9341 31268
rect 11203 31228 11212 31268
rect 11252 31228 13324 31268
rect 13364 31228 13373 31268
rect 4483 31227 4541 31228
rect 9283 31227 9341 31228
rect 8803 31184 8861 31185
rect 12163 31184 12221 31185
rect 4099 31144 4108 31184
rect 4148 31144 4780 31184
rect 4820 31144 4829 31184
rect 5731 31144 5740 31184
rect 5780 31144 6316 31184
rect 6356 31144 6365 31184
rect 6499 31144 6508 31184
rect 6548 31144 6700 31184
rect 6740 31144 6749 31184
rect 7747 31144 7756 31184
rect 7796 31144 8812 31184
rect 8852 31144 8861 31184
rect 12078 31144 12172 31184
rect 12212 31144 12221 31184
rect 14188 31184 14228 31396
rect 14563 31395 14621 31396
rect 17251 31395 17309 31396
rect 14275 31312 14284 31352
rect 14324 31312 14572 31352
rect 14612 31312 14865 31352
rect 14905 31312 15148 31352
rect 15188 31312 15197 31352
rect 16483 31312 16492 31352
rect 16532 31312 17164 31352
rect 17204 31312 17213 31352
rect 17347 31312 17356 31352
rect 17396 31312 18124 31352
rect 18164 31312 18173 31352
rect 18499 31312 18508 31352
rect 18548 31312 19372 31352
rect 19412 31312 19421 31352
rect 17356 31268 17396 31312
rect 18211 31268 18269 31269
rect 16867 31228 16876 31268
rect 16916 31228 17396 31268
rect 17620 31228 18220 31268
rect 18260 31228 18269 31268
rect 17620 31184 17660 31228
rect 18211 31227 18269 31228
rect 19459 31184 19517 31185
rect 14188 31144 14764 31184
rect 14804 31144 14813 31184
rect 16675 31144 16684 31184
rect 16724 31144 17660 31184
rect 18979 31144 18988 31184
rect 19028 31144 19468 31184
rect 19508 31144 19517 31184
rect 8803 31143 8861 31144
rect 12163 31143 12221 31144
rect 19459 31143 19517 31144
rect 3427 31100 3485 31101
rect 3331 31060 3340 31100
rect 3380 31060 3436 31100
rect 3476 31060 7508 31100
rect 7555 31060 7564 31100
rect 7604 31060 8524 31100
rect 8564 31060 8573 31100
rect 14659 31060 14668 31100
rect 14708 31060 15052 31100
rect 15092 31060 15101 31100
rect 16003 31060 16012 31100
rect 16052 31060 17068 31100
rect 17108 31060 17452 31100
rect 17492 31060 17501 31100
rect 3427 31059 3485 31060
rect 0 31016 80 31036
rect 7468 31016 7508 31060
rect 16483 31016 16541 31017
rect 21424 31016 21504 31036
rect 0 30976 2668 31016
rect 2708 30976 2717 31016
rect 4919 30976 4928 31016
rect 4968 30976 5010 31016
rect 5050 30976 5092 31016
rect 5132 30976 5174 31016
rect 5214 30976 5256 31016
rect 5296 30976 5305 31016
rect 6691 30976 6700 31016
rect 6740 30976 7372 31016
rect 7412 30976 7421 31016
rect 7468 30976 10540 31016
rect 10580 30976 10589 31016
rect 15139 30976 15148 31016
rect 15188 30976 16108 31016
rect 16148 30976 16157 31016
rect 16483 30976 16492 31016
rect 16532 30976 19660 31016
rect 19700 30976 19709 31016
rect 20039 30976 20048 31016
rect 20088 30976 20130 31016
rect 20170 30976 20212 31016
rect 20252 30976 20294 31016
rect 20334 30976 20376 31016
rect 20416 30976 20425 31016
rect 20707 30976 20716 31016
rect 20756 30976 21504 31016
rect 0 30956 80 30976
rect 16483 30975 16541 30976
rect 21424 30956 21504 30976
rect 7747 30892 7756 30932
rect 7796 30892 8620 30932
rect 8660 30892 8669 30932
rect 9091 30892 9100 30932
rect 9140 30892 11360 30932
rect 13315 30892 13324 30932
rect 13364 30892 15724 30932
rect 15764 30892 15773 30932
rect 11320 30848 11360 30892
rect 5539 30808 5548 30848
rect 5588 30808 11212 30848
rect 11252 30808 11261 30848
rect 11320 30808 13844 30848
rect 13987 30808 13996 30848
rect 14036 30808 14228 30848
rect 18307 30808 18316 30848
rect 18356 30808 18796 30848
rect 18836 30808 18845 30848
rect 5539 30764 5597 30765
rect 5347 30724 5356 30764
rect 5396 30724 5548 30764
rect 5588 30724 6604 30764
rect 6644 30724 8620 30764
rect 8660 30724 9772 30764
rect 9812 30724 9821 30764
rect 10243 30724 10252 30764
rect 10292 30724 12076 30764
rect 12116 30724 13420 30764
rect 13460 30724 13469 30764
rect 5539 30723 5597 30724
rect 0 30680 80 30700
rect 8995 30680 9053 30681
rect 0 30640 1708 30680
rect 1748 30640 4820 30680
rect 4867 30640 4876 30680
rect 4916 30640 6124 30680
rect 6164 30640 6173 30680
rect 8910 30640 9004 30680
rect 9044 30640 9053 30680
rect 0 30620 80 30640
rect 4780 30596 4820 30640
rect 8995 30639 9053 30640
rect 9004 30596 9044 30639
rect 1603 30556 1612 30596
rect 1652 30556 2860 30596
rect 2900 30556 2909 30596
rect 4780 30556 5260 30596
rect 5300 30556 5309 30596
rect 9004 30556 12940 30596
rect 12980 30556 12989 30596
rect 4099 30512 4157 30513
rect 4099 30472 4108 30512
rect 4148 30472 9100 30512
rect 9140 30472 9149 30512
rect 4099 30471 4157 30472
rect 13804 30428 13844 30808
rect 13891 30680 13949 30681
rect 13891 30640 13900 30680
rect 13940 30640 13996 30680
rect 14036 30640 14045 30680
rect 13891 30639 13949 30640
rect 14188 30512 14228 30808
rect 14371 30680 14429 30681
rect 19555 30680 19613 30681
rect 14371 30640 14380 30680
rect 14420 30640 14476 30680
rect 14516 30640 14525 30680
rect 16579 30640 16588 30680
rect 16628 30640 16876 30680
rect 16916 30640 17204 30680
rect 17251 30640 17260 30680
rect 17300 30640 17932 30680
rect 17972 30640 17981 30680
rect 19555 30640 19564 30680
rect 19604 30640 20044 30680
rect 20084 30640 20093 30680
rect 14371 30639 14429 30640
rect 17164 30596 17204 30640
rect 15523 30556 15532 30596
rect 15572 30556 15581 30596
rect 15715 30556 15724 30596
rect 15764 30556 16340 30596
rect 17155 30556 17164 30596
rect 17204 30556 17213 30596
rect 14179 30472 14188 30512
rect 14228 30472 14237 30512
rect 15532 30428 15572 30556
rect 16300 30512 16340 30556
rect 17260 30512 17300 30640
rect 19555 30639 19613 30640
rect 17539 30596 17597 30597
rect 17443 30556 17452 30596
rect 17492 30556 17548 30596
rect 17588 30556 17597 30596
rect 17539 30555 17597 30556
rect 16291 30472 16300 30512
rect 16340 30472 16349 30512
rect 16867 30472 16876 30512
rect 16916 30472 17300 30512
rect 18595 30512 18653 30513
rect 21424 30512 21504 30532
rect 18595 30472 18604 30512
rect 18644 30472 18892 30512
rect 18932 30472 18941 30512
rect 20611 30472 20620 30512
rect 20660 30472 21504 30512
rect 18595 30471 18653 30472
rect 21424 30452 21504 30472
rect 12547 30388 12556 30428
rect 12596 30388 12940 30428
rect 12980 30388 12989 30428
rect 13804 30388 16012 30428
rect 16052 30388 19756 30428
rect 19796 30388 19805 30428
rect 0 30344 80 30364
rect 16387 30344 16445 30345
rect 0 30304 1324 30344
rect 1364 30304 1373 30344
rect 10435 30304 10444 30344
rect 10484 30304 12364 30344
rect 12404 30304 12413 30344
rect 16302 30304 16396 30344
rect 16436 30304 16445 30344
rect 17059 30304 17068 30344
rect 17108 30304 17260 30344
rect 17300 30304 17309 30344
rect 0 30284 80 30304
rect 16387 30303 16445 30304
rect 19267 30260 19325 30261
rect 2275 30220 2284 30260
rect 2324 30220 2764 30260
rect 2804 30220 2813 30260
rect 3679 30220 3688 30260
rect 3728 30220 3770 30260
rect 3810 30220 3852 30260
rect 3892 30220 3934 30260
rect 3974 30220 4016 30260
rect 4056 30220 4065 30260
rect 7459 30220 7468 30260
rect 7508 30220 7852 30260
rect 7892 30220 7901 30260
rect 8515 30220 8524 30260
rect 8564 30220 8812 30260
rect 8852 30220 8861 30260
rect 10915 30220 10924 30260
rect 10964 30220 11596 30260
rect 11636 30220 13516 30260
rect 13556 30220 13565 30260
rect 14947 30220 14956 30260
rect 14996 30220 15628 30260
rect 15668 30220 15677 30260
rect 18799 30220 18808 30260
rect 18848 30220 18890 30260
rect 18930 30220 18972 30260
rect 19012 30220 19054 30260
rect 19094 30220 19136 30260
rect 19176 30220 19185 30260
rect 19267 30220 19276 30260
rect 19316 30220 21100 30260
rect 21140 30220 21149 30260
rect 19267 30219 19325 30220
rect 3139 30176 3197 30177
rect 3053 30136 3148 30176
rect 3188 30136 3532 30176
rect 3572 30136 10348 30176
rect 10388 30136 10397 30176
rect 3139 30135 3197 30136
rect 3043 30092 3101 30093
rect 13987 30092 14045 30093
rect 2563 30052 2572 30092
rect 2612 30052 3052 30092
rect 3092 30052 3101 30092
rect 5251 30052 5260 30092
rect 5300 30052 6220 30092
rect 6260 30052 10676 30092
rect 11875 30052 11884 30092
rect 11924 30052 12460 30092
rect 12500 30052 12509 30092
rect 13603 30052 13612 30092
rect 13652 30052 13996 30092
rect 14036 30052 14045 30092
rect 18403 30052 18412 30092
rect 18452 30052 18892 30092
rect 18932 30052 18941 30092
rect 19459 30052 19468 30092
rect 19508 30052 19660 30092
rect 19700 30052 19709 30092
rect 3043 30051 3101 30052
rect 0 30008 80 30028
rect 0 29968 3244 30008
rect 3284 29968 5492 30008
rect 8803 29968 8812 30008
rect 8852 29968 9388 30008
rect 9428 29968 9437 30008
rect 0 29948 80 29968
rect 1315 29840 1373 29841
rect 1230 29800 1324 29840
rect 1364 29800 1373 29840
rect 4579 29800 4588 29840
rect 4628 29800 4780 29840
rect 4820 29800 4829 29840
rect 1315 29799 1373 29800
rect 0 29672 80 29692
rect 0 29632 212 29672
rect 2755 29632 2764 29672
rect 2804 29632 2956 29672
rect 2996 29632 3005 29672
rect 0 29612 80 29632
rect 172 29504 212 29632
rect 3043 29588 3101 29589
rect 5452 29588 5492 29968
rect 10636 29924 10676 30052
rect 13987 30051 14045 30052
rect 21424 30008 21504 30028
rect 11395 29968 11404 30008
rect 11444 29968 11692 30008
rect 11732 29968 11741 30008
rect 13507 29968 13516 30008
rect 13556 29968 13804 30008
rect 13844 29968 13853 30008
rect 16963 29968 16972 30008
rect 17012 29968 17021 30008
rect 17827 29968 17836 30008
rect 17876 29968 21504 30008
rect 11779 29924 11837 29925
rect 16972 29924 17012 29968
rect 21424 29948 21504 29968
rect 8716 29884 10540 29924
rect 10580 29884 10589 29924
rect 10636 29884 11788 29924
rect 11828 29884 11837 29924
rect 15331 29884 15340 29924
rect 15380 29884 15916 29924
rect 15956 29884 15965 29924
rect 16876 29884 17012 29924
rect 8716 29840 8756 29884
rect 11779 29883 11837 29884
rect 12643 29840 12701 29841
rect 5539 29800 5548 29840
rect 5588 29800 5932 29840
rect 5972 29800 5981 29840
rect 8707 29800 8716 29840
rect 8756 29800 8765 29840
rect 8995 29800 9004 29840
rect 9044 29800 9236 29840
rect 9475 29800 9484 29840
rect 9524 29800 9868 29840
rect 9908 29800 9917 29840
rect 10051 29800 10060 29840
rect 10100 29800 11884 29840
rect 11924 29800 11933 29840
rect 12067 29800 12076 29840
rect 12116 29800 12652 29840
rect 12692 29800 12701 29840
rect 14371 29800 14380 29840
rect 14420 29800 14572 29840
rect 14612 29800 14621 29840
rect 6019 29716 6028 29756
rect 6068 29716 6604 29756
rect 6644 29716 6653 29756
rect 7363 29716 7372 29756
rect 7412 29716 8812 29756
rect 8852 29716 8861 29756
rect 9196 29672 9236 29800
rect 12643 29799 12701 29800
rect 16876 29756 16916 29884
rect 19555 29840 19613 29841
rect 16963 29800 16972 29840
rect 17012 29800 17164 29840
rect 17204 29800 17213 29840
rect 18691 29800 18700 29840
rect 18740 29800 19564 29840
rect 19604 29800 19756 29840
rect 19796 29800 19805 29840
rect 9571 29716 9580 29756
rect 9620 29716 15532 29756
rect 15572 29716 15581 29756
rect 16876 29716 17068 29756
rect 17108 29716 17117 29756
rect 16963 29672 17021 29673
rect 18700 29672 18740 29800
rect 19555 29799 19613 29800
rect 19171 29716 19180 29756
rect 19220 29716 20236 29756
rect 20276 29716 20285 29756
rect 5635 29632 5644 29672
rect 5684 29632 6316 29672
rect 6356 29632 6365 29672
rect 9187 29632 9196 29672
rect 9236 29632 9245 29672
rect 10339 29632 10348 29672
rect 10388 29632 13132 29672
rect 13172 29632 15092 29672
rect 15052 29588 15092 29632
rect 16963 29632 16972 29672
rect 17012 29632 17356 29672
rect 17396 29632 17405 29672
rect 17827 29632 17836 29672
rect 17876 29632 18740 29672
rect 16963 29631 17021 29632
rect 3043 29548 3052 29588
rect 3092 29548 5396 29588
rect 5452 29548 14324 29588
rect 15052 29548 17492 29588
rect 18019 29548 18028 29588
rect 18068 29548 18412 29588
rect 18452 29548 18461 29588
rect 19843 29548 19852 29588
rect 19892 29548 20852 29588
rect 3043 29547 3101 29548
rect 5356 29504 5396 29548
rect 6499 29504 6557 29505
rect 14284 29504 14324 29548
rect 17452 29504 17492 29548
rect 20812 29504 20852 29548
rect 21424 29504 21504 29524
rect 172 29464 2860 29504
rect 2900 29464 2909 29504
rect 4919 29464 4928 29504
rect 4968 29464 5010 29504
rect 5050 29464 5092 29504
rect 5132 29464 5174 29504
rect 5214 29464 5256 29504
rect 5296 29464 5305 29504
rect 5356 29464 6508 29504
rect 6548 29464 6557 29504
rect 6691 29464 6700 29504
rect 6740 29464 12076 29504
rect 12116 29464 12125 29504
rect 14275 29464 14284 29504
rect 14324 29464 17356 29504
rect 17396 29464 17405 29504
rect 17452 29464 19948 29504
rect 19988 29464 19997 29504
rect 20039 29464 20048 29504
rect 20088 29464 20130 29504
rect 20170 29464 20212 29504
rect 20252 29464 20294 29504
rect 20334 29464 20376 29504
rect 20416 29464 20425 29504
rect 20812 29464 21504 29504
rect 6499 29463 6557 29464
rect 21424 29444 21504 29464
rect 12259 29420 12317 29421
rect 3331 29380 3340 29420
rect 3380 29380 4588 29420
rect 4628 29380 7084 29420
rect 7124 29380 7133 29420
rect 7564 29380 10444 29420
rect 10484 29380 10493 29420
rect 12259 29380 12268 29420
rect 12308 29380 18700 29420
rect 18740 29380 18749 29420
rect 0 29336 80 29356
rect 5164 29336 5204 29380
rect 0 29296 3052 29336
rect 3092 29296 3101 29336
rect 5155 29296 5164 29336
rect 5204 29296 5213 29336
rect 5443 29296 5452 29336
rect 5492 29296 7468 29336
rect 7508 29296 7517 29336
rect 0 29276 80 29296
rect 5443 29252 5501 29253
rect 6499 29252 6557 29253
rect 7564 29252 7604 29380
rect 12259 29379 12317 29380
rect 11971 29336 12029 29337
rect 18403 29336 18461 29337
rect 7651 29296 7660 29336
rect 7700 29296 7709 29336
rect 8131 29296 8140 29336
rect 8180 29296 8812 29336
rect 8852 29296 8861 29336
rect 11971 29296 11980 29336
rect 12020 29296 15820 29336
rect 15860 29296 18068 29336
rect 5347 29212 5356 29252
rect 5396 29212 5452 29252
rect 5492 29212 5501 29252
rect 5443 29211 5501 29212
rect 5836 29212 6220 29252
rect 6260 29212 6269 29252
rect 6499 29212 6508 29252
rect 6548 29212 7604 29252
rect 7660 29252 7700 29296
rect 11971 29295 12029 29296
rect 14179 29252 14237 29253
rect 15427 29252 15485 29253
rect 18028 29252 18068 29296
rect 18403 29296 18412 29336
rect 18452 29296 18508 29336
rect 18548 29296 18557 29336
rect 18883 29296 18892 29336
rect 18932 29296 20620 29336
rect 20660 29296 20669 29336
rect 18403 29295 18461 29296
rect 7660 29212 8908 29252
rect 8948 29212 8957 29252
rect 14083 29212 14092 29252
rect 14132 29212 14188 29252
rect 14228 29212 14237 29252
rect 14467 29212 14476 29252
rect 14516 29212 14764 29252
rect 14804 29212 14813 29252
rect 15427 29212 15436 29252
rect 15476 29212 15724 29252
rect 15764 29212 15773 29252
rect 16771 29212 16780 29252
rect 16820 29212 17972 29252
rect 18028 29212 18988 29252
rect 19028 29212 19037 29252
rect 20515 29212 20524 29252
rect 20564 29212 21388 29252
rect 21428 29212 21437 29252
rect 4099 29168 4157 29169
rect 5836 29168 5876 29212
rect 6499 29211 6557 29212
rect 14179 29211 14237 29212
rect 15427 29211 15485 29212
rect 14947 29168 15005 29169
rect 17932 29168 17972 29212
rect 3907 29128 3916 29168
rect 3956 29128 4108 29168
rect 4148 29128 4157 29168
rect 4771 29128 4780 29168
rect 4820 29128 5836 29168
rect 5876 29128 5885 29168
rect 6019 29128 6028 29168
rect 6068 29128 6412 29168
rect 6452 29128 6461 29168
rect 8611 29128 8620 29168
rect 8660 29128 9292 29168
rect 9332 29128 9341 29168
rect 9667 29128 9676 29168
rect 9716 29128 11404 29168
rect 11444 29128 14956 29168
rect 14996 29128 15005 29168
rect 17155 29128 17164 29168
rect 17204 29128 17836 29168
rect 17876 29128 17885 29168
rect 17932 29128 18499 29168
rect 18539 29128 18548 29168
rect 18595 29128 18604 29168
rect 18644 29128 19468 29168
rect 19508 29128 19517 29168
rect 4099 29127 4157 29128
rect 14947 29127 15005 29128
rect 3427 29044 3436 29084
rect 3476 29044 5740 29084
rect 5780 29044 5789 29084
rect 5836 29044 6548 29084
rect 6595 29044 6604 29084
rect 6644 29044 8756 29084
rect 9763 29044 9772 29084
rect 9812 29044 11692 29084
rect 11732 29044 11741 29084
rect 11971 29044 11980 29084
rect 12020 29044 18644 29084
rect 18979 29044 18988 29084
rect 19028 29044 19412 29084
rect 20515 29044 20524 29084
rect 20564 29044 20812 29084
rect 20852 29044 20861 29084
rect 0 29001 80 29020
rect 0 29000 125 29001
rect 5836 29000 5876 29044
rect 6508 29000 6548 29044
rect 8515 29000 8573 29001
rect 8716 29000 8756 29044
rect 9763 29000 9821 29001
rect 11011 29000 11069 29001
rect 11779 29000 11837 29001
rect 18604 29000 18644 29044
rect 19372 29000 19412 29044
rect 19843 29000 19901 29001
rect 21424 29000 21504 29020
rect 0 28960 76 29000
rect 116 28960 125 29000
rect 5796 28960 5836 29000
rect 5876 28960 5885 29000
rect 6468 28960 6508 29000
rect 6548 28960 6557 29000
rect 8419 28960 8428 29000
rect 8468 28960 8524 29000
rect 8564 28960 8573 29000
rect 8676 28960 8716 29000
rect 8756 28960 8765 29000
rect 9283 28960 9292 29000
rect 9332 28960 9772 29000
rect 9812 28960 9821 29000
rect 10926 28960 11020 29000
rect 11060 28960 11069 29000
rect 11587 28960 11596 29000
rect 11636 28960 11788 29000
rect 11828 28960 11837 29000
rect 0 28959 125 28960
rect 8515 28959 8573 28960
rect 9763 28959 9821 28960
rect 11011 28959 11069 28960
rect 11779 28959 11837 28960
rect 11884 28960 16588 29000
rect 16628 28960 16637 29000
rect 18564 28960 18604 29000
rect 18644 28960 18653 29000
rect 19267 28960 19276 29000
rect 19316 28960 19412 29000
rect 19758 28960 19852 29000
rect 19892 28960 19901 29000
rect 21379 28960 21388 29000
rect 21428 28960 21504 29000
rect 0 28940 80 28959
rect 8899 28916 8957 28917
rect 11884 28916 11924 28960
rect 19843 28959 19901 28960
rect 21424 28940 21504 28960
rect 16195 28916 16253 28917
rect 3523 28876 3532 28916
rect 3572 28876 5644 28916
rect 5684 28876 5693 28916
rect 6595 28876 6604 28916
rect 6644 28876 7180 28916
rect 7220 28876 7229 28916
rect 8899 28876 8908 28916
rect 8948 28876 11924 28916
rect 11971 28876 11980 28916
rect 12020 28876 13132 28916
rect 13172 28876 13181 28916
rect 16110 28876 16204 28916
rect 16244 28876 16253 28916
rect 8899 28875 8957 28876
rect 16195 28875 16253 28876
rect 13987 28832 14045 28833
rect 8227 28792 8236 28832
rect 8276 28792 10732 28832
rect 10772 28792 10781 28832
rect 13795 28792 13804 28832
rect 13844 28792 13996 28832
rect 14036 28792 17452 28832
rect 17492 28792 17501 28832
rect 13987 28791 14045 28792
rect 14563 28748 14621 28749
rect 3679 28708 3688 28748
rect 3728 28708 3770 28748
rect 3810 28708 3852 28748
rect 3892 28708 3934 28748
rect 3974 28708 4016 28748
rect 4056 28708 4065 28748
rect 7171 28708 7180 28748
rect 7220 28708 7372 28748
rect 7412 28708 7421 28748
rect 11320 28708 14572 28748
rect 14612 28708 14621 28748
rect 18799 28708 18808 28748
rect 18848 28708 18890 28748
rect 18930 28708 18972 28748
rect 19012 28708 19054 28748
rect 19094 28708 19136 28748
rect 19176 28708 19185 28748
rect 0 28664 80 28684
rect 11320 28664 11360 28708
rect 14563 28707 14621 28708
rect 17635 28664 17693 28665
rect 0 28624 11360 28664
rect 12835 28624 12844 28664
rect 12884 28624 13228 28664
rect 13268 28624 13277 28664
rect 17443 28624 17452 28664
rect 17492 28624 17644 28664
rect 17684 28624 17693 28664
rect 0 28604 80 28624
rect 17635 28623 17693 28624
rect 8131 28580 8189 28581
rect 11779 28580 11837 28581
rect 2179 28540 2188 28580
rect 2228 28540 2476 28580
rect 2516 28540 2525 28580
rect 3139 28540 3148 28580
rect 3188 28540 8140 28580
rect 8180 28540 8189 28580
rect 9379 28540 9388 28580
rect 9428 28540 9580 28580
rect 9620 28540 9629 28580
rect 10723 28540 10732 28580
rect 10772 28540 11444 28580
rect 11694 28540 11788 28580
rect 11828 28540 11837 28580
rect 15523 28540 15532 28580
rect 15572 28540 16108 28580
rect 16148 28540 16157 28580
rect 8131 28539 8189 28540
rect 11404 28496 11444 28540
rect 11779 28539 11837 28540
rect 12355 28496 12413 28497
rect 17059 28496 17117 28497
rect 21424 28496 21504 28516
rect 1507 28456 1516 28496
rect 1556 28456 4684 28496
rect 4724 28456 4733 28496
rect 5731 28456 5740 28496
rect 5780 28456 5932 28496
rect 5972 28456 5981 28496
rect 6979 28456 6988 28496
rect 7028 28456 7037 28496
rect 7459 28456 7468 28496
rect 7508 28456 10100 28496
rect 10339 28456 10348 28496
rect 10388 28456 11116 28496
rect 11156 28456 11165 28496
rect 11395 28456 11404 28496
rect 11444 28456 11453 28496
rect 11683 28456 11692 28496
rect 11732 28456 12364 28496
rect 12404 28456 12413 28496
rect 16974 28456 17068 28496
rect 17108 28456 17117 28496
rect 20227 28456 20236 28496
rect 20276 28456 21504 28496
rect 1699 28372 1708 28412
rect 1748 28372 1996 28412
rect 2036 28372 2045 28412
rect 2500 28372 3916 28412
rect 3956 28372 3965 28412
rect 0 28328 80 28348
rect 2500 28328 2540 28372
rect 0 28288 1612 28328
rect 1652 28288 1661 28328
rect 1891 28288 1900 28328
rect 1940 28288 2540 28328
rect 3523 28288 3532 28328
rect 3572 28288 3581 28328
rect 4579 28288 4588 28328
rect 4628 28288 5740 28328
rect 5780 28288 5789 28328
rect 0 28268 80 28288
rect 3532 28244 3572 28288
rect 6988 28244 7028 28456
rect 8995 28372 9004 28412
rect 9044 28372 9196 28412
rect 9236 28372 9245 28412
rect 10060 28328 10100 28456
rect 12355 28455 12413 28456
rect 17059 28455 17117 28456
rect 21424 28436 21504 28456
rect 16963 28412 17021 28413
rect 11020 28372 11308 28412
rect 11348 28372 11788 28412
rect 11828 28372 11837 28412
rect 16878 28372 16972 28412
rect 17012 28372 17021 28412
rect 11020 28328 11060 28372
rect 16963 28371 17021 28372
rect 17539 28328 17597 28329
rect 8515 28288 8524 28328
rect 8564 28288 9676 28328
rect 9716 28288 9725 28328
rect 10051 28288 10060 28328
rect 10100 28288 10348 28328
rect 10388 28288 10397 28328
rect 11011 28288 11020 28328
rect 11060 28288 11069 28328
rect 11116 28288 12364 28328
rect 12404 28288 12413 28328
rect 17454 28288 17548 28328
rect 17588 28288 17597 28328
rect 9475 28244 9533 28245
rect 11116 28244 11156 28288
rect 17539 28287 17597 28288
rect 1507 28204 1516 28244
rect 1556 28204 2380 28244
rect 2420 28204 3572 28244
rect 5155 28204 5164 28244
rect 5204 28204 5644 28244
rect 5684 28204 5693 28244
rect 6988 28204 7084 28244
rect 7124 28204 7133 28244
rect 8323 28204 8332 28244
rect 8372 28204 9196 28244
rect 9236 28204 9245 28244
rect 9390 28204 9484 28244
rect 9524 28204 9533 28244
rect 10243 28204 10252 28244
rect 10292 28204 11156 28244
rect 11320 28204 14668 28244
rect 14708 28204 14717 28244
rect 9475 28203 9533 28204
rect 11320 28160 11360 28204
rect 12451 28160 12509 28161
rect 4483 28120 4492 28160
rect 4532 28120 9964 28160
rect 10004 28120 10013 28160
rect 10435 28120 10444 28160
rect 10484 28120 11360 28160
rect 11491 28120 11500 28160
rect 11540 28120 11692 28160
rect 11732 28120 11741 28160
rect 12366 28120 12460 28160
rect 12500 28120 12509 28160
rect 12643 28120 12652 28160
rect 12692 28120 12940 28160
rect 12980 28120 12989 28160
rect 18211 28120 18220 28160
rect 18260 28120 19468 28160
rect 19508 28120 19517 28160
rect 1891 28036 1900 28076
rect 1940 28036 2188 28076
rect 2228 28036 2237 28076
rect 0 27992 80 28012
rect 4492 27992 4532 28120
rect 12451 28119 12509 28120
rect 15907 28076 15965 28077
rect 4771 28036 4780 28076
rect 4820 28036 7468 28076
rect 7508 28036 9580 28076
rect 9620 28036 9629 28076
rect 10051 28036 10060 28076
rect 10100 28036 10540 28076
rect 10580 28036 10589 28076
rect 11203 28036 11212 28076
rect 11252 28036 15916 28076
rect 15956 28036 16588 28076
rect 16628 28036 16637 28076
rect 15907 28035 15965 28036
rect 9283 27992 9341 27993
rect 21424 27992 21504 28012
rect 0 27952 3436 27992
rect 3476 27952 4532 27992
rect 4919 27952 4928 27992
rect 4968 27952 5010 27992
rect 5050 27952 5092 27992
rect 5132 27952 5174 27992
rect 5214 27952 5256 27992
rect 5296 27952 5305 27992
rect 6979 27952 6988 27992
rect 7028 27952 7852 27992
rect 7892 27952 7901 27992
rect 8035 27952 8044 27992
rect 8084 27952 9196 27992
rect 9236 27952 9292 27992
rect 9332 27952 9360 27992
rect 20039 27952 20048 27992
rect 20088 27952 20130 27992
rect 20170 27952 20212 27992
rect 20252 27952 20294 27992
rect 20334 27952 20376 27992
rect 20416 27952 20425 27992
rect 20611 27952 20620 27992
rect 20660 27952 21504 27992
rect 0 27932 80 27952
rect 9283 27951 9341 27952
rect 21424 27932 21504 27952
rect 18211 27908 18269 27909
rect 1411 27868 1420 27908
rect 1460 27868 3340 27908
rect 3380 27868 3389 27908
rect 4387 27868 4396 27908
rect 4436 27868 10444 27908
rect 10484 27868 10493 27908
rect 18126 27868 18220 27908
rect 18260 27868 18269 27908
rect 18211 27867 18269 27868
rect 9475 27824 9533 27825
rect 18595 27824 18653 27825
rect 1603 27784 1612 27824
rect 1652 27784 1996 27824
rect 2036 27784 2045 27824
rect 3619 27784 3628 27824
rect 3668 27784 4588 27824
rect 4628 27784 4637 27824
rect 9475 27784 9484 27824
rect 9524 27784 12460 27824
rect 12500 27784 12509 27824
rect 12835 27784 12844 27824
rect 12884 27784 13804 27824
rect 13844 27784 13853 27824
rect 18499 27784 18508 27824
rect 18548 27784 18604 27824
rect 18644 27784 18653 27824
rect 9475 27783 9533 27784
rect 18595 27783 18653 27784
rect 2563 27740 2621 27741
rect 19459 27740 19517 27741
rect 2477 27700 2572 27740
rect 2612 27700 3532 27740
rect 3572 27700 3581 27740
rect 8803 27700 8812 27740
rect 8852 27700 9580 27740
rect 9620 27700 9629 27740
rect 9763 27700 9772 27740
rect 9812 27700 10348 27740
rect 10388 27700 10397 27740
rect 11971 27700 11980 27740
rect 12020 27700 13036 27740
rect 13076 27700 13085 27740
rect 13987 27700 13996 27740
rect 14036 27700 14476 27740
rect 14516 27700 15340 27740
rect 15380 27700 15389 27740
rect 16483 27700 16492 27740
rect 16532 27700 17164 27740
rect 17204 27700 18356 27740
rect 2563 27699 2621 27700
rect 0 27656 80 27676
rect 1603 27656 1661 27657
rect 4579 27656 4637 27657
rect 4771 27656 4829 27657
rect 18316 27656 18356 27700
rect 19459 27700 19468 27740
rect 19508 27700 19564 27740
rect 19604 27700 19613 27740
rect 19459 27699 19517 27700
rect 18403 27656 18461 27657
rect 0 27616 1364 27656
rect 0 27596 80 27616
rect 1324 27404 1364 27616
rect 1603 27616 1612 27656
rect 1652 27616 1708 27656
rect 1748 27616 4532 27656
rect 1603 27615 1661 27616
rect 4492 27572 4532 27616
rect 4579 27616 4588 27656
rect 4628 27616 4780 27656
rect 4820 27616 4829 27656
rect 6115 27616 6124 27656
rect 6164 27616 9524 27656
rect 14179 27616 14188 27656
rect 14228 27616 15148 27656
rect 15188 27616 15197 27656
rect 15427 27616 15436 27656
rect 15476 27616 16108 27656
rect 16148 27616 16157 27656
rect 17827 27616 17836 27656
rect 17876 27616 18124 27656
rect 18164 27616 18173 27656
rect 18307 27616 18316 27656
rect 18356 27616 18412 27656
rect 18452 27616 18461 27656
rect 19171 27616 19180 27656
rect 19220 27616 19948 27656
rect 19988 27616 19997 27656
rect 4579 27615 4637 27616
rect 4771 27615 4829 27616
rect 1411 27532 1420 27572
rect 1460 27532 4396 27572
rect 4436 27532 4445 27572
rect 4492 27532 4588 27572
rect 4628 27532 4637 27572
rect 8131 27532 8140 27572
rect 8180 27532 9004 27572
rect 9044 27532 9053 27572
rect 9379 27532 9388 27572
rect 9428 27532 9437 27572
rect 5539 27488 5597 27489
rect 9388 27488 9428 27532
rect 5443 27448 5452 27488
rect 5492 27448 5548 27488
rect 5588 27448 5597 27488
rect 8803 27448 8812 27488
rect 8852 27448 9428 27488
rect 9484 27488 9524 27616
rect 18403 27615 18461 27616
rect 9667 27532 9676 27572
rect 9716 27532 12172 27572
rect 12212 27532 12556 27572
rect 12596 27532 12605 27572
rect 15724 27532 21196 27572
rect 21236 27532 21245 27572
rect 15724 27488 15764 27532
rect 15907 27488 15965 27489
rect 21424 27488 21504 27508
rect 9484 27448 15764 27488
rect 15811 27448 15820 27488
rect 15860 27448 15916 27488
rect 15956 27448 15965 27488
rect 18883 27448 18892 27488
rect 18932 27448 21504 27488
rect 5539 27447 5597 27448
rect 15907 27447 15965 27448
rect 21424 27428 21504 27448
rect 8707 27404 8765 27405
rect 12355 27404 12413 27405
rect 1324 27364 6932 27404
rect 8622 27364 8716 27404
rect 8756 27364 8765 27404
rect 9379 27364 9388 27404
rect 9428 27364 11404 27404
rect 11444 27364 11453 27404
rect 12355 27364 12364 27404
rect 12404 27364 12460 27404
rect 12500 27364 12509 27404
rect 14659 27364 14668 27404
rect 14708 27364 15916 27404
rect 15956 27364 15965 27404
rect 19843 27364 19852 27404
rect 19892 27364 20812 27404
rect 20852 27364 20861 27404
rect 0 27320 80 27340
rect 6499 27320 6557 27321
rect 6892 27320 6932 27364
rect 8707 27363 8765 27364
rect 12355 27363 12413 27364
rect 0 27280 4628 27320
rect 0 27260 80 27280
rect 4588 27236 4628 27280
rect 6499 27280 6508 27320
rect 6548 27280 6700 27320
rect 6740 27280 6749 27320
rect 6892 27280 16876 27320
rect 16916 27280 17548 27320
rect 17588 27280 17597 27320
rect 6499 27279 6557 27280
rect 11491 27236 11549 27237
rect 15523 27236 15581 27237
rect 3679 27196 3688 27236
rect 3728 27196 3770 27236
rect 3810 27196 3852 27236
rect 3892 27196 3934 27236
rect 3974 27196 4016 27236
rect 4056 27196 4065 27236
rect 4588 27196 8812 27236
rect 8852 27196 8861 27236
rect 10915 27196 10924 27236
rect 10964 27196 11500 27236
rect 11540 27196 11549 27236
rect 12067 27196 12076 27236
rect 12116 27196 15052 27236
rect 15092 27196 15101 27236
rect 15235 27196 15244 27236
rect 15284 27196 15532 27236
rect 15572 27196 15581 27236
rect 15715 27196 15724 27236
rect 15764 27196 16204 27236
rect 16244 27196 16253 27236
rect 18799 27196 18808 27236
rect 18848 27196 18890 27236
rect 18930 27196 18972 27236
rect 19012 27196 19054 27236
rect 19094 27196 19136 27236
rect 19176 27196 19185 27236
rect 11491 27195 11549 27196
rect 15523 27195 15581 27196
rect 7075 27152 7133 27153
rect 2659 27112 2668 27152
rect 2708 27112 3052 27152
rect 3092 27112 3101 27152
rect 5347 27112 5356 27152
rect 5396 27112 5740 27152
rect 5780 27112 6604 27152
rect 6644 27112 6653 27152
rect 7075 27112 7084 27152
rect 7124 27112 13516 27152
rect 13556 27112 18700 27152
rect 18740 27112 18749 27152
rect 7075 27111 7133 27112
rect 3331 27068 3389 27069
rect 5731 27068 5789 27069
rect 1219 27028 1228 27068
rect 1268 27028 3340 27068
rect 3380 27028 5740 27068
rect 5780 27028 5789 27068
rect 14563 27028 14572 27068
rect 14612 27028 14860 27068
rect 14900 27028 18028 27068
rect 18068 27028 18077 27068
rect 3331 27027 3389 27028
rect 5731 27027 5789 27028
rect 0 26984 80 27004
rect 14179 26984 14237 26985
rect 21424 26984 21504 27004
rect 0 26944 6988 26984
rect 7028 26944 7037 26984
rect 8323 26944 8332 26984
rect 8372 26944 10252 26984
rect 10292 26944 11360 26984
rect 0 26924 80 26944
rect 11320 26900 11360 26944
rect 14179 26944 14188 26984
rect 14228 26944 15052 26984
rect 15092 26944 15101 26984
rect 15715 26944 15724 26984
rect 15764 26944 16396 26984
rect 16436 26944 16445 26984
rect 18115 26944 18124 26984
rect 18164 26944 18412 26984
rect 18452 26944 18461 26984
rect 19939 26944 19948 26984
rect 19988 26944 21504 26984
rect 14179 26943 14237 26944
rect 21424 26924 21504 26944
rect 12259 26900 12317 26901
rect 15715 26900 15773 26901
rect 1315 26860 1324 26900
rect 1364 26860 3092 26900
rect 3427 26860 3436 26900
rect 3476 26860 3628 26900
rect 3668 26860 3677 26900
rect 5923 26860 5932 26900
rect 5972 26860 8236 26900
rect 8276 26860 8285 26900
rect 9859 26860 9868 26900
rect 9908 26860 10828 26900
rect 10868 26860 10877 26900
rect 11320 26860 12076 26900
rect 12116 26860 12125 26900
rect 12259 26860 12268 26900
rect 12308 26860 12364 26900
rect 12404 26860 12413 26900
rect 15715 26860 15724 26900
rect 15764 26860 18452 26900
rect 3052 26732 3092 26860
rect 12259 26859 12317 26860
rect 15715 26859 15773 26860
rect 18412 26816 18452 26860
rect 3139 26776 3148 26816
rect 3188 26776 3916 26816
rect 3956 26776 5644 26816
rect 5684 26776 5836 26816
rect 5876 26776 5885 26816
rect 6211 26776 6220 26816
rect 6260 26776 6604 26816
rect 6644 26776 6653 26816
rect 7075 26776 7084 26816
rect 7124 26776 7133 26816
rect 8515 26776 8524 26816
rect 8564 26776 8908 26816
rect 8948 26776 9580 26816
rect 9620 26776 10732 26816
rect 10772 26776 10781 26816
rect 11107 26776 11116 26816
rect 11156 26776 11500 26816
rect 11540 26776 11549 26816
rect 11779 26776 11788 26816
rect 11828 26776 12268 26816
rect 12308 26776 12317 26816
rect 13795 26776 13804 26816
rect 13844 26776 14092 26816
rect 14132 26776 14476 26816
rect 14516 26776 14525 26816
rect 15139 26776 15148 26816
rect 15188 26776 16684 26816
rect 16724 26776 16733 26816
rect 18403 26776 18412 26816
rect 18452 26776 18461 26816
rect 18787 26776 18796 26816
rect 18836 26776 18988 26816
rect 19028 26776 19037 26816
rect 6499 26732 6557 26733
rect 7084 26732 7124 26776
rect 8995 26732 9053 26733
rect 11875 26732 11933 26733
rect 15907 26732 15965 26733
rect 3052 26692 4108 26732
rect 4148 26692 6260 26732
rect 0 26648 80 26668
rect 6220 26648 6260 26692
rect 6499 26692 6508 26732
rect 6548 26692 6892 26732
rect 6932 26692 6941 26732
rect 7084 26692 9004 26732
rect 9044 26692 11884 26732
rect 11924 26692 11933 26732
rect 15331 26692 15340 26732
rect 15380 26692 15916 26732
rect 15956 26692 15965 26732
rect 6499 26691 6557 26692
rect 8995 26691 9053 26692
rect 11875 26691 11933 26692
rect 15907 26691 15965 26692
rect 17635 26732 17693 26733
rect 18403 26732 18461 26733
rect 17635 26692 17644 26732
rect 17684 26692 18412 26732
rect 18452 26692 19756 26732
rect 19796 26692 19805 26732
rect 17635 26691 17693 26692
rect 18403 26691 18461 26692
rect 16963 26648 17021 26649
rect 0 26608 2540 26648
rect 3811 26608 3820 26648
rect 3860 26608 5356 26648
rect 5396 26608 5405 26648
rect 6211 26608 6220 26648
rect 6260 26608 6269 26648
rect 7171 26608 7180 26648
rect 7220 26608 10388 26648
rect 10435 26608 10444 26648
rect 10484 26608 10924 26648
rect 10964 26608 11348 26648
rect 11395 26608 11404 26648
rect 11444 26608 16972 26648
rect 17012 26608 17021 26648
rect 19555 26608 19564 26648
rect 19604 26608 21332 26648
rect 0 26588 80 26608
rect 2500 26564 2540 26608
rect 2500 26524 8756 26564
rect 2563 26480 2621 26481
rect 2851 26480 2909 26481
rect 7075 26480 7133 26481
rect 2478 26440 2572 26480
rect 2612 26440 2621 26480
rect 2766 26440 2860 26480
rect 2900 26440 2909 26480
rect 4919 26440 4928 26480
rect 4968 26440 5010 26480
rect 5050 26440 5092 26480
rect 5132 26440 5174 26480
rect 5214 26440 5256 26480
rect 5296 26440 5305 26480
rect 6019 26440 6028 26480
rect 6068 26440 6412 26480
rect 6452 26440 6461 26480
rect 6990 26440 7084 26480
rect 7124 26440 7133 26480
rect 8716 26480 8756 26524
rect 8716 26440 9428 26480
rect 2563 26439 2621 26440
rect 2851 26439 2909 26440
rect 6028 26396 6068 26440
rect 7075 26439 7133 26440
rect 9388 26396 9428 26440
rect 9955 26396 10013 26397
rect 4771 26356 4780 26396
rect 4820 26356 5548 26396
rect 5588 26356 6068 26396
rect 9091 26356 9100 26396
rect 9140 26356 9292 26396
rect 9332 26356 9341 26396
rect 9388 26356 9964 26396
rect 10004 26356 10013 26396
rect 10348 26396 10388 26608
rect 11308 26564 11348 26608
rect 16963 26607 17021 26608
rect 11299 26524 11308 26564
rect 11348 26524 11357 26564
rect 11491 26480 11549 26481
rect 18019 26480 18077 26481
rect 21292 26480 21332 26608
rect 21424 26480 21504 26500
rect 11406 26440 11500 26480
rect 11540 26440 11549 26480
rect 11491 26439 11549 26440
rect 14188 26440 14668 26480
rect 14708 26440 14717 26480
rect 14947 26440 14956 26480
rect 14996 26440 15820 26480
rect 15860 26440 15869 26480
rect 16291 26440 16300 26480
rect 16340 26440 17068 26480
rect 17108 26440 17117 26480
rect 17934 26440 18028 26480
rect 18068 26440 18077 26480
rect 18595 26440 18604 26480
rect 18644 26440 18892 26480
rect 18932 26440 18941 26480
rect 20039 26440 20048 26480
rect 20088 26440 20130 26480
rect 20170 26440 20212 26480
rect 20252 26440 20294 26480
rect 20334 26440 20376 26480
rect 20416 26440 20425 26480
rect 21292 26440 21504 26480
rect 12739 26396 12797 26397
rect 14188 26396 14228 26440
rect 18019 26439 18077 26440
rect 21424 26420 21504 26440
rect 14371 26396 14429 26397
rect 10348 26356 10828 26396
rect 10868 26356 10877 26396
rect 12739 26356 12748 26396
rect 12788 26356 13612 26396
rect 13652 26356 13804 26396
rect 13844 26356 14228 26396
rect 14286 26356 14380 26396
rect 14420 26356 16588 26396
rect 16628 26356 16637 26396
rect 9955 26355 10013 26356
rect 12739 26355 12797 26356
rect 14371 26355 14429 26356
rect 0 26312 80 26332
rect 8995 26312 9053 26313
rect 0 26272 1036 26312
rect 1076 26272 1085 26312
rect 4963 26272 4972 26312
rect 5012 26272 6028 26312
rect 6068 26272 6077 26312
rect 8910 26272 9004 26312
rect 9044 26272 9053 26312
rect 0 26252 80 26272
rect 8995 26271 9053 26272
rect 14179 26312 14237 26313
rect 16963 26312 17021 26313
rect 14179 26272 14188 26312
rect 14228 26272 14284 26312
rect 14324 26272 14333 26312
rect 14467 26272 14476 26312
rect 14516 26272 15244 26312
rect 15284 26272 15293 26312
rect 15715 26272 15724 26312
rect 15764 26272 16396 26312
rect 16436 26272 16445 26312
rect 16878 26272 16972 26312
rect 17012 26272 17021 26312
rect 18403 26272 18412 26312
rect 18452 26272 19180 26312
rect 19220 26272 19229 26312
rect 14179 26271 14237 26272
rect 16963 26271 17021 26272
rect 1315 26228 1373 26229
rect 1315 26188 1324 26228
rect 1364 26188 5108 26228
rect 6115 26188 6124 26228
rect 6164 26188 6700 26228
rect 6740 26188 6749 26228
rect 10819 26188 10828 26228
rect 10868 26188 13036 26228
rect 13076 26188 16204 26228
rect 16244 26188 16253 26228
rect 1315 26187 1373 26188
rect 1507 26144 1565 26145
rect 5068 26144 5108 26188
rect 1422 26104 1516 26144
rect 1556 26104 1565 26144
rect 2467 26104 2476 26144
rect 2516 26104 2764 26144
rect 2804 26104 2813 26144
rect 3331 26104 3340 26144
rect 3380 26104 5012 26144
rect 5068 26104 7660 26144
rect 7700 26104 7709 26144
rect 11683 26104 11692 26144
rect 11732 26104 11741 26144
rect 12547 26104 12556 26144
rect 12596 26104 12844 26144
rect 12884 26104 12893 26144
rect 15043 26104 15052 26144
rect 15092 26104 16396 26144
rect 16436 26104 16972 26144
rect 17012 26104 17021 26144
rect 18979 26104 18988 26144
rect 19028 26104 19372 26144
rect 19412 26104 19421 26144
rect 1507 26103 1565 26104
rect 4972 26060 5012 26104
rect 11692 26060 11732 26104
rect 12259 26060 12317 26061
rect 16195 26060 16253 26061
rect 2500 26020 3724 26060
rect 3764 26020 3773 26060
rect 4972 26020 7372 26060
rect 7412 26020 7421 26060
rect 11692 26020 12268 26060
rect 12308 26020 14996 26060
rect 16110 26020 16204 26060
rect 16244 26020 16253 26060
rect 0 25976 80 25996
rect 2500 25976 2540 26020
rect 12259 26019 12317 26020
rect 14956 25977 14996 26020
rect 16195 26019 16253 26020
rect 16771 26060 16829 26061
rect 16771 26020 16780 26060
rect 16820 26020 19660 26060
rect 19700 26020 19709 26060
rect 16771 26019 16829 26020
rect 14947 25976 15005 25977
rect 21424 25976 21504 25996
rect 0 25936 1940 25976
rect 2371 25936 2380 25976
rect 2420 25936 2540 25976
rect 5155 25936 5164 25976
rect 5204 25936 6508 25976
rect 6548 25936 6557 25976
rect 14947 25936 14956 25976
rect 14996 25936 17164 25976
rect 17204 25936 17836 25976
rect 17876 25936 18796 25976
rect 18836 25936 18845 25976
rect 20227 25936 20236 25976
rect 20276 25936 21504 25976
rect 0 25916 80 25936
rect 1900 25892 1940 25936
rect 14947 25935 15005 25936
rect 21424 25916 21504 25936
rect 1900 25852 2708 25892
rect 2755 25852 2764 25892
rect 2804 25852 3820 25892
rect 3860 25852 3869 25892
rect 14275 25852 14284 25892
rect 14324 25852 15724 25892
rect 15764 25852 15773 25892
rect 16867 25852 16876 25892
rect 16916 25852 17356 25892
rect 17396 25852 18700 25892
rect 18740 25852 18749 25892
rect 2668 25808 2708 25852
rect 15724 25808 15764 25852
rect 1507 25768 1516 25808
rect 1556 25768 2540 25808
rect 2668 25768 8428 25808
rect 8468 25768 8477 25808
rect 15724 25768 19372 25808
rect 19412 25768 19421 25808
rect 2500 25724 2540 25768
rect 5443 25724 5501 25725
rect 15523 25724 15581 25725
rect 2500 25684 3436 25724
rect 3476 25684 3485 25724
rect 3679 25684 3688 25724
rect 3728 25684 3770 25724
rect 3810 25684 3852 25724
rect 3892 25684 3934 25724
rect 3974 25684 4016 25724
rect 4056 25684 4065 25724
rect 5347 25684 5356 25724
rect 5396 25684 5452 25724
rect 5492 25684 12844 25724
rect 12884 25684 12893 25724
rect 13795 25684 13804 25724
rect 13844 25684 14188 25724
rect 14228 25684 14237 25724
rect 15427 25684 15436 25724
rect 15476 25684 15532 25724
rect 15572 25684 15581 25724
rect 18799 25684 18808 25724
rect 18848 25684 18890 25724
rect 18930 25684 18972 25724
rect 19012 25684 19054 25724
rect 19094 25684 19136 25724
rect 19176 25684 19185 25724
rect 19843 25684 19852 25724
rect 19892 25684 21388 25724
rect 21428 25684 21437 25724
rect 5443 25683 5501 25684
rect 15523 25683 15581 25684
rect 0 25640 80 25660
rect 14755 25640 14813 25641
rect 0 25600 1036 25640
rect 1076 25600 1085 25640
rect 2083 25600 2092 25640
rect 2132 25600 4396 25640
rect 4436 25600 4445 25640
rect 11587 25600 11596 25640
rect 11636 25600 12268 25640
rect 12308 25600 12317 25640
rect 14755 25600 14764 25640
rect 14804 25600 14860 25640
rect 14900 25600 14909 25640
rect 15724 25600 17356 25640
rect 17396 25600 17405 25640
rect 0 25580 80 25600
rect 14755 25599 14813 25600
rect 4771 25556 4829 25557
rect 15724 25556 15764 25600
rect 2851 25516 2860 25556
rect 2900 25516 3340 25556
rect 3380 25516 4780 25556
rect 4820 25516 4829 25556
rect 8803 25516 8812 25556
rect 8852 25516 15764 25556
rect 15811 25516 15820 25556
rect 15860 25516 20044 25556
rect 20084 25516 20093 25556
rect 4771 25515 4829 25516
rect 1795 25472 1853 25473
rect 21424 25472 21504 25492
rect 1795 25432 1804 25472
rect 1844 25432 2380 25472
rect 2420 25432 2429 25472
rect 2500 25432 4300 25472
rect 4340 25432 4349 25472
rect 9571 25432 9580 25472
rect 9620 25432 9868 25472
rect 9908 25432 9917 25472
rect 10627 25432 10636 25472
rect 10676 25432 11884 25472
rect 11924 25432 11933 25472
rect 15043 25432 15052 25472
rect 15092 25432 18548 25472
rect 21379 25432 21388 25472
rect 21428 25432 21504 25472
rect 1795 25431 1853 25432
rect 2500 25388 2540 25432
rect 14371 25388 14429 25389
rect 2188 25348 2540 25388
rect 2947 25348 2956 25388
rect 2996 25348 3820 25388
rect 3860 25348 3869 25388
rect 7267 25348 7276 25388
rect 7316 25348 8908 25388
rect 8948 25348 8957 25388
rect 14083 25348 14092 25388
rect 14132 25348 14380 25388
rect 14420 25348 15340 25388
rect 15380 25348 15389 25388
rect 0 25304 80 25324
rect 2188 25304 2228 25348
rect 14371 25347 14429 25348
rect 3235 25304 3293 25305
rect 13315 25304 13373 25305
rect 0 25264 2228 25304
rect 2275 25264 2284 25304
rect 2324 25264 2668 25304
rect 2708 25264 2717 25304
rect 2851 25264 2860 25304
rect 2900 25264 3052 25304
rect 3092 25264 3244 25304
rect 3284 25264 3293 25304
rect 3427 25264 3436 25304
rect 3476 25264 4340 25304
rect 4387 25264 4396 25304
rect 4436 25264 7180 25304
rect 7220 25264 7229 25304
rect 9091 25264 9100 25304
rect 9140 25264 9580 25304
rect 9620 25264 10060 25304
rect 10100 25264 10444 25304
rect 10484 25264 10493 25304
rect 13315 25264 13324 25304
rect 13364 25264 13516 25304
rect 13556 25264 13565 25304
rect 16291 25264 16300 25304
rect 16340 25264 17932 25304
rect 17972 25264 17981 25304
rect 0 25244 80 25264
rect 3235 25263 3293 25264
rect 2371 25220 2429 25221
rect 4003 25220 4061 25221
rect 2371 25180 2380 25220
rect 2420 25180 2764 25220
rect 2804 25180 2813 25220
rect 3918 25180 4012 25220
rect 4052 25180 4061 25220
rect 4300 25220 4340 25264
rect 13315 25263 13373 25264
rect 7747 25220 7805 25221
rect 10147 25220 10205 25221
rect 4300 25180 7756 25220
rect 7796 25180 7805 25220
rect 8035 25180 8044 25220
rect 8084 25180 9484 25220
rect 9524 25180 9533 25220
rect 10062 25180 10156 25220
rect 10196 25180 10205 25220
rect 2371 25179 2429 25180
rect 4003 25179 4061 25180
rect 7747 25179 7805 25180
rect 10147 25179 10205 25180
rect 10339 25220 10397 25221
rect 12355 25220 12413 25221
rect 15619 25220 15677 25221
rect 16579 25220 16637 25221
rect 18508 25220 18548 25432
rect 21424 25412 21504 25432
rect 18883 25348 18892 25388
rect 18932 25348 19660 25388
rect 19700 25348 19709 25388
rect 18691 25264 18700 25304
rect 18740 25264 20044 25304
rect 20084 25264 20093 25304
rect 10339 25180 10348 25220
rect 10388 25180 11020 25220
rect 11060 25180 11069 25220
rect 12270 25180 12364 25220
rect 12404 25180 12413 25220
rect 13603 25180 13612 25220
rect 13652 25180 13900 25220
rect 13940 25180 13949 25220
rect 14371 25180 14380 25220
rect 14420 25180 14860 25220
rect 14900 25180 14909 25220
rect 15043 25180 15052 25220
rect 15092 25180 15572 25220
rect 10339 25179 10397 25180
rect 12355 25179 12413 25180
rect 11779 25136 11837 25137
rect 15532 25136 15572 25180
rect 15619 25180 15628 25220
rect 15668 25180 16588 25220
rect 16628 25180 16637 25220
rect 18019 25180 18028 25220
rect 18068 25180 18412 25220
rect 18452 25180 18461 25220
rect 18508 25180 19180 25220
rect 19220 25180 19796 25220
rect 15619 25179 15677 25180
rect 16579 25179 16637 25180
rect 19756 25136 19796 25180
rect 172 25096 2540 25136
rect 7459 25096 7468 25136
rect 7508 25096 7660 25136
rect 7700 25096 7709 25136
rect 10819 25096 10828 25136
rect 10868 25096 11116 25136
rect 11156 25096 11165 25136
rect 11779 25096 11788 25136
rect 11828 25096 13132 25136
rect 13172 25096 13181 25136
rect 15532 25096 15628 25136
rect 15668 25096 15677 25136
rect 18499 25096 18508 25136
rect 18548 25096 18796 25136
rect 18836 25096 18845 25136
rect 19747 25096 19756 25136
rect 19796 25096 19805 25136
rect 0 24968 80 24988
rect 172 24968 212 25096
rect 2500 25052 2540 25096
rect 11779 25095 11837 25096
rect 17539 25052 17597 25053
rect 2500 25012 17548 25052
rect 17588 25012 17597 25052
rect 17539 25011 17597 25012
rect 21424 24968 21504 24988
rect 0 24928 212 24968
rect 4919 24928 4928 24968
rect 4968 24928 5010 24968
rect 5050 24928 5092 24968
rect 5132 24928 5174 24968
rect 5214 24928 5256 24968
rect 5296 24928 5305 24968
rect 5827 24928 5836 24968
rect 5876 24928 6028 24968
rect 6068 24928 6077 24968
rect 9955 24928 9964 24968
rect 10004 24928 10924 24968
rect 10964 24928 10973 24968
rect 20039 24928 20048 24968
rect 20088 24928 20130 24968
rect 20170 24928 20212 24968
rect 20252 24928 20294 24968
rect 20334 24928 20376 24968
rect 20416 24928 20425 24968
rect 20812 24928 21504 24968
rect 0 24908 80 24928
rect 16387 24884 16445 24885
rect 6403 24844 6412 24884
rect 6452 24844 16396 24884
rect 16436 24844 16445 24884
rect 16387 24843 16445 24844
rect 3331 24800 3389 24801
rect 20812 24800 20852 24928
rect 21424 24908 21504 24928
rect 3331 24760 3340 24800
rect 3380 24760 3532 24800
rect 3572 24760 3581 24800
rect 14563 24760 14572 24800
rect 14612 24760 14621 24800
rect 14755 24760 14764 24800
rect 14804 24760 15340 24800
rect 15380 24760 15389 24800
rect 20227 24760 20236 24800
rect 20276 24760 20852 24800
rect 3331 24759 3389 24760
rect 9955 24716 10013 24717
rect 14572 24716 14612 24760
rect 9955 24676 9964 24716
rect 10004 24676 10060 24716
rect 10100 24676 10109 24716
rect 10723 24676 10732 24716
rect 10772 24676 11692 24716
rect 11732 24676 11741 24716
rect 12067 24676 12076 24716
rect 12116 24676 12125 24716
rect 14572 24676 14996 24716
rect 9955 24675 10013 24676
rect 0 24632 80 24652
rect 5443 24632 5501 24633
rect 12076 24632 12116 24676
rect 14563 24632 14621 24633
rect 14956 24632 14996 24676
rect 16483 24632 16541 24633
rect 19651 24632 19709 24633
rect 0 24592 2036 24632
rect 4579 24592 4588 24632
rect 4628 24592 4780 24632
rect 4820 24592 5452 24632
rect 5492 24592 5501 24632
rect 6115 24592 6124 24632
rect 6164 24592 8332 24632
rect 8372 24592 8381 24632
rect 11203 24592 11212 24632
rect 11252 24592 11884 24632
rect 11924 24592 11933 24632
rect 12076 24592 13900 24632
rect 13940 24592 14420 24632
rect 14478 24592 14572 24632
rect 14612 24592 14621 24632
rect 14947 24592 14956 24632
rect 14996 24592 16300 24632
rect 16340 24592 16349 24632
rect 16483 24592 16492 24632
rect 16532 24592 16588 24632
rect 16628 24592 16637 24632
rect 19171 24592 19180 24632
rect 19220 24592 19660 24632
rect 19700 24592 19709 24632
rect 19843 24592 19852 24632
rect 19892 24592 19901 24632
rect 0 24572 80 24592
rect 1996 24464 2036 24592
rect 5443 24591 5501 24592
rect 2083 24548 2141 24549
rect 7171 24548 7229 24549
rect 13219 24548 13277 24549
rect 2083 24508 2092 24548
rect 2132 24508 7180 24548
rect 7220 24508 7229 24548
rect 8803 24508 8812 24548
rect 8852 24508 9484 24548
rect 9524 24508 9676 24548
rect 9716 24508 9725 24548
rect 13219 24508 13228 24548
rect 13268 24508 13708 24548
rect 13748 24508 13757 24548
rect 2083 24507 2141 24508
rect 7171 24507 7229 24508
rect 13219 24507 13277 24508
rect 14380 24464 14420 24592
rect 14563 24591 14621 24592
rect 16483 24591 16541 24592
rect 19651 24591 19709 24592
rect 19852 24548 19892 24592
rect 14851 24508 14860 24548
rect 14900 24508 16012 24548
rect 16052 24508 16061 24548
rect 16867 24508 16876 24548
rect 16916 24508 17260 24548
rect 17300 24508 17309 24548
rect 18604 24508 19892 24548
rect 18019 24464 18077 24465
rect 18604 24464 18644 24508
rect 21424 24464 21504 24484
rect 1996 24424 2540 24464
rect 6019 24424 6028 24464
rect 6068 24424 6220 24464
rect 6260 24424 6796 24464
rect 6836 24424 7948 24464
rect 7988 24424 7997 24464
rect 8044 24424 10540 24464
rect 10580 24424 10589 24464
rect 13219 24424 13228 24464
rect 13268 24424 13900 24464
rect 13940 24424 13949 24464
rect 14371 24424 14380 24464
rect 14420 24424 14429 24464
rect 18019 24424 18028 24464
rect 18068 24424 18604 24464
rect 18644 24424 18653 24464
rect 19843 24424 19852 24464
rect 19892 24424 21504 24464
rect 2500 24380 2540 24424
rect 8044 24380 8084 24424
rect 18019 24423 18077 24424
rect 21424 24404 21504 24424
rect 11107 24380 11165 24381
rect 2500 24340 8084 24380
rect 8323 24340 8332 24380
rect 8372 24340 11116 24380
rect 11156 24340 11165 24380
rect 11107 24339 11165 24340
rect 13507 24380 13565 24381
rect 13507 24340 13516 24380
rect 13556 24340 14956 24380
rect 14996 24340 15005 24380
rect 13507 24339 13565 24340
rect 0 24296 80 24316
rect 14755 24296 14813 24297
rect 0 24256 6508 24296
rect 6548 24256 9100 24296
rect 9140 24256 9149 24296
rect 14563 24256 14572 24296
rect 14612 24256 14764 24296
rect 14804 24256 14813 24296
rect 0 24236 80 24256
rect 14755 24255 14813 24256
rect 14860 24256 21388 24296
rect 21428 24256 21437 24296
rect 12067 24212 12125 24213
rect 14860 24212 14900 24256
rect 18019 24212 18077 24213
rect 3679 24172 3688 24212
rect 3728 24172 3770 24212
rect 3810 24172 3852 24212
rect 3892 24172 3934 24212
rect 3974 24172 4016 24212
rect 4056 24172 4065 24212
rect 5827 24172 5836 24212
rect 5876 24172 11360 24212
rect 8899 24128 8957 24129
rect 11320 24128 11360 24172
rect 12067 24172 12076 24212
rect 12116 24172 14900 24212
rect 16483 24172 16492 24212
rect 16532 24172 16780 24212
rect 16820 24172 16829 24212
rect 17347 24172 17356 24212
rect 17396 24172 18028 24212
rect 18068 24172 18077 24212
rect 18799 24172 18808 24212
rect 18848 24172 18890 24212
rect 18930 24172 18972 24212
rect 19012 24172 19054 24212
rect 19094 24172 19136 24212
rect 19176 24172 19185 24212
rect 12067 24171 12125 24172
rect 18019 24171 18077 24172
rect 6691 24088 6700 24128
rect 6740 24088 8908 24128
rect 8948 24088 10060 24128
rect 10100 24088 10109 24128
rect 11320 24088 19660 24128
rect 19700 24088 19709 24128
rect 8899 24087 8957 24088
rect 2500 24004 9580 24044
rect 9620 24004 9629 24044
rect 16675 24004 16684 24044
rect 16724 24004 17452 24044
rect 17492 24004 17501 24044
rect 18307 24004 18316 24044
rect 18356 24004 18988 24044
rect 19028 24004 19037 24044
rect 0 23960 80 23980
rect 0 23920 500 23960
rect 0 23900 80 23920
rect 460 23876 500 23920
rect 2500 23876 2540 24004
rect 17347 23960 17405 23961
rect 21424 23960 21504 23980
rect 3523 23920 3532 23960
rect 3572 23920 4012 23960
rect 4052 23920 4061 23960
rect 5251 23920 5260 23960
rect 5300 23920 5452 23960
rect 5492 23920 5501 23960
rect 6595 23920 6604 23960
rect 6644 23920 7564 23960
rect 7604 23920 7613 23960
rect 11395 23920 11404 23960
rect 11444 23920 11596 23960
rect 11636 23920 11645 23960
rect 12643 23920 12652 23960
rect 12692 23920 12701 23960
rect 13315 23920 13324 23960
rect 13364 23920 13708 23960
rect 13748 23920 13757 23960
rect 17347 23920 17356 23960
rect 17396 23920 17548 23960
rect 17588 23920 17597 23960
rect 19267 23920 19276 23960
rect 19316 23920 19660 23960
rect 19700 23920 19709 23960
rect 21379 23920 21388 23960
rect 21428 23920 21504 23960
rect 460 23836 2540 23876
rect 5827 23876 5885 23877
rect 5827 23836 5836 23876
rect 5876 23836 6892 23876
rect 6932 23836 6941 23876
rect 8899 23836 8908 23876
rect 8948 23836 10636 23876
rect 10676 23836 10685 23876
rect 5827 23835 5885 23836
rect 1699 23792 1757 23793
rect 1315 23752 1324 23792
rect 1364 23752 1708 23792
rect 1748 23752 1757 23792
rect 1699 23751 1757 23752
rect 2851 23792 2909 23793
rect 12652 23792 12692 23920
rect 17347 23919 17405 23920
rect 21424 23900 21504 23920
rect 12835 23836 12844 23876
rect 12884 23836 13132 23876
rect 13172 23836 15244 23876
rect 15284 23836 15293 23876
rect 16483 23792 16541 23793
rect 16771 23792 16829 23793
rect 2851 23752 2860 23792
rect 2900 23752 3532 23792
rect 3572 23752 4972 23792
rect 5012 23752 5021 23792
rect 5251 23752 5260 23792
rect 5300 23752 5644 23792
rect 5684 23752 6412 23792
rect 6452 23752 6461 23792
rect 6979 23752 6988 23792
rect 7028 23752 8140 23792
rect 8180 23752 8189 23792
rect 10339 23752 10348 23792
rect 10388 23752 13804 23792
rect 13844 23752 13853 23792
rect 14083 23752 14092 23792
rect 14132 23752 14668 23792
rect 14708 23752 15436 23792
rect 15476 23752 15485 23792
rect 15715 23752 15724 23792
rect 15764 23752 16492 23792
rect 16532 23752 16780 23792
rect 16820 23752 16829 23792
rect 18499 23752 18508 23792
rect 18548 23752 18892 23792
rect 18932 23752 18941 23792
rect 19555 23752 19564 23792
rect 19604 23752 19613 23792
rect 2851 23751 2909 23752
rect 0 23624 80 23644
rect 4972 23624 5012 23752
rect 16483 23751 16541 23752
rect 16771 23751 16829 23752
rect 19564 23708 19604 23752
rect 5539 23668 5548 23708
rect 5588 23668 8044 23708
rect 8084 23668 8093 23708
rect 8419 23668 8428 23708
rect 8468 23668 14188 23708
rect 14228 23668 14237 23708
rect 14851 23668 14860 23708
rect 14900 23668 15532 23708
rect 15572 23668 15581 23708
rect 18403 23668 18412 23708
rect 18452 23668 19604 23708
rect 0 23584 76 23624
rect 116 23584 125 23624
rect 2659 23584 2668 23624
rect 2708 23584 3436 23624
rect 3476 23584 4684 23624
rect 4724 23584 4733 23624
rect 4972 23584 6508 23624
rect 6548 23584 6557 23624
rect 10627 23584 10636 23624
rect 10676 23584 11212 23624
rect 11252 23584 11924 23624
rect 13795 23584 13804 23624
rect 13844 23584 14092 23624
rect 14132 23584 14141 23624
rect 17635 23584 17644 23624
rect 17684 23584 18796 23624
rect 18836 23584 18845 23624
rect 20131 23584 20140 23624
rect 20180 23584 21332 23624
rect 0 23564 80 23584
rect 6499 23540 6557 23541
rect 1699 23500 1708 23540
rect 1748 23500 6124 23540
rect 6164 23500 6173 23540
rect 6499 23500 6508 23540
rect 6548 23500 6604 23540
rect 6644 23500 6653 23540
rect 7660 23500 8840 23540
rect 6124 23456 6164 23500
rect 6499 23499 6557 23500
rect 7171 23456 7229 23457
rect 4919 23416 4928 23456
rect 4968 23416 5010 23456
rect 5050 23416 5092 23456
rect 5132 23416 5174 23456
rect 5214 23416 5256 23456
rect 5296 23416 5305 23456
rect 5635 23416 5644 23456
rect 5684 23416 5836 23456
rect 5876 23416 5885 23456
rect 6124 23416 6988 23456
rect 7028 23416 7037 23456
rect 7086 23416 7180 23456
rect 7220 23416 7229 23456
rect 7171 23415 7229 23416
rect 1699 23372 1757 23373
rect 1699 23332 1708 23372
rect 1748 23332 5548 23372
rect 5588 23332 5597 23372
rect 6403 23332 6412 23372
rect 6452 23332 7564 23372
rect 7604 23332 7613 23372
rect 1699 23331 1757 23332
rect 0 23288 80 23308
rect 7660 23288 7700 23500
rect 8800 23372 8840 23500
rect 11884 23456 11924 23584
rect 18403 23540 18461 23541
rect 12643 23500 12652 23540
rect 12692 23500 14380 23540
rect 14420 23500 14429 23540
rect 18403 23500 18412 23540
rect 18452 23500 18604 23540
rect 18644 23500 18653 23540
rect 18403 23499 18461 23500
rect 16963 23456 17021 23457
rect 18211 23456 18269 23457
rect 21292 23456 21332 23584
rect 21424 23456 21504 23476
rect 11875 23416 11884 23456
rect 11924 23416 16972 23456
rect 17012 23416 17021 23456
rect 18115 23416 18124 23456
rect 18164 23416 18220 23456
rect 18260 23416 18269 23456
rect 20039 23416 20048 23456
rect 20088 23416 20130 23456
rect 20170 23416 20212 23456
rect 20252 23416 20294 23456
rect 20334 23416 20376 23456
rect 20416 23416 20425 23456
rect 21292 23416 21504 23456
rect 16963 23415 17021 23416
rect 18211 23415 18269 23416
rect 21424 23396 21504 23416
rect 13315 23372 13373 23373
rect 13507 23372 13565 23373
rect 8800 23332 13324 23372
rect 13364 23332 13516 23372
rect 13556 23332 13612 23372
rect 13652 23332 13661 23372
rect 15907 23332 15916 23372
rect 15956 23332 16204 23372
rect 16244 23332 16253 23372
rect 17452 23332 17836 23372
rect 17876 23332 17885 23372
rect 13315 23331 13373 23332
rect 13507 23331 13565 23332
rect 0 23248 7700 23288
rect 7747 23288 7805 23289
rect 8419 23288 8477 23289
rect 17059 23288 17117 23289
rect 17452 23288 17492 23332
rect 7747 23248 7756 23288
rect 7796 23248 8140 23288
rect 8180 23248 8428 23288
rect 8468 23248 10772 23288
rect 11491 23248 11500 23288
rect 11540 23248 12076 23288
rect 12116 23248 12125 23288
rect 13516 23248 17068 23288
rect 17108 23248 17492 23288
rect 17539 23248 17548 23288
rect 17588 23248 18124 23288
rect 18164 23248 18173 23288
rect 18499 23248 18508 23288
rect 18548 23248 18740 23288
rect 0 23228 80 23248
rect 7747 23247 7805 23248
rect 8419 23247 8477 23248
rect 4387 23204 4445 23205
rect 4387 23164 4396 23204
rect 4436 23164 7412 23204
rect 7747 23164 7756 23204
rect 7796 23164 8908 23204
rect 8948 23164 9388 23204
rect 9428 23164 9437 23204
rect 9571 23164 9580 23204
rect 9620 23164 9964 23204
rect 10004 23164 10013 23204
rect 4387 23163 4445 23164
rect 4675 23120 4733 23121
rect 2467 23080 2476 23120
rect 2516 23080 2572 23120
rect 2612 23080 4300 23120
rect 4340 23080 4349 23120
rect 4675 23080 4684 23120
rect 4724 23080 4972 23120
rect 5012 23080 5021 23120
rect 4675 23079 4733 23080
rect 7372 23036 7412 23164
rect 10732 23120 10772 23248
rect 13516 23204 13556 23248
rect 17059 23247 17117 23248
rect 18700 23204 18740 23248
rect 11011 23164 11020 23204
rect 11060 23164 13556 23204
rect 17251 23164 17260 23204
rect 17300 23164 17932 23204
rect 17972 23164 17981 23204
rect 18691 23164 18700 23204
rect 18740 23164 19084 23204
rect 19124 23164 19133 23204
rect 7459 23080 7468 23120
rect 7508 23080 7852 23120
rect 7892 23080 8044 23120
rect 8084 23080 10156 23120
rect 10196 23080 10205 23120
rect 10339 23080 10348 23120
rect 10388 23080 10636 23120
rect 10676 23080 10685 23120
rect 10732 23080 13900 23120
rect 13940 23080 13949 23120
rect 14371 23080 14380 23120
rect 14420 23080 15244 23120
rect 15284 23080 16492 23120
rect 16532 23080 16541 23120
rect 17155 23080 17164 23120
rect 17204 23080 17644 23120
rect 17684 23080 17693 23120
rect 19843 23080 19852 23120
rect 19892 23080 19901 23120
rect 10339 23036 10397 23037
rect 19852 23036 19892 23080
rect 4099 22996 4108 23036
rect 4148 22996 5836 23036
rect 5876 22996 5885 23036
rect 6883 22996 6892 23036
rect 6932 22996 7180 23036
rect 7220 22996 7229 23036
rect 7372 22996 8908 23036
rect 8948 22996 9292 23036
rect 9332 22996 9341 23036
rect 10339 22996 10348 23036
rect 10388 22996 19892 23036
rect 10339 22995 10397 22996
rect 0 22952 80 22972
rect 16963 22952 17021 22953
rect 21424 22952 21504 22972
rect 0 22912 1132 22952
rect 1172 22912 1181 22952
rect 2755 22912 2764 22952
rect 2804 22912 3148 22952
rect 3188 22912 8140 22952
rect 8180 22912 8189 22952
rect 16963 22912 16972 22952
rect 17012 22912 17356 22952
rect 17396 22912 18604 22952
rect 18644 22912 18653 22952
rect 18787 22912 18796 22952
rect 18836 22912 21504 22952
rect 0 22892 80 22912
rect 16963 22911 17021 22912
rect 21424 22892 21504 22912
rect 9091 22868 9149 22869
rect 9571 22868 9629 22869
rect 5539 22828 5548 22868
rect 5588 22828 8180 22868
rect 2179 22784 2237 22785
rect 6211 22784 6269 22785
rect 2179 22744 2188 22784
rect 2228 22744 6220 22784
rect 6260 22744 6269 22784
rect 2179 22743 2237 22744
rect 6211 22743 6269 22744
rect 2851 22700 2909 22701
rect 3331 22700 3389 22701
rect 8140 22700 8180 22828
rect 9091 22828 9100 22868
rect 9140 22828 9580 22868
rect 9620 22828 17548 22868
rect 17588 22828 17597 22868
rect 18412 22828 18892 22868
rect 18932 22828 18941 22868
rect 9091 22827 9149 22828
rect 9571 22827 9629 22828
rect 16867 22784 16925 22785
rect 18412 22784 18452 22828
rect 11779 22744 11788 22784
rect 11828 22744 12556 22784
rect 12596 22744 12605 22784
rect 15139 22744 15148 22784
rect 15188 22744 15628 22784
rect 15668 22744 15677 22784
rect 15811 22744 15820 22784
rect 15860 22744 16876 22784
rect 16916 22744 16925 22784
rect 17635 22744 17644 22784
rect 17684 22744 17932 22784
rect 17972 22744 17981 22784
rect 18403 22744 18412 22784
rect 18452 22744 18461 22784
rect 16867 22743 16925 22744
rect 11875 22700 11933 22701
rect 12067 22700 12125 22701
rect 15235 22700 15293 22701
rect 2851 22660 2860 22700
rect 2900 22660 3052 22700
rect 3092 22660 3340 22700
rect 3380 22660 3389 22700
rect 3679 22660 3688 22700
rect 3728 22660 3770 22700
rect 3810 22660 3852 22700
rect 3892 22660 3934 22700
rect 3974 22660 4016 22700
rect 4056 22660 4065 22700
rect 4195 22660 4204 22700
rect 4244 22660 6316 22700
rect 6356 22660 6365 22700
rect 6499 22660 6508 22700
rect 6548 22660 7084 22700
rect 7124 22660 7133 22700
rect 7555 22660 7564 22700
rect 7604 22660 8044 22700
rect 8084 22660 8093 22700
rect 8140 22660 10348 22700
rect 10388 22660 10397 22700
rect 11875 22660 11884 22700
rect 11924 22660 12076 22700
rect 12116 22660 12125 22700
rect 14467 22660 14476 22700
rect 14516 22660 15244 22700
rect 15284 22660 15293 22700
rect 2851 22659 2909 22660
rect 3331 22659 3389 22660
rect 11875 22659 11933 22660
rect 12067 22659 12125 22660
rect 15235 22659 15293 22660
rect 16387 22700 16445 22701
rect 16387 22660 16396 22700
rect 16436 22660 18356 22700
rect 18799 22660 18808 22700
rect 18848 22660 18890 22700
rect 18930 22660 18972 22700
rect 19012 22660 19054 22700
rect 19094 22660 19136 22700
rect 19176 22660 19185 22700
rect 16387 22659 16445 22660
rect 0 22616 80 22636
rect 2371 22616 2429 22617
rect 7171 22616 7229 22617
rect 0 22576 2380 22616
rect 2420 22576 2429 22616
rect 2851 22576 2860 22616
rect 2900 22576 5740 22616
rect 5780 22576 5789 22616
rect 5923 22576 5932 22616
rect 5972 22576 7180 22616
rect 7220 22576 7852 22616
rect 7892 22576 7901 22616
rect 10531 22576 10540 22616
rect 10580 22576 18220 22616
rect 18260 22576 18269 22616
rect 0 22556 80 22576
rect 2371 22575 2429 22576
rect 7171 22575 7229 22576
rect 4291 22532 4349 22533
rect 6307 22532 6365 22533
rect 11011 22532 11069 22533
rect 18211 22532 18269 22533
rect 4291 22492 4300 22532
rect 4340 22492 6316 22532
rect 6356 22492 9292 22532
rect 9332 22492 9341 22532
rect 9388 22492 11020 22532
rect 11060 22492 17780 22532
rect 18019 22492 18028 22532
rect 18068 22492 18220 22532
rect 18260 22492 18269 22532
rect 18316 22532 18356 22660
rect 18316 22492 20180 22532
rect 4291 22491 4349 22492
rect 6307 22491 6365 22492
rect 4483 22408 4492 22448
rect 4532 22408 6452 22448
rect 6499 22408 6508 22448
rect 6548 22408 6796 22448
rect 6836 22408 6845 22448
rect 6979 22408 6988 22448
rect 7028 22408 8521 22448
rect 8561 22408 8716 22448
rect 8756 22408 8765 22448
rect 3139 22364 3197 22365
rect 6412 22364 6452 22408
rect 9388 22364 9428 22492
rect 11011 22491 11069 22492
rect 9763 22408 9772 22448
rect 9812 22408 10580 22448
rect 11395 22408 11404 22448
rect 11444 22408 12556 22448
rect 12596 22408 12605 22448
rect 3139 22324 3148 22364
rect 3188 22324 5068 22364
rect 5108 22324 5117 22364
rect 6412 22324 9428 22364
rect 3139 22323 3197 22324
rect 0 22280 80 22300
rect 1891 22280 1949 22281
rect 2371 22280 2429 22281
rect 6499 22280 6557 22281
rect 10540 22280 10580 22408
rect 11011 22364 11069 22365
rect 13507 22364 13565 22365
rect 15523 22364 15581 22365
rect 11011 22324 11020 22364
rect 11060 22324 11308 22364
rect 11348 22324 11357 22364
rect 11491 22324 11500 22364
rect 11540 22324 11692 22364
rect 11732 22324 11741 22364
rect 13507 22324 13516 22364
rect 13556 22324 13708 22364
rect 13748 22324 13757 22364
rect 15331 22324 15340 22364
rect 15380 22324 15532 22364
rect 15572 22324 15581 22364
rect 11011 22323 11069 22324
rect 13507 22323 13565 22324
rect 15523 22323 15581 22324
rect 15907 22280 15965 22281
rect 16099 22280 16157 22281
rect 17740 22280 17780 22492
rect 18211 22491 18269 22492
rect 20140 22448 20180 22492
rect 21424 22448 21504 22468
rect 18883 22408 18892 22448
rect 18932 22408 19468 22448
rect 19508 22408 19517 22448
rect 19651 22408 19660 22448
rect 19700 22408 19948 22448
rect 19988 22408 19997 22448
rect 20140 22408 21504 22448
rect 21424 22388 21504 22408
rect 0 22240 1900 22280
rect 1940 22240 2380 22280
rect 2420 22240 2429 22280
rect 2563 22240 2572 22280
rect 2612 22240 4012 22280
rect 4052 22240 4684 22280
rect 4724 22240 4733 22280
rect 6499 22240 6508 22280
rect 6548 22240 8620 22280
rect 8660 22240 8669 22280
rect 9283 22240 9292 22280
rect 9332 22240 10156 22280
rect 10196 22240 10205 22280
rect 10540 22240 11980 22280
rect 12020 22240 12029 22280
rect 13219 22240 13228 22280
rect 13268 22240 14380 22280
rect 14420 22240 14429 22280
rect 14755 22240 14764 22280
rect 14804 22240 15244 22280
rect 15284 22240 15293 22280
rect 15822 22240 15916 22280
rect 15956 22240 15965 22280
rect 16014 22240 16108 22280
rect 16148 22240 16157 22280
rect 16387 22240 16396 22280
rect 16436 22240 17260 22280
rect 17300 22240 17309 22280
rect 17731 22240 17740 22280
rect 17780 22240 17932 22280
rect 17972 22240 17981 22280
rect 18211 22240 18220 22280
rect 18260 22240 18508 22280
rect 18548 22240 18557 22280
rect 19171 22240 19180 22280
rect 19220 22240 19948 22280
rect 19988 22240 19997 22280
rect 0 22220 80 22240
rect 1891 22239 1949 22240
rect 2371 22239 2429 22240
rect 6499 22239 6557 22240
rect 14380 22196 14420 22240
rect 15907 22239 15965 22240
rect 16099 22239 16157 22240
rect 3619 22156 3628 22196
rect 3668 22156 7180 22196
rect 7220 22156 7229 22196
rect 14380 22156 15436 22196
rect 15476 22156 15485 22196
rect 7180 22112 7220 22156
rect 20707 22112 20765 22113
rect 2284 22072 4492 22112
rect 4532 22072 4541 22112
rect 7180 22072 7948 22112
rect 7988 22072 8620 22112
rect 8660 22072 8669 22112
rect 12259 22072 12268 22112
rect 12308 22072 20716 22112
rect 20756 22072 20765 22112
rect 0 21944 80 21964
rect 2284 21944 2324 22072
rect 20707 22071 20765 22072
rect 2371 22028 2429 22029
rect 2371 21988 2380 22028
rect 2420 21988 11596 22028
rect 11636 21988 11645 22028
rect 13987 21988 13996 22028
rect 14036 21988 14284 22028
rect 14324 21988 14333 22028
rect 2371 21987 2429 21988
rect 0 21904 2324 21944
rect 3235 21944 3293 21945
rect 4483 21944 4541 21945
rect 21424 21944 21504 21964
rect 3235 21904 3244 21944
rect 3284 21904 3724 21944
rect 3764 21904 4492 21944
rect 4532 21904 4541 21944
rect 4919 21904 4928 21944
rect 4968 21904 5010 21944
rect 5050 21904 5092 21944
rect 5132 21904 5174 21944
rect 5214 21904 5256 21944
rect 5296 21904 5305 21944
rect 20039 21904 20048 21944
rect 20088 21904 20130 21944
rect 20170 21904 20212 21944
rect 20252 21904 20294 21944
rect 20334 21904 20376 21944
rect 20416 21904 20425 21944
rect 20803 21904 20812 21944
rect 20852 21904 21504 21944
rect 0 21884 80 21904
rect 3235 21903 3293 21904
rect 4483 21903 4541 21904
rect 21424 21884 21504 21904
rect 5731 21860 5789 21861
rect 16771 21860 16829 21861
rect 3235 21820 3244 21860
rect 3284 21820 5684 21860
rect 5644 21776 5684 21820
rect 5731 21820 5740 21860
rect 5780 21820 9004 21860
rect 9044 21820 12556 21860
rect 12596 21820 16780 21860
rect 16820 21820 16829 21860
rect 5731 21819 5789 21820
rect 16771 21819 16829 21820
rect 18019 21860 18077 21861
rect 18019 21820 18028 21860
rect 18068 21820 18124 21860
rect 18164 21820 18173 21860
rect 18019 21819 18077 21820
rect 7075 21776 7133 21777
rect 12067 21776 12125 21777
rect 5644 21736 6028 21776
rect 6068 21736 6077 21776
rect 6691 21736 6700 21776
rect 6740 21736 6749 21776
rect 7075 21736 7084 21776
rect 7124 21736 7276 21776
rect 7316 21736 7325 21776
rect 12067 21736 12076 21776
rect 12116 21736 18700 21776
rect 18740 21736 18749 21776
rect 6499 21692 6557 21693
rect 844 21652 6508 21692
rect 6548 21652 6557 21692
rect 0 21608 80 21628
rect 844 21608 884 21652
rect 6499 21651 6557 21652
rect 0 21568 884 21608
rect 931 21568 940 21608
rect 980 21568 1228 21608
rect 1268 21568 1277 21608
rect 2659 21568 2668 21608
rect 2708 21568 2956 21608
rect 2996 21568 3148 21608
rect 3188 21568 4588 21608
rect 4628 21568 4637 21608
rect 5059 21568 5068 21608
rect 5108 21568 5932 21608
rect 5972 21568 5981 21608
rect 0 21548 80 21568
rect 6700 21524 6740 21736
rect 7075 21735 7133 21736
rect 12067 21735 12125 21736
rect 7363 21692 7421 21693
rect 7278 21652 7372 21692
rect 7412 21652 7421 21692
rect 7363 21651 7421 21652
rect 12643 21692 12701 21693
rect 12643 21652 12652 21692
rect 12692 21652 12748 21692
rect 12788 21652 12797 21692
rect 17155 21652 17164 21692
rect 17204 21652 17548 21692
rect 17588 21652 18412 21692
rect 18452 21652 18461 21692
rect 12643 21651 12701 21652
rect 16099 21608 16157 21609
rect 19939 21608 19997 21609
rect 7075 21568 7084 21608
rect 7124 21568 7852 21608
rect 7892 21568 7901 21608
rect 11587 21568 11596 21608
rect 11636 21568 14572 21608
rect 14612 21568 14621 21608
rect 14947 21568 14956 21608
rect 14996 21568 15532 21608
rect 15572 21568 15581 21608
rect 16014 21568 16108 21608
rect 16148 21568 16157 21608
rect 17827 21568 17836 21608
rect 17876 21568 18508 21608
rect 18548 21568 18557 21608
rect 19854 21568 19948 21608
rect 19988 21568 19997 21608
rect 16099 21567 16157 21568
rect 19939 21567 19997 21568
rect 15523 21524 15581 21525
rect 2563 21484 2572 21524
rect 2612 21484 3340 21524
rect 3380 21484 3389 21524
rect 3628 21484 4340 21524
rect 5539 21484 5548 21524
rect 5588 21484 6508 21524
rect 6548 21484 7276 21524
rect 7316 21484 7325 21524
rect 7651 21484 7660 21524
rect 7700 21484 9484 21524
rect 9524 21484 9533 21524
rect 12067 21484 12076 21524
rect 12116 21484 15532 21524
rect 15572 21484 15628 21524
rect 15668 21484 15677 21524
rect 3628 21440 3668 21484
rect 2755 21400 2764 21440
rect 2804 21400 3668 21440
rect 3715 21400 3724 21440
rect 3764 21400 4204 21440
rect 4244 21400 4253 21440
rect 4300 21356 4340 21484
rect 15523 21483 15581 21484
rect 9475 21440 9533 21441
rect 6115 21400 6124 21440
rect 6164 21400 6604 21440
rect 6644 21400 6653 21440
rect 6883 21400 6892 21440
rect 6932 21400 9484 21440
rect 9524 21400 9533 21440
rect 9475 21399 9533 21400
rect 9667 21440 9725 21441
rect 12739 21440 12797 21441
rect 9667 21400 9676 21440
rect 9716 21400 10156 21440
rect 10196 21400 10205 21440
rect 10531 21400 10540 21440
rect 10580 21400 12748 21440
rect 12788 21400 12797 21440
rect 9667 21399 9725 21400
rect 10540 21356 10580 21400
rect 12739 21399 12797 21400
rect 13603 21440 13661 21441
rect 19267 21440 19325 21441
rect 21424 21440 21504 21460
rect 13603 21400 13612 21440
rect 13652 21400 14668 21440
rect 14708 21400 14717 21440
rect 15907 21400 15916 21440
rect 15956 21400 19276 21440
rect 19316 21400 19325 21440
rect 19843 21400 19852 21440
rect 19892 21400 21504 21440
rect 13603 21399 13661 21400
rect 19267 21399 19325 21400
rect 21424 21380 21504 21400
rect 3523 21316 3532 21356
rect 3572 21316 3916 21356
rect 3956 21316 3965 21356
rect 4300 21316 7084 21356
rect 7124 21316 7133 21356
rect 7363 21316 7372 21356
rect 7412 21316 7660 21356
rect 7700 21316 7709 21356
rect 9859 21316 9868 21356
rect 9908 21316 10580 21356
rect 0 21272 80 21292
rect 4483 21272 4541 21273
rect 11683 21272 11741 21273
rect 16963 21272 17021 21273
rect 0 21232 2540 21272
rect 4195 21232 4204 21272
rect 4244 21232 4492 21272
rect 4532 21232 4541 21272
rect 0 21212 80 21232
rect 2500 21104 2540 21232
rect 4483 21231 4541 21232
rect 6316 21232 8716 21272
rect 8756 21232 8765 21272
rect 11683 21232 11692 21272
rect 11732 21232 16972 21272
rect 17012 21232 17021 21272
rect 3679 21148 3688 21188
rect 3728 21148 3770 21188
rect 3810 21148 3852 21188
rect 3892 21148 3934 21188
rect 3974 21148 4016 21188
rect 4056 21148 4065 21188
rect 6316 21104 6356 21232
rect 11683 21231 11741 21232
rect 16963 21231 17021 21232
rect 9667 21188 9725 21189
rect 6403 21148 6412 21188
rect 6452 21148 6461 21188
rect 6691 21148 6700 21188
rect 6740 21148 6892 21188
rect 6932 21148 6941 21188
rect 7075 21148 7084 21188
rect 7124 21148 9676 21188
rect 9716 21148 9725 21188
rect 11587 21148 11596 21188
rect 11636 21148 13612 21188
rect 13652 21148 13661 21188
rect 14947 21148 14956 21188
rect 14996 21148 15244 21188
rect 15284 21148 15293 21188
rect 18799 21148 18808 21188
rect 18848 21148 18890 21188
rect 18930 21148 18972 21188
rect 19012 21148 19054 21188
rect 19094 21148 19136 21188
rect 19176 21148 19185 21188
rect 2500 21064 6356 21104
rect 4099 21020 4157 21021
rect 6211 21020 6269 21021
rect 1219 20980 1228 21020
rect 1268 20980 4108 21020
rect 4148 20980 4157 21020
rect 5731 20980 5740 21020
rect 5780 20980 6220 21020
rect 6260 20980 6269 21020
rect 4099 20979 4157 20980
rect 6211 20979 6269 20980
rect 0 20936 80 20956
rect 6307 20936 6365 20937
rect 0 20896 2764 20936
rect 2804 20896 2813 20936
rect 3043 20896 3052 20936
rect 3092 20896 3101 20936
rect 3235 20896 3244 20936
rect 3284 20896 3572 20936
rect 0 20876 80 20896
rect 3052 20852 3092 20896
rect 3532 20852 3572 20896
rect 4588 20896 4684 20936
rect 4724 20896 4733 20936
rect 5635 20896 5644 20936
rect 5684 20896 6316 20936
rect 6356 20896 6365 20936
rect 1123 20812 1132 20852
rect 1172 20812 2956 20852
rect 2996 20812 3005 20852
rect 3052 20812 3476 20852
rect 3523 20812 3532 20852
rect 3572 20812 3581 20852
rect 3436 20768 3476 20812
rect 4588 20768 4628 20896
rect 6307 20895 6365 20896
rect 4771 20852 4829 20853
rect 6412 20852 6452 21148
rect 9667 21147 9725 21148
rect 12259 21064 12268 21104
rect 12308 21064 16108 21104
rect 16148 21064 16157 21104
rect 17347 21064 17356 21104
rect 17396 21064 17740 21104
rect 17780 21064 17789 21104
rect 17356 21020 17396 21064
rect 13411 20980 13420 21020
rect 13460 20980 13612 21020
rect 13652 20980 13661 21020
rect 14179 20980 14188 21020
rect 14228 20980 14572 21020
rect 14612 20980 15148 21020
rect 15188 20980 17396 21020
rect 21424 20936 21504 20956
rect 12355 20896 12364 20936
rect 12404 20896 21504 20936
rect 21424 20876 21504 20896
rect 7363 20852 7421 20853
rect 4771 20812 4780 20852
rect 4820 20812 5068 20852
rect 5108 20812 5117 20852
rect 5731 20812 5740 20852
rect 5780 20812 6028 20852
rect 6068 20812 6700 20852
rect 6740 20812 6749 20852
rect 6793 20812 6802 20852
rect 6842 20812 7372 20852
rect 7412 20812 7421 20852
rect 4771 20811 4829 20812
rect 7363 20811 7421 20812
rect 19180 20812 19756 20852
rect 19796 20812 19805 20852
rect 6211 20768 6269 20769
rect 12739 20768 12797 20769
rect 14179 20768 14237 20769
rect 1219 20728 1228 20768
rect 1268 20728 1612 20768
rect 1652 20728 1661 20768
rect 2659 20728 2668 20768
rect 2708 20728 3052 20768
rect 3092 20728 3101 20768
rect 3436 20728 3628 20768
rect 3668 20728 3677 20768
rect 3811 20728 3820 20768
rect 3860 20728 4204 20768
rect 4244 20728 4253 20768
rect 4588 20728 5644 20768
rect 5684 20728 5693 20768
rect 6211 20728 6220 20768
rect 6260 20728 7084 20768
rect 7124 20728 7133 20768
rect 11299 20728 11308 20768
rect 11348 20728 12268 20768
rect 12308 20728 12317 20768
rect 12547 20728 12556 20768
rect 12596 20728 12748 20768
rect 12788 20728 12797 20768
rect 13315 20728 13324 20768
rect 13364 20728 14188 20768
rect 14228 20728 14237 20768
rect 18115 20728 18124 20768
rect 18164 20728 18412 20768
rect 18452 20728 18461 20768
rect 4588 20684 4628 20728
rect 6211 20727 6269 20728
rect 12739 20727 12797 20728
rect 14179 20727 14237 20728
rect 8323 20684 8381 20685
rect 16579 20684 16637 20685
rect 3340 20644 4628 20684
rect 6979 20644 6988 20684
rect 7028 20644 8140 20684
rect 8180 20644 8332 20684
rect 8372 20644 8381 20684
rect 0 20600 80 20620
rect 3340 20600 3380 20644
rect 8323 20643 8381 20644
rect 9580 20644 11116 20684
rect 11156 20644 11165 20684
rect 12931 20644 12940 20684
rect 12980 20644 16588 20684
rect 16628 20644 16637 20684
rect 9580 20600 9620 20644
rect 16579 20643 16637 20644
rect 19180 20600 19220 20812
rect 19555 20728 19564 20768
rect 19604 20728 19948 20768
rect 19988 20728 19997 20768
rect 0 20560 2540 20600
rect 3331 20560 3340 20600
rect 3380 20560 3389 20600
rect 3907 20560 3916 20600
rect 3956 20560 9620 20600
rect 9667 20560 9676 20600
rect 9716 20560 11980 20600
rect 12020 20560 12029 20600
rect 14755 20560 14764 20600
rect 14804 20560 15148 20600
rect 15188 20560 15197 20600
rect 19171 20560 19180 20600
rect 19220 20560 19229 20600
rect 19747 20560 19756 20600
rect 19796 20560 20140 20600
rect 20180 20560 20189 20600
rect 0 20540 80 20560
rect 2500 20516 2540 20560
rect 2500 20476 11360 20516
rect 12163 20476 12172 20516
rect 12212 20476 20852 20516
rect 11320 20432 11360 20476
rect 20812 20432 20852 20476
rect 21424 20432 21504 20452
rect 4919 20392 4928 20432
rect 4968 20392 5010 20432
rect 5050 20392 5092 20432
rect 5132 20392 5174 20432
rect 5214 20392 5256 20432
rect 5296 20392 5305 20432
rect 6115 20392 6124 20432
rect 6164 20392 8428 20432
rect 8468 20392 8477 20432
rect 11320 20392 11596 20432
rect 11636 20392 11645 20432
rect 16396 20392 17452 20432
rect 17492 20392 17501 20432
rect 20039 20392 20048 20432
rect 20088 20392 20130 20432
rect 20170 20392 20212 20432
rect 20252 20392 20294 20432
rect 20334 20392 20376 20432
rect 20416 20392 20425 20432
rect 20812 20392 21504 20432
rect 5539 20348 5597 20349
rect 5539 20308 5548 20348
rect 5588 20308 11360 20348
rect 14755 20308 14764 20348
rect 14804 20308 15052 20348
rect 15092 20308 15101 20348
rect 5539 20307 5597 20308
rect 0 20264 80 20284
rect 11320 20264 11360 20308
rect 16396 20264 16436 20392
rect 21424 20372 21504 20392
rect 0 20224 2284 20264
rect 2324 20224 2333 20264
rect 2659 20224 2668 20264
rect 2708 20224 4108 20264
rect 4148 20224 5836 20264
rect 5876 20224 5885 20264
rect 10627 20224 10636 20264
rect 10676 20224 11252 20264
rect 11320 20224 16436 20264
rect 16483 20224 16492 20264
rect 16532 20224 16541 20264
rect 0 20204 80 20224
rect 11011 20180 11069 20181
rect 11212 20180 11252 20224
rect 11395 20180 11453 20181
rect 14083 20180 14141 20181
rect 15907 20180 15965 20181
rect 1123 20140 1132 20180
rect 1172 20140 3916 20180
rect 3956 20140 3965 20180
rect 4387 20140 4396 20180
rect 4436 20140 5932 20180
rect 5972 20140 5981 20180
rect 10212 20140 10252 20180
rect 10292 20140 10301 20180
rect 11011 20140 11020 20180
rect 11060 20140 11116 20180
rect 11156 20140 11165 20180
rect 11212 20140 11404 20180
rect 11444 20140 11453 20180
rect 13998 20140 14092 20180
rect 14132 20140 14141 20180
rect 15043 20140 15052 20180
rect 15092 20140 15916 20180
rect 15956 20140 15965 20180
rect 2851 20096 2909 20097
rect 9763 20096 9821 20097
rect 10252 20096 10292 20140
rect 11011 20139 11069 20140
rect 11395 20139 11453 20140
rect 14083 20139 14141 20140
rect 15907 20139 15965 20140
rect 2766 20056 2860 20096
rect 2900 20056 2909 20096
rect 4195 20056 4204 20096
rect 4244 20056 5260 20096
rect 5300 20056 5309 20096
rect 5539 20056 5548 20096
rect 5588 20056 6796 20096
rect 6836 20056 6845 20096
rect 7363 20056 7372 20096
rect 7412 20056 7756 20096
rect 7796 20056 7805 20096
rect 9763 20056 9772 20096
rect 9812 20056 10292 20096
rect 11875 20096 11933 20097
rect 16387 20096 16445 20097
rect 16492 20096 16532 20224
rect 16644 20140 16684 20180
rect 16724 20140 16733 20180
rect 19555 20140 19564 20180
rect 19604 20140 19613 20180
rect 11875 20056 11884 20096
rect 11924 20056 12748 20096
rect 12788 20056 12797 20096
rect 14371 20056 14380 20096
rect 14420 20056 14860 20096
rect 14900 20056 14909 20096
rect 16387 20056 16396 20096
rect 16436 20056 16532 20096
rect 16684 20096 16724 20140
rect 19459 20096 19517 20097
rect 16684 20056 18124 20096
rect 18164 20056 18173 20096
rect 18403 20056 18412 20096
rect 18452 20056 18892 20096
rect 18932 20056 18941 20096
rect 19171 20056 19180 20096
rect 19220 20056 19468 20096
rect 19508 20056 19517 20096
rect 2851 20055 2909 20056
rect 9763 20055 9821 20056
rect 11875 20055 11933 20056
rect 16387 20055 16445 20056
rect 19459 20055 19517 20056
rect 14083 20012 14141 20013
rect 19564 20012 19604 20140
rect 19939 20096 19997 20097
rect 19854 20056 19948 20096
rect 19988 20056 19997 20096
rect 19939 20055 19997 20056
rect 2467 19972 2476 20012
rect 2516 19972 4012 20012
rect 4052 19972 4061 20012
rect 4291 19972 4300 20012
rect 4340 19972 4684 20012
rect 4724 19972 4733 20012
rect 6211 19972 6220 20012
rect 6260 19972 6892 20012
rect 6932 19972 6941 20012
rect 11875 19972 11884 20012
rect 11924 19972 13364 20012
rect 13891 19972 13900 20012
rect 13940 19972 14092 20012
rect 14132 19972 14141 20012
rect 17347 19972 17356 20012
rect 17396 19972 17932 20012
rect 17972 19972 19604 20012
rect 0 19928 80 19948
rect 1795 19928 1853 19929
rect 13324 19928 13364 19972
rect 14083 19971 14141 19972
rect 21424 19928 21504 19948
rect 0 19888 1804 19928
rect 1844 19888 1853 19928
rect 11491 19888 11500 19928
rect 11540 19888 12172 19928
rect 12212 19888 13228 19928
rect 13268 19888 13277 19928
rect 13324 19888 16396 19928
rect 16436 19888 16445 19928
rect 21283 19888 21292 19928
rect 21332 19888 21504 19928
rect 0 19868 80 19888
rect 1795 19887 1853 19888
rect 21424 19868 21504 19888
rect 6211 19844 6269 19845
rect 7075 19844 7133 19845
rect 4099 19804 4108 19844
rect 4148 19804 4157 19844
rect 4771 19804 4780 19844
rect 4820 19804 5932 19844
rect 5972 19804 5981 19844
rect 6126 19804 6220 19844
rect 6260 19804 6269 19844
rect 6787 19804 6796 19844
rect 6836 19804 7084 19844
rect 7124 19804 7133 19844
rect 4108 19760 4148 19804
rect 6211 19803 6269 19804
rect 7075 19803 7133 19804
rect 10147 19844 10205 19845
rect 10147 19804 10156 19844
rect 10196 19804 11596 19844
rect 11636 19804 11645 19844
rect 12067 19804 12076 19844
rect 12116 19804 18220 19844
rect 18260 19804 18269 19844
rect 10147 19803 10205 19804
rect 13219 19760 13277 19761
rect 16387 19760 16445 19761
rect 4108 19720 4876 19760
rect 4916 19720 7660 19760
rect 7700 19720 7709 19760
rect 13134 19720 13228 19760
rect 13268 19720 13277 19760
rect 13987 19720 13996 19760
rect 14036 19720 14420 19760
rect 16302 19720 16396 19760
rect 16436 19720 16445 19760
rect 13219 19719 13277 19720
rect 8899 19676 8957 19677
rect 13891 19676 13949 19677
rect 14380 19676 14420 19720
rect 16387 19719 16445 19720
rect 16483 19676 16541 19677
rect 1219 19636 1228 19676
rect 1268 19636 3572 19676
rect 3679 19636 3688 19676
rect 3728 19636 3770 19676
rect 3810 19636 3852 19676
rect 3892 19636 3934 19676
rect 3974 19636 4016 19676
rect 4056 19636 4065 19676
rect 6307 19636 6316 19676
rect 6356 19636 8908 19676
rect 8948 19636 9292 19676
rect 9332 19636 9484 19676
rect 9524 19636 9533 19676
rect 13891 19636 13900 19676
rect 13940 19636 14092 19676
rect 14132 19636 14141 19676
rect 14371 19636 14380 19676
rect 14420 19636 14429 19676
rect 16398 19636 16492 19676
rect 16532 19636 16541 19676
rect 18799 19636 18808 19676
rect 18848 19636 18890 19676
rect 18930 19636 18972 19676
rect 19012 19636 19054 19676
rect 19094 19636 19136 19676
rect 19176 19636 19185 19676
rect 19267 19636 19276 19676
rect 19316 19636 19852 19676
rect 19892 19636 19901 19676
rect 0 19592 80 19612
rect 0 19552 1132 19592
rect 1172 19552 1181 19592
rect 0 19532 80 19552
rect 3532 19508 3572 19636
rect 8899 19635 8957 19636
rect 13891 19635 13949 19636
rect 16483 19635 16541 19636
rect 5827 19592 5885 19593
rect 4387 19552 4396 19592
rect 4436 19552 4972 19592
rect 5012 19552 5021 19592
rect 5827 19552 5836 19592
rect 5876 19552 17164 19592
rect 17204 19552 17213 19592
rect 19555 19552 19564 19592
rect 19604 19552 20140 19592
rect 20180 19552 20189 19592
rect 5827 19551 5885 19552
rect 19267 19508 19325 19509
rect 3532 19468 9580 19508
rect 9620 19468 9629 19508
rect 11320 19468 12076 19508
rect 12116 19468 16492 19508
rect 16532 19468 16541 19508
rect 19267 19468 19276 19508
rect 19316 19468 20756 19508
rect 4099 19424 4157 19425
rect 11320 19424 11360 19468
rect 19267 19467 19325 19468
rect 20716 19424 20756 19468
rect 21424 19424 21504 19444
rect 4099 19384 4108 19424
rect 4148 19384 9196 19424
rect 9236 19384 11360 19424
rect 15811 19384 15820 19424
rect 15860 19384 16300 19424
rect 16340 19384 16349 19424
rect 19084 19384 19948 19424
rect 19988 19384 19997 19424
rect 20227 19384 20236 19424
rect 20276 19384 20620 19424
rect 20660 19384 20669 19424
rect 20716 19384 21504 19424
rect 4099 19383 4157 19384
rect 12259 19340 12317 19341
rect 4387 19300 4396 19340
rect 4436 19300 4780 19340
rect 4820 19300 4829 19340
rect 8803 19300 8812 19340
rect 8852 19300 9100 19340
rect 9140 19300 9149 19340
rect 10531 19300 10540 19340
rect 10580 19300 11308 19340
rect 11348 19300 12268 19340
rect 12308 19300 12364 19340
rect 12404 19300 12413 19340
rect 14275 19300 14284 19340
rect 14324 19300 15148 19340
rect 15188 19300 16108 19340
rect 16148 19300 16972 19340
rect 17012 19300 17021 19340
rect 12259 19299 12317 19300
rect 0 19256 80 19276
rect 1603 19256 1661 19257
rect 5827 19256 5885 19257
rect 14563 19256 14621 19257
rect 19084 19256 19124 19384
rect 21424 19364 21504 19384
rect 0 19216 1612 19256
rect 1652 19216 1661 19256
rect 1795 19216 1804 19256
rect 1844 19216 2572 19256
rect 2612 19216 2621 19256
rect 2755 19216 2764 19256
rect 2804 19216 3532 19256
rect 3572 19216 3581 19256
rect 4579 19216 4588 19256
rect 4628 19216 4876 19256
rect 4916 19216 4925 19256
rect 5742 19216 5836 19256
rect 5876 19216 5885 19256
rect 6307 19216 6316 19256
rect 6356 19216 7468 19256
rect 7508 19216 12308 19256
rect 14478 19216 14572 19256
rect 14612 19216 14621 19256
rect 15523 19216 15532 19256
rect 15572 19216 15724 19256
rect 15764 19216 15773 19256
rect 17731 19216 17740 19256
rect 17780 19216 19084 19256
rect 19124 19216 19133 19256
rect 0 19196 80 19216
rect 1603 19215 1661 19216
rect 5827 19215 5885 19216
rect 2851 19172 2909 19173
rect 5443 19172 5501 19173
rect 8323 19172 8381 19173
rect 11683 19172 11741 19173
rect 2851 19132 2860 19172
rect 2900 19132 3284 19172
rect 2851 19131 2909 19132
rect 3244 19088 3284 19132
rect 5443 19132 5452 19172
rect 5492 19132 6548 19172
rect 8238 19132 8332 19172
rect 8372 19132 8381 19172
rect 10339 19132 10348 19172
rect 10388 19132 11116 19172
rect 11156 19132 11692 19172
rect 11732 19132 11741 19172
rect 12268 19172 12308 19216
rect 14563 19215 14621 19216
rect 17347 19172 17405 19173
rect 12268 19132 17356 19172
rect 17396 19132 17405 19172
rect 5443 19131 5501 19132
rect 6508 19088 6548 19132
rect 8323 19131 8381 19132
rect 11683 19131 11741 19132
rect 17347 19131 17405 19132
rect 9955 19088 10013 19089
rect 2179 19048 2188 19088
rect 2228 19048 3148 19088
rect 3188 19048 3197 19088
rect 3244 19048 6316 19088
rect 6356 19048 6365 19088
rect 6499 19048 6508 19088
rect 6548 19048 9292 19088
rect 9332 19048 9341 19088
rect 9870 19048 9964 19088
rect 10004 19048 10013 19088
rect 10531 19048 10540 19088
rect 10580 19048 17836 19088
rect 17876 19048 19660 19088
rect 19700 19048 19709 19088
rect 9955 19047 10013 19048
rect 940 18964 1708 19004
rect 1748 18964 1757 19004
rect 5635 18964 5644 19004
rect 5684 18964 20564 19004
rect 0 18920 80 18940
rect 940 18920 980 18964
rect 6019 18920 6077 18921
rect 12067 18920 12125 18921
rect 19459 18920 19517 18921
rect 20524 18920 20564 18964
rect 21424 18920 21504 18940
rect 0 18880 980 18920
rect 1027 18880 1036 18920
rect 1076 18880 2764 18920
rect 2804 18880 2813 18920
rect 4919 18880 4928 18920
rect 4968 18880 5010 18920
rect 5050 18880 5092 18920
rect 5132 18880 5174 18920
rect 5214 18880 5256 18920
rect 5296 18880 5305 18920
rect 6019 18880 6028 18920
rect 6068 18880 6604 18920
rect 6644 18880 6653 18920
rect 9763 18880 9772 18920
rect 9812 18880 11636 18920
rect 11779 18880 11788 18920
rect 11828 18880 12076 18920
rect 12116 18880 12125 18920
rect 14179 18880 14188 18920
rect 14228 18880 15052 18920
rect 15092 18880 15101 18920
rect 19075 18880 19084 18920
rect 19124 18880 19468 18920
rect 19508 18880 19517 18920
rect 20039 18880 20048 18920
rect 20088 18880 20130 18920
rect 20170 18880 20212 18920
rect 20252 18880 20294 18920
rect 20334 18880 20376 18920
rect 20416 18880 20425 18920
rect 20524 18880 21504 18920
rect 0 18860 80 18880
rect 6019 18879 6077 18880
rect 2179 18796 2188 18836
rect 2228 18796 2956 18836
rect 2996 18796 3005 18836
rect 5635 18796 5644 18836
rect 5684 18796 10924 18836
rect 10964 18796 11360 18836
rect 8995 18752 9053 18753
rect 11320 18752 11360 18796
rect 11491 18752 11549 18753
rect 4291 18712 4300 18752
rect 4340 18712 4588 18752
rect 4628 18712 4637 18752
rect 4867 18712 4876 18752
rect 4916 18712 5356 18752
rect 5396 18712 5405 18752
rect 6499 18712 6508 18752
rect 6548 18712 8428 18752
rect 8468 18712 8477 18752
rect 8995 18712 9004 18752
rect 9044 18712 9964 18752
rect 10004 18712 10013 18752
rect 11320 18712 11500 18752
rect 11540 18712 11549 18752
rect 11596 18752 11636 18880
rect 12067 18879 12125 18880
rect 19459 18879 19517 18880
rect 21424 18860 21504 18880
rect 14275 18796 14284 18836
rect 14324 18796 14476 18836
rect 14516 18796 14525 18836
rect 14572 18796 17260 18836
rect 17300 18796 17309 18836
rect 14572 18752 14612 18796
rect 16291 18752 16349 18753
rect 16675 18752 16733 18753
rect 11596 18712 14612 18752
rect 14659 18712 14668 18752
rect 14708 18712 14860 18752
rect 14900 18712 14909 18752
rect 16206 18712 16300 18752
rect 16340 18712 16349 18752
rect 16483 18712 16492 18752
rect 16532 18712 16684 18752
rect 16724 18712 16733 18752
rect 8995 18711 9053 18712
rect 11491 18711 11549 18712
rect 16291 18711 16349 18712
rect 16675 18711 16733 18712
rect 16867 18752 16925 18753
rect 16867 18712 16876 18752
rect 16916 18712 18700 18752
rect 18740 18712 18749 18752
rect 18883 18712 18892 18752
rect 18932 18712 19756 18752
rect 19796 18712 19805 18752
rect 16867 18711 16925 18712
rect 3427 18668 3485 18669
rect 18403 18668 18461 18669
rect 2275 18628 2284 18668
rect 2324 18628 3052 18668
rect 3092 18628 3101 18668
rect 3342 18628 3436 18668
rect 3476 18628 3485 18668
rect 3427 18627 3485 18628
rect 4012 18628 8812 18668
rect 8852 18628 8861 18668
rect 15523 18628 15532 18668
rect 15572 18628 15916 18668
rect 15956 18628 18412 18668
rect 18452 18628 18461 18668
rect 0 18584 80 18604
rect 4012 18584 4052 18628
rect 18403 18627 18461 18628
rect 4771 18584 4829 18585
rect 16867 18584 16925 18585
rect 0 18544 4052 18584
rect 4099 18544 4108 18584
rect 4148 18544 4780 18584
rect 4820 18544 4829 18584
rect 5059 18544 5068 18584
rect 5108 18544 7756 18584
rect 7796 18544 9676 18584
rect 9716 18544 11980 18584
rect 12020 18544 12029 18584
rect 12835 18544 12844 18584
rect 12884 18544 13324 18584
rect 13364 18544 13373 18584
rect 13891 18544 13900 18584
rect 13940 18544 14092 18584
rect 14132 18544 14141 18584
rect 14188 18544 16876 18584
rect 16916 18544 16925 18584
rect 17155 18544 17164 18584
rect 17204 18544 18124 18584
rect 18164 18544 18173 18584
rect 0 18524 80 18544
rect 4771 18543 4829 18544
rect 11491 18500 11549 18501
rect 12355 18500 12413 18501
rect 14188 18500 14228 18544
rect 16867 18543 16925 18544
rect 14563 18500 14621 18501
rect 2947 18460 2956 18500
rect 2996 18460 7660 18500
rect 7700 18460 7709 18500
rect 11491 18460 11500 18500
rect 11540 18460 12364 18500
rect 12404 18460 12413 18500
rect 12643 18460 12652 18500
rect 12692 18460 12940 18500
rect 12980 18460 12989 18500
rect 14179 18460 14188 18500
rect 14228 18460 14237 18500
rect 14371 18460 14380 18500
rect 14420 18460 14572 18500
rect 14612 18460 14621 18500
rect 16099 18460 16108 18500
rect 16148 18460 16157 18500
rect 16387 18460 16396 18500
rect 16436 18460 18412 18500
rect 18452 18460 18461 18500
rect 11491 18459 11549 18460
rect 12355 18459 12413 18460
rect 4675 18416 4733 18417
rect 11683 18416 11741 18417
rect 14188 18416 14228 18460
rect 14563 18459 14621 18460
rect 2755 18376 2764 18416
rect 2804 18376 3244 18416
rect 3284 18376 3820 18416
rect 3860 18376 3869 18416
rect 4675 18376 4684 18416
rect 4724 18376 8140 18416
rect 8180 18376 8428 18416
rect 8468 18376 8477 18416
rect 11683 18376 11692 18416
rect 11732 18376 14228 18416
rect 16108 18416 16148 18460
rect 21424 18416 21504 18436
rect 16108 18376 16300 18416
rect 16340 18376 16349 18416
rect 21187 18376 21196 18416
rect 21236 18376 21504 18416
rect 4675 18375 4733 18376
rect 11683 18375 11741 18376
rect 21424 18356 21504 18376
rect 2851 18292 2860 18332
rect 2900 18292 3628 18332
rect 3668 18292 3677 18332
rect 4195 18292 4204 18332
rect 4244 18292 4588 18332
rect 4628 18292 4637 18332
rect 6787 18292 6796 18332
rect 6836 18292 10060 18332
rect 10100 18292 10540 18332
rect 10580 18292 10589 18332
rect 16099 18292 16108 18332
rect 16148 18292 17740 18332
rect 17780 18292 17789 18332
rect 0 18248 80 18268
rect 4579 18248 4637 18249
rect 14179 18248 14237 18249
rect 0 18208 1268 18248
rect 1315 18208 1324 18248
rect 1364 18208 4588 18248
rect 4628 18208 12364 18248
rect 12404 18208 12413 18248
rect 14179 18208 14188 18248
rect 14228 18208 15532 18248
rect 15572 18208 15581 18248
rect 17932 18208 19468 18248
rect 19508 18208 19517 18248
rect 0 18188 80 18208
rect 1228 18164 1268 18208
rect 4579 18207 4637 18208
rect 14179 18207 14237 18208
rect 1987 18164 2045 18165
rect 2371 18164 2429 18165
rect 8323 18164 8381 18165
rect 17932 18164 17972 18208
rect 1228 18124 1996 18164
rect 2036 18124 2380 18164
rect 2420 18124 2429 18164
rect 3679 18124 3688 18164
rect 3728 18124 3770 18164
rect 3810 18124 3852 18164
rect 3892 18124 3934 18164
rect 3974 18124 4016 18164
rect 4056 18124 4065 18164
rect 4195 18124 4204 18164
rect 4244 18124 4492 18164
rect 4532 18124 4541 18164
rect 4771 18124 4780 18164
rect 4820 18124 8332 18164
rect 8372 18124 8381 18164
rect 10723 18124 10732 18164
rect 10772 18124 17932 18164
rect 17972 18124 17981 18164
rect 18799 18124 18808 18164
rect 18848 18124 18890 18164
rect 18930 18124 18972 18164
rect 19012 18124 19054 18164
rect 19094 18124 19136 18164
rect 19176 18124 19185 18164
rect 1987 18123 2045 18124
rect 2371 18123 2429 18124
rect 8323 18123 8381 18124
rect 4579 18080 4637 18081
rect 2500 18040 4396 18080
rect 4436 18040 4445 18080
rect 4579 18040 4588 18080
rect 4628 18040 5356 18080
rect 5396 18040 5405 18080
rect 9571 18040 9580 18080
rect 9620 18040 10828 18080
rect 10868 18040 12652 18080
rect 12692 18040 12701 18080
rect 12835 18040 12844 18080
rect 12884 18040 14668 18080
rect 14708 18040 15436 18080
rect 15476 18040 15485 18080
rect 2500 17996 2540 18040
rect 4579 18039 4637 18040
rect 2371 17956 2380 17996
rect 2420 17956 2540 17996
rect 3811 17956 3820 17996
rect 3860 17956 11884 17996
rect 11924 17956 11933 17996
rect 15523 17956 15532 17996
rect 15572 17956 20236 17996
rect 20276 17956 20285 17996
rect 0 17912 80 17932
rect 12355 17912 12413 17913
rect 12739 17912 12797 17913
rect 19843 17912 19901 17913
rect 21424 17912 21504 17932
rect 0 17872 12076 17912
rect 12116 17872 12125 17912
rect 12355 17872 12364 17912
rect 12404 17872 12460 17912
rect 12500 17872 12509 17912
rect 12654 17872 12748 17912
rect 12788 17872 12797 17912
rect 12931 17872 12940 17912
rect 12980 17872 13804 17912
rect 13844 17872 15244 17912
rect 15284 17872 15293 17912
rect 19843 17872 19852 17912
rect 19892 17872 21504 17912
rect 0 17852 80 17872
rect 12355 17871 12413 17872
rect 12739 17871 12797 17872
rect 19843 17871 19901 17872
rect 21424 17852 21504 17872
rect 3331 17788 3340 17828
rect 3380 17788 3628 17828
rect 3668 17788 3677 17828
rect 4099 17788 4108 17828
rect 4148 17788 4492 17828
rect 4532 17788 4541 17828
rect 6883 17788 6892 17828
rect 6932 17788 6941 17828
rect 12163 17788 12172 17828
rect 12212 17788 13900 17828
rect 13940 17788 13949 17828
rect 16291 17788 16300 17828
rect 16340 17788 19028 17828
rect 1699 17704 1708 17744
rect 1748 17704 2668 17744
rect 2708 17704 3532 17744
rect 3572 17704 3581 17744
rect 4387 17704 4396 17744
rect 4436 17704 5068 17744
rect 5108 17704 5117 17744
rect 3235 17660 3293 17661
rect 3427 17660 3485 17661
rect 6892 17660 6932 17788
rect 8803 17744 8861 17745
rect 10147 17744 10205 17745
rect 18988 17744 19028 17788
rect 8515 17704 8524 17744
rect 8564 17704 8812 17744
rect 8852 17704 8861 17744
rect 10062 17704 10156 17744
rect 10196 17704 10205 17744
rect 12451 17704 12460 17744
rect 12500 17704 12844 17744
rect 12884 17704 12893 17744
rect 13123 17704 13132 17744
rect 13172 17704 14668 17744
rect 14708 17704 14860 17744
rect 14900 17704 14909 17744
rect 16579 17704 16588 17744
rect 16628 17704 17452 17744
rect 17492 17704 17501 17744
rect 18211 17704 18220 17744
rect 18260 17704 18269 17744
rect 18979 17704 18988 17744
rect 19028 17704 19852 17744
rect 19892 17704 19901 17744
rect 8803 17703 8861 17704
rect 10147 17703 10205 17704
rect 7459 17660 7517 17661
rect 8899 17660 8957 17661
rect 3150 17620 3244 17660
rect 3284 17620 3293 17660
rect 3342 17620 3436 17660
rect 3476 17620 3485 17660
rect 5251 17620 5260 17660
rect 5300 17620 6412 17660
rect 6452 17620 6461 17660
rect 6691 17620 6700 17660
rect 6740 17620 6932 17660
rect 7374 17620 7468 17660
rect 7508 17620 7517 17660
rect 8814 17620 8908 17660
rect 8948 17620 8957 17660
rect 3235 17619 3293 17620
rect 3427 17619 3485 17620
rect 7459 17619 7517 17620
rect 8899 17619 8957 17620
rect 11395 17660 11453 17661
rect 18220 17660 18260 17704
rect 11395 17620 11404 17660
rect 11444 17620 11538 17660
rect 11875 17620 11884 17660
rect 11924 17620 12500 17660
rect 12547 17620 12556 17660
rect 12596 17620 14092 17660
rect 14132 17620 14284 17660
rect 14324 17620 14333 17660
rect 15619 17620 15628 17660
rect 15668 17620 15916 17660
rect 15956 17620 15965 17660
rect 16963 17620 16972 17660
rect 17012 17620 17260 17660
rect 17300 17620 17309 17660
rect 17356 17620 19084 17660
rect 19124 17620 19133 17660
rect 11395 17619 11453 17620
rect 0 17576 80 17596
rect 12460 17576 12500 17620
rect 17356 17576 17396 17620
rect 0 17536 1804 17576
rect 1844 17536 2572 17576
rect 2612 17536 7756 17576
rect 7796 17536 7805 17576
rect 12460 17536 12844 17576
rect 12884 17536 12893 17576
rect 17347 17536 17356 17576
rect 17396 17536 17405 17576
rect 0 17516 80 17536
rect 16003 17492 16061 17493
rect 6595 17452 6604 17492
rect 6644 17452 6988 17492
rect 7028 17452 7037 17492
rect 11971 17452 11980 17492
rect 12020 17452 16012 17492
rect 16052 17452 16061 17492
rect 16003 17451 16061 17452
rect 21424 17408 21504 17428
rect 4919 17368 4928 17408
rect 4968 17368 5010 17408
rect 5050 17368 5092 17408
rect 5132 17368 5174 17408
rect 5214 17368 5256 17408
rect 5296 17368 5305 17408
rect 12739 17368 12748 17408
rect 12788 17368 14380 17408
rect 14420 17368 14429 17408
rect 20039 17368 20048 17408
rect 20088 17368 20130 17408
rect 20170 17368 20212 17408
rect 20252 17368 20294 17408
rect 20334 17368 20376 17408
rect 20416 17368 20425 17408
rect 20611 17368 20620 17408
rect 20660 17368 21504 17408
rect 21424 17348 21504 17368
rect 0 17240 80 17260
rect 0 17200 7276 17240
rect 7316 17200 7325 17240
rect 0 17180 80 17200
rect 6211 17116 6220 17156
rect 6260 17116 8332 17156
rect 8372 17116 8381 17156
rect 11683 17116 11692 17156
rect 11732 17116 11741 17156
rect 1315 17072 1373 17073
rect 1230 17032 1324 17072
rect 1364 17032 2380 17072
rect 2420 17032 2429 17072
rect 9187 17032 9196 17072
rect 9236 17032 9580 17072
rect 9620 17032 11116 17072
rect 11156 17032 11165 17072
rect 1315 17031 1373 17032
rect 10339 16988 10397 16989
rect 10339 16948 10348 16988
rect 10388 16948 10444 16988
rect 10484 16948 10493 16988
rect 10339 16947 10397 16948
rect 0 16904 80 16924
rect 0 16864 11020 16904
rect 11060 16864 11069 16904
rect 0 16844 80 16864
rect 11692 16820 11732 17116
rect 16099 17072 16157 17073
rect 16099 17032 16108 17072
rect 16148 17032 16396 17072
rect 16436 17032 16780 17072
rect 16820 17032 16829 17072
rect 16099 17031 16157 17032
rect 18691 16948 18700 16988
rect 18740 16948 19660 16988
rect 19700 16948 19709 16988
rect 20899 16904 20957 16905
rect 21424 16904 21504 16924
rect 15811 16864 15820 16904
rect 15860 16864 19564 16904
rect 19604 16864 19613 16904
rect 20899 16864 20908 16904
rect 20948 16864 21504 16904
rect 20899 16863 20957 16864
rect 21424 16844 21504 16864
rect 11683 16780 11692 16820
rect 11732 16780 11741 16820
rect 8323 16736 8381 16737
rect 5443 16696 5452 16736
rect 5492 16696 8332 16736
rect 8372 16696 8620 16736
rect 8660 16696 8669 16736
rect 8323 16695 8381 16696
rect 2947 16612 2956 16652
rect 2996 16612 3340 16652
rect 3380 16612 3389 16652
rect 3679 16612 3688 16652
rect 3728 16612 3770 16652
rect 3810 16612 3852 16652
rect 3892 16612 3934 16652
rect 3974 16612 4016 16652
rect 4056 16612 4065 16652
rect 7459 16612 7468 16652
rect 7508 16612 9908 16652
rect 9955 16612 9964 16652
rect 10004 16612 12172 16652
rect 12212 16612 12221 16652
rect 18799 16612 18808 16652
rect 18848 16612 18890 16652
rect 18930 16612 18972 16652
rect 19012 16612 19054 16652
rect 19094 16612 19136 16652
rect 19176 16612 19185 16652
rect 0 16568 80 16588
rect 9868 16568 9908 16612
rect 12547 16568 12605 16569
rect 0 16528 9772 16568
rect 9812 16528 9821 16568
rect 9868 16528 12556 16568
rect 12596 16528 12605 16568
rect 0 16508 80 16528
rect 12547 16527 12605 16528
rect 6019 16484 6077 16485
rect 3139 16444 3148 16484
rect 3188 16444 3724 16484
rect 3764 16444 3773 16484
rect 5934 16444 6028 16484
rect 6068 16444 6077 16484
rect 6691 16444 6700 16484
rect 6740 16444 8620 16484
rect 8660 16444 9196 16484
rect 9236 16444 9245 16484
rect 12067 16444 12076 16484
rect 12116 16444 12460 16484
rect 12500 16444 12509 16484
rect 15331 16444 15340 16484
rect 15380 16444 19276 16484
rect 19316 16444 19325 16484
rect 6019 16443 6077 16444
rect 11971 16400 12029 16401
rect 17347 16400 17405 16401
rect 18595 16400 18653 16401
rect 1420 16360 2540 16400
rect 2947 16360 2956 16400
rect 2996 16360 3244 16400
rect 3284 16360 3293 16400
rect 4012 16360 4972 16400
rect 5012 16360 5021 16400
rect 5347 16360 5356 16400
rect 5396 16360 6220 16400
rect 6260 16360 6269 16400
rect 7363 16360 7372 16400
rect 7412 16360 11980 16400
rect 12020 16360 12029 16400
rect 13123 16360 13132 16400
rect 13172 16360 13324 16400
rect 13364 16360 15148 16400
rect 15188 16360 15197 16400
rect 17262 16360 17356 16400
rect 17396 16360 17405 16400
rect 18211 16360 18220 16400
rect 18260 16360 18508 16400
rect 18548 16360 18604 16400
rect 18644 16360 18653 16400
rect 0 16232 80 16252
rect 1420 16232 1460 16360
rect 2500 16316 2540 16360
rect 4012 16316 4052 16360
rect 11971 16359 12029 16360
rect 17347 16359 17405 16360
rect 18595 16359 18653 16360
rect 19555 16400 19613 16401
rect 20707 16400 20765 16401
rect 21424 16400 21504 16420
rect 19555 16360 19564 16400
rect 19604 16360 20044 16400
rect 20084 16360 20093 16400
rect 20707 16360 20716 16400
rect 20756 16360 21504 16400
rect 19555 16359 19613 16360
rect 20707 16359 20765 16360
rect 21424 16340 21504 16360
rect 14179 16316 14237 16317
rect 2500 16276 4052 16316
rect 4108 16276 9004 16316
rect 9044 16276 11360 16316
rect 13603 16276 13612 16316
rect 13652 16276 13661 16316
rect 14094 16276 14188 16316
rect 14228 16276 14380 16316
rect 14420 16276 14429 16316
rect 4108 16232 4148 16276
rect 4291 16232 4349 16233
rect 0 16192 1460 16232
rect 1507 16192 1516 16232
rect 1556 16192 4148 16232
rect 4206 16192 4300 16232
rect 4340 16192 4349 16232
rect 0 16172 80 16192
rect 4291 16191 4349 16192
rect 7939 16232 7997 16233
rect 7939 16192 7948 16232
rect 7988 16192 10156 16232
rect 10196 16192 10205 16232
rect 7939 16191 7997 16192
rect 7267 16148 7325 16149
rect 11320 16148 11360 16276
rect 11875 16192 11884 16232
rect 11924 16192 12460 16232
rect 12500 16192 12509 16232
rect 13315 16201 13324 16241
rect 13364 16232 13373 16241
rect 13612 16232 13652 16276
rect 14179 16275 14237 16276
rect 13364 16201 13652 16232
rect 13324 16192 13652 16201
rect 13795 16192 13804 16232
rect 13844 16192 14092 16232
rect 14132 16192 14141 16232
rect 16579 16192 16588 16232
rect 16628 16192 16780 16232
rect 16820 16192 17356 16232
rect 17396 16192 17405 16232
rect 18115 16192 18124 16232
rect 18164 16192 18604 16232
rect 18644 16192 18796 16232
rect 18836 16192 18845 16232
rect 12067 16148 12125 16149
rect 7267 16108 7276 16148
rect 7316 16108 9676 16148
rect 9716 16108 10252 16148
rect 10292 16108 10301 16148
rect 11320 16108 12076 16148
rect 12116 16108 12125 16148
rect 7267 16107 7325 16108
rect 12067 16107 12125 16108
rect 12451 16064 12509 16065
rect 5827 16024 5836 16064
rect 5876 16024 6220 16064
rect 6260 16024 6269 16064
rect 9283 16024 9292 16064
rect 9332 16024 9772 16064
rect 9812 16024 9821 16064
rect 12451 16024 12460 16064
rect 12500 16024 12652 16064
rect 12692 16024 12701 16064
rect 14083 16024 14092 16064
rect 14132 16024 14668 16064
rect 14708 16024 14717 16064
rect 12451 16023 12509 16024
rect 5827 15980 5885 15981
rect 17539 15980 17597 15981
rect 2659 15940 2668 15980
rect 2708 15940 3148 15980
rect 3188 15940 3197 15980
rect 3811 15940 3820 15980
rect 3860 15940 5836 15980
rect 5876 15940 11360 15980
rect 13315 15940 13324 15980
rect 13364 15940 13708 15980
rect 13748 15940 13757 15980
rect 17347 15940 17356 15980
rect 17396 15940 17548 15980
rect 17588 15940 19756 15980
rect 19796 15940 19805 15980
rect 5827 15939 5885 15940
rect 0 15896 80 15916
rect 0 15856 1900 15896
rect 1940 15856 1949 15896
rect 4919 15856 4928 15896
rect 4968 15856 5010 15896
rect 5050 15856 5092 15896
rect 5132 15856 5174 15896
rect 5214 15856 5256 15896
rect 5296 15856 5305 15896
rect 5443 15856 5452 15896
rect 5492 15856 5740 15896
rect 5780 15856 5789 15896
rect 6019 15856 6028 15896
rect 6068 15856 6077 15896
rect 10531 15856 10540 15896
rect 10580 15856 11116 15896
rect 11156 15856 11165 15896
rect 0 15836 80 15856
rect 6028 15812 6068 15856
rect 11320 15812 11360 15940
rect 17539 15939 17597 15940
rect 21424 15896 21504 15916
rect 20039 15856 20048 15896
rect 20088 15856 20130 15896
rect 20170 15856 20212 15896
rect 20252 15856 20294 15896
rect 20334 15856 20376 15896
rect 20416 15856 20425 15896
rect 21091 15856 21100 15896
rect 21140 15856 21504 15896
rect 21424 15836 21504 15856
rect 17347 15812 17405 15813
rect 2083 15772 2092 15812
rect 2132 15772 6068 15812
rect 8899 15772 8908 15812
rect 8948 15772 9388 15812
rect 9428 15772 9437 15812
rect 10627 15772 10636 15812
rect 10676 15772 10828 15812
rect 10868 15772 10877 15812
rect 11320 15772 12268 15812
rect 12308 15772 12317 15812
rect 17262 15772 17356 15812
rect 17396 15772 17405 15812
rect 17347 15771 17405 15772
rect 5251 15688 5260 15728
rect 5300 15688 5932 15728
rect 5972 15688 5981 15728
rect 6028 15688 12076 15728
rect 12116 15688 12125 15728
rect 17827 15688 17836 15728
rect 17876 15688 18124 15728
rect 18164 15688 18173 15728
rect 6028 15644 6068 15688
rect 1603 15604 1612 15644
rect 1652 15604 2540 15644
rect 2851 15604 2860 15644
rect 2900 15604 3340 15644
rect 3380 15604 3389 15644
rect 5059 15604 5068 15644
rect 5108 15604 5548 15644
rect 5588 15604 6068 15644
rect 6883 15604 6892 15644
rect 6932 15604 7180 15644
rect 7220 15604 7229 15644
rect 11011 15604 11020 15644
rect 11060 15604 11596 15644
rect 11636 15604 11788 15644
rect 11828 15604 13132 15644
rect 13172 15604 13181 15644
rect 0 15560 80 15580
rect 2500 15560 2540 15604
rect 5731 15560 5789 15561
rect 0 15520 1516 15560
rect 1556 15520 1565 15560
rect 2500 15520 5396 15560
rect 5443 15520 5452 15560
rect 5492 15520 5740 15560
rect 5780 15520 5789 15560
rect 0 15500 80 15520
rect 5356 15476 5396 15520
rect 5731 15519 5789 15520
rect 6019 15560 6077 15561
rect 7267 15560 7325 15561
rect 7939 15560 7997 15561
rect 6019 15520 6028 15560
rect 6068 15520 6700 15560
rect 6740 15520 6749 15560
rect 7182 15520 7276 15560
rect 7316 15520 7325 15560
rect 7747 15520 7756 15560
rect 7796 15520 7948 15560
rect 7988 15520 7997 15560
rect 6019 15519 6077 15520
rect 7267 15519 7325 15520
rect 7939 15519 7997 15520
rect 8044 15520 8812 15560
rect 8852 15520 13900 15560
rect 13940 15520 13949 15560
rect 16291 15520 16300 15560
rect 16340 15520 16972 15560
rect 17012 15520 17021 15560
rect 17155 15520 17164 15560
rect 17204 15520 17836 15560
rect 17876 15520 17885 15560
rect 2371 15436 2380 15476
rect 2420 15436 2540 15476
rect 5356 15436 7372 15476
rect 7412 15436 7421 15476
rect 2500 15392 2540 15436
rect 8044 15392 8084 15520
rect 19555 15476 19613 15477
rect 10339 15436 10348 15476
rect 10388 15436 10635 15476
rect 10675 15436 10684 15476
rect 16867 15436 16876 15476
rect 16916 15436 17260 15476
rect 17300 15436 19564 15476
rect 19604 15436 19613 15476
rect 19555 15435 19613 15436
rect 21424 15392 21504 15412
rect 2500 15352 8084 15392
rect 10147 15352 10156 15392
rect 10196 15352 10732 15392
rect 10772 15352 10781 15392
rect 16195 15352 16204 15392
rect 16244 15352 21504 15392
rect 21424 15332 21504 15352
rect 7075 15308 7133 15309
rect 6691 15268 6700 15308
rect 6740 15268 7084 15308
rect 7124 15268 7756 15308
rect 7796 15268 9388 15308
rect 9428 15268 9964 15308
rect 10004 15268 11020 15308
rect 11060 15268 11069 15308
rect 7075 15267 7133 15268
rect 0 15224 80 15244
rect 0 15184 17932 15224
rect 17972 15184 17981 15224
rect 0 15164 80 15184
rect 3679 15100 3688 15140
rect 3728 15100 3770 15140
rect 3810 15100 3852 15140
rect 3892 15100 3934 15140
rect 3974 15100 4016 15140
rect 4056 15100 4065 15140
rect 6883 15100 6892 15140
rect 6932 15100 7660 15140
rect 7700 15100 10060 15140
rect 10100 15100 10636 15140
rect 10676 15100 10685 15140
rect 12835 15100 12844 15140
rect 12884 15100 14284 15140
rect 14324 15100 14333 15140
rect 16387 15100 16396 15140
rect 16436 15100 18316 15140
rect 18356 15100 18365 15140
rect 18799 15100 18808 15140
rect 18848 15100 18890 15140
rect 18930 15100 18972 15140
rect 19012 15100 19054 15140
rect 19094 15100 19136 15140
rect 19176 15100 19185 15140
rect 15811 15016 15820 15056
rect 15860 15016 16300 15056
rect 16340 15016 16349 15056
rect 12739 14972 12797 14973
rect 7939 14932 7948 14972
rect 7988 14932 8716 14972
rect 8756 14932 8765 14972
rect 12739 14932 12748 14972
rect 12788 14932 12844 14972
rect 12884 14932 12893 14972
rect 14659 14932 14668 14972
rect 14708 14932 18124 14972
rect 18164 14932 18173 14972
rect 12739 14931 12797 14932
rect 0 14888 80 14908
rect 21424 14888 21504 14908
rect 0 14848 2284 14888
rect 2324 14848 2333 14888
rect 4099 14848 4108 14888
rect 4148 14848 21504 14888
rect 0 14828 80 14848
rect 21424 14828 21504 14848
rect 8419 14804 8477 14805
rect 2083 14764 2092 14804
rect 2132 14764 4396 14804
rect 4436 14764 4445 14804
rect 6499 14764 6508 14804
rect 6548 14764 8428 14804
rect 8468 14764 8477 14804
rect 14179 14764 14188 14804
rect 14228 14764 16684 14804
rect 16724 14764 18892 14804
rect 18932 14764 18941 14804
rect 8419 14763 8477 14764
rect 3235 14720 3293 14721
rect 16099 14720 16157 14721
rect 19363 14720 19421 14721
rect 3150 14680 3244 14720
rect 3284 14680 3293 14720
rect 5059 14680 5068 14720
rect 5108 14680 5452 14720
rect 5492 14680 5501 14720
rect 5923 14680 5932 14720
rect 5972 14680 6412 14720
rect 6452 14680 6461 14720
rect 7267 14680 7276 14720
rect 7316 14680 8236 14720
rect 8276 14680 10828 14720
rect 10868 14680 11212 14720
rect 11252 14680 11261 14720
rect 16014 14680 16108 14720
rect 16148 14680 16157 14720
rect 19278 14680 19372 14720
rect 19412 14680 19421 14720
rect 3235 14679 3293 14680
rect 16099 14679 16157 14680
rect 19363 14679 19421 14680
rect 11971 14636 12029 14637
rect 3715 14596 3724 14636
rect 3764 14596 8332 14636
rect 8372 14596 9100 14636
rect 9140 14596 9149 14636
rect 11971 14596 11980 14636
rect 12020 14596 17356 14636
rect 17396 14596 19084 14636
rect 19124 14596 19133 14636
rect 11971 14595 12029 14596
rect 0 14552 80 14572
rect 0 14512 1516 14552
rect 1556 14512 1565 14552
rect 2500 14512 15340 14552
rect 15380 14512 15389 14552
rect 16483 14512 16492 14552
rect 16532 14512 17452 14552
rect 17492 14512 17501 14552
rect 0 14492 80 14512
rect 2500 14468 2540 14512
rect 5827 14468 5885 14469
rect 9571 14468 9629 14469
rect 1987 14428 1996 14468
rect 2036 14428 2540 14468
rect 5742 14428 5836 14468
rect 5876 14428 5885 14468
rect 8131 14428 8140 14468
rect 8180 14428 9580 14468
rect 9620 14428 9629 14468
rect 5827 14427 5885 14428
rect 9571 14427 9629 14428
rect 6499 14384 6557 14385
rect 8419 14384 8477 14385
rect 10915 14384 10973 14385
rect 21424 14384 21504 14404
rect 4919 14344 4928 14384
rect 4968 14344 5010 14384
rect 5050 14344 5092 14384
rect 5132 14344 5174 14384
rect 5214 14344 5256 14384
rect 5296 14344 5305 14384
rect 6499 14344 6508 14384
rect 6548 14344 6604 14384
rect 6644 14344 6653 14384
rect 8419 14344 8428 14384
rect 8468 14344 10924 14384
rect 10964 14344 10973 14384
rect 20039 14344 20048 14384
rect 20088 14344 20130 14384
rect 20170 14344 20212 14384
rect 20252 14344 20294 14384
rect 20334 14344 20376 14384
rect 20416 14344 20425 14384
rect 20524 14344 21504 14384
rect 6499 14343 6557 14344
rect 8419 14343 8477 14344
rect 10915 14343 10973 14344
rect 4387 14300 4445 14301
rect 20524 14300 20564 14344
rect 21424 14324 21504 14344
rect 4387 14260 4396 14300
rect 4436 14260 20564 14300
rect 4387 14259 4445 14260
rect 0 14216 80 14236
rect 12355 14216 12413 14217
rect 0 14176 1324 14216
rect 1364 14176 1373 14216
rect 11875 14176 11884 14216
rect 11924 14176 12364 14216
rect 12404 14176 12413 14216
rect 17635 14176 17644 14216
rect 17684 14176 18316 14216
rect 18356 14176 18365 14216
rect 0 14156 80 14176
rect 12355 14175 12413 14176
rect 3043 14132 3101 14133
rect 2659 14092 2668 14132
rect 2708 14092 3052 14132
rect 3092 14092 3101 14132
rect 4291 14092 4300 14132
rect 4340 14092 7372 14132
rect 7412 14092 7421 14132
rect 3043 14091 3101 14092
rect 8323 14048 8381 14049
rect 10147 14048 10205 14049
rect 1699 14008 1708 14048
rect 1748 14008 5548 14048
rect 5588 14008 5597 14048
rect 5923 14008 5932 14048
rect 5972 14008 6892 14048
rect 6932 14008 6941 14048
rect 7843 14008 7852 14048
rect 7892 14008 8332 14048
rect 8372 14008 8381 14048
rect 10062 14008 10156 14048
rect 10196 14008 10205 14048
rect 11683 14008 11692 14048
rect 11732 14008 12364 14048
rect 12404 14008 12413 14048
rect 13027 14008 13036 14048
rect 13076 14008 13804 14048
rect 13844 14008 13853 14048
rect 17251 14008 17260 14048
rect 17300 14008 19276 14048
rect 19316 14008 19325 14048
rect 8323 14007 8381 14008
rect 10147 14007 10205 14008
rect 13315 13964 13373 13965
rect 17539 13964 17597 13965
rect 2083 13924 2092 13964
rect 2132 13924 2141 13964
rect 2563 13924 2572 13964
rect 2612 13924 3340 13964
rect 3380 13924 3916 13964
rect 3956 13924 5260 13964
rect 5300 13924 6412 13964
rect 6452 13924 8236 13964
rect 8276 13924 8285 13964
rect 13315 13924 13324 13964
rect 13364 13924 13420 13964
rect 13460 13924 15052 13964
rect 15092 13924 17548 13964
rect 17588 13924 17836 13964
rect 17876 13924 17885 13964
rect 0 13880 80 13900
rect 2092 13880 2132 13924
rect 13315 13923 13373 13924
rect 17539 13923 17597 13924
rect 20707 13880 20765 13881
rect 21424 13880 21504 13900
rect 0 13840 1900 13880
rect 1940 13840 1949 13880
rect 2092 13840 15628 13880
rect 15668 13840 15677 13880
rect 18700 13840 19084 13880
rect 19124 13840 19133 13880
rect 20707 13840 20716 13880
rect 20756 13840 21504 13880
rect 0 13820 80 13840
rect 6691 13796 6749 13797
rect 5059 13756 5068 13796
rect 5108 13756 5644 13796
rect 5684 13756 5693 13796
rect 6691 13756 6700 13796
rect 6740 13756 7756 13796
rect 7796 13756 7805 13796
rect 8035 13756 8044 13796
rect 8084 13756 11692 13796
rect 11732 13756 11741 13796
rect 6691 13755 6749 13756
rect 7651 13672 7660 13712
rect 7700 13672 11788 13712
rect 11828 13672 11837 13712
rect 10147 13628 10205 13629
rect 3679 13588 3688 13628
rect 3728 13588 3770 13628
rect 3810 13588 3852 13628
rect 3892 13588 3934 13628
rect 3974 13588 4016 13628
rect 4056 13588 4065 13628
rect 10051 13588 10060 13628
rect 10100 13588 10156 13628
rect 10196 13588 10205 13628
rect 10147 13587 10205 13588
rect 0 13544 80 13564
rect 0 13504 1804 13544
rect 1844 13504 1853 13544
rect 8707 13504 8716 13544
rect 8756 13504 12844 13544
rect 12884 13504 12893 13544
rect 0 13484 80 13504
rect 14083 13420 14092 13460
rect 14132 13420 15532 13460
rect 15572 13420 15581 13460
rect 16387 13420 16396 13460
rect 16436 13420 17356 13460
rect 17396 13420 17405 13460
rect 17635 13420 17644 13460
rect 17684 13420 18028 13460
rect 18068 13420 18077 13460
rect 2500 13336 17396 13376
rect 2500 13292 2540 13336
rect 17356 13292 17396 13336
rect 18700 13292 18740 13840
rect 20707 13839 20765 13840
rect 21424 13820 21504 13840
rect 18799 13588 18808 13628
rect 18848 13588 18890 13628
rect 18930 13588 18972 13628
rect 19012 13588 19054 13628
rect 19094 13588 19136 13628
rect 19176 13588 19185 13628
rect 18892 13504 19372 13544
rect 19412 13504 19421 13544
rect 18892 13460 18932 13504
rect 18883 13420 18892 13460
rect 18932 13420 18941 13460
rect 21424 13376 21504 13396
rect 20707 13336 20716 13376
rect 20756 13336 21504 13376
rect 21424 13316 21504 13336
rect 1507 13252 1516 13292
rect 1556 13252 2540 13292
rect 3523 13252 3532 13292
rect 3572 13252 8716 13292
rect 8756 13252 8765 13292
rect 12931 13252 12940 13292
rect 12980 13252 13556 13292
rect 14947 13252 14956 13292
rect 14996 13252 16724 13292
rect 17347 13252 17356 13292
rect 17396 13252 17405 13292
rect 18211 13252 18220 13292
rect 18260 13252 18269 13292
rect 18691 13252 18700 13292
rect 18740 13252 18749 13292
rect 0 13208 80 13228
rect 6115 13208 6173 13209
rect 13516 13208 13556 13252
rect 16684 13208 16724 13252
rect 18220 13208 18260 13252
rect 0 13168 1940 13208
rect 3139 13168 3148 13208
rect 3188 13168 4396 13208
rect 4436 13168 6124 13208
rect 6164 13168 6173 13208
rect 10915 13168 10924 13208
rect 10964 13168 13420 13208
rect 13460 13168 13469 13208
rect 13516 13168 13612 13208
rect 13652 13168 15244 13208
rect 15284 13168 15293 13208
rect 16675 13168 16684 13208
rect 16724 13168 18260 13208
rect 0 13148 80 13168
rect 1900 13124 1940 13168
rect 6115 13167 6173 13168
rect 4195 13124 4253 13125
rect 1891 13084 1900 13124
rect 1940 13084 1949 13124
rect 2083 13084 2092 13124
rect 2132 13084 4204 13124
rect 4244 13084 4253 13124
rect 4195 13083 4253 13084
rect 2500 13000 20140 13040
rect 20180 13000 20189 13040
rect 2500 12956 2540 13000
rect 6499 12956 6557 12957
rect 1987 12916 1996 12956
rect 2036 12916 2540 12956
rect 6403 12916 6412 12956
rect 6452 12916 6508 12956
rect 6548 12916 6557 12956
rect 6499 12915 6557 12916
rect 0 12872 80 12892
rect 21424 12872 21504 12892
rect 0 12832 1516 12872
rect 1556 12832 1565 12872
rect 4919 12832 4928 12872
rect 4968 12832 5010 12872
rect 5050 12832 5092 12872
rect 5132 12832 5174 12872
rect 5214 12832 5256 12872
rect 5296 12832 5305 12872
rect 20039 12832 20048 12872
rect 20088 12832 20130 12872
rect 20170 12832 20212 12872
rect 20252 12832 20294 12872
rect 20334 12832 20376 12872
rect 20416 12832 20425 12872
rect 20524 12832 21504 12872
rect 0 12812 80 12832
rect 11971 12788 12029 12789
rect 20524 12788 20564 12832
rect 21424 12812 21504 12832
rect 11971 12748 11980 12788
rect 12020 12748 20564 12788
rect 11971 12747 12029 12748
rect 2467 12664 2476 12704
rect 2516 12664 10924 12704
rect 10964 12664 10973 12704
rect 15427 12664 15436 12704
rect 15476 12664 15820 12704
rect 15860 12664 15869 12704
rect 3139 12620 3197 12621
rect 1699 12580 1708 12620
rect 1748 12580 1757 12620
rect 2947 12580 2956 12620
rect 2996 12580 3148 12620
rect 3188 12580 4108 12620
rect 4148 12580 4157 12620
rect 8899 12580 8908 12620
rect 8948 12580 9196 12620
rect 9236 12580 9245 12620
rect 9763 12580 9772 12620
rect 9812 12580 11360 12620
rect 11779 12580 11788 12620
rect 11828 12580 16780 12620
rect 16820 12580 16829 12620
rect 0 12536 80 12556
rect 1708 12536 1748 12580
rect 3139 12579 3197 12580
rect 3043 12536 3101 12537
rect 8707 12536 8765 12537
rect 11320 12536 11360 12580
rect 14371 12536 14429 12537
rect 0 12496 1748 12536
rect 2467 12496 2476 12536
rect 2516 12496 3052 12536
rect 3092 12496 3101 12536
rect 3907 12496 3916 12536
rect 3956 12496 4492 12536
rect 4532 12496 4541 12536
rect 8227 12496 8236 12536
rect 8276 12496 8716 12536
rect 8756 12496 8765 12536
rect 0 12476 80 12496
rect 3043 12495 3101 12496
rect 8707 12495 8765 12496
rect 8908 12496 9868 12536
rect 9908 12496 10252 12536
rect 10292 12496 10301 12536
rect 11320 12496 13228 12536
rect 13268 12496 13516 12536
rect 13556 12496 13565 12536
rect 14371 12496 14380 12536
rect 14420 12496 14476 12536
rect 14516 12496 14525 12536
rect 16387 12496 16396 12536
rect 16436 12496 17164 12536
rect 17204 12496 17213 12536
rect 19747 12496 19756 12536
rect 19796 12496 19948 12536
rect 19988 12496 19997 12536
rect 8908 12452 8948 12496
rect 14371 12495 14429 12496
rect 2083 12412 2092 12452
rect 2132 12412 8524 12452
rect 8564 12412 8573 12452
rect 8899 12412 8908 12452
rect 8948 12412 8957 12452
rect 9763 12412 9772 12452
rect 9812 12412 11404 12452
rect 11444 12412 11692 12452
rect 11732 12412 11741 12452
rect 12931 12412 12940 12452
rect 12980 12412 15052 12452
rect 15092 12412 15101 12452
rect 20995 12368 21053 12369
rect 21424 12368 21504 12388
rect 1603 12328 1612 12368
rect 1652 12328 17068 12368
rect 17108 12328 17117 12368
rect 20995 12328 21004 12368
rect 21044 12328 21504 12368
rect 20995 12327 21053 12328
rect 21424 12308 21504 12328
rect 1699 12244 1708 12284
rect 1748 12244 14764 12284
rect 14804 12244 14813 12284
rect 18700 12244 18892 12284
rect 18932 12244 18941 12284
rect 0 12200 80 12220
rect 7459 12200 7517 12201
rect 0 12160 1516 12200
rect 1556 12160 1565 12200
rect 7459 12160 7468 12200
rect 7508 12160 7564 12200
rect 7604 12160 7613 12200
rect 7939 12160 7948 12200
rect 7988 12160 8716 12200
rect 8756 12160 8765 12200
rect 13123 12160 13132 12200
rect 13172 12160 13708 12200
rect 13748 12160 13757 12200
rect 0 12140 80 12160
rect 7459 12159 7517 12160
rect 13315 12116 13373 12117
rect 14371 12116 14429 12117
rect 3679 12076 3688 12116
rect 3728 12076 3770 12116
rect 3810 12076 3852 12116
rect 3892 12076 3934 12116
rect 3974 12076 4016 12116
rect 4056 12076 4065 12116
rect 12835 12076 12844 12116
rect 12884 12076 13324 12116
rect 13364 12076 14380 12116
rect 14420 12076 14429 12116
rect 13315 12075 13373 12076
rect 14371 12075 14429 12076
rect 16867 11992 16876 12032
rect 16916 11992 17260 12032
rect 17300 11992 17309 12032
rect 18700 11948 18740 12244
rect 18799 12076 18808 12116
rect 18848 12076 18890 12116
rect 18930 12076 18972 12116
rect 19012 12076 19054 12116
rect 19094 12076 19136 12116
rect 19176 12076 19185 12116
rect 16579 11908 16588 11948
rect 16628 11908 18988 11948
rect 19028 11908 19037 11948
rect 0 11865 80 11884
rect 0 11864 125 11865
rect 10147 11864 10205 11865
rect 10339 11864 10397 11865
rect 21424 11864 21504 11884
rect 0 11824 76 11864
rect 116 11824 125 11864
rect 5059 11824 5068 11864
rect 5108 11824 10156 11864
rect 10196 11824 10348 11864
rect 10388 11824 10397 11864
rect 18883 11824 18892 11864
rect 18932 11824 19276 11864
rect 19316 11824 21504 11864
rect 0 11823 125 11824
rect 10147 11823 10205 11824
rect 10339 11823 10397 11824
rect 0 11804 80 11823
rect 21424 11804 21504 11824
rect 1699 11740 1708 11780
rect 1748 11740 8524 11780
rect 8564 11740 8573 11780
rect 9763 11740 9772 11780
rect 9812 11740 9964 11780
rect 10004 11740 12076 11780
rect 12116 11740 12125 11780
rect 15043 11740 15052 11780
rect 15092 11740 15820 11780
rect 15860 11740 16972 11780
rect 17012 11740 17021 11780
rect 19267 11696 19325 11697
rect 3523 11656 3532 11696
rect 3572 11656 6316 11696
rect 6356 11656 6365 11696
rect 7843 11656 7852 11696
rect 7892 11656 11252 11696
rect 11587 11656 11596 11696
rect 11636 11656 12844 11696
rect 12884 11656 12893 11696
rect 13891 11656 13900 11696
rect 13940 11656 14284 11696
rect 14324 11656 14333 11696
rect 15139 11656 15148 11696
rect 15188 11656 16204 11696
rect 16244 11656 17068 11696
rect 17108 11656 17396 11696
rect 6316 11612 6356 11656
rect 9955 11612 10013 11613
rect 11212 11612 11252 11656
rect 12844 11612 12884 11656
rect 17356 11612 17396 11656
rect 19267 11656 19276 11696
rect 19316 11656 19468 11696
rect 19508 11656 19517 11696
rect 19267 11655 19325 11656
rect 2500 11572 3916 11612
rect 3956 11572 3965 11612
rect 6316 11572 8428 11612
rect 8468 11572 8477 11612
rect 9955 11572 9964 11612
rect 10004 11572 10924 11612
rect 10964 11572 10973 11612
rect 11212 11572 11884 11612
rect 11924 11572 11933 11612
rect 12844 11572 17300 11612
rect 17347 11572 17356 11612
rect 17396 11572 17405 11612
rect 0 11528 80 11548
rect 0 11488 1804 11528
rect 1844 11488 1853 11528
rect 0 11468 80 11488
rect 2500 11360 2540 11572
rect 9955 11571 10013 11572
rect 17260 11528 17300 11572
rect 4387 11488 4396 11528
rect 4436 11488 4445 11528
rect 7363 11488 7372 11528
rect 7412 11488 8236 11528
rect 8276 11488 8285 11528
rect 8995 11488 9004 11528
rect 9044 11488 9868 11528
rect 9908 11488 9917 11528
rect 15715 11488 15724 11528
rect 15764 11488 16204 11528
rect 16244 11488 16253 11528
rect 17260 11488 17932 11528
rect 17972 11488 18316 11528
rect 18356 11488 19756 11528
rect 19796 11488 19805 11528
rect 4396 11444 4436 11488
rect 3139 11404 3148 11444
rect 3188 11404 4436 11444
rect 9475 11444 9533 11445
rect 9475 11404 9484 11444
rect 9524 11404 14092 11444
rect 14132 11404 14141 11444
rect 18691 11404 18700 11444
rect 18740 11404 20564 11444
rect 9475 11403 9533 11404
rect 8803 11360 8861 11361
rect 20524 11360 20564 11404
rect 21424 11360 21504 11380
rect 1507 11320 1516 11360
rect 1556 11320 2476 11360
rect 2516 11320 2540 11360
rect 4919 11320 4928 11360
rect 4968 11320 5010 11360
rect 5050 11320 5092 11360
rect 5132 11320 5174 11360
rect 5214 11320 5256 11360
rect 5296 11320 5305 11360
rect 6691 11320 6700 11360
rect 6740 11320 7276 11360
rect 7316 11320 7468 11360
rect 7508 11320 7517 11360
rect 8803 11320 8812 11360
rect 8852 11320 8908 11360
rect 8948 11320 8957 11360
rect 20039 11320 20048 11360
rect 20088 11320 20130 11360
rect 20170 11320 20212 11360
rect 20252 11320 20294 11360
rect 20334 11320 20376 11360
rect 20416 11320 20425 11360
rect 20524 11320 21504 11360
rect 8803 11319 8861 11320
rect 21424 11300 21504 11320
rect 1699 11236 1708 11276
rect 1748 11236 16012 11276
rect 16052 11236 16061 11276
rect 0 11192 80 11212
rect 6115 11192 6173 11193
rect 9571 11192 9629 11193
rect 0 11152 2188 11192
rect 2228 11152 2237 11192
rect 6115 11152 6124 11192
rect 6164 11152 7372 11192
rect 7412 11152 7421 11192
rect 8323 11152 8332 11192
rect 8372 11152 9004 11192
rect 9044 11152 9053 11192
rect 9486 11152 9580 11192
rect 9620 11152 9629 11192
rect 14275 11152 14284 11192
rect 14324 11152 14668 11192
rect 14708 11152 14717 11192
rect 14851 11152 14860 11192
rect 14900 11152 15436 11192
rect 15476 11152 18220 11192
rect 18260 11152 18269 11192
rect 19555 11152 19564 11192
rect 19604 11152 19852 11192
rect 19892 11152 19901 11192
rect 0 11132 80 11152
rect 6115 11151 6173 11152
rect 9571 11151 9629 11152
rect 7459 11108 7517 11109
rect 5347 11068 5356 11108
rect 5396 11068 5644 11108
rect 5684 11068 5693 11108
rect 5827 11068 5836 11108
rect 5876 11068 6124 11108
rect 6164 11068 6173 11108
rect 7459 11068 7468 11108
rect 7508 11068 10060 11108
rect 10100 11068 10109 11108
rect 7459 11067 7517 11068
rect 3043 11024 3101 11025
rect 2467 10984 2476 11024
rect 2516 10984 3052 11024
rect 3092 10984 3532 11024
rect 3572 10984 3581 11024
rect 6211 10984 6220 11024
rect 6260 10984 6892 11024
rect 6932 10984 6941 11024
rect 9187 10984 9196 11024
rect 9236 10984 9580 11024
rect 9620 10984 10348 11024
rect 10388 10984 10397 11024
rect 13891 10984 13900 11024
rect 13940 10984 18700 11024
rect 18740 10984 18749 11024
rect 3043 10983 3101 10984
rect 8707 10940 8765 10941
rect 6115 10900 6124 10940
rect 6164 10900 6796 10940
rect 6836 10900 6845 10940
rect 8707 10900 8716 10940
rect 8756 10900 10828 10940
rect 10868 10900 10877 10940
rect 14755 10900 14764 10940
rect 14804 10900 15532 10940
rect 15572 10900 16108 10940
rect 16148 10900 16157 10940
rect 8707 10899 8765 10900
rect 0 10856 80 10876
rect 21424 10856 21504 10876
rect 0 10816 1324 10856
rect 1364 10816 1373 10856
rect 11203 10816 11212 10856
rect 11252 10816 11788 10856
rect 11828 10816 11837 10856
rect 12259 10816 12268 10856
rect 12308 10816 16972 10856
rect 17012 10816 17021 10856
rect 18019 10816 18028 10856
rect 18068 10816 18412 10856
rect 18452 10816 18461 10856
rect 20140 10816 21504 10856
rect 0 10796 80 10816
rect 20140 10772 20180 10816
rect 21424 10796 21504 10816
rect 3715 10732 3724 10772
rect 3764 10732 4204 10772
rect 4244 10732 4253 10772
rect 8419 10732 8428 10772
rect 8468 10732 8812 10772
rect 8852 10732 8861 10772
rect 11683 10732 11692 10772
rect 11732 10732 20180 10772
rect 4483 10688 4541 10689
rect 4398 10648 4492 10688
rect 4532 10648 10540 10688
rect 10580 10648 10589 10688
rect 14371 10648 14380 10688
rect 14420 10648 19660 10688
rect 19700 10648 19709 10688
rect 4483 10647 4541 10648
rect 8803 10604 8861 10605
rect 3679 10564 3688 10604
rect 3728 10564 3770 10604
rect 3810 10564 3852 10604
rect 3892 10564 3934 10604
rect 3974 10564 4016 10604
rect 4056 10564 4065 10604
rect 6595 10564 6604 10604
rect 6644 10564 6988 10604
rect 7028 10564 7037 10604
rect 8718 10564 8812 10604
rect 8852 10564 8861 10604
rect 8995 10564 9004 10604
rect 9044 10564 10156 10604
rect 10196 10564 11020 10604
rect 11060 10564 11069 10604
rect 13315 10564 13324 10604
rect 13364 10564 13373 10604
rect 13795 10564 13804 10604
rect 13844 10564 15148 10604
rect 15188 10564 15197 10604
rect 17923 10564 17932 10604
rect 17972 10564 18124 10604
rect 18164 10564 18173 10604
rect 18799 10564 18808 10604
rect 18848 10564 18890 10604
rect 18930 10564 18972 10604
rect 19012 10564 19054 10604
rect 19094 10564 19136 10604
rect 19176 10564 19185 10604
rect 8803 10563 8861 10564
rect 0 10520 80 10540
rect 13324 10520 13364 10564
rect 0 10480 2860 10520
rect 2900 10480 2909 10520
rect 8899 10480 8908 10520
rect 8948 10480 9580 10520
rect 9620 10480 9629 10520
rect 9964 10480 12268 10520
rect 12308 10480 12317 10520
rect 13324 10480 13516 10520
rect 13556 10480 13565 10520
rect 16195 10480 16204 10520
rect 16244 10480 18700 10520
rect 18740 10480 18749 10520
rect 0 10460 80 10480
rect 2755 10396 2764 10436
rect 2804 10396 3916 10436
rect 3956 10396 3965 10436
rect 4195 10396 4204 10436
rect 4244 10396 8812 10436
rect 8852 10396 8861 10436
rect 9964 10352 10004 10480
rect 14179 10436 14237 10437
rect 10051 10396 10060 10436
rect 10100 10396 11596 10436
rect 11636 10396 11645 10436
rect 13795 10396 13804 10436
rect 13844 10396 14188 10436
rect 14228 10396 14237 10436
rect 14467 10396 14476 10436
rect 14516 10396 14764 10436
rect 14804 10396 14813 10436
rect 16387 10396 16396 10436
rect 16436 10396 16684 10436
rect 16724 10396 16733 10436
rect 18499 10396 18508 10436
rect 18548 10396 20716 10436
rect 20756 10396 20765 10436
rect 14179 10395 14237 10396
rect 21424 10352 21504 10372
rect 1411 10312 1420 10352
rect 1460 10312 3532 10352
rect 3572 10312 5548 10352
rect 5588 10312 5597 10352
rect 6979 10312 6988 10352
rect 7028 10312 7180 10352
rect 7220 10312 7229 10352
rect 8611 10312 8620 10352
rect 8660 10312 8908 10352
rect 8948 10312 8957 10352
rect 9091 10312 9100 10352
rect 9140 10312 9964 10352
rect 10004 10312 10013 10352
rect 10531 10312 10540 10352
rect 10580 10312 21504 10352
rect 21424 10292 21504 10312
rect 7075 10268 7133 10269
rect 12931 10268 12989 10269
rect 14371 10268 14429 10269
rect 3811 10228 3820 10268
rect 3860 10228 4684 10268
rect 4724 10228 4733 10268
rect 5155 10228 5164 10268
rect 5204 10228 7084 10268
rect 7124 10228 7133 10268
rect 8323 10228 8332 10268
rect 8372 10228 9388 10268
rect 9428 10228 9676 10268
rect 9716 10228 9725 10268
rect 11320 10228 12172 10268
rect 12212 10228 12221 10268
rect 12846 10228 12940 10268
rect 12980 10228 12989 10268
rect 14275 10228 14284 10268
rect 14324 10228 14380 10268
rect 14420 10228 14429 10268
rect 15235 10228 15244 10268
rect 15284 10228 16012 10268
rect 16052 10228 19180 10268
rect 19220 10228 19229 10268
rect 0 10184 80 10204
rect 6796 10184 6836 10228
rect 7075 10227 7133 10228
rect 7459 10184 7517 10185
rect 0 10144 1420 10184
rect 1460 10144 1469 10184
rect 2371 10144 2380 10184
rect 2420 10144 5012 10184
rect 6787 10144 6796 10184
rect 6836 10144 6988 10184
rect 7028 10144 7037 10184
rect 7171 10144 7180 10184
rect 7220 10144 7468 10184
rect 7508 10144 7517 10184
rect 0 10124 80 10144
rect 4972 10100 5012 10144
rect 7459 10143 7517 10144
rect 8899 10184 8957 10185
rect 11320 10184 11360 10228
rect 12931 10227 12989 10228
rect 14371 10227 14429 10228
rect 8899 10144 8908 10184
rect 8948 10144 9292 10184
rect 9332 10144 9341 10184
rect 9475 10144 9484 10184
rect 9524 10144 11308 10184
rect 11348 10144 11360 10184
rect 13123 10144 13132 10184
rect 13172 10144 13900 10184
rect 13940 10144 13949 10184
rect 14179 10144 14188 10184
rect 14228 10144 17452 10184
rect 17492 10144 17501 10184
rect 18211 10144 18220 10184
rect 18260 10144 19948 10184
rect 19988 10144 19997 10184
rect 8899 10143 8957 10144
rect 20707 10100 20765 10101
rect 1891 10060 1900 10100
rect 1940 10060 2572 10100
rect 2612 10060 2860 10100
rect 2900 10060 2909 10100
rect 3715 10060 3724 10100
rect 3764 10060 4204 10100
rect 4244 10060 4253 10100
rect 4963 10060 4972 10100
rect 5012 10060 5021 10100
rect 6892 10060 18028 10100
rect 18068 10060 18077 10100
rect 18787 10060 18796 10100
rect 18836 10060 20716 10100
rect 20756 10060 20765 10100
rect 6892 10016 6932 10060
rect 20707 10059 20765 10060
rect 1603 9976 1612 10016
rect 1652 9976 6932 10016
rect 8419 9976 8428 10016
rect 8468 9976 10444 10016
rect 10484 9976 10493 10016
rect 10627 9976 10636 10016
rect 10676 9976 10685 10016
rect 16387 9976 16396 10016
rect 16436 9976 16588 10016
rect 16628 9976 16637 10016
rect 10636 9932 10676 9976
rect 2467 9892 2476 9932
rect 2516 9892 10676 9932
rect 15532 9892 16012 9932
rect 16052 9892 16061 9932
rect 0 9848 80 9868
rect 9571 9848 9629 9849
rect 0 9808 4684 9848
rect 4724 9808 4733 9848
rect 4919 9808 4928 9848
rect 4968 9808 5010 9848
rect 5050 9808 5092 9848
rect 5132 9808 5174 9848
rect 5214 9808 5256 9848
rect 5296 9808 5305 9848
rect 9475 9808 9484 9848
rect 9524 9808 9580 9848
rect 9620 9808 9629 9848
rect 0 9788 80 9808
rect 9571 9807 9629 9808
rect 15532 9764 15572 9892
rect 21424 9848 21504 9868
rect 15715 9808 15724 9848
rect 15764 9808 17836 9848
rect 17876 9808 17885 9848
rect 20039 9808 20048 9848
rect 20088 9808 20130 9848
rect 20170 9808 20212 9848
rect 20252 9808 20294 9848
rect 20334 9808 20376 9848
rect 20416 9808 20425 9848
rect 20524 9808 21504 9848
rect 20524 9764 20564 9808
rect 21424 9788 21504 9808
rect 2083 9724 2092 9764
rect 2132 9724 7180 9764
rect 7220 9724 7229 9764
rect 8707 9724 8716 9764
rect 8756 9724 15572 9764
rect 15619 9724 15628 9764
rect 15668 9724 20564 9764
rect 7843 9640 7852 9680
rect 7892 9640 11788 9680
rect 11828 9640 12172 9680
rect 12212 9640 12221 9680
rect 17155 9640 17164 9680
rect 17204 9640 17452 9680
rect 17492 9640 17501 9680
rect 19075 9640 19084 9680
rect 19124 9640 19756 9680
rect 19796 9640 19805 9680
rect 6211 9596 6269 9597
rect 2851 9556 2860 9596
rect 2900 9556 5452 9596
rect 5492 9556 5501 9596
rect 6211 9556 6220 9596
rect 6260 9556 12748 9596
rect 12788 9556 12797 9596
rect 6211 9555 6269 9556
rect 0 9512 80 9532
rect 3043 9512 3101 9513
rect 0 9472 2284 9512
rect 2324 9472 2333 9512
rect 2958 9472 3052 9512
rect 3092 9472 3101 9512
rect 3427 9472 3436 9512
rect 3476 9472 3724 9512
rect 3764 9472 3773 9512
rect 4483 9472 4492 9512
rect 4532 9472 4780 9512
rect 4820 9472 7852 9512
rect 7892 9472 7901 9512
rect 8227 9472 8236 9512
rect 8276 9472 8428 9512
rect 8468 9472 11596 9512
rect 11636 9472 11645 9512
rect 14275 9472 14284 9512
rect 14324 9472 15052 9512
rect 15092 9472 15101 9512
rect 16003 9472 16012 9512
rect 16052 9472 17644 9512
rect 17684 9472 17693 9512
rect 0 9452 80 9472
rect 3043 9471 3101 9472
rect 4291 9388 4300 9428
rect 4340 9388 8044 9428
rect 8084 9388 8093 9428
rect 11203 9388 11212 9428
rect 11252 9388 11788 9428
rect 11828 9388 12076 9428
rect 12116 9388 12125 9428
rect 15139 9388 15148 9428
rect 15188 9388 16108 9428
rect 16148 9388 16157 9428
rect 18019 9388 18028 9428
rect 18068 9388 19372 9428
rect 19412 9388 20180 9428
rect 3235 9344 3293 9345
rect 3139 9304 3148 9344
rect 3188 9304 3244 9344
rect 3284 9304 3293 9344
rect 3235 9303 3293 9304
rect 9379 9344 9437 9345
rect 20140 9344 20180 9388
rect 21424 9344 21504 9364
rect 9379 9304 9388 9344
rect 9428 9304 10540 9344
rect 10580 9304 10589 9344
rect 15523 9304 15532 9344
rect 15572 9304 15916 9344
rect 15956 9304 15965 9344
rect 20140 9304 21504 9344
rect 9379 9303 9437 9304
rect 21424 9284 21504 9304
rect 547 9220 556 9260
rect 596 9220 19372 9260
rect 19412 9220 19421 9260
rect 0 9176 80 9196
rect 20995 9176 21053 9177
rect 0 9136 2668 9176
rect 2708 9136 2717 9176
rect 4195 9136 4204 9176
rect 4244 9136 21004 9176
rect 21044 9136 21053 9176
rect 0 9116 80 9136
rect 20995 9135 21053 9136
rect 8515 9092 8573 9093
rect 15811 9092 15869 9093
rect 3679 9052 3688 9092
rect 3728 9052 3770 9092
rect 3810 9052 3852 9092
rect 3892 9052 3934 9092
rect 3974 9052 4016 9092
rect 4056 9052 4065 9092
rect 8515 9052 8524 9092
rect 8564 9052 13612 9092
rect 13652 9052 13661 9092
rect 14275 9052 14284 9092
rect 14324 9052 15820 9092
rect 15860 9052 15869 9092
rect 8515 9051 8573 9052
rect 15811 9051 15869 9052
rect 16003 9092 16061 9093
rect 16003 9052 16012 9092
rect 16052 9052 17452 9092
rect 17492 9052 17501 9092
rect 18799 9052 18808 9092
rect 18848 9052 18890 9092
rect 18930 9052 18972 9092
rect 19012 9052 19054 9092
rect 19094 9052 19136 9092
rect 19176 9052 19185 9092
rect 16003 9051 16061 9052
rect 16675 9008 16733 9009
rect 4675 8968 4684 9008
rect 4724 8968 14188 9008
rect 14228 8968 14237 9008
rect 15523 8968 15532 9008
rect 15572 8968 16012 9008
rect 16052 8968 16061 9008
rect 16590 8968 16684 9008
rect 16724 8968 16733 9008
rect 16675 8967 16733 8968
rect 18403 9008 18461 9009
rect 18403 8968 18412 9008
rect 18452 8968 18508 9008
rect 18548 8968 18557 9008
rect 18403 8967 18461 8968
rect 1987 8884 1996 8924
rect 2036 8884 2045 8924
rect 11683 8884 11692 8924
rect 11732 8884 20180 8924
rect 0 8840 80 8860
rect 1996 8840 2036 8884
rect 11971 8840 12029 8841
rect 16099 8840 16157 8841
rect 17539 8840 17597 8841
rect 19459 8840 19517 8841
rect 0 8800 1516 8840
rect 1556 8800 1565 8840
rect 1804 8800 2036 8840
rect 4675 8800 4684 8840
rect 4724 8800 5548 8840
rect 5588 8800 5597 8840
rect 5731 8800 5740 8840
rect 5780 8800 6220 8840
rect 6260 8800 6269 8840
rect 7075 8800 7084 8840
rect 7124 8800 8908 8840
rect 8948 8800 8957 8840
rect 11886 8800 11980 8840
rect 12020 8800 12029 8840
rect 12547 8800 12556 8840
rect 12596 8800 13036 8840
rect 13076 8800 13085 8840
rect 14851 8800 14860 8840
rect 14900 8800 15436 8840
rect 15476 8800 15485 8840
rect 15811 8800 15820 8840
rect 15860 8800 15869 8840
rect 16014 8800 16108 8840
rect 16148 8800 16157 8840
rect 17454 8800 17548 8840
rect 17588 8800 17597 8840
rect 17731 8800 17740 8840
rect 17780 8800 19468 8840
rect 19508 8800 19517 8840
rect 20140 8840 20180 8884
rect 21424 8840 21504 8860
rect 20140 8800 21504 8840
rect 0 8780 80 8800
rect 1804 8672 1844 8800
rect 11971 8799 12029 8800
rect 6211 8756 6269 8757
rect 11683 8756 11741 8757
rect 15820 8756 15860 8800
rect 16099 8799 16157 8800
rect 17539 8799 17597 8800
rect 19459 8799 19517 8800
rect 21424 8780 21504 8800
rect 1987 8716 1996 8756
rect 2036 8716 6220 8756
rect 6260 8716 6269 8756
rect 7843 8716 7852 8756
rect 7892 8716 8716 8756
rect 8756 8716 9868 8756
rect 9908 8716 9917 8756
rect 11587 8716 11596 8756
rect 11636 8716 11692 8756
rect 11732 8716 11741 8756
rect 12067 8716 12076 8756
rect 12116 8716 12844 8756
rect 12884 8716 14380 8756
rect 14420 8716 14429 8756
rect 15619 8716 15628 8756
rect 15668 8716 15860 8756
rect 16771 8756 16829 8757
rect 16771 8716 16780 8756
rect 16820 8716 18508 8756
rect 18548 8716 18557 8756
rect 6211 8715 6269 8716
rect 11683 8715 11741 8716
rect 16771 8715 16829 8716
rect 1795 8632 1804 8672
rect 1844 8632 1853 8672
rect 2500 8632 16916 8672
rect 17251 8632 17260 8672
rect 17300 8632 19276 8672
rect 19316 8632 19948 8672
rect 19988 8632 19997 8672
rect 2500 8588 2540 8632
rect 16675 8588 16733 8589
rect 2083 8548 2092 8588
rect 2132 8548 2540 8588
rect 2755 8548 2764 8588
rect 2804 8548 4780 8588
rect 4820 8548 4829 8588
rect 10627 8548 10636 8588
rect 10676 8548 11020 8588
rect 11060 8548 12076 8588
rect 12116 8548 12125 8588
rect 16675 8548 16684 8588
rect 16724 8548 16780 8588
rect 16820 8548 16829 8588
rect 16675 8547 16733 8548
rect 0 8504 80 8524
rect 16876 8504 16916 8632
rect 18211 8504 18269 8505
rect 0 8464 556 8504
rect 596 8464 605 8504
rect 6883 8464 6892 8504
rect 6932 8464 7468 8504
rect 7508 8464 10828 8504
rect 10868 8464 14668 8504
rect 14708 8464 14717 8504
rect 16867 8464 16876 8504
rect 16916 8464 16925 8504
rect 18126 8464 18220 8504
rect 18260 8464 18269 8504
rect 0 8444 80 8464
rect 18211 8463 18269 8464
rect 18403 8504 18461 8505
rect 18403 8464 18412 8504
rect 18452 8464 18508 8504
rect 18548 8464 18557 8504
rect 18403 8463 18461 8464
rect 19267 8420 19325 8421
rect 14563 8380 14572 8420
rect 14612 8380 15340 8420
rect 15380 8380 19276 8420
rect 19316 8380 19325 8420
rect 19267 8379 19325 8380
rect 21424 8336 21504 8356
rect 4919 8296 4928 8336
rect 4968 8296 5010 8336
rect 5050 8296 5092 8336
rect 5132 8296 5174 8336
rect 5214 8296 5256 8336
rect 5296 8296 5305 8336
rect 13411 8296 13420 8336
rect 13460 8296 18700 8336
rect 18740 8296 18749 8336
rect 20039 8296 20048 8336
rect 20088 8296 20130 8336
rect 20170 8296 20212 8336
rect 20252 8296 20294 8336
rect 20334 8296 20376 8336
rect 20416 8296 20425 8336
rect 20524 8296 21504 8336
rect 20524 8252 20564 8296
rect 21424 8276 21504 8296
rect 3235 8212 3244 8252
rect 3284 8212 4300 8252
rect 4340 8212 20564 8252
rect 0 8168 80 8188
rect 4195 8168 4253 8169
rect 4675 8168 4733 8169
rect 0 8128 1804 8168
rect 1844 8128 1853 8168
rect 4110 8128 4204 8168
rect 4244 8128 4684 8168
rect 4724 8128 4733 8168
rect 5731 8128 5740 8168
rect 5780 8128 6124 8168
rect 6164 8128 11596 8168
rect 11636 8128 11645 8168
rect 14659 8128 14668 8168
rect 14708 8128 16876 8168
rect 16916 8128 17356 8168
rect 17396 8128 17405 8168
rect 17635 8128 17644 8168
rect 17684 8128 17932 8168
rect 17972 8128 17981 8168
rect 18115 8128 18124 8168
rect 18164 8128 21484 8168
rect 0 8108 80 8128
rect 4195 8127 4253 8128
rect 4675 8127 4733 8128
rect 18124 8084 18164 8128
rect 10819 8044 10828 8084
rect 10868 8044 11116 8084
rect 11156 8044 11165 8084
rect 12835 8044 12844 8084
rect 12884 8044 12893 8084
rect 15052 8044 18164 8084
rect 4771 7960 4780 8000
rect 4820 7960 7372 8000
rect 7412 7960 9004 8000
rect 9044 7960 9053 8000
rect 12844 7916 12884 8044
rect 15052 8000 15092 8044
rect 18403 8000 18461 8001
rect 19267 8000 19325 8001
rect 21444 8000 21484 8128
rect 15043 7960 15052 8000
rect 15092 7960 15101 8000
rect 15235 7960 15244 8000
rect 15284 7960 15820 8000
rect 15860 7960 18316 8000
rect 18356 7960 18412 8000
rect 18452 7960 18461 8000
rect 19182 7960 19276 8000
rect 19316 7960 19325 8000
rect 18403 7959 18461 7960
rect 19267 7959 19325 7960
rect 21292 7960 21484 8000
rect 15235 7916 15293 7917
rect 1603 7876 1612 7916
rect 1652 7876 12884 7916
rect 14371 7876 14380 7916
rect 14420 7876 14860 7916
rect 14900 7876 15244 7916
rect 15284 7876 15916 7916
rect 15956 7876 17260 7916
rect 17300 7876 17309 7916
rect 18316 7876 18700 7916
rect 18740 7876 18749 7916
rect 15235 7875 15293 7876
rect 0 7832 80 7852
rect 18316 7832 18356 7876
rect 21292 7832 21332 7960
rect 21424 7832 21504 7852
rect 0 7792 1324 7832
rect 1364 7792 1373 7832
rect 3043 7792 3052 7832
rect 3092 7792 3436 7832
rect 3476 7792 5452 7832
rect 5492 7792 5501 7832
rect 9379 7792 9388 7832
rect 9428 7792 9580 7832
rect 9620 7792 9772 7832
rect 9812 7792 9821 7832
rect 18307 7792 18316 7832
rect 18356 7792 18365 7832
rect 21292 7792 21504 7832
rect 0 7772 80 7792
rect 21424 7772 21504 7792
rect 12259 7748 12317 7749
rect 2179 7708 2188 7748
rect 2228 7708 4108 7748
rect 4148 7708 4684 7748
rect 4724 7708 4733 7748
rect 7555 7708 7564 7748
rect 7604 7708 9964 7748
rect 10004 7708 10013 7748
rect 12174 7708 12268 7748
rect 12308 7708 12317 7748
rect 14083 7708 14092 7748
rect 14132 7708 15244 7748
rect 15284 7708 15293 7748
rect 17827 7708 17836 7748
rect 17876 7708 18796 7748
rect 18836 7708 18845 7748
rect 12259 7707 12317 7708
rect 11491 7664 11549 7665
rect 11491 7624 11500 7664
rect 11540 7624 13324 7664
rect 13364 7624 13373 7664
rect 14851 7624 14860 7664
rect 14900 7624 15436 7664
rect 15476 7624 15485 7664
rect 11491 7623 11549 7624
rect 11875 7580 11933 7581
rect 2467 7540 2476 7580
rect 2516 7540 2764 7580
rect 2804 7540 2813 7580
rect 3679 7540 3688 7580
rect 3728 7540 3770 7580
rect 3810 7540 3852 7580
rect 3892 7540 3934 7580
rect 3974 7540 4016 7580
rect 4056 7540 4065 7580
rect 8803 7540 8812 7580
rect 8852 7540 9388 7580
rect 9428 7540 10060 7580
rect 10100 7540 11692 7580
rect 11732 7540 11741 7580
rect 11875 7540 11884 7580
rect 11924 7540 12268 7580
rect 12308 7540 12317 7580
rect 18799 7540 18808 7580
rect 18848 7540 18890 7580
rect 18930 7540 18972 7580
rect 19012 7540 19054 7580
rect 19094 7540 19136 7580
rect 19176 7540 19185 7580
rect 11875 7539 11933 7540
rect 0 7496 80 7516
rect 0 7456 1804 7496
rect 1844 7456 1853 7496
rect 4483 7456 4492 7496
rect 4532 7456 4780 7496
rect 4820 7456 4829 7496
rect 6595 7456 6604 7496
rect 6644 7456 6892 7496
rect 6932 7456 6941 7496
rect 7555 7456 7564 7496
rect 7604 7456 9868 7496
rect 9908 7456 9917 7496
rect 17923 7456 17932 7496
rect 17972 7456 18124 7496
rect 18164 7456 18173 7496
rect 0 7436 80 7456
rect 1987 7372 1996 7412
rect 2036 7372 19948 7412
rect 19988 7372 19997 7412
rect 18211 7328 18269 7329
rect 4483 7288 4492 7328
rect 4532 7288 7948 7328
rect 7988 7288 7997 7328
rect 18115 7288 18124 7328
rect 18164 7288 18220 7328
rect 18260 7288 18269 7328
rect 18211 7287 18269 7288
rect 19267 7328 19325 7329
rect 19555 7328 19613 7329
rect 21424 7328 21504 7348
rect 19267 7288 19276 7328
rect 19316 7288 19564 7328
rect 19604 7288 21504 7328
rect 19267 7287 19325 7288
rect 19555 7287 19613 7288
rect 21424 7268 21504 7288
rect 4387 7244 4445 7245
rect 1603 7204 1612 7244
rect 1652 7204 4148 7244
rect 4302 7204 4396 7244
rect 4436 7204 4445 7244
rect 4963 7204 4972 7244
rect 5012 7204 5780 7244
rect 7843 7204 7852 7244
rect 7892 7204 8044 7244
rect 8084 7204 8093 7244
rect 8419 7204 8428 7244
rect 8468 7204 9196 7244
rect 9236 7204 9245 7244
rect 11320 7204 11788 7244
rect 11828 7204 12172 7244
rect 12212 7204 12221 7244
rect 16579 7204 16588 7244
rect 16628 7204 18028 7244
rect 18068 7204 18077 7244
rect 0 7160 80 7180
rect 4108 7160 4148 7204
rect 4387 7203 4445 7204
rect 5740 7160 5780 7204
rect 0 7120 2132 7160
rect 3523 7120 3532 7160
rect 3572 7120 3916 7160
rect 3956 7120 3965 7160
rect 4108 7120 5684 7160
rect 5740 7120 8812 7160
rect 8852 7120 8861 7160
rect 9859 7120 9868 7160
rect 9908 7120 10156 7160
rect 10196 7120 10444 7160
rect 10484 7120 10493 7160
rect 0 7100 80 7120
rect 2092 7076 2132 7120
rect 4387 7076 4445 7077
rect 2092 7036 4396 7076
rect 4436 7036 4445 7076
rect 4387 7035 4445 7036
rect 5644 6992 5684 7120
rect 11320 7076 11360 7204
rect 11587 7120 11596 7160
rect 11636 7120 12460 7160
rect 12500 7120 12509 7160
rect 12835 7120 12844 7160
rect 12884 7120 14380 7160
rect 14420 7120 14429 7160
rect 15427 7120 15436 7160
rect 15476 7120 16012 7160
rect 16052 7120 16061 7160
rect 16675 7120 16684 7160
rect 16724 7120 19372 7160
rect 19412 7120 19421 7160
rect 12259 7076 12317 7077
rect 9379 7036 9388 7076
rect 9428 7036 11360 7076
rect 12163 7036 12172 7076
rect 12212 7036 12268 7076
rect 12308 7036 12317 7076
rect 15139 7036 15148 7076
rect 15188 7036 16396 7076
rect 16436 7036 17068 7076
rect 17108 7036 18604 7076
rect 18644 7036 18653 7076
rect 12259 7035 12317 7036
rect 2179 6952 2188 6992
rect 2228 6952 2860 6992
rect 2900 6952 2909 6992
rect 3331 6952 3340 6992
rect 3380 6952 4972 6992
rect 5012 6952 5021 6992
rect 5635 6952 5644 6992
rect 5684 6952 5693 6992
rect 8035 6952 8044 6992
rect 8084 6952 8236 6992
rect 8276 6952 8285 6992
rect 8803 6952 8812 6992
rect 8852 6952 19564 6992
rect 19604 6952 19613 6992
rect 10243 6908 10301 6909
rect 1987 6868 1996 6908
rect 2036 6868 8428 6908
rect 8468 6868 8477 6908
rect 8899 6868 8908 6908
rect 8948 6868 10252 6908
rect 10292 6868 10301 6908
rect 12163 6868 12172 6908
rect 12212 6868 20564 6908
rect 10243 6867 10301 6868
rect 0 6824 80 6844
rect 20524 6824 20564 6868
rect 21424 6824 21504 6844
rect 0 6784 1516 6824
rect 1556 6784 1565 6824
rect 4919 6784 4928 6824
rect 4968 6784 5010 6824
rect 5050 6784 5092 6824
rect 5132 6784 5174 6824
rect 5214 6784 5256 6824
rect 5296 6784 5305 6824
rect 5644 6784 13228 6824
rect 13268 6784 13277 6824
rect 16387 6784 16396 6824
rect 16436 6784 16876 6824
rect 16916 6784 16925 6824
rect 20039 6784 20048 6824
rect 20088 6784 20130 6824
rect 20170 6784 20212 6824
rect 20252 6784 20294 6824
rect 20334 6784 20376 6824
rect 20416 6784 20425 6824
rect 20524 6784 21504 6824
rect 0 6764 80 6784
rect 5644 6740 5684 6784
rect 21424 6764 21504 6784
rect 172 6700 2956 6740
rect 2996 6700 3005 6740
rect 3811 6700 3820 6740
rect 3860 6700 4300 6740
rect 4340 6700 4349 6740
rect 5635 6700 5644 6740
rect 5684 6700 5693 6740
rect 5827 6700 5836 6740
rect 5876 6700 6316 6740
rect 6356 6700 6365 6740
rect 11320 6700 17740 6740
rect 17780 6700 17789 6740
rect 0 6488 80 6508
rect 0 6446 116 6488
rect 172 6446 212 6700
rect 11320 6656 11360 6700
rect 2083 6616 2092 6656
rect 2132 6616 11360 6656
rect 12547 6616 12556 6656
rect 12596 6616 13460 6656
rect 14659 6616 14668 6656
rect 14708 6616 15628 6656
rect 15668 6616 15677 6656
rect 13420 6572 13460 6616
rect 1795 6532 1804 6572
rect 1844 6532 2668 6572
rect 2708 6532 2717 6572
rect 3907 6532 3916 6572
rect 3956 6532 4588 6572
rect 4628 6532 9388 6572
rect 9428 6532 9620 6572
rect 9667 6532 9676 6572
rect 9716 6532 11788 6572
rect 11828 6532 11837 6572
rect 13027 6532 13036 6572
rect 13076 6532 13085 6572
rect 13420 6532 21484 6572
rect 9580 6488 9620 6532
rect 2755 6448 2764 6488
rect 2804 6448 4396 6488
rect 4436 6448 4445 6488
rect 5923 6448 5932 6488
rect 5972 6448 7564 6488
rect 7604 6448 7613 6488
rect 9571 6448 9580 6488
rect 9620 6448 9629 6488
rect 0 6428 212 6446
rect 76 6406 212 6428
rect 1699 6364 1708 6404
rect 1748 6364 1757 6404
rect 2275 6364 2284 6404
rect 2324 6364 2516 6404
rect 4003 6364 4012 6404
rect 4052 6364 4300 6404
rect 4340 6364 4349 6404
rect 1708 6236 1748 6364
rect 2476 6320 2516 6364
rect 13036 6320 13076 6532
rect 17059 6488 17117 6489
rect 21444 6488 21484 6532
rect 14467 6448 14476 6488
rect 14516 6448 14860 6488
rect 14900 6448 14909 6488
rect 16974 6448 17068 6488
rect 17108 6448 17117 6488
rect 17059 6447 17117 6448
rect 21388 6448 21484 6488
rect 21388 6340 21428 6448
rect 19939 6320 19997 6321
rect 2467 6280 2476 6320
rect 2516 6280 2525 6320
rect 2572 6280 13076 6320
rect 19854 6280 19948 6320
rect 19988 6280 19997 6320
rect 21388 6280 21504 6340
rect 2572 6236 2612 6280
rect 19939 6279 19997 6280
rect 21424 6260 21504 6280
rect 12067 6236 12125 6237
rect 1708 6196 2612 6236
rect 4483 6196 4492 6236
rect 4532 6196 6316 6236
rect 6356 6196 6892 6236
rect 6932 6196 6941 6236
rect 7459 6196 7468 6236
rect 7508 6196 9676 6236
rect 9716 6196 9725 6236
rect 12067 6196 12076 6236
rect 12116 6196 15820 6236
rect 15860 6196 16300 6236
rect 16340 6196 16349 6236
rect 12067 6195 12125 6196
rect 0 6152 80 6172
rect 0 6112 17356 6152
rect 17396 6112 17405 6152
rect 0 6092 80 6112
rect 3679 6028 3688 6068
rect 3728 6028 3770 6068
rect 3810 6028 3852 6068
rect 3892 6028 3934 6068
rect 3974 6028 4016 6068
rect 4056 6028 4065 6068
rect 6691 6028 6700 6068
rect 6740 6028 11596 6068
rect 11636 6028 11645 6068
rect 18799 6028 18808 6068
rect 18848 6028 18890 6068
rect 18930 6028 18972 6068
rect 19012 6028 19054 6068
rect 19094 6028 19136 6068
rect 19176 6028 19185 6068
rect 12931 5984 12989 5985
rect 2500 5944 12940 5984
rect 12980 5944 12989 5984
rect 2500 5900 2540 5944
rect 12931 5943 12989 5944
rect 2179 5860 2188 5900
rect 2228 5860 2540 5900
rect 5539 5860 5548 5900
rect 5588 5860 5932 5900
rect 5972 5860 5981 5900
rect 7363 5860 7372 5900
rect 7412 5860 7948 5900
rect 7988 5860 7997 5900
rect 8131 5860 8140 5900
rect 8180 5860 10156 5900
rect 10196 5860 10205 5900
rect 0 5816 80 5836
rect 21424 5816 21504 5836
rect 0 5776 8812 5816
rect 8852 5776 8861 5816
rect 14371 5776 14380 5816
rect 14420 5776 19756 5816
rect 19796 5776 21504 5816
rect 0 5756 80 5776
rect 21424 5756 21504 5776
rect 18211 5732 18269 5733
rect 1411 5692 1420 5732
rect 1460 5692 13900 5732
rect 13940 5692 13949 5732
rect 17539 5692 17548 5732
rect 17588 5692 17932 5732
rect 17972 5692 18220 5732
rect 18260 5692 18269 5732
rect 18211 5691 18269 5692
rect 10147 5648 10205 5649
rect 12931 5648 12989 5649
rect 1315 5608 1324 5648
rect 1364 5608 4492 5648
rect 4532 5608 4541 5648
rect 7555 5608 7564 5648
rect 7604 5608 8140 5648
rect 8180 5608 8189 5648
rect 9955 5608 9964 5648
rect 10004 5608 10156 5648
rect 10196 5608 11404 5648
rect 11444 5608 11453 5648
rect 11683 5608 11692 5648
rect 11732 5608 11741 5648
rect 12846 5608 12940 5648
rect 12980 5608 12989 5648
rect 13411 5608 13420 5648
rect 13460 5608 13556 5648
rect 16003 5608 16012 5648
rect 16052 5608 16972 5648
rect 17012 5608 18124 5648
rect 18164 5608 18173 5648
rect 10147 5607 10205 5608
rect 11692 5564 11732 5608
rect 12931 5607 12989 5608
rect 7939 5524 7948 5564
rect 7988 5524 8524 5564
rect 8564 5524 8573 5564
rect 9667 5524 9676 5564
rect 9716 5524 11732 5564
rect 0 5480 80 5500
rect 8524 5480 8564 5524
rect 12931 5480 12989 5481
rect 0 5440 1708 5480
rect 1748 5440 1757 5480
rect 8524 5440 11212 5480
rect 11252 5440 12940 5480
rect 12980 5440 12989 5480
rect 0 5420 80 5440
rect 12931 5439 12989 5440
rect 1987 5356 1996 5396
rect 2036 5356 8044 5396
rect 8084 5356 8093 5396
rect 13516 5312 13556 5608
rect 15811 5524 15820 5564
rect 15860 5524 17644 5564
rect 17684 5524 20180 5564
rect 15235 5480 15293 5481
rect 17059 5480 17117 5481
rect 15150 5440 15244 5480
rect 15284 5440 17068 5480
rect 17108 5440 17117 5480
rect 19939 5440 19948 5480
rect 19988 5440 19997 5480
rect 15235 5439 15293 5440
rect 17059 5439 17117 5440
rect 16483 5356 16492 5396
rect 16532 5356 17548 5396
rect 17588 5356 17597 5396
rect 4919 5272 4928 5312
rect 4968 5272 5010 5312
rect 5050 5272 5092 5312
rect 5132 5272 5174 5312
rect 5214 5272 5256 5312
rect 5296 5272 5305 5312
rect 11395 5272 11404 5312
rect 11444 5272 11692 5312
rect 11732 5272 11741 5312
rect 13507 5272 13516 5312
rect 13556 5272 13565 5312
rect 2467 5228 2525 5229
rect 19948 5228 19988 5440
rect 20140 5396 20180 5524
rect 20140 5356 21428 5396
rect 21388 5332 21428 5356
rect 20039 5272 20048 5312
rect 20088 5272 20130 5312
rect 20170 5272 20212 5312
rect 20252 5272 20294 5312
rect 20334 5272 20376 5312
rect 20416 5272 20425 5312
rect 21388 5272 21504 5332
rect 21424 5252 21504 5272
rect 2467 5188 2476 5228
rect 2516 5188 19988 5228
rect 2467 5187 2525 5188
rect 0 5144 80 5164
rect 0 5104 2284 5144
rect 2324 5104 2333 5144
rect 10723 5104 10732 5144
rect 10772 5104 16012 5144
rect 16052 5104 16061 5144
rect 0 5084 80 5104
rect 4483 5060 4541 5061
rect 12067 5060 12125 5061
rect 2467 5020 2476 5060
rect 2516 5020 3340 5060
rect 3380 5020 3389 5060
rect 3523 5020 3532 5060
rect 3572 5020 3916 5060
rect 3956 5020 3965 5060
rect 4099 5020 4108 5060
rect 4148 5020 4492 5060
rect 4532 5020 4541 5060
rect 5827 5020 5836 5060
rect 5876 5020 6124 5060
rect 6164 5020 7468 5060
rect 7508 5020 7517 5060
rect 11587 5020 11596 5060
rect 11636 5020 12076 5060
rect 12116 5020 12125 5060
rect 18211 5020 18220 5060
rect 18260 5020 18700 5060
rect 18740 5020 18749 5060
rect 4483 5019 4541 5020
rect 12067 5019 12125 5020
rect 67 4976 125 4977
rect 67 4936 76 4976
rect 116 4936 1324 4976
rect 1364 4936 1373 4976
rect 2083 4936 2092 4976
rect 2132 4936 2141 4976
rect 3043 4936 3052 4976
rect 3092 4936 5644 4976
rect 5684 4936 5693 4976
rect 6691 4936 6700 4976
rect 6740 4936 7084 4976
rect 7124 4936 7276 4976
rect 7316 4936 7325 4976
rect 7372 4936 8332 4976
rect 8372 4936 8381 4976
rect 9571 4936 9580 4976
rect 9620 4936 11020 4976
rect 11060 4936 11212 4976
rect 11252 4936 12748 4976
rect 12788 4936 12797 4976
rect 12931 4936 12940 4976
rect 12980 4936 13708 4976
rect 13748 4936 18604 4976
rect 18644 4936 18653 4976
rect 67 4935 125 4936
rect 2092 4892 2132 4936
rect 4291 4892 4349 4893
rect 7372 4892 7412 4936
rect 2092 4852 4300 4892
rect 4340 4852 7412 4892
rect 7747 4852 7756 4892
rect 7796 4852 9772 4892
rect 9812 4852 9821 4892
rect 13891 4852 13900 4892
rect 13940 4852 20524 4892
rect 20564 4852 20573 4892
rect 4291 4851 4349 4852
rect 0 4808 80 4828
rect 2467 4808 2525 4809
rect 14947 4808 15005 4809
rect 21424 4808 21504 4828
rect 0 4768 2476 4808
rect 2516 4768 2525 4808
rect 3043 4768 3052 4808
rect 3092 4768 3628 4808
rect 3668 4768 3677 4808
rect 4195 4768 4204 4808
rect 4244 4768 4396 4808
rect 4436 4768 8428 4808
rect 8468 4768 8477 4808
rect 14755 4768 14764 4808
rect 14804 4768 14956 4808
rect 14996 4768 15005 4808
rect 17827 4768 17836 4808
rect 17876 4768 19852 4808
rect 19892 4768 19901 4808
rect 21379 4768 21388 4808
rect 21428 4768 21504 4808
rect 0 4748 80 4768
rect 2467 4767 2525 4768
rect 14947 4767 15005 4768
rect 21424 4748 21504 4768
rect 18403 4724 18461 4725
rect 3523 4684 3532 4724
rect 3572 4684 4492 4724
rect 4532 4684 4541 4724
rect 7939 4684 7948 4724
rect 7988 4684 18412 4724
rect 18452 4684 18461 4724
rect 18403 4683 18461 4684
rect 1315 4600 1324 4640
rect 1364 4600 4204 4640
rect 4244 4600 4253 4640
rect 5635 4600 5644 4640
rect 5684 4600 5932 4640
rect 5972 4600 9964 4640
rect 10004 4600 10013 4640
rect 3679 4516 3688 4556
rect 3728 4516 3770 4556
rect 3810 4516 3852 4556
rect 3892 4516 3934 4556
rect 3974 4516 4016 4556
rect 4056 4516 4065 4556
rect 4291 4516 4300 4556
rect 4340 4516 4492 4556
rect 4532 4516 13900 4556
rect 13940 4516 13949 4556
rect 14371 4516 14380 4556
rect 14420 4516 15148 4556
rect 15188 4516 15197 4556
rect 18799 4516 18808 4556
rect 18848 4516 18890 4556
rect 18930 4516 18972 4556
rect 19012 4516 19054 4556
rect 19094 4516 19136 4556
rect 19176 4516 19185 4556
rect 0 4472 80 4492
rect 0 4432 17740 4472
rect 17780 4432 17789 4472
rect 20428 4432 21388 4472
rect 21428 4432 21437 4472
rect 0 4412 80 4432
rect 4099 4388 4157 4389
rect 4014 4348 4108 4388
rect 4148 4348 4157 4388
rect 4099 4347 4157 4348
rect 4204 4348 5740 4388
rect 5780 4348 5789 4388
rect 7075 4348 7084 4388
rect 7124 4348 7564 4388
rect 7604 4348 7613 4388
rect 11395 4348 11404 4388
rect 11444 4348 11692 4388
rect 11732 4348 11741 4388
rect 14371 4348 14380 4388
rect 14420 4348 15052 4388
rect 15092 4348 15101 4388
rect 16099 4348 16108 4388
rect 16148 4348 17164 4388
rect 17204 4348 18796 4388
rect 18836 4348 18845 4388
rect 4204 4304 4244 4348
rect 20428 4304 20468 4432
rect 21424 4304 21504 4324
rect 2860 4264 3052 4304
rect 3092 4264 4244 4304
rect 4291 4264 4300 4304
rect 4340 4264 5644 4304
rect 5684 4264 5693 4304
rect 5923 4264 5932 4304
rect 5972 4264 6604 4304
rect 6644 4264 7852 4304
rect 7892 4264 7901 4304
rect 10435 4264 10444 4304
rect 10484 4264 11212 4304
rect 11252 4264 20468 4304
rect 20515 4264 20524 4304
rect 20564 4264 21504 4304
rect 0 4136 80 4156
rect 2860 4137 2900 4264
rect 21424 4244 21504 4264
rect 3139 4180 3148 4220
rect 3188 4180 4108 4220
rect 4148 4180 4157 4220
rect 5059 4180 5068 4220
rect 5108 4180 11884 4220
rect 11924 4180 11933 4220
rect 15436 4180 16108 4220
rect 16148 4180 16157 4220
rect 16483 4180 16492 4220
rect 16532 4180 16684 4220
rect 16724 4180 16733 4220
rect 17539 4180 17548 4220
rect 17588 4180 19948 4220
rect 19988 4180 19997 4220
rect 2851 4136 2909 4137
rect 0 4096 1900 4136
rect 1940 4096 1949 4136
rect 2467 4096 2476 4136
rect 2516 4096 2860 4136
rect 2900 4096 2909 4136
rect 4108 4136 4148 4180
rect 15436 4136 15476 4180
rect 4108 4096 7220 4136
rect 9763 4096 9772 4136
rect 9812 4096 10156 4136
rect 10196 4096 10205 4136
rect 12739 4096 12748 4136
rect 12788 4096 14476 4136
rect 14516 4096 14525 4136
rect 15427 4096 15436 4136
rect 15476 4096 15485 4136
rect 16003 4096 16012 4136
rect 16052 4096 16780 4136
rect 16820 4096 17740 4136
rect 17780 4096 19276 4136
rect 19316 4096 19325 4136
rect 0 4076 80 4096
rect 2851 4095 2909 4096
rect 7180 4052 7220 4096
rect 19651 4052 19709 4053
rect 2659 4012 2668 4052
rect 2708 4012 4588 4052
rect 4628 4012 4637 4052
rect 7171 4012 7180 4052
rect 7220 4012 7229 4052
rect 15523 4012 15532 4052
rect 15572 4012 18316 4052
rect 18356 4012 18365 4052
rect 18499 4012 18508 4052
rect 18548 4012 19660 4052
rect 19700 4012 19709 4052
rect 19651 4011 19709 4012
rect 4291 3968 4349 3969
rect 1507 3928 1516 3968
rect 1556 3928 2860 3968
rect 2900 3928 2909 3968
rect 4099 3928 4108 3968
rect 4148 3928 4300 3968
rect 4340 3928 4684 3968
rect 4724 3928 4733 3968
rect 4867 3928 4876 3968
rect 4916 3928 4925 3968
rect 8419 3928 8428 3968
rect 8468 3928 12556 3968
rect 12596 3928 12605 3968
rect 13219 3928 13228 3968
rect 13268 3928 13996 3968
rect 14036 3928 18604 3968
rect 18644 3928 18653 3968
rect 4291 3927 4349 3928
rect 4876 3884 4916 3928
rect 355 3844 364 3884
rect 404 3844 4916 3884
rect 18403 3884 18461 3885
rect 18403 3844 18412 3884
rect 18452 3844 20564 3884
rect 18403 3843 18461 3844
rect 0 3800 80 3820
rect 2851 3800 2909 3801
rect 20524 3800 20564 3844
rect 21424 3800 21504 3820
rect 0 3760 2188 3800
rect 2228 3760 2237 3800
rect 2851 3760 2860 3800
rect 2900 3760 2956 3800
rect 2996 3760 3005 3800
rect 3331 3760 3340 3800
rect 3380 3760 4396 3800
rect 4436 3760 4445 3800
rect 4919 3760 4928 3800
rect 4968 3760 5010 3800
rect 5050 3760 5092 3800
rect 5132 3760 5174 3800
rect 5214 3760 5256 3800
rect 5296 3760 5305 3800
rect 20039 3760 20048 3800
rect 20088 3760 20130 3800
rect 20170 3760 20212 3800
rect 20252 3760 20294 3800
rect 20334 3760 20376 3800
rect 20416 3760 20425 3800
rect 20524 3760 21504 3800
rect 0 3740 80 3760
rect 2851 3759 2909 3760
rect 21424 3740 21504 3760
rect 12931 3716 12989 3717
rect 5443 3676 5452 3716
rect 5492 3676 5740 3716
rect 5780 3676 5789 3716
rect 12931 3676 12940 3716
rect 12980 3676 14764 3716
rect 14804 3676 17836 3716
rect 17876 3676 18028 3716
rect 18068 3676 18077 3716
rect 12931 3675 12989 3676
rect 2467 3592 2476 3632
rect 2516 3592 16684 3632
rect 16724 3592 16733 3632
rect 19459 3592 19468 3632
rect 19508 3592 20044 3632
rect 20084 3592 20093 3632
rect 6019 3508 6028 3548
rect 6068 3508 6796 3548
rect 6836 3508 6845 3548
rect 17923 3508 17932 3548
rect 17972 3508 18412 3548
rect 18452 3508 18461 3548
rect 0 3464 80 3484
rect 19267 3464 19325 3465
rect 0 3424 2284 3464
rect 2324 3424 2333 3464
rect 4387 3424 4396 3464
rect 4436 3424 5548 3464
rect 5588 3424 5597 3464
rect 6403 3424 6412 3464
rect 6452 3424 7468 3464
rect 7508 3424 7517 3464
rect 8800 3424 9004 3464
rect 9044 3424 10828 3464
rect 10868 3424 10877 3464
rect 16771 3424 16780 3464
rect 16820 3424 16972 3464
rect 17012 3424 17021 3464
rect 17251 3424 17260 3464
rect 17300 3424 19276 3464
rect 19316 3424 19325 3464
rect 0 3404 80 3424
rect 8800 3380 8840 3424
rect 15427 3380 15485 3381
rect 7267 3340 7276 3380
rect 7316 3340 8840 3380
rect 9859 3340 9868 3380
rect 9908 3340 11788 3380
rect 11828 3340 11837 3380
rect 15342 3340 15436 3380
rect 15476 3340 15485 3380
rect 15427 3339 15485 3340
rect 14947 3296 15005 3297
rect 16972 3296 17012 3424
rect 19267 3423 19325 3424
rect 19747 3340 19756 3380
rect 19796 3340 19948 3380
rect 19988 3340 19997 3380
rect 21424 3296 21504 3316
rect 14179 3256 14188 3296
rect 14228 3256 14804 3296
rect 14764 3212 14804 3256
rect 14947 3256 14956 3296
rect 14996 3256 15090 3296
rect 16972 3256 21504 3296
rect 14947 3255 15005 3256
rect 21424 3236 21504 3256
rect 1507 3172 1516 3212
rect 1556 3172 1565 3212
rect 2500 3172 13420 3212
rect 13460 3172 13469 3212
rect 14755 3172 14764 3212
rect 14804 3172 14813 3212
rect 0 3128 80 3148
rect 1516 3128 1556 3172
rect 2500 3128 2540 3172
rect 0 3088 1556 3128
rect 2371 3088 2380 3128
rect 2420 3088 2540 3128
rect 11395 3088 11404 3128
rect 11444 3088 15436 3128
rect 15476 3088 15485 3128
rect 0 3068 80 3088
rect 3679 3004 3688 3044
rect 3728 3004 3770 3044
rect 3810 3004 3852 3044
rect 3892 3004 3934 3044
rect 3974 3004 4016 3044
rect 4056 3004 4065 3044
rect 18799 3004 18808 3044
rect 18848 3004 18890 3044
rect 18930 3004 18972 3044
rect 19012 3004 19054 3044
rect 19094 3004 19136 3044
rect 19176 3004 19185 3044
rect 4108 2920 4780 2960
rect 4820 2920 12364 2960
rect 12404 2920 12413 2960
rect 4108 2876 4148 2920
rect 7651 2876 7709 2877
rect 8035 2876 8093 2877
rect 4099 2836 4108 2876
rect 4148 2836 4157 2876
rect 5923 2836 5932 2876
rect 5972 2836 6508 2876
rect 6548 2836 6557 2876
rect 7566 2836 7660 2876
rect 7700 2836 7709 2876
rect 7950 2836 8044 2876
rect 8084 2836 8093 2876
rect 19555 2836 19564 2876
rect 19604 2836 20044 2876
rect 20084 2836 20093 2876
rect 7651 2835 7709 2836
rect 8035 2835 8093 2836
rect 0 2792 80 2812
rect 21424 2792 21504 2812
rect 0 2752 1900 2792
rect 1940 2752 1949 2792
rect 3139 2752 3148 2792
rect 3188 2752 4492 2792
rect 4532 2752 4541 2792
rect 5164 2752 14380 2792
rect 14420 2752 14429 2792
rect 15427 2752 15436 2792
rect 15476 2752 21504 2792
rect 0 2732 80 2752
rect 5164 2708 5204 2752
rect 21424 2732 21504 2752
rect 9763 2708 9821 2709
rect 11395 2708 11453 2709
rect 13699 2708 13757 2709
rect 2467 2668 2476 2708
rect 2516 2668 4780 2708
rect 4820 2668 4829 2708
rect 5155 2668 5164 2708
rect 5204 2668 5213 2708
rect 5539 2668 5548 2708
rect 5588 2668 5836 2708
rect 5876 2668 5885 2708
rect 9678 2668 9772 2708
rect 9812 2668 9821 2708
rect 11107 2668 11116 2708
rect 11156 2668 11404 2708
rect 11444 2668 11453 2708
rect 12739 2668 12748 2708
rect 12788 2668 13132 2708
rect 13172 2668 13181 2708
rect 13614 2668 13708 2708
rect 13748 2668 13757 2708
rect 9763 2667 9821 2668
rect 11395 2667 11453 2668
rect 4099 2624 4157 2625
rect 8227 2624 8285 2625
rect 12163 2624 12221 2625
rect 3619 2584 3628 2624
rect 3668 2584 4108 2624
rect 4148 2584 4157 2624
rect 4483 2584 4492 2624
rect 4532 2584 5452 2624
rect 5492 2584 5501 2624
rect 5635 2584 5644 2624
rect 5684 2584 5932 2624
rect 5972 2584 5981 2624
rect 8227 2584 8236 2624
rect 8276 2584 8756 2624
rect 4099 2583 4157 2584
rect 8227 2583 8285 2584
rect 8716 2540 8756 2584
rect 11320 2584 12172 2624
rect 12212 2584 12221 2624
rect 1987 2500 1996 2540
rect 2036 2500 2380 2540
rect 2420 2500 2429 2540
rect 3427 2500 3436 2540
rect 3476 2500 3724 2540
rect 3764 2500 3773 2540
rect 4195 2500 4204 2540
rect 4244 2500 4876 2540
rect 4916 2500 4925 2540
rect 8707 2500 8716 2540
rect 8756 2500 8765 2540
rect 10147 2500 10156 2540
rect 10196 2500 10205 2540
rect 0 2456 80 2476
rect 0 2416 1516 2456
rect 1556 2416 1565 2456
rect 1795 2416 1804 2456
rect 1844 2416 5548 2456
rect 5588 2416 5597 2456
rect 8611 2416 8620 2456
rect 8660 2416 9292 2456
rect 9332 2416 9341 2456
rect 0 2396 80 2416
rect 10156 2372 10196 2500
rect 11320 2456 11360 2584
rect 12163 2583 12221 2584
rect 13132 2624 13172 2668
rect 13699 2667 13757 2668
rect 13987 2708 14045 2709
rect 14467 2708 14525 2709
rect 14851 2708 14909 2709
rect 16099 2708 16157 2709
rect 13987 2668 13996 2708
rect 14036 2668 14092 2708
rect 14132 2668 14141 2708
rect 14382 2668 14476 2708
rect 14516 2668 14525 2708
rect 14766 2668 14860 2708
rect 14900 2668 14909 2708
rect 15331 2668 15340 2708
rect 15380 2668 16108 2708
rect 16148 2668 18604 2708
rect 18644 2668 18653 2708
rect 13987 2667 14045 2668
rect 14467 2667 14525 2668
rect 14851 2667 14909 2668
rect 16099 2667 16157 2668
rect 13132 2584 16588 2624
rect 16628 2584 18220 2624
rect 18260 2584 18269 2624
rect 11011 2416 11020 2456
rect 11060 2416 11360 2456
rect 1411 2332 1420 2372
rect 1460 2332 2092 2372
rect 2132 2332 2141 2372
rect 2947 2332 2956 2372
rect 2996 2332 3148 2372
rect 3188 2332 6412 2372
rect 6452 2332 6461 2372
rect 8707 2332 8716 2372
rect 8756 2332 10196 2372
rect 13132 2372 13172 2584
rect 16684 2540 16724 2584
rect 16675 2500 16684 2540
rect 16724 2500 16733 2540
rect 13795 2416 13804 2456
rect 13844 2416 14284 2456
rect 14324 2416 14333 2456
rect 14659 2416 14668 2456
rect 14708 2416 14717 2456
rect 14668 2372 14708 2416
rect 13132 2332 13708 2372
rect 13748 2332 13757 2372
rect 13987 2332 13996 2372
rect 14036 2332 14708 2372
rect 16771 2288 16829 2289
rect 4919 2248 4928 2288
rect 4968 2248 5010 2288
rect 5050 2248 5092 2288
rect 5132 2248 5174 2288
rect 5214 2248 5256 2288
rect 5296 2248 5305 2288
rect 6892 2248 8236 2288
rect 8276 2248 8285 2288
rect 9571 2248 9580 2288
rect 9620 2248 10156 2288
rect 10196 2248 10205 2288
rect 12451 2248 12460 2288
rect 12500 2248 16780 2288
rect 16820 2248 16829 2288
rect 20039 2248 20048 2288
rect 20088 2248 20130 2288
rect 20170 2248 20212 2288
rect 20252 2248 20294 2288
rect 20334 2248 20376 2288
rect 20416 2248 20425 2288
rect 6892 2205 6932 2248
rect 16771 2247 16829 2248
rect 6883 2204 6941 2205
rect 2563 2164 2572 2204
rect 2612 2164 6892 2204
rect 6932 2164 6941 2204
rect 7651 2164 7660 2204
rect 7700 2164 8140 2204
rect 8180 2164 8189 2204
rect 13315 2164 13324 2204
rect 13364 2164 13900 2204
rect 13940 2164 13949 2204
rect 6883 2163 6941 2164
rect 0 2120 80 2140
rect 0 2080 1900 2120
rect 1940 2080 1949 2120
rect 2467 2080 2476 2120
rect 2516 2080 12748 2120
rect 12788 2080 12797 2120
rect 0 2060 80 2080
rect 2371 2036 2429 2037
rect 2371 1996 2380 2036
rect 2420 1996 4876 2036
rect 4916 1996 4925 2036
rect 6508 1996 16588 2036
rect 16628 1996 16637 2036
rect 2371 1995 2429 1996
rect 2659 1912 2668 1952
rect 2708 1912 4396 1952
rect 4436 1912 4445 1952
rect 0 1784 80 1804
rect 6508 1784 6548 1996
rect 9187 1952 9245 1953
rect 9102 1912 9196 1952
rect 9236 1912 9245 1952
rect 9187 1911 9245 1912
rect 9955 1952 10013 1953
rect 15331 1952 15389 1953
rect 16771 1952 16829 1953
rect 9955 1912 9964 1952
rect 10004 1912 10252 1952
rect 10292 1912 10301 1952
rect 13603 1912 13612 1952
rect 13652 1912 15148 1952
rect 15188 1912 15197 1952
rect 15331 1912 15340 1952
rect 15380 1912 15474 1952
rect 16686 1912 16780 1952
rect 16820 1912 16829 1952
rect 9955 1911 10013 1912
rect 15331 1911 15389 1912
rect 16771 1911 16829 1912
rect 10051 1868 10109 1869
rect 10435 1868 10493 1869
rect 11299 1868 11357 1869
rect 11587 1868 11645 1869
rect 15043 1868 15101 1869
rect 9966 1828 10060 1868
rect 10100 1828 10109 1868
rect 10350 1828 10444 1868
rect 10484 1828 10493 1868
rect 11203 1828 11212 1868
rect 11252 1828 11308 1868
rect 11348 1828 11357 1868
rect 11502 1828 11596 1868
rect 11636 1828 11645 1868
rect 14083 1828 14092 1868
rect 14132 1828 14284 1868
rect 14324 1828 15052 1868
rect 15092 1828 15101 1868
rect 16291 1828 16300 1868
rect 16340 1828 16876 1868
rect 16916 1828 16925 1868
rect 10051 1827 10109 1828
rect 10435 1827 10493 1828
rect 11299 1827 11357 1828
rect 11587 1827 11645 1828
rect 15043 1827 15101 1828
rect 17059 1784 17117 1785
rect 0 1744 1516 1784
rect 1556 1744 1565 1784
rect 3715 1744 3724 1784
rect 3764 1744 6548 1784
rect 13891 1744 13900 1784
rect 13940 1744 14860 1784
rect 14900 1744 14909 1784
rect 16579 1744 16588 1784
rect 16628 1744 17068 1784
rect 17108 1744 17117 1784
rect 0 1724 80 1744
rect 17059 1743 17117 1744
rect 2851 1660 2860 1700
rect 2900 1660 9100 1700
rect 9140 1660 9149 1700
rect 9859 1660 9868 1700
rect 9908 1660 10828 1700
rect 10868 1660 10877 1700
rect 12643 1660 12652 1700
rect 12692 1660 14380 1700
rect 14420 1660 14429 1700
rect 14563 1660 14572 1700
rect 14612 1660 15340 1700
rect 15380 1660 15389 1700
rect 16771 1660 16780 1700
rect 16820 1660 18028 1700
rect 18068 1660 18077 1700
rect 4675 1616 4733 1617
rect 1411 1576 1420 1616
rect 1460 1576 4684 1616
rect 4724 1576 4733 1616
rect 4675 1575 4733 1576
rect 4780 1576 7028 1616
rect 10051 1576 10060 1616
rect 10100 1576 10732 1616
rect 10772 1576 10781 1616
rect 4780 1532 4820 1576
rect 3679 1492 3688 1532
rect 3728 1492 3770 1532
rect 3810 1492 3852 1532
rect 3892 1492 3934 1532
rect 3974 1492 4016 1532
rect 4056 1492 4065 1532
rect 4204 1492 4820 1532
rect 6988 1532 7028 1576
rect 6988 1492 14956 1532
rect 14996 1492 15005 1532
rect 18799 1492 18808 1532
rect 18848 1492 18890 1532
rect 18930 1492 18972 1532
rect 19012 1492 19054 1532
rect 19094 1492 19136 1532
rect 19176 1492 19185 1532
rect 0 1448 80 1468
rect 0 1408 2284 1448
rect 2324 1408 2333 1448
rect 0 1388 80 1408
rect 4204 1364 4244 1492
rect 4291 1408 4300 1448
rect 4340 1408 5932 1448
rect 5972 1408 6604 1448
rect 6644 1408 16012 1448
rect 16052 1408 16061 1448
rect 8515 1364 8573 1365
rect 20611 1364 20669 1365
rect 2179 1324 2188 1364
rect 2228 1324 4244 1364
rect 7651 1324 7660 1364
rect 7700 1324 7988 1364
rect 8430 1324 8524 1364
rect 8564 1324 8573 1364
rect 10723 1324 10732 1364
rect 10772 1324 12076 1364
rect 12116 1324 12125 1364
rect 18883 1324 18892 1364
rect 18932 1324 20620 1364
rect 20660 1324 20669 1364
rect 2755 1280 2813 1281
rect 2670 1240 2764 1280
rect 2804 1240 2813 1280
rect 2755 1239 2813 1240
rect 2947 1280 3005 1281
rect 3139 1280 3197 1281
rect 3523 1280 3581 1281
rect 6403 1280 6461 1281
rect 6979 1280 7037 1281
rect 7843 1280 7901 1281
rect 2947 1240 2956 1280
rect 2996 1240 3090 1280
rect 3139 1240 3148 1280
rect 3188 1240 3282 1280
rect 3438 1240 3532 1280
rect 3572 1240 3581 1280
rect 6318 1240 6412 1280
rect 6452 1240 6461 1280
rect 6894 1240 6988 1280
rect 7028 1240 7037 1280
rect 7758 1240 7852 1280
rect 7892 1240 7901 1280
rect 7948 1280 7988 1324
rect 8515 1323 8573 1324
rect 20611 1323 20669 1324
rect 7948 1240 9484 1280
rect 9524 1240 9533 1280
rect 10627 1240 10636 1280
rect 10676 1240 11788 1280
rect 11828 1240 11837 1280
rect 15139 1240 15148 1280
rect 15188 1240 15436 1280
rect 15476 1240 18508 1280
rect 18548 1240 18557 1280
rect 19075 1240 19084 1280
rect 19124 1240 20620 1280
rect 20660 1240 20669 1280
rect 2947 1239 3005 1240
rect 3139 1239 3197 1240
rect 3523 1239 3581 1240
rect 6403 1239 6461 1240
rect 6979 1239 7037 1240
rect 7843 1239 7901 1240
rect 2275 1196 2333 1197
rect 6691 1196 6749 1197
rect 8611 1196 8669 1197
rect 10819 1196 10877 1197
rect 11203 1196 11261 1197
rect 12643 1196 12701 1197
rect 13027 1196 13085 1197
rect 13411 1196 13469 1197
rect 13795 1196 13853 1197
rect 17251 1196 17309 1197
rect 20515 1196 20573 1197
rect 2275 1156 2284 1196
rect 2324 1156 3916 1196
rect 3956 1156 3965 1196
rect 6691 1156 6700 1196
rect 6740 1156 7372 1196
rect 7412 1156 7421 1196
rect 7939 1156 7948 1196
rect 7988 1156 8620 1196
rect 8660 1156 8669 1196
rect 10734 1156 10828 1196
rect 10868 1156 10877 1196
rect 11118 1156 11212 1196
rect 11252 1156 11261 1196
rect 12558 1156 12652 1196
rect 12692 1156 12701 1196
rect 12942 1156 13036 1196
rect 13076 1156 13085 1196
rect 13326 1156 13420 1196
rect 13460 1156 13469 1196
rect 13710 1156 13804 1196
rect 13844 1156 13853 1196
rect 14755 1156 14764 1196
rect 14804 1156 15052 1196
rect 15092 1156 15101 1196
rect 17251 1156 17260 1196
rect 17300 1156 17356 1196
rect 17396 1156 17405 1196
rect 17731 1156 17740 1196
rect 17780 1156 20524 1196
rect 20564 1156 20573 1196
rect 2275 1155 2333 1156
rect 6691 1155 6749 1156
rect 8611 1155 8669 1156
rect 10819 1155 10877 1156
rect 11203 1155 11261 1156
rect 12643 1155 12701 1156
rect 13027 1155 13085 1156
rect 13411 1155 13469 1156
rect 13795 1155 13853 1156
rect 17251 1155 17309 1156
rect 20515 1155 20573 1156
rect 0 1112 80 1132
rect 1123 1112 1181 1113
rect 0 1072 364 1112
rect 404 1072 413 1112
rect 1123 1072 1132 1112
rect 1172 1072 4300 1112
rect 4340 1072 4349 1112
rect 5059 1072 5068 1112
rect 5108 1072 9388 1112
rect 9428 1072 9437 1112
rect 10243 1072 10252 1112
rect 10292 1072 11308 1112
rect 11348 1072 11357 1112
rect 16675 1072 16684 1112
rect 16724 1072 16972 1112
rect 17012 1072 17021 1112
rect 0 1052 80 1072
rect 1123 1071 1181 1072
rect 1699 988 1708 1028
rect 1748 988 17932 1028
rect 17972 988 17981 1028
rect 6595 944 6653 945
rect 17539 944 17597 945
rect 4483 904 4492 944
rect 4532 904 5260 944
rect 5300 904 5309 944
rect 6510 904 6604 944
rect 6644 904 6653 944
rect 7651 904 7660 944
rect 7700 904 8716 944
rect 8756 904 8765 944
rect 10627 904 10636 944
rect 10676 904 11212 944
rect 11252 904 11261 944
rect 11395 904 11404 944
rect 11444 904 11980 944
rect 12020 904 12029 944
rect 12547 904 12556 944
rect 12596 904 13228 944
rect 13268 904 13277 944
rect 13507 904 13516 944
rect 13556 904 14092 944
rect 14132 904 14141 944
rect 15139 904 15148 944
rect 15188 904 17164 944
rect 17204 904 17213 944
rect 17347 904 17356 944
rect 17396 904 17548 944
rect 17588 904 17597 944
rect 6595 903 6653 904
rect 17539 903 17597 904
rect 15139 860 15197 861
rect 4099 820 4108 860
rect 4148 820 8620 860
rect 8660 820 8669 860
rect 10435 820 10444 860
rect 10484 820 10924 860
rect 10964 820 10973 860
rect 11491 820 11500 860
rect 11540 820 12172 860
rect 12212 820 12221 860
rect 14659 820 14668 860
rect 14708 820 15148 860
rect 15188 820 15197 860
rect 15139 819 15197 820
rect 17443 860 17501 861
rect 17443 820 17452 860
rect 17492 820 17548 860
rect 17588 820 17597 860
rect 17443 819 17501 820
rect 0 776 80 796
rect 6787 776 6845 777
rect 0 736 3340 776
rect 3380 736 3389 776
rect 4919 736 4928 776
rect 4968 736 5010 776
rect 5050 736 5092 776
rect 5132 736 5174 776
rect 5214 736 5256 776
rect 5296 736 5305 776
rect 5347 736 5356 776
rect 5396 736 6068 776
rect 6702 736 6796 776
rect 6836 736 6845 776
rect 0 716 80 736
rect 4675 692 4733 693
rect 5356 692 5396 736
rect 5923 692 5981 693
rect 2371 652 2380 692
rect 2420 652 4628 692
rect 1027 608 1085 609
rect 4588 608 4628 652
rect 4675 652 4684 692
rect 4724 652 5396 692
rect 5443 652 5452 692
rect 5492 652 5932 692
rect 5972 652 5981 692
rect 6028 692 6068 736
rect 6787 735 6845 736
rect 6892 736 8236 776
rect 8276 736 8285 776
rect 8899 736 8908 776
rect 8948 736 15244 776
rect 15284 736 15293 776
rect 20039 736 20048 776
rect 20088 736 20130 776
rect 20170 736 20212 776
rect 20252 736 20294 776
rect 20334 736 20376 776
rect 20416 736 20425 776
rect 6892 692 6932 736
rect 15619 692 15677 693
rect 17923 692 17981 693
rect 6028 652 6932 692
rect 7747 652 7756 692
rect 7796 652 8812 692
rect 8852 652 8861 692
rect 9475 652 9484 692
rect 9524 652 12980 692
rect 14083 652 14092 692
rect 14132 652 14956 692
rect 14996 652 15005 692
rect 15534 652 15628 692
rect 15668 652 15677 692
rect 17838 652 17932 692
rect 17972 652 17981 692
rect 4675 651 4733 652
rect 5923 651 5981 652
rect 5347 608 5405 609
rect 12940 608 12980 652
rect 15619 651 15677 652
rect 17923 651 17981 652
rect 18115 692 18173 693
rect 18307 692 18365 693
rect 18499 692 18557 693
rect 19459 692 19517 693
rect 18115 652 18124 692
rect 18164 652 18258 692
rect 18307 652 18316 692
rect 18356 652 18450 692
rect 18499 652 18508 692
rect 18548 652 18642 692
rect 19374 652 19468 692
rect 19508 652 19517 692
rect 18115 651 18173 652
rect 18307 651 18365 652
rect 18499 651 18557 652
rect 19459 651 19517 652
rect 16963 608 17021 609
rect 1027 568 1036 608
rect 1076 568 3340 608
rect 3380 568 3389 608
rect 4588 568 4916 608
rect 5059 568 5068 608
rect 5108 568 5356 608
rect 5396 568 5405 608
rect 8035 568 8044 608
rect 8084 568 8332 608
rect 8372 568 8381 608
rect 9091 568 9100 608
rect 9140 568 12844 608
rect 12884 568 12893 608
rect 12940 568 15820 608
rect 15860 568 15869 608
rect 16963 568 16972 608
rect 17012 568 19276 608
rect 19316 568 19325 608
rect 1027 567 1085 568
rect 4876 524 4916 568
rect 5347 567 5405 568
rect 16963 567 17021 568
rect 9955 524 10013 525
rect 18691 524 18749 525
rect 4876 484 9964 524
rect 10004 484 10013 524
rect 10147 484 10156 524
rect 10196 484 10828 524
rect 10868 484 10877 524
rect 11011 484 11020 524
rect 11060 484 11596 524
rect 11636 484 11645 524
rect 12739 484 12748 524
rect 12788 484 13612 524
rect 13652 484 13661 524
rect 18606 484 18700 524
rect 18740 484 18749 524
rect 9955 483 10013 484
rect 18691 483 18749 484
rect 0 440 80 460
rect 7555 440 7613 441
rect 0 400 4204 440
rect 4244 400 4253 440
rect 4675 400 4684 440
rect 4724 400 7564 440
rect 7604 400 7613 440
rect 9667 400 9676 440
rect 9716 400 12460 440
rect 12500 400 12509 440
rect 13123 400 13132 440
rect 13172 400 14476 440
rect 14516 400 14525 440
rect 0 380 80 400
rect 7555 399 7613 400
rect 8515 356 8573 357
rect 14275 356 14333 357
rect 3715 316 3724 356
rect 3764 316 8524 356
rect 8564 316 8573 356
rect 10339 316 10348 356
rect 10388 316 11020 356
rect 11060 316 11069 356
rect 14190 316 14284 356
rect 14324 316 14333 356
rect 15043 316 15052 356
rect 15092 316 18220 356
rect 18260 316 18269 356
rect 8515 315 8573 316
rect 14275 315 14333 316
rect 1219 272 1277 273
rect 5251 272 5309 273
rect 11491 272 11549 273
rect 1219 232 1228 272
rect 1268 232 4876 272
rect 4916 232 4925 272
rect 5166 232 5260 272
rect 5300 232 5309 272
rect 6019 232 6028 272
rect 6068 232 11500 272
rect 11540 232 11549 272
rect 1219 231 1277 232
rect 5251 231 5309 232
rect 11491 231 11549 232
rect 2500 148 2668 188
rect 2708 148 2717 188
rect 0 104 80 124
rect 2500 104 2540 148
rect 0 64 2540 104
rect 0 44 80 64
<< via3 >>
rect 1612 42736 1652 42776
rect 11404 42652 11444 42692
rect 4780 42568 4820 42608
rect 7756 42232 7796 42272
rect 14668 42148 14708 42188
rect 8044 41728 8084 41768
rect 13612 41728 13652 41768
rect 7852 41644 7892 41684
rect 13804 41644 13844 41684
rect 15052 41644 15092 41684
rect 18700 41644 18740 41684
rect 4928 41560 4968 41600
rect 5010 41560 5050 41600
rect 5092 41560 5132 41600
rect 5174 41560 5214 41600
rect 5256 41560 5296 41600
rect 7468 41560 7508 41600
rect 9484 41560 9524 41600
rect 11212 41560 11252 41600
rect 12556 41560 12596 41600
rect 13420 41560 13460 41600
rect 13708 41560 13748 41600
rect 14092 41560 14132 41600
rect 14476 41560 14516 41600
rect 14860 41560 14900 41600
rect 16684 41560 16724 41600
rect 20048 41560 20088 41600
rect 20130 41560 20170 41600
rect 20212 41560 20252 41600
rect 20294 41560 20334 41600
rect 20376 41560 20416 41600
rect 11788 41476 11828 41516
rect 5548 41140 5588 41180
rect 13996 41224 14036 41264
rect 10252 41140 10292 41180
rect 11692 41140 11732 41180
rect 3436 41056 3476 41096
rect 4204 41056 4244 41096
rect 4780 41056 4820 41096
rect 14284 40972 14324 41012
rect 15148 40972 15188 41012
rect 3688 40804 3728 40844
rect 3770 40804 3810 40844
rect 3852 40804 3892 40844
rect 3934 40804 3974 40844
rect 4016 40804 4056 40844
rect 12364 40804 12404 40844
rect 17740 40804 17780 40844
rect 18808 40804 18848 40844
rect 18890 40804 18930 40844
rect 18972 40804 19012 40844
rect 19054 40804 19094 40844
rect 19136 40804 19176 40844
rect 2284 40636 2324 40676
rect 4780 40636 4820 40676
rect 18700 40636 18740 40676
rect 6316 40552 6356 40592
rect 13516 40552 13556 40592
rect 15820 40552 15860 40592
rect 20524 40552 20564 40592
rect 8620 40468 8660 40508
rect 18316 40468 18356 40508
rect 2956 40384 2996 40424
rect 3244 40300 3284 40340
rect 9196 40300 9236 40340
rect 16300 40300 16340 40340
rect 18124 40300 18164 40340
rect 3532 40216 3572 40256
rect 1324 40048 1364 40088
rect 4928 40048 4968 40088
rect 5010 40048 5050 40088
rect 5092 40048 5132 40088
rect 5174 40048 5214 40088
rect 5256 40048 5296 40088
rect 8716 40048 8756 40088
rect 20048 40048 20088 40088
rect 20130 40048 20170 40088
rect 20212 40048 20252 40088
rect 20294 40048 20334 40088
rect 20376 40048 20416 40088
rect 1420 39964 1460 40004
rect 7372 39964 7412 40004
rect 17548 39964 17588 40004
rect 8140 39880 8180 39920
rect 17644 39880 17684 39920
rect 5068 39628 5108 39668
rect 6796 39628 6836 39668
rect 2764 39544 2804 39584
rect 3820 39544 3860 39584
rect 2284 39376 2324 39416
rect 6604 39544 6644 39584
rect 11212 39544 11252 39584
rect 19852 39712 19892 39752
rect 20620 39712 20660 39752
rect 15724 39544 15764 39584
rect 17932 39544 17972 39584
rect 4012 39460 4052 39500
rect 4396 39460 4436 39500
rect 8908 39460 8948 39500
rect 3688 39292 3728 39332
rect 3770 39292 3810 39332
rect 3852 39292 3892 39332
rect 3934 39292 3974 39332
rect 4016 39292 4056 39332
rect 18808 39292 18848 39332
rect 18890 39292 18930 39332
rect 18972 39292 19012 39332
rect 19054 39292 19094 39332
rect 19136 39292 19176 39332
rect 76 39208 116 39248
rect 19468 39208 19508 39248
rect 2188 39124 2228 39164
rect 8236 39040 8276 39080
rect 11308 39040 11348 39080
rect 4684 38956 4724 38996
rect 4972 38956 5012 38996
rect 6700 38956 6740 38996
rect 6892 38956 6932 38996
rect 10636 38872 10676 38912
rect 10924 38872 10964 38912
rect 6220 38788 6260 38828
rect 19948 38788 19988 38828
rect 1420 38704 1460 38744
rect 17452 38704 17492 38744
rect 18508 38704 18548 38744
rect 2188 38620 2228 38660
rect 4928 38536 4968 38576
rect 5010 38536 5050 38576
rect 5092 38536 5132 38576
rect 5174 38536 5214 38576
rect 5256 38536 5296 38576
rect 19948 38536 19988 38576
rect 20048 38536 20088 38576
rect 20130 38536 20170 38576
rect 20212 38536 20252 38576
rect 20294 38536 20334 38576
rect 20376 38536 20416 38576
rect 19468 38452 19508 38492
rect 7948 38368 7988 38408
rect 17644 38368 17684 38408
rect 20428 38368 20468 38408
rect 2668 38116 2708 38156
rect 4396 38116 4436 38156
rect 3820 37948 3860 37988
rect 11596 38200 11636 38240
rect 5932 38116 5972 38156
rect 17164 38116 17204 38156
rect 17356 38116 17396 38156
rect 19852 38116 19892 38156
rect 6028 38032 6068 38072
rect 18700 38032 18740 38072
rect 20524 38032 20564 38072
rect 17356 37948 17396 37988
rect 19276 37948 19316 37988
rect 17260 37864 17300 37904
rect 2476 37780 2516 37820
rect 2668 37780 2708 37820
rect 3436 37780 3476 37820
rect 3688 37780 3728 37820
rect 3770 37780 3810 37820
rect 3852 37780 3892 37820
rect 3934 37780 3974 37820
rect 4016 37780 4056 37820
rect 13996 37780 14036 37820
rect 17548 37864 17588 37904
rect 18808 37780 18848 37820
rect 18890 37780 18930 37820
rect 18972 37780 19012 37820
rect 19054 37780 19094 37820
rect 19136 37780 19176 37820
rect 2476 37528 2516 37568
rect 4588 37528 4628 37568
rect 11788 37528 11828 37568
rect 18700 37528 18740 37568
rect 5548 37360 5588 37400
rect 10828 37276 10868 37316
rect 4780 37192 4820 37232
rect 5644 37192 5684 37232
rect 20908 37192 20948 37232
rect 5836 37108 5876 37148
rect 4928 37024 4968 37064
rect 5010 37024 5050 37064
rect 5092 37024 5132 37064
rect 5174 37024 5214 37064
rect 5256 37024 5296 37064
rect 9004 37024 9044 37064
rect 20048 37024 20088 37064
rect 20130 37024 20170 37064
rect 20212 37024 20252 37064
rect 20294 37024 20334 37064
rect 20376 37024 20416 37064
rect 10732 36940 10772 36980
rect 17836 36940 17876 36980
rect 16492 36772 16532 36812
rect 7180 36688 7220 36728
rect 17260 36688 17300 36728
rect 17740 36688 17780 36728
rect 7084 36604 7124 36644
rect 1324 36520 1364 36560
rect 1804 36520 1844 36560
rect 10444 36604 10484 36644
rect 4684 36520 4724 36560
rect 12652 36352 12692 36392
rect 3688 36268 3728 36308
rect 3770 36268 3810 36308
rect 3852 36268 3892 36308
rect 3934 36268 3974 36308
rect 4016 36268 4056 36308
rect 18808 36268 18848 36308
rect 18890 36268 18930 36308
rect 18972 36268 19012 36308
rect 19054 36268 19094 36308
rect 19136 36268 19176 36308
rect 19372 36268 19412 36308
rect 9388 36184 9428 36224
rect 17260 36184 17300 36224
rect 6316 36016 6356 36056
rect 4876 35848 4916 35888
rect 19372 35848 19412 35888
rect 4012 35680 4052 35720
rect 9580 35680 9620 35720
rect 13036 35680 13076 35720
rect 17356 35680 17396 35720
rect 4928 35512 4968 35552
rect 5010 35512 5050 35552
rect 5092 35512 5132 35552
rect 5174 35512 5214 35552
rect 5256 35512 5296 35552
rect 4108 35344 4148 35384
rect 19372 35344 19412 35384
rect 20048 35512 20088 35552
rect 20130 35512 20170 35552
rect 20212 35512 20252 35552
rect 20294 35512 20334 35552
rect 20376 35512 20416 35552
rect 20908 35512 20948 35552
rect 7468 35008 7508 35048
rect 10060 35260 10100 35300
rect 10732 35260 10772 35300
rect 8812 35176 8852 35216
rect 9100 35176 9140 35216
rect 17836 35092 17876 35132
rect 18700 35008 18740 35048
rect 8908 34924 8948 34964
rect 9676 34924 9716 34964
rect 17164 34840 17204 34880
rect 3340 34756 3380 34796
rect 3688 34756 3728 34796
rect 3770 34756 3810 34796
rect 3852 34756 3892 34796
rect 3934 34756 3974 34796
rect 4016 34756 4056 34796
rect 9868 34756 9908 34796
rect 18808 34756 18848 34796
rect 18890 34756 18930 34796
rect 18972 34756 19012 34796
rect 19054 34756 19094 34796
rect 19136 34756 19176 34796
rect 9292 34672 9332 34712
rect 9964 34588 10004 34628
rect 4492 34336 4532 34376
rect 7084 34252 7124 34292
rect 8332 34252 8372 34292
rect 9004 34252 9044 34292
rect 9772 34252 9812 34292
rect 15244 34252 15284 34292
rect 6316 34168 6356 34208
rect 8524 34168 8564 34208
rect 4928 34000 4968 34040
rect 5010 34000 5050 34040
rect 5092 34000 5132 34040
rect 5174 34000 5214 34040
rect 5256 34000 5296 34040
rect 8428 34000 8468 34040
rect 9484 34000 9524 34040
rect 12076 34000 12116 34040
rect 20048 34000 20088 34040
rect 20130 34000 20170 34040
rect 20212 34000 20252 34040
rect 20294 34000 20334 34040
rect 20376 34000 20416 34040
rect 11980 33832 12020 33872
rect 1612 33748 1652 33788
rect 8428 33664 8468 33704
rect 19564 33664 19604 33704
rect 7756 33580 7796 33620
rect 7948 33580 7988 33620
rect 9676 33580 9716 33620
rect 7276 33496 7316 33536
rect 1708 33328 1748 33368
rect 12268 33328 12308 33368
rect 3688 33244 3728 33284
rect 3770 33244 3810 33284
rect 3852 33244 3892 33284
rect 3934 33244 3974 33284
rect 4016 33244 4056 33284
rect 18808 33244 18848 33284
rect 18890 33244 18930 33284
rect 18972 33244 19012 33284
rect 19054 33244 19094 33284
rect 19136 33244 19176 33284
rect 1900 33160 1940 33200
rect 19372 33160 19412 33200
rect 12652 32908 12692 32948
rect 9964 32824 10004 32864
rect 14956 32824 14996 32864
rect 15916 32824 15956 32864
rect 4300 32740 4340 32780
rect 4684 32740 4724 32780
rect 9292 32740 9332 32780
rect 9580 32656 9620 32696
rect 8332 32572 8372 32612
rect 4928 32488 4968 32528
rect 5010 32488 5050 32528
rect 5092 32488 5132 32528
rect 5174 32488 5214 32528
rect 5256 32488 5296 32528
rect 20048 32488 20088 32528
rect 20130 32488 20170 32528
rect 20212 32488 20252 32528
rect 20294 32488 20334 32528
rect 20376 32488 20416 32528
rect 4396 32152 4436 32192
rect 8716 32152 8756 32192
rect 14668 32152 14708 32192
rect 16588 32152 16628 32192
rect 15340 32068 15380 32108
rect 16396 32068 16436 32108
rect 3688 31732 3728 31772
rect 3770 31732 3810 31772
rect 3852 31732 3892 31772
rect 3934 31732 3974 31772
rect 4016 31732 4056 31772
rect 14380 31732 14420 31772
rect 18808 31732 18848 31772
rect 18890 31732 18930 31772
rect 18972 31732 19012 31772
rect 19054 31732 19094 31772
rect 19136 31732 19176 31772
rect 14572 31396 14612 31436
rect 17260 31396 17300 31436
rect 5452 31312 5492 31352
rect 6412 31312 6452 31352
rect 8716 31312 8756 31352
rect 12364 31312 12404 31352
rect 4492 31228 4532 31268
rect 9292 31228 9332 31268
rect 8812 31144 8852 31184
rect 12172 31144 12212 31184
rect 18220 31228 18260 31268
rect 19468 31144 19508 31184
rect 3436 31060 3476 31100
rect 4928 30976 4968 31016
rect 5010 30976 5050 31016
rect 5092 30976 5132 31016
rect 5174 30976 5214 31016
rect 5256 30976 5296 31016
rect 16492 30976 16532 31016
rect 20048 30976 20088 31016
rect 20130 30976 20170 31016
rect 20212 30976 20252 31016
rect 20294 30976 20334 31016
rect 20376 30976 20416 31016
rect 5548 30724 5588 30764
rect 9004 30640 9044 30680
rect 4108 30472 4148 30512
rect 13900 30640 13940 30680
rect 14380 30640 14420 30680
rect 19564 30640 19604 30680
rect 17548 30556 17588 30596
rect 18604 30472 18644 30512
rect 16396 30304 16436 30344
rect 3688 30220 3728 30260
rect 3770 30220 3810 30260
rect 3852 30220 3892 30260
rect 3934 30220 3974 30260
rect 4016 30220 4056 30260
rect 18808 30220 18848 30260
rect 18890 30220 18930 30260
rect 18972 30220 19012 30260
rect 19054 30220 19094 30260
rect 19136 30220 19176 30260
rect 19276 30220 19316 30260
rect 3148 30136 3188 30176
rect 3052 30052 3092 30092
rect 13996 30052 14036 30092
rect 1324 29800 1364 29840
rect 11788 29884 11828 29924
rect 12652 29800 12692 29840
rect 19564 29800 19604 29840
rect 16972 29632 17012 29672
rect 3052 29548 3092 29588
rect 4928 29464 4968 29504
rect 5010 29464 5050 29504
rect 5092 29464 5132 29504
rect 5174 29464 5214 29504
rect 5256 29464 5296 29504
rect 6508 29464 6548 29504
rect 20048 29464 20088 29504
rect 20130 29464 20170 29504
rect 20212 29464 20252 29504
rect 20294 29464 20334 29504
rect 20376 29464 20416 29504
rect 12268 29380 12308 29420
rect 11980 29296 12020 29336
rect 5452 29212 5492 29252
rect 6508 29212 6548 29252
rect 18412 29296 18452 29336
rect 14188 29212 14228 29252
rect 15436 29212 15476 29252
rect 4108 29128 4148 29168
rect 14956 29128 14996 29168
rect 76 28960 116 29000
rect 8524 28960 8564 29000
rect 9772 28960 9812 29000
rect 11020 28960 11060 29000
rect 11788 28960 11828 29000
rect 19852 28960 19892 29000
rect 8908 28876 8948 28916
rect 16204 28876 16244 28916
rect 13996 28792 14036 28832
rect 3688 28708 3728 28748
rect 3770 28708 3810 28748
rect 3852 28708 3892 28748
rect 3934 28708 3974 28748
rect 4016 28708 4056 28748
rect 14572 28708 14612 28748
rect 18808 28708 18848 28748
rect 18890 28708 18930 28748
rect 18972 28708 19012 28748
rect 19054 28708 19094 28748
rect 19136 28708 19176 28748
rect 17644 28624 17684 28664
rect 8140 28540 8180 28580
rect 11788 28540 11828 28580
rect 12364 28456 12404 28496
rect 17068 28456 17108 28496
rect 16972 28372 17012 28412
rect 17548 28288 17588 28328
rect 9484 28204 9524 28244
rect 12460 28120 12500 28160
rect 15916 28036 15956 28076
rect 4928 27952 4968 27992
rect 5010 27952 5050 27992
rect 5092 27952 5132 27992
rect 5174 27952 5214 27992
rect 5256 27952 5296 27992
rect 9292 27952 9332 27992
rect 20048 27952 20088 27992
rect 20130 27952 20170 27992
rect 20212 27952 20252 27992
rect 20294 27952 20334 27992
rect 20376 27952 20416 27992
rect 18220 27868 18260 27908
rect 9484 27784 9524 27824
rect 18604 27784 18644 27824
rect 2572 27700 2612 27740
rect 19468 27700 19508 27740
rect 1612 27616 1652 27656
rect 4588 27616 4628 27656
rect 4780 27616 4820 27656
rect 18412 27616 18452 27656
rect 5548 27448 5588 27488
rect 15916 27448 15956 27488
rect 8716 27364 8756 27404
rect 12364 27364 12404 27404
rect 6508 27280 6548 27320
rect 3688 27196 3728 27236
rect 3770 27196 3810 27236
rect 3852 27196 3892 27236
rect 3934 27196 3974 27236
rect 4016 27196 4056 27236
rect 11500 27196 11540 27236
rect 15532 27196 15572 27236
rect 18808 27196 18848 27236
rect 18890 27196 18930 27236
rect 18972 27196 19012 27236
rect 19054 27196 19094 27236
rect 19136 27196 19176 27236
rect 7084 27112 7124 27152
rect 3340 27028 3380 27068
rect 5740 27028 5780 27068
rect 14188 26944 14228 26984
rect 12268 26860 12308 26900
rect 15724 26860 15764 26900
rect 6508 26692 6548 26732
rect 9004 26692 9044 26732
rect 11884 26692 11924 26732
rect 15916 26692 15956 26732
rect 17644 26692 17684 26732
rect 18412 26692 18452 26732
rect 16972 26608 17012 26648
rect 2572 26440 2612 26480
rect 2860 26440 2900 26480
rect 4928 26440 4968 26480
rect 5010 26440 5050 26480
rect 5092 26440 5132 26480
rect 5174 26440 5214 26480
rect 5256 26440 5296 26480
rect 7084 26440 7124 26480
rect 9964 26356 10004 26396
rect 11500 26440 11540 26480
rect 18028 26440 18068 26480
rect 20048 26440 20088 26480
rect 20130 26440 20170 26480
rect 20212 26440 20252 26480
rect 20294 26440 20334 26480
rect 20376 26440 20416 26480
rect 12748 26356 12788 26396
rect 14380 26356 14420 26396
rect 9004 26272 9044 26312
rect 14188 26272 14228 26312
rect 16972 26272 17012 26312
rect 1324 26188 1364 26228
rect 1516 26104 1556 26144
rect 12268 26020 12308 26060
rect 16204 26020 16244 26060
rect 16780 26020 16820 26060
rect 14956 25936 14996 25976
rect 3688 25684 3728 25724
rect 3770 25684 3810 25724
rect 3852 25684 3892 25724
rect 3934 25684 3974 25724
rect 4016 25684 4056 25724
rect 5452 25684 5492 25724
rect 15532 25684 15572 25724
rect 18808 25684 18848 25724
rect 18890 25684 18930 25724
rect 18972 25684 19012 25724
rect 19054 25684 19094 25724
rect 19136 25684 19176 25724
rect 14764 25600 14804 25640
rect 4780 25516 4820 25556
rect 1804 25432 1844 25472
rect 14380 25348 14420 25388
rect 3244 25264 3284 25304
rect 13324 25264 13364 25304
rect 2380 25180 2420 25220
rect 4012 25180 4052 25220
rect 7756 25180 7796 25220
rect 10156 25180 10196 25220
rect 10348 25180 10388 25220
rect 12364 25180 12404 25220
rect 15628 25180 15668 25220
rect 16588 25180 16628 25220
rect 11788 25096 11828 25136
rect 17548 25012 17588 25052
rect 4928 24928 4968 24968
rect 5010 24928 5050 24968
rect 5092 24928 5132 24968
rect 5174 24928 5214 24968
rect 5256 24928 5296 24968
rect 20048 24928 20088 24968
rect 20130 24928 20170 24968
rect 20212 24928 20252 24968
rect 20294 24928 20334 24968
rect 20376 24928 20416 24968
rect 16396 24844 16436 24884
rect 3340 24760 3380 24800
rect 9964 24676 10004 24716
rect 5452 24592 5492 24632
rect 14572 24592 14612 24632
rect 16492 24592 16532 24632
rect 19660 24592 19700 24632
rect 2092 24508 2132 24548
rect 7180 24508 7220 24548
rect 13228 24508 13268 24548
rect 18028 24424 18068 24464
rect 11116 24340 11156 24380
rect 13516 24340 13556 24380
rect 14764 24256 14804 24296
rect 3688 24172 3728 24212
rect 3770 24172 3810 24212
rect 3852 24172 3892 24212
rect 3934 24172 3974 24212
rect 4016 24172 4056 24212
rect 12076 24172 12116 24212
rect 18028 24172 18068 24212
rect 18808 24172 18848 24212
rect 18890 24172 18930 24212
rect 18972 24172 19012 24212
rect 19054 24172 19094 24212
rect 19136 24172 19176 24212
rect 8908 24088 8948 24128
rect 17356 23920 17396 23960
rect 5836 23836 5876 23876
rect 1708 23752 1748 23792
rect 2860 23752 2900 23792
rect 16492 23752 16532 23792
rect 16780 23752 16820 23792
rect 6508 23500 6548 23540
rect 4928 23416 4968 23456
rect 5010 23416 5050 23456
rect 5092 23416 5132 23456
rect 5174 23416 5214 23456
rect 5256 23416 5296 23456
rect 7180 23416 7220 23456
rect 1708 23332 1748 23372
rect 18412 23500 18452 23540
rect 16972 23416 17012 23456
rect 18220 23416 18260 23456
rect 20048 23416 20088 23456
rect 20130 23416 20170 23456
rect 20212 23416 20252 23456
rect 20294 23416 20334 23456
rect 20376 23416 20416 23456
rect 13324 23332 13364 23372
rect 13516 23332 13556 23372
rect 7756 23248 7796 23288
rect 8428 23248 8468 23288
rect 17068 23248 17108 23288
rect 4396 23164 4436 23204
rect 4684 23080 4724 23120
rect 10348 22996 10388 23036
rect 16972 22912 17012 22952
rect 2188 22744 2228 22784
rect 6220 22744 6260 22784
rect 9100 22828 9140 22868
rect 9580 22828 9620 22868
rect 16876 22744 16916 22784
rect 2860 22660 2900 22700
rect 3340 22660 3380 22700
rect 3688 22660 3728 22700
rect 3770 22660 3810 22700
rect 3852 22660 3892 22700
rect 3934 22660 3974 22700
rect 4016 22660 4056 22700
rect 11884 22660 11924 22700
rect 12076 22660 12116 22700
rect 15244 22660 15284 22700
rect 16396 22660 16436 22700
rect 18808 22660 18848 22700
rect 18890 22660 18930 22700
rect 18972 22660 19012 22700
rect 19054 22660 19094 22700
rect 19136 22660 19176 22700
rect 2380 22576 2420 22616
rect 7180 22576 7220 22616
rect 4300 22492 4340 22532
rect 6316 22492 6356 22532
rect 11020 22492 11060 22532
rect 18220 22492 18260 22532
rect 3148 22324 3188 22364
rect 11020 22324 11060 22364
rect 13516 22324 13556 22364
rect 15532 22324 15572 22364
rect 1900 22240 1940 22280
rect 2380 22240 2420 22280
rect 6508 22240 6548 22280
rect 15916 22240 15956 22280
rect 16108 22240 16148 22280
rect 20716 22072 20756 22112
rect 2380 21988 2420 22028
rect 3244 21904 3284 21944
rect 4492 21904 4532 21944
rect 4928 21904 4968 21944
rect 5010 21904 5050 21944
rect 5092 21904 5132 21944
rect 5174 21904 5214 21944
rect 5256 21904 5296 21944
rect 20048 21904 20088 21944
rect 20130 21904 20170 21944
rect 20212 21904 20252 21944
rect 20294 21904 20334 21944
rect 20376 21904 20416 21944
rect 5740 21820 5780 21860
rect 16780 21820 16820 21860
rect 18028 21820 18068 21860
rect 7084 21736 7124 21776
rect 12076 21736 12116 21776
rect 6508 21652 6548 21692
rect 7372 21652 7412 21692
rect 12652 21652 12692 21692
rect 16108 21568 16148 21608
rect 19948 21568 19988 21608
rect 15532 21484 15572 21524
rect 9484 21400 9524 21440
rect 9676 21400 9716 21440
rect 12748 21400 12788 21440
rect 13612 21400 13652 21440
rect 19276 21400 19316 21440
rect 4492 21232 4532 21272
rect 11692 21232 11732 21272
rect 16972 21232 17012 21272
rect 3688 21148 3728 21188
rect 3770 21148 3810 21188
rect 3852 21148 3892 21188
rect 3934 21148 3974 21188
rect 4016 21148 4056 21188
rect 9676 21148 9716 21188
rect 18808 21148 18848 21188
rect 18890 21148 18930 21188
rect 18972 21148 19012 21188
rect 19054 21148 19094 21188
rect 19136 21148 19176 21188
rect 4108 20980 4148 21020
rect 6220 20980 6260 21020
rect 6316 20896 6356 20936
rect 4780 20812 4820 20852
rect 7372 20812 7412 20852
rect 6220 20728 6260 20768
rect 12748 20728 12788 20768
rect 14188 20728 14228 20768
rect 8332 20644 8372 20684
rect 16588 20644 16628 20684
rect 4928 20392 4968 20432
rect 5010 20392 5050 20432
rect 5092 20392 5132 20432
rect 5174 20392 5214 20432
rect 5256 20392 5296 20432
rect 20048 20392 20088 20432
rect 20130 20392 20170 20432
rect 20212 20392 20252 20432
rect 20294 20392 20334 20432
rect 20376 20392 20416 20432
rect 5548 20308 5588 20348
rect 11020 20140 11060 20180
rect 11404 20140 11444 20180
rect 14092 20140 14132 20180
rect 15916 20140 15956 20180
rect 2860 20056 2900 20096
rect 9772 20056 9812 20096
rect 11884 20056 11924 20096
rect 16396 20056 16436 20096
rect 19468 20056 19508 20096
rect 19948 20056 19988 20096
rect 14092 19972 14132 20012
rect 1804 19888 1844 19928
rect 6220 19804 6260 19844
rect 7084 19804 7124 19844
rect 10156 19804 10196 19844
rect 13228 19720 13268 19760
rect 16396 19720 16436 19760
rect 3688 19636 3728 19676
rect 3770 19636 3810 19676
rect 3852 19636 3892 19676
rect 3934 19636 3974 19676
rect 4016 19636 4056 19676
rect 8908 19636 8948 19676
rect 13900 19636 13940 19676
rect 16492 19636 16532 19676
rect 18808 19636 18848 19676
rect 18890 19636 18930 19676
rect 18972 19636 19012 19676
rect 19054 19636 19094 19676
rect 19136 19636 19176 19676
rect 5836 19552 5876 19592
rect 19276 19468 19316 19508
rect 4108 19384 4148 19424
rect 12268 19300 12308 19340
rect 1612 19216 1652 19256
rect 5836 19216 5876 19256
rect 14572 19216 14612 19256
rect 2860 19132 2900 19172
rect 5452 19132 5492 19172
rect 8332 19132 8372 19172
rect 11692 19132 11732 19172
rect 17356 19132 17396 19172
rect 9964 19048 10004 19088
rect 4928 18880 4968 18920
rect 5010 18880 5050 18920
rect 5092 18880 5132 18920
rect 5174 18880 5214 18920
rect 5256 18880 5296 18920
rect 6028 18880 6068 18920
rect 12076 18880 12116 18920
rect 19468 18880 19508 18920
rect 20048 18880 20088 18920
rect 20130 18880 20170 18920
rect 20212 18880 20252 18920
rect 20294 18880 20334 18920
rect 20376 18880 20416 18920
rect 9004 18712 9044 18752
rect 11500 18712 11540 18752
rect 16300 18712 16340 18752
rect 16684 18712 16724 18752
rect 16876 18712 16916 18752
rect 3436 18628 3476 18668
rect 18412 18628 18452 18668
rect 4780 18544 4820 18584
rect 16876 18544 16916 18584
rect 11500 18460 11540 18500
rect 12364 18460 12404 18500
rect 14572 18460 14612 18500
rect 4684 18376 4724 18416
rect 11692 18376 11732 18416
rect 4588 18208 4628 18248
rect 14188 18208 14228 18248
rect 1996 18124 2036 18164
rect 2380 18124 2420 18164
rect 3688 18124 3728 18164
rect 3770 18124 3810 18164
rect 3852 18124 3892 18164
rect 3934 18124 3974 18164
rect 4016 18124 4056 18164
rect 8332 18124 8372 18164
rect 18808 18124 18848 18164
rect 18890 18124 18930 18164
rect 18972 18124 19012 18164
rect 19054 18124 19094 18164
rect 19136 18124 19176 18164
rect 4588 18040 4628 18080
rect 12364 17872 12404 17912
rect 12748 17872 12788 17912
rect 19852 17872 19892 17912
rect 8812 17704 8852 17744
rect 10156 17704 10196 17744
rect 3244 17620 3284 17660
rect 3436 17620 3476 17660
rect 7468 17620 7508 17660
rect 8908 17620 8948 17660
rect 11404 17620 11444 17660
rect 16012 17452 16052 17492
rect 4928 17368 4968 17408
rect 5010 17368 5050 17408
rect 5092 17368 5132 17408
rect 5174 17368 5214 17408
rect 5256 17368 5296 17408
rect 20048 17368 20088 17408
rect 20130 17368 20170 17408
rect 20212 17368 20252 17408
rect 20294 17368 20334 17408
rect 20376 17368 20416 17408
rect 1324 17032 1364 17072
rect 10348 16948 10388 16988
rect 16108 17032 16148 17072
rect 20908 16864 20948 16904
rect 8332 16696 8372 16736
rect 3688 16612 3728 16652
rect 3770 16612 3810 16652
rect 3852 16612 3892 16652
rect 3934 16612 3974 16652
rect 4016 16612 4056 16652
rect 18808 16612 18848 16652
rect 18890 16612 18930 16652
rect 18972 16612 19012 16652
rect 19054 16612 19094 16652
rect 19136 16612 19176 16652
rect 12556 16528 12596 16568
rect 6028 16444 6068 16484
rect 11980 16360 12020 16400
rect 17356 16360 17396 16400
rect 18604 16360 18644 16400
rect 19564 16360 19604 16400
rect 20716 16360 20756 16400
rect 14188 16276 14228 16316
rect 4300 16192 4340 16232
rect 7948 16192 7988 16232
rect 7276 16108 7316 16148
rect 12076 16108 12116 16148
rect 12460 16024 12500 16064
rect 5836 15940 5876 15980
rect 17548 15940 17588 15980
rect 4928 15856 4968 15896
rect 5010 15856 5050 15896
rect 5092 15856 5132 15896
rect 5174 15856 5214 15896
rect 5256 15856 5296 15896
rect 20048 15856 20088 15896
rect 20130 15856 20170 15896
rect 20212 15856 20252 15896
rect 20294 15856 20334 15896
rect 20376 15856 20416 15896
rect 17356 15772 17396 15812
rect 5740 15520 5780 15560
rect 6028 15520 6068 15560
rect 7276 15520 7316 15560
rect 7948 15520 7988 15560
rect 19564 15436 19604 15476
rect 7084 15268 7124 15308
rect 3688 15100 3728 15140
rect 3770 15100 3810 15140
rect 3852 15100 3892 15140
rect 3934 15100 3974 15140
rect 4016 15100 4056 15140
rect 18808 15100 18848 15140
rect 18890 15100 18930 15140
rect 18972 15100 19012 15140
rect 19054 15100 19094 15140
rect 19136 15100 19176 15140
rect 12748 14932 12788 14972
rect 8428 14764 8468 14804
rect 3244 14680 3284 14720
rect 16108 14680 16148 14720
rect 19372 14680 19412 14720
rect 11980 14596 12020 14636
rect 5836 14428 5876 14468
rect 9580 14428 9620 14468
rect 4928 14344 4968 14384
rect 5010 14344 5050 14384
rect 5092 14344 5132 14384
rect 5174 14344 5214 14384
rect 5256 14344 5296 14384
rect 6508 14344 6548 14384
rect 8428 14344 8468 14384
rect 10924 14344 10964 14384
rect 20048 14344 20088 14384
rect 20130 14344 20170 14384
rect 20212 14344 20252 14384
rect 20294 14344 20334 14384
rect 20376 14344 20416 14384
rect 4396 14260 4436 14300
rect 12364 14176 12404 14216
rect 3052 14092 3092 14132
rect 8332 14008 8372 14048
rect 10156 14008 10196 14048
rect 13324 13924 13364 13964
rect 17548 13924 17588 13964
rect 20716 13840 20756 13880
rect 6700 13756 6740 13796
rect 3688 13588 3728 13628
rect 3770 13588 3810 13628
rect 3852 13588 3892 13628
rect 3934 13588 3974 13628
rect 4016 13588 4056 13628
rect 10156 13588 10196 13628
rect 18808 13588 18848 13628
rect 18890 13588 18930 13628
rect 18972 13588 19012 13628
rect 19054 13588 19094 13628
rect 19136 13588 19176 13628
rect 6124 13168 6164 13208
rect 4204 13084 4244 13124
rect 6508 12916 6548 12956
rect 4928 12832 4968 12872
rect 5010 12832 5050 12872
rect 5092 12832 5132 12872
rect 5174 12832 5214 12872
rect 5256 12832 5296 12872
rect 20048 12832 20088 12872
rect 20130 12832 20170 12872
rect 20212 12832 20252 12872
rect 20294 12832 20334 12872
rect 20376 12832 20416 12872
rect 11980 12748 12020 12788
rect 3148 12580 3188 12620
rect 3052 12496 3092 12536
rect 8716 12496 8756 12536
rect 14380 12496 14420 12536
rect 21004 12328 21044 12368
rect 7468 12160 7508 12200
rect 3688 12076 3728 12116
rect 3770 12076 3810 12116
rect 3852 12076 3892 12116
rect 3934 12076 3974 12116
rect 4016 12076 4056 12116
rect 13324 12076 13364 12116
rect 14380 12076 14420 12116
rect 18808 12076 18848 12116
rect 18890 12076 18930 12116
rect 18972 12076 19012 12116
rect 19054 12076 19094 12116
rect 19136 12076 19176 12116
rect 76 11824 116 11864
rect 10156 11824 10196 11864
rect 10348 11824 10388 11864
rect 19276 11656 19316 11696
rect 9964 11572 10004 11612
rect 9484 11404 9524 11444
rect 4928 11320 4968 11360
rect 5010 11320 5050 11360
rect 5092 11320 5132 11360
rect 5174 11320 5214 11360
rect 5256 11320 5296 11360
rect 8812 11320 8852 11360
rect 20048 11320 20088 11360
rect 20130 11320 20170 11360
rect 20212 11320 20252 11360
rect 20294 11320 20334 11360
rect 20376 11320 20416 11360
rect 6124 11152 6164 11192
rect 9580 11152 9620 11192
rect 7468 11068 7508 11108
rect 3052 10984 3092 11024
rect 8716 10900 8756 10940
rect 4492 10648 4532 10688
rect 3688 10564 3728 10604
rect 3770 10564 3810 10604
rect 3852 10564 3892 10604
rect 3934 10564 3974 10604
rect 4016 10564 4056 10604
rect 8812 10564 8852 10604
rect 18808 10564 18848 10604
rect 18890 10564 18930 10604
rect 18972 10564 19012 10604
rect 19054 10564 19094 10604
rect 19136 10564 19176 10604
rect 14188 10396 14228 10436
rect 7084 10228 7124 10268
rect 12940 10228 12980 10268
rect 14380 10228 14420 10268
rect 7468 10144 7508 10184
rect 8908 10144 8948 10184
rect 20716 10060 20756 10100
rect 4928 9808 4968 9848
rect 5010 9808 5050 9848
rect 5092 9808 5132 9848
rect 5174 9808 5214 9848
rect 5256 9808 5296 9848
rect 9580 9808 9620 9848
rect 20048 9808 20088 9848
rect 20130 9808 20170 9848
rect 20212 9808 20252 9848
rect 20294 9808 20334 9848
rect 20376 9808 20416 9848
rect 6220 9556 6260 9596
rect 3052 9472 3092 9512
rect 3244 9304 3284 9344
rect 9388 9304 9428 9344
rect 21004 9136 21044 9176
rect 3688 9052 3728 9092
rect 3770 9052 3810 9092
rect 3852 9052 3892 9092
rect 3934 9052 3974 9092
rect 4016 9052 4056 9092
rect 8524 9052 8564 9092
rect 15820 9052 15860 9092
rect 16012 9052 16052 9092
rect 18808 9052 18848 9092
rect 18890 9052 18930 9092
rect 18972 9052 19012 9092
rect 19054 9052 19094 9092
rect 19136 9052 19176 9092
rect 16684 8968 16724 9008
rect 18412 8968 18452 9008
rect 11980 8800 12020 8840
rect 16108 8800 16148 8840
rect 17548 8800 17588 8840
rect 19468 8800 19508 8840
rect 6220 8716 6260 8756
rect 11692 8716 11732 8756
rect 16780 8716 16820 8756
rect 16684 8548 16724 8588
rect 18220 8464 18260 8504
rect 18412 8464 18452 8504
rect 19276 8380 19316 8420
rect 4928 8296 4968 8336
rect 5010 8296 5050 8336
rect 5092 8296 5132 8336
rect 5174 8296 5214 8336
rect 5256 8296 5296 8336
rect 20048 8296 20088 8336
rect 20130 8296 20170 8336
rect 20212 8296 20252 8336
rect 20294 8296 20334 8336
rect 20376 8296 20416 8336
rect 4204 8128 4244 8168
rect 4684 8128 4724 8168
rect 18412 7960 18452 8000
rect 19276 7960 19316 8000
rect 15244 7876 15284 7916
rect 12268 7708 12308 7748
rect 11500 7624 11540 7664
rect 3688 7540 3728 7580
rect 3770 7540 3810 7580
rect 3852 7540 3892 7580
rect 3934 7540 3974 7580
rect 4016 7540 4056 7580
rect 11884 7540 11924 7580
rect 18808 7540 18848 7580
rect 18890 7540 18930 7580
rect 18972 7540 19012 7580
rect 19054 7540 19094 7580
rect 19136 7540 19176 7580
rect 18220 7288 18260 7328
rect 19276 7288 19316 7328
rect 19564 7288 19604 7328
rect 4396 7204 4436 7244
rect 4396 7036 4436 7076
rect 12268 7036 12308 7076
rect 10252 6868 10292 6908
rect 4928 6784 4968 6824
rect 5010 6784 5050 6824
rect 5092 6784 5132 6824
rect 5174 6784 5214 6824
rect 5256 6784 5296 6824
rect 20048 6784 20088 6824
rect 20130 6784 20170 6824
rect 20212 6784 20252 6824
rect 20294 6784 20334 6824
rect 20376 6784 20416 6824
rect 17068 6448 17108 6488
rect 19948 6280 19988 6320
rect 12076 6196 12116 6236
rect 3688 6028 3728 6068
rect 3770 6028 3810 6068
rect 3852 6028 3892 6068
rect 3934 6028 3974 6068
rect 4016 6028 4056 6068
rect 18808 6028 18848 6068
rect 18890 6028 18930 6068
rect 18972 6028 19012 6068
rect 19054 6028 19094 6068
rect 19136 6028 19176 6068
rect 12940 5944 12980 5984
rect 18220 5692 18260 5732
rect 10156 5608 10196 5648
rect 12940 5608 12980 5648
rect 12940 5440 12980 5480
rect 15244 5440 15284 5480
rect 17068 5440 17108 5480
rect 4928 5272 4968 5312
rect 5010 5272 5050 5312
rect 5092 5272 5132 5312
rect 5174 5272 5214 5312
rect 5256 5272 5296 5312
rect 20048 5272 20088 5312
rect 20130 5272 20170 5312
rect 20212 5272 20252 5312
rect 20294 5272 20334 5312
rect 20376 5272 20416 5312
rect 2476 5188 2516 5228
rect 4492 5020 4532 5060
rect 12076 5020 12116 5060
rect 76 4936 116 4976
rect 4300 4852 4340 4892
rect 2476 4768 2516 4808
rect 14956 4768 14996 4808
rect 18412 4684 18452 4724
rect 3688 4516 3728 4556
rect 3770 4516 3810 4556
rect 3852 4516 3892 4556
rect 3934 4516 3974 4556
rect 4016 4516 4056 4556
rect 18808 4516 18848 4556
rect 18890 4516 18930 4556
rect 18972 4516 19012 4556
rect 19054 4516 19094 4556
rect 19136 4516 19176 4556
rect 4108 4348 4148 4388
rect 2860 4096 2900 4136
rect 19660 4012 19700 4052
rect 4300 3928 4340 3968
rect 18412 3844 18452 3884
rect 2860 3760 2900 3800
rect 4928 3760 4968 3800
rect 5010 3760 5050 3800
rect 5092 3760 5132 3800
rect 5174 3760 5214 3800
rect 5256 3760 5296 3800
rect 20048 3760 20088 3800
rect 20130 3760 20170 3800
rect 20212 3760 20252 3800
rect 20294 3760 20334 3800
rect 20376 3760 20416 3800
rect 12940 3676 12980 3716
rect 19276 3424 19316 3464
rect 15436 3340 15476 3380
rect 14956 3256 14996 3296
rect 3688 3004 3728 3044
rect 3770 3004 3810 3044
rect 3852 3004 3892 3044
rect 3934 3004 3974 3044
rect 4016 3004 4056 3044
rect 18808 3004 18848 3044
rect 18890 3004 18930 3044
rect 18972 3004 19012 3044
rect 19054 3004 19094 3044
rect 19136 3004 19176 3044
rect 7660 2836 7700 2876
rect 8044 2836 8084 2876
rect 9772 2668 9812 2708
rect 11404 2668 11444 2708
rect 13708 2668 13748 2708
rect 4108 2584 4148 2624
rect 8236 2584 8276 2624
rect 12172 2584 12212 2624
rect 13996 2668 14036 2708
rect 14476 2668 14516 2708
rect 14860 2668 14900 2708
rect 16108 2668 16148 2708
rect 4928 2248 4968 2288
rect 5010 2248 5050 2288
rect 5092 2248 5132 2288
rect 5174 2248 5214 2288
rect 5256 2248 5296 2288
rect 16780 2248 16820 2288
rect 20048 2248 20088 2288
rect 20130 2248 20170 2288
rect 20212 2248 20252 2288
rect 20294 2248 20334 2288
rect 20376 2248 20416 2288
rect 6892 2164 6932 2204
rect 2380 1996 2420 2036
rect 9196 1912 9236 1952
rect 9964 1912 10004 1952
rect 15340 1912 15380 1952
rect 16780 1912 16820 1952
rect 10060 1828 10100 1868
rect 10444 1828 10484 1868
rect 11308 1828 11348 1868
rect 11596 1828 11636 1868
rect 15052 1828 15092 1868
rect 17068 1744 17108 1784
rect 4684 1576 4724 1616
rect 3688 1492 3728 1532
rect 3770 1492 3810 1532
rect 3852 1492 3892 1532
rect 3934 1492 3974 1532
rect 4016 1492 4056 1532
rect 18808 1492 18848 1532
rect 18890 1492 18930 1532
rect 18972 1492 19012 1532
rect 19054 1492 19094 1532
rect 19136 1492 19176 1532
rect 8524 1324 8564 1364
rect 20620 1324 20660 1364
rect 2764 1240 2804 1280
rect 2956 1240 2996 1280
rect 3148 1240 3188 1280
rect 3532 1240 3572 1280
rect 6412 1240 6452 1280
rect 6988 1240 7028 1280
rect 7852 1240 7892 1280
rect 2284 1156 2324 1196
rect 6700 1156 6740 1196
rect 8620 1156 8660 1196
rect 10828 1156 10868 1196
rect 11212 1156 11252 1196
rect 12652 1156 12692 1196
rect 13036 1156 13076 1196
rect 13420 1156 13460 1196
rect 13804 1156 13844 1196
rect 17260 1156 17300 1196
rect 20524 1156 20564 1196
rect 1132 1072 1172 1112
rect 6604 904 6644 944
rect 17548 904 17588 944
rect 15148 820 15188 860
rect 17452 820 17492 860
rect 4928 736 4968 776
rect 5010 736 5050 776
rect 5092 736 5132 776
rect 5174 736 5214 776
rect 5256 736 5296 776
rect 6796 736 6836 776
rect 4684 652 4724 692
rect 5932 652 5972 692
rect 20048 736 20088 776
rect 20130 736 20170 776
rect 20212 736 20252 776
rect 20294 736 20334 776
rect 20376 736 20416 776
rect 15628 652 15668 692
rect 17932 652 17972 692
rect 18124 652 18164 692
rect 18316 652 18356 692
rect 18508 652 18548 692
rect 19468 652 19508 692
rect 1036 568 1076 608
rect 5356 568 5396 608
rect 16972 568 17012 608
rect 9964 484 10004 524
rect 18700 484 18740 524
rect 7564 400 7604 440
rect 8524 316 8564 356
rect 14284 316 14324 356
rect 1228 232 1268 272
rect 5260 232 5300 272
rect 11500 232 11540 272
<< metal4 >>
rect 1612 42776 1652 42785
rect 1324 40088 1364 40097
rect 76 39248 116 39257
rect 76 29000 116 39208
rect 1227 36560 1269 36569
rect 1227 36520 1228 36560
rect 1268 36520 1269 36560
rect 1227 36511 1269 36520
rect 1324 36560 1364 40048
rect 1324 36511 1364 36520
rect 1420 40004 1460 40013
rect 1420 38744 1460 39964
rect 1131 35888 1173 35897
rect 1131 35848 1132 35888
rect 1172 35848 1173 35888
rect 1131 35839 1173 35848
rect 1035 33872 1077 33881
rect 1035 33832 1036 33872
rect 1076 33832 1077 33872
rect 1035 33823 1077 33832
rect 76 28951 116 28960
rect 76 11864 116 11873
rect 76 4976 116 11824
rect 76 4927 116 4936
rect 1036 608 1076 33823
rect 1132 1112 1172 35839
rect 1132 1063 1172 1072
rect 1036 559 1076 568
rect 1228 272 1268 36511
rect 1420 31520 1460 38704
rect 1324 31480 1460 31520
rect 1612 33788 1652 42736
rect 11404 42692 11444 42701
rect 4780 42608 4820 42617
rect 3436 41096 3476 41105
rect 2284 40676 2324 40685
rect 2284 39416 2324 40636
rect 2956 40424 2996 40433
rect 2284 39367 2324 39376
rect 2764 39584 2804 39593
rect 2188 39164 2228 39173
rect 2188 38660 2228 39124
rect 1324 29840 1364 31480
rect 1324 26228 1364 29800
rect 1515 28832 1557 28841
rect 1515 28792 1516 28832
rect 1556 28792 1557 28832
rect 1515 28783 1557 28792
rect 1324 17072 1364 26188
rect 1516 26144 1556 28783
rect 1612 27656 1652 33748
rect 1804 36560 1844 36569
rect 1612 27607 1652 27616
rect 1708 33368 1748 33377
rect 1516 26095 1556 26104
rect 1708 23792 1748 33328
rect 1804 28841 1844 36520
rect 1900 33200 1940 33209
rect 1803 28832 1845 28841
rect 1803 28792 1804 28832
rect 1844 28792 1845 28832
rect 1803 28783 1845 28792
rect 1708 23372 1748 23752
rect 1708 23323 1748 23332
rect 1804 25472 1844 25481
rect 1804 19928 1844 25432
rect 1900 22280 1940 33160
rect 2188 29000 2228 38620
rect 2668 38156 2708 38165
rect 2476 37820 2516 37829
rect 2476 37568 2516 37780
rect 2668 37820 2708 38116
rect 2668 37771 2708 37780
rect 2476 37519 2516 37528
rect 2764 35729 2804 39544
rect 2956 38417 2996 40384
rect 3243 40340 3285 40349
rect 3243 40300 3244 40340
rect 3284 40300 3285 40340
rect 3243 40291 3285 40300
rect 3244 40206 3284 40291
rect 2955 38408 2997 38417
rect 2955 38368 2956 38408
rect 2996 38368 2997 38408
rect 2955 38359 2997 38368
rect 2763 35720 2805 35729
rect 2763 35680 2764 35720
rect 2804 35680 2805 35720
rect 2763 35671 2805 35680
rect 1900 22231 1940 22240
rect 1996 28960 2228 29000
rect 1804 19879 1844 19888
rect 1611 19256 1653 19265
rect 1611 19216 1612 19256
rect 1652 19216 1653 19256
rect 1611 19207 1653 19216
rect 1612 19122 1652 19207
rect 1996 18164 2036 28960
rect 2572 27740 2612 27749
rect 2572 26480 2612 27700
rect 2572 26431 2612 26440
rect 2380 25220 2420 25229
rect 1996 18115 2036 18124
rect 2092 24548 2132 24557
rect 1324 17023 1364 17032
rect 2092 15140 2132 24508
rect 2188 22784 2228 22793
rect 2188 17408 2228 22744
rect 2380 22616 2420 25180
rect 2475 25220 2517 25229
rect 2475 25180 2476 25220
rect 2516 25180 2517 25220
rect 2475 25171 2517 25180
rect 2380 22567 2420 22576
rect 2380 22280 2420 22289
rect 2380 22028 2420 22240
rect 2380 21979 2420 21988
rect 2380 18164 2420 18173
rect 2380 17753 2420 18124
rect 2379 17744 2421 17753
rect 2379 17704 2380 17744
rect 2420 17704 2421 17744
rect 2379 17695 2421 17704
rect 2188 17368 2420 17408
rect 2380 15140 2420 17368
rect 2092 15100 2228 15140
rect 2188 1289 2228 15100
rect 2284 15100 2420 15140
rect 2187 1280 2229 1289
rect 2187 1240 2188 1280
rect 2228 1240 2229 1280
rect 2187 1231 2229 1240
rect 2284 1196 2324 15100
rect 2476 6320 2516 25171
rect 2380 6280 2516 6320
rect 2380 2036 2420 6280
rect 2476 5228 2516 5237
rect 2476 4808 2516 5188
rect 2476 4759 2516 4768
rect 2380 1987 2420 1996
rect 2764 1280 2804 35671
rect 2860 26480 2900 26489
rect 2860 23792 2900 26440
rect 2860 23743 2900 23752
rect 2860 22700 2900 22709
rect 2860 20096 2900 22660
rect 2860 19172 2900 20056
rect 2860 19123 2900 19132
rect 2860 4136 2900 4145
rect 2860 3800 2900 4096
rect 2860 3751 2900 3760
rect 2764 1231 2804 1240
rect 2956 1280 2996 38359
rect 3436 37820 3476 41056
rect 4204 41096 4244 41105
rect 3688 40844 4056 40853
rect 3728 40804 3770 40844
rect 3810 40804 3852 40844
rect 3892 40804 3934 40844
rect 3974 40804 4016 40844
rect 3688 40795 4056 40804
rect 3532 40256 3572 40265
rect 3532 39677 3572 40216
rect 3531 39668 3573 39677
rect 3531 39628 3532 39668
rect 3572 39628 3573 39668
rect 3531 39619 3573 39628
rect 3436 37771 3476 37780
rect 3340 34796 3380 34805
rect 3148 30176 3188 30185
rect 3052 30092 3092 30101
rect 3052 29588 3092 30052
rect 3052 14132 3092 29548
rect 3052 12536 3092 14092
rect 3148 22364 3188 30136
rect 3340 27068 3380 34756
rect 3340 27019 3380 27028
rect 3436 31100 3476 31109
rect 3148 12620 3188 22324
rect 3244 25304 3284 25313
rect 3244 21944 3284 25264
rect 3340 24800 3380 24809
rect 3340 22700 3380 24760
rect 3340 22651 3380 22660
rect 3244 21895 3284 21904
rect 3436 19265 3476 31060
rect 3435 19256 3477 19265
rect 3435 19216 3436 19256
rect 3476 19216 3477 19256
rect 3435 19207 3477 19216
rect 3436 18668 3476 18677
rect 3148 12571 3188 12580
rect 3244 17660 3284 17669
rect 3244 14720 3284 17620
rect 3436 17660 3476 18628
rect 3436 17611 3476 17620
rect 3052 12487 3092 12496
rect 3052 11024 3092 11033
rect 3052 9512 3092 10984
rect 3052 9463 3092 9472
rect 3244 9344 3284 14680
rect 3244 9295 3284 9304
rect 2956 1231 2996 1240
rect 3147 1280 3189 1289
rect 3147 1240 3148 1280
rect 3188 1240 3189 1280
rect 3147 1231 3189 1240
rect 3532 1280 3572 39619
rect 3820 39584 3860 39593
rect 3820 39500 3860 39544
rect 4012 39500 4052 39509
rect 3820 39460 4012 39500
rect 4012 39451 4052 39460
rect 3688 39332 4056 39341
rect 3728 39292 3770 39332
rect 3810 39292 3852 39332
rect 3892 39292 3934 39332
rect 3974 39292 4016 39332
rect 3688 39283 4056 39292
rect 3820 37997 3860 38082
rect 3819 37988 3861 37997
rect 3819 37948 3820 37988
rect 3860 37948 3861 37988
rect 3819 37939 3861 37948
rect 3688 37820 4056 37829
rect 3728 37780 3770 37820
rect 3810 37780 3852 37820
rect 3892 37780 3934 37820
rect 3974 37780 4016 37820
rect 4204 37820 4244 41056
rect 4780 41096 4820 42568
rect 7756 42272 7796 42281
rect 4928 41600 5296 41609
rect 4968 41560 5010 41600
rect 5050 41560 5092 41600
rect 5132 41560 5174 41600
rect 5214 41560 5256 41600
rect 4928 41551 5296 41560
rect 7468 41600 7508 41609
rect 4780 41047 4820 41056
rect 5548 41180 5588 41189
rect 4780 40676 4820 40685
rect 4396 39500 4436 39509
rect 4396 38156 4436 39460
rect 4204 37780 4340 37820
rect 3688 37771 4056 37780
rect 3688 36308 4056 36317
rect 3728 36268 3770 36308
rect 3810 36268 3852 36308
rect 3892 36268 3934 36308
rect 3974 36268 4016 36308
rect 3688 36259 4056 36268
rect 4011 35720 4053 35729
rect 4011 35680 4012 35720
rect 4052 35680 4053 35720
rect 4011 35671 4053 35680
rect 4012 35586 4052 35671
rect 4108 35384 4148 35393
rect 3688 34796 4056 34805
rect 3728 34756 3770 34796
rect 3810 34756 3852 34796
rect 3892 34756 3934 34796
rect 3974 34756 4016 34796
rect 3688 34747 4056 34756
rect 3688 33284 4056 33293
rect 3728 33244 3770 33284
rect 3810 33244 3852 33284
rect 3892 33244 3934 33284
rect 3974 33244 4016 33284
rect 3688 33235 4056 33244
rect 3688 31772 4056 31781
rect 3728 31732 3770 31772
rect 3810 31732 3852 31772
rect 3892 31732 3934 31772
rect 3974 31732 4016 31772
rect 3688 31723 4056 31732
rect 4108 30512 4148 35344
rect 4300 32780 4340 37780
rect 4300 32731 4340 32740
rect 3688 30260 4056 30269
rect 3728 30220 3770 30260
rect 3810 30220 3852 30260
rect 3892 30220 3934 30260
rect 3974 30220 4016 30260
rect 3688 30211 4056 30220
rect 4108 29168 4148 30472
rect 4108 29000 4148 29128
rect 4396 32192 4436 38116
rect 4684 38996 4724 39005
rect 4587 37568 4629 37577
rect 4587 37528 4588 37568
rect 4628 37528 4629 37568
rect 4587 37519 4629 37528
rect 4588 37434 4628 37519
rect 4684 36560 4724 38956
rect 4780 37232 4820 40636
rect 4928 40088 5296 40097
rect 4968 40048 5010 40088
rect 5050 40048 5092 40088
rect 5132 40048 5174 40088
rect 5214 40048 5256 40088
rect 4928 40039 5296 40048
rect 5067 39668 5109 39677
rect 5067 39628 5068 39668
rect 5108 39628 5109 39668
rect 5067 39619 5109 39628
rect 5355 39668 5397 39677
rect 5355 39628 5356 39668
rect 5396 39628 5397 39668
rect 5355 39619 5397 39628
rect 5068 39534 5108 39619
rect 4971 38996 5013 39005
rect 4971 38956 4972 38996
rect 5012 38956 5013 38996
rect 4971 38947 5013 38956
rect 4972 38862 5012 38947
rect 4928 38576 5296 38585
rect 4968 38536 5010 38576
rect 5050 38536 5092 38576
rect 5132 38536 5174 38576
rect 5214 38536 5256 38576
rect 4928 38527 5296 38536
rect 4780 36653 4820 37192
rect 4928 37064 5296 37073
rect 4968 37024 5010 37064
rect 5050 37024 5092 37064
rect 5132 37024 5174 37064
rect 5214 37024 5256 37064
rect 4928 37015 5296 37024
rect 4779 36644 4821 36653
rect 4779 36604 4780 36644
rect 4820 36604 4821 36644
rect 4779 36595 4821 36604
rect 4684 36476 4724 36520
rect 4684 36436 4820 36476
rect 4684 36425 4724 36436
rect 4108 28960 4244 29000
rect 3688 28748 4056 28757
rect 3728 28708 3770 28748
rect 3810 28708 3852 28748
rect 3892 28708 3934 28748
rect 3974 28708 4016 28748
rect 3688 28699 4056 28708
rect 3688 27236 4056 27245
rect 3728 27196 3770 27236
rect 3810 27196 3852 27236
rect 3892 27196 3934 27236
rect 3974 27196 4016 27236
rect 3688 27187 4056 27196
rect 3688 25724 4056 25733
rect 3728 25684 3770 25724
rect 3810 25684 3852 25724
rect 3892 25684 3934 25724
rect 3974 25684 4016 25724
rect 3688 25675 4056 25684
rect 4011 25220 4053 25229
rect 4011 25180 4012 25220
rect 4052 25180 4053 25220
rect 4011 25171 4053 25180
rect 4012 25086 4052 25171
rect 3688 24212 4056 24221
rect 3728 24172 3770 24212
rect 3810 24172 3852 24212
rect 3892 24172 3934 24212
rect 3974 24172 4016 24212
rect 3688 24163 4056 24172
rect 3688 22700 4056 22709
rect 3728 22660 3770 22700
rect 3810 22660 3852 22700
rect 3892 22660 3934 22700
rect 3974 22660 4016 22700
rect 3688 22651 4056 22660
rect 3688 21188 4056 21197
rect 3728 21148 3770 21188
rect 3810 21148 3852 21188
rect 3892 21148 3934 21188
rect 3974 21148 4016 21188
rect 3688 21139 4056 21148
rect 4108 21020 4148 21029
rect 3688 19676 4056 19685
rect 3728 19636 3770 19676
rect 3810 19636 3852 19676
rect 3892 19636 3934 19676
rect 3974 19636 4016 19676
rect 3688 19627 4056 19636
rect 4108 19424 4148 20980
rect 4108 19375 4148 19384
rect 3688 18164 4056 18173
rect 3728 18124 3770 18164
rect 3810 18124 3852 18164
rect 3892 18124 3934 18164
rect 3974 18124 4016 18164
rect 3688 18115 4056 18124
rect 3688 16652 4056 16661
rect 3728 16612 3770 16652
rect 3810 16612 3852 16652
rect 3892 16612 3934 16652
rect 3974 16612 4016 16652
rect 3688 16603 4056 16612
rect 3688 15140 4056 15149
rect 3728 15100 3770 15140
rect 3810 15100 3852 15140
rect 3892 15100 3934 15140
rect 3974 15100 4016 15140
rect 3688 15091 4056 15100
rect 3688 13628 4056 13637
rect 3728 13588 3770 13628
rect 3810 13588 3852 13628
rect 3892 13588 3934 13628
rect 3974 13588 4016 13628
rect 3688 13579 4056 13588
rect 4204 13124 4244 28960
rect 4396 23204 4436 32152
rect 4492 34376 4532 34385
rect 4492 31268 4532 34336
rect 4492 31219 4532 31228
rect 4684 32780 4724 32789
rect 4396 23155 4436 23164
rect 4588 27656 4628 27665
rect 3688 12116 4056 12125
rect 3728 12076 3770 12116
rect 3810 12076 3852 12116
rect 3892 12076 3934 12116
rect 3974 12076 4016 12116
rect 3688 12067 4056 12076
rect 3688 10604 4056 10613
rect 3728 10564 3770 10604
rect 3810 10564 3852 10604
rect 3892 10564 3934 10604
rect 3974 10564 4016 10604
rect 3688 10555 4056 10564
rect 3688 9092 4056 9101
rect 3728 9052 3770 9092
rect 3810 9052 3852 9092
rect 3892 9052 3934 9092
rect 3974 9052 4016 9092
rect 3688 9043 4056 9052
rect 4204 8168 4244 13084
rect 4204 8119 4244 8128
rect 4300 22532 4340 22541
rect 4300 16232 4340 22492
rect 4492 21944 4532 21953
rect 4492 21272 4532 21904
rect 4492 18080 4532 21232
rect 4588 18248 4628 27616
rect 4684 23120 4724 32740
rect 4780 27656 4820 36436
rect 4875 35888 4917 35897
rect 4875 35848 4876 35888
rect 4916 35848 4917 35888
rect 4875 35839 4917 35848
rect 4876 35754 4916 35839
rect 4928 35552 5296 35561
rect 4968 35512 5010 35552
rect 5050 35512 5092 35552
rect 5132 35512 5174 35552
rect 5214 35512 5256 35552
rect 4928 35503 5296 35512
rect 4928 34040 5296 34049
rect 4968 34000 5010 34040
rect 5050 34000 5092 34040
rect 5132 34000 5174 34040
rect 5214 34000 5256 34040
rect 4928 33991 5296 34000
rect 4928 32528 5296 32537
rect 4968 32488 5010 32528
rect 5050 32488 5092 32528
rect 5132 32488 5174 32528
rect 5214 32488 5256 32528
rect 4928 32479 5296 32488
rect 4928 31016 5296 31025
rect 4968 30976 5010 31016
rect 5050 30976 5092 31016
rect 5132 30976 5174 31016
rect 5214 30976 5256 31016
rect 4928 30967 5296 30976
rect 4928 29504 5296 29513
rect 4968 29464 5010 29504
rect 5050 29464 5092 29504
rect 5132 29464 5174 29504
rect 5214 29464 5256 29504
rect 4928 29455 5296 29464
rect 4928 27992 5296 28001
rect 4968 27952 5010 27992
rect 5050 27952 5092 27992
rect 5132 27952 5174 27992
rect 5214 27952 5256 27992
rect 4928 27943 5296 27952
rect 4780 27607 4820 27616
rect 4928 26480 5296 26489
rect 4968 26440 5010 26480
rect 5050 26440 5092 26480
rect 5132 26440 5174 26480
rect 5214 26440 5256 26480
rect 4928 26431 5296 26440
rect 4684 18416 4724 23080
rect 4780 25556 4820 25565
rect 4780 20852 4820 25516
rect 4928 24968 5296 24977
rect 4968 24928 5010 24968
rect 5050 24928 5092 24968
rect 5132 24928 5174 24968
rect 5214 24928 5256 24968
rect 4928 24919 5296 24928
rect 4928 23456 5296 23465
rect 4968 23416 5010 23456
rect 5050 23416 5092 23456
rect 5132 23416 5174 23456
rect 5214 23416 5256 23456
rect 4928 23407 5296 23416
rect 4928 21944 5296 21953
rect 4968 21904 5010 21944
rect 5050 21904 5092 21944
rect 5132 21904 5174 21944
rect 5214 21904 5256 21944
rect 4928 21895 5296 21904
rect 4780 18584 4820 20812
rect 4928 20432 5296 20441
rect 4968 20392 5010 20432
rect 5050 20392 5092 20432
rect 5132 20392 5174 20432
rect 5214 20392 5256 20432
rect 4928 20383 5296 20392
rect 4928 18920 5296 18929
rect 4968 18880 5010 18920
rect 5050 18880 5092 18920
rect 5132 18880 5174 18920
rect 5214 18880 5256 18920
rect 4928 18871 5296 18880
rect 4780 18535 4820 18544
rect 4684 18367 4724 18376
rect 4588 18199 4628 18208
rect 4588 18080 4628 18089
rect 4492 18040 4588 18080
rect 4588 18031 4628 18040
rect 4928 17408 5296 17417
rect 4968 17368 5010 17408
rect 5050 17368 5092 17408
rect 5132 17368 5174 17408
rect 5214 17368 5256 17408
rect 4928 17359 5296 17368
rect 3688 7580 4056 7589
rect 3728 7540 3770 7580
rect 3810 7540 3852 7580
rect 3892 7540 3934 7580
rect 3974 7540 4016 7580
rect 3688 7531 4056 7540
rect 3688 6068 4056 6077
rect 3728 6028 3770 6068
rect 3810 6028 3852 6068
rect 3892 6028 3934 6068
rect 3974 6028 4016 6068
rect 3688 6019 4056 6028
rect 4300 4892 4340 16192
rect 4928 15896 5296 15905
rect 4968 15856 5010 15896
rect 5050 15856 5092 15896
rect 5132 15856 5174 15896
rect 5214 15856 5256 15896
rect 4928 15847 5296 15856
rect 4928 14384 5296 14393
rect 4968 14344 5010 14384
rect 5050 14344 5092 14384
rect 5132 14344 5174 14384
rect 5214 14344 5256 14384
rect 4928 14335 5296 14344
rect 4396 14300 4436 14309
rect 4396 7244 4436 14260
rect 4928 12872 5296 12881
rect 4968 12832 5010 12872
rect 5050 12832 5092 12872
rect 5132 12832 5174 12872
rect 5214 12832 5256 12872
rect 4928 12823 5296 12832
rect 4928 11360 5296 11369
rect 4968 11320 5010 11360
rect 5050 11320 5092 11360
rect 5132 11320 5174 11360
rect 5214 11320 5256 11360
rect 4928 11311 5296 11320
rect 4396 7195 4436 7204
rect 4492 10688 4532 10697
rect 4396 7076 4436 7085
rect 4396 6329 4436 7036
rect 4395 6320 4437 6329
rect 4395 6280 4396 6320
rect 4436 6280 4437 6320
rect 4395 6271 4437 6280
rect 4492 5060 4532 10648
rect 4928 9848 5296 9857
rect 4968 9808 5010 9848
rect 5050 9808 5092 9848
rect 5132 9808 5174 9848
rect 5214 9808 5256 9848
rect 4928 9799 5296 9808
rect 4928 8336 5296 8345
rect 4968 8296 5010 8336
rect 5050 8296 5092 8336
rect 5132 8296 5174 8336
rect 5214 8296 5256 8336
rect 4928 8287 5296 8296
rect 4492 5011 4532 5020
rect 4684 8168 4724 8177
rect 3688 4556 4056 4565
rect 3728 4516 3770 4556
rect 3810 4516 3852 4556
rect 3892 4516 3934 4556
rect 3974 4516 4016 4556
rect 3688 4507 4056 4516
rect 4108 4388 4148 4397
rect 3688 3044 4056 3053
rect 3728 3004 3770 3044
rect 3810 3004 3852 3044
rect 3892 3004 3934 3044
rect 3974 3004 4016 3044
rect 3688 2995 4056 3004
rect 4108 2624 4148 4348
rect 4300 3968 4340 4852
rect 4300 3919 4340 3928
rect 4108 2575 4148 2584
rect 4684 1616 4724 8128
rect 4928 6824 5296 6833
rect 4968 6784 5010 6824
rect 5050 6784 5092 6824
rect 5132 6784 5174 6824
rect 5214 6784 5256 6824
rect 4928 6775 5296 6784
rect 4928 5312 5296 5321
rect 4968 5272 5010 5312
rect 5050 5272 5092 5312
rect 5132 5272 5174 5312
rect 5214 5272 5256 5312
rect 4928 5263 5296 5272
rect 4928 3800 5296 3809
rect 4968 3760 5010 3800
rect 5050 3760 5092 3800
rect 5132 3760 5174 3800
rect 5214 3760 5256 3800
rect 4928 3751 5296 3760
rect 4928 2288 5296 2297
rect 4968 2248 5010 2288
rect 5050 2248 5092 2288
rect 5132 2248 5174 2288
rect 5214 2248 5256 2288
rect 4928 2239 5296 2248
rect 3688 1532 4056 1541
rect 3728 1492 3770 1532
rect 3810 1492 3852 1532
rect 3892 1492 3934 1532
rect 3974 1492 4016 1532
rect 3688 1483 4056 1492
rect 3532 1231 3572 1240
rect 2284 1147 2324 1156
rect 3148 1146 3188 1231
rect 4684 692 4724 1576
rect 4928 776 5296 785
rect 4968 736 5010 776
rect 5050 736 5092 776
rect 5132 736 5174 776
rect 5214 736 5256 776
rect 4928 727 5296 736
rect 4684 643 4724 652
rect 5356 608 5396 39619
rect 5548 37577 5588 41140
rect 6316 40592 6356 40601
rect 5739 38996 5781 39005
rect 5739 38956 5740 38996
rect 5780 38956 5781 38996
rect 5739 38947 5781 38956
rect 5547 37568 5589 37577
rect 5547 37528 5548 37568
rect 5588 37528 5589 37568
rect 5547 37519 5589 37528
rect 5548 37400 5588 37409
rect 5451 36644 5493 36653
rect 5451 36604 5452 36644
rect 5492 36604 5493 36644
rect 5451 36595 5493 36604
rect 5452 31352 5492 36595
rect 5548 36569 5588 37360
rect 5643 37232 5685 37241
rect 5643 37192 5644 37232
rect 5684 37192 5685 37232
rect 5643 37183 5685 37192
rect 5547 36560 5589 36569
rect 5547 36520 5548 36560
rect 5588 36520 5589 36560
rect 5547 36511 5589 36520
rect 5644 33881 5684 37183
rect 5643 33872 5685 33881
rect 5643 33832 5644 33872
rect 5684 33832 5685 33872
rect 5643 33823 5685 33832
rect 5740 32789 5780 38947
rect 6220 38828 6260 38837
rect 5932 38156 5972 38165
rect 5835 37148 5877 37157
rect 5835 37108 5836 37148
rect 5876 37108 5877 37148
rect 5835 37099 5877 37108
rect 5836 37014 5876 37099
rect 5739 32780 5781 32789
rect 5739 32740 5740 32780
rect 5780 32740 5781 32780
rect 5739 32731 5781 32740
rect 5452 31303 5492 31312
rect 5548 30764 5588 30773
rect 5452 29252 5492 29261
rect 5452 25724 5492 29212
rect 5548 27488 5588 30724
rect 5548 27439 5588 27448
rect 5452 25675 5492 25684
rect 5740 27068 5780 27077
rect 5452 24632 5492 24641
rect 5452 19172 5492 24592
rect 5740 21860 5780 27028
rect 5548 20348 5588 20357
rect 5548 19265 5588 20308
rect 5547 19256 5589 19265
rect 5547 19216 5548 19256
rect 5588 19216 5589 19256
rect 5547 19207 5589 19216
rect 5452 19123 5492 19132
rect 5740 15560 5780 21820
rect 5836 23876 5876 23885
rect 5836 19592 5876 23836
rect 5836 19256 5876 19552
rect 5836 19207 5876 19216
rect 5740 15511 5780 15520
rect 5836 15980 5876 15989
rect 5836 14468 5876 15940
rect 5836 14419 5876 14428
rect 5932 692 5972 38116
rect 6028 38072 6068 38081
rect 6028 18920 6068 38032
rect 6220 22784 6260 38788
rect 6220 22735 6260 22744
rect 6316 36056 6356 40552
rect 6891 40340 6933 40349
rect 6891 40300 6892 40340
rect 6932 40300 6933 40340
rect 6891 40291 6933 40300
rect 7371 40340 7413 40349
rect 7371 40300 7372 40340
rect 7412 40300 7413 40340
rect 7371 40291 7413 40300
rect 6795 39668 6837 39677
rect 6795 39628 6796 39668
rect 6836 39628 6837 39668
rect 6795 39619 6837 39628
rect 6316 34208 6356 36016
rect 6316 22532 6356 34168
rect 6604 39584 6644 39593
rect 6316 22483 6356 22492
rect 6412 31352 6452 31361
rect 6220 21020 6260 21029
rect 6220 20768 6260 20980
rect 6028 18871 6068 18880
rect 6124 20728 6220 20768
rect 6028 16484 6068 16493
rect 6028 15560 6068 16444
rect 6028 15511 6068 15520
rect 6124 13208 6164 20728
rect 6220 20719 6260 20728
rect 6316 20936 6356 20945
rect 6316 20180 6356 20896
rect 6220 20140 6356 20180
rect 6220 19844 6260 20140
rect 6220 19795 6260 19804
rect 6124 11192 6164 13168
rect 6124 11143 6164 11152
rect 6220 9596 6260 9605
rect 6220 8756 6260 9556
rect 6220 8707 6260 8716
rect 6412 1280 6452 31312
rect 6508 29504 6548 29513
rect 6508 29252 6548 29464
rect 6508 29203 6548 29212
rect 6508 27320 6548 27329
rect 6508 26732 6548 27280
rect 6508 26683 6548 26692
rect 6508 23540 6548 23549
rect 6508 22280 6548 23500
rect 6508 21692 6548 22240
rect 6508 21643 6548 21652
rect 6508 14384 6548 14393
rect 6508 12956 6548 14344
rect 6508 12907 6548 12916
rect 6604 11360 6644 39544
rect 6796 39534 6836 39619
rect 6892 39332 6932 40291
rect 7372 40004 7412 40291
rect 7372 39955 7412 39964
rect 6796 39292 6932 39332
rect 6700 38996 6740 39005
rect 6700 13796 6740 38956
rect 6700 13747 6740 13756
rect 6604 11320 6740 11360
rect 6412 1231 6452 1240
rect 6700 1196 6740 11320
rect 6700 1147 6740 1156
rect 6603 944 6645 953
rect 6603 904 6604 944
rect 6644 904 6645 944
rect 6603 895 6645 904
rect 6604 810 6644 895
rect 6796 776 6836 39292
rect 6892 38996 6932 39005
rect 6892 2204 6932 38956
rect 6987 37568 7029 37577
rect 6987 37528 6988 37568
rect 7028 37528 7029 37568
rect 6987 37519 7029 37528
rect 6892 2155 6932 2164
rect 6988 1280 7028 37519
rect 7180 36728 7220 36737
rect 7083 36644 7125 36653
rect 7083 36604 7084 36644
rect 7124 36604 7125 36644
rect 7083 36595 7125 36604
rect 7084 36510 7124 36595
rect 7084 34292 7124 34301
rect 7084 27152 7124 34252
rect 7084 26480 7124 27112
rect 7084 26431 7124 26440
rect 7180 24548 7220 36688
rect 7468 35300 7508 41560
rect 7468 35260 7604 35300
rect 7468 35048 7508 35057
rect 7180 24499 7220 24508
rect 7276 33536 7316 33545
rect 7180 23456 7220 23465
rect 7180 22616 7220 23416
rect 7180 22567 7220 22576
rect 7084 21776 7124 21785
rect 7084 19844 7124 21736
rect 7084 19795 7124 19804
rect 7276 16148 7316 33496
rect 7468 26480 7508 35008
rect 7564 29000 7604 35260
rect 7756 33620 7796 42232
rect 8044 41768 8084 41777
rect 7756 33571 7796 33580
rect 7852 41684 7892 41693
rect 7564 28960 7700 29000
rect 7468 26440 7604 26480
rect 7372 21692 7412 21701
rect 7372 20852 7412 21652
rect 7372 20803 7412 20812
rect 7276 15560 7316 16108
rect 7276 15511 7316 15520
rect 7468 17660 7508 17669
rect 7084 15308 7124 15317
rect 7084 10268 7124 15268
rect 7084 10219 7124 10228
rect 7468 12200 7508 17620
rect 7468 11108 7508 12160
rect 7468 10184 7508 11068
rect 7468 10135 7508 10144
rect 6988 1231 7028 1240
rect 6796 727 6836 736
rect 5932 643 5972 652
rect 5356 559 5396 568
rect 7564 440 7604 26440
rect 7660 2876 7700 28960
rect 7756 25220 7796 25229
rect 7756 23288 7796 25180
rect 7756 23239 7796 23248
rect 7660 2827 7700 2836
rect 7852 1280 7892 41644
rect 7947 38408 7989 38417
rect 7947 38368 7948 38408
rect 7988 38368 7989 38408
rect 7947 38359 7989 38368
rect 7948 38274 7988 38359
rect 7948 33620 7988 33629
rect 7948 16232 7988 33580
rect 7948 15560 7988 16192
rect 7948 15511 7988 15520
rect 8044 2876 8084 41728
rect 9484 41600 9524 41609
rect 8620 40508 8660 40517
rect 8140 39920 8180 39929
rect 8140 37241 8180 39880
rect 8236 39080 8276 39089
rect 8139 37232 8181 37241
rect 8139 37192 8140 37232
rect 8180 37192 8181 37232
rect 8139 37183 8181 37192
rect 8236 32696 8276 39040
rect 8140 32656 8276 32696
rect 8332 34292 8372 34301
rect 8140 28580 8180 32656
rect 8332 32612 8372 34252
rect 8524 34208 8564 34217
rect 8332 32563 8372 32572
rect 8428 34040 8468 34049
rect 8428 33704 8468 34000
rect 8428 29000 8468 33664
rect 8140 28531 8180 28540
rect 8236 28960 8468 29000
rect 8524 29000 8564 34168
rect 8044 2827 8084 2836
rect 8236 2624 8276 28960
rect 8524 28951 8564 28960
rect 8428 23288 8468 23297
rect 8332 20684 8372 20693
rect 8332 19172 8372 20644
rect 8332 18164 8372 19132
rect 8332 18115 8372 18124
rect 8332 16736 8372 16745
rect 8332 14048 8372 16696
rect 8428 14804 8468 23248
rect 8468 14764 8564 14804
rect 8428 14755 8468 14764
rect 8332 13999 8372 14008
rect 8428 14384 8468 14393
rect 8236 2575 8276 2584
rect 7852 1231 7892 1240
rect 7564 391 7604 400
rect 8428 281 8468 14344
rect 8524 9092 8564 14764
rect 8524 9043 8564 9052
rect 8524 1364 8564 1373
rect 8524 356 8564 1324
rect 8620 1196 8660 40468
rect 9196 40340 9236 40349
rect 8716 40088 8756 40097
rect 8716 32192 8756 40048
rect 8908 39500 8948 39509
rect 8811 37988 8853 37997
rect 8811 37948 8812 37988
rect 8852 37948 8853 37988
rect 8811 37939 8853 37948
rect 8812 35216 8852 37939
rect 8812 35167 8852 35176
rect 8908 34964 8948 39460
rect 8908 34915 8948 34924
rect 9004 37064 9044 37073
rect 9004 34292 9044 37024
rect 9004 34243 9044 34252
rect 9100 35216 9140 35225
rect 8716 31520 8756 32152
rect 8716 31480 8948 31520
rect 8716 31352 8756 31361
rect 8716 27404 8756 31312
rect 8716 27355 8756 27364
rect 8812 31184 8852 31193
rect 8812 17744 8852 31144
rect 8908 28916 8948 31480
rect 8908 28867 8948 28876
rect 9004 30680 9044 30689
rect 9004 26732 9044 30640
rect 9004 26683 9044 26692
rect 9004 26312 9044 26321
rect 8908 24128 8948 24137
rect 8908 19676 8948 24088
rect 8908 19627 8948 19636
rect 9004 18752 9044 26272
rect 9100 22868 9140 35176
rect 9100 22819 9140 22828
rect 9004 18703 9044 18712
rect 8812 17695 8852 17704
rect 8908 17660 8948 17669
rect 8716 12536 8756 12545
rect 8716 10940 8756 12496
rect 8716 10891 8756 10900
rect 8812 11360 8852 11369
rect 8812 10604 8852 11320
rect 8812 10555 8852 10564
rect 8908 10184 8948 17620
rect 8908 10135 8948 10144
rect 9196 1952 9236 40300
rect 9388 36224 9428 36233
rect 9292 34712 9332 34721
rect 9292 32780 9332 34672
rect 9292 32731 9332 32740
rect 9292 31268 9332 31277
rect 9292 27992 9332 31228
rect 9292 27943 9332 27952
rect 9388 9344 9428 36184
rect 9484 34040 9524 41560
rect 11212 41600 11252 41609
rect 10252 41180 10292 41189
rect 9484 33991 9524 34000
rect 9580 35720 9620 35729
rect 9580 32696 9620 35680
rect 10060 35300 10100 35309
rect 9580 32647 9620 32656
rect 9676 34964 9716 34973
rect 9676 34796 9716 34924
rect 9868 34796 9908 34805
rect 9676 34756 9868 34796
rect 9676 33620 9716 34756
rect 9868 34747 9908 34756
rect 9964 34628 10004 34637
rect 9484 28244 9524 28253
rect 9484 27824 9524 28204
rect 9484 27775 9524 27784
rect 9580 22868 9620 22877
rect 9484 21440 9524 21449
rect 9484 11444 9524 21400
rect 9580 14468 9620 22828
rect 9676 21440 9716 33580
rect 9772 34292 9812 34301
rect 9772 29000 9812 34252
rect 9964 32864 10004 34588
rect 9964 32815 10004 32824
rect 9772 28951 9812 28960
rect 9964 26396 10004 26405
rect 9964 24716 10004 26356
rect 9964 24667 10004 24676
rect 9676 21188 9716 21400
rect 9676 21139 9716 21148
rect 9580 14419 9620 14428
rect 9772 20096 9812 20105
rect 9484 11395 9524 11404
rect 9580 11192 9620 11201
rect 9580 9848 9620 11152
rect 9580 9799 9620 9808
rect 9388 9295 9428 9304
rect 9772 2708 9812 20056
rect 9964 19088 10004 19097
rect 9964 11612 10004 19048
rect 9964 11563 10004 11572
rect 9772 2659 9812 2668
rect 9196 1903 9236 1912
rect 9964 1952 10004 1961
rect 8620 1147 8660 1156
rect 9964 524 10004 1912
rect 10060 1868 10100 35260
rect 10156 25220 10196 25229
rect 10156 19844 10196 25180
rect 10156 19795 10196 19804
rect 10155 17744 10197 17753
rect 10155 17704 10156 17744
rect 10196 17704 10197 17744
rect 10155 17695 10197 17704
rect 10156 17610 10196 17695
rect 10156 14048 10196 14057
rect 10156 13628 10196 14008
rect 10156 13579 10196 13588
rect 10156 11864 10196 11873
rect 10156 5648 10196 11824
rect 10252 6908 10292 41140
rect 11212 39584 11252 41560
rect 10636 38912 10676 38921
rect 10636 37997 10676 38872
rect 10924 38912 10964 38921
rect 10635 37988 10677 37997
rect 10635 37948 10636 37988
rect 10676 37948 10677 37988
rect 10635 37939 10677 37948
rect 10828 37316 10868 37325
rect 10443 37148 10485 37157
rect 10443 37108 10444 37148
rect 10484 37108 10485 37148
rect 10443 37099 10485 37108
rect 10444 36644 10484 37099
rect 10348 25220 10388 25229
rect 10348 23036 10388 25180
rect 10348 16988 10388 22996
rect 10348 11864 10388 16948
rect 10348 11815 10388 11824
rect 10252 6859 10292 6868
rect 10156 5599 10196 5608
rect 10060 1819 10100 1828
rect 10444 1868 10484 36604
rect 10732 36980 10772 36989
rect 10732 35300 10772 36940
rect 10828 36653 10868 37276
rect 10827 36644 10869 36653
rect 10827 36604 10828 36644
rect 10868 36604 10869 36644
rect 10827 36595 10869 36604
rect 10732 35251 10772 35260
rect 10444 1819 10484 1828
rect 10828 1196 10868 36595
rect 10924 14384 10964 38872
rect 11020 29000 11060 29009
rect 11020 22532 11060 28960
rect 11020 22483 11060 22492
rect 11116 24380 11156 24389
rect 11020 22364 11060 22373
rect 11020 20180 11060 22324
rect 11020 20131 11060 20140
rect 11116 18341 11156 24340
rect 11115 18332 11157 18341
rect 11115 18292 11116 18332
rect 11156 18292 11157 18332
rect 11115 18283 11157 18292
rect 10924 14335 10964 14344
rect 10828 1147 10868 1156
rect 11212 1196 11252 39544
rect 11308 39080 11348 39089
rect 11308 1868 11348 39040
rect 11404 35300 11444 42652
rect 14668 42188 14708 42197
rect 13612 41768 13652 41777
rect 12556 41600 12596 41609
rect 11788 41516 11828 41525
rect 11692 41180 11732 41189
rect 11596 38240 11636 38249
rect 11404 35260 11540 35300
rect 11500 29000 11540 35260
rect 11404 28960 11540 29000
rect 11404 20180 11444 28960
rect 11500 27236 11540 27245
rect 11500 26480 11540 27196
rect 11500 26431 11540 26440
rect 11404 20131 11444 20140
rect 11500 18752 11540 18761
rect 11500 18500 11540 18712
rect 11500 18451 11540 18460
rect 11404 17660 11444 17669
rect 11404 2708 11444 17620
rect 11404 2659 11444 2668
rect 11500 7664 11540 7673
rect 11308 1819 11348 1828
rect 11212 1147 11252 1156
rect 9964 475 10004 484
rect 8524 307 8564 316
rect 1228 223 1268 232
rect 5259 272 5301 281
rect 5259 232 5260 272
rect 5300 232 5301 272
rect 5259 223 5301 232
rect 8427 272 8469 281
rect 8427 232 8428 272
rect 8468 232 8469 272
rect 8427 223 8469 232
rect 11500 272 11540 7624
rect 11596 1868 11636 38200
rect 11692 21272 11732 41140
rect 11788 37568 11828 41476
rect 11788 37519 11828 37528
rect 12364 40844 12404 40853
rect 12076 34040 12116 34049
rect 11980 33872 12020 33881
rect 11788 29924 11828 29933
rect 11788 29000 11828 29884
rect 11788 28951 11828 28960
rect 11980 29336 12020 33832
rect 11788 28580 11828 28589
rect 11788 25136 11828 28540
rect 11788 25087 11828 25096
rect 11884 26732 11924 26741
rect 11884 22700 11924 26692
rect 11884 22651 11924 22660
rect 11692 21223 11732 21232
rect 11884 20096 11924 20105
rect 11692 19172 11732 19181
rect 11692 18416 11732 19132
rect 11692 8756 11732 18376
rect 11692 8707 11732 8716
rect 11884 7580 11924 20056
rect 11980 16400 12020 29296
rect 12076 24212 12116 34000
rect 12268 33368 12308 33377
rect 12076 24163 12116 24172
rect 12172 31184 12212 31193
rect 12076 22700 12116 22709
rect 12076 21776 12116 22660
rect 12076 18920 12116 21736
rect 12076 18871 12116 18880
rect 11980 14636 12020 16360
rect 11980 14587 12020 14596
rect 12076 16148 12116 16157
rect 11980 12788 12020 12797
rect 11980 8840 12020 12748
rect 11980 8791 12020 8800
rect 11884 7531 11924 7540
rect 12076 6236 12116 16108
rect 12076 5060 12116 6196
rect 12076 5011 12116 5020
rect 12172 2624 12212 31144
rect 12268 29420 12308 33328
rect 12364 31352 12404 40804
rect 12364 31303 12404 31312
rect 12268 26900 12308 29380
rect 12364 28496 12404 28505
rect 12364 27404 12404 28456
rect 12364 27355 12404 27364
rect 12460 28160 12500 28169
rect 12268 26851 12308 26860
rect 12268 26060 12308 26069
rect 12268 19340 12308 26020
rect 12268 19291 12308 19300
rect 12364 25220 12404 25229
rect 12364 18500 12404 25180
rect 12364 18451 12404 18460
rect 12364 17912 12404 17921
rect 12364 14216 12404 17872
rect 12460 16064 12500 28120
rect 12556 16568 12596 41560
rect 13420 41600 13460 41609
rect 12652 36392 12692 36401
rect 12652 32948 12692 36352
rect 12652 29840 12692 32908
rect 12652 29791 12692 29800
rect 13036 35720 13076 35729
rect 12748 26396 12788 26405
rect 12556 16519 12596 16528
rect 12652 21692 12692 21701
rect 12460 16015 12500 16024
rect 12364 14167 12404 14176
rect 12268 7748 12308 7757
rect 12268 7076 12308 7708
rect 12268 7027 12308 7036
rect 12172 2575 12212 2584
rect 11596 1819 11636 1828
rect 12652 1196 12692 21652
rect 12748 21440 12788 26356
rect 12748 20768 12788 21400
rect 12748 20719 12788 20728
rect 12748 17912 12788 17921
rect 12748 14972 12788 17872
rect 12748 14923 12788 14932
rect 12940 10268 12980 10277
rect 12940 5984 12980 10228
rect 12940 5935 12980 5944
rect 12940 5648 12980 5657
rect 12940 5480 12980 5608
rect 12940 3716 12980 5440
rect 12940 3667 12980 3676
rect 12652 1147 12692 1156
rect 13036 1196 13076 35680
rect 13324 25304 13364 25313
rect 13228 24548 13268 24557
rect 13228 19760 13268 24508
rect 13324 23372 13364 25264
rect 13324 23323 13364 23332
rect 13228 19711 13268 19720
rect 13324 13964 13364 13973
rect 13324 12116 13364 13924
rect 13324 12067 13364 12076
rect 13036 1147 13076 1156
rect 13420 1196 13460 41560
rect 13516 40592 13556 40601
rect 13516 24380 13556 40552
rect 13516 24331 13556 24340
rect 13516 23372 13556 23381
rect 13516 22364 13556 23332
rect 13516 22315 13556 22324
rect 13612 21440 13652 41728
rect 13804 41684 13844 41693
rect 13612 21391 13652 21400
rect 13708 41600 13748 41609
rect 13708 2708 13748 41560
rect 13708 2659 13748 2668
rect 13420 1147 13460 1156
rect 13804 1196 13844 41644
rect 14092 41600 14132 41609
rect 13996 41264 14036 41273
rect 13996 37820 14036 41224
rect 13996 37771 14036 37780
rect 13900 30680 13940 30689
rect 13900 19676 13940 30640
rect 13996 30092 14036 30101
rect 13996 28832 14036 30052
rect 13996 28783 14036 28792
rect 14092 21692 14132 41560
rect 14476 41600 14516 41609
rect 14284 41012 14324 41021
rect 14188 29252 14228 29261
rect 14188 26984 14228 29212
rect 14188 26935 14228 26944
rect 13900 19627 13940 19636
rect 13996 21652 14132 21692
rect 14188 26312 14228 26321
rect 13996 2708 14036 21652
rect 14188 20768 14228 26272
rect 14092 20180 14132 20189
rect 14092 20012 14132 20140
rect 14092 19963 14132 19972
rect 14188 18248 14228 20728
rect 14188 18199 14228 18208
rect 14188 16316 14228 16325
rect 14188 10436 14228 16276
rect 14188 10387 14228 10396
rect 13996 2659 14036 2668
rect 13804 1147 13844 1156
rect 14284 356 14324 40972
rect 14380 31772 14420 31781
rect 14380 30680 14420 31732
rect 14380 30631 14420 30640
rect 14380 26396 14420 26405
rect 14380 25388 14420 26356
rect 14380 25339 14420 25348
rect 14380 12536 14420 12545
rect 14380 12116 14420 12496
rect 14380 10268 14420 12076
rect 14380 10219 14420 10228
rect 14476 2708 14516 41560
rect 14668 32192 14708 42148
rect 15052 41684 15092 41693
rect 14572 31436 14612 31445
rect 14572 28748 14612 31396
rect 14572 24632 14612 28708
rect 14572 24583 14612 24592
rect 14668 20180 14708 32152
rect 14860 41600 14900 41609
rect 14764 25640 14804 25649
rect 14764 24296 14804 25600
rect 14764 24247 14804 24256
rect 14572 20140 14708 20180
rect 14572 19256 14612 20140
rect 14572 18500 14612 19216
rect 14572 18451 14612 18460
rect 14476 2659 14516 2668
rect 14860 2708 14900 41560
rect 14956 32864 14996 32873
rect 14956 29168 14996 32824
rect 14956 25976 14996 29128
rect 14956 25927 14996 25936
rect 14956 4808 14996 4817
rect 14956 3296 14996 4768
rect 14956 3247 14996 3256
rect 14860 2659 14900 2668
rect 15052 1868 15092 41644
rect 18700 41684 18740 41693
rect 16684 41600 16724 41609
rect 15052 1819 15092 1828
rect 15148 41012 15188 41021
rect 15148 860 15188 40972
rect 15820 40592 15860 40601
rect 15724 39584 15764 39593
rect 15244 34292 15284 34301
rect 15244 22700 15284 34252
rect 15244 22651 15284 22660
rect 15340 32108 15380 32117
rect 15244 7916 15284 7925
rect 15244 5480 15284 7876
rect 15244 5431 15284 5440
rect 15340 1952 15380 32068
rect 15436 29252 15476 29261
rect 15436 3380 15476 29212
rect 15532 27236 15572 27245
rect 15532 25724 15572 27196
rect 15724 26900 15764 39544
rect 15724 26851 15764 26860
rect 15532 25675 15572 25684
rect 15628 25220 15668 25229
rect 15532 22364 15572 22373
rect 15532 21524 15572 22324
rect 15532 21475 15572 21484
rect 15436 3331 15476 3340
rect 15340 1903 15380 1912
rect 15148 811 15188 820
rect 15628 692 15668 25180
rect 15820 9092 15860 40552
rect 16300 40340 16340 40349
rect 15916 32864 15956 32873
rect 15916 28076 15956 32824
rect 15916 28027 15956 28036
rect 16204 28916 16244 28925
rect 15916 27488 15956 27497
rect 15916 26732 15956 27448
rect 15916 26683 15956 26692
rect 16204 26060 16244 28876
rect 16204 26011 16244 26020
rect 15916 22280 15956 22289
rect 15916 20180 15956 22240
rect 16108 22280 16148 22289
rect 16108 21608 16148 22240
rect 16108 21559 16148 21568
rect 15916 20131 15956 20140
rect 16300 18752 16340 40300
rect 16492 36812 16532 36821
rect 16396 32108 16436 32117
rect 16396 30344 16436 32068
rect 16396 30295 16436 30304
rect 16492 31016 16532 36772
rect 16396 24884 16436 24893
rect 16396 22700 16436 24844
rect 16492 24632 16532 30976
rect 16588 32192 16628 32201
rect 16588 25220 16628 32152
rect 16588 25171 16628 25180
rect 16532 24592 16628 24632
rect 16492 24583 16532 24592
rect 16396 22651 16436 22660
rect 16492 23792 16532 23801
rect 16396 20096 16436 20105
rect 16396 19760 16436 20056
rect 16396 19711 16436 19720
rect 16492 19676 16532 23752
rect 16588 20684 16628 24592
rect 16588 20635 16628 20644
rect 16492 19627 16532 19636
rect 16300 18703 16340 18712
rect 16684 18752 16724 41560
rect 17740 40844 17780 40853
rect 17548 40004 17588 40013
rect 17452 38744 17492 38753
rect 17164 38156 17204 38165
rect 17356 38156 17396 38165
rect 17164 34880 17204 38116
rect 17260 38116 17356 38156
rect 17260 37904 17300 38116
rect 17356 38107 17396 38116
rect 17260 37855 17300 37864
rect 17356 37988 17396 37997
rect 17260 36728 17300 36737
rect 17260 36224 17300 36688
rect 17260 36175 17300 36184
rect 17356 35720 17396 37948
rect 17356 35671 17396 35680
rect 17164 34831 17204 34840
rect 17260 31436 17300 31445
rect 16972 29672 17012 29681
rect 16972 28412 17012 29632
rect 16972 26648 17012 28372
rect 16972 26599 17012 26608
rect 17068 28496 17108 28505
rect 16972 26312 17012 26321
rect 16780 26060 16820 26069
rect 16780 23792 16820 26020
rect 16780 23743 16820 23752
rect 16972 23456 17012 26272
rect 16972 22952 17012 23416
rect 17068 23288 17108 28456
rect 17068 23239 17108 23248
rect 16972 22903 17012 22912
rect 16876 22784 16916 22793
rect 16684 18703 16724 18712
rect 16780 21860 16820 21869
rect 15820 9043 15860 9052
rect 16012 17492 16052 17501
rect 16012 9092 16052 17452
rect 16108 17072 16148 17081
rect 16108 14720 16148 17032
rect 16108 14671 16148 14680
rect 16012 9043 16052 9052
rect 16684 9008 16724 9017
rect 16108 8840 16148 8849
rect 16108 2708 16148 8800
rect 16684 8588 16724 8968
rect 16684 8539 16724 8548
rect 16780 8756 16820 21820
rect 16876 18752 16916 22744
rect 16876 18584 16916 18712
rect 16876 18535 16916 18544
rect 16972 21272 17012 21281
rect 16108 2659 16148 2668
rect 16780 2288 16820 8716
rect 16780 1952 16820 2248
rect 16780 1903 16820 1912
rect 15628 643 15668 652
rect 16972 608 17012 21232
rect 17068 6488 17108 6497
rect 17068 5480 17108 6448
rect 17068 1784 17108 5440
rect 17068 1735 17108 1744
rect 17260 1196 17300 31396
rect 17356 23960 17396 23969
rect 17356 19172 17396 23920
rect 17356 19123 17396 19132
rect 17356 16400 17396 16409
rect 17356 15812 17396 16360
rect 17356 15763 17396 15772
rect 17260 1147 17300 1156
rect 17452 860 17492 38704
rect 17548 37904 17588 39964
rect 17644 39920 17684 39929
rect 17644 38408 17684 39880
rect 17644 38359 17684 38368
rect 17548 37855 17588 37864
rect 17740 36728 17780 40804
rect 18700 40676 18740 41644
rect 20048 41600 20416 41609
rect 20088 41560 20130 41600
rect 20170 41560 20212 41600
rect 20252 41560 20294 41600
rect 20334 41560 20376 41600
rect 20048 41551 20416 41560
rect 18808 40844 19176 40853
rect 18848 40804 18890 40844
rect 18930 40804 18972 40844
rect 19012 40804 19054 40844
rect 19094 40804 19136 40844
rect 18808 40795 19176 40804
rect 18700 40627 18740 40636
rect 20524 40592 20564 40601
rect 18316 40508 18356 40517
rect 18124 40340 18164 40349
rect 17932 39584 17972 39593
rect 17740 36679 17780 36688
rect 17836 36980 17876 36989
rect 17836 35132 17876 36940
rect 17836 35083 17876 35092
rect 17548 30596 17588 30605
rect 17548 28328 17588 30556
rect 17548 25052 17588 28288
rect 17644 28664 17684 28673
rect 17644 26732 17684 28624
rect 17644 26683 17684 26692
rect 17548 25003 17588 25012
rect 17548 15980 17588 15989
rect 17548 13964 17588 15940
rect 17548 13915 17588 13924
rect 17548 8840 17588 8849
rect 17548 944 17588 8800
rect 17548 895 17588 904
rect 17452 811 17492 820
rect 17932 692 17972 39544
rect 18028 26480 18068 26489
rect 18028 24464 18068 26440
rect 18028 24415 18068 24424
rect 18028 24212 18068 24221
rect 18028 21860 18068 24172
rect 18028 21811 18068 21820
rect 17932 643 17972 652
rect 18124 692 18164 40300
rect 18220 31268 18260 31277
rect 18220 27908 18260 31228
rect 18220 27859 18260 27868
rect 18220 23456 18260 23465
rect 18220 22532 18260 23416
rect 18220 22483 18260 22492
rect 18220 8504 18260 8513
rect 18220 7328 18260 8464
rect 18220 5732 18260 7288
rect 18220 5683 18260 5692
rect 18124 643 18164 652
rect 18316 692 18356 40468
rect 20048 40088 20416 40097
rect 20088 40048 20130 40088
rect 20170 40048 20212 40088
rect 20252 40048 20294 40088
rect 20334 40048 20376 40088
rect 20048 40039 20416 40048
rect 19852 39752 19892 39761
rect 18808 39332 19176 39341
rect 18848 39292 18890 39332
rect 18930 39292 18972 39332
rect 19012 39292 19054 39332
rect 19094 39292 19136 39332
rect 18808 39283 19176 39292
rect 19468 39248 19508 39257
rect 18508 38744 18548 38753
rect 18412 29336 18452 29345
rect 18412 27656 18452 29296
rect 18412 27607 18452 27616
rect 18412 26732 18452 26741
rect 18412 24305 18452 26692
rect 18411 24296 18453 24305
rect 18411 24256 18412 24296
rect 18452 24256 18453 24296
rect 18411 24247 18453 24256
rect 18412 23540 18452 23549
rect 18412 18668 18452 23500
rect 18412 18619 18452 18628
rect 18412 9008 18452 9017
rect 18412 8504 18452 8968
rect 18412 8455 18452 8464
rect 18412 8000 18452 8009
rect 18412 4724 18452 7960
rect 18412 3884 18452 4684
rect 18412 3835 18452 3844
rect 18316 643 18356 652
rect 18508 692 18548 38704
rect 19468 38492 19508 39208
rect 19468 38443 19508 38452
rect 19852 38156 19892 39712
rect 19948 38828 19988 38837
rect 19948 38576 19988 38788
rect 19948 38527 19988 38536
rect 20048 38576 20416 38585
rect 20088 38536 20130 38576
rect 20170 38536 20212 38576
rect 20252 38536 20294 38576
rect 20334 38536 20376 38576
rect 20048 38527 20416 38536
rect 19852 38107 19892 38116
rect 20428 38408 20468 38417
rect 18700 38072 18740 38081
rect 18700 37568 18740 38032
rect 19276 37988 19316 37997
rect 18808 37820 19176 37829
rect 18848 37780 18890 37820
rect 18930 37780 18972 37820
rect 19012 37780 19054 37820
rect 19094 37780 19136 37820
rect 18808 37771 19176 37780
rect 18700 37519 18740 37528
rect 18808 36308 19176 36317
rect 18848 36268 18890 36308
rect 18930 36268 18972 36308
rect 19012 36268 19054 36308
rect 19094 36268 19136 36308
rect 18808 36259 19176 36268
rect 18700 35048 18740 35057
rect 18604 30512 18644 30521
rect 18604 27824 18644 30472
rect 18604 27775 18644 27784
rect 18603 24296 18645 24305
rect 18603 24256 18604 24296
rect 18644 24256 18645 24296
rect 18603 24247 18645 24256
rect 18604 16400 18644 24247
rect 18604 16351 18644 16360
rect 18508 643 18548 652
rect 16972 559 17012 568
rect 18700 524 18740 35008
rect 18808 34796 19176 34805
rect 18848 34756 18890 34796
rect 18930 34756 18972 34796
rect 19012 34756 19054 34796
rect 19094 34756 19136 34796
rect 18808 34747 19176 34756
rect 18808 33284 19176 33293
rect 18848 33244 18890 33284
rect 18930 33244 18972 33284
rect 19012 33244 19054 33284
rect 19094 33244 19136 33284
rect 18808 33235 19176 33244
rect 18808 31772 19176 31781
rect 18848 31732 18890 31772
rect 18930 31732 18972 31772
rect 19012 31732 19054 31772
rect 19094 31732 19136 31772
rect 18808 31723 19176 31732
rect 18808 30260 19176 30269
rect 18848 30220 18890 30260
rect 18930 30220 18972 30260
rect 19012 30220 19054 30260
rect 19094 30220 19136 30260
rect 18808 30211 19176 30220
rect 19276 30260 19316 37948
rect 20428 37904 20468 38368
rect 20524 38072 20564 40552
rect 20524 38023 20564 38032
rect 20620 39752 20660 39761
rect 20428 37864 20564 37904
rect 20048 37064 20416 37073
rect 20088 37024 20130 37064
rect 20170 37024 20212 37064
rect 20252 37024 20294 37064
rect 20334 37024 20376 37064
rect 20048 37015 20416 37024
rect 19276 30211 19316 30220
rect 19372 36308 19412 36317
rect 19372 35888 19412 36268
rect 19372 35384 19412 35848
rect 20048 35552 20416 35561
rect 20088 35512 20130 35552
rect 20170 35512 20212 35552
rect 20252 35512 20294 35552
rect 20334 35512 20376 35552
rect 20048 35503 20416 35512
rect 19372 33200 19412 35344
rect 20048 34040 20416 34049
rect 20088 34000 20130 34040
rect 20170 34000 20212 34040
rect 20252 34000 20294 34040
rect 20334 34000 20376 34040
rect 20048 33991 20416 34000
rect 18808 28748 19176 28757
rect 18848 28708 18890 28748
rect 18930 28708 18972 28748
rect 19012 28708 19054 28748
rect 19094 28708 19136 28748
rect 18808 28699 19176 28708
rect 18808 27236 19176 27245
rect 18848 27196 18890 27236
rect 18930 27196 18972 27236
rect 19012 27196 19054 27236
rect 19094 27196 19136 27236
rect 18808 27187 19176 27196
rect 18808 25724 19176 25733
rect 18848 25684 18890 25724
rect 18930 25684 18972 25724
rect 19012 25684 19054 25724
rect 19094 25684 19136 25724
rect 18808 25675 19176 25684
rect 18808 24212 19176 24221
rect 18848 24172 18890 24212
rect 18930 24172 18972 24212
rect 19012 24172 19054 24212
rect 19094 24172 19136 24212
rect 18808 24163 19176 24172
rect 18808 22700 19176 22709
rect 18848 22660 18890 22700
rect 18930 22660 18972 22700
rect 19012 22660 19054 22700
rect 19094 22660 19136 22700
rect 18808 22651 19176 22660
rect 19276 21440 19316 21449
rect 18808 21188 19176 21197
rect 18848 21148 18890 21188
rect 18930 21148 18972 21188
rect 19012 21148 19054 21188
rect 19094 21148 19136 21188
rect 18808 21139 19176 21148
rect 18808 19676 19176 19685
rect 18848 19636 18890 19676
rect 18930 19636 18972 19676
rect 19012 19636 19054 19676
rect 19094 19636 19136 19676
rect 18808 19627 19176 19636
rect 19276 19508 19316 21400
rect 19276 19459 19316 19468
rect 18808 18164 19176 18173
rect 18848 18124 18890 18164
rect 18930 18124 18972 18164
rect 19012 18124 19054 18164
rect 19094 18124 19136 18164
rect 18808 18115 19176 18124
rect 18808 16652 19176 16661
rect 18848 16612 18890 16652
rect 18930 16612 18972 16652
rect 19012 16612 19054 16652
rect 19094 16612 19136 16652
rect 18808 16603 19176 16612
rect 18808 15140 19176 15149
rect 18848 15100 18890 15140
rect 18930 15100 18972 15140
rect 19012 15100 19054 15140
rect 19094 15100 19136 15140
rect 18808 15091 19176 15100
rect 19372 14720 19412 33160
rect 19564 33704 19604 33713
rect 19468 31184 19508 31193
rect 19468 27740 19508 31144
rect 19564 30680 19604 33664
rect 20048 32528 20416 32537
rect 20088 32488 20130 32528
rect 20170 32488 20212 32528
rect 20252 32488 20294 32528
rect 20334 32488 20376 32528
rect 20048 32479 20416 32488
rect 20048 31016 20416 31025
rect 20088 30976 20130 31016
rect 20170 30976 20212 31016
rect 20252 30976 20294 31016
rect 20334 30976 20376 31016
rect 20048 30967 20416 30976
rect 19564 29840 19604 30640
rect 19564 29791 19604 29800
rect 20048 29504 20416 29513
rect 20088 29464 20130 29504
rect 20170 29464 20212 29504
rect 20252 29464 20294 29504
rect 20334 29464 20376 29504
rect 20048 29455 20416 29464
rect 19468 27691 19508 27700
rect 19852 29000 19892 29009
rect 19660 24632 19700 24641
rect 19468 20096 19508 20105
rect 19468 18920 19508 20056
rect 19468 18871 19508 18880
rect 19372 14671 19412 14680
rect 19564 16400 19604 16409
rect 19564 15476 19604 16360
rect 18808 13628 19176 13637
rect 18848 13588 18890 13628
rect 18930 13588 18972 13628
rect 19012 13588 19054 13628
rect 19094 13588 19136 13628
rect 18808 13579 19176 13588
rect 18808 12116 19176 12125
rect 18848 12076 18890 12116
rect 18930 12076 18972 12116
rect 19012 12076 19054 12116
rect 19094 12076 19136 12116
rect 18808 12067 19176 12076
rect 19276 11696 19316 11705
rect 18808 10604 19176 10613
rect 18848 10564 18890 10604
rect 18930 10564 18972 10604
rect 19012 10564 19054 10604
rect 19094 10564 19136 10604
rect 18808 10555 19176 10564
rect 18808 9092 19176 9101
rect 18848 9052 18890 9092
rect 18930 9052 18972 9092
rect 19012 9052 19054 9092
rect 19094 9052 19136 9092
rect 18808 9043 19176 9052
rect 19276 8420 19316 11656
rect 19276 8000 19316 8380
rect 19276 7951 19316 7960
rect 19468 8840 19508 8849
rect 18808 7580 19176 7589
rect 18848 7540 18890 7580
rect 18930 7540 18972 7580
rect 19012 7540 19054 7580
rect 19094 7540 19136 7580
rect 18808 7531 19176 7540
rect 19276 7328 19316 7337
rect 18808 6068 19176 6077
rect 18848 6028 18890 6068
rect 18930 6028 18972 6068
rect 19012 6028 19054 6068
rect 19094 6028 19136 6068
rect 18808 6019 19176 6028
rect 18808 4556 19176 4565
rect 18848 4516 18890 4556
rect 18930 4516 18972 4556
rect 19012 4516 19054 4556
rect 19094 4516 19136 4556
rect 18808 4507 19176 4516
rect 19276 3464 19316 7288
rect 19276 3415 19316 3424
rect 18808 3044 19176 3053
rect 18848 3004 18890 3044
rect 18930 3004 18972 3044
rect 19012 3004 19054 3044
rect 19094 3004 19136 3044
rect 18808 2995 19176 3004
rect 18808 1532 19176 1541
rect 18848 1492 18890 1532
rect 18930 1492 18972 1532
rect 19012 1492 19054 1532
rect 19094 1492 19136 1532
rect 18808 1483 19176 1492
rect 19468 692 19508 8800
rect 19564 7328 19604 15436
rect 19564 7279 19604 7288
rect 19660 4052 19700 24592
rect 19852 17912 19892 28960
rect 20048 27992 20416 28001
rect 20088 27952 20130 27992
rect 20170 27952 20212 27992
rect 20252 27952 20294 27992
rect 20334 27952 20376 27992
rect 20048 27943 20416 27952
rect 20048 26480 20416 26489
rect 20088 26440 20130 26480
rect 20170 26440 20212 26480
rect 20252 26440 20294 26480
rect 20334 26440 20376 26480
rect 20048 26431 20416 26440
rect 20048 24968 20416 24977
rect 20088 24928 20130 24968
rect 20170 24928 20212 24968
rect 20252 24928 20294 24968
rect 20334 24928 20376 24968
rect 20048 24919 20416 24928
rect 20048 23456 20416 23465
rect 20088 23416 20130 23456
rect 20170 23416 20212 23456
rect 20252 23416 20294 23456
rect 20334 23416 20376 23456
rect 20048 23407 20416 23416
rect 20048 21944 20416 21953
rect 20088 21904 20130 21944
rect 20170 21904 20212 21944
rect 20252 21904 20294 21944
rect 20334 21904 20376 21944
rect 20048 21895 20416 21904
rect 19948 21608 19988 21617
rect 19948 20096 19988 21568
rect 20048 20432 20416 20441
rect 20088 20392 20130 20432
rect 20170 20392 20212 20432
rect 20252 20392 20294 20432
rect 20334 20392 20376 20432
rect 20048 20383 20416 20392
rect 19948 20047 19988 20056
rect 20048 18920 20416 18929
rect 20088 18880 20130 18920
rect 20170 18880 20212 18920
rect 20252 18880 20294 18920
rect 20334 18880 20376 18920
rect 20048 18871 20416 18880
rect 19852 17863 19892 17872
rect 20048 17408 20416 17417
rect 20088 17368 20130 17408
rect 20170 17368 20212 17408
rect 20252 17368 20294 17408
rect 20334 17368 20376 17408
rect 20048 17359 20416 17368
rect 20048 15896 20416 15905
rect 20088 15856 20130 15896
rect 20170 15856 20212 15896
rect 20252 15856 20294 15896
rect 20334 15856 20376 15896
rect 20048 15847 20416 15856
rect 20048 14384 20416 14393
rect 20088 14344 20130 14384
rect 20170 14344 20212 14384
rect 20252 14344 20294 14384
rect 20334 14344 20376 14384
rect 20048 14335 20416 14344
rect 20048 12872 20416 12881
rect 20088 12832 20130 12872
rect 20170 12832 20212 12872
rect 20252 12832 20294 12872
rect 20334 12832 20376 12872
rect 20048 12823 20416 12832
rect 20048 11360 20416 11369
rect 20088 11320 20130 11360
rect 20170 11320 20212 11360
rect 20252 11320 20294 11360
rect 20334 11320 20376 11360
rect 20048 11311 20416 11320
rect 20048 9848 20416 9857
rect 20088 9808 20130 9848
rect 20170 9808 20212 9848
rect 20252 9808 20294 9848
rect 20334 9808 20376 9848
rect 20048 9799 20416 9808
rect 20048 8336 20416 8345
rect 20088 8296 20130 8336
rect 20170 8296 20212 8336
rect 20252 8296 20294 8336
rect 20334 8296 20376 8336
rect 20048 8287 20416 8296
rect 20048 6824 20416 6833
rect 20088 6784 20130 6824
rect 20170 6784 20212 6824
rect 20252 6784 20294 6824
rect 20334 6784 20376 6824
rect 20048 6775 20416 6784
rect 19947 6320 19989 6329
rect 19947 6280 19948 6320
rect 19988 6280 19989 6320
rect 19947 6271 19989 6280
rect 19948 6186 19988 6271
rect 20048 5312 20416 5321
rect 20088 5272 20130 5312
rect 20170 5272 20212 5312
rect 20252 5272 20294 5312
rect 20334 5272 20376 5312
rect 20048 5263 20416 5272
rect 19660 4003 19700 4012
rect 20048 3800 20416 3809
rect 20088 3760 20130 3800
rect 20170 3760 20212 3800
rect 20252 3760 20294 3800
rect 20334 3760 20376 3800
rect 20048 3751 20416 3760
rect 20048 2288 20416 2297
rect 20088 2248 20130 2288
rect 20170 2248 20212 2288
rect 20252 2248 20294 2288
rect 20334 2248 20376 2288
rect 20048 2239 20416 2248
rect 20524 1196 20564 37864
rect 20620 1364 20660 39712
rect 20908 37232 20948 37241
rect 20908 35552 20948 37192
rect 20908 35503 20948 35512
rect 20716 22112 20756 22121
rect 20716 16400 20756 22072
rect 20907 18332 20949 18341
rect 20907 18292 20908 18332
rect 20948 18292 20949 18332
rect 20907 18283 20949 18292
rect 20908 16904 20948 18283
rect 20908 16855 20948 16864
rect 20716 16351 20756 16360
rect 20716 13880 20756 13889
rect 20716 10100 20756 13840
rect 20716 10051 20756 10060
rect 21004 12368 21044 12377
rect 21004 9176 21044 12328
rect 21004 9127 21044 9136
rect 20620 1315 20660 1324
rect 20524 1147 20564 1156
rect 20048 776 20416 785
rect 20088 736 20130 776
rect 20170 736 20212 776
rect 20252 736 20294 776
rect 20334 736 20376 776
rect 20048 727 20416 736
rect 19468 643 19508 652
rect 18700 475 18740 484
rect 14284 307 14324 316
rect 11500 223 11540 232
rect 5260 138 5300 223
<< via4 >>
rect 1228 36520 1268 36560
rect 1132 35848 1172 35888
rect 1036 33832 1076 33872
rect 1516 28792 1556 28832
rect 1804 28792 1844 28832
rect 3244 40300 3284 40340
rect 2956 38368 2996 38408
rect 2764 35680 2804 35720
rect 1612 19216 1652 19256
rect 2476 25180 2516 25220
rect 2380 17704 2420 17744
rect 2188 1240 2228 1280
rect 3688 40804 3728 40844
rect 3770 40804 3810 40844
rect 3852 40804 3892 40844
rect 3934 40804 3974 40844
rect 4016 40804 4056 40844
rect 3532 39628 3572 39668
rect 3436 19216 3476 19256
rect 3148 1240 3188 1280
rect 3688 39292 3728 39332
rect 3770 39292 3810 39332
rect 3852 39292 3892 39332
rect 3934 39292 3974 39332
rect 4016 39292 4056 39332
rect 3820 37948 3860 37988
rect 3688 37780 3728 37820
rect 3770 37780 3810 37820
rect 3852 37780 3892 37820
rect 3934 37780 3974 37820
rect 4016 37780 4056 37820
rect 4928 41560 4968 41600
rect 5010 41560 5050 41600
rect 5092 41560 5132 41600
rect 5174 41560 5214 41600
rect 5256 41560 5296 41600
rect 3688 36268 3728 36308
rect 3770 36268 3810 36308
rect 3852 36268 3892 36308
rect 3934 36268 3974 36308
rect 4016 36268 4056 36308
rect 4012 35680 4052 35720
rect 3688 34756 3728 34796
rect 3770 34756 3810 34796
rect 3852 34756 3892 34796
rect 3934 34756 3974 34796
rect 4016 34756 4056 34796
rect 3688 33244 3728 33284
rect 3770 33244 3810 33284
rect 3852 33244 3892 33284
rect 3934 33244 3974 33284
rect 4016 33244 4056 33284
rect 3688 31732 3728 31772
rect 3770 31732 3810 31772
rect 3852 31732 3892 31772
rect 3934 31732 3974 31772
rect 4016 31732 4056 31772
rect 3688 30220 3728 30260
rect 3770 30220 3810 30260
rect 3852 30220 3892 30260
rect 3934 30220 3974 30260
rect 4016 30220 4056 30260
rect 4588 37528 4628 37568
rect 4928 40048 4968 40088
rect 5010 40048 5050 40088
rect 5092 40048 5132 40088
rect 5174 40048 5214 40088
rect 5256 40048 5296 40088
rect 5068 39628 5108 39668
rect 5356 39628 5396 39668
rect 4972 38956 5012 38996
rect 4928 38536 4968 38576
rect 5010 38536 5050 38576
rect 5092 38536 5132 38576
rect 5174 38536 5214 38576
rect 5256 38536 5296 38576
rect 4928 37024 4968 37064
rect 5010 37024 5050 37064
rect 5092 37024 5132 37064
rect 5174 37024 5214 37064
rect 5256 37024 5296 37064
rect 4780 36604 4820 36644
rect 3688 28708 3728 28748
rect 3770 28708 3810 28748
rect 3852 28708 3892 28748
rect 3934 28708 3974 28748
rect 4016 28708 4056 28748
rect 3688 27196 3728 27236
rect 3770 27196 3810 27236
rect 3852 27196 3892 27236
rect 3934 27196 3974 27236
rect 4016 27196 4056 27236
rect 3688 25684 3728 25724
rect 3770 25684 3810 25724
rect 3852 25684 3892 25724
rect 3934 25684 3974 25724
rect 4016 25684 4056 25724
rect 4012 25180 4052 25220
rect 3688 24172 3728 24212
rect 3770 24172 3810 24212
rect 3852 24172 3892 24212
rect 3934 24172 3974 24212
rect 4016 24172 4056 24212
rect 3688 22660 3728 22700
rect 3770 22660 3810 22700
rect 3852 22660 3892 22700
rect 3934 22660 3974 22700
rect 4016 22660 4056 22700
rect 3688 21148 3728 21188
rect 3770 21148 3810 21188
rect 3852 21148 3892 21188
rect 3934 21148 3974 21188
rect 4016 21148 4056 21188
rect 3688 19636 3728 19676
rect 3770 19636 3810 19676
rect 3852 19636 3892 19676
rect 3934 19636 3974 19676
rect 4016 19636 4056 19676
rect 3688 18124 3728 18164
rect 3770 18124 3810 18164
rect 3852 18124 3892 18164
rect 3934 18124 3974 18164
rect 4016 18124 4056 18164
rect 3688 16612 3728 16652
rect 3770 16612 3810 16652
rect 3852 16612 3892 16652
rect 3934 16612 3974 16652
rect 4016 16612 4056 16652
rect 3688 15100 3728 15140
rect 3770 15100 3810 15140
rect 3852 15100 3892 15140
rect 3934 15100 3974 15140
rect 4016 15100 4056 15140
rect 3688 13588 3728 13628
rect 3770 13588 3810 13628
rect 3852 13588 3892 13628
rect 3934 13588 3974 13628
rect 4016 13588 4056 13628
rect 3688 12076 3728 12116
rect 3770 12076 3810 12116
rect 3852 12076 3892 12116
rect 3934 12076 3974 12116
rect 4016 12076 4056 12116
rect 3688 10564 3728 10604
rect 3770 10564 3810 10604
rect 3852 10564 3892 10604
rect 3934 10564 3974 10604
rect 4016 10564 4056 10604
rect 3688 9052 3728 9092
rect 3770 9052 3810 9092
rect 3852 9052 3892 9092
rect 3934 9052 3974 9092
rect 4016 9052 4056 9092
rect 4876 35848 4916 35888
rect 4928 35512 4968 35552
rect 5010 35512 5050 35552
rect 5092 35512 5132 35552
rect 5174 35512 5214 35552
rect 5256 35512 5296 35552
rect 4928 34000 4968 34040
rect 5010 34000 5050 34040
rect 5092 34000 5132 34040
rect 5174 34000 5214 34040
rect 5256 34000 5296 34040
rect 4928 32488 4968 32528
rect 5010 32488 5050 32528
rect 5092 32488 5132 32528
rect 5174 32488 5214 32528
rect 5256 32488 5296 32528
rect 4928 30976 4968 31016
rect 5010 30976 5050 31016
rect 5092 30976 5132 31016
rect 5174 30976 5214 31016
rect 5256 30976 5296 31016
rect 4928 29464 4968 29504
rect 5010 29464 5050 29504
rect 5092 29464 5132 29504
rect 5174 29464 5214 29504
rect 5256 29464 5296 29504
rect 4928 27952 4968 27992
rect 5010 27952 5050 27992
rect 5092 27952 5132 27992
rect 5174 27952 5214 27992
rect 5256 27952 5296 27992
rect 4928 26440 4968 26480
rect 5010 26440 5050 26480
rect 5092 26440 5132 26480
rect 5174 26440 5214 26480
rect 5256 26440 5296 26480
rect 4928 24928 4968 24968
rect 5010 24928 5050 24968
rect 5092 24928 5132 24968
rect 5174 24928 5214 24968
rect 5256 24928 5296 24968
rect 4928 23416 4968 23456
rect 5010 23416 5050 23456
rect 5092 23416 5132 23456
rect 5174 23416 5214 23456
rect 5256 23416 5296 23456
rect 4928 21904 4968 21944
rect 5010 21904 5050 21944
rect 5092 21904 5132 21944
rect 5174 21904 5214 21944
rect 5256 21904 5296 21944
rect 4928 20392 4968 20432
rect 5010 20392 5050 20432
rect 5092 20392 5132 20432
rect 5174 20392 5214 20432
rect 5256 20392 5296 20432
rect 4928 18880 4968 18920
rect 5010 18880 5050 18920
rect 5092 18880 5132 18920
rect 5174 18880 5214 18920
rect 5256 18880 5296 18920
rect 4928 17368 4968 17408
rect 5010 17368 5050 17408
rect 5092 17368 5132 17408
rect 5174 17368 5214 17408
rect 5256 17368 5296 17408
rect 3688 7540 3728 7580
rect 3770 7540 3810 7580
rect 3852 7540 3892 7580
rect 3934 7540 3974 7580
rect 4016 7540 4056 7580
rect 3688 6028 3728 6068
rect 3770 6028 3810 6068
rect 3852 6028 3892 6068
rect 3934 6028 3974 6068
rect 4016 6028 4056 6068
rect 4928 15856 4968 15896
rect 5010 15856 5050 15896
rect 5092 15856 5132 15896
rect 5174 15856 5214 15896
rect 5256 15856 5296 15896
rect 4928 14344 4968 14384
rect 5010 14344 5050 14384
rect 5092 14344 5132 14384
rect 5174 14344 5214 14384
rect 5256 14344 5296 14384
rect 4928 12832 4968 12872
rect 5010 12832 5050 12872
rect 5092 12832 5132 12872
rect 5174 12832 5214 12872
rect 5256 12832 5296 12872
rect 4928 11320 4968 11360
rect 5010 11320 5050 11360
rect 5092 11320 5132 11360
rect 5174 11320 5214 11360
rect 5256 11320 5296 11360
rect 4396 6280 4436 6320
rect 4928 9808 4968 9848
rect 5010 9808 5050 9848
rect 5092 9808 5132 9848
rect 5174 9808 5214 9848
rect 5256 9808 5296 9848
rect 4928 8296 4968 8336
rect 5010 8296 5050 8336
rect 5092 8296 5132 8336
rect 5174 8296 5214 8336
rect 5256 8296 5296 8336
rect 3688 4516 3728 4556
rect 3770 4516 3810 4556
rect 3852 4516 3892 4556
rect 3934 4516 3974 4556
rect 4016 4516 4056 4556
rect 3688 3004 3728 3044
rect 3770 3004 3810 3044
rect 3852 3004 3892 3044
rect 3934 3004 3974 3044
rect 4016 3004 4056 3044
rect 4928 6784 4968 6824
rect 5010 6784 5050 6824
rect 5092 6784 5132 6824
rect 5174 6784 5214 6824
rect 5256 6784 5296 6824
rect 4928 5272 4968 5312
rect 5010 5272 5050 5312
rect 5092 5272 5132 5312
rect 5174 5272 5214 5312
rect 5256 5272 5296 5312
rect 4928 3760 4968 3800
rect 5010 3760 5050 3800
rect 5092 3760 5132 3800
rect 5174 3760 5214 3800
rect 5256 3760 5296 3800
rect 4928 2248 4968 2288
rect 5010 2248 5050 2288
rect 5092 2248 5132 2288
rect 5174 2248 5214 2288
rect 5256 2248 5296 2288
rect 3688 1492 3728 1532
rect 3770 1492 3810 1532
rect 3852 1492 3892 1532
rect 3934 1492 3974 1532
rect 4016 1492 4056 1532
rect 4928 736 4968 776
rect 5010 736 5050 776
rect 5092 736 5132 776
rect 5174 736 5214 776
rect 5256 736 5296 776
rect 5740 38956 5780 38996
rect 5548 37528 5588 37568
rect 5452 36604 5492 36644
rect 5644 37192 5684 37232
rect 5548 36520 5588 36560
rect 5644 33832 5684 33872
rect 5836 37108 5876 37148
rect 5740 32740 5780 32780
rect 5548 19216 5588 19256
rect 6892 40300 6932 40340
rect 7372 40300 7412 40340
rect 6796 39628 6836 39668
rect 6604 904 6644 944
rect 6988 37528 7028 37568
rect 7084 36604 7124 36644
rect 7948 38368 7988 38408
rect 8140 37192 8180 37232
rect 8812 37948 8852 37988
rect 10156 17704 10196 17744
rect 10636 37948 10676 37988
rect 10444 37108 10484 37148
rect 10828 36604 10868 36644
rect 11116 18292 11156 18332
rect 5260 232 5300 272
rect 8428 232 8468 272
rect 20048 41560 20088 41600
rect 20130 41560 20170 41600
rect 20212 41560 20252 41600
rect 20294 41560 20334 41600
rect 20376 41560 20416 41600
rect 18808 40804 18848 40844
rect 18890 40804 18930 40844
rect 18972 40804 19012 40844
rect 19054 40804 19094 40844
rect 19136 40804 19176 40844
rect 20048 40048 20088 40088
rect 20130 40048 20170 40088
rect 20212 40048 20252 40088
rect 20294 40048 20334 40088
rect 20376 40048 20416 40088
rect 18808 39292 18848 39332
rect 18890 39292 18930 39332
rect 18972 39292 19012 39332
rect 19054 39292 19094 39332
rect 19136 39292 19176 39332
rect 18412 24256 18452 24296
rect 20048 38536 20088 38576
rect 20130 38536 20170 38576
rect 20212 38536 20252 38576
rect 20294 38536 20334 38576
rect 20376 38536 20416 38576
rect 18808 37780 18848 37820
rect 18890 37780 18930 37820
rect 18972 37780 19012 37820
rect 19054 37780 19094 37820
rect 19136 37780 19176 37820
rect 18808 36268 18848 36308
rect 18890 36268 18930 36308
rect 18972 36268 19012 36308
rect 19054 36268 19094 36308
rect 19136 36268 19176 36308
rect 18604 24256 18644 24296
rect 18808 34756 18848 34796
rect 18890 34756 18930 34796
rect 18972 34756 19012 34796
rect 19054 34756 19094 34796
rect 19136 34756 19176 34796
rect 18808 33244 18848 33284
rect 18890 33244 18930 33284
rect 18972 33244 19012 33284
rect 19054 33244 19094 33284
rect 19136 33244 19176 33284
rect 18808 31732 18848 31772
rect 18890 31732 18930 31772
rect 18972 31732 19012 31772
rect 19054 31732 19094 31772
rect 19136 31732 19176 31772
rect 18808 30220 18848 30260
rect 18890 30220 18930 30260
rect 18972 30220 19012 30260
rect 19054 30220 19094 30260
rect 19136 30220 19176 30260
rect 20048 37024 20088 37064
rect 20130 37024 20170 37064
rect 20212 37024 20252 37064
rect 20294 37024 20334 37064
rect 20376 37024 20416 37064
rect 20048 35512 20088 35552
rect 20130 35512 20170 35552
rect 20212 35512 20252 35552
rect 20294 35512 20334 35552
rect 20376 35512 20416 35552
rect 20048 34000 20088 34040
rect 20130 34000 20170 34040
rect 20212 34000 20252 34040
rect 20294 34000 20334 34040
rect 20376 34000 20416 34040
rect 18808 28708 18848 28748
rect 18890 28708 18930 28748
rect 18972 28708 19012 28748
rect 19054 28708 19094 28748
rect 19136 28708 19176 28748
rect 18808 27196 18848 27236
rect 18890 27196 18930 27236
rect 18972 27196 19012 27236
rect 19054 27196 19094 27236
rect 19136 27196 19176 27236
rect 18808 25684 18848 25724
rect 18890 25684 18930 25724
rect 18972 25684 19012 25724
rect 19054 25684 19094 25724
rect 19136 25684 19176 25724
rect 18808 24172 18848 24212
rect 18890 24172 18930 24212
rect 18972 24172 19012 24212
rect 19054 24172 19094 24212
rect 19136 24172 19176 24212
rect 18808 22660 18848 22700
rect 18890 22660 18930 22700
rect 18972 22660 19012 22700
rect 19054 22660 19094 22700
rect 19136 22660 19176 22700
rect 18808 21148 18848 21188
rect 18890 21148 18930 21188
rect 18972 21148 19012 21188
rect 19054 21148 19094 21188
rect 19136 21148 19176 21188
rect 18808 19636 18848 19676
rect 18890 19636 18930 19676
rect 18972 19636 19012 19676
rect 19054 19636 19094 19676
rect 19136 19636 19176 19676
rect 18808 18124 18848 18164
rect 18890 18124 18930 18164
rect 18972 18124 19012 18164
rect 19054 18124 19094 18164
rect 19136 18124 19176 18164
rect 18808 16612 18848 16652
rect 18890 16612 18930 16652
rect 18972 16612 19012 16652
rect 19054 16612 19094 16652
rect 19136 16612 19176 16652
rect 18808 15100 18848 15140
rect 18890 15100 18930 15140
rect 18972 15100 19012 15140
rect 19054 15100 19094 15140
rect 19136 15100 19176 15140
rect 20048 32488 20088 32528
rect 20130 32488 20170 32528
rect 20212 32488 20252 32528
rect 20294 32488 20334 32528
rect 20376 32488 20416 32528
rect 20048 30976 20088 31016
rect 20130 30976 20170 31016
rect 20212 30976 20252 31016
rect 20294 30976 20334 31016
rect 20376 30976 20416 31016
rect 20048 29464 20088 29504
rect 20130 29464 20170 29504
rect 20212 29464 20252 29504
rect 20294 29464 20334 29504
rect 20376 29464 20416 29504
rect 18808 13588 18848 13628
rect 18890 13588 18930 13628
rect 18972 13588 19012 13628
rect 19054 13588 19094 13628
rect 19136 13588 19176 13628
rect 18808 12076 18848 12116
rect 18890 12076 18930 12116
rect 18972 12076 19012 12116
rect 19054 12076 19094 12116
rect 19136 12076 19176 12116
rect 18808 10564 18848 10604
rect 18890 10564 18930 10604
rect 18972 10564 19012 10604
rect 19054 10564 19094 10604
rect 19136 10564 19176 10604
rect 18808 9052 18848 9092
rect 18890 9052 18930 9092
rect 18972 9052 19012 9092
rect 19054 9052 19094 9092
rect 19136 9052 19176 9092
rect 18808 7540 18848 7580
rect 18890 7540 18930 7580
rect 18972 7540 19012 7580
rect 19054 7540 19094 7580
rect 19136 7540 19176 7580
rect 18808 6028 18848 6068
rect 18890 6028 18930 6068
rect 18972 6028 19012 6068
rect 19054 6028 19094 6068
rect 19136 6028 19176 6068
rect 18808 4516 18848 4556
rect 18890 4516 18930 4556
rect 18972 4516 19012 4556
rect 19054 4516 19094 4556
rect 19136 4516 19176 4556
rect 18808 3004 18848 3044
rect 18890 3004 18930 3044
rect 18972 3004 19012 3044
rect 19054 3004 19094 3044
rect 19136 3004 19176 3044
rect 18808 1492 18848 1532
rect 18890 1492 18930 1532
rect 18972 1492 19012 1532
rect 19054 1492 19094 1532
rect 19136 1492 19176 1532
rect 20048 27952 20088 27992
rect 20130 27952 20170 27992
rect 20212 27952 20252 27992
rect 20294 27952 20334 27992
rect 20376 27952 20416 27992
rect 20048 26440 20088 26480
rect 20130 26440 20170 26480
rect 20212 26440 20252 26480
rect 20294 26440 20334 26480
rect 20376 26440 20416 26480
rect 20048 24928 20088 24968
rect 20130 24928 20170 24968
rect 20212 24928 20252 24968
rect 20294 24928 20334 24968
rect 20376 24928 20416 24968
rect 20048 23416 20088 23456
rect 20130 23416 20170 23456
rect 20212 23416 20252 23456
rect 20294 23416 20334 23456
rect 20376 23416 20416 23456
rect 20048 21904 20088 21944
rect 20130 21904 20170 21944
rect 20212 21904 20252 21944
rect 20294 21904 20334 21944
rect 20376 21904 20416 21944
rect 20048 20392 20088 20432
rect 20130 20392 20170 20432
rect 20212 20392 20252 20432
rect 20294 20392 20334 20432
rect 20376 20392 20416 20432
rect 20048 18880 20088 18920
rect 20130 18880 20170 18920
rect 20212 18880 20252 18920
rect 20294 18880 20334 18920
rect 20376 18880 20416 18920
rect 20048 17368 20088 17408
rect 20130 17368 20170 17408
rect 20212 17368 20252 17408
rect 20294 17368 20334 17408
rect 20376 17368 20416 17408
rect 20048 15856 20088 15896
rect 20130 15856 20170 15896
rect 20212 15856 20252 15896
rect 20294 15856 20334 15896
rect 20376 15856 20416 15896
rect 20048 14344 20088 14384
rect 20130 14344 20170 14384
rect 20212 14344 20252 14384
rect 20294 14344 20334 14384
rect 20376 14344 20416 14384
rect 20048 12832 20088 12872
rect 20130 12832 20170 12872
rect 20212 12832 20252 12872
rect 20294 12832 20334 12872
rect 20376 12832 20416 12872
rect 20048 11320 20088 11360
rect 20130 11320 20170 11360
rect 20212 11320 20252 11360
rect 20294 11320 20334 11360
rect 20376 11320 20416 11360
rect 20048 9808 20088 9848
rect 20130 9808 20170 9848
rect 20212 9808 20252 9848
rect 20294 9808 20334 9848
rect 20376 9808 20416 9848
rect 20048 8296 20088 8336
rect 20130 8296 20170 8336
rect 20212 8296 20252 8336
rect 20294 8296 20334 8336
rect 20376 8296 20416 8336
rect 20048 6784 20088 6824
rect 20130 6784 20170 6824
rect 20212 6784 20252 6824
rect 20294 6784 20334 6824
rect 20376 6784 20416 6824
rect 19948 6280 19988 6320
rect 20048 5272 20088 5312
rect 20130 5272 20170 5312
rect 20212 5272 20252 5312
rect 20294 5272 20334 5312
rect 20376 5272 20416 5312
rect 20048 3760 20088 3800
rect 20130 3760 20170 3800
rect 20212 3760 20252 3800
rect 20294 3760 20334 3800
rect 20376 3760 20416 3800
rect 20048 2248 20088 2288
rect 20130 2248 20170 2288
rect 20212 2248 20252 2288
rect 20294 2248 20334 2288
rect 20376 2248 20416 2288
rect 20908 18292 20948 18332
rect 20048 736 20088 776
rect 20130 736 20170 776
rect 20212 736 20252 776
rect 20294 736 20334 776
rect 20376 736 20416 776
<< metal5 >>
rect 4919 41623 5305 41642
rect 4919 41600 4985 41623
rect 5071 41600 5153 41623
rect 5239 41600 5305 41623
rect 4919 41560 4928 41600
rect 4968 41560 4985 41600
rect 5071 41560 5092 41600
rect 5132 41560 5153 41600
rect 5239 41560 5256 41600
rect 5296 41560 5305 41600
rect 4919 41537 4985 41560
rect 5071 41537 5153 41560
rect 5239 41537 5305 41560
rect 4919 41518 5305 41537
rect 20039 41623 20425 41642
rect 20039 41600 20105 41623
rect 20191 41600 20273 41623
rect 20359 41600 20425 41623
rect 20039 41560 20048 41600
rect 20088 41560 20105 41600
rect 20191 41560 20212 41600
rect 20252 41560 20273 41600
rect 20359 41560 20376 41600
rect 20416 41560 20425 41600
rect 20039 41537 20105 41560
rect 20191 41537 20273 41560
rect 20359 41537 20425 41560
rect 20039 41518 20425 41537
rect 3679 40867 4065 40886
rect 3679 40844 3745 40867
rect 3831 40844 3913 40867
rect 3999 40844 4065 40867
rect 3679 40804 3688 40844
rect 3728 40804 3745 40844
rect 3831 40804 3852 40844
rect 3892 40804 3913 40844
rect 3999 40804 4016 40844
rect 4056 40804 4065 40844
rect 3679 40781 3745 40804
rect 3831 40781 3913 40804
rect 3999 40781 4065 40804
rect 3679 40762 4065 40781
rect 18799 40867 19185 40886
rect 18799 40844 18865 40867
rect 18951 40844 19033 40867
rect 19119 40844 19185 40867
rect 18799 40804 18808 40844
rect 18848 40804 18865 40844
rect 18951 40804 18972 40844
rect 19012 40804 19033 40844
rect 19119 40804 19136 40844
rect 19176 40804 19185 40844
rect 18799 40781 18865 40804
rect 18951 40781 19033 40804
rect 19119 40781 19185 40804
rect 18799 40762 19185 40781
rect 3235 40300 3244 40340
rect 3284 40300 6892 40340
rect 6932 40300 7372 40340
rect 7412 40300 7421 40340
rect 4919 40111 5305 40130
rect 4919 40088 4985 40111
rect 5071 40088 5153 40111
rect 5239 40088 5305 40111
rect 4919 40048 4928 40088
rect 4968 40048 4985 40088
rect 5071 40048 5092 40088
rect 5132 40048 5153 40088
rect 5239 40048 5256 40088
rect 5296 40048 5305 40088
rect 4919 40025 4985 40048
rect 5071 40025 5153 40048
rect 5239 40025 5305 40048
rect 4919 40006 5305 40025
rect 20039 40111 20425 40130
rect 20039 40088 20105 40111
rect 20191 40088 20273 40111
rect 20359 40088 20425 40111
rect 20039 40048 20048 40088
rect 20088 40048 20105 40088
rect 20191 40048 20212 40088
rect 20252 40048 20273 40088
rect 20359 40048 20376 40088
rect 20416 40048 20425 40088
rect 20039 40025 20105 40048
rect 20191 40025 20273 40048
rect 20359 40025 20425 40048
rect 20039 40006 20425 40025
rect 3523 39628 3532 39668
rect 3572 39628 5068 39668
rect 5108 39628 5117 39668
rect 5347 39628 5356 39668
rect 5396 39628 6796 39668
rect 6836 39628 6845 39668
rect 3679 39355 4065 39374
rect 3679 39332 3745 39355
rect 3831 39332 3913 39355
rect 3999 39332 4065 39355
rect 3679 39292 3688 39332
rect 3728 39292 3745 39332
rect 3831 39292 3852 39332
rect 3892 39292 3913 39332
rect 3999 39292 4016 39332
rect 4056 39292 4065 39332
rect 3679 39269 3745 39292
rect 3831 39269 3913 39292
rect 3999 39269 4065 39292
rect 3679 39250 4065 39269
rect 18799 39355 19185 39374
rect 18799 39332 18865 39355
rect 18951 39332 19033 39355
rect 19119 39332 19185 39355
rect 18799 39292 18808 39332
rect 18848 39292 18865 39332
rect 18951 39292 18972 39332
rect 19012 39292 19033 39332
rect 19119 39292 19136 39332
rect 19176 39292 19185 39332
rect 18799 39269 18865 39292
rect 18951 39269 19033 39292
rect 19119 39269 19185 39292
rect 18799 39250 19185 39269
rect 4963 38956 4972 38996
rect 5012 38956 5740 38996
rect 5780 38956 5789 38996
rect 4919 38599 5305 38618
rect 4919 38576 4985 38599
rect 5071 38576 5153 38599
rect 5239 38576 5305 38599
rect 4919 38536 4928 38576
rect 4968 38536 4985 38576
rect 5071 38536 5092 38576
rect 5132 38536 5153 38576
rect 5239 38536 5256 38576
rect 5296 38536 5305 38576
rect 4919 38513 4985 38536
rect 5071 38513 5153 38536
rect 5239 38513 5305 38536
rect 4919 38494 5305 38513
rect 20039 38599 20425 38618
rect 20039 38576 20105 38599
rect 20191 38576 20273 38599
rect 20359 38576 20425 38599
rect 20039 38536 20048 38576
rect 20088 38536 20105 38576
rect 20191 38536 20212 38576
rect 20252 38536 20273 38576
rect 20359 38536 20376 38576
rect 20416 38536 20425 38576
rect 20039 38513 20105 38536
rect 20191 38513 20273 38536
rect 20359 38513 20425 38536
rect 20039 38494 20425 38513
rect 2947 38368 2956 38408
rect 2996 38368 7948 38408
rect 7988 38368 7997 38408
rect 3811 37948 3820 37988
rect 3860 37948 8812 37988
rect 8852 37948 10636 37988
rect 10676 37948 10685 37988
rect 3679 37843 4065 37862
rect 3679 37820 3745 37843
rect 3831 37820 3913 37843
rect 3999 37820 4065 37843
rect 3679 37780 3688 37820
rect 3728 37780 3745 37820
rect 3831 37780 3852 37820
rect 3892 37780 3913 37820
rect 3999 37780 4016 37820
rect 4056 37780 4065 37820
rect 3679 37757 3745 37780
rect 3831 37757 3913 37780
rect 3999 37757 4065 37780
rect 3679 37738 4065 37757
rect 18799 37843 19185 37862
rect 18799 37820 18865 37843
rect 18951 37820 19033 37843
rect 19119 37820 19185 37843
rect 18799 37780 18808 37820
rect 18848 37780 18865 37820
rect 18951 37780 18972 37820
rect 19012 37780 19033 37820
rect 19119 37780 19136 37820
rect 19176 37780 19185 37820
rect 18799 37757 18865 37780
rect 18951 37757 19033 37780
rect 19119 37757 19185 37780
rect 18799 37738 19185 37757
rect 4579 37528 4588 37568
rect 4628 37528 5548 37568
rect 5588 37528 6988 37568
rect 7028 37528 7037 37568
rect 5635 37192 5644 37232
rect 5684 37192 8140 37232
rect 8180 37192 8189 37232
rect 5827 37108 5836 37148
rect 5876 37108 10444 37148
rect 10484 37108 10493 37148
rect 4919 37087 5305 37106
rect 4919 37064 4985 37087
rect 5071 37064 5153 37087
rect 5239 37064 5305 37087
rect 4919 37024 4928 37064
rect 4968 37024 4985 37064
rect 5071 37024 5092 37064
rect 5132 37024 5153 37064
rect 5239 37024 5256 37064
rect 5296 37024 5305 37064
rect 4919 37001 4985 37024
rect 5071 37001 5153 37024
rect 5239 37001 5305 37024
rect 4919 36982 5305 37001
rect 20039 37087 20425 37106
rect 20039 37064 20105 37087
rect 20191 37064 20273 37087
rect 20359 37064 20425 37087
rect 20039 37024 20048 37064
rect 20088 37024 20105 37064
rect 20191 37024 20212 37064
rect 20252 37024 20273 37064
rect 20359 37024 20376 37064
rect 20416 37024 20425 37064
rect 20039 37001 20105 37024
rect 20191 37001 20273 37024
rect 20359 37001 20425 37024
rect 20039 36982 20425 37001
rect 4771 36604 4780 36644
rect 4820 36604 5452 36644
rect 5492 36604 5501 36644
rect 7075 36604 7084 36644
rect 7124 36604 10828 36644
rect 10868 36604 10877 36644
rect 1219 36520 1228 36560
rect 1268 36520 5548 36560
rect 5588 36520 5597 36560
rect 3679 36331 4065 36350
rect 3679 36308 3745 36331
rect 3831 36308 3913 36331
rect 3999 36308 4065 36331
rect 3679 36268 3688 36308
rect 3728 36268 3745 36308
rect 3831 36268 3852 36308
rect 3892 36268 3913 36308
rect 3999 36268 4016 36308
rect 4056 36268 4065 36308
rect 3679 36245 3745 36268
rect 3831 36245 3913 36268
rect 3999 36245 4065 36268
rect 3679 36226 4065 36245
rect 18799 36331 19185 36350
rect 18799 36308 18865 36331
rect 18951 36308 19033 36331
rect 19119 36308 19185 36331
rect 18799 36268 18808 36308
rect 18848 36268 18865 36308
rect 18951 36268 18972 36308
rect 19012 36268 19033 36308
rect 19119 36268 19136 36308
rect 19176 36268 19185 36308
rect 18799 36245 18865 36268
rect 18951 36245 19033 36268
rect 19119 36245 19185 36268
rect 18799 36226 19185 36245
rect 1123 35848 1132 35888
rect 1172 35848 4876 35888
rect 4916 35848 4925 35888
rect 2755 35680 2764 35720
rect 2804 35680 4012 35720
rect 4052 35680 4061 35720
rect 4919 35575 5305 35594
rect 4919 35552 4985 35575
rect 5071 35552 5153 35575
rect 5239 35552 5305 35575
rect 4919 35512 4928 35552
rect 4968 35512 4985 35552
rect 5071 35512 5092 35552
rect 5132 35512 5153 35552
rect 5239 35512 5256 35552
rect 5296 35512 5305 35552
rect 4919 35489 4985 35512
rect 5071 35489 5153 35512
rect 5239 35489 5305 35512
rect 4919 35470 5305 35489
rect 20039 35575 20425 35594
rect 20039 35552 20105 35575
rect 20191 35552 20273 35575
rect 20359 35552 20425 35575
rect 20039 35512 20048 35552
rect 20088 35512 20105 35552
rect 20191 35512 20212 35552
rect 20252 35512 20273 35552
rect 20359 35512 20376 35552
rect 20416 35512 20425 35552
rect 20039 35489 20105 35512
rect 20191 35489 20273 35512
rect 20359 35489 20425 35512
rect 20039 35470 20425 35489
rect 3679 34819 4065 34838
rect 3679 34796 3745 34819
rect 3831 34796 3913 34819
rect 3999 34796 4065 34819
rect 3679 34756 3688 34796
rect 3728 34756 3745 34796
rect 3831 34756 3852 34796
rect 3892 34756 3913 34796
rect 3999 34756 4016 34796
rect 4056 34756 4065 34796
rect 3679 34733 3745 34756
rect 3831 34733 3913 34756
rect 3999 34733 4065 34756
rect 3679 34714 4065 34733
rect 18799 34819 19185 34838
rect 18799 34796 18865 34819
rect 18951 34796 19033 34819
rect 19119 34796 19185 34819
rect 18799 34756 18808 34796
rect 18848 34756 18865 34796
rect 18951 34756 18972 34796
rect 19012 34756 19033 34796
rect 19119 34756 19136 34796
rect 19176 34756 19185 34796
rect 18799 34733 18865 34756
rect 18951 34733 19033 34756
rect 19119 34733 19185 34756
rect 18799 34714 19185 34733
rect 4919 34063 5305 34082
rect 4919 34040 4985 34063
rect 5071 34040 5153 34063
rect 5239 34040 5305 34063
rect 4919 34000 4928 34040
rect 4968 34000 4985 34040
rect 5071 34000 5092 34040
rect 5132 34000 5153 34040
rect 5239 34000 5256 34040
rect 5296 34000 5305 34040
rect 4919 33977 4985 34000
rect 5071 33977 5153 34000
rect 5239 33977 5305 34000
rect 4919 33958 5305 33977
rect 20039 34063 20425 34082
rect 20039 34040 20105 34063
rect 20191 34040 20273 34063
rect 20359 34040 20425 34063
rect 20039 34000 20048 34040
rect 20088 34000 20105 34040
rect 20191 34000 20212 34040
rect 20252 34000 20273 34040
rect 20359 34000 20376 34040
rect 20416 34000 20425 34040
rect 20039 33977 20105 34000
rect 20191 33977 20273 34000
rect 20359 33977 20425 34000
rect 20039 33958 20425 33977
rect 1027 33832 1036 33872
rect 1076 33832 5644 33872
rect 5684 33832 5693 33872
rect 3679 33307 4065 33326
rect 3679 33284 3745 33307
rect 3831 33284 3913 33307
rect 3999 33284 4065 33307
rect 3679 33244 3688 33284
rect 3728 33244 3745 33284
rect 3831 33244 3852 33284
rect 3892 33244 3913 33284
rect 3999 33244 4016 33284
rect 4056 33244 4065 33284
rect 3679 33221 3745 33244
rect 3831 33221 3913 33244
rect 3999 33221 4065 33244
rect 3679 33202 4065 33221
rect 18799 33307 19185 33326
rect 18799 33284 18865 33307
rect 18951 33284 19033 33307
rect 19119 33284 19185 33307
rect 18799 33244 18808 33284
rect 18848 33244 18865 33284
rect 18951 33244 18972 33284
rect 19012 33244 19033 33284
rect 19119 33244 19136 33284
rect 19176 33244 19185 33284
rect 18799 33221 18865 33244
rect 18951 33221 19033 33244
rect 19119 33221 19185 33244
rect 18799 33202 19185 33221
rect 6650 32803 6774 32822
rect 6650 32780 6669 32803
rect 5731 32740 5740 32780
rect 5780 32740 6669 32780
rect 6650 32717 6669 32740
rect 6755 32717 6774 32803
rect 6650 32698 6774 32717
rect 4919 32551 5305 32570
rect 4919 32528 4985 32551
rect 5071 32528 5153 32551
rect 5239 32528 5305 32551
rect 4919 32488 4928 32528
rect 4968 32488 4985 32528
rect 5071 32488 5092 32528
rect 5132 32488 5153 32528
rect 5239 32488 5256 32528
rect 5296 32488 5305 32528
rect 4919 32465 4985 32488
rect 5071 32465 5153 32488
rect 5239 32465 5305 32488
rect 4919 32446 5305 32465
rect 20039 32551 20425 32570
rect 20039 32528 20105 32551
rect 20191 32528 20273 32551
rect 20359 32528 20425 32551
rect 20039 32488 20048 32528
rect 20088 32488 20105 32528
rect 20191 32488 20212 32528
rect 20252 32488 20273 32528
rect 20359 32488 20376 32528
rect 20416 32488 20425 32528
rect 20039 32465 20105 32488
rect 20191 32465 20273 32488
rect 20359 32465 20425 32488
rect 20039 32446 20425 32465
rect 3679 31795 4065 31814
rect 3679 31772 3745 31795
rect 3831 31772 3913 31795
rect 3999 31772 4065 31795
rect 3679 31732 3688 31772
rect 3728 31732 3745 31772
rect 3831 31732 3852 31772
rect 3892 31732 3913 31772
rect 3999 31732 4016 31772
rect 4056 31732 4065 31772
rect 3679 31709 3745 31732
rect 3831 31709 3913 31732
rect 3999 31709 4065 31732
rect 3679 31690 4065 31709
rect 18799 31795 19185 31814
rect 18799 31772 18865 31795
rect 18951 31772 19033 31795
rect 19119 31772 19185 31795
rect 18799 31732 18808 31772
rect 18848 31732 18865 31772
rect 18951 31732 18972 31772
rect 19012 31732 19033 31772
rect 19119 31732 19136 31772
rect 19176 31732 19185 31772
rect 18799 31709 18865 31732
rect 18951 31709 19033 31732
rect 19119 31709 19185 31732
rect 18799 31690 19185 31709
rect 4919 31039 5305 31058
rect 4919 31016 4985 31039
rect 5071 31016 5153 31039
rect 5239 31016 5305 31039
rect 4919 30976 4928 31016
rect 4968 30976 4985 31016
rect 5071 30976 5092 31016
rect 5132 30976 5153 31016
rect 5239 30976 5256 31016
rect 5296 30976 5305 31016
rect 4919 30953 4985 30976
rect 5071 30953 5153 30976
rect 5239 30953 5305 30976
rect 4919 30934 5305 30953
rect 20039 31039 20425 31058
rect 20039 31016 20105 31039
rect 20191 31016 20273 31039
rect 20359 31016 20425 31039
rect 20039 30976 20048 31016
rect 20088 30976 20105 31016
rect 20191 30976 20212 31016
rect 20252 30976 20273 31016
rect 20359 30976 20376 31016
rect 20416 30976 20425 31016
rect 20039 30953 20105 30976
rect 20191 30953 20273 30976
rect 20359 30953 20425 30976
rect 20039 30934 20425 30953
rect 3679 30283 4065 30302
rect 3679 30260 3745 30283
rect 3831 30260 3913 30283
rect 3999 30260 4065 30283
rect 3679 30220 3688 30260
rect 3728 30220 3745 30260
rect 3831 30220 3852 30260
rect 3892 30220 3913 30260
rect 3999 30220 4016 30260
rect 4056 30220 4065 30260
rect 3679 30197 3745 30220
rect 3831 30197 3913 30220
rect 3999 30197 4065 30220
rect 3679 30178 4065 30197
rect 18799 30283 19185 30302
rect 18799 30260 18865 30283
rect 18951 30260 19033 30283
rect 19119 30260 19185 30283
rect 18799 30220 18808 30260
rect 18848 30220 18865 30260
rect 18951 30220 18972 30260
rect 19012 30220 19033 30260
rect 19119 30220 19136 30260
rect 19176 30220 19185 30260
rect 18799 30197 18865 30220
rect 18951 30197 19033 30220
rect 19119 30197 19185 30220
rect 18799 30178 19185 30197
rect 4919 29527 5305 29546
rect 4919 29504 4985 29527
rect 5071 29504 5153 29527
rect 5239 29504 5305 29527
rect 4919 29464 4928 29504
rect 4968 29464 4985 29504
rect 5071 29464 5092 29504
rect 5132 29464 5153 29504
rect 5239 29464 5256 29504
rect 5296 29464 5305 29504
rect 4919 29441 4985 29464
rect 5071 29441 5153 29464
rect 5239 29441 5305 29464
rect 4919 29422 5305 29441
rect 20039 29527 20425 29546
rect 20039 29504 20105 29527
rect 20191 29504 20273 29527
rect 20359 29504 20425 29527
rect 20039 29464 20048 29504
rect 20088 29464 20105 29504
rect 20191 29464 20212 29504
rect 20252 29464 20273 29504
rect 20359 29464 20376 29504
rect 20416 29464 20425 29504
rect 20039 29441 20105 29464
rect 20191 29441 20273 29464
rect 20359 29441 20425 29464
rect 20039 29422 20425 29441
rect 1507 28792 1516 28832
rect 1556 28792 1804 28832
rect 1844 28792 1853 28832
rect 3679 28771 4065 28790
rect 3679 28748 3745 28771
rect 3831 28748 3913 28771
rect 3999 28748 4065 28771
rect 3679 28708 3688 28748
rect 3728 28708 3745 28748
rect 3831 28708 3852 28748
rect 3892 28708 3913 28748
rect 3999 28708 4016 28748
rect 4056 28708 4065 28748
rect 3679 28685 3745 28708
rect 3831 28685 3913 28708
rect 3999 28685 4065 28708
rect 3679 28666 4065 28685
rect 18799 28771 19185 28790
rect 18799 28748 18865 28771
rect 18951 28748 19033 28771
rect 19119 28748 19185 28771
rect 18799 28708 18808 28748
rect 18848 28708 18865 28748
rect 18951 28708 18972 28748
rect 19012 28708 19033 28748
rect 19119 28708 19136 28748
rect 19176 28708 19185 28748
rect 18799 28685 18865 28708
rect 18951 28685 19033 28708
rect 19119 28685 19185 28708
rect 18799 28666 19185 28685
rect 4919 28015 5305 28034
rect 4919 27992 4985 28015
rect 5071 27992 5153 28015
rect 5239 27992 5305 28015
rect 4919 27952 4928 27992
rect 4968 27952 4985 27992
rect 5071 27952 5092 27992
rect 5132 27952 5153 27992
rect 5239 27952 5256 27992
rect 5296 27952 5305 27992
rect 4919 27929 4985 27952
rect 5071 27929 5153 27952
rect 5239 27929 5305 27952
rect 4919 27910 5305 27929
rect 20039 28015 20425 28034
rect 20039 27992 20105 28015
rect 20191 27992 20273 28015
rect 20359 27992 20425 28015
rect 20039 27952 20048 27992
rect 20088 27952 20105 27992
rect 20191 27952 20212 27992
rect 20252 27952 20273 27992
rect 20359 27952 20376 27992
rect 20416 27952 20425 27992
rect 20039 27929 20105 27952
rect 20191 27929 20273 27952
rect 20359 27929 20425 27952
rect 20039 27910 20425 27929
rect 3679 27259 4065 27278
rect 3679 27236 3745 27259
rect 3831 27236 3913 27259
rect 3999 27236 4065 27259
rect 3679 27196 3688 27236
rect 3728 27196 3745 27236
rect 3831 27196 3852 27236
rect 3892 27196 3913 27236
rect 3999 27196 4016 27236
rect 4056 27196 4065 27236
rect 3679 27173 3745 27196
rect 3831 27173 3913 27196
rect 3999 27173 4065 27196
rect 3679 27154 4065 27173
rect 18799 27259 19185 27278
rect 18799 27236 18865 27259
rect 18951 27236 19033 27259
rect 19119 27236 19185 27259
rect 18799 27196 18808 27236
rect 18848 27196 18865 27236
rect 18951 27196 18972 27236
rect 19012 27196 19033 27236
rect 19119 27196 19136 27236
rect 19176 27196 19185 27236
rect 18799 27173 18865 27196
rect 18951 27173 19033 27196
rect 19119 27173 19185 27196
rect 18799 27154 19185 27173
rect 4919 26503 5305 26522
rect 4919 26480 4985 26503
rect 5071 26480 5153 26503
rect 5239 26480 5305 26503
rect 4919 26440 4928 26480
rect 4968 26440 4985 26480
rect 5071 26440 5092 26480
rect 5132 26440 5153 26480
rect 5239 26440 5256 26480
rect 5296 26440 5305 26480
rect 4919 26417 4985 26440
rect 5071 26417 5153 26440
rect 5239 26417 5305 26440
rect 4919 26398 5305 26417
rect 20039 26503 20425 26522
rect 20039 26480 20105 26503
rect 20191 26480 20273 26503
rect 20359 26480 20425 26503
rect 20039 26440 20048 26480
rect 20088 26440 20105 26480
rect 20191 26440 20212 26480
rect 20252 26440 20273 26480
rect 20359 26440 20376 26480
rect 20416 26440 20425 26480
rect 20039 26417 20105 26440
rect 20191 26417 20273 26440
rect 20359 26417 20425 26440
rect 20039 26398 20425 26417
rect 3679 25747 4065 25766
rect 3679 25724 3745 25747
rect 3831 25724 3913 25747
rect 3999 25724 4065 25747
rect 3679 25684 3688 25724
rect 3728 25684 3745 25724
rect 3831 25684 3852 25724
rect 3892 25684 3913 25724
rect 3999 25684 4016 25724
rect 4056 25684 4065 25724
rect 3679 25661 3745 25684
rect 3831 25661 3913 25684
rect 3999 25661 4065 25684
rect 3679 25642 4065 25661
rect 18799 25747 19185 25766
rect 18799 25724 18865 25747
rect 18951 25724 19033 25747
rect 19119 25724 19185 25747
rect 18799 25684 18808 25724
rect 18848 25684 18865 25724
rect 18951 25684 18972 25724
rect 19012 25684 19033 25724
rect 19119 25684 19136 25724
rect 19176 25684 19185 25724
rect 18799 25661 18865 25684
rect 18951 25661 19033 25684
rect 19119 25661 19185 25684
rect 18799 25642 19185 25661
rect 2467 25180 2476 25220
rect 2516 25180 4012 25220
rect 4052 25180 4061 25220
rect 4919 24991 5305 25010
rect 4919 24968 4985 24991
rect 5071 24968 5153 24991
rect 5239 24968 5305 24991
rect 4919 24928 4928 24968
rect 4968 24928 4985 24968
rect 5071 24928 5092 24968
rect 5132 24928 5153 24968
rect 5239 24928 5256 24968
rect 5296 24928 5305 24968
rect 4919 24905 4985 24928
rect 5071 24905 5153 24928
rect 5239 24905 5305 24928
rect 4919 24886 5305 24905
rect 20039 24991 20425 25010
rect 20039 24968 20105 24991
rect 20191 24968 20273 24991
rect 20359 24968 20425 24991
rect 20039 24928 20048 24968
rect 20088 24928 20105 24968
rect 20191 24928 20212 24968
rect 20252 24928 20273 24968
rect 20359 24928 20376 24968
rect 20416 24928 20425 24968
rect 20039 24905 20105 24928
rect 20191 24905 20273 24928
rect 20359 24905 20425 24928
rect 20039 24886 20425 24905
rect 18403 24256 18412 24296
rect 18452 24256 18604 24296
rect 18644 24256 18653 24296
rect 3679 24235 4065 24254
rect 3679 24212 3745 24235
rect 3831 24212 3913 24235
rect 3999 24212 4065 24235
rect 3679 24172 3688 24212
rect 3728 24172 3745 24212
rect 3831 24172 3852 24212
rect 3892 24172 3913 24212
rect 3999 24172 4016 24212
rect 4056 24172 4065 24212
rect 3679 24149 3745 24172
rect 3831 24149 3913 24172
rect 3999 24149 4065 24172
rect 3679 24130 4065 24149
rect 18799 24235 19185 24254
rect 18799 24212 18865 24235
rect 18951 24212 19033 24235
rect 19119 24212 19185 24235
rect 18799 24172 18808 24212
rect 18848 24172 18865 24212
rect 18951 24172 18972 24212
rect 19012 24172 19033 24212
rect 19119 24172 19136 24212
rect 19176 24172 19185 24212
rect 18799 24149 18865 24172
rect 18951 24149 19033 24172
rect 19119 24149 19185 24172
rect 18799 24130 19185 24149
rect 4919 23479 5305 23498
rect 4919 23456 4985 23479
rect 5071 23456 5153 23479
rect 5239 23456 5305 23479
rect 4919 23416 4928 23456
rect 4968 23416 4985 23456
rect 5071 23416 5092 23456
rect 5132 23416 5153 23456
rect 5239 23416 5256 23456
rect 5296 23416 5305 23456
rect 4919 23393 4985 23416
rect 5071 23393 5153 23416
rect 5239 23393 5305 23416
rect 4919 23374 5305 23393
rect 20039 23479 20425 23498
rect 20039 23456 20105 23479
rect 20191 23456 20273 23479
rect 20359 23456 20425 23479
rect 20039 23416 20048 23456
rect 20088 23416 20105 23456
rect 20191 23416 20212 23456
rect 20252 23416 20273 23456
rect 20359 23416 20376 23456
rect 20416 23416 20425 23456
rect 20039 23393 20105 23416
rect 20191 23393 20273 23416
rect 20359 23393 20425 23416
rect 20039 23374 20425 23393
rect 3679 22723 4065 22742
rect 3679 22700 3745 22723
rect 3831 22700 3913 22723
rect 3999 22700 4065 22723
rect 3679 22660 3688 22700
rect 3728 22660 3745 22700
rect 3831 22660 3852 22700
rect 3892 22660 3913 22700
rect 3999 22660 4016 22700
rect 4056 22660 4065 22700
rect 3679 22637 3745 22660
rect 3831 22637 3913 22660
rect 3999 22637 4065 22660
rect 3679 22618 4065 22637
rect 18799 22723 19185 22742
rect 18799 22700 18865 22723
rect 18951 22700 19033 22723
rect 19119 22700 19185 22723
rect 18799 22660 18808 22700
rect 18848 22660 18865 22700
rect 18951 22660 18972 22700
rect 19012 22660 19033 22700
rect 19119 22660 19136 22700
rect 19176 22660 19185 22700
rect 18799 22637 18865 22660
rect 18951 22637 19033 22660
rect 19119 22637 19185 22660
rect 18799 22618 19185 22637
rect 4919 21967 5305 21986
rect 4919 21944 4985 21967
rect 5071 21944 5153 21967
rect 5239 21944 5305 21967
rect 4919 21904 4928 21944
rect 4968 21904 4985 21944
rect 5071 21904 5092 21944
rect 5132 21904 5153 21944
rect 5239 21904 5256 21944
rect 5296 21904 5305 21944
rect 4919 21881 4985 21904
rect 5071 21881 5153 21904
rect 5239 21881 5305 21904
rect 4919 21862 5305 21881
rect 20039 21967 20425 21986
rect 20039 21944 20105 21967
rect 20191 21944 20273 21967
rect 20359 21944 20425 21967
rect 20039 21904 20048 21944
rect 20088 21904 20105 21944
rect 20191 21904 20212 21944
rect 20252 21904 20273 21944
rect 20359 21904 20376 21944
rect 20416 21904 20425 21944
rect 20039 21881 20105 21904
rect 20191 21881 20273 21904
rect 20359 21881 20425 21904
rect 20039 21862 20425 21881
rect 3679 21211 4065 21230
rect 3679 21188 3745 21211
rect 3831 21188 3913 21211
rect 3999 21188 4065 21211
rect 3679 21148 3688 21188
rect 3728 21148 3745 21188
rect 3831 21148 3852 21188
rect 3892 21148 3913 21188
rect 3999 21148 4016 21188
rect 4056 21148 4065 21188
rect 3679 21125 3745 21148
rect 3831 21125 3913 21148
rect 3999 21125 4065 21148
rect 3679 21106 4065 21125
rect 18799 21211 19185 21230
rect 18799 21188 18865 21211
rect 18951 21188 19033 21211
rect 19119 21188 19185 21211
rect 18799 21148 18808 21188
rect 18848 21148 18865 21188
rect 18951 21148 18972 21188
rect 19012 21148 19033 21188
rect 19119 21148 19136 21188
rect 19176 21148 19185 21188
rect 18799 21125 18865 21148
rect 18951 21125 19033 21148
rect 19119 21125 19185 21148
rect 18799 21106 19185 21125
rect 4919 20455 5305 20474
rect 4919 20432 4985 20455
rect 5071 20432 5153 20455
rect 5239 20432 5305 20455
rect 4919 20392 4928 20432
rect 4968 20392 4985 20432
rect 5071 20392 5092 20432
rect 5132 20392 5153 20432
rect 5239 20392 5256 20432
rect 5296 20392 5305 20432
rect 4919 20369 4985 20392
rect 5071 20369 5153 20392
rect 5239 20369 5305 20392
rect 4919 20350 5305 20369
rect 20039 20455 20425 20474
rect 20039 20432 20105 20455
rect 20191 20432 20273 20455
rect 20359 20432 20425 20455
rect 20039 20392 20048 20432
rect 20088 20392 20105 20432
rect 20191 20392 20212 20432
rect 20252 20392 20273 20432
rect 20359 20392 20376 20432
rect 20416 20392 20425 20432
rect 20039 20369 20105 20392
rect 20191 20369 20273 20392
rect 20359 20369 20425 20392
rect 20039 20350 20425 20369
rect 3679 19699 4065 19718
rect 3679 19676 3745 19699
rect 3831 19676 3913 19699
rect 3999 19676 4065 19699
rect 3679 19636 3688 19676
rect 3728 19636 3745 19676
rect 3831 19636 3852 19676
rect 3892 19636 3913 19676
rect 3999 19636 4016 19676
rect 4056 19636 4065 19676
rect 3679 19613 3745 19636
rect 3831 19613 3913 19636
rect 3999 19613 4065 19636
rect 3679 19594 4065 19613
rect 18799 19699 19185 19718
rect 18799 19676 18865 19699
rect 18951 19676 19033 19699
rect 19119 19676 19185 19699
rect 18799 19636 18808 19676
rect 18848 19636 18865 19676
rect 18951 19636 18972 19676
rect 19012 19636 19033 19676
rect 19119 19636 19136 19676
rect 19176 19636 19185 19676
rect 18799 19613 18865 19636
rect 18951 19613 19033 19636
rect 19119 19613 19185 19636
rect 18799 19594 19185 19613
rect 1603 19216 1612 19256
rect 1652 19216 3436 19256
rect 3476 19216 5548 19256
rect 5588 19216 5597 19256
rect 4919 18943 5305 18962
rect 4919 18920 4985 18943
rect 5071 18920 5153 18943
rect 5239 18920 5305 18943
rect 4919 18880 4928 18920
rect 4968 18880 4985 18920
rect 5071 18880 5092 18920
rect 5132 18880 5153 18920
rect 5239 18880 5256 18920
rect 5296 18880 5305 18920
rect 4919 18857 4985 18880
rect 5071 18857 5153 18880
rect 5239 18857 5305 18880
rect 4919 18838 5305 18857
rect 20039 18943 20425 18962
rect 20039 18920 20105 18943
rect 20191 18920 20273 18943
rect 20359 18920 20425 18943
rect 20039 18880 20048 18920
rect 20088 18880 20105 18920
rect 20191 18880 20212 18920
rect 20252 18880 20273 18920
rect 20359 18880 20376 18920
rect 20416 18880 20425 18920
rect 20039 18857 20105 18880
rect 20191 18857 20273 18880
rect 20359 18857 20425 18880
rect 20039 18838 20425 18857
rect 11107 18292 11116 18332
rect 11156 18292 20908 18332
rect 20948 18292 20957 18332
rect 3679 18187 4065 18206
rect 3679 18164 3745 18187
rect 3831 18164 3913 18187
rect 3999 18164 4065 18187
rect 3679 18124 3688 18164
rect 3728 18124 3745 18164
rect 3831 18124 3852 18164
rect 3892 18124 3913 18164
rect 3999 18124 4016 18164
rect 4056 18124 4065 18164
rect 3679 18101 3745 18124
rect 3831 18101 3913 18124
rect 3999 18101 4065 18124
rect 3679 18082 4065 18101
rect 18799 18187 19185 18206
rect 18799 18164 18865 18187
rect 18951 18164 19033 18187
rect 19119 18164 19185 18187
rect 18799 18124 18808 18164
rect 18848 18124 18865 18164
rect 18951 18124 18972 18164
rect 19012 18124 19033 18164
rect 19119 18124 19136 18164
rect 19176 18124 19185 18164
rect 18799 18101 18865 18124
rect 18951 18101 19033 18124
rect 19119 18101 19185 18124
rect 18799 18082 19185 18101
rect 2371 17704 2380 17744
rect 2420 17704 10156 17744
rect 10196 17704 10205 17744
rect 4919 17431 5305 17450
rect 4919 17408 4985 17431
rect 5071 17408 5153 17431
rect 5239 17408 5305 17431
rect 4919 17368 4928 17408
rect 4968 17368 4985 17408
rect 5071 17368 5092 17408
rect 5132 17368 5153 17408
rect 5239 17368 5256 17408
rect 5296 17368 5305 17408
rect 4919 17345 4985 17368
rect 5071 17345 5153 17368
rect 5239 17345 5305 17368
rect 4919 17326 5305 17345
rect 20039 17431 20425 17450
rect 20039 17408 20105 17431
rect 20191 17408 20273 17431
rect 20359 17408 20425 17431
rect 20039 17368 20048 17408
rect 20088 17368 20105 17408
rect 20191 17368 20212 17408
rect 20252 17368 20273 17408
rect 20359 17368 20376 17408
rect 20416 17368 20425 17408
rect 20039 17345 20105 17368
rect 20191 17345 20273 17368
rect 20359 17345 20425 17368
rect 20039 17326 20425 17345
rect 3679 16675 4065 16694
rect 3679 16652 3745 16675
rect 3831 16652 3913 16675
rect 3999 16652 4065 16675
rect 3679 16612 3688 16652
rect 3728 16612 3745 16652
rect 3831 16612 3852 16652
rect 3892 16612 3913 16652
rect 3999 16612 4016 16652
rect 4056 16612 4065 16652
rect 3679 16589 3745 16612
rect 3831 16589 3913 16612
rect 3999 16589 4065 16612
rect 3679 16570 4065 16589
rect 18799 16675 19185 16694
rect 18799 16652 18865 16675
rect 18951 16652 19033 16675
rect 19119 16652 19185 16675
rect 18799 16612 18808 16652
rect 18848 16612 18865 16652
rect 18951 16612 18972 16652
rect 19012 16612 19033 16652
rect 19119 16612 19136 16652
rect 19176 16612 19185 16652
rect 18799 16589 18865 16612
rect 18951 16589 19033 16612
rect 19119 16589 19185 16612
rect 18799 16570 19185 16589
rect 4919 15919 5305 15938
rect 4919 15896 4985 15919
rect 5071 15896 5153 15919
rect 5239 15896 5305 15919
rect 4919 15856 4928 15896
rect 4968 15856 4985 15896
rect 5071 15856 5092 15896
rect 5132 15856 5153 15896
rect 5239 15856 5256 15896
rect 5296 15856 5305 15896
rect 4919 15833 4985 15856
rect 5071 15833 5153 15856
rect 5239 15833 5305 15856
rect 4919 15814 5305 15833
rect 20039 15919 20425 15938
rect 20039 15896 20105 15919
rect 20191 15896 20273 15919
rect 20359 15896 20425 15919
rect 20039 15856 20048 15896
rect 20088 15856 20105 15896
rect 20191 15856 20212 15896
rect 20252 15856 20273 15896
rect 20359 15856 20376 15896
rect 20416 15856 20425 15896
rect 20039 15833 20105 15856
rect 20191 15833 20273 15856
rect 20359 15833 20425 15856
rect 20039 15814 20425 15833
rect 3679 15163 4065 15182
rect 3679 15140 3745 15163
rect 3831 15140 3913 15163
rect 3999 15140 4065 15163
rect 3679 15100 3688 15140
rect 3728 15100 3745 15140
rect 3831 15100 3852 15140
rect 3892 15100 3913 15140
rect 3999 15100 4016 15140
rect 4056 15100 4065 15140
rect 3679 15077 3745 15100
rect 3831 15077 3913 15100
rect 3999 15077 4065 15100
rect 3679 15058 4065 15077
rect 18799 15163 19185 15182
rect 18799 15140 18865 15163
rect 18951 15140 19033 15163
rect 19119 15140 19185 15163
rect 18799 15100 18808 15140
rect 18848 15100 18865 15140
rect 18951 15100 18972 15140
rect 19012 15100 19033 15140
rect 19119 15100 19136 15140
rect 19176 15100 19185 15140
rect 18799 15077 18865 15100
rect 18951 15077 19033 15100
rect 19119 15077 19185 15100
rect 18799 15058 19185 15077
rect 4919 14407 5305 14426
rect 4919 14384 4985 14407
rect 5071 14384 5153 14407
rect 5239 14384 5305 14407
rect 4919 14344 4928 14384
rect 4968 14344 4985 14384
rect 5071 14344 5092 14384
rect 5132 14344 5153 14384
rect 5239 14344 5256 14384
rect 5296 14344 5305 14384
rect 4919 14321 4985 14344
rect 5071 14321 5153 14344
rect 5239 14321 5305 14344
rect 4919 14302 5305 14321
rect 20039 14407 20425 14426
rect 20039 14384 20105 14407
rect 20191 14384 20273 14407
rect 20359 14384 20425 14407
rect 20039 14344 20048 14384
rect 20088 14344 20105 14384
rect 20191 14344 20212 14384
rect 20252 14344 20273 14384
rect 20359 14344 20376 14384
rect 20416 14344 20425 14384
rect 20039 14321 20105 14344
rect 20191 14321 20273 14344
rect 20359 14321 20425 14344
rect 20039 14302 20425 14321
rect 3679 13651 4065 13670
rect 3679 13628 3745 13651
rect 3831 13628 3913 13651
rect 3999 13628 4065 13651
rect 3679 13588 3688 13628
rect 3728 13588 3745 13628
rect 3831 13588 3852 13628
rect 3892 13588 3913 13628
rect 3999 13588 4016 13628
rect 4056 13588 4065 13628
rect 3679 13565 3745 13588
rect 3831 13565 3913 13588
rect 3999 13565 4065 13588
rect 3679 13546 4065 13565
rect 18799 13651 19185 13670
rect 18799 13628 18865 13651
rect 18951 13628 19033 13651
rect 19119 13628 19185 13651
rect 18799 13588 18808 13628
rect 18848 13588 18865 13628
rect 18951 13588 18972 13628
rect 19012 13588 19033 13628
rect 19119 13588 19136 13628
rect 19176 13588 19185 13628
rect 18799 13565 18865 13588
rect 18951 13565 19033 13588
rect 19119 13565 19185 13588
rect 18799 13546 19185 13565
rect 4919 12895 5305 12914
rect 4919 12872 4985 12895
rect 5071 12872 5153 12895
rect 5239 12872 5305 12895
rect 4919 12832 4928 12872
rect 4968 12832 4985 12872
rect 5071 12832 5092 12872
rect 5132 12832 5153 12872
rect 5239 12832 5256 12872
rect 5296 12832 5305 12872
rect 4919 12809 4985 12832
rect 5071 12809 5153 12832
rect 5239 12809 5305 12832
rect 4919 12790 5305 12809
rect 20039 12895 20425 12914
rect 20039 12872 20105 12895
rect 20191 12872 20273 12895
rect 20359 12872 20425 12895
rect 20039 12832 20048 12872
rect 20088 12832 20105 12872
rect 20191 12832 20212 12872
rect 20252 12832 20273 12872
rect 20359 12832 20376 12872
rect 20416 12832 20425 12872
rect 20039 12809 20105 12832
rect 20191 12809 20273 12832
rect 20359 12809 20425 12832
rect 20039 12790 20425 12809
rect 3679 12139 4065 12158
rect 3679 12116 3745 12139
rect 3831 12116 3913 12139
rect 3999 12116 4065 12139
rect 3679 12076 3688 12116
rect 3728 12076 3745 12116
rect 3831 12076 3852 12116
rect 3892 12076 3913 12116
rect 3999 12076 4016 12116
rect 4056 12076 4065 12116
rect 3679 12053 3745 12076
rect 3831 12053 3913 12076
rect 3999 12053 4065 12076
rect 3679 12034 4065 12053
rect 18799 12139 19185 12158
rect 18799 12116 18865 12139
rect 18951 12116 19033 12139
rect 19119 12116 19185 12139
rect 18799 12076 18808 12116
rect 18848 12076 18865 12116
rect 18951 12076 18972 12116
rect 19012 12076 19033 12116
rect 19119 12076 19136 12116
rect 19176 12076 19185 12116
rect 18799 12053 18865 12076
rect 18951 12053 19033 12076
rect 19119 12053 19185 12076
rect 18799 12034 19185 12053
rect 4919 11383 5305 11402
rect 4919 11360 4985 11383
rect 5071 11360 5153 11383
rect 5239 11360 5305 11383
rect 4919 11320 4928 11360
rect 4968 11320 4985 11360
rect 5071 11320 5092 11360
rect 5132 11320 5153 11360
rect 5239 11320 5256 11360
rect 5296 11320 5305 11360
rect 4919 11297 4985 11320
rect 5071 11297 5153 11320
rect 5239 11297 5305 11320
rect 4919 11278 5305 11297
rect 20039 11383 20425 11402
rect 20039 11360 20105 11383
rect 20191 11360 20273 11383
rect 20359 11360 20425 11383
rect 20039 11320 20048 11360
rect 20088 11320 20105 11360
rect 20191 11320 20212 11360
rect 20252 11320 20273 11360
rect 20359 11320 20376 11360
rect 20416 11320 20425 11360
rect 20039 11297 20105 11320
rect 20191 11297 20273 11320
rect 20359 11297 20425 11320
rect 20039 11278 20425 11297
rect 3679 10627 4065 10646
rect 3679 10604 3745 10627
rect 3831 10604 3913 10627
rect 3999 10604 4065 10627
rect 3679 10564 3688 10604
rect 3728 10564 3745 10604
rect 3831 10564 3852 10604
rect 3892 10564 3913 10604
rect 3999 10564 4016 10604
rect 4056 10564 4065 10604
rect 3679 10541 3745 10564
rect 3831 10541 3913 10564
rect 3999 10541 4065 10564
rect 3679 10522 4065 10541
rect 18799 10627 19185 10646
rect 18799 10604 18865 10627
rect 18951 10604 19033 10627
rect 19119 10604 19185 10627
rect 18799 10564 18808 10604
rect 18848 10564 18865 10604
rect 18951 10564 18972 10604
rect 19012 10564 19033 10604
rect 19119 10564 19136 10604
rect 19176 10564 19185 10604
rect 18799 10541 18865 10564
rect 18951 10541 19033 10564
rect 19119 10541 19185 10564
rect 18799 10522 19185 10541
rect 4919 9871 5305 9890
rect 4919 9848 4985 9871
rect 5071 9848 5153 9871
rect 5239 9848 5305 9871
rect 4919 9808 4928 9848
rect 4968 9808 4985 9848
rect 5071 9808 5092 9848
rect 5132 9808 5153 9848
rect 5239 9808 5256 9848
rect 5296 9808 5305 9848
rect 4919 9785 4985 9808
rect 5071 9785 5153 9808
rect 5239 9785 5305 9808
rect 4919 9766 5305 9785
rect 20039 9871 20425 9890
rect 20039 9848 20105 9871
rect 20191 9848 20273 9871
rect 20359 9848 20425 9871
rect 20039 9808 20048 9848
rect 20088 9808 20105 9848
rect 20191 9808 20212 9848
rect 20252 9808 20273 9848
rect 20359 9808 20376 9848
rect 20416 9808 20425 9848
rect 20039 9785 20105 9808
rect 20191 9785 20273 9808
rect 20359 9785 20425 9808
rect 20039 9766 20425 9785
rect 3679 9115 4065 9134
rect 3679 9092 3745 9115
rect 3831 9092 3913 9115
rect 3999 9092 4065 9115
rect 3679 9052 3688 9092
rect 3728 9052 3745 9092
rect 3831 9052 3852 9092
rect 3892 9052 3913 9092
rect 3999 9052 4016 9092
rect 4056 9052 4065 9092
rect 3679 9029 3745 9052
rect 3831 9029 3913 9052
rect 3999 9029 4065 9052
rect 3679 9010 4065 9029
rect 18799 9115 19185 9134
rect 18799 9092 18865 9115
rect 18951 9092 19033 9115
rect 19119 9092 19185 9115
rect 18799 9052 18808 9092
rect 18848 9052 18865 9092
rect 18951 9052 18972 9092
rect 19012 9052 19033 9092
rect 19119 9052 19136 9092
rect 19176 9052 19185 9092
rect 18799 9029 18865 9052
rect 18951 9029 19033 9052
rect 19119 9029 19185 9052
rect 18799 9010 19185 9029
rect 4919 8359 5305 8378
rect 4919 8336 4985 8359
rect 5071 8336 5153 8359
rect 5239 8336 5305 8359
rect 4919 8296 4928 8336
rect 4968 8296 4985 8336
rect 5071 8296 5092 8336
rect 5132 8296 5153 8336
rect 5239 8296 5256 8336
rect 5296 8296 5305 8336
rect 4919 8273 4985 8296
rect 5071 8273 5153 8296
rect 5239 8273 5305 8296
rect 4919 8254 5305 8273
rect 20039 8359 20425 8378
rect 20039 8336 20105 8359
rect 20191 8336 20273 8359
rect 20359 8336 20425 8359
rect 20039 8296 20048 8336
rect 20088 8296 20105 8336
rect 20191 8296 20212 8336
rect 20252 8296 20273 8336
rect 20359 8296 20376 8336
rect 20416 8296 20425 8336
rect 20039 8273 20105 8296
rect 20191 8273 20273 8296
rect 20359 8273 20425 8296
rect 20039 8254 20425 8273
rect 3679 7603 4065 7622
rect 3679 7580 3745 7603
rect 3831 7580 3913 7603
rect 3999 7580 4065 7603
rect 3679 7540 3688 7580
rect 3728 7540 3745 7580
rect 3831 7540 3852 7580
rect 3892 7540 3913 7580
rect 3999 7540 4016 7580
rect 4056 7540 4065 7580
rect 3679 7517 3745 7540
rect 3831 7517 3913 7540
rect 3999 7517 4065 7540
rect 3679 7498 4065 7517
rect 18799 7603 19185 7622
rect 18799 7580 18865 7603
rect 18951 7580 19033 7603
rect 19119 7580 19185 7603
rect 18799 7540 18808 7580
rect 18848 7540 18865 7580
rect 18951 7540 18972 7580
rect 19012 7540 19033 7580
rect 19119 7540 19136 7580
rect 19176 7540 19185 7580
rect 18799 7517 18865 7540
rect 18951 7517 19033 7540
rect 19119 7517 19185 7540
rect 18799 7498 19185 7517
rect 4919 6847 5305 6866
rect 4919 6824 4985 6847
rect 5071 6824 5153 6847
rect 5239 6824 5305 6847
rect 4919 6784 4928 6824
rect 4968 6784 4985 6824
rect 5071 6784 5092 6824
rect 5132 6784 5153 6824
rect 5239 6784 5256 6824
rect 5296 6784 5305 6824
rect 4919 6761 4985 6784
rect 5071 6761 5153 6784
rect 5239 6761 5305 6784
rect 4919 6742 5305 6761
rect 20039 6847 20425 6866
rect 20039 6824 20105 6847
rect 20191 6824 20273 6847
rect 20359 6824 20425 6847
rect 20039 6784 20048 6824
rect 20088 6784 20105 6824
rect 20191 6784 20212 6824
rect 20252 6784 20273 6824
rect 20359 6784 20376 6824
rect 20416 6784 20425 6824
rect 20039 6761 20105 6784
rect 20191 6761 20273 6784
rect 20359 6761 20425 6784
rect 20039 6742 20425 6761
rect 4387 6280 4396 6320
rect 4436 6280 19948 6320
rect 19988 6280 19997 6320
rect 3679 6091 4065 6110
rect 3679 6068 3745 6091
rect 3831 6068 3913 6091
rect 3999 6068 4065 6091
rect 3679 6028 3688 6068
rect 3728 6028 3745 6068
rect 3831 6028 3852 6068
rect 3892 6028 3913 6068
rect 3999 6028 4016 6068
rect 4056 6028 4065 6068
rect 3679 6005 3745 6028
rect 3831 6005 3913 6028
rect 3999 6005 4065 6028
rect 3679 5986 4065 6005
rect 18799 6091 19185 6110
rect 18799 6068 18865 6091
rect 18951 6068 19033 6091
rect 19119 6068 19185 6091
rect 18799 6028 18808 6068
rect 18848 6028 18865 6068
rect 18951 6028 18972 6068
rect 19012 6028 19033 6068
rect 19119 6028 19136 6068
rect 19176 6028 19185 6068
rect 18799 6005 18865 6028
rect 18951 6005 19033 6028
rect 19119 6005 19185 6028
rect 18799 5986 19185 6005
rect 4919 5335 5305 5354
rect 4919 5312 4985 5335
rect 5071 5312 5153 5335
rect 5239 5312 5305 5335
rect 4919 5272 4928 5312
rect 4968 5272 4985 5312
rect 5071 5272 5092 5312
rect 5132 5272 5153 5312
rect 5239 5272 5256 5312
rect 5296 5272 5305 5312
rect 4919 5249 4985 5272
rect 5071 5249 5153 5272
rect 5239 5249 5305 5272
rect 4919 5230 5305 5249
rect 20039 5335 20425 5354
rect 20039 5312 20105 5335
rect 20191 5312 20273 5335
rect 20359 5312 20425 5335
rect 20039 5272 20048 5312
rect 20088 5272 20105 5312
rect 20191 5272 20212 5312
rect 20252 5272 20273 5312
rect 20359 5272 20376 5312
rect 20416 5272 20425 5312
rect 20039 5249 20105 5272
rect 20191 5249 20273 5272
rect 20359 5249 20425 5272
rect 20039 5230 20425 5249
rect 3679 4579 4065 4598
rect 3679 4556 3745 4579
rect 3831 4556 3913 4579
rect 3999 4556 4065 4579
rect 3679 4516 3688 4556
rect 3728 4516 3745 4556
rect 3831 4516 3852 4556
rect 3892 4516 3913 4556
rect 3999 4516 4016 4556
rect 4056 4516 4065 4556
rect 3679 4493 3745 4516
rect 3831 4493 3913 4516
rect 3999 4493 4065 4516
rect 3679 4474 4065 4493
rect 18799 4579 19185 4598
rect 18799 4556 18865 4579
rect 18951 4556 19033 4579
rect 19119 4556 19185 4579
rect 18799 4516 18808 4556
rect 18848 4516 18865 4556
rect 18951 4516 18972 4556
rect 19012 4516 19033 4556
rect 19119 4516 19136 4556
rect 19176 4516 19185 4556
rect 18799 4493 18865 4516
rect 18951 4493 19033 4516
rect 19119 4493 19185 4516
rect 18799 4474 19185 4493
rect 4919 3823 5305 3842
rect 4919 3800 4985 3823
rect 5071 3800 5153 3823
rect 5239 3800 5305 3823
rect 4919 3760 4928 3800
rect 4968 3760 4985 3800
rect 5071 3760 5092 3800
rect 5132 3760 5153 3800
rect 5239 3760 5256 3800
rect 5296 3760 5305 3800
rect 4919 3737 4985 3760
rect 5071 3737 5153 3760
rect 5239 3737 5305 3760
rect 4919 3718 5305 3737
rect 20039 3823 20425 3842
rect 20039 3800 20105 3823
rect 20191 3800 20273 3823
rect 20359 3800 20425 3823
rect 20039 3760 20048 3800
rect 20088 3760 20105 3800
rect 20191 3760 20212 3800
rect 20252 3760 20273 3800
rect 20359 3760 20376 3800
rect 20416 3760 20425 3800
rect 20039 3737 20105 3760
rect 20191 3737 20273 3760
rect 20359 3737 20425 3760
rect 20039 3718 20425 3737
rect 3679 3067 4065 3086
rect 3679 3044 3745 3067
rect 3831 3044 3913 3067
rect 3999 3044 4065 3067
rect 3679 3004 3688 3044
rect 3728 3004 3745 3044
rect 3831 3004 3852 3044
rect 3892 3004 3913 3044
rect 3999 3004 4016 3044
rect 4056 3004 4065 3044
rect 3679 2981 3745 3004
rect 3831 2981 3913 3004
rect 3999 2981 4065 3004
rect 3679 2962 4065 2981
rect 18799 3067 19185 3086
rect 18799 3044 18865 3067
rect 18951 3044 19033 3067
rect 19119 3044 19185 3067
rect 18799 3004 18808 3044
rect 18848 3004 18865 3044
rect 18951 3004 18972 3044
rect 19012 3004 19033 3044
rect 19119 3004 19136 3044
rect 19176 3004 19185 3044
rect 18799 2981 18865 3004
rect 18951 2981 19033 3004
rect 19119 2981 19185 3004
rect 18799 2962 19185 2981
rect 4919 2311 5305 2330
rect 4919 2288 4985 2311
rect 5071 2288 5153 2311
rect 5239 2288 5305 2311
rect 4919 2248 4928 2288
rect 4968 2248 4985 2288
rect 5071 2248 5092 2288
rect 5132 2248 5153 2288
rect 5239 2248 5256 2288
rect 5296 2248 5305 2288
rect 4919 2225 4985 2248
rect 5071 2225 5153 2248
rect 5239 2225 5305 2248
rect 4919 2206 5305 2225
rect 20039 2311 20425 2330
rect 20039 2288 20105 2311
rect 20191 2288 20273 2311
rect 20359 2288 20425 2311
rect 20039 2248 20048 2288
rect 20088 2248 20105 2288
rect 20191 2248 20212 2288
rect 20252 2248 20273 2288
rect 20359 2248 20376 2288
rect 20416 2248 20425 2288
rect 20039 2225 20105 2248
rect 20191 2225 20273 2248
rect 20359 2225 20425 2248
rect 20039 2206 20425 2225
rect 3679 1555 4065 1574
rect 3679 1532 3745 1555
rect 3831 1532 3913 1555
rect 3999 1532 4065 1555
rect 3679 1492 3688 1532
rect 3728 1492 3745 1532
rect 3831 1492 3852 1532
rect 3892 1492 3913 1532
rect 3999 1492 4016 1532
rect 4056 1492 4065 1532
rect 3679 1469 3745 1492
rect 3831 1469 3913 1492
rect 3999 1469 4065 1492
rect 3679 1450 4065 1469
rect 18799 1555 19185 1574
rect 18799 1532 18865 1555
rect 18951 1532 19033 1555
rect 19119 1532 19185 1555
rect 18799 1492 18808 1532
rect 18848 1492 18865 1532
rect 18951 1492 18972 1532
rect 19012 1492 19033 1532
rect 19119 1492 19136 1532
rect 19176 1492 19185 1532
rect 18799 1469 18865 1492
rect 18951 1469 19033 1492
rect 19119 1469 19185 1492
rect 18799 1450 19185 1469
rect 2179 1240 2188 1280
rect 2228 1240 3148 1280
rect 3188 1240 3197 1280
rect 6650 967 6774 986
rect 6650 944 6669 967
rect 6595 904 6604 944
rect 6644 904 6669 944
rect 6650 881 6669 904
rect 6755 881 6774 967
rect 6650 862 6774 881
rect 4919 799 5305 818
rect 4919 776 4985 799
rect 5071 776 5153 799
rect 5239 776 5305 799
rect 4919 736 4928 776
rect 4968 736 4985 776
rect 5071 736 5092 776
rect 5132 736 5153 776
rect 5239 736 5256 776
rect 5296 736 5305 776
rect 4919 713 4985 736
rect 5071 713 5153 736
rect 5239 713 5305 736
rect 4919 694 5305 713
rect 20039 799 20425 818
rect 20039 776 20105 799
rect 20191 776 20273 799
rect 20359 776 20425 799
rect 20039 736 20048 776
rect 20088 736 20105 776
rect 20191 736 20212 776
rect 20252 736 20273 776
rect 20359 736 20376 776
rect 20416 736 20425 776
rect 20039 713 20105 736
rect 20191 713 20273 736
rect 20359 713 20425 736
rect 20039 694 20425 713
rect 5251 232 5260 272
rect 5300 232 8428 272
rect 8468 232 8477 272
<< via5 >>
rect 4985 41600 5071 41623
rect 5153 41600 5239 41623
rect 4985 41560 5010 41600
rect 5010 41560 5050 41600
rect 5050 41560 5071 41600
rect 5153 41560 5174 41600
rect 5174 41560 5214 41600
rect 5214 41560 5239 41600
rect 4985 41537 5071 41560
rect 5153 41537 5239 41560
rect 20105 41600 20191 41623
rect 20273 41600 20359 41623
rect 20105 41560 20130 41600
rect 20130 41560 20170 41600
rect 20170 41560 20191 41600
rect 20273 41560 20294 41600
rect 20294 41560 20334 41600
rect 20334 41560 20359 41600
rect 20105 41537 20191 41560
rect 20273 41537 20359 41560
rect 3745 40844 3831 40867
rect 3913 40844 3999 40867
rect 3745 40804 3770 40844
rect 3770 40804 3810 40844
rect 3810 40804 3831 40844
rect 3913 40804 3934 40844
rect 3934 40804 3974 40844
rect 3974 40804 3999 40844
rect 3745 40781 3831 40804
rect 3913 40781 3999 40804
rect 18865 40844 18951 40867
rect 19033 40844 19119 40867
rect 18865 40804 18890 40844
rect 18890 40804 18930 40844
rect 18930 40804 18951 40844
rect 19033 40804 19054 40844
rect 19054 40804 19094 40844
rect 19094 40804 19119 40844
rect 18865 40781 18951 40804
rect 19033 40781 19119 40804
rect 4985 40088 5071 40111
rect 5153 40088 5239 40111
rect 4985 40048 5010 40088
rect 5010 40048 5050 40088
rect 5050 40048 5071 40088
rect 5153 40048 5174 40088
rect 5174 40048 5214 40088
rect 5214 40048 5239 40088
rect 4985 40025 5071 40048
rect 5153 40025 5239 40048
rect 20105 40088 20191 40111
rect 20273 40088 20359 40111
rect 20105 40048 20130 40088
rect 20130 40048 20170 40088
rect 20170 40048 20191 40088
rect 20273 40048 20294 40088
rect 20294 40048 20334 40088
rect 20334 40048 20359 40088
rect 20105 40025 20191 40048
rect 20273 40025 20359 40048
rect 3745 39332 3831 39355
rect 3913 39332 3999 39355
rect 3745 39292 3770 39332
rect 3770 39292 3810 39332
rect 3810 39292 3831 39332
rect 3913 39292 3934 39332
rect 3934 39292 3974 39332
rect 3974 39292 3999 39332
rect 3745 39269 3831 39292
rect 3913 39269 3999 39292
rect 18865 39332 18951 39355
rect 19033 39332 19119 39355
rect 18865 39292 18890 39332
rect 18890 39292 18930 39332
rect 18930 39292 18951 39332
rect 19033 39292 19054 39332
rect 19054 39292 19094 39332
rect 19094 39292 19119 39332
rect 18865 39269 18951 39292
rect 19033 39269 19119 39292
rect 4985 38576 5071 38599
rect 5153 38576 5239 38599
rect 4985 38536 5010 38576
rect 5010 38536 5050 38576
rect 5050 38536 5071 38576
rect 5153 38536 5174 38576
rect 5174 38536 5214 38576
rect 5214 38536 5239 38576
rect 4985 38513 5071 38536
rect 5153 38513 5239 38536
rect 20105 38576 20191 38599
rect 20273 38576 20359 38599
rect 20105 38536 20130 38576
rect 20130 38536 20170 38576
rect 20170 38536 20191 38576
rect 20273 38536 20294 38576
rect 20294 38536 20334 38576
rect 20334 38536 20359 38576
rect 20105 38513 20191 38536
rect 20273 38513 20359 38536
rect 3745 37820 3831 37843
rect 3913 37820 3999 37843
rect 3745 37780 3770 37820
rect 3770 37780 3810 37820
rect 3810 37780 3831 37820
rect 3913 37780 3934 37820
rect 3934 37780 3974 37820
rect 3974 37780 3999 37820
rect 3745 37757 3831 37780
rect 3913 37757 3999 37780
rect 18865 37820 18951 37843
rect 19033 37820 19119 37843
rect 18865 37780 18890 37820
rect 18890 37780 18930 37820
rect 18930 37780 18951 37820
rect 19033 37780 19054 37820
rect 19054 37780 19094 37820
rect 19094 37780 19119 37820
rect 18865 37757 18951 37780
rect 19033 37757 19119 37780
rect 4985 37064 5071 37087
rect 5153 37064 5239 37087
rect 4985 37024 5010 37064
rect 5010 37024 5050 37064
rect 5050 37024 5071 37064
rect 5153 37024 5174 37064
rect 5174 37024 5214 37064
rect 5214 37024 5239 37064
rect 4985 37001 5071 37024
rect 5153 37001 5239 37024
rect 20105 37064 20191 37087
rect 20273 37064 20359 37087
rect 20105 37024 20130 37064
rect 20130 37024 20170 37064
rect 20170 37024 20191 37064
rect 20273 37024 20294 37064
rect 20294 37024 20334 37064
rect 20334 37024 20359 37064
rect 20105 37001 20191 37024
rect 20273 37001 20359 37024
rect 3745 36308 3831 36331
rect 3913 36308 3999 36331
rect 3745 36268 3770 36308
rect 3770 36268 3810 36308
rect 3810 36268 3831 36308
rect 3913 36268 3934 36308
rect 3934 36268 3974 36308
rect 3974 36268 3999 36308
rect 3745 36245 3831 36268
rect 3913 36245 3999 36268
rect 18865 36308 18951 36331
rect 19033 36308 19119 36331
rect 18865 36268 18890 36308
rect 18890 36268 18930 36308
rect 18930 36268 18951 36308
rect 19033 36268 19054 36308
rect 19054 36268 19094 36308
rect 19094 36268 19119 36308
rect 18865 36245 18951 36268
rect 19033 36245 19119 36268
rect 4985 35552 5071 35575
rect 5153 35552 5239 35575
rect 4985 35512 5010 35552
rect 5010 35512 5050 35552
rect 5050 35512 5071 35552
rect 5153 35512 5174 35552
rect 5174 35512 5214 35552
rect 5214 35512 5239 35552
rect 4985 35489 5071 35512
rect 5153 35489 5239 35512
rect 20105 35552 20191 35575
rect 20273 35552 20359 35575
rect 20105 35512 20130 35552
rect 20130 35512 20170 35552
rect 20170 35512 20191 35552
rect 20273 35512 20294 35552
rect 20294 35512 20334 35552
rect 20334 35512 20359 35552
rect 20105 35489 20191 35512
rect 20273 35489 20359 35512
rect 3745 34796 3831 34819
rect 3913 34796 3999 34819
rect 3745 34756 3770 34796
rect 3770 34756 3810 34796
rect 3810 34756 3831 34796
rect 3913 34756 3934 34796
rect 3934 34756 3974 34796
rect 3974 34756 3999 34796
rect 3745 34733 3831 34756
rect 3913 34733 3999 34756
rect 18865 34796 18951 34819
rect 19033 34796 19119 34819
rect 18865 34756 18890 34796
rect 18890 34756 18930 34796
rect 18930 34756 18951 34796
rect 19033 34756 19054 34796
rect 19054 34756 19094 34796
rect 19094 34756 19119 34796
rect 18865 34733 18951 34756
rect 19033 34733 19119 34756
rect 4985 34040 5071 34063
rect 5153 34040 5239 34063
rect 4985 34000 5010 34040
rect 5010 34000 5050 34040
rect 5050 34000 5071 34040
rect 5153 34000 5174 34040
rect 5174 34000 5214 34040
rect 5214 34000 5239 34040
rect 4985 33977 5071 34000
rect 5153 33977 5239 34000
rect 20105 34040 20191 34063
rect 20273 34040 20359 34063
rect 20105 34000 20130 34040
rect 20130 34000 20170 34040
rect 20170 34000 20191 34040
rect 20273 34000 20294 34040
rect 20294 34000 20334 34040
rect 20334 34000 20359 34040
rect 20105 33977 20191 34000
rect 20273 33977 20359 34000
rect 3745 33284 3831 33307
rect 3913 33284 3999 33307
rect 3745 33244 3770 33284
rect 3770 33244 3810 33284
rect 3810 33244 3831 33284
rect 3913 33244 3934 33284
rect 3934 33244 3974 33284
rect 3974 33244 3999 33284
rect 3745 33221 3831 33244
rect 3913 33221 3999 33244
rect 18865 33284 18951 33307
rect 19033 33284 19119 33307
rect 18865 33244 18890 33284
rect 18890 33244 18930 33284
rect 18930 33244 18951 33284
rect 19033 33244 19054 33284
rect 19054 33244 19094 33284
rect 19094 33244 19119 33284
rect 18865 33221 18951 33244
rect 19033 33221 19119 33244
rect 6669 32717 6755 32803
rect 4985 32528 5071 32551
rect 5153 32528 5239 32551
rect 4985 32488 5010 32528
rect 5010 32488 5050 32528
rect 5050 32488 5071 32528
rect 5153 32488 5174 32528
rect 5174 32488 5214 32528
rect 5214 32488 5239 32528
rect 4985 32465 5071 32488
rect 5153 32465 5239 32488
rect 20105 32528 20191 32551
rect 20273 32528 20359 32551
rect 20105 32488 20130 32528
rect 20130 32488 20170 32528
rect 20170 32488 20191 32528
rect 20273 32488 20294 32528
rect 20294 32488 20334 32528
rect 20334 32488 20359 32528
rect 20105 32465 20191 32488
rect 20273 32465 20359 32488
rect 3745 31772 3831 31795
rect 3913 31772 3999 31795
rect 3745 31732 3770 31772
rect 3770 31732 3810 31772
rect 3810 31732 3831 31772
rect 3913 31732 3934 31772
rect 3934 31732 3974 31772
rect 3974 31732 3999 31772
rect 3745 31709 3831 31732
rect 3913 31709 3999 31732
rect 18865 31772 18951 31795
rect 19033 31772 19119 31795
rect 18865 31732 18890 31772
rect 18890 31732 18930 31772
rect 18930 31732 18951 31772
rect 19033 31732 19054 31772
rect 19054 31732 19094 31772
rect 19094 31732 19119 31772
rect 18865 31709 18951 31732
rect 19033 31709 19119 31732
rect 4985 31016 5071 31039
rect 5153 31016 5239 31039
rect 4985 30976 5010 31016
rect 5010 30976 5050 31016
rect 5050 30976 5071 31016
rect 5153 30976 5174 31016
rect 5174 30976 5214 31016
rect 5214 30976 5239 31016
rect 4985 30953 5071 30976
rect 5153 30953 5239 30976
rect 20105 31016 20191 31039
rect 20273 31016 20359 31039
rect 20105 30976 20130 31016
rect 20130 30976 20170 31016
rect 20170 30976 20191 31016
rect 20273 30976 20294 31016
rect 20294 30976 20334 31016
rect 20334 30976 20359 31016
rect 20105 30953 20191 30976
rect 20273 30953 20359 30976
rect 3745 30260 3831 30283
rect 3913 30260 3999 30283
rect 3745 30220 3770 30260
rect 3770 30220 3810 30260
rect 3810 30220 3831 30260
rect 3913 30220 3934 30260
rect 3934 30220 3974 30260
rect 3974 30220 3999 30260
rect 3745 30197 3831 30220
rect 3913 30197 3999 30220
rect 18865 30260 18951 30283
rect 19033 30260 19119 30283
rect 18865 30220 18890 30260
rect 18890 30220 18930 30260
rect 18930 30220 18951 30260
rect 19033 30220 19054 30260
rect 19054 30220 19094 30260
rect 19094 30220 19119 30260
rect 18865 30197 18951 30220
rect 19033 30197 19119 30220
rect 4985 29504 5071 29527
rect 5153 29504 5239 29527
rect 4985 29464 5010 29504
rect 5010 29464 5050 29504
rect 5050 29464 5071 29504
rect 5153 29464 5174 29504
rect 5174 29464 5214 29504
rect 5214 29464 5239 29504
rect 4985 29441 5071 29464
rect 5153 29441 5239 29464
rect 20105 29504 20191 29527
rect 20273 29504 20359 29527
rect 20105 29464 20130 29504
rect 20130 29464 20170 29504
rect 20170 29464 20191 29504
rect 20273 29464 20294 29504
rect 20294 29464 20334 29504
rect 20334 29464 20359 29504
rect 20105 29441 20191 29464
rect 20273 29441 20359 29464
rect 3745 28748 3831 28771
rect 3913 28748 3999 28771
rect 3745 28708 3770 28748
rect 3770 28708 3810 28748
rect 3810 28708 3831 28748
rect 3913 28708 3934 28748
rect 3934 28708 3974 28748
rect 3974 28708 3999 28748
rect 3745 28685 3831 28708
rect 3913 28685 3999 28708
rect 18865 28748 18951 28771
rect 19033 28748 19119 28771
rect 18865 28708 18890 28748
rect 18890 28708 18930 28748
rect 18930 28708 18951 28748
rect 19033 28708 19054 28748
rect 19054 28708 19094 28748
rect 19094 28708 19119 28748
rect 18865 28685 18951 28708
rect 19033 28685 19119 28708
rect 4985 27992 5071 28015
rect 5153 27992 5239 28015
rect 4985 27952 5010 27992
rect 5010 27952 5050 27992
rect 5050 27952 5071 27992
rect 5153 27952 5174 27992
rect 5174 27952 5214 27992
rect 5214 27952 5239 27992
rect 4985 27929 5071 27952
rect 5153 27929 5239 27952
rect 20105 27992 20191 28015
rect 20273 27992 20359 28015
rect 20105 27952 20130 27992
rect 20130 27952 20170 27992
rect 20170 27952 20191 27992
rect 20273 27952 20294 27992
rect 20294 27952 20334 27992
rect 20334 27952 20359 27992
rect 20105 27929 20191 27952
rect 20273 27929 20359 27952
rect 3745 27236 3831 27259
rect 3913 27236 3999 27259
rect 3745 27196 3770 27236
rect 3770 27196 3810 27236
rect 3810 27196 3831 27236
rect 3913 27196 3934 27236
rect 3934 27196 3974 27236
rect 3974 27196 3999 27236
rect 3745 27173 3831 27196
rect 3913 27173 3999 27196
rect 18865 27236 18951 27259
rect 19033 27236 19119 27259
rect 18865 27196 18890 27236
rect 18890 27196 18930 27236
rect 18930 27196 18951 27236
rect 19033 27196 19054 27236
rect 19054 27196 19094 27236
rect 19094 27196 19119 27236
rect 18865 27173 18951 27196
rect 19033 27173 19119 27196
rect 4985 26480 5071 26503
rect 5153 26480 5239 26503
rect 4985 26440 5010 26480
rect 5010 26440 5050 26480
rect 5050 26440 5071 26480
rect 5153 26440 5174 26480
rect 5174 26440 5214 26480
rect 5214 26440 5239 26480
rect 4985 26417 5071 26440
rect 5153 26417 5239 26440
rect 20105 26480 20191 26503
rect 20273 26480 20359 26503
rect 20105 26440 20130 26480
rect 20130 26440 20170 26480
rect 20170 26440 20191 26480
rect 20273 26440 20294 26480
rect 20294 26440 20334 26480
rect 20334 26440 20359 26480
rect 20105 26417 20191 26440
rect 20273 26417 20359 26440
rect 3745 25724 3831 25747
rect 3913 25724 3999 25747
rect 3745 25684 3770 25724
rect 3770 25684 3810 25724
rect 3810 25684 3831 25724
rect 3913 25684 3934 25724
rect 3934 25684 3974 25724
rect 3974 25684 3999 25724
rect 3745 25661 3831 25684
rect 3913 25661 3999 25684
rect 18865 25724 18951 25747
rect 19033 25724 19119 25747
rect 18865 25684 18890 25724
rect 18890 25684 18930 25724
rect 18930 25684 18951 25724
rect 19033 25684 19054 25724
rect 19054 25684 19094 25724
rect 19094 25684 19119 25724
rect 18865 25661 18951 25684
rect 19033 25661 19119 25684
rect 4985 24968 5071 24991
rect 5153 24968 5239 24991
rect 4985 24928 5010 24968
rect 5010 24928 5050 24968
rect 5050 24928 5071 24968
rect 5153 24928 5174 24968
rect 5174 24928 5214 24968
rect 5214 24928 5239 24968
rect 4985 24905 5071 24928
rect 5153 24905 5239 24928
rect 20105 24968 20191 24991
rect 20273 24968 20359 24991
rect 20105 24928 20130 24968
rect 20130 24928 20170 24968
rect 20170 24928 20191 24968
rect 20273 24928 20294 24968
rect 20294 24928 20334 24968
rect 20334 24928 20359 24968
rect 20105 24905 20191 24928
rect 20273 24905 20359 24928
rect 3745 24212 3831 24235
rect 3913 24212 3999 24235
rect 3745 24172 3770 24212
rect 3770 24172 3810 24212
rect 3810 24172 3831 24212
rect 3913 24172 3934 24212
rect 3934 24172 3974 24212
rect 3974 24172 3999 24212
rect 3745 24149 3831 24172
rect 3913 24149 3999 24172
rect 18865 24212 18951 24235
rect 19033 24212 19119 24235
rect 18865 24172 18890 24212
rect 18890 24172 18930 24212
rect 18930 24172 18951 24212
rect 19033 24172 19054 24212
rect 19054 24172 19094 24212
rect 19094 24172 19119 24212
rect 18865 24149 18951 24172
rect 19033 24149 19119 24172
rect 4985 23456 5071 23479
rect 5153 23456 5239 23479
rect 4985 23416 5010 23456
rect 5010 23416 5050 23456
rect 5050 23416 5071 23456
rect 5153 23416 5174 23456
rect 5174 23416 5214 23456
rect 5214 23416 5239 23456
rect 4985 23393 5071 23416
rect 5153 23393 5239 23416
rect 20105 23456 20191 23479
rect 20273 23456 20359 23479
rect 20105 23416 20130 23456
rect 20130 23416 20170 23456
rect 20170 23416 20191 23456
rect 20273 23416 20294 23456
rect 20294 23416 20334 23456
rect 20334 23416 20359 23456
rect 20105 23393 20191 23416
rect 20273 23393 20359 23416
rect 3745 22700 3831 22723
rect 3913 22700 3999 22723
rect 3745 22660 3770 22700
rect 3770 22660 3810 22700
rect 3810 22660 3831 22700
rect 3913 22660 3934 22700
rect 3934 22660 3974 22700
rect 3974 22660 3999 22700
rect 3745 22637 3831 22660
rect 3913 22637 3999 22660
rect 18865 22700 18951 22723
rect 19033 22700 19119 22723
rect 18865 22660 18890 22700
rect 18890 22660 18930 22700
rect 18930 22660 18951 22700
rect 19033 22660 19054 22700
rect 19054 22660 19094 22700
rect 19094 22660 19119 22700
rect 18865 22637 18951 22660
rect 19033 22637 19119 22660
rect 4985 21944 5071 21967
rect 5153 21944 5239 21967
rect 4985 21904 5010 21944
rect 5010 21904 5050 21944
rect 5050 21904 5071 21944
rect 5153 21904 5174 21944
rect 5174 21904 5214 21944
rect 5214 21904 5239 21944
rect 4985 21881 5071 21904
rect 5153 21881 5239 21904
rect 20105 21944 20191 21967
rect 20273 21944 20359 21967
rect 20105 21904 20130 21944
rect 20130 21904 20170 21944
rect 20170 21904 20191 21944
rect 20273 21904 20294 21944
rect 20294 21904 20334 21944
rect 20334 21904 20359 21944
rect 20105 21881 20191 21904
rect 20273 21881 20359 21904
rect 3745 21188 3831 21211
rect 3913 21188 3999 21211
rect 3745 21148 3770 21188
rect 3770 21148 3810 21188
rect 3810 21148 3831 21188
rect 3913 21148 3934 21188
rect 3934 21148 3974 21188
rect 3974 21148 3999 21188
rect 3745 21125 3831 21148
rect 3913 21125 3999 21148
rect 18865 21188 18951 21211
rect 19033 21188 19119 21211
rect 18865 21148 18890 21188
rect 18890 21148 18930 21188
rect 18930 21148 18951 21188
rect 19033 21148 19054 21188
rect 19054 21148 19094 21188
rect 19094 21148 19119 21188
rect 18865 21125 18951 21148
rect 19033 21125 19119 21148
rect 4985 20432 5071 20455
rect 5153 20432 5239 20455
rect 4985 20392 5010 20432
rect 5010 20392 5050 20432
rect 5050 20392 5071 20432
rect 5153 20392 5174 20432
rect 5174 20392 5214 20432
rect 5214 20392 5239 20432
rect 4985 20369 5071 20392
rect 5153 20369 5239 20392
rect 20105 20432 20191 20455
rect 20273 20432 20359 20455
rect 20105 20392 20130 20432
rect 20130 20392 20170 20432
rect 20170 20392 20191 20432
rect 20273 20392 20294 20432
rect 20294 20392 20334 20432
rect 20334 20392 20359 20432
rect 20105 20369 20191 20392
rect 20273 20369 20359 20392
rect 3745 19676 3831 19699
rect 3913 19676 3999 19699
rect 3745 19636 3770 19676
rect 3770 19636 3810 19676
rect 3810 19636 3831 19676
rect 3913 19636 3934 19676
rect 3934 19636 3974 19676
rect 3974 19636 3999 19676
rect 3745 19613 3831 19636
rect 3913 19613 3999 19636
rect 18865 19676 18951 19699
rect 19033 19676 19119 19699
rect 18865 19636 18890 19676
rect 18890 19636 18930 19676
rect 18930 19636 18951 19676
rect 19033 19636 19054 19676
rect 19054 19636 19094 19676
rect 19094 19636 19119 19676
rect 18865 19613 18951 19636
rect 19033 19613 19119 19636
rect 4985 18920 5071 18943
rect 5153 18920 5239 18943
rect 4985 18880 5010 18920
rect 5010 18880 5050 18920
rect 5050 18880 5071 18920
rect 5153 18880 5174 18920
rect 5174 18880 5214 18920
rect 5214 18880 5239 18920
rect 4985 18857 5071 18880
rect 5153 18857 5239 18880
rect 20105 18920 20191 18943
rect 20273 18920 20359 18943
rect 20105 18880 20130 18920
rect 20130 18880 20170 18920
rect 20170 18880 20191 18920
rect 20273 18880 20294 18920
rect 20294 18880 20334 18920
rect 20334 18880 20359 18920
rect 20105 18857 20191 18880
rect 20273 18857 20359 18880
rect 3745 18164 3831 18187
rect 3913 18164 3999 18187
rect 3745 18124 3770 18164
rect 3770 18124 3810 18164
rect 3810 18124 3831 18164
rect 3913 18124 3934 18164
rect 3934 18124 3974 18164
rect 3974 18124 3999 18164
rect 3745 18101 3831 18124
rect 3913 18101 3999 18124
rect 18865 18164 18951 18187
rect 19033 18164 19119 18187
rect 18865 18124 18890 18164
rect 18890 18124 18930 18164
rect 18930 18124 18951 18164
rect 19033 18124 19054 18164
rect 19054 18124 19094 18164
rect 19094 18124 19119 18164
rect 18865 18101 18951 18124
rect 19033 18101 19119 18124
rect 4985 17408 5071 17431
rect 5153 17408 5239 17431
rect 4985 17368 5010 17408
rect 5010 17368 5050 17408
rect 5050 17368 5071 17408
rect 5153 17368 5174 17408
rect 5174 17368 5214 17408
rect 5214 17368 5239 17408
rect 4985 17345 5071 17368
rect 5153 17345 5239 17368
rect 20105 17408 20191 17431
rect 20273 17408 20359 17431
rect 20105 17368 20130 17408
rect 20130 17368 20170 17408
rect 20170 17368 20191 17408
rect 20273 17368 20294 17408
rect 20294 17368 20334 17408
rect 20334 17368 20359 17408
rect 20105 17345 20191 17368
rect 20273 17345 20359 17368
rect 3745 16652 3831 16675
rect 3913 16652 3999 16675
rect 3745 16612 3770 16652
rect 3770 16612 3810 16652
rect 3810 16612 3831 16652
rect 3913 16612 3934 16652
rect 3934 16612 3974 16652
rect 3974 16612 3999 16652
rect 3745 16589 3831 16612
rect 3913 16589 3999 16612
rect 18865 16652 18951 16675
rect 19033 16652 19119 16675
rect 18865 16612 18890 16652
rect 18890 16612 18930 16652
rect 18930 16612 18951 16652
rect 19033 16612 19054 16652
rect 19054 16612 19094 16652
rect 19094 16612 19119 16652
rect 18865 16589 18951 16612
rect 19033 16589 19119 16612
rect 4985 15896 5071 15919
rect 5153 15896 5239 15919
rect 4985 15856 5010 15896
rect 5010 15856 5050 15896
rect 5050 15856 5071 15896
rect 5153 15856 5174 15896
rect 5174 15856 5214 15896
rect 5214 15856 5239 15896
rect 4985 15833 5071 15856
rect 5153 15833 5239 15856
rect 20105 15896 20191 15919
rect 20273 15896 20359 15919
rect 20105 15856 20130 15896
rect 20130 15856 20170 15896
rect 20170 15856 20191 15896
rect 20273 15856 20294 15896
rect 20294 15856 20334 15896
rect 20334 15856 20359 15896
rect 20105 15833 20191 15856
rect 20273 15833 20359 15856
rect 3745 15140 3831 15163
rect 3913 15140 3999 15163
rect 3745 15100 3770 15140
rect 3770 15100 3810 15140
rect 3810 15100 3831 15140
rect 3913 15100 3934 15140
rect 3934 15100 3974 15140
rect 3974 15100 3999 15140
rect 3745 15077 3831 15100
rect 3913 15077 3999 15100
rect 18865 15140 18951 15163
rect 19033 15140 19119 15163
rect 18865 15100 18890 15140
rect 18890 15100 18930 15140
rect 18930 15100 18951 15140
rect 19033 15100 19054 15140
rect 19054 15100 19094 15140
rect 19094 15100 19119 15140
rect 18865 15077 18951 15100
rect 19033 15077 19119 15100
rect 4985 14384 5071 14407
rect 5153 14384 5239 14407
rect 4985 14344 5010 14384
rect 5010 14344 5050 14384
rect 5050 14344 5071 14384
rect 5153 14344 5174 14384
rect 5174 14344 5214 14384
rect 5214 14344 5239 14384
rect 4985 14321 5071 14344
rect 5153 14321 5239 14344
rect 20105 14384 20191 14407
rect 20273 14384 20359 14407
rect 20105 14344 20130 14384
rect 20130 14344 20170 14384
rect 20170 14344 20191 14384
rect 20273 14344 20294 14384
rect 20294 14344 20334 14384
rect 20334 14344 20359 14384
rect 20105 14321 20191 14344
rect 20273 14321 20359 14344
rect 3745 13628 3831 13651
rect 3913 13628 3999 13651
rect 3745 13588 3770 13628
rect 3770 13588 3810 13628
rect 3810 13588 3831 13628
rect 3913 13588 3934 13628
rect 3934 13588 3974 13628
rect 3974 13588 3999 13628
rect 3745 13565 3831 13588
rect 3913 13565 3999 13588
rect 18865 13628 18951 13651
rect 19033 13628 19119 13651
rect 18865 13588 18890 13628
rect 18890 13588 18930 13628
rect 18930 13588 18951 13628
rect 19033 13588 19054 13628
rect 19054 13588 19094 13628
rect 19094 13588 19119 13628
rect 18865 13565 18951 13588
rect 19033 13565 19119 13588
rect 4985 12872 5071 12895
rect 5153 12872 5239 12895
rect 4985 12832 5010 12872
rect 5010 12832 5050 12872
rect 5050 12832 5071 12872
rect 5153 12832 5174 12872
rect 5174 12832 5214 12872
rect 5214 12832 5239 12872
rect 4985 12809 5071 12832
rect 5153 12809 5239 12832
rect 20105 12872 20191 12895
rect 20273 12872 20359 12895
rect 20105 12832 20130 12872
rect 20130 12832 20170 12872
rect 20170 12832 20191 12872
rect 20273 12832 20294 12872
rect 20294 12832 20334 12872
rect 20334 12832 20359 12872
rect 20105 12809 20191 12832
rect 20273 12809 20359 12832
rect 3745 12116 3831 12139
rect 3913 12116 3999 12139
rect 3745 12076 3770 12116
rect 3770 12076 3810 12116
rect 3810 12076 3831 12116
rect 3913 12076 3934 12116
rect 3934 12076 3974 12116
rect 3974 12076 3999 12116
rect 3745 12053 3831 12076
rect 3913 12053 3999 12076
rect 18865 12116 18951 12139
rect 19033 12116 19119 12139
rect 18865 12076 18890 12116
rect 18890 12076 18930 12116
rect 18930 12076 18951 12116
rect 19033 12076 19054 12116
rect 19054 12076 19094 12116
rect 19094 12076 19119 12116
rect 18865 12053 18951 12076
rect 19033 12053 19119 12076
rect 4985 11360 5071 11383
rect 5153 11360 5239 11383
rect 4985 11320 5010 11360
rect 5010 11320 5050 11360
rect 5050 11320 5071 11360
rect 5153 11320 5174 11360
rect 5174 11320 5214 11360
rect 5214 11320 5239 11360
rect 4985 11297 5071 11320
rect 5153 11297 5239 11320
rect 20105 11360 20191 11383
rect 20273 11360 20359 11383
rect 20105 11320 20130 11360
rect 20130 11320 20170 11360
rect 20170 11320 20191 11360
rect 20273 11320 20294 11360
rect 20294 11320 20334 11360
rect 20334 11320 20359 11360
rect 20105 11297 20191 11320
rect 20273 11297 20359 11320
rect 3745 10604 3831 10627
rect 3913 10604 3999 10627
rect 3745 10564 3770 10604
rect 3770 10564 3810 10604
rect 3810 10564 3831 10604
rect 3913 10564 3934 10604
rect 3934 10564 3974 10604
rect 3974 10564 3999 10604
rect 3745 10541 3831 10564
rect 3913 10541 3999 10564
rect 18865 10604 18951 10627
rect 19033 10604 19119 10627
rect 18865 10564 18890 10604
rect 18890 10564 18930 10604
rect 18930 10564 18951 10604
rect 19033 10564 19054 10604
rect 19054 10564 19094 10604
rect 19094 10564 19119 10604
rect 18865 10541 18951 10564
rect 19033 10541 19119 10564
rect 4985 9848 5071 9871
rect 5153 9848 5239 9871
rect 4985 9808 5010 9848
rect 5010 9808 5050 9848
rect 5050 9808 5071 9848
rect 5153 9808 5174 9848
rect 5174 9808 5214 9848
rect 5214 9808 5239 9848
rect 4985 9785 5071 9808
rect 5153 9785 5239 9808
rect 20105 9848 20191 9871
rect 20273 9848 20359 9871
rect 20105 9808 20130 9848
rect 20130 9808 20170 9848
rect 20170 9808 20191 9848
rect 20273 9808 20294 9848
rect 20294 9808 20334 9848
rect 20334 9808 20359 9848
rect 20105 9785 20191 9808
rect 20273 9785 20359 9808
rect 3745 9092 3831 9115
rect 3913 9092 3999 9115
rect 3745 9052 3770 9092
rect 3770 9052 3810 9092
rect 3810 9052 3831 9092
rect 3913 9052 3934 9092
rect 3934 9052 3974 9092
rect 3974 9052 3999 9092
rect 3745 9029 3831 9052
rect 3913 9029 3999 9052
rect 18865 9092 18951 9115
rect 19033 9092 19119 9115
rect 18865 9052 18890 9092
rect 18890 9052 18930 9092
rect 18930 9052 18951 9092
rect 19033 9052 19054 9092
rect 19054 9052 19094 9092
rect 19094 9052 19119 9092
rect 18865 9029 18951 9052
rect 19033 9029 19119 9052
rect 4985 8336 5071 8359
rect 5153 8336 5239 8359
rect 4985 8296 5010 8336
rect 5010 8296 5050 8336
rect 5050 8296 5071 8336
rect 5153 8296 5174 8336
rect 5174 8296 5214 8336
rect 5214 8296 5239 8336
rect 4985 8273 5071 8296
rect 5153 8273 5239 8296
rect 20105 8336 20191 8359
rect 20273 8336 20359 8359
rect 20105 8296 20130 8336
rect 20130 8296 20170 8336
rect 20170 8296 20191 8336
rect 20273 8296 20294 8336
rect 20294 8296 20334 8336
rect 20334 8296 20359 8336
rect 20105 8273 20191 8296
rect 20273 8273 20359 8296
rect 3745 7580 3831 7603
rect 3913 7580 3999 7603
rect 3745 7540 3770 7580
rect 3770 7540 3810 7580
rect 3810 7540 3831 7580
rect 3913 7540 3934 7580
rect 3934 7540 3974 7580
rect 3974 7540 3999 7580
rect 3745 7517 3831 7540
rect 3913 7517 3999 7540
rect 18865 7580 18951 7603
rect 19033 7580 19119 7603
rect 18865 7540 18890 7580
rect 18890 7540 18930 7580
rect 18930 7540 18951 7580
rect 19033 7540 19054 7580
rect 19054 7540 19094 7580
rect 19094 7540 19119 7580
rect 18865 7517 18951 7540
rect 19033 7517 19119 7540
rect 4985 6824 5071 6847
rect 5153 6824 5239 6847
rect 4985 6784 5010 6824
rect 5010 6784 5050 6824
rect 5050 6784 5071 6824
rect 5153 6784 5174 6824
rect 5174 6784 5214 6824
rect 5214 6784 5239 6824
rect 4985 6761 5071 6784
rect 5153 6761 5239 6784
rect 20105 6824 20191 6847
rect 20273 6824 20359 6847
rect 20105 6784 20130 6824
rect 20130 6784 20170 6824
rect 20170 6784 20191 6824
rect 20273 6784 20294 6824
rect 20294 6784 20334 6824
rect 20334 6784 20359 6824
rect 20105 6761 20191 6784
rect 20273 6761 20359 6784
rect 3745 6068 3831 6091
rect 3913 6068 3999 6091
rect 3745 6028 3770 6068
rect 3770 6028 3810 6068
rect 3810 6028 3831 6068
rect 3913 6028 3934 6068
rect 3934 6028 3974 6068
rect 3974 6028 3999 6068
rect 3745 6005 3831 6028
rect 3913 6005 3999 6028
rect 18865 6068 18951 6091
rect 19033 6068 19119 6091
rect 18865 6028 18890 6068
rect 18890 6028 18930 6068
rect 18930 6028 18951 6068
rect 19033 6028 19054 6068
rect 19054 6028 19094 6068
rect 19094 6028 19119 6068
rect 18865 6005 18951 6028
rect 19033 6005 19119 6028
rect 4985 5312 5071 5335
rect 5153 5312 5239 5335
rect 4985 5272 5010 5312
rect 5010 5272 5050 5312
rect 5050 5272 5071 5312
rect 5153 5272 5174 5312
rect 5174 5272 5214 5312
rect 5214 5272 5239 5312
rect 4985 5249 5071 5272
rect 5153 5249 5239 5272
rect 20105 5312 20191 5335
rect 20273 5312 20359 5335
rect 20105 5272 20130 5312
rect 20130 5272 20170 5312
rect 20170 5272 20191 5312
rect 20273 5272 20294 5312
rect 20294 5272 20334 5312
rect 20334 5272 20359 5312
rect 20105 5249 20191 5272
rect 20273 5249 20359 5272
rect 3745 4556 3831 4579
rect 3913 4556 3999 4579
rect 3745 4516 3770 4556
rect 3770 4516 3810 4556
rect 3810 4516 3831 4556
rect 3913 4516 3934 4556
rect 3934 4516 3974 4556
rect 3974 4516 3999 4556
rect 3745 4493 3831 4516
rect 3913 4493 3999 4516
rect 18865 4556 18951 4579
rect 19033 4556 19119 4579
rect 18865 4516 18890 4556
rect 18890 4516 18930 4556
rect 18930 4516 18951 4556
rect 19033 4516 19054 4556
rect 19054 4516 19094 4556
rect 19094 4516 19119 4556
rect 18865 4493 18951 4516
rect 19033 4493 19119 4516
rect 4985 3800 5071 3823
rect 5153 3800 5239 3823
rect 4985 3760 5010 3800
rect 5010 3760 5050 3800
rect 5050 3760 5071 3800
rect 5153 3760 5174 3800
rect 5174 3760 5214 3800
rect 5214 3760 5239 3800
rect 4985 3737 5071 3760
rect 5153 3737 5239 3760
rect 20105 3800 20191 3823
rect 20273 3800 20359 3823
rect 20105 3760 20130 3800
rect 20130 3760 20170 3800
rect 20170 3760 20191 3800
rect 20273 3760 20294 3800
rect 20294 3760 20334 3800
rect 20334 3760 20359 3800
rect 20105 3737 20191 3760
rect 20273 3737 20359 3760
rect 3745 3044 3831 3067
rect 3913 3044 3999 3067
rect 3745 3004 3770 3044
rect 3770 3004 3810 3044
rect 3810 3004 3831 3044
rect 3913 3004 3934 3044
rect 3934 3004 3974 3044
rect 3974 3004 3999 3044
rect 3745 2981 3831 3004
rect 3913 2981 3999 3004
rect 18865 3044 18951 3067
rect 19033 3044 19119 3067
rect 18865 3004 18890 3044
rect 18890 3004 18930 3044
rect 18930 3004 18951 3044
rect 19033 3004 19054 3044
rect 19054 3004 19094 3044
rect 19094 3004 19119 3044
rect 18865 2981 18951 3004
rect 19033 2981 19119 3004
rect 4985 2288 5071 2311
rect 5153 2288 5239 2311
rect 4985 2248 5010 2288
rect 5010 2248 5050 2288
rect 5050 2248 5071 2288
rect 5153 2248 5174 2288
rect 5174 2248 5214 2288
rect 5214 2248 5239 2288
rect 4985 2225 5071 2248
rect 5153 2225 5239 2248
rect 20105 2288 20191 2311
rect 20273 2288 20359 2311
rect 20105 2248 20130 2288
rect 20130 2248 20170 2288
rect 20170 2248 20191 2288
rect 20273 2248 20294 2288
rect 20294 2248 20334 2288
rect 20334 2248 20359 2288
rect 20105 2225 20191 2248
rect 20273 2225 20359 2248
rect 3745 1532 3831 1555
rect 3913 1532 3999 1555
rect 3745 1492 3770 1532
rect 3770 1492 3810 1532
rect 3810 1492 3831 1532
rect 3913 1492 3934 1532
rect 3934 1492 3974 1532
rect 3974 1492 3999 1532
rect 3745 1469 3831 1492
rect 3913 1469 3999 1492
rect 18865 1532 18951 1555
rect 19033 1532 19119 1555
rect 18865 1492 18890 1532
rect 18890 1492 18930 1532
rect 18930 1492 18951 1532
rect 19033 1492 19054 1532
rect 19054 1492 19094 1532
rect 19094 1492 19119 1532
rect 18865 1469 18951 1492
rect 19033 1469 19119 1492
rect 6669 881 6755 967
rect 4985 776 5071 799
rect 5153 776 5239 799
rect 4985 736 5010 776
rect 5010 736 5050 776
rect 5050 736 5071 776
rect 5153 736 5174 776
rect 5174 736 5214 776
rect 5214 736 5239 776
rect 4985 713 5071 736
rect 5153 713 5239 736
rect 20105 776 20191 799
rect 20273 776 20359 799
rect 20105 736 20130 776
rect 20130 736 20170 776
rect 20170 736 20191 776
rect 20273 736 20294 776
rect 20294 736 20334 776
rect 20334 736 20359 776
rect 20105 713 20191 736
rect 20273 713 20359 736
<< metal6 >>
rect 3652 40867 4092 43008
rect 3652 40781 3745 40867
rect 3831 40781 3913 40867
rect 3999 40781 4092 40867
rect 3652 39355 4092 40781
rect 3652 39269 3745 39355
rect 3831 39269 3913 39355
rect 3999 39269 4092 39355
rect 3652 37843 4092 39269
rect 3652 37757 3745 37843
rect 3831 37757 3913 37843
rect 3999 37757 4092 37843
rect 3652 36331 4092 37757
rect 3652 36245 3745 36331
rect 3831 36245 3913 36331
rect 3999 36245 4092 36331
rect 3652 34819 4092 36245
rect 3652 34733 3745 34819
rect 3831 34733 3913 34819
rect 3999 34733 4092 34819
rect 3652 33307 4092 34733
rect 3652 33221 3745 33307
rect 3831 33221 3913 33307
rect 3999 33221 4092 33307
rect 3652 31795 4092 33221
rect 3652 31709 3745 31795
rect 3831 31709 3913 31795
rect 3999 31709 4092 31795
rect 3652 30283 4092 31709
rect 3652 30197 3745 30283
rect 3831 30197 3913 30283
rect 3999 30197 4092 30283
rect 3652 28771 4092 30197
rect 3652 28685 3745 28771
rect 3831 28685 3913 28771
rect 3999 28685 4092 28771
rect 3652 27259 4092 28685
rect 3652 27173 3745 27259
rect 3831 27173 3913 27259
rect 3999 27173 4092 27259
rect 3652 25747 4092 27173
rect 3652 25661 3745 25747
rect 3831 25661 3913 25747
rect 3999 25661 4092 25747
rect 3652 24235 4092 25661
rect 3652 24149 3745 24235
rect 3831 24149 3913 24235
rect 3999 24149 4092 24235
rect 3652 22723 4092 24149
rect 3652 22637 3745 22723
rect 3831 22637 3913 22723
rect 3999 22637 4092 22723
rect 3652 21211 4092 22637
rect 3652 21125 3745 21211
rect 3831 21125 3913 21211
rect 3999 21125 4092 21211
rect 3652 19699 4092 21125
rect 3652 19613 3745 19699
rect 3831 19613 3913 19699
rect 3999 19613 4092 19699
rect 3652 18187 4092 19613
rect 3652 18101 3745 18187
rect 3831 18101 3913 18187
rect 3999 18101 4092 18187
rect 3652 16675 4092 18101
rect 3652 16589 3745 16675
rect 3831 16589 3913 16675
rect 3999 16589 4092 16675
rect 3652 15163 4092 16589
rect 3652 15077 3745 15163
rect 3831 15077 3913 15163
rect 3999 15077 4092 15163
rect 3652 13651 4092 15077
rect 3652 13565 3745 13651
rect 3831 13565 3913 13651
rect 3999 13565 4092 13651
rect 3652 12139 4092 13565
rect 3652 12053 3745 12139
rect 3831 12053 3913 12139
rect 3999 12053 4092 12139
rect 3652 10627 4092 12053
rect 3652 10541 3745 10627
rect 3831 10541 3913 10627
rect 3999 10541 4092 10627
rect 3652 9115 4092 10541
rect 3652 9029 3745 9115
rect 3831 9029 3913 9115
rect 3999 9029 4092 9115
rect 3652 7603 4092 9029
rect 3652 7517 3745 7603
rect 3831 7517 3913 7603
rect 3999 7517 4092 7603
rect 3652 6091 4092 7517
rect 3652 6005 3745 6091
rect 3831 6005 3913 6091
rect 3999 6005 4092 6091
rect 3652 4579 4092 6005
rect 3652 4493 3745 4579
rect 3831 4493 3913 4579
rect 3999 4493 4092 4579
rect 3652 3067 4092 4493
rect 3652 2981 3745 3067
rect 3831 2981 3913 3067
rect 3999 2981 4092 3067
rect 3652 1555 4092 2981
rect 3652 1469 3745 1555
rect 3831 1469 3913 1555
rect 3999 1469 4092 1555
rect 3652 0 4092 1469
rect 4892 41623 5332 43008
rect 4892 41537 4985 41623
rect 5071 41537 5153 41623
rect 5239 41537 5332 41623
rect 4892 40111 5332 41537
rect 4892 40025 4985 40111
rect 5071 40025 5153 40111
rect 5239 40025 5332 40111
rect 4892 38599 5332 40025
rect 4892 38513 4985 38599
rect 5071 38513 5153 38599
rect 5239 38513 5332 38599
rect 4892 37087 5332 38513
rect 4892 37001 4985 37087
rect 5071 37001 5153 37087
rect 5239 37001 5332 37087
rect 4892 35575 5332 37001
rect 4892 35489 4985 35575
rect 5071 35489 5153 35575
rect 5239 35489 5332 35575
rect 4892 34063 5332 35489
rect 4892 33977 4985 34063
rect 5071 33977 5153 34063
rect 5239 33977 5332 34063
rect 4892 32551 5332 33977
rect 18772 40867 19212 43008
rect 18772 40781 18865 40867
rect 18951 40781 19033 40867
rect 19119 40781 19212 40867
rect 18772 39355 19212 40781
rect 18772 39269 18865 39355
rect 18951 39269 19033 39355
rect 19119 39269 19212 39355
rect 18772 37843 19212 39269
rect 18772 37757 18865 37843
rect 18951 37757 19033 37843
rect 19119 37757 19212 37843
rect 18772 36331 19212 37757
rect 18772 36245 18865 36331
rect 18951 36245 19033 36331
rect 19119 36245 19212 36331
rect 18772 34819 19212 36245
rect 18772 34733 18865 34819
rect 18951 34733 19033 34819
rect 19119 34733 19212 34819
rect 18772 33307 19212 34733
rect 18772 33221 18865 33307
rect 18951 33221 19033 33307
rect 19119 33221 19212 33307
rect 4892 32465 4985 32551
rect 5071 32465 5153 32551
rect 5239 32465 5332 32551
rect 4892 31039 5332 32465
rect 4892 30953 4985 31039
rect 5071 30953 5153 31039
rect 5239 30953 5332 31039
rect 4892 29527 5332 30953
rect 4892 29441 4985 29527
rect 5071 29441 5153 29527
rect 5239 29441 5332 29527
rect 4892 28015 5332 29441
rect 4892 27929 4985 28015
rect 5071 27929 5153 28015
rect 5239 27929 5332 28015
rect 4892 26503 5332 27929
rect 4892 26417 4985 26503
rect 5071 26417 5153 26503
rect 5239 26417 5332 26503
rect 4892 24991 5332 26417
rect 4892 24905 4985 24991
rect 5071 24905 5153 24991
rect 5239 24905 5332 24991
rect 4892 23479 5332 24905
rect 4892 23393 4985 23479
rect 5071 23393 5153 23479
rect 5239 23393 5332 23479
rect 4892 21967 5332 23393
rect 4892 21881 4985 21967
rect 5071 21881 5153 21967
rect 5239 21881 5332 21967
rect 4892 20455 5332 21881
rect 4892 20369 4985 20455
rect 5071 20369 5153 20455
rect 5239 20369 5332 20455
rect 4892 18943 5332 20369
rect 4892 18857 4985 18943
rect 5071 18857 5153 18943
rect 5239 18857 5332 18943
rect 4892 17431 5332 18857
rect 4892 17345 4985 17431
rect 5071 17345 5153 17431
rect 5239 17345 5332 17431
rect 4892 15919 5332 17345
rect 4892 15833 4985 15919
rect 5071 15833 5153 15919
rect 5239 15833 5332 15919
rect 4892 14407 5332 15833
rect 4892 14321 4985 14407
rect 5071 14321 5153 14407
rect 5239 14321 5332 14407
rect 4892 12895 5332 14321
rect 4892 12809 4985 12895
rect 5071 12809 5153 12895
rect 5239 12809 5332 12895
rect 4892 11383 5332 12809
rect 4892 11297 4985 11383
rect 5071 11297 5153 11383
rect 5239 11297 5332 11383
rect 4892 9871 5332 11297
rect 4892 9785 4985 9871
rect 5071 9785 5153 9871
rect 5239 9785 5332 9871
rect 4892 8359 5332 9785
rect 4892 8273 4985 8359
rect 5071 8273 5153 8359
rect 5239 8273 5332 8359
rect 4892 6847 5332 8273
rect 4892 6761 4985 6847
rect 5071 6761 5153 6847
rect 5239 6761 5332 6847
rect 4892 5335 5332 6761
rect 4892 5249 4985 5335
rect 5071 5249 5153 5335
rect 5239 5249 5332 5335
rect 4892 3823 5332 5249
rect 4892 3737 4985 3823
rect 5071 3737 5153 3823
rect 5239 3737 5332 3823
rect 4892 2311 5332 3737
rect 4892 2225 4985 2311
rect 5071 2225 5153 2311
rect 5239 2225 5332 2311
rect 4892 799 5332 2225
rect 4892 713 4985 799
rect 5071 713 5153 799
rect 5239 713 5332 799
rect 6548 32803 6876 32924
rect 6548 32717 6669 32803
rect 6755 32717 6876 32803
rect 6548 967 6876 32717
rect 6548 881 6669 967
rect 6755 881 6876 967
rect 6548 760 6876 881
rect 18772 31795 19212 33221
rect 18772 31709 18865 31795
rect 18951 31709 19033 31795
rect 19119 31709 19212 31795
rect 18772 30283 19212 31709
rect 18772 30197 18865 30283
rect 18951 30197 19033 30283
rect 19119 30197 19212 30283
rect 18772 28771 19212 30197
rect 18772 28685 18865 28771
rect 18951 28685 19033 28771
rect 19119 28685 19212 28771
rect 18772 27259 19212 28685
rect 18772 27173 18865 27259
rect 18951 27173 19033 27259
rect 19119 27173 19212 27259
rect 18772 25747 19212 27173
rect 18772 25661 18865 25747
rect 18951 25661 19033 25747
rect 19119 25661 19212 25747
rect 18772 24235 19212 25661
rect 18772 24149 18865 24235
rect 18951 24149 19033 24235
rect 19119 24149 19212 24235
rect 18772 22723 19212 24149
rect 18772 22637 18865 22723
rect 18951 22637 19033 22723
rect 19119 22637 19212 22723
rect 18772 21211 19212 22637
rect 18772 21125 18865 21211
rect 18951 21125 19033 21211
rect 19119 21125 19212 21211
rect 18772 19699 19212 21125
rect 18772 19613 18865 19699
rect 18951 19613 19033 19699
rect 19119 19613 19212 19699
rect 18772 18187 19212 19613
rect 18772 18101 18865 18187
rect 18951 18101 19033 18187
rect 19119 18101 19212 18187
rect 18772 16675 19212 18101
rect 18772 16589 18865 16675
rect 18951 16589 19033 16675
rect 19119 16589 19212 16675
rect 18772 15163 19212 16589
rect 18772 15077 18865 15163
rect 18951 15077 19033 15163
rect 19119 15077 19212 15163
rect 18772 13651 19212 15077
rect 18772 13565 18865 13651
rect 18951 13565 19033 13651
rect 19119 13565 19212 13651
rect 18772 12139 19212 13565
rect 18772 12053 18865 12139
rect 18951 12053 19033 12139
rect 19119 12053 19212 12139
rect 18772 10627 19212 12053
rect 18772 10541 18865 10627
rect 18951 10541 19033 10627
rect 19119 10541 19212 10627
rect 18772 9115 19212 10541
rect 18772 9029 18865 9115
rect 18951 9029 19033 9115
rect 19119 9029 19212 9115
rect 18772 7603 19212 9029
rect 18772 7517 18865 7603
rect 18951 7517 19033 7603
rect 19119 7517 19212 7603
rect 18772 6091 19212 7517
rect 18772 6005 18865 6091
rect 18951 6005 19033 6091
rect 19119 6005 19212 6091
rect 18772 4579 19212 6005
rect 18772 4493 18865 4579
rect 18951 4493 19033 4579
rect 19119 4493 19212 4579
rect 18772 3067 19212 4493
rect 18772 2981 18865 3067
rect 18951 2981 19033 3067
rect 19119 2981 19212 3067
rect 18772 1555 19212 2981
rect 18772 1469 18865 1555
rect 18951 1469 19033 1555
rect 19119 1469 19212 1555
rect 4892 0 5332 713
rect 18772 0 19212 1469
rect 20012 41623 20452 43008
rect 20012 41537 20105 41623
rect 20191 41537 20273 41623
rect 20359 41537 20452 41623
rect 20012 40111 20452 41537
rect 20012 40025 20105 40111
rect 20191 40025 20273 40111
rect 20359 40025 20452 40111
rect 20012 38599 20452 40025
rect 20012 38513 20105 38599
rect 20191 38513 20273 38599
rect 20359 38513 20452 38599
rect 20012 37087 20452 38513
rect 20012 37001 20105 37087
rect 20191 37001 20273 37087
rect 20359 37001 20452 37087
rect 20012 35575 20452 37001
rect 20012 35489 20105 35575
rect 20191 35489 20273 35575
rect 20359 35489 20452 35575
rect 20012 34063 20452 35489
rect 20012 33977 20105 34063
rect 20191 33977 20273 34063
rect 20359 33977 20452 34063
rect 20012 32551 20452 33977
rect 20012 32465 20105 32551
rect 20191 32465 20273 32551
rect 20359 32465 20452 32551
rect 20012 31039 20452 32465
rect 20012 30953 20105 31039
rect 20191 30953 20273 31039
rect 20359 30953 20452 31039
rect 20012 29527 20452 30953
rect 20012 29441 20105 29527
rect 20191 29441 20273 29527
rect 20359 29441 20452 29527
rect 20012 28015 20452 29441
rect 20012 27929 20105 28015
rect 20191 27929 20273 28015
rect 20359 27929 20452 28015
rect 20012 26503 20452 27929
rect 20012 26417 20105 26503
rect 20191 26417 20273 26503
rect 20359 26417 20452 26503
rect 20012 24991 20452 26417
rect 20012 24905 20105 24991
rect 20191 24905 20273 24991
rect 20359 24905 20452 24991
rect 20012 23479 20452 24905
rect 20012 23393 20105 23479
rect 20191 23393 20273 23479
rect 20359 23393 20452 23479
rect 20012 21967 20452 23393
rect 20012 21881 20105 21967
rect 20191 21881 20273 21967
rect 20359 21881 20452 21967
rect 20012 20455 20452 21881
rect 20012 20369 20105 20455
rect 20191 20369 20273 20455
rect 20359 20369 20452 20455
rect 20012 18943 20452 20369
rect 20012 18857 20105 18943
rect 20191 18857 20273 18943
rect 20359 18857 20452 18943
rect 20012 17431 20452 18857
rect 20012 17345 20105 17431
rect 20191 17345 20273 17431
rect 20359 17345 20452 17431
rect 20012 15919 20452 17345
rect 20012 15833 20105 15919
rect 20191 15833 20273 15919
rect 20359 15833 20452 15919
rect 20012 14407 20452 15833
rect 20012 14321 20105 14407
rect 20191 14321 20273 14407
rect 20359 14321 20452 14407
rect 20012 12895 20452 14321
rect 20012 12809 20105 12895
rect 20191 12809 20273 12895
rect 20359 12809 20452 12895
rect 20012 11383 20452 12809
rect 20012 11297 20105 11383
rect 20191 11297 20273 11383
rect 20359 11297 20452 11383
rect 20012 9871 20452 11297
rect 20012 9785 20105 9871
rect 20191 9785 20273 9871
rect 20359 9785 20452 9871
rect 20012 8359 20452 9785
rect 20012 8273 20105 8359
rect 20191 8273 20273 8359
rect 20359 8273 20452 8359
rect 20012 6847 20452 8273
rect 20012 6761 20105 6847
rect 20191 6761 20273 6847
rect 20359 6761 20452 6847
rect 20012 5335 20452 6761
rect 20012 5249 20105 5335
rect 20191 5249 20273 5335
rect 20359 5249 20452 5335
rect 20012 3823 20452 5249
rect 20012 3737 20105 3823
rect 20191 3737 20273 3823
rect 20359 3737 20452 3823
rect 20012 2311 20452 3737
rect 20012 2225 20105 2311
rect 20191 2225 20273 2311
rect 20359 2225 20452 2311
rect 20012 799 20452 2225
rect 20012 713 20105 799
rect 20191 713 20273 799
rect 20359 713 20452 799
rect 20012 0 20452 713
use sg13g2_inv_1  _209_
timestamp 1676382929
transform -1 0 9984 0 1 34020
box -48 -56 336 834
use sg13g2_inv_1  _210_
timestamp 1676382929
transform 1 0 8640 0 1 32508
box -48 -56 336 834
use sg13g2_inv_1  _211_
timestamp 1676382929
transform -1 0 7776 0 -1 34020
box -48 -56 336 834
use sg13g2_inv_1  _212_
timestamp 1676382929
transform -1 0 12672 0 1 38556
box -48 -56 336 834
use sg13g2_inv_1  _213_
timestamp 1676382929
transform 1 0 14496 0 -1 32508
box -48 -56 336 834
use sg13g2_inv_1  _214_
timestamp 1676382929
transform -1 0 6624 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _215_
timestamp 1676382929
transform 1 0 13440 0 1 24948
box -48 -56 336 834
use sg13g2_inv_1  _216_
timestamp 1676382929
transform 1 0 5760 0 -1 20412
box -48 -56 336 834
use sg13g2_inv_1  _217_
timestamp 1676382929
transform 1 0 3456 0 1 17388
box -48 -56 336 834
use sg13g2_inv_1  _218_
timestamp 1676382929
transform 1 0 11712 0 1 26460
box -48 -56 336 834
use sg13g2_inv_1  _219_
timestamp 1676382929
transform 1 0 12384 0 -1 30996
box -48 -56 336 834
use sg13g2_inv_1  _220_
timestamp 1676382929
transform 1 0 7200 0 -1 21924
box -48 -56 336 834
use sg13g2_inv_1  _221_
timestamp 1676382929
transform 1 0 7680 0 -1 20412
box -48 -56 336 834
use sg13g2_inv_1  _222_
timestamp 1676382929
transform 1 0 8928 0 -1 27972
box -48 -56 336 834
use sg13g2_inv_1  _223_
timestamp 1676382929
transform 1 0 8256 0 1 29484
box -48 -56 336 834
use sg13g2_inv_1  _224_
timestamp 1676382929
transform -1 0 14592 0 1 27972
box -48 -56 336 834
use sg13g2_inv_1  _225_
timestamp 1676382929
transform 1 0 15552 0 -1 26460
box -48 -56 336 834
use sg13g2_inv_1  _226_
timestamp 1676382929
transform 1 0 14016 0 1 26460
box -48 -56 336 834
use sg13g2_inv_1  _227_
timestamp 1676382929
transform 1 0 2880 0 -1 21924
box -48 -56 336 834
use sg13g2_inv_1  _228_
timestamp 1676382929
transform 1 0 4608 0 -1 23436
box -48 -56 336 834
use sg13g2_mux2_1  _229_
timestamp 1677247768
transform 1 0 8352 0 -1 34020
box -48 -56 1008 834
use sg13g2_nand2_1  _230_
timestamp 1676557249
transform 1 0 9888 0 1 32508
box -48 -56 432 834
use sg13g2_mux2_1  _231_
timestamp 1677247768
transform 1 0 8736 0 1 34020
box -48 -56 1008 834
use sg13g2_a21oi_1  _232_
timestamp 1683973020
transform 1 0 9408 0 1 32508
box -48 -56 528 834
use sg13g2_mux2_1  _233_
timestamp 1677247768
transform -1 0 9312 0 -1 35532
box -48 -56 1008 834
use sg13g2_nand2b_1  _234_
timestamp 1676567195
transform 1 0 7872 0 -1 32508
box -48 -56 528 834
use sg13g2_o21ai_1  _235_
timestamp 1685175443
transform -1 0 6720 0 1 35532
box -48 -56 538 834
use sg13g2_nand2b_1  _236_
timestamp 1676567195
transform -1 0 6432 0 1 34020
box -48 -56 528 834
use sg13g2_a21oi_1  _237_
timestamp 1683973020
transform 1 0 7872 0 -1 35532
box -48 -56 528 834
use sg13g2_a221oi_1  _238_
timestamp 1685197497
transform -1 0 10080 0 -1 35532
box -48 -56 816 834
use sg13g2_nor2_1  _239_
timestamp 1676627187
transform -1 0 11616 0 -1 35532
box -48 -56 432 834
use sg13g2_nor2b_1  _240_
timestamp 1685181386
transform 1 0 8544 0 -1 37044
box -54 -56 528 834
use sg13g2_nor2b_1  _241_
timestamp 1685181386
transform -1 0 7776 0 1 37044
box -54 -56 528 834
use sg13g2_a22oi_1  _242_
timestamp 1685173987
transform 1 0 8928 0 1 35532
box -48 -56 624 834
use sg13g2_a21oi_1  _243_
timestamp 1683973020
transform -1 0 9408 0 1 32508
box -48 -56 528 834
use sg13g2_o21ai_1  _244_
timestamp 1685175443
transform -1 0 11232 0 -1 35532
box -48 -56 538 834
use sg13g2_a22oi_1  _245_
timestamp 1685173987
transform 1 0 7776 0 -1 34020
box -48 -56 624 834
use sg13g2_and2_1  _246_
timestamp 1676901763
transform 1 0 7776 0 1 37044
box -48 -56 528 834
use sg13g2_a22oi_1  _247_
timestamp 1685173987
transform -1 0 9888 0 -1 34020
box -48 -56 624 834
use sg13g2_a21o_1  _248_
timestamp 1677175127
transform -1 0 10752 0 -1 35532
box -48 -56 720 834
use sg13g2_mux4_1  _249_
timestamp 1677257233
transform 1 0 8256 0 1 40068
box -48 -56 2064 834
use sg13g2_inv_1  _250_
timestamp 1676382929
transform 1 0 11328 0 1 27972
box -48 -56 336 834
use sg13g2_mux4_1  _251_
timestamp 1677257233
transform 1 0 9984 0 -1 14364
box -48 -56 2064 834
use sg13g2_nor2b_1  _252_
timestamp 1685181386
transform 1 0 3552 0 1 26460
box -54 -56 528 834
use sg13g2_a21oi_1  _253_
timestamp 1683973020
transform 1 0 5088 0 -1 26460
box -48 -56 528 834
use sg13g2_nand3b_1  _254_
timestamp 1676573470
transform 1 0 5664 0 1 26460
box -48 -56 720 834
use sg13g2_o21ai_1  _255_
timestamp 1685175443
transform 1 0 6336 0 1 26460
box -48 -56 538 834
use sg13g2_mux4_1  _256_
timestamp 1677257233
transform 1 0 3072 0 -1 26460
box -48 -56 2064 834
use sg13g2_mux2_1  _257_
timestamp 1677247768
transform 1 0 5568 0 -1 26460
box -48 -56 1008 834
use sg13g2_mux4_1  _258_
timestamp 1677257233
transform 1 0 10368 0 1 38556
box -48 -56 2064 834
use sg13g2_mux4_1  _259_
timestamp 1677257233
transform 1 0 13248 0 1 34020
box -48 -56 2064 834
use sg13g2_nor2b_1  _260_
timestamp 1685181386
transform 1 0 17472 0 -1 27972
box -54 -56 528 834
use sg13g2_a21oi_1  _261_
timestamp 1683973020
transform 1 0 18144 0 -1 29484
box -48 -56 528 834
use sg13g2_nand3b_1  _262_
timestamp 1676573470
transform 1 0 17952 0 -1 27972
box -48 -56 720 834
use sg13g2_o21ai_1  _263_
timestamp 1685175443
transform 1 0 18624 0 1 30996
box -48 -56 538 834
use sg13g2_mux4_1  _264_
timestamp 1677257233
transform 1 0 16320 0 1 27972
box -48 -56 2064 834
use sg13g2_mux2_1  _265_
timestamp 1677247768
transform 1 0 19008 0 -1 27972
box -48 -56 1008 834
use sg13g2_mux4_1  _266_
timestamp 1677257233
transform 1 0 13632 0 -1 18900
box -48 -56 2064 834
use sg13g2_mux4_1  _267_
timestamp 1677257233
transform 1 0 6144 0 -1 40068
box -48 -56 2064 834
use sg13g2_mux4_1  _268_
timestamp 1677257233
transform 1 0 16992 0 1 21924
box -48 -56 2064 834
use sg13g2_nand3b_1  _269_
timestamp 1676573470
transform 1 0 18720 0 1 23436
box -48 -56 720 834
use sg13g2_nor2b_1  _270_
timestamp 1685181386
transform 1 0 18048 0 -1 21924
box -54 -56 528 834
use sg13g2_a21oi_1  _271_
timestamp 1683973020
transform 1 0 18240 0 1 23436
box -48 -56 528 834
use sg13g2_o21ai_1  _272_
timestamp 1685175443
transform 1 0 19392 0 1 23436
box -48 -56 538 834
use sg13g2_mux2_1  _273_
timestamp 1677247768
transform 1 0 19008 0 1 21924
box -48 -56 1008 834
use sg13g2_mux4_1  _274_
timestamp 1677257233
transform 1 0 6048 0 1 6804
box -48 -56 2064 834
use sg13g2_mux4_1  _275_
timestamp 1677257233
transform 1 0 4896 0 1 37044
box -48 -56 2064 834
use sg13g2_inv_1  _276_
timestamp 1676382929
transform 1 0 6240 0 -1 20412
box -48 -56 336 834
use sg13g2_nor2b_1  _277_
timestamp 1685181386
transform 1 0 7104 0 -1 23436
box -54 -56 528 834
use sg13g2_a21oi_1  _278_
timestamp 1683973020
transform 1 0 7584 0 -1 23436
box -48 -56 528 834
use sg13g2_nand3b_1  _279_
timestamp 1676573470
transform -1 0 10368 0 -1 23436
box -48 -56 720 834
use sg13g2_o21ai_1  _280_
timestamp 1685175443
transform 1 0 9312 0 1 20412
box -48 -56 538 834
use sg13g2_mux4_1  _281_
timestamp 1677257233
transform 1 0 7872 0 1 21924
box -48 -56 2064 834
use sg13g2_mux2_1  _282_
timestamp 1677247768
transform 1 0 11520 0 1 21924
box -48 -56 1008 834
use sg13g2_mux4_1  _283_
timestamp 1677257233
transform 1 0 9408 0 1 15876
box -48 -56 2064 834
use sg13g2_mux4_1  _284_
timestamp 1677257233
transform 1 0 6240 0 -1 37044
box -48 -56 2064 834
use sg13g2_nand3b_1  _285_
timestamp 1676573470
transform 1 0 10272 0 1 24948
box -48 -56 720 834
use sg13g2_nor2b_1  _286_
timestamp 1685181386
transform 1 0 9216 0 1 24948
box -54 -56 528 834
use sg13g2_a21oi_1  _287_
timestamp 1683973020
transform 1 0 9792 0 1 24948
box -48 -56 528 834
use sg13g2_o21ai_1  _288_
timestamp 1685175443
transform 1 0 10848 0 -1 24948
box -48 -56 538 834
use sg13g2_mux4_1  _289_
timestamp 1677257233
transform 1 0 8832 0 -1 24948
box -48 -56 2064 834
use sg13g2_mux2_1  _290_
timestamp 1677247768
transform 1 0 11328 0 -1 24948
box -48 -56 1008 834
use sg13g2_mux4_1  _291_
timestamp 1677257233
transform 1 0 13152 0 -1 40068
box -48 -56 2064 834
use sg13g2_mux4_1  _292_
timestamp 1677257233
transform 1 0 8256 0 1 37044
box -48 -56 2064 834
use sg13g2_mux4_1  _293_
timestamp 1677257233
transform 1 0 17856 0 -1 35532
box -48 -56 2064 834
use sg13g2_nand3b_1  _294_
timestamp 1676573470
transform 1 0 19584 0 1 35532
box -48 -56 720 834
use sg13g2_nor2b_1  _295_
timestamp 1685181386
transform 1 0 17760 0 1 34020
box -54 -56 528 834
use sg13g2_a21oi_1  _296_
timestamp 1683973020
transform -1 0 17760 0 -1 37044
box -48 -56 528 834
use sg13g2_o21ai_1  _297_
timestamp 1685175443
transform 1 0 19872 0 -1 35532
box -48 -56 538 834
use sg13g2_mux2_1  _298_
timestamp 1677247768
transform 1 0 19296 0 1 32508
box -48 -56 1008 834
use sg13g2_mux4_1  _299_
timestamp 1677257233
transform 1 0 11904 0 1 17388
box -48 -56 2064 834
use sg13g2_mux4_1  _300_
timestamp 1677257233
transform 1 0 4224 0 1 35532
box -48 -56 2064 834
use sg13g2_nor2b_1  _301_
timestamp 1685181386
transform 1 0 14496 0 -1 21924
box -54 -56 528 834
use sg13g2_a21oi_1  _302_
timestamp 1683973020
transform 1 0 14880 0 -1 20412
box -48 -56 528 834
use sg13g2_nand3b_1  _303_
timestamp 1676573470
transform 1 0 15072 0 1 21924
box -48 -56 720 834
use sg13g2_o21ai_1  _304_
timestamp 1685175443
transform 1 0 15744 0 1 21924
box -48 -56 538 834
use sg13g2_mux4_1  _305_
timestamp 1677257233
transform 1 0 13056 0 1 21924
box -48 -56 2064 834
use sg13g2_mux2_1  _306_
timestamp 1677247768
transform 1 0 15072 0 -1 21924
box -48 -56 1008 834
use sg13g2_mux4_1  _307_
timestamp 1677257233
transform 1 0 7968 0 -1 2268
box -48 -56 2064 834
use sg13g2_inv_1  _308_
timestamp 1676382929
transform -1 0 5184 0 1 20412
box -48 -56 336 834
use sg13g2_mux4_1  _309_
timestamp 1677257233
transform 1 0 5856 0 -1 5292
box -48 -56 2064 834
use sg13g2_inv_1  _310_
timestamp 1676382929
transform -1 0 4704 0 -1 20412
box -48 -56 336 834
use sg13g2_nand3_1  _311_
timestamp 1683988354
transform 1 0 4032 0 -1 18900
box -48 -56 528 834
use sg13g2_or2_1  _312_
timestamp 1684236171
transform 1 0 3936 0 1 20412
box -48 -56 528 834
use sg13g2_o21ai_1  _313_
timestamp 1685175443
transform -1 0 4896 0 1 20412
box -48 -56 538 834
use sg13g2_o21ai_1  _314_
timestamp 1685175443
transform 1 0 4512 0 -1 18900
box -48 -56 538 834
use sg13g2_mux4_1  _315_
timestamp 1677257233
transform 1 0 2304 0 1 18900
box -48 -56 2064 834
use sg13g2_mux2_1  _316_
timestamp 1677247768
transform 1 0 4800 0 -1 20412
box -48 -56 1008 834
use sg13g2_mux4_1  _317_
timestamp 1677257233
transform 1 0 7008 0 -1 15876
box -48 -56 2064 834
use sg13g2_mux4_1  _318_
timestamp 1677257233
transform 1 0 3264 0 1 27972
box -48 -56 2064 834
use sg13g2_nand3b_1  _319_
timestamp 1676573470
transform 1 0 5472 0 -1 29484
box -48 -56 720 834
use sg13g2_nor2b_1  _320_
timestamp 1685181386
transform -1 0 6336 0 1 29484
box -54 -56 528 834
use sg13g2_a21oi_1  _321_
timestamp 1683973020
transform -1 0 5856 0 1 29484
box -48 -56 528 834
use sg13g2_o21ai_1  _322_
timestamp 1685175443
transform 1 0 6144 0 -1 29484
box -48 -56 538 834
use sg13g2_mux2_1  _323_
timestamp 1677247768
transform 1 0 5280 0 -1 27972
box -48 -56 1008 834
use sg13g2_mux4_1  _324_
timestamp 1677257233
transform 1 0 13920 0 1 38556
box -48 -56 2064 834
use sg13g2_mux4_1  _325_
timestamp 1677257233
transform 1 0 16704 0 -1 30996
box -48 -56 2064 834
use sg13g2_nand3b_1  _326_
timestamp 1676573470
transform 1 0 17952 0 1 30996
box -48 -56 720 834
use sg13g2_nor2b_1  _327_
timestamp 1685181386
transform 1 0 16224 0 -1 30996
box -54 -56 528 834
use sg13g2_a21oi_1  _328_
timestamp 1683973020
transform 1 0 17088 0 1 30996
box -48 -56 528 834
use sg13g2_o21ai_1  _329_
timestamp 1685175443
transform 1 0 19104 0 1 30996
box -48 -56 538 834
use sg13g2_mux2_1  _330_
timestamp 1677247768
transform 1 0 19008 0 -1 29484
box -48 -56 1008 834
use sg13g2_mux4_1  _331_
timestamp 1677257233
transform 1 0 13440 0 1 15876
box -48 -56 2064 834
use sg13g2_nor2b_1  _332_
timestamp 1685181386
transform 1 0 18048 0 -1 20412
box -54 -56 528 834
use sg13g2_a21oi_1  _333_
timestamp 1683973020
transform 1 0 18720 0 -1 18900
box -48 -56 528 834
use sg13g2_nand3b_1  _334_
timestamp 1676573470
transform 1 0 19200 0 1 20412
box -48 -56 720 834
use sg13g2_o21ai_1  _335_
timestamp 1685175443
transform 1 0 19872 0 1 20412
box -48 -56 538 834
use sg13g2_mux4_1  _336_
timestamp 1677257233
transform 1 0 17184 0 1 20412
box -48 -56 2064 834
use sg13g2_mux2_1  _337_
timestamp 1677247768
transform 1 0 19392 0 1 18900
box -48 -56 1008 834
use sg13g2_mux4_1  _338_
timestamp 1677257233
transform 1 0 5472 0 -1 11340
box -48 -56 2064 834
use sg13g2_nor2b_1  _339_
timestamp 1685181386
transform 1 0 4896 0 1 23436
box -54 -56 528 834
use sg13g2_a21oi_1  _340_
timestamp 1683973020
transform 1 0 5376 0 1 23436
box -48 -56 528 834
use sg13g2_nand3b_1  _341_
timestamp 1676573470
transform 1 0 6432 0 -1 24948
box -48 -56 720 834
use sg13g2_o21ai_1  _342_
timestamp 1685175443
transform 1 0 7872 0 1 23436
box -48 -56 538 834
use sg13g2_mux4_1  _343_
timestamp 1677257233
transform 1 0 5856 0 1 23436
box -48 -56 2064 834
use sg13g2_mux2_1  _344_
timestamp 1677247768
transform 1 0 7488 0 -1 24948
box -48 -56 1008 834
use sg13g2_mux4_1  _345_
timestamp 1677257233
transform 1 0 9984 0 1 14364
box -48 -56 2064 834
use sg13g2_mux4_1  _346_
timestamp 1677257233
transform 1 0 8736 0 -1 26460
box -48 -56 2064 834
use sg13g2_nand3b_1  _347_
timestamp 1676573470
transform 1 0 10560 0 1 26460
box -48 -56 720 834
use sg13g2_nor2b_1  _348_
timestamp 1685181386
transform 1 0 8448 0 -1 27972
box -54 -56 528 834
use sg13g2_a21oi_1  _349_
timestamp 1683973020
transform 1 0 9312 0 -1 27972
box -48 -56 528 834
use sg13g2_o21ai_1  _350_
timestamp 1685175443
transform 1 0 11232 0 1 26460
box -48 -56 538 834
use sg13g2_mux2_1  _351_
timestamp 1677247768
transform 1 0 11424 0 1 24948
box -48 -56 1008 834
use sg13g2_mux4_1  _352_
timestamp 1677257233
transform 1 0 13920 0 1 37044
box -48 -56 2064 834
use sg13g2_mux4_1  _353_
timestamp 1677257233
transform 1 0 16416 0 -1 38556
box -48 -56 2064 834
use sg13g2_nand3b_1  _354_
timestamp 1676573470
transform 1 0 17376 0 -1 40068
box -48 -56 720 834
use sg13g2_nor2b_1  _355_
timestamp 1685181386
transform 1 0 15936 0 1 38556
box -54 -56 528 834
use sg13g2_a21oi_1  _356_
timestamp 1683973020
transform 1 0 16896 0 -1 40068
box -48 -56 528 834
use sg13g2_o21ai_1  _357_
timestamp 1685175443
transform 1 0 18720 0 1 38556
box -48 -56 538 834
use sg13g2_mux2_1  _358_
timestamp 1677247768
transform 1 0 18432 0 -1 38556
box -48 -56 1008 834
use sg13g2_mux4_1  _359_
timestamp 1677257233
transform 1 0 13824 0 1 18900
box -48 -56 2064 834
use sg13g2_nor2b_1  _360_
timestamp 1685181386
transform -1 0 14688 0 -1 24948
box -54 -56 528 834
use sg13g2_a21oi_1  _361_
timestamp 1683973020
transform 1 0 14208 0 1 24948
box -48 -56 528 834
use sg13g2_nand3b_1  _362_
timestamp 1676573470
transform -1 0 15648 0 1 23436
box -48 -56 720 834
use sg13g2_o21ai_1  _363_
timestamp 1685175443
transform 1 0 14688 0 1 24948
box -48 -56 538 834
use sg13g2_mux4_1  _364_
timestamp 1677257233
transform 1 0 12960 0 1 23436
box -48 -56 2064 834
use sg13g2_mux2_1  _365_
timestamp 1677247768
transform 1 0 15072 0 -1 24948
box -48 -56 1008 834
use sg13g2_mux4_1  _366_
timestamp 1677257233
transform 1 0 5280 0 1 2268
box -48 -56 2064 834
use sg13g2_nand3_1  _367_
timestamp 1683988354
transform -1 0 4032 0 -1 18900
box -48 -56 528 834
use sg13g2_or2_1  _368_
timestamp 1684236171
transform 1 0 1824 0 1 18900
box -48 -56 528 834
use sg13g2_o21ai_1  _369_
timestamp 1685175443
transform -1 0 3456 0 1 17388
box -48 -56 538 834
use sg13g2_o21ai_1  _370_
timestamp 1685175443
transform 1 0 3072 0 -1 15876
box -48 -56 538 834
use sg13g2_mux4_1  _371_
timestamp 1677257233
transform 1 0 1536 0 -1 18900
box -48 -56 2064 834
use sg13g2_mux2_1  _372_
timestamp 1677247768
transform 1 0 3072 0 1 15876
box -48 -56 1008 834
use sg13g2_o21ai_1  _373_
timestamp 1685175443
transform 1 0 12000 0 -1 27972
box -48 -56 538 834
use sg13g2_a21o_1  _374_
timestamp 1677175127
transform -1 0 12288 0 1 27972
box -48 -56 720 834
use sg13g2_mux2_1  _375_
timestamp 1677247768
transform 1 0 11136 0 -1 29484
box -48 -56 1008 834
use sg13g2_a21oi_1  _376_
timestamp 1683973020
transform 1 0 12768 0 1 27972
box -48 -56 528 834
use sg13g2_mux4_1  _377_
timestamp 1677257233
transform 1 0 9312 0 1 27972
box -48 -56 2064 834
use sg13g2_nor2_1  _378_
timestamp 1676627187
transform 1 0 9984 0 1 29484
box -48 -56 432 834
use sg13g2_a21oi_1  _379_
timestamp 1683973020
transform 1 0 12288 0 1 27972
box -48 -56 528 834
use sg13g2_mux4_1  _380_
timestamp 1677257233
transform 1 0 15648 0 1 32508
box -48 -56 2064 834
use sg13g2_mux4_1  _381_
timestamp 1677257233
transform 1 0 15744 0 -1 32508
box -48 -56 2064 834
use sg13g2_mux2_1  _382_
timestamp 1677247768
transform 1 0 16992 0 -1 34020
box -48 -56 1008 834
use sg13g2_mux4_1  _383_
timestamp 1677257233
transform 1 0 16704 0 1 24948
box -48 -56 2064 834
use sg13g2_nand2b_1  _384_
timestamp 1676567195
transform 1 0 18720 0 1 26460
box -48 -56 528 834
use sg13g2_mux2_1  _385_
timestamp 1677247768
transform 1 0 18720 0 1 24948
box -48 -56 1008 834
use sg13g2_nand2b_1  _386_
timestamp 1676567195
transform 1 0 19680 0 1 24948
box -48 -56 528 834
use sg13g2_nand2_1  _387_
timestamp 1676557249
transform 1 0 18336 0 1 26460
box -48 -56 432 834
use sg13g2_and3_1  _388_
timestamp 1676971669
transform 1 0 18432 0 -1 24948
box -48 -56 720 834
use sg13g2_o21ai_1  _389_
timestamp 1685175443
transform 1 0 19104 0 -1 26460
box -48 -56 538 834
use sg13g2_o21ai_1  _390_
timestamp 1685175443
transform -1 0 19584 0 -1 24948
box -48 -56 538 834
use sg13g2_o21ai_1  _391_
timestamp 1685175443
transform -1 0 5856 0 1 20412
box -48 -56 538 834
use sg13g2_a21o_1  _392_
timestamp 1677175127
transform -1 0 7200 0 -1 20412
box -48 -56 720 834
use sg13g2_mux2_1  _393_
timestamp 1677247768
transform 1 0 6624 0 1 21924
box -48 -56 1008 834
use sg13g2_a21oi_1  _394_
timestamp 1683973020
transform -1 0 7968 0 1 20412
box -48 -56 528 834
use sg13g2_o21ai_1  _395_
timestamp 1685175443
transform -1 0 7008 0 -1 23436
box -48 -56 538 834
use sg13g2_a21o_1  _396_
timestamp 1677175127
transform -1 0 6528 0 1 20412
box -48 -56 720 834
use sg13g2_mux2_1  _397_
timestamp 1677247768
transform 1 0 6528 0 1 20412
box -48 -56 1008 834
use sg13g2_a21oi_1  _398_
timestamp 1683973020
transform 1 0 7200 0 -1 20412
box -48 -56 528 834
use sg13g2_a22oi_1  _399_
timestamp 1685173987
transform 1 0 6624 0 -1 21924
box -48 -56 624 834
use sg13g2_mux4_1  _400_
timestamp 1677257233
transform 1 0 7296 0 1 27972
box -48 -56 2064 834
use sg13g2_nand2b_1  _401_
timestamp 1676567195
transform 1 0 7296 0 -1 29484
box -48 -56 528 834
use sg13g2_a21oi_1  _402_
timestamp 1683973020
transform -1 0 9120 0 1 29484
box -48 -56 528 834
use sg13g2_nand2b_1  _403_
timestamp 1676567195
transform 1 0 8448 0 -1 30996
box -48 -56 528 834
use sg13g2_a21oi_1  _404_
timestamp 1683973020
transform 1 0 9120 0 1 29484
box -48 -56 528 834
use sg13g2_a221oi_1  _405_
timestamp 1685197497
transform 1 0 8448 0 -1 29484
box -48 -56 816 834
use sg13g2_a21o_1  _406_
timestamp 1677175127
transform 1 0 7776 0 -1 29484
box -48 -56 720 834
use sg13g2_mux4_1  _407_
timestamp 1677257233
transform 1 0 15168 0 1 35532
box -48 -56 2064 834
use sg13g2_mux4_1  _408_
timestamp 1677257233
transform 1 0 15264 0 -1 35532
box -48 -56 2064 834
use sg13g2_mux2_1  _409_
timestamp 1677247768
transform -1 0 20352 0 -1 38556
box -48 -56 1008 834
use sg13g2_nor2_1  _410_
timestamp 1676627187
transform 1 0 14688 0 -1 24948
box -48 -56 432 834
use sg13g2_o21ai_1  _411_
timestamp 1685175443
transform 1 0 15072 0 -1 27972
box -48 -56 538 834
use sg13g2_or2_1  _412_
timestamp 1684236171
transform -1 0 16320 0 1 26460
box -48 -56 528 834
use sg13g2_mux2_1  _413_
timestamp 1677247768
transform 1 0 14304 0 1 26460
box -48 -56 1008 834
use sg13g2_a21oi_1  _414_
timestamp 1683973020
transform 1 0 16320 0 1 26460
box -48 -56 528 834
use sg13g2_a21oi_1  _415_
timestamp 1683973020
transform -1 0 14208 0 1 24948
box -48 -56 528 834
use sg13g2_o21ai_1  _416_
timestamp 1685175443
transform 1 0 14112 0 -1 26460
box -48 -56 538 834
use sg13g2_mux2_1  _417_
timestamp 1677247768
transform 1 0 14592 0 -1 26460
box -48 -56 1008 834
use sg13g2_a21oi_1  _418_
timestamp 1683973020
transform -1 0 15648 0 1 24948
box -48 -56 528 834
use sg13g2_a22oi_1  _419_
timestamp 1685173987
transform 1 0 15264 0 1 26460
box -48 -56 624 834
use sg13g2_o21ai_1  _420_
timestamp 1685175443
transform -1 0 4896 0 -1 21924
box -48 -56 538 834
use sg13g2_a21o_1  _421_
timestamp 1677175127
transform 1 0 4224 0 1 21924
box -48 -56 720 834
use sg13g2_mux2_1  _422_
timestamp 1677247768
transform -1 0 4224 0 1 21924
box -48 -56 1008 834
use sg13g2_a21oi_1  _423_
timestamp 1683973020
transform -1 0 3936 0 1 20412
box -48 -56 528 834
use sg13g2_mux2_1  _424_
timestamp 1677247768
transform 1 0 2304 0 1 21924
box -48 -56 1008 834
use sg13g2_o21ai_1  _425_
timestamp 1685175443
transform 1 0 2880 0 1 20412
box -48 -56 538 834
use sg13g2_a21o_1  _426_
timestamp 1677175127
transform -1 0 3840 0 -1 21924
box -48 -56 720 834
use sg13g2_a21oi_1  _427_
timestamp 1683973020
transform -1 0 3744 0 -1 24948
box -48 -56 528 834
use sg13g2_a22oi_1  _428_
timestamp 1685173987
transform -1 0 4416 0 -1 21924
box -48 -56 624 834
use sg13g2_o21ai_1  _429_
timestamp 1685175443
transform 1 0 17760 0 -1 23436
box -48 -56 538 834
use sg13g2_nand2b_1  _430_
timestamp 1676567195
transform -1 0 17760 0 -1 23436
box -48 -56 528 834
use sg13g2_o21ai_1  _431_
timestamp 1685175443
transform 1 0 17280 0 1 23436
box -48 -56 538 834
use sg13g2_mux4_1  _432_
timestamp 1677257233
transform 1 0 2496 0 1 14364
box -48 -56 2064 834
use sg13g2_mux4_1  _433_
timestamp 1677257233
transform 1 0 15168 0 -1 12852
box -48 -56 2064 834
use sg13g2_mux4_1  _434_
timestamp 1677257233
transform 1 0 16704 0 1 17388
box -48 -56 2064 834
use sg13g2_mux4_1  _435_
timestamp 1677257233
transform 1 0 9024 0 -1 12852
box -48 -56 2064 834
use sg13g2_mux4_1  _436_
timestamp 1677257233
transform 1 0 3648 0 1 12852
box -48 -56 2064 834
use sg13g2_mux4_1  _437_
timestamp 1677257233
transform 1 0 15360 0 1 9828
box -48 -56 2064 834
use sg13g2_mux4_1  _438_
timestamp 1677257233
transform -1 0 17568 0 -1 14364
box -48 -56 2064 834
use sg13g2_mux4_1  _439_
timestamp 1677257233
transform -1 0 9120 0 -1 9828
box -48 -56 2064 834
use sg13g2_mux4_1  _440_
timestamp 1677257233
transform 1 0 6624 0 -1 14364
box -48 -56 2064 834
use sg13g2_mux4_1  _441_
timestamp 1677257233
transform 1 0 12864 0 1 12852
box -48 -56 2064 834
use sg13g2_mux4_1  _442_
timestamp 1677257233
transform 1 0 13440 0 1 14364
box -48 -56 2064 834
use sg13g2_mux4_1  _443_
timestamp 1677257233
transform 1 0 6624 0 1 11340
box -48 -56 2064 834
use sg13g2_mux4_1  _444_
timestamp 1677257233
transform -1 0 4800 0 1 3780
box -48 -56 2064 834
use sg13g2_mux4_1  _445_
timestamp 1677257233
transform 1 0 14976 0 1 8316
box -48 -56 2064 834
use sg13g2_mux4_1  _446_
timestamp 1677257233
transform 1 0 15840 0 1 6804
box -48 -56 2064 834
use sg13g2_mux4_1  _447_
timestamp 1677257233
transform 1 0 10944 0 -1 8316
box -48 -56 2064 834
use sg13g2_mux4_1  _448_
timestamp 1677257233
transform 1 0 2496 0 1 11340
box -48 -56 2064 834
use sg13g2_mux4_1  _449_
timestamp 1677257233
transform 1 0 14112 0 -1 11340
box -48 -56 2064 834
use sg13g2_mux4_1  _450_
timestamp 1677257233
transform 1 0 16128 0 -1 15876
box -48 -56 2064 834
use sg13g2_mux4_1  _451_
timestamp 1677257233
transform 1 0 8736 0 1 9828
box -48 -56 2064 834
use sg13g2_mux4_1  _452_
timestamp 1677257233
transform 1 0 3552 0 -1 9828
box -48 -56 2064 834
use sg13g2_mux4_1  _453_
timestamp 1677257233
transform -1 0 19968 0 1 9828
box -48 -56 2064 834
use sg13g2_mux4_1  _454_
timestamp 1677257233
transform 1 0 18144 0 1 14364
box -48 -56 2064 834
use sg13g2_mux4_1  _455_
timestamp 1677257233
transform 1 0 10848 0 -1 9828
box -48 -56 2064 834
use sg13g2_mux4_1  _456_
timestamp 1677257233
transform 1 0 3744 0 1 6804
box -48 -56 2064 834
use sg13g2_mux4_1  _457_
timestamp 1677257233
transform 1 0 18048 0 -1 8316
box -48 -56 2064 834
use sg13g2_mux4_1  _458_
timestamp 1677257233
transform 1 0 17856 0 1 5292
box -48 -56 2064 834
use sg13g2_mux4_1  _459_
timestamp 1677257233
transform 1 0 11136 0 -1 6804
box -48 -56 2064 834
use sg13g2_mux4_1  _460_
timestamp 1677257233
transform 1 0 3744 0 -1 5292
box -48 -56 2064 834
use sg13g2_mux4_1  _461_
timestamp 1677257233
transform 1 0 18048 0 1 3780
box -48 -56 2064 834
use sg13g2_mux4_1  _462_
timestamp 1677257233
transform 1 0 17856 0 -1 6804
box -48 -56 2064 834
use sg13g2_mux4_1  _463_
timestamp 1677257233
transform -1 0 10368 0 -1 6804
box -48 -56 2064 834
use sg13g2_mux4_1  _464_
timestamp 1677257233
transform 1 0 3072 0 1 9828
box -48 -56 2064 834
use sg13g2_mux4_1  _465_
timestamp 1677257233
transform 1 0 18240 0 1 11340
box -48 -56 2064 834
use sg13g2_mux4_1  _466_
timestamp 1677257233
transform -1 0 20352 0 -1 17388
box -48 -56 2064 834
use sg13g2_mux4_1  _467_
timestamp 1677257233
transform 1 0 11040 0 1 9828
box -48 -56 2064 834
use sg13g2_mux4_1  _468_
timestamp 1677257233
transform 1 0 2880 0 1 2268
box -48 -56 2064 834
use sg13g2_mux4_1  _469_
timestamp 1677257233
transform 1 0 14784 0 1 3780
box -48 -56 2064 834
use sg13g2_mux4_1  _470_
timestamp 1677257233
transform 1 0 18240 0 1 12852
box -48 -56 2064 834
use sg13g2_mux4_1  _471_
timestamp 1677257233
transform -1 0 10176 0 1 6804
box -48 -56 2064 834
use sg13g2_mux4_1  _472_
timestamp 1677257233
transform -1 0 4608 0 -1 6804
box -48 -56 2064 834
use sg13g2_mux4_1  _473_
timestamp 1677257233
transform -1 0 15840 0 1 6804
box -48 -56 2064 834
use sg13g2_mux4_1  _474_
timestamp 1677257233
transform 1 0 16512 0 -1 3780
box -48 -56 2064 834
use sg13g2_mux4_1  _475_
timestamp 1677257233
transform 1 0 11136 0 -1 3780
box -48 -56 2064 834
use sg13g2_mux4_1  _476_
timestamp 1677257233
transform 1 0 9984 0 1 3780
box -48 -56 2064 834
use sg13g2_mux4_1  _477_
timestamp 1677257233
transform 1 0 14688 0 -1 2268
box -48 -56 2064 834
use sg13g2_mux4_1  _478_
timestamp 1677257233
transform 1 0 13152 0 -1 5292
box -48 -56 2064 834
use sg13g2_mux4_1  _479_
timestamp 1677257233
transform 1 0 7200 0 1 3780
box -48 -56 2064 834
use sg13g2_mux4_1  _480_
timestamp 1677257233
transform 1 0 7008 0 1 17388
box -48 -56 2064 834
use sg13g2_mux4_1  _481_
timestamp 1677257233
transform 1 0 10848 0 -1 20412
box -48 -56 2064 834
use sg13g2_mux4_1  _482_
timestamp 1677257233
transform 1 0 9504 0 1 17388
box -48 -56 2064 834
use sg13g2_mux4_1  _483_
timestamp 1677257233
transform 1 0 8064 0 1 18900
box -48 -56 2064 834
use sg13g2_mux4_1  _484_
timestamp 1677257233
transform 1 0 8160 0 1 30996
box -48 -56 2064 834
use sg13g2_mux4_1  _485_
timestamp 1677257233
transform 1 0 10272 0 1 30996
box -48 -56 2064 834
use sg13g2_mux4_1  _486_
timestamp 1677257233
transform 1 0 10848 0 -1 21924
box -48 -56 2064 834
use sg13g2_mux4_1  _487_
timestamp 1677257233
transform 1 0 2112 0 1 24948
box -48 -56 2064 834
use sg13g2_nor3_1  _488_
timestamp 1676639442
transform 1 0 3744 0 -1 34020
box -48 -56 528 834
use sg13g2_nand2b_1  _489_
timestamp 1676567195
transform 1 0 5760 0 -1 32508
box -48 -56 528 834
use sg13g2_a221oi_1  _490_
timestamp 1685197497
transform 1 0 6048 0 1 32508
box -48 -56 816 834
use sg13g2_mux4_1  _491_
timestamp 1677257233
transform 1 0 5856 0 1 30996
box -48 -56 2064 834
use sg13g2_nor3_1  _492_
timestamp 1676639442
transform -1 0 12384 0 1 40068
box -48 -56 528 834
use sg13g2_nand2b_1  _493_
timestamp 1676567195
transform 1 0 12576 0 -1 40068
box -48 -56 528 834
use sg13g2_a221oi_1  _494_
timestamp 1685197497
transform 1 0 11808 0 -1 40068
box -48 -56 816 834
use sg13g2_mux4_1  _495_
timestamp 1677257233
transform 1 0 11136 0 1 35532
box -48 -56 2064 834
use sg13g2_nor3_1  _496_
timestamp 1676639442
transform 1 0 13920 0 -1 30996
box -48 -56 528 834
use sg13g2_nand2b_1  _497_
timestamp 1676567195
transform 1 0 15072 0 1 30996
box -48 -56 528 834
use sg13g2_a221oi_1  _498_
timestamp 1685197497
transform 1 0 14304 0 1 30996
box -48 -56 816 834
use sg13g2_mux4_1  _499_
timestamp 1677257233
transform 1 0 13824 0 -1 29484
box -48 -56 2064 834
use sg13g2_nor3_1  _500_
timestamp 1676639442
transform 1 0 4992 0 1 14364
box -48 -56 528 834
use sg13g2_nand2b_1  _501_
timestamp 1676567195
transform 1 0 5856 0 1 15876
box -48 -56 528 834
use sg13g2_a221oi_1  _502_
timestamp 1685197497
transform 1 0 5472 0 1 14364
box -48 -56 816 834
use sg13g2_mux4_1  _503_
timestamp 1677257233
transform 1 0 4704 0 -1 17388
box -48 -56 2064 834
use sg13g2_mux4_1  _504_
timestamp 1677257233
transform 1 0 2112 0 -1 30996
box -48 -56 2064 834
use sg13g2_mux4_1  _505_
timestamp 1677257233
transform 1 0 11520 0 -1 34020
box -48 -56 2064 834
use sg13g2_mux4_1  _506_
timestamp 1677257233
transform 1 0 1824 0 -1 40068
box -48 -56 2064 834
use sg13g2_mux4_1  _507_
timestamp 1677257233
transform 1 0 2112 0 1 37044
box -48 -56 2064 834
use sg13g2_mux4_1  _508_
timestamp 1677257233
transform 1 0 2208 0 1 34020
box -48 -56 2064 834
use sg13g2_mux4_1  _509_
timestamp 1677257233
transform -1 0 3936 0 1 32508
box -48 -56 2064 834
use sg13g2_mux4_1  _510_
timestamp 1677257233
transform 1 0 1728 0 1 35532
box -48 -56 2064 834
use sg13g2_mux4_1  _511_
timestamp 1677257233
transform 1 0 1248 0 1 27972
box -48 -56 2064 834
use sg13g2_mux4_1  _512_
timestamp 1677257233
transform 1 0 4608 0 -1 30996
box -48 -56 2064 834
use sg13g2_mux4_1  _513_
timestamp 1677257233
transform 1 0 11040 0 -1 37044
box -48 -56 2064 834
use sg13g2_mux4_1  _514_
timestamp 1677257233
transform 1 0 13632 0 1 29484
box -48 -56 2064 834
use sg13g2_mux4_1  _515_
timestamp 1677257233
transform 1 0 2880 0 1 23436
box -48 -56 2064 834
use sg13g2_dlhq_1  _516_
timestamp 1678805552
transform 1 0 1152 0 -1 23436
box -50 -56 1692 834
use sg13g2_dlhq_1  _517_
timestamp 1678805552
transform 1 0 2976 0 -1 23436
box -50 -56 1692 834
use sg13g2_dlhq_1  _518_
timestamp 1678805552
transform 1 0 12000 0 1 29484
box -50 -56 1692 834
use sg13g2_dlhq_1  _519_
timestamp 1678805552
transform 1 0 14400 0 -1 30996
box -50 -56 1692 834
use sg13g2_dlhq_1  _520_
timestamp 1678805552
transform 1 0 9504 0 1 35532
box -50 -56 1692 834
use sg13g2_dlhq_1  _521_
timestamp 1678805552
transform 1 0 11424 0 1 37044
box -50 -56 1692 834
use sg13g2_dlhq_1  _522_
timestamp 1678805552
transform 1 0 2592 0 1 30996
box -50 -56 1692 834
use sg13g2_dlhq_1  _523_
timestamp 1678805552
transform 1 0 4224 0 1 30996
box -50 -56 1692 834
use sg13g2_dlhq_1  _524_
timestamp 1678805552
transform -1 0 4896 0 -1 27972
box -50 -56 1692 834
use sg13g2_dlhq_1  _525_
timestamp 1678805552
transform 1 0 1248 0 1 29484
box -50 -56 1692 834
use sg13g2_dlhq_1  _526_
timestamp 1678805552
transform -1 0 5760 0 -1 38556
box -50 -56 1692 834
use sg13g2_dlhq_1  _527_
timestamp 1678805552
transform 1 0 2208 0 -1 41580
box -50 -56 1692 834
use sg13g2_dlhq_1  _528_
timestamp 1678805552
transform -1 0 3456 0 -1 35532
box -50 -56 1692 834
use sg13g2_dlhq_1  _529_
timestamp 1678805552
transform 1 0 1152 0 -1 37044
box -50 -56 1692 834
use sg13g2_dlhq_1  _530_
timestamp 1678805552
transform -1 0 5856 0 1 34020
box -50 -56 1692 834
use sg13g2_dlhq_1  _531_
timestamp 1678805552
transform 1 0 1152 0 -1 38556
box -50 -56 1692 834
use sg13g2_dlhq_1  _532_
timestamp 1678805552
transform -1 0 7872 0 -1 41580
box -50 -56 1692 834
use sg13g2_dlhq_1  _533_
timestamp 1678805552
transform -1 0 9504 0 -1 41580
box -50 -56 1692 834
use sg13g2_dlhq_1  _534_
timestamp 1678805552
transform -1 0 5184 0 1 40068
box -50 -56 1692 834
use sg13g2_dlhq_1  _535_
timestamp 1678805552
transform -1 0 5472 0 -1 41580
box -50 -56 1692 834
use sg13g2_dlhq_1  _536_
timestamp 1678805552
transform 1 0 11808 0 1 32508
box -50 -56 1692 834
use sg13g2_dlhq_1  _537_
timestamp 1678805552
transform 1 0 9888 0 -1 34020
box -50 -56 1692 834
use sg13g2_dlhq_1  _538_
timestamp 1678805552
transform 1 0 1152 0 -1 34020
box -50 -56 1692 834
use sg13g2_dlhq_1  _539_
timestamp 1678805552
transform 1 0 2016 0 -1 32508
box -50 -56 1692 834
use sg13g2_dlhq_1  _540_
timestamp 1678805552
transform 1 0 1152 0 -1 21924
box -50 -56 1692 834
use sg13g2_dlhq_1  _541_
timestamp 1678805552
transform 1 0 1152 0 1 23436
box -50 -56 1692 834
use sg13g2_dlhq_1  _542_
timestamp 1678805552
transform 1 0 1152 0 1 20412
box -50 -56 1692 834
use sg13g2_dlhq_1  _543_
timestamp 1678805552
transform 1 0 12480 0 -1 26460
box -50 -56 1692 834
use sg13g2_dlhq_1  _544_
timestamp 1678805552
transform 1 0 13440 0 -1 27972
box -50 -56 1692 834
use sg13g2_dlhq_1  _545_
timestamp 1678805552
transform 1 0 12288 0 1 26460
box -50 -56 1692 834
use sg13g2_dlhq_1  _546_
timestamp 1678805552
transform 1 0 13632 0 -1 35532
box -50 -56 1692 834
use sg13g2_dlhq_1  _547_
timestamp 1678805552
transform 1 0 15456 0 1 34020
box -50 -56 1692 834
use sg13g2_dlhq_1  _548_
timestamp 1678805552
transform 1 0 15072 0 -1 37044
box -50 -56 1692 834
use sg13g2_dlhq_1  _549_
timestamp 1678805552
transform 1 0 5664 0 1 27972
box -50 -56 1692 834
use sg13g2_dlhq_1  _550_
timestamp 1678805552
transform 1 0 6624 0 -1 27972
box -50 -56 1692 834
use sg13g2_dlhq_1  _551_
timestamp 1678805552
transform 1 0 6624 0 1 29484
box -50 -56 1692 834
use sg13g2_dlhq_1  _552_
timestamp 1678805552
transform 1 0 3072 0 -1 17388
box -50 -56 1692 834
use sg13g2_dlhq_1  _553_
timestamp 1678805552
transform 1 0 3744 0 1 17388
box -50 -56 1692 834
use sg13g2_dlhq_1  _554_
timestamp 1678805552
transform 1 0 12192 0 -1 29484
box -50 -56 1692 834
use sg13g2_dlhq_1  _555_
timestamp 1678805552
transform 1 0 14592 0 1 27972
box -50 -56 1692 834
use sg13g2_dlhq_1  _556_
timestamp 1678805552
transform 1 0 9408 0 -1 37044
box -50 -56 1692 834
use sg13g2_dlhq_1  _557_
timestamp 1678805552
transform 1 0 11808 0 -1 35532
box -50 -56 1692 834
use sg13g2_dlhq_1  _558_
timestamp 1678805552
transform 1 0 4128 0 -1 32508
box -50 -56 1692 834
use sg13g2_dlhq_1  _559_
timestamp 1678805552
transform 1 0 6240 0 -1 32508
box -50 -56 1692 834
use sg13g2_dlhq_1  _560_
timestamp 1678805552
transform 1 0 1152 0 1 26460
box -50 -56 1692 834
use sg13g2_dlhq_1  _561_
timestamp 1678805552
transform 1 0 1440 0 -1 26460
box -50 -56 1692 834
use sg13g2_dlhq_1  _562_
timestamp 1678805552
transform 1 0 9216 0 -1 21924
box -50 -56 1692 834
use sg13g2_dlhq_1  _563_
timestamp 1678805552
transform 1 0 11232 0 1 20412
box -50 -56 1692 834
use sg13g2_dlhq_1  _564_
timestamp 1678805552
transform 1 0 10752 0 -1 30996
box -50 -56 1692 834
use sg13g2_dlhq_1  _565_
timestamp 1678805552
transform 1 0 8928 0 -1 30996
box -50 -56 1692 834
use sg13g2_dlhq_1  _566_
timestamp 1678805552
transform 1 0 8640 0 -1 32508
box -50 -56 1692 834
use sg13g2_dlhq_1  _567_
timestamp 1678805552
transform 1 0 6912 0 1 32508
box -50 -56 1692 834
use sg13g2_dlhq_1  _568_
timestamp 1678805552
transform 1 0 8352 0 -1 18900
box -50 -56 1692 834
use sg13g2_dlhq_1  _569_
timestamp 1678805552
transform 1 0 6432 0 1 18900
box -50 -56 1692 834
use sg13g2_dlhq_1  _570_
timestamp 1678805552
transform 1 0 8256 0 -1 17388
box -50 -56 1692 834
use sg13g2_dlhq_1  _571_
timestamp 1678805552
transform 1 0 9984 0 -1 18900
box -50 -56 1692 834
use sg13g2_dlhq_1  _572_
timestamp 1678805552
transform 1 0 9216 0 -1 20412
box -50 -56 1692 834
use sg13g2_dlhq_1  _573_
timestamp 1678805552
transform 1 0 11040 0 1 18900
box -50 -56 1692 834
use sg13g2_dlhq_1  _574_
timestamp 1678805552
transform 1 0 7296 0 1 15876
box -50 -56 1692 834
use sg13g2_dlhq_1  _575_
timestamp 1678805552
transform 1 0 5376 0 1 17388
box -50 -56 1692 834
use sg13g2_dlhq_1  _576_
timestamp 1678805552
transform 1 0 4992 0 -1 21924
box -50 -56 1692 834
use sg13g2_dlhq_1  _577_
timestamp 1678805552
transform 1 0 5568 0 -1 18900
box -50 -56 1692 834
use sg13g2_dlhq_1  _578_
timestamp 1678805552
transform 1 0 4992 0 1 21924
box -50 -56 1692 834
use sg13g2_dlhq_1  _579_
timestamp 1678805552
transform 1 0 15840 0 -1 26460
box -50 -56 1692 834
use sg13g2_dlhq_1  _580_
timestamp 1678805552
transform 1 0 16512 0 -1 24948
box -50 -56 1692 834
use sg13g2_dlhq_1  _581_
timestamp 1678805552
transform 1 0 17472 0 -1 26460
box -50 -56 1692 834
use sg13g2_dlhq_1  _582_
timestamp 1678805552
transform 1 0 14016 0 1 32508
box -50 -56 1692 834
use sg13g2_dlhq_1  _583_
timestamp 1678805552
transform -1 0 19296 0 1 32508
box -50 -56 1692 834
use sg13g2_dlhq_1  _584_
timestamp 1678805552
transform 1 0 15360 0 -1 34020
box -50 -56 1692 834
use sg13g2_dlhq_1  _585_
timestamp 1678805552
transform -1 0 11040 0 -1 29484
box -50 -56 1692 834
use sg13g2_dlhq_1  _586_
timestamp 1678805552
transform 1 0 10368 0 1 29484
box -50 -56 1692 834
use sg13g2_dlhq_1  _587_
timestamp 1678805552
transform 1 0 10368 0 -1 27972
box -50 -56 1692 834
use sg13g2_dlhq_1  _588_
timestamp 1678805552
transform 1 0 5952 0 -1 3780
box -50 -56 1692 834
use sg13g2_dlhq_1  _589_
timestamp 1678805552
transform 1 0 7680 0 -1 3780
box -50 -56 1692 834
use sg13g2_dlhq_1  _590_
timestamp 1678805552
transform 1 0 11520 0 -1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _591_
timestamp 1678805552
transform 1 0 13152 0 1 3780
box -50 -56 1692 834
use sg13g2_dlhq_1  _592_
timestamp 1678805552
transform 1 0 12384 0 -1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _593_
timestamp 1678805552
transform 1 0 15360 0 1 756
box -50 -56 1692 834
use sg13g2_dlhq_1  _594_
timestamp 1678805552
transform 1 0 8256 0 -1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _595_
timestamp 1678805552
transform 1 0 9888 0 -1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _596_
timestamp 1678805552
transform 1 0 11808 0 1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _597_
timestamp 1678805552
transform 1 0 9504 0 -1 3780
box -50 -56 1692 834
use sg13g2_dlhq_1  _598_
timestamp 1678805552
transform 1 0 16896 0 1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _599_
timestamp 1678805552
transform 1 0 15264 0 1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _600_
timestamp 1678805552
transform -1 0 16800 0 -1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _601_
timestamp 1678805552
transform 1 0 13152 0 -1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _602_
timestamp 1678805552
transform -1 0 3744 0 1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _603_
timestamp 1678805552
transform 1 0 1152 0 1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _604_
timestamp 1678805552
transform 1 0 7680 0 -1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _605_
timestamp 1678805552
transform 1 0 6048 0 -1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _606_
timestamp 1678805552
transform 1 0 18624 0 -1 12852
box -50 -56 1692 834
use sg13g2_dlhq_1  _607_
timestamp 1678805552
transform 1 0 16608 0 1 12852
box -50 -56 1692 834
use sg13g2_dlhq_1  _608_
timestamp 1678805552
transform 1 0 15168 0 -1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _609_
timestamp 1678805552
transform 1 0 13440 0 -1 3780
box -50 -56 1692 834
use sg13g2_dlhq_1  _610_
timestamp 1678805552
transform 1 0 3168 0 1 756
box -50 -56 1692 834
use sg13g2_dlhq_1  _611_
timestamp 1678805552
transform 1 0 1344 0 -1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _612_
timestamp 1678805552
transform 1 0 10272 0 1 11340
box -50 -56 1692 834
use sg13g2_dlhq_1  _613_
timestamp 1678805552
transform 1 0 11520 0 -1 11340
box -50 -56 1692 834
use sg13g2_dlhq_1  _614_
timestamp 1678805552
transform 1 0 18720 0 1 15876
box -50 -56 1692 834
use sg13g2_dlhq_1  _615_
timestamp 1678805552
transform -1 0 20352 0 1 17388
box -50 -56 1692 834
use sg13g2_dlhq_1  _616_
timestamp 1678805552
transform 1 0 16992 0 -1 11340
box -50 -56 1692 834
use sg13g2_dlhq_1  _617_
timestamp 1678805552
transform 1 0 18624 0 -1 11340
box -50 -56 1692 834
use sg13g2_dlhq_1  _618_
timestamp 1678805552
transform 1 0 1440 0 1 9828
box -50 -56 1692 834
use sg13g2_dlhq_1  _619_
timestamp 1678805552
transform 1 0 3456 0 1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _620_
timestamp 1678805552
transform 1 0 6624 0 1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _621_
timestamp 1678805552
transform -1 0 9888 0 1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _622_
timestamp 1678805552
transform 1 0 16224 0 1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _623_
timestamp 1678805552
transform 1 0 18528 0 -1 3780
box -50 -56 1692 834
use sg13g2_dlhq_1  _624_
timestamp 1678805552
transform 1 0 16704 0 -1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _625_
timestamp 1678805552
transform 1 0 18432 0 -1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _626_
timestamp 1678805552
transform 1 0 2016 0 -1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _627_
timestamp 1678805552
transform 1 0 4224 0 -1 3780
box -50 -56 1692 834
use sg13g2_dlhq_1  _628_
timestamp 1678805552
transform 1 0 9888 0 1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _629_
timestamp 1678805552
transform 1 0 11616 0 1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _630_
timestamp 1678805552
transform 1 0 16800 0 -1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _631_
timestamp 1678805552
transform 1 0 18528 0 1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _632_
timestamp 1678805552
transform -1 0 19488 0 1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _633_
timestamp 1678805552
transform 1 0 18528 0 -1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _634_
timestamp 1678805552
transform 1 0 2112 0 -1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _635_
timestamp 1678805552
transform 1 0 4416 0 1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _636_
timestamp 1678805552
transform 1 0 9696 0 1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _637_
timestamp 1678805552
transform 1 0 11520 0 1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _638_
timestamp 1678805552
transform -1 0 19200 0 -1 14364
box -50 -56 1692 834
use sg13g2_dlhq_1  _639_
timestamp 1678805552
transform 1 0 18432 0 -1 15876
box -50 -56 1692 834
use sg13g2_dlhq_1  _640_
timestamp 1678805552
transform 1 0 17568 0 -1 9828
box -50 -56 1692 834
use sg13g2_dlhq_1  _641_
timestamp 1678805552
transform 1 0 18624 0 1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _642_
timestamp 1678805552
transform 1 0 1824 0 -1 9828
box -50 -56 1692 834
use sg13g2_dlhq_1  _643_
timestamp 1678805552
transform 1 0 4128 0 -1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _644_
timestamp 1678805552
transform 1 0 9120 0 -1 9828
box -50 -56 1692 834
use sg13g2_dlhq_1  _645_
timestamp 1678805552
transform 1 0 7104 0 1 9828
box -50 -56 1692 834
use sg13g2_dlhq_1  _646_
timestamp 1678805552
transform -1 0 18720 0 1 15876
box -50 -56 1692 834
use sg13g2_dlhq_1  _647_
timestamp 1678805552
transform 1 0 15456 0 1 15876
box -50 -56 1692 834
use sg13g2_dlhq_1  _648_
timestamp 1678805552
transform 1 0 14208 0 -1 9828
box -50 -56 1692 834
use sg13g2_dlhq_1  _649_
timestamp 1678805552
transform 1 0 13056 0 1 9828
box -50 -56 1692 834
use sg13g2_dlhq_1  _650_
timestamp 1678805552
transform 1 0 2400 0 -1 12852
box -50 -56 1692 834
use sg13g2_dlhq_1  _651_
timestamp 1678805552
transform 1 0 1152 0 -1 11340
box -50 -56 1692 834
use sg13g2_dlhq_1  _652_
timestamp 1678805552
transform 1 0 11520 0 1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _653_
timestamp 1678805552
transform 1 0 9312 0 -1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _654_
timestamp 1678805552
transform 1 0 15744 0 -1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _655_
timestamp 1678805552
transform 1 0 13920 0 1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _656_
timestamp 1678805552
transform -1 0 18624 0 1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _657_
timestamp 1678805552
transform 1 0 13536 0 -1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _658_
timestamp 1678805552
transform -1 0 4224 0 -1 3780
box -50 -56 1692 834
use sg13g2_dlhq_1  _659_
timestamp 1678805552
transform 1 0 1152 0 1 3780
box -50 -56 1692 834
use sg13g2_dlhq_1  _660_
timestamp 1678805552
transform 1 0 4992 0 1 11340
box -50 -56 1692 834
use sg13g2_dlhq_1  _661_
timestamp 1678805552
transform 1 0 7488 0 -1 11340
box -50 -56 1692 834
use sg13g2_dlhq_1  _662_
timestamp 1678805552
transform 1 0 12096 0 -1 14364
box -50 -56 1692 834
use sg13g2_dlhq_1  _663_
timestamp 1678805552
transform 1 0 13728 0 -1 14364
box -50 -56 1692 834
use sg13g2_dlhq_1  _664_
timestamp 1678805552
transform 1 0 11520 0 -1 12852
box -50 -56 1692 834
use sg13g2_dlhq_1  _665_
timestamp 1678805552
transform 1 0 13152 0 -1 12852
box -50 -56 1692 834
use sg13g2_dlhq_1  _666_
timestamp 1678805552
transform 1 0 4992 0 -1 14364
box -50 -56 1692 834
use sg13g2_dlhq_1  _667_
timestamp 1678805552
transform 1 0 6912 0 1 12852
box -50 -56 1692 834
use sg13g2_dlhq_1  _668_
timestamp 1678805552
transform -1 0 8832 0 1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _669_
timestamp 1678805552
transform 1 0 5568 0 1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _670_
timestamp 1678805552
transform -1 0 17472 0 1 14364
box -50 -56 1692 834
use sg13g2_dlhq_1  _671_
timestamp 1678805552
transform 1 0 14880 0 1 12852
box -50 -56 1692 834
use sg13g2_dlhq_1  _672_
timestamp 1678805552
transform 1 0 15936 0 -1 9828
box -50 -56 1692 834
use sg13g2_dlhq_1  _673_
timestamp 1678805552
transform 1 0 13344 0 1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _674_
timestamp 1678805552
transform 1 0 4032 0 -1 12852
box -50 -56 1692 834
use sg13g2_dlhq_1  _675_
timestamp 1678805552
transform 1 0 2016 0 1 12852
box -50 -56 1692 834
use sg13g2_dlhq_1  _676_
timestamp 1678805552
transform 1 0 9504 0 -1 11340
box -50 -56 1692 834
use sg13g2_dlhq_1  _677_
timestamp 1678805552
transform 1 0 7392 0 -1 12852
box -50 -56 1692 834
use sg13g2_dlhq_1  _678_
timestamp 1678805552
transform 1 0 17088 0 -1 18900
box -50 -56 1692 834
use sg13g2_dlhq_1  _679_
timestamp 1678805552
transform 1 0 15456 0 -1 17388
box -50 -56 1692 834
use sg13g2_dlhq_1  _680_
timestamp 1678805552
transform 1 0 15744 0 1 11340
box -50 -56 1692 834
use sg13g2_dlhq_1  _681_
timestamp 1678805552
transform 1 0 13824 0 1 11340
box -50 -56 1692 834
use sg13g2_dlhq_1  _682_
timestamp 1678805552
transform 1 0 2592 0 -1 14364
box -50 -56 1692 834
use sg13g2_dlhq_1  _683_
timestamp 1678805552
transform 1 0 1152 0 -1 15876
box -50 -56 1692 834
use sg13g2_dlhq_1  _684_
timestamp 1678805552
transform 1 0 1152 0 1 17388
box -50 -56 1692 834
use sg13g2_dlhq_1  _685_
timestamp 1678805552
transform 1 0 1248 0 -1 17388
box -50 -56 1692 834
use sg13g2_dlhq_1  _686_
timestamp 1678805552
transform 1 0 1440 0 1 15876
box -50 -56 1692 834
use sg13g2_dlhq_1  _687_
timestamp 1678805552
transform 1 0 12576 0 -1 24948
box -50 -56 1692 834
use sg13g2_dlhq_1  _688_
timestamp 1678805552
transform 1 0 11328 0 1 23436
box -50 -56 1692 834
use sg13g2_dlhq_1  _689_
timestamp 1678805552
transform 1 0 13824 0 -1 23436
box -50 -56 1692 834
use sg13g2_dlhq_1  _690_
timestamp 1678805552
transform 1 0 16416 0 1 38556
box -50 -56 1692 834
use sg13g2_dlhq_1  _691_
timestamp 1678805552
transform 1 0 16128 0 1 37044
box -50 -56 1692 834
use sg13g2_dlhq_1  _692_
timestamp 1678805552
transform -1 0 19968 0 -1 37044
box -50 -56 1692 834
use sg13g2_dlhq_1  _693_
timestamp 1678805552
transform 1 0 7008 0 1 26460
box -50 -56 1692 834
use sg13g2_dlhq_1  _694_
timestamp 1678805552
transform 1 0 8928 0 1 26460
box -50 -56 1692 834
use sg13g2_dlhq_1  _695_
timestamp 1678805552
transform 1 0 10752 0 -1 26460
box -50 -56 1692 834
use sg13g2_dlhq_1  _696_
timestamp 1678805552
transform 1 0 4896 0 -1 23436
box -50 -56 1692 834
use sg13g2_dlhq_1  _697_
timestamp 1678805552
transform 1 0 4704 0 -1 24948
box -50 -56 1692 834
use sg13g2_dlhq_1  _698_
timestamp 1678805552
transform 1 0 5952 0 1 24948
box -50 -56 1692 834
use sg13g2_dlhq_1  _699_
timestamp 1678805552
transform 1 0 17760 0 1 18900
box -50 -56 1692 834
use sg13g2_dlhq_1  _700_
timestamp 1678805552
transform 1 0 16416 0 -1 20412
box -50 -56 1692 834
use sg13g2_dlhq_1  _701_
timestamp 1678805552
transform 1 0 18624 0 -1 20412
box -50 -56 1692 834
use sg13g2_dlhq_1  _702_
timestamp 1678805552
transform 1 0 15648 0 1 29484
box -50 -56 1692 834
use sg13g2_dlhq_1  _703_
timestamp 1678805552
transform 1 0 17376 0 1 29484
box -50 -56 1692 834
use sg13g2_dlhq_1  _704_
timestamp 1678805552
transform 1 0 18720 0 -1 30996
box -50 -56 1692 834
use sg13g2_dlhq_1  _705_
timestamp 1678805552
transform 1 0 2016 0 -1 29484
box -50 -56 1692 834
use sg13g2_dlhq_1  _706_
timestamp 1678805552
transform 1 0 3456 0 1 29484
box -50 -56 1692 834
use sg13g2_dlhq_1  _707_
timestamp 1678805552
transform 1 0 3840 0 -1 29484
box -50 -56 1692 834
use sg13g2_dlhq_1  _708_
timestamp 1678805552
transform 1 0 1152 0 -1 20412
box -50 -56 1692 834
use sg13g2_dlhq_1  _709_
timestamp 1678805552
transform 1 0 2784 0 -1 20412
box -50 -56 1692 834
use sg13g2_dlhq_1  _710_
timestamp 1678805552
transform -1 0 5952 0 1 18900
box -50 -56 1692 834
use sg13g2_dlhq_1  _711_
timestamp 1678805552
transform 1 0 13248 0 1 20412
box -50 -56 1692 834
use sg13g2_dlhq_1  _712_
timestamp 1678805552
transform 1 0 12864 0 -1 21924
box -50 -56 1692 834
use sg13g2_dlhq_1  _713_
timestamp 1678805552
transform -1 0 16512 0 1 20412
box -50 -56 1692 834
use sg13g2_dlhq_1  _714_
timestamp 1678805552
transform 1 0 17952 0 1 35532
box -50 -56 1692 834
use sg13g2_dlhq_1  _715_
timestamp 1678805552
transform 1 0 18240 0 1 34020
box -50 -56 1692 834
use sg13g2_dlhq_1  _716_
timestamp 1678805552
transform 1 0 18240 0 -1 34020
box -50 -56 1692 834
use sg13g2_dlhq_1  _717_
timestamp 1678805552
transform 1 0 7584 0 1 24948
box -50 -56 1692 834
use sg13g2_dlhq_1  _718_
timestamp 1678805552
transform 1 0 9312 0 1 23436
box -50 -56 1692 834
use sg13g2_dlhq_1  _719_
timestamp 1678805552
transform 1 0 10560 0 -1 23436
box -50 -56 1692 834
use sg13g2_dlhq_1  _720_
timestamp 1678805552
transform -1 0 9120 0 -1 21924
box -50 -56 1692 834
use sg13g2_dlhq_1  _721_
timestamp 1678805552
transform 1 0 8064 0 -1 23436
box -50 -56 1692 834
use sg13g2_dlhq_1  _722_
timestamp 1678805552
transform 1 0 9888 0 1 21924
box -50 -56 1692 834
use sg13g2_dlhq_1  _723_
timestamp 1678805552
transform 1 0 16032 0 -1 21924
box -50 -56 1692 834
use sg13g2_dlhq_1  _724_
timestamp 1678805552
transform -1 0 19968 0 -1 23436
box -50 -56 1692 834
use sg13g2_dlhq_1  _725_
timestamp 1678805552
transform 1 0 18624 0 -1 21924
box -50 -56 1692 834
use sg13g2_dlhq_1  _726_
timestamp 1678805552
transform 1 0 16512 0 -1 29484
box -50 -56 1692 834
use sg13g2_dlhq_1  _727_
timestamp 1678805552
transform 1 0 15648 0 -1 27972
box -50 -56 1692 834
use sg13g2_dlhq_1  _728_
timestamp 1678805552
transform 1 0 18432 0 1 27972
box -50 -56 1692 834
use sg13g2_dlhq_1  _729_
timestamp 1678805552
transform 1 0 1632 0 -1 27972
box -50 -56 1692 834
use sg13g2_dlhq_1  _730_
timestamp 1678805552
transform 1 0 4032 0 1 26460
box -50 -56 1692 834
use sg13g2_dlhq_1  _731_
timestamp 1678805552
transform 1 0 4320 0 1 24948
box -50 -56 1692 834
use sg13g2_dlhq_1  _732_
timestamp 1678805552
transform 1 0 15648 0 1 23436
box -50 -56 1692 834
use sg13g2_dlhq_1  _733_
timestamp 1678805552
transform 1 0 15648 0 -1 23436
box -50 -56 1692 834
use sg13g2_dlhq_1  _734_
timestamp 1678805552
transform 1 0 5856 0 -1 34020
box -50 -56 1692 834
use sg13g2_dlhq_1  _735_
timestamp 1678805552
transform 1 0 5952 0 -1 35532
box -50 -56 1692 834
use sg13g2_dlhq_1  _736_
timestamp 1678805552
transform 1 0 6432 0 1 34020
box -50 -56 1692 834
use sg13g2_dlhq_1  _737_
timestamp 1678805552
transform -1 0 11616 0 1 34020
box -50 -56 1692 834
use sg13g2_dlhq_1  _738_
timestamp 1678805552
transform 1 0 2976 0 -1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _739_
timestamp 1678805552
transform 1 0 5280 0 1 756
box -50 -56 1692 834
use sg13g2_dlhq_1  _740_
timestamp 1678805552
transform 1 0 12864 0 -1 20412
box -50 -56 1692 834
use sg13g2_dlhq_1  _741_
timestamp 1678805552
transform -1 0 17472 0 1 18900
box -50 -56 1692 834
use sg13g2_dlhq_1  _742_
timestamp 1678805552
transform 1 0 12768 0 -1 38556
box -50 -56 1692 834
use sg13g2_dlhq_1  _743_
timestamp 1678805552
transform 1 0 14400 0 -1 38556
box -50 -56 1692 834
use sg13g2_dlhq_1  _744_
timestamp 1678805552
transform 1 0 8640 0 1 12852
box -50 -56 1692 834
use sg13g2_dlhq_1  _745_
timestamp 1678805552
transform -1 0 12960 0 -1 15876
box -50 -56 1692 834
use sg13g2_dlhq_1  _746_
timestamp 1678805552
transform 1 0 3840 0 -1 11340
box -50 -56 1692 834
use sg13g2_dlhq_1  _747_
timestamp 1678805552
transform 1 0 5472 0 1 9828
box -50 -56 1692 834
use sg13g2_dlhq_1  _748_
timestamp 1678805552
transform 1 0 11808 0 1 15876
box -50 -56 1692 834
use sg13g2_dlhq_1  _749_
timestamp 1678805552
transform 1 0 13824 0 -1 15876
box -50 -56 1692 834
use sg13g2_dlhq_1  _750_
timestamp 1678805552
transform 1 0 12480 0 1 40068
box -50 -56 1692 834
use sg13g2_dlhq_1  _751_
timestamp 1678805552
transform -1 0 16800 0 -1 40068
box -50 -56 1692 834
use sg13g2_dlhq_1  _752_
timestamp 1678805552
transform 1 0 5376 0 -1 15876
box -50 -56 1692 834
use sg13g2_dlhq_1  _753_
timestamp 1678805552
transform 1 0 6432 0 1 14364
box -50 -56 1692 834
use sg13g2_dlhq_1  _754_
timestamp 1678805552
transform 1 0 4608 0 -1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _755_
timestamp 1678805552
transform 1 0 5568 0 1 3780
box -50 -56 1692 834
use sg13g2_dlhq_1  _756_
timestamp 1678805552
transform 1 0 10368 0 -1 17388
box -50 -56 1692 834
use sg13g2_dlhq_1  _757_
timestamp 1678805552
transform 1 0 12000 0 -1 17388
box -50 -56 1692 834
use sg13g2_dlhq_1  _758_
timestamp 1678805552
transform 1 0 11904 0 -1 41580
box -50 -56 1692 834
use sg13g2_dlhq_1  _759_
timestamp 1678805552
transform -1 0 15744 0 1 40068
box -50 -56 1692 834
use sg13g2_dlhq_1  _760_
timestamp 1678805552
transform 1 0 8064 0 1 14364
box -50 -56 1692 834
use sg13g2_dlhq_1  _761_
timestamp 1678805552
transform 1 0 9696 0 -1 15876
box -50 -56 1692 834
use sg13g2_dlhq_1  _762_
timestamp 1678805552
transform 1 0 4608 0 -1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _763_
timestamp 1678805552
transform 1 0 6240 0 -1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _764_
timestamp 1678805552
transform 1 0 12000 0 -1 18900
box -50 -56 1692 834
use sg13g2_dlhq_1  _765_
timestamp 1678805552
transform 1 0 14112 0 1 17388
box -50 -56 1692 834
use sg13g2_dlhq_1  _766_
timestamp 1678805552
transform 1 0 11616 0 1 34020
box -50 -56 1692 834
use sg13g2_dlhq_1  _767_
timestamp 1678805552
transform 1 0 13536 0 -1 34020
box -50 -56 1692 834
use sg13g2_dlhq_1  _768_
timestamp 1678805552
transform 1 0 8640 0 1 11340
box -50 -56 1692 834
use sg13g2_dlhq_1  _769_
timestamp 1678805552
transform 1 0 10848 0 1 12852
box -50 -56 1692 834
use sg13g2_dlhq_1  _770_
timestamp 1678805552
transform 1 0 6336 0 -1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _771_
timestamp 1678805552
transform 1 0 8160 0 1 756
box -50 -56 1692 834
use sg13g2_dlhq_1  _772_
timestamp 1678805552
transform 1 0 2976 0 -1 37044
box -50 -56 1692 834
use sg13g2_dlhq_1  _773_
timestamp 1678805552
transform 1 0 4320 0 -1 35532
box -50 -56 1692 834
use sg13g2_dlhq_1  _774_
timestamp 1678805552
transform 1 0 8544 0 -1 38556
box -50 -56 1692 834
use sg13g2_dlhq_1  _775_
timestamp 1678805552
transform 1 0 6336 0 -1 38556
box -50 -56 1692 834
use sg13g2_dlhq_1  _776_
timestamp 1678805552
transform 1 0 6720 0 1 35532
box -50 -56 1692 834
use sg13g2_dlhq_1  _777_
timestamp 1678805552
transform 1 0 4608 0 -1 37044
box -50 -56 1692 834
use sg13g2_dlhq_1  _778_
timestamp 1678805552
transform 1 0 3264 0 1 38556
box -50 -56 1692 834
use sg13g2_dlhq_1  _779_
timestamp 1678805552
transform 1 0 3936 0 -1 40068
box -50 -56 1692 834
use sg13g2_dlhq_1  _780_
timestamp 1678805552
transform 1 0 1632 0 1 38556
box -50 -56 1692 834
use sg13g2_dlhq_1  _781_
timestamp 1678805552
transform 1 0 5952 0 1 40068
box -50 -56 1692 834
use sg13g2_dlhq_1  _782_
timestamp 1678805552
transform 1 0 8736 0 1 38556
box -50 -56 1692 834
use sg13g2_dlhq_1  _783_
timestamp 1678805552
transform 1 0 10560 0 -1 38556
box -50 -56 1692 834
use sg13g2_dlhq_1  _784_
timestamp 1678805552
transform 1 0 7104 0 1 38556
box -50 -56 1692 834
use sg13g2_dlhq_1  _785_
timestamp 1678805552
transform 1 0 8448 0 -1 40068
box -50 -56 1692 834
use sg13g2_dlhq_1  _786_
timestamp 1678805552
transform 1 0 4224 0 1 15876
box -50 -56 1692 834
use sg13g2_dlhq_1  _787_
timestamp 1678805552
transform 1 0 3744 0 -1 15876
box -50 -56 1692 834
use sg13g2_dlhq_1  _788_
timestamp 1678805552
transform 1 0 12672 0 1 30996
box -50 -56 1692 834
use sg13g2_dlhq_1  _789_
timestamp 1678805552
transform 1 0 12864 0 -1 32508
box -50 -56 1692 834
use sg13g2_dlhq_1  _790_
timestamp 1678805552
transform 1 0 10176 0 -1 40068
box -50 -56 1692 834
use sg13g2_dlhq_1  _791_
timestamp 1678805552
transform 1 0 10272 0 1 40068
box -50 -56 1692 834
use sg13g2_dlhq_1  _792_
timestamp 1678805552
transform 1 0 4320 0 1 32508
box -50 -56 1692 834
use sg13g2_dlhq_1  _793_
timestamp 1678805552
transform 1 0 4224 0 -1 34020
box -50 -56 1692 834
use sg13g2_buf_1  _794_
timestamp 1676381911
transform 1 0 19872 0 1 23436
box -48 -56 432 834
use sg13g2_buf_1  _795_
timestamp 1676381911
transform 1 0 19584 0 -1 24948
box -48 -56 432 834
use sg13g2_buf_1  _796_
timestamp 1676381911
transform 1 0 19968 0 -1 24948
box -48 -56 432 834
use sg13g2_buf_1  _797_
timestamp 1676381911
transform 1 0 19584 0 -1 26460
box -48 -56 432 834
use sg13g2_buf_1  _798_
timestamp 1676381911
transform 1 0 19968 0 -1 26460
box -48 -56 432 834
use sg13g2_buf_1  _799_
timestamp 1676381911
transform 1 0 19296 0 1 26460
box -48 -56 432 834
use sg13g2_buf_1  _800_
timestamp 1676381911
transform 1 0 19680 0 1 26460
box -48 -56 432 834
use sg13g2_buf_1  _801_
timestamp 1676381911
transform 1 0 18624 0 -1 27972
box -48 -56 432 834
use sg13g2_buf_1  _802_
timestamp 1676381911
transform 1 0 18624 0 -1 29484
box -48 -56 432 834
use sg13g2_buf_1  _803_
timestamp 1676381911
transform 1 0 19968 0 -1 29484
box -48 -56 432 834
use sg13g2_buf_1  _804_
timestamp 1676381911
transform 1 0 19968 0 1 30996
box -48 -56 432 834
use sg13g2_buf_1  _805_
timestamp 1676381911
transform 1 0 19584 0 1 30996
box -48 -56 432 834
use sg13g2_buf_1  _806_
timestamp 1676381911
transform 1 0 17568 0 1 30996
box -48 -56 432 834
use sg13g2_buf_1  _807_
timestamp 1676381911
transform 1 0 19872 0 -1 34020
box -48 -56 432 834
use sg13g2_buf_1  _808_
timestamp 1676381911
transform 1 0 19872 0 1 34020
box -48 -56 432 834
use sg13g2_buf_1  _809_
timestamp 1676381911
transform 1 0 19968 0 -1 32508
box -48 -56 432 834
use sg13g2_buf_1  _810_
timestamp 1676381911
transform 1 0 19584 0 -1 32508
box -48 -56 432 834
use sg13g2_buf_1  _811_
timestamp 1676381911
transform 1 0 19968 0 -1 37044
box -48 -56 432 834
use sg13g2_buf_1  _812_
timestamp 1676381911
transform 1 0 19200 0 -1 32508
box -48 -56 432 834
use sg13g2_buf_1  _813_
timestamp 1676381911
transform 1 0 19968 0 1 37044
box -48 -56 432 834
use sg13g2_buf_1  _814_
timestamp 1676381911
transform 1 0 19968 0 -1 40068
box -48 -56 432 834
use sg13g2_buf_1  _815_
timestamp 1676381911
transform 1 0 17376 0 1 34020
box -48 -56 432 834
use sg13g2_buf_1  _816_
timestamp 1676381911
transform 1 0 19968 0 1 38556
box -48 -56 432 834
use sg13g2_buf_1  _817_
timestamp 1676381911
transform 1 0 19584 0 1 38556
box -48 -56 432 834
use sg13g2_buf_1  _818_
timestamp 1676381911
transform 1 0 19392 0 -1 40068
box -48 -56 432 834
use sg13g2_buf_1  _819_
timestamp 1676381911
transform 1 0 16896 0 -1 37044
box -48 -56 432 834
use sg13g2_buf_1  _820_
timestamp 1676381911
transform 1 0 19776 0 1 40068
box -48 -56 432 834
use sg13g2_buf_1  _821_
timestamp 1676381911
transform 1 0 17664 0 1 40068
box -48 -56 432 834
use sg13g2_buf_1  _822_
timestamp 1676381911
transform 1 0 19296 0 1 40068
box -48 -56 432 834
use sg13g2_buf_1  _823_
timestamp 1676381911
transform 1 0 19200 0 1 38556
box -48 -56 432 834
use sg13g2_buf_1  _824_
timestamp 1676381911
transform 1 0 16032 0 -1 38556
box -48 -56 432 834
use sg13g2_buf_1  _825_
timestamp 1676381911
transform 1 0 19296 0 -1 41580
box -48 -56 432 834
use sg13g2_buf_1  _826_
timestamp 1676381911
transform 1 0 17184 0 1 35532
box -48 -56 432 834
use sg13g2_buf_1  _827_
timestamp 1676381911
transform -1 0 16512 0 1 40068
box -48 -56 432 834
use sg13g2_buf_1  _828_
timestamp 1676381911
transform -1 0 16896 0 1 40068
box -48 -56 432 834
use sg13g2_buf_1  _829_
timestamp 1676381911
transform -1 0 16416 0 -1 41580
box -48 -56 432 834
use sg13g2_buf_1  _830_
timestamp 1676381911
transform -1 0 17280 0 1 40068
box -48 -56 432 834
use sg13g2_buf_1  _831_
timestamp 1676381911
transform -1 0 16800 0 -1 18900
box -48 -56 432 834
use sg13g2_buf_1  _832_
timestamp 1676381911
transform 1 0 16032 0 -1 18900
box -48 -56 432 834
use sg13g2_buf_1  _833_
timestamp 1676381911
transform -1 0 17568 0 -1 41580
box -48 -56 432 834
use sg13g2_buf_1  _834_
timestamp 1676381911
transform -1 0 19200 0 1 40068
box -48 -56 432 834
use sg13g2_buf_1  _835_
timestamp 1676381911
transform -1 0 19200 0 -1 41580
box -48 -56 432 834
use sg13g2_buf_1  _836_
timestamp 1676381911
transform -1 0 18432 0 1 40068
box -48 -56 432 834
use sg13g2_buf_1  _837_
timestamp 1676381911
transform 1 0 17568 0 -1 41580
box -48 -56 432 834
use sg13g2_buf_1  _838_
timestamp 1676381911
transform -1 0 18816 0 1 40068
box -48 -56 432 834
use sg13g2_buf_1  _839_
timestamp 1676381911
transform -1 0 18432 0 -1 41580
box -48 -56 432 834
use sg13g2_buf_1  _840_
timestamp 1676381911
transform -1 0 20064 0 -1 41580
box -48 -56 432 834
use sg13g2_buf_1  _841_
timestamp 1676381911
transform -1 0 18816 0 -1 40068
box -48 -56 432 834
use sg13g2_buf_1  _842_
timestamp 1676381911
transform 1 0 17568 0 1 35532
box -48 -56 432 834
use sg13g2_buf_1  _843_
timestamp 1676381911
transform -1 0 19200 0 -1 40068
box -48 -56 432 834
use sg13g2_buf_1  _844_
timestamp 1676381911
transform 1 0 18048 0 1 37044
box -48 -56 432 834
use sg13g2_buf_1  _845_
timestamp 1676381911
transform 1 0 11520 0 -1 41580
box -48 -56 432 834
use sg13g2_buf_1  _846_
timestamp 1676381911
transform 1 0 18432 0 -1 41580
box -48 -56 432 834
use sg13g2_buf_1  _847_
timestamp 1676381911
transform 1 0 1440 0 1 34020
box -48 -56 432 834
use sg13g2_buf_1  _848_
timestamp 1676381911
transform -1 0 2208 0 1 34020
box -48 -56 432 834
use sg13g2_buf_1  _849_
timestamp 1676381911
transform 1 0 1440 0 -1 35532
box -48 -56 432 834
use sg13g2_buf_1  _850_
timestamp 1676381911
transform 1 0 1344 0 1 35532
box -48 -56 432 834
use sg13g2_buf_1  _851_
timestamp 1676381911
transform -1 0 10656 0 -1 41580
box -48 -56 432 834
use sg13g2_buf_1  _852_
timestamp 1676381911
transform -1 0 4128 0 -1 35532
box -48 -56 432 834
use sg13g2_buf_1  _853_
timestamp 1676381911
transform 1 0 1344 0 1 37044
box -48 -56 432 834
use sg13g2_buf_1  _854_
timestamp 1676381911
transform 1 0 1728 0 1 37044
box -48 -56 432 834
use sg13g2_buf_1  _855_
timestamp 1676381911
transform 1 0 2880 0 -1 38556
box -48 -56 432 834
use sg13g2_buf_1  _856_
timestamp 1676381911
transform 1 0 3264 0 -1 38556
box -48 -56 432 834
use sg13g2_buf_1  _857_
timestamp 1676381911
transform -1 0 13152 0 1 38556
box -48 -56 432 834
use sg13g2_buf_1  _858_
timestamp 1676381911
transform 1 0 1248 0 1 38556
box -48 -56 432 834
use sg13g2_buf_1  _859_
timestamp 1676381911
transform -1 0 7104 0 1 38556
box -48 -56 432 834
use sg13g2_buf_1  _860_
timestamp 1676381911
transform 1 0 1440 0 -1 40068
box -48 -56 432 834
use sg13g2_buf_1  _861_
timestamp 1676381911
transform 1 0 1440 0 1 40068
box -48 -56 432 834
use sg13g2_buf_1  _862_
timestamp 1676381911
transform -1 0 7296 0 1 37044
box -48 -56 432 834
use sg13g2_buf_1  _863_
timestamp 1676381911
transform -1 0 9888 0 -1 41580
box -48 -56 432 834
use sg13g2_buf_1  _864_
timestamp 1676381911
transform 1 0 1824 0 -1 41580
box -48 -56 432 834
use sg13g2_buf_1  _865_
timestamp 1676381911
transform 1 0 3744 0 -1 38556
box -48 -56 432 834
use sg13g2_buf_1  _866_
timestamp 1676381911
transform -1 0 5664 0 1 38556
box -48 -56 432 834
use sg13g2_buf_1  _867_
timestamp 1676381911
transform 1 0 2784 0 1 40068
box -48 -56 432 834
use sg13g2_buf_1  _868_
timestamp 1676381911
transform 1 0 4896 0 1 38556
box -48 -56 432 834
use sg13g2_buf_1  _869_
timestamp 1676381911
transform 1 0 3168 0 1 40068
box -48 -56 432 834
use sg13g2_buf_1  _870_
timestamp 1676381911
transform 1 0 5472 0 -1 41580
box -48 -56 432 834
use sg13g2_buf_1  _871_
timestamp 1676381911
transform 1 0 5952 0 1 38556
box -48 -56 432 834
use sg13g2_buf_1  _872_
timestamp 1676381911
transform 1 0 5184 0 1 40068
box -48 -56 432 834
use sg13g2_buf_1  _873_
timestamp 1676381911
transform 1 0 6336 0 1 38556
box -48 -56 432 834
use sg13g2_buf_1  _874_
timestamp 1676381911
transform -1 0 10272 0 -1 41580
box -48 -56 432 834
use sg13g2_buf_1  _875_
timestamp 1676381911
transform -1 0 8256 0 1 40068
box -48 -56 432 834
use sg13g2_buf_1  _876_
timestamp 1676381911
transform -1 0 7968 0 1 2268
box -48 -56 432 834
use sg13g2_buf_1  _877_
timestamp 1676381911
transform -1 0 8160 0 1 756
box -48 -56 432 834
use sg13g2_buf_1  _878_
timestamp 1676381911
transform -1 0 8352 0 1 2268
box -48 -56 432 834
use sg13g2_buf_1  _879_
timestamp 1676381911
transform 1 0 5568 0 1 40068
box -48 -56 432 834
use sg13g2_buf_1  _880_
timestamp 1676381911
transform -1 0 14112 0 -1 41580
box -48 -56 432 834
use sg13g2_buf_1  _881_
timestamp 1676381911
transform -1 0 17088 0 -1 41580
box -48 -56 432 834
use sg13g2_buf_1  _882_
timestamp 1676381911
transform 1 0 5856 0 -1 41580
box -48 -56 432 834
use sg13g2_buf_1  _883_
timestamp 1676381911
transform 1 0 7392 0 1 756
box -48 -56 432 834
use sg13g2_buf_1  _884_
timestamp 1676381911
transform -1 0 15552 0 -1 3780
box -48 -56 432 834
use sg13g2_buf_1  _885_
timestamp 1676381911
transform -1 0 13152 0 1 756
box -48 -56 432 834
use sg13g2_buf_1  _886_
timestamp 1676381911
transform 1 0 8352 0 1 2268
box -48 -56 432 834
use sg13g2_buf_1  _887_
timestamp 1676381911
transform 1 0 4800 0 1 756
box -48 -56 432 834
use sg13g2_buf_1  _888_
timestamp 1676381911
transform -1 0 12768 0 1 756
box -48 -56 432 834
use sg13g2_buf_1  _889_
timestamp 1676381911
transform -1 0 11136 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _890_
timestamp 1676381911
transform 1 0 9696 0 1 2268
box -48 -56 432 834
use sg13g2_buf_1  _891_
timestamp 1676381911
transform 1 0 9984 0 1 756
box -48 -56 432 834
use sg13g2_buf_1  _892_
timestamp 1676381911
transform -1 0 11232 0 1 2268
box -48 -56 432 834
use sg13g2_buf_1  _893_
timestamp 1676381911
transform -1 0 12384 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _894_
timestamp 1676381911
transform 1 0 9312 0 1 2268
box -48 -56 432 834
use sg13g2_buf_1  _895_
timestamp 1676381911
transform 1 0 10080 0 1 2268
box -48 -56 432 834
use sg13g2_buf_1  _896_
timestamp 1676381911
transform 1 0 10368 0 1 756
box -48 -56 432 834
use sg13g2_buf_1  _897_
timestamp 1676381911
transform 1 0 9984 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _898_
timestamp 1676381911
transform 1 0 10752 0 1 756
box -48 -56 432 834
use sg13g2_buf_1  _899_
timestamp 1676381911
transform 1 0 10368 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _900_
timestamp 1676381911
transform 1 0 11136 0 1 756
box -48 -56 432 834
use sg13g2_buf_1  _901_
timestamp 1676381911
transform 1 0 11136 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _902_
timestamp 1676381911
transform 1 0 11520 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _903_
timestamp 1676381911
transform -1 0 13536 0 1 756
box -48 -56 432 834
use sg13g2_buf_1  _904_
timestamp 1676381911
transform -1 0 13920 0 1 756
box -48 -56 432 834
use sg13g2_buf_1  _905_
timestamp 1676381911
transform -1 0 13824 0 1 2268
box -48 -56 432 834
use sg13g2_buf_1  _906_
timestamp 1676381911
transform -1 0 14784 0 1 756
box -48 -56 432 834
use sg13g2_buf_1  _907_
timestamp 1676381911
transform -1 0 14208 0 1 2268
box -48 -56 432 834
use sg13g2_buf_1  _908_
timestamp 1676381911
transform -1 0 14400 0 1 756
box -48 -56 432 834
use sg13g2_buf_1  _909_
timestamp 1676381911
transform -1 0 14592 0 1 2268
box -48 -56 432 834
use sg13g2_buf_1  _910_
timestamp 1676381911
transform -1 0 14976 0 1 2268
box -48 -56 432 834
use sg13g2_buf_1  _911_
timestamp 1676381911
transform -1 0 14688 0 -1 41580
box -48 -56 432 834
use sg13g2_buf_1  _912_
timestamp 1676381911
transform -1 0 15072 0 -1 41580
box -48 -56 432 834
use sg13g2_buf_1  _913_
timestamp 1676381911
transform -1 0 16128 0 1 40068
box -48 -56 432 834
use sg13g2_buf_1  _914_
timestamp 1676381911
transform -1 0 15456 0 -1 41580
box -48 -56 432 834
use sg13g2_buf_1  _915_
timestamp 1676381911
transform -1 0 15168 0 1 756
box -48 -56 432 834
use sg13g2_buf_1  _916_
timestamp 1676381911
transform -1 0 18528 0 1 756
box -48 -56 432 834
use sg13g2_buf_1  _917_
timestamp 1676381911
transform -1 0 17472 0 1 756
box -48 -56 432 834
use sg13g2_buf_1  _918_
timestamp 1676381911
transform 1 0 14304 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _919_
timestamp 1676381911
transform -1 0 16032 0 -1 41580
box -48 -56 432 834
use sg13g2_buf_1  _920_
timestamp 1676381911
transform -1 0 2976 0 1 756
box -48 -56 432 834
use sg13g2_buf_1  _921_
timestamp 1676381911
transform -1 0 5280 0 1 2268
box -48 -56 432 834
use sg13g2_buf_1  _922_
timestamp 1676381911
transform -1 0 3552 0 1 5292
box -48 -56 432 834
use sg13g2_buf_1  _923_
timestamp 1676381911
transform -1 0 5184 0 1 3780
box -48 -56 432 834
use sg13g2_buf_1  _924_
timestamp 1676381911
transform -1 0 2592 0 1 756
box -48 -56 432 834
use sg13g2_buf_1  _925_
timestamp 1676381911
transform -1 0 1824 0 1 756
box -48 -56 432 834
use sg13g2_buf_1  _926_
timestamp 1676381911
transform -1 0 2208 0 1 756
box -48 -56 432 834
use sg13g2_buf_1  _927_
timestamp 1676381911
transform -1 0 1824 0 1 2268
box -48 -56 432 834
use sg13g2_buf_1  _928_
timestamp 1676381911
transform -1 0 2208 0 1 2268
box -48 -56 432 834
use sg13g2_buf_1  _929_
timestamp 1676381911
transform -1 0 1824 0 -1 3780
box -48 -56 432 834
use sg13g2_buf_1  _930_
timestamp 1676381911
transform -1 0 2592 0 -1 3780
box -48 -56 432 834
use sg13g2_buf_1  _931_
timestamp 1676381911
transform -1 0 2592 0 1 2268
box -48 -56 432 834
use sg13g2_buf_1  _932_
timestamp 1676381911
transform -1 0 2208 0 -1 3780
box -48 -56 432 834
use sg13g2_buf_1  _933_
timestamp 1676381911
transform -1 0 18048 0 1 3780
box -48 -56 432 834
use sg13g2_buf_1  _934_
timestamp 1676381911
transform -1 0 20256 0 1 5292
box -48 -56 432 834
use sg13g2_buf_1  _935_
timestamp 1676381911
transform -1 0 2592 0 -1 6804
box -48 -56 432 834
use sg13g2_buf_1  _936_
timestamp 1676381911
transform -1 0 2016 0 -1 5292
box -48 -56 432 834
use sg13g2_buf_1  _937_
timestamp 1676381911
transform -1 0 19872 0 1 6804
box -48 -56 432 834
use sg13g2_buf_1  _938_
timestamp 1676381911
transform -1 0 17664 0 1 3780
box -48 -56 432 834
use sg13g2_buf_1  _939_
timestamp 1676381911
transform -1 0 3168 0 1 5292
box -48 -56 432 834
use sg13g2_buf_1  _940_
timestamp 1676381911
transform -1 0 1824 0 1 11340
box -48 -56 432 834
use sg13g2_buf_1  _941_
timestamp 1676381911
transform -1 0 2016 0 1 12852
box -48 -56 432 834
use sg13g2_buf_1  _942_
timestamp 1676381911
transform -1 0 1824 0 -1 12852
box -48 -56 432 834
use sg13g2_buf_1  _943_
timestamp 1676381911
transform -1 0 2208 0 -1 12852
box -48 -56 432 834
use sg13g2_buf_1  _944_
timestamp 1676381911
transform -1 0 2208 0 1 11340
box -48 -56 432 834
use sg13g2_buf_1  _945_
timestamp 1676381911
transform -1 0 2208 0 -1 14364
box -48 -56 432 834
use sg13g2_buf_1  _946_
timestamp 1676381911
transform -1 0 1632 0 1 12852
box -48 -56 432 834
use sg13g2_buf_1  _947_
timestamp 1676381911
transform -1 0 1824 0 -1 14364
box -48 -56 432 834
use sg13g2_buf_1  _948_
timestamp 1676381911
transform -1 0 2592 0 -1 14364
box -48 -56 432 834
use sg13g2_buf_1  _949_
timestamp 1676381911
transform -1 0 18336 0 -1 17388
box -48 -56 432 834
use sg13g2_buf_1  _950_
timestamp 1676381911
transform -1 0 1824 0 1 14364
box -48 -56 432 834
use sg13g2_buf_1  _951_
timestamp 1676381911
transform -1 0 2208 0 1 14364
box -48 -56 432 834
use sg13g2_buf_1  _952_
timestamp 1676381911
transform -1 0 1824 0 -1 6804
box -48 -56 432 834
use sg13g2_buf_1  _953_
timestamp 1676381911
transform -1 0 20256 0 -1 6804
box -48 -56 432 834
use sg13g2_buf_1  _954_
timestamp 1676381911
transform -1 0 2112 0 1 6804
box -48 -56 432 834
use sg13g2_buf_1  _955_
timestamp 1676381911
transform -1 0 1728 0 1 6804
box -48 -56 432 834
use sg13g2_buf_1  _956_
timestamp 1676381911
transform -1 0 2112 0 -1 8316
box -48 -56 432 834
use sg13g2_buf_1  _957_
timestamp 1676381911
transform -1 0 19680 0 -1 9828
box -48 -56 432 834
use sg13g2_buf_1  _958_
timestamp 1676381911
transform -1 0 1824 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  _959_
timestamp 1676381911
transform -1 0 2976 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  _960_
timestamp 1676381911
transform -1 0 2592 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  _961_
timestamp 1676381911
transform -1 0 17760 0 1 9828
box -48 -56 432 834
use sg13g2_buf_1  _962_
timestamp 1676381911
transform -1 0 1824 0 -1 9828
box -48 -56 432 834
use sg13g2_buf_1  _963_
timestamp 1676381911
transform -1 0 3168 0 -1 11340
box -48 -56 432 834
use sg13g2_buf_1  _964_
timestamp 1676381911
transform -1 0 1728 0 -1 8316
box -48 -56 432 834
use sg13g2_buf_1  _965_
timestamp 1676381911
transform -1 0 2208 0 -1 6804
box -48 -56 432 834
use sg13g2_buf_1  _966_
timestamp 1676381911
transform -1 0 2208 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  _967_
timestamp 1676381911
transform -1 0 1632 0 -1 5292
box -48 -56 432 834
use sg13g2_antennanp  ANTENNA_1
timestamp 1679999689
transform -1 0 16704 0 -1 41580
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_2
timestamp 1679999689
transform 1 0 18144 0 -1 40068
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_3
timestamp 1679999689
transform -1 0 17664 0 1 40068
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_4
timestamp 1679999689
transform 1 0 18432 0 1 38556
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_5
timestamp 1679999689
transform 1 0 18432 0 1 37044
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_6
timestamp 1679999689
transform 1 0 18048 0 1 38556
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_7
timestamp 1679999689
transform 1 0 7584 0 1 40068
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_8
timestamp 1679999689
transform -1 0 1440 0 -1 40068
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_9
timestamp 1679999689
transform 1 0 3936 0 1 35532
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_10
timestamp 1679999689
transform -1 0 1440 0 1 40068
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_11
timestamp 1679999689
transform 1 0 2112 0 1 40068
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_12
timestamp 1679999689
transform 1 0 7968 0 -1 38556
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_13
timestamp 1679999689
transform -1 0 1440 0 -1 41580
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_14
timestamp 1679999689
transform 1 0 4608 0 1 37044
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_15
timestamp 1679999689
transform 1 0 8160 0 -1 40068
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_16
timestamp 1679999689
transform -1 0 4608 0 1 37044
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_17
timestamp 1679999689
transform 1 0 5568 0 -1 40068
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_18
timestamp 1679999689
transform 1 0 14016 0 -1 2268
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_19
timestamp 1679999689
transform 1 0 17568 0 -1 35532
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_20
timestamp 1679999689
transform 1 0 18048 0 -1 37044
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_21
timestamp 1679999689
transform 1 0 8352 0 1 34020
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_22
timestamp 1679999689
transform 1 0 8256 0 -1 37044
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_23
timestamp 1679999689
transform 1 0 8352 0 1 35532
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_24
timestamp 1679999689
transform -1 0 8544 0 -1 38556
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_25
timestamp 1679999689
transform 1 0 1824 0 1 40068
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_26
timestamp 1679999689
transform 1 0 5856 0 -1 40068
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_27
timestamp 1679999689
transform -1 0 1824 0 -1 41580
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_28
timestamp 1679999689
transform 1 0 5952 0 -1 38556
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_29
timestamp 1679999689
transform -1 0 5952 0 1 38556
box -48 -56 336 834
use sg13g2_buf_8  clkbuf_0_UserCLK
timestamp 1676451365
transform 1 0 17952 0 -1 32508
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_1_0__f_UserCLK
timestamp 1676451365
transform 1 0 19008 0 1 29484
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_1_1__f_UserCLK
timestamp 1676451365
transform 1 0 18720 0 1 37044
box -48 -56 1296 834
use sg13g2_fill_2  FILLER_0_0
timestamp 1677580104
transform 1 0 1152 0 1 756
box -48 -56 240 834
use sg13g2_fill_1  FILLER_0_2
timestamp 1677579658
transform 1 0 1344 0 1 756
box -48 -56 144 834
use sg13g2_fill_2  FILLER_0_19
timestamp 1677580104
transform 1 0 2976 0 1 756
box -48 -56 240 834
use sg13g2_fill_1  FILLER_0_42
timestamp 1677579658
transform 1 0 5184 0 1 756
box -48 -56 144 834
use sg13g2_decap_4  FILLER_0_60
timestamp 1679577901
transform 1 0 6912 0 1 756
box -48 -56 432 834
use sg13g2_fill_1  FILLER_0_64
timestamp 1677579658
transform 1 0 7296 0 1 756
box -48 -56 144 834
use sg13g2_fill_2  FILLER_0_90
timestamp 1677580104
transform 1 0 9792 0 1 756
box -48 -56 240 834
use sg13g2_decap_8  FILLER_0_108
timestamp 1679581782
transform 1 0 11520 0 1 756
box -48 -56 720 834
use sg13g2_fill_2  FILLER_0_115
timestamp 1677580104
transform 1 0 12192 0 1 756
box -48 -56 240 834
use sg13g2_fill_1  FILLER_0_133
timestamp 1677579658
transform 1 0 13920 0 1 756
box -48 -56 144 834
use sg13g2_fill_2  FILLER_0_146
timestamp 1677580104
transform 1 0 15168 0 1 756
box -48 -56 240 834
use sg13g2_fill_1  FILLER_0_165
timestamp 1677579658
transform 1 0 16992 0 1 756
box -48 -56 144 834
use sg13g2_decap_8  FILLER_0_170
timestamp 1679581782
transform 1 0 17472 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_181
timestamp 1679581782
transform 1 0 18528 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_188
timestamp 1679581782
transform 1 0 19200 0 1 756
box -48 -56 720 834
use sg13g2_decap_4  FILLER_0_195
timestamp 1679577901
transform 1 0 19872 0 1 756
box -48 -56 432 834
use sg13g2_fill_1  FILLER_0_199
timestamp 1677579658
transform 1 0 20256 0 1 756
box -48 -56 144 834
use sg13g2_fill_2  FILLER_1_0
timestamp 1677580104
transform 1 0 1152 0 -1 2268
box -48 -56 240 834
use sg13g2_fill_1  FILLER_1_53
timestamp 1677579658
transform 1 0 6240 0 -1 2268
box -48 -56 144 834
use sg13g2_fill_1  FILLER_1_112
timestamp 1677579658
transform 1 0 11904 0 -1 2268
box -48 -56 144 834
use sg13g2_fill_1  FILLER_1_179
timestamp 1677579658
transform 1 0 18336 0 -1 2268
box -48 -56 144 834
use sg13g2_fill_2  FILLER_1_197
timestamp 1677580104
transform 1 0 20064 0 -1 2268
box -48 -56 240 834
use sg13g2_fill_1  FILLER_1_199
timestamp 1677579658
transform 1 0 20256 0 -1 2268
box -48 -56 144 834
use sg13g2_fill_2  FILLER_2_0
timestamp 1677580104
transform 1 0 1152 0 1 2268
box -48 -56 240 834
use sg13g2_fill_1  FILLER_2_2
timestamp 1677579658
transform 1 0 1344 0 1 2268
box -48 -56 144 834
use sg13g2_fill_2  FILLER_2_15
timestamp 1677580104
transform 1 0 2592 0 1 2268
box -48 -56 240 834
use sg13g2_fill_1  FILLER_2_17
timestamp 1677579658
transform 1 0 2784 0 1 2268
box -48 -56 144 834
use sg13g2_fill_2  FILLER_2_64
timestamp 1677580104
transform 1 0 7296 0 1 2268
box -48 -56 240 834
use sg13g2_fill_1  FILLER_2_66
timestamp 1677579658
transform 1 0 7488 0 1 2268
box -48 -56 144 834
use sg13g2_decap_4  FILLER_2_79
timestamp 1679577901
transform 1 0 8736 0 1 2268
box -48 -56 432 834
use sg13g2_fill_2  FILLER_2_83
timestamp 1677580104
transform 1 0 9120 0 1 2268
box -48 -56 240 834
use sg13g2_decap_4  FILLER_2_97
timestamp 1679577901
transform 1 0 10464 0 1 2268
box -48 -56 432 834
use sg13g2_decap_4  FILLER_2_105
timestamp 1679577901
transform 1 0 11232 0 1 2268
box -48 -56 432 834
use sg13g2_fill_2  FILLER_2_109
timestamp 1677580104
transform 1 0 11616 0 1 2268
box -48 -56 240 834
use sg13g2_fill_2  FILLER_2_144
timestamp 1677580104
transform 1 0 14976 0 1 2268
box -48 -56 240 834
use sg13g2_fill_1  FILLER_2_146
timestamp 1677579658
transform 1 0 15168 0 1 2268
box -48 -56 144 834
use sg13g2_fill_2  FILLER_2_198
timestamp 1677580104
transform 1 0 20160 0 1 2268
box -48 -56 240 834
use sg13g2_fill_2  FILLER_3_0
timestamp 1677580104
transform 1 0 1152 0 -1 3780
box -48 -56 240 834
use sg13g2_fill_1  FILLER_3_2
timestamp 1677579658
transform 1 0 1344 0 -1 3780
box -48 -56 144 834
use sg13g2_fill_1  FILLER_3_49
timestamp 1677579658
transform 1 0 5856 0 -1 3780
box -48 -56 144 834
use sg13g2_fill_1  FILLER_3_67
timestamp 1677579658
transform 1 0 7584 0 -1 3780
box -48 -56 144 834
use sg13g2_fill_2  FILLER_3_85
timestamp 1677580104
transform 1 0 9312 0 -1 3780
box -48 -56 240 834
use sg13g2_fill_2  FILLER_3_125
timestamp 1677580104
transform 1 0 13152 0 -1 3780
box -48 -56 240 834
use sg13g2_fill_1  FILLER_3_127
timestamp 1677579658
transform 1 0 13344 0 -1 3780
box -48 -56 144 834
use sg13g2_fill_1  FILLER_3_145
timestamp 1677579658
transform 1 0 15072 0 -1 3780
box -48 -56 144 834
use sg13g2_decap_8  FILLER_3_150
timestamp 1679581782
transform 1 0 15552 0 -1 3780
box -48 -56 720 834
use sg13g2_fill_2  FILLER_3_157
timestamp 1677580104
transform 1 0 16224 0 -1 3780
box -48 -56 240 834
use sg13g2_fill_1  FILLER_3_159
timestamp 1677579658
transform 1 0 16416 0 -1 3780
box -48 -56 144 834
use sg13g2_fill_2  FILLER_3_198
timestamp 1677580104
transform 1 0 20160 0 -1 3780
box -48 -56 240 834
use sg13g2_decap_4  FILLER_4_42
timestamp 1679577901
transform 1 0 5184 0 1 3780
box -48 -56 432 834
use sg13g2_decap_8  FILLER_4_84
timestamp 1679581782
transform 1 0 9216 0 1 3780
box -48 -56 720 834
use sg13g2_fill_1  FILLER_4_91
timestamp 1677579658
transform 1 0 9888 0 1 3780
box -48 -56 144 834
use sg13g2_decap_8  FILLER_4_113
timestamp 1679581782
transform 1 0 12000 0 1 3780
box -48 -56 720 834
use sg13g2_decap_4  FILLER_4_120
timestamp 1679577901
transform 1 0 12672 0 1 3780
box -48 -56 432 834
use sg13g2_fill_1  FILLER_4_124
timestamp 1677579658
transform 1 0 13056 0 1 3780
box -48 -56 144 834
use sg13g2_decap_4  FILLER_4_163
timestamp 1679577901
transform 1 0 16800 0 1 3780
box -48 -56 432 834
use sg13g2_fill_1  FILLER_4_167
timestamp 1677579658
transform 1 0 17184 0 1 3780
box -48 -56 144 834
use sg13g2_fill_2  FILLER_4_197
timestamp 1677580104
transform 1 0 20064 0 1 3780
box -48 -56 240 834
use sg13g2_fill_1  FILLER_4_199
timestamp 1677579658
transform 1 0 20256 0 1 3780
box -48 -56 144 834
use sg13g2_fill_1  FILLER_5_0
timestamp 1677579658
transform 1 0 1152 0 -1 5292
box -48 -56 144 834
use sg13g2_fill_1  FILLER_5_26
timestamp 1677579658
transform 1 0 3648 0 -1 5292
box -48 -56 144 834
use sg13g2_fill_1  FILLER_5_48
timestamp 1677579658
transform 1 0 5760 0 -1 5292
box -48 -56 144 834
use sg13g2_decap_4  FILLER_5_70
timestamp 1679577901
transform 1 0 7872 0 -1 5292
box -48 -56 432 834
use sg13g2_fill_1  FILLER_5_180
timestamp 1677579658
transform 1 0 18432 0 -1 5292
box -48 -56 144 834
use sg13g2_fill_2  FILLER_5_198
timestamp 1677580104
transform 1 0 20160 0 -1 5292
box -48 -56 240 834
use sg13g2_decap_8  FILLER_6_25
timestamp 1679581782
transform 1 0 3552 0 1 5292
box -48 -56 720 834
use sg13g2_fill_2  FILLER_6_32
timestamp 1677580104
transform 1 0 4224 0 1 5292
box -48 -56 240 834
use sg13g2_decap_4  FILLER_6_51
timestamp 1679577901
transform 1 0 6048 0 1 5292
box -48 -56 432 834
use sg13g2_fill_2  FILLER_6_55
timestamp 1677580104
transform 1 0 6432 0 1 5292
box -48 -56 240 834
use sg13g2_fill_1  FILLER_6_108
timestamp 1677579658
transform 1 0 11520 0 1 5292
box -48 -56 144 834
use sg13g2_decap_8  FILLER_6_126
timestamp 1679581782
transform 1 0 13248 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_150
timestamp 1679581782
transform 1 0 15552 0 1 5292
box -48 -56 720 834
use sg13g2_fill_1  FILLER_6_199
timestamp 1677579658
transform 1 0 20256 0 1 5292
box -48 -56 144 834
use sg13g2_fill_2  FILLER_7_0
timestamp 1677580104
transform 1 0 1152 0 -1 6804
box -48 -56 240 834
use sg13g2_fill_1  FILLER_7_2
timestamp 1677579658
transform 1 0 1344 0 -1 6804
box -48 -56 144 834
use sg13g2_decap_4  FILLER_7_70
timestamp 1679577901
transform 1 0 7872 0 -1 6804
box -48 -56 432 834
use sg13g2_fill_1  FILLER_7_74
timestamp 1677579658
transform 1 0 8256 0 -1 6804
box -48 -56 144 834
use sg13g2_decap_8  FILLER_7_96
timestamp 1679581782
transform 1 0 10368 0 -1 6804
box -48 -56 720 834
use sg13g2_fill_1  FILLER_7_103
timestamp 1677579658
transform 1 0 11040 0 -1 6804
box -48 -56 144 834
use sg13g2_decap_8  FILLER_7_142
timestamp 1679581782
transform 1 0 14784 0 -1 6804
box -48 -56 720 834
use sg13g2_fill_2  FILLER_7_149
timestamp 1677580104
transform 1 0 15456 0 -1 6804
box -48 -56 240 834
use sg13g2_fill_1  FILLER_7_151
timestamp 1677579658
transform 1 0 15648 0 -1 6804
box -48 -56 144 834
use sg13g2_decap_4  FILLER_7_169
timestamp 1679577901
transform 1 0 17376 0 -1 6804
box -48 -56 432 834
use sg13g2_fill_1  FILLER_7_173
timestamp 1677579658
transform 1 0 17760 0 -1 6804
box -48 -56 144 834
use sg13g2_fill_1  FILLER_7_199
timestamp 1677579658
transform 1 0 20256 0 -1 6804
box -48 -56 144 834
use sg13g2_fill_2  FILLER_8_0
timestamp 1677580104
transform 1 0 1152 0 1 6804
box -48 -56 240 834
use sg13g2_fill_2  FILLER_8_48
timestamp 1677580104
transform 1 0 5760 0 1 6804
box -48 -56 240 834
use sg13g2_fill_1  FILLER_8_50
timestamp 1677579658
transform 1 0 5952 0 1 6804
box -48 -56 144 834
use sg13g2_fill_1  FILLER_8_72
timestamp 1677579658
transform 1 0 8064 0 1 6804
box -48 -56 144 834
use sg13g2_decap_8  FILLER_8_94
timestamp 1679581782
transform 1 0 10176 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_101
timestamp 1679581782
transform 1 0 10848 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_125
timestamp 1679581782
transform 1 0 13152 0 1 6804
box -48 -56 720 834
use sg13g2_decap_4  FILLER_8_195
timestamp 1679577901
transform 1 0 19872 0 1 6804
box -48 -56 432 834
use sg13g2_fill_1  FILLER_8_199
timestamp 1677579658
transform 1 0 20256 0 1 6804
box -48 -56 144 834
use sg13g2_fill_2  FILLER_9_0
timestamp 1677580104
transform 1 0 1152 0 -1 8316
box -48 -56 240 834
use sg13g2_decap_4  FILLER_9_27
timestamp 1679577901
transform 1 0 3744 0 -1 8316
box -48 -56 432 834
use sg13g2_fill_2  FILLER_9_48
timestamp 1677580104
transform 1 0 5760 0 -1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_9_50
timestamp 1677579658
transform 1 0 5952 0 -1 8316
box -48 -56 144 834
use sg13g2_decap_4  FILLER_9_123
timestamp 1679577901
transform 1 0 12960 0 -1 8316
box -48 -56 432 834
use sg13g2_fill_2  FILLER_9_127
timestamp 1677580104
transform 1 0 13344 0 -1 8316
box -48 -56 240 834
use sg13g2_decap_8  FILLER_9_163
timestamp 1679581782
transform 1 0 16800 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_4  FILLER_9_170
timestamp 1679577901
transform 1 0 17472 0 -1 8316
box -48 -56 432 834
use sg13g2_fill_2  FILLER_9_174
timestamp 1677580104
transform 1 0 17856 0 -1 8316
box -48 -56 240 834
use sg13g2_fill_2  FILLER_9_197
timestamp 1677580104
transform 1 0 20064 0 -1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_9_199
timestamp 1677579658
transform 1 0 20256 0 -1 8316
box -48 -56 144 834
use sg13g2_fill_2  FILLER_10_0
timestamp 1677580104
transform 1 0 1152 0 1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_10_2
timestamp 1677579658
transform 1 0 1344 0 1 8316
box -48 -56 144 834
use sg13g2_decap_4  FILLER_10_19
timestamp 1679577901
transform 1 0 2976 0 1 8316
box -48 -56 432 834
use sg13g2_fill_1  FILLER_10_23
timestamp 1677579658
transform 1 0 3360 0 1 8316
box -48 -56 144 834
use sg13g2_decap_4  FILLER_10_41
timestamp 1679577901
transform 1 0 5088 0 1 8316
box -48 -56 432 834
use sg13g2_fill_1  FILLER_10_45
timestamp 1677579658
transform 1 0 5472 0 1 8316
box -48 -56 144 834
use sg13g2_decap_8  FILLER_10_80
timestamp 1679581782
transform 1 0 8832 0 1 8316
box -48 -56 720 834
use sg13g2_fill_2  FILLER_10_87
timestamp 1677580104
transform 1 0 9504 0 1 8316
box -48 -56 240 834
use sg13g2_fill_2  FILLER_10_106
timestamp 1677580104
transform 1 0 11328 0 1 8316
box -48 -56 240 834
use sg13g2_fill_2  FILLER_10_125
timestamp 1677580104
transform 1 0 13152 0 1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_10_199
timestamp 1677579658
transform 1 0 20256 0 1 8316
box -48 -56 144 834
use sg13g2_fill_2  FILLER_11_0
timestamp 1677580104
transform 1 0 1152 0 -1 9828
box -48 -56 240 834
use sg13g2_fill_1  FILLER_11_2
timestamp 1677579658
transform 1 0 1344 0 -1 9828
box -48 -56 144 834
use sg13g2_fill_1  FILLER_11_24
timestamp 1677579658
transform 1 0 3456 0 -1 9828
box -48 -56 144 834
use sg13g2_decap_8  FILLER_11_46
timestamp 1679581782
transform 1 0 5568 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_53
timestamp 1679581782
transform 1 0 6240 0 -1 9828
box -48 -56 720 834
use sg13g2_fill_2  FILLER_11_60
timestamp 1677580104
transform 1 0 6912 0 -1 9828
box -48 -56 240 834
use sg13g2_fill_1  FILLER_11_100
timestamp 1677579658
transform 1 0 10752 0 -1 9828
box -48 -56 144 834
use sg13g2_decap_8  FILLER_11_122
timestamp 1679581782
transform 1 0 12864 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_129
timestamp 1679581782
transform 1 0 13536 0 -1 9828
box -48 -56 720 834
use sg13g2_fill_1  FILLER_11_153
timestamp 1677579658
transform 1 0 15840 0 -1 9828
box -48 -56 144 834
use sg13g2_fill_1  FILLER_11_188
timestamp 1677579658
transform 1 0 19200 0 -1 9828
box -48 -56 144 834
use sg13g2_decap_8  FILLER_11_193
timestamp 1679581782
transform 1 0 19680 0 -1 9828
box -48 -56 720 834
use sg13g2_fill_2  FILLER_12_0
timestamp 1677580104
transform 1 0 1152 0 1 9828
box -48 -56 240 834
use sg13g2_fill_1  FILLER_12_2
timestamp 1677579658
transform 1 0 1344 0 1 9828
box -48 -56 144 834
use sg13g2_decap_4  FILLER_12_41
timestamp 1679577901
transform 1 0 5088 0 1 9828
box -48 -56 432 834
use sg13g2_fill_2  FILLER_12_100
timestamp 1677580104
transform 1 0 10752 0 1 9828
box -48 -56 240 834
use sg13g2_fill_1  FILLER_12_102
timestamp 1677579658
transform 1 0 10944 0 1 9828
box -48 -56 144 834
use sg13g2_decap_8  FILLER_12_141
timestamp 1679581782
transform 1 0 14688 0 1 9828
box -48 -56 720 834
use sg13g2_fill_2  FILLER_12_173
timestamp 1677580104
transform 1 0 17760 0 1 9828
box -48 -56 240 834
use sg13g2_decap_4  FILLER_12_196
timestamp 1679577901
transform 1 0 19968 0 1 9828
box -48 -56 432 834
use sg13g2_decap_8  FILLER_13_21
timestamp 1679581782
transform 1 0 3168 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_4  FILLER_13_83
timestamp 1679577901
transform 1 0 9120 0 -1 11340
box -48 -56 432 834
use sg13g2_decap_4  FILLER_13_104
timestamp 1679577901
transform 1 0 11136 0 -1 11340
box -48 -56 432 834
use sg13g2_decap_8  FILLER_13_125
timestamp 1679581782
transform 1 0 13152 0 -1 11340
box -48 -56 720 834
use sg13g2_fill_2  FILLER_13_132
timestamp 1677580104
transform 1 0 13824 0 -1 11340
box -48 -56 240 834
use sg13g2_fill_1  FILLER_13_134
timestamp 1677579658
transform 1 0 14016 0 -1 11340
box -48 -56 144 834
use sg13g2_decap_8  FILLER_13_156
timestamp 1679581782
transform 1 0 16128 0 -1 11340
box -48 -56 720 834
use sg13g2_fill_2  FILLER_13_163
timestamp 1677580104
transform 1 0 16800 0 -1 11340
box -48 -56 240 834
use sg13g2_fill_1  FILLER_13_199
timestamp 1677579658
transform 1 0 20256 0 -1 11340
box -48 -56 144 834
use sg13g2_fill_2  FILLER_14_0
timestamp 1677580104
transform 1 0 1152 0 1 11340
box -48 -56 240 834
use sg13g2_fill_1  FILLER_14_2
timestamp 1677579658
transform 1 0 1344 0 1 11340
box -48 -56 144 834
use sg13g2_fill_2  FILLER_14_11
timestamp 1677580104
transform 1 0 2208 0 1 11340
box -48 -56 240 834
use sg13g2_fill_1  FILLER_14_13
timestamp 1677579658
transform 1 0 2400 0 1 11340
box -48 -56 144 834
use sg13g2_decap_4  FILLER_14_35
timestamp 1679577901
transform 1 0 4512 0 1 11340
box -48 -56 432 834
use sg13g2_fill_1  FILLER_14_39
timestamp 1677579658
transform 1 0 4896 0 1 11340
box -48 -56 144 834
use sg13g2_decap_8  FILLER_14_112
timestamp 1679581782
transform 1 0 11904 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_119
timestamp 1679581782
transform 1 0 12576 0 1 11340
box -48 -56 720 834
use sg13g2_decap_4  FILLER_14_126
timestamp 1679577901
transform 1 0 13248 0 1 11340
box -48 -56 432 834
use sg13g2_fill_2  FILLER_14_130
timestamp 1677580104
transform 1 0 13632 0 1 11340
box -48 -56 240 834
use sg13g2_fill_2  FILLER_14_149
timestamp 1677580104
transform 1 0 15456 0 1 11340
box -48 -56 240 834
use sg13g2_fill_1  FILLER_14_151
timestamp 1677579658
transform 1 0 15648 0 1 11340
box -48 -56 144 834
use sg13g2_decap_8  FILLER_14_169
timestamp 1679581782
transform 1 0 17376 0 1 11340
box -48 -56 720 834
use sg13g2_fill_2  FILLER_14_176
timestamp 1677580104
transform 1 0 18048 0 1 11340
box -48 -56 240 834
use sg13g2_fill_1  FILLER_14_199
timestamp 1677579658
transform 1 0 20256 0 1 11340
box -48 -56 144 834
use sg13g2_fill_2  FILLER_15_0
timestamp 1677580104
transform 1 0 1152 0 -1 12852
box -48 -56 240 834
use sg13g2_fill_1  FILLER_15_2
timestamp 1677579658
transform 1 0 1344 0 -1 12852
box -48 -56 144 834
use sg13g2_fill_2  FILLER_15_11
timestamp 1677580104
transform 1 0 2208 0 -1 12852
box -48 -56 240 834
use sg13g2_decap_8  FILLER_15_47
timestamp 1679581782
transform 1 0 5664 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_54
timestamp 1679581782
transform 1 0 6336 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_4  FILLER_15_61
timestamp 1679577901
transform 1 0 7008 0 -1 12852
box -48 -56 432 834
use sg13g2_decap_4  FILLER_15_103
timestamp 1679577901
transform 1 0 11040 0 -1 12852
box -48 -56 432 834
use sg13g2_fill_1  FILLER_15_107
timestamp 1677579658
transform 1 0 11424 0 -1 12852
box -48 -56 144 834
use sg13g2_decap_4  FILLER_15_142
timestamp 1679577901
transform 1 0 14784 0 -1 12852
box -48 -56 432 834
use sg13g2_decap_8  FILLER_15_167
timestamp 1679581782
transform 1 0 17184 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_174
timestamp 1679581782
transform 1 0 17856 0 -1 12852
box -48 -56 720 834
use sg13g2_fill_1  FILLER_15_181
timestamp 1677579658
transform 1 0 18528 0 -1 12852
box -48 -56 144 834
use sg13g2_fill_1  FILLER_15_199
timestamp 1677579658
transform 1 0 20256 0 -1 12852
box -48 -56 144 834
use sg13g2_fill_1  FILLER_16_0
timestamp 1677579658
transform 1 0 1152 0 1 12852
box -48 -56 144 834
use sg13g2_decap_8  FILLER_16_47
timestamp 1679581782
transform 1 0 5664 0 1 12852
box -48 -56 720 834
use sg13g2_decap_4  FILLER_16_54
timestamp 1679577901
transform 1 0 6336 0 1 12852
box -48 -56 432 834
use sg13g2_fill_2  FILLER_16_58
timestamp 1677580104
transform 1 0 6720 0 1 12852
box -48 -56 240 834
use sg13g2_fill_1  FILLER_16_77
timestamp 1677579658
transform 1 0 8544 0 1 12852
box -48 -56 144 834
use sg13g2_decap_4  FILLER_16_95
timestamp 1679577901
transform 1 0 10272 0 1 12852
box -48 -56 432 834
use sg13g2_fill_2  FILLER_16_99
timestamp 1677580104
transform 1 0 10656 0 1 12852
box -48 -56 240 834
use sg13g2_decap_4  FILLER_16_118
timestamp 1679577901
transform 1 0 12480 0 1 12852
box -48 -56 432 834
use sg13g2_fill_1  FILLER_16_160
timestamp 1677579658
transform 1 0 16512 0 1 12852
box -48 -56 144 834
use sg13g2_fill_1  FILLER_16_199
timestamp 1677579658
transform 1 0 20256 0 1 12852
box -48 -56 144 834
use sg13g2_fill_2  FILLER_17_0
timestamp 1677580104
transform 1 0 1152 0 -1 14364
box -48 -56 240 834
use sg13g2_fill_1  FILLER_17_2
timestamp 1677579658
transform 1 0 1344 0 -1 14364
box -48 -56 144 834
use sg13g2_decap_8  FILLER_17_32
timestamp 1679581782
transform 1 0 4224 0 -1 14364
box -48 -56 720 834
use sg13g2_fill_1  FILLER_17_39
timestamp 1677579658
transform 1 0 4896 0 -1 14364
box -48 -56 144 834
use sg13g2_decap_8  FILLER_17_78
timestamp 1679581782
transform 1 0 8640 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_85
timestamp 1679581782
transform 1 0 9312 0 -1 14364
box -48 -56 720 834
use sg13g2_fill_1  FILLER_17_113
timestamp 1677579658
transform 1 0 12000 0 -1 14364
box -48 -56 144 834
use sg13g2_fill_2  FILLER_17_148
timestamp 1677580104
transform 1 0 15360 0 -1 14364
box -48 -56 240 834
use sg13g2_decap_8  FILLER_17_188
timestamp 1679581782
transform 1 0 19200 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_4  FILLER_17_195
timestamp 1679577901
transform 1 0 19872 0 -1 14364
box -48 -56 432 834
use sg13g2_fill_1  FILLER_17_199
timestamp 1677579658
transform 1 0 20256 0 -1 14364
box -48 -56 144 834
use sg13g2_fill_2  FILLER_18_0
timestamp 1677580104
transform 1 0 1152 0 1 14364
box -48 -56 240 834
use sg13g2_fill_1  FILLER_18_2
timestamp 1677579658
transform 1 0 1344 0 1 14364
box -48 -56 144 834
use sg13g2_fill_2  FILLER_18_11
timestamp 1677580104
transform 1 0 2208 0 1 14364
box -48 -56 240 834
use sg13g2_fill_1  FILLER_18_13
timestamp 1677579658
transform 1 0 2400 0 1 14364
box -48 -56 144 834
use sg13g2_decap_4  FILLER_18_35
timestamp 1679577901
transform 1 0 4512 0 1 14364
box -48 -56 432 834
use sg13g2_fill_1  FILLER_18_39
timestamp 1677579658
transform 1 0 4896 0 1 14364
box -48 -56 144 834
use sg13g2_fill_2  FILLER_18_53
timestamp 1677580104
transform 1 0 6240 0 1 14364
box -48 -56 240 834
use sg13g2_fill_2  FILLER_18_89
timestamp 1677580104
transform 1 0 9696 0 1 14364
box -48 -56 240 834
use sg13g2_fill_1  FILLER_18_91
timestamp 1677579658
transform 1 0 9888 0 1 14364
box -48 -56 144 834
use sg13g2_decap_8  FILLER_18_113
timestamp 1679581782
transform 1 0 12000 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_120
timestamp 1679581782
transform 1 0 12672 0 1 14364
box -48 -56 720 834
use sg13g2_fill_1  FILLER_18_127
timestamp 1677579658
transform 1 0 13344 0 1 14364
box -48 -56 144 834
use sg13g2_decap_4  FILLER_18_149
timestamp 1679577901
transform 1 0 15456 0 1 14364
box -48 -56 432 834
use sg13g2_decap_8  FILLER_18_170
timestamp 1679581782
transform 1 0 17472 0 1 14364
box -48 -56 720 834
use sg13g2_fill_2  FILLER_18_198
timestamp 1677580104
transform 1 0 20160 0 1 14364
box -48 -56 240 834
use sg13g2_fill_2  FILLER_19_17
timestamp 1677580104
transform 1 0 2784 0 -1 15876
box -48 -56 240 834
use sg13g2_fill_1  FILLER_19_19
timestamp 1677579658
transform 1 0 2976 0 -1 15876
box -48 -56 144 834
use sg13g2_fill_2  FILLER_19_25
timestamp 1677580104
transform 1 0 3552 0 -1 15876
box -48 -56 240 834
use sg13g2_decap_8  FILLER_19_82
timestamp 1679581782
transform 1 0 9024 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_123
timestamp 1679581782
transform 1 0 12960 0 -1 15876
box -48 -56 720 834
use sg13g2_fill_2  FILLER_19_130
timestamp 1677580104
transform 1 0 13632 0 -1 15876
box -48 -56 240 834
use sg13g2_decap_8  FILLER_19_149
timestamp 1679581782
transform 1 0 15456 0 -1 15876
box -48 -56 720 834
use sg13g2_fill_2  FILLER_19_177
timestamp 1677580104
transform 1 0 18144 0 -1 15876
box -48 -56 240 834
use sg13g2_fill_1  FILLER_19_179
timestamp 1677579658
transform 1 0 18336 0 -1 15876
box -48 -56 144 834
use sg13g2_fill_2  FILLER_19_197
timestamp 1677580104
transform 1 0 20064 0 -1 15876
box -48 -56 240 834
use sg13g2_fill_1  FILLER_19_199
timestamp 1677579658
transform 1 0 20256 0 -1 15876
box -48 -56 144 834
use sg13g2_fill_2  FILLER_20_0
timestamp 1677580104
transform 1 0 1152 0 1 15876
box -48 -56 240 834
use sg13g2_fill_1  FILLER_20_2
timestamp 1677579658
transform 1 0 1344 0 1 15876
box -48 -56 144 834
use sg13g2_fill_2  FILLER_20_30
timestamp 1677580104
transform 1 0 4032 0 1 15876
box -48 -56 240 834
use sg13g2_decap_8  FILLER_20_57
timestamp 1679581782
transform 1 0 6624 0 1 15876
box -48 -56 720 834
use sg13g2_decap_4  FILLER_20_81
timestamp 1679577901
transform 1 0 8928 0 1 15876
box -48 -56 432 834
use sg13g2_fill_1  FILLER_20_85
timestamp 1677579658
transform 1 0 9312 0 1 15876
box -48 -56 144 834
use sg13g2_decap_4  FILLER_20_107
timestamp 1679577901
transform 1 0 11424 0 1 15876
box -48 -56 432 834
use sg13g2_fill_1  FILLER_21_0
timestamp 1677579658
transform 1 0 1152 0 -1 17388
box -48 -56 144 834
use sg13g2_fill_2  FILLER_21_18
timestamp 1677580104
transform 1 0 2880 0 -1 17388
box -48 -56 240 834
use sg13g2_decap_8  FILLER_21_58
timestamp 1679581782
transform 1 0 6720 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_65
timestamp 1679581782
transform 1 0 7392 0 -1 17388
box -48 -56 720 834
use sg13g2_fill_2  FILLER_21_72
timestamp 1677580104
transform 1 0 8064 0 -1 17388
box -48 -56 240 834
use sg13g2_decap_4  FILLER_21_91
timestamp 1679577901
transform 1 0 9888 0 -1 17388
box -48 -56 432 834
use sg13g2_fill_1  FILLER_21_95
timestamp 1677579658
transform 1 0 10272 0 -1 17388
box -48 -56 144 834
use sg13g2_decap_8  FILLER_21_130
timestamp 1679581782
transform 1 0 13632 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_137
timestamp 1679581782
transform 1 0 14304 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_4  FILLER_21_144
timestamp 1679577901
transform 1 0 14976 0 -1 17388
box -48 -56 432 834
use sg13g2_fill_1  FILLER_21_148
timestamp 1677579658
transform 1 0 15360 0 -1 17388
box -48 -56 144 834
use sg13g2_decap_8  FILLER_21_166
timestamp 1679581782
transform 1 0 17088 0 -1 17388
box -48 -56 720 834
use sg13g2_fill_2  FILLER_21_173
timestamp 1677580104
transform 1 0 17760 0 -1 17388
box -48 -56 240 834
use sg13g2_fill_2  FILLER_22_17
timestamp 1677580104
transform 1 0 2784 0 1 17388
box -48 -56 240 834
use sg13g2_decap_4  FILLER_22_82
timestamp 1679577901
transform 1 0 9024 0 1 17388
box -48 -56 432 834
use sg13g2_fill_1  FILLER_22_86
timestamp 1677579658
transform 1 0 9408 0 1 17388
box -48 -56 144 834
use sg13g2_decap_4  FILLER_22_108
timestamp 1679577901
transform 1 0 11520 0 1 17388
box -48 -56 432 834
use sg13g2_fill_2  FILLER_22_133
timestamp 1677580104
transform 1 0 13920 0 1 17388
box -48 -56 240 834
use sg13g2_decap_8  FILLER_22_152
timestamp 1679581782
transform 1 0 15744 0 1 17388
box -48 -56 720 834
use sg13g2_fill_2  FILLER_22_159
timestamp 1677580104
transform 1 0 16416 0 1 17388
box -48 -56 240 834
use sg13g2_fill_1  FILLER_22_161
timestamp 1677579658
transform 1 0 16608 0 1 17388
box -48 -56 144 834
use sg13g2_decap_4  FILLER_23_0
timestamp 1679577901
transform 1 0 1152 0 -1 18900
box -48 -56 432 834
use sg13g2_decap_4  FILLER_23_40
timestamp 1679577901
transform 1 0 4992 0 -1 18900
box -48 -56 432 834
use sg13g2_fill_2  FILLER_23_44
timestamp 1677580104
transform 1 0 5376 0 -1 18900
box -48 -56 240 834
use sg13g2_decap_8  FILLER_23_63
timestamp 1679581782
transform 1 0 7200 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_4  FILLER_23_70
timestamp 1679577901
transform 1 0 7872 0 -1 18900
box -48 -56 432 834
use sg13g2_fill_1  FILLER_23_74
timestamp 1677579658
transform 1 0 8256 0 -1 18900
box -48 -56 144 834
use sg13g2_decap_4  FILLER_23_109
timestamp 1679577901
transform 1 0 11616 0 -1 18900
box -48 -56 432 834
use sg13g2_decap_4  FILLER_23_151
timestamp 1679577901
transform 1 0 15648 0 -1 18900
box -48 -56 432 834
use sg13g2_fill_2  FILLER_23_163
timestamp 1677580104
transform 1 0 16800 0 -1 18900
box -48 -56 240 834
use sg13g2_fill_1  FILLER_23_165
timestamp 1677579658
transform 1 0 16992 0 -1 18900
box -48 -56 144 834
use sg13g2_decap_8  FILLER_23_188
timestamp 1679581782
transform 1 0 19200 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_4  FILLER_23_195
timestamp 1679577901
transform 1 0 19872 0 -1 18900
box -48 -56 432 834
use sg13g2_fill_1  FILLER_23_199
timestamp 1677579658
transform 1 0 20256 0 -1 18900
box -48 -56 144 834
use sg13g2_decap_8  FILLER_24_0
timestamp 1679581782
transform 1 0 1152 0 1 18900
box -48 -56 720 834
use sg13g2_decap_4  FILLER_24_50
timestamp 1679577901
transform 1 0 5952 0 1 18900
box -48 -56 432 834
use sg13g2_fill_1  FILLER_24_54
timestamp 1677579658
transform 1 0 6336 0 1 18900
box -48 -56 144 834
use sg13g2_decap_8  FILLER_24_93
timestamp 1679581782
transform 1 0 10080 0 1 18900
box -48 -56 720 834
use sg13g2_fill_2  FILLER_24_100
timestamp 1677580104
transform 1 0 10752 0 1 18900
box -48 -56 240 834
use sg13g2_fill_1  FILLER_24_102
timestamp 1677579658
transform 1 0 10944 0 1 18900
box -48 -56 144 834
use sg13g2_decap_8  FILLER_24_120
timestamp 1679581782
transform 1 0 12672 0 1 18900
box -48 -56 720 834
use sg13g2_decap_4  FILLER_24_127
timestamp 1679577901
transform 1 0 13344 0 1 18900
box -48 -56 432 834
use sg13g2_fill_1  FILLER_24_131
timestamp 1677579658
transform 1 0 13728 0 1 18900
box -48 -56 144 834
use sg13g2_fill_2  FILLER_24_170
timestamp 1677580104
transform 1 0 17472 0 1 18900
box -48 -56 240 834
use sg13g2_fill_1  FILLER_24_172
timestamp 1677579658
transform 1 0 17664 0 1 18900
box -48 -56 144 834
use sg13g2_fill_1  FILLER_25_37
timestamp 1677579658
transform 1 0 4704 0 -1 20412
box -48 -56 144 834
use sg13g2_fill_2  FILLER_25_51
timestamp 1677580104
transform 1 0 6048 0 -1 20412
box -48 -56 240 834
use sg13g2_decap_8  FILLER_25_71
timestamp 1679581782
transform 1 0 7968 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_4  FILLER_25_78
timestamp 1679577901
transform 1 0 8640 0 -1 20412
box -48 -56 432 834
use sg13g2_fill_2  FILLER_25_82
timestamp 1677580104
transform 1 0 9024 0 -1 20412
box -48 -56 240 834
use sg13g2_decap_4  FILLER_25_139
timestamp 1679577901
transform 1 0 14496 0 -1 20412
box -48 -56 432 834
use sg13g2_decap_8  FILLER_25_148
timestamp 1679581782
transform 1 0 15360 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_4  FILLER_25_155
timestamp 1679577901
transform 1 0 16032 0 -1 20412
box -48 -56 432 834
use sg13g2_fill_1  FILLER_25_181
timestamp 1677579658
transform 1 0 18528 0 -1 20412
box -48 -56 144 834
use sg13g2_fill_1  FILLER_25_199
timestamp 1677579658
transform 1 0 20256 0 -1 20412
box -48 -56 144 834
use sg13g2_fill_1  FILLER_26_17
timestamp 1677579658
transform 1 0 2784 0 1 20412
box -48 -56 144 834
use sg13g2_fill_1  FILLER_26_23
timestamp 1677579658
transform 1 0 3360 0 1 20412
box -48 -56 144 834
use sg13g2_fill_2  FILLER_26_42
timestamp 1677580104
transform 1 0 5184 0 1 20412
box -48 -56 240 834
use sg13g2_decap_8  FILLER_26_71
timestamp 1679581782
transform 1 0 7968 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_78
timestamp 1679581782
transform 1 0 8640 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_90
timestamp 1679581782
transform 1 0 9792 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_97
timestamp 1679581782
transform 1 0 10464 0 1 20412
box -48 -56 720 834
use sg13g2_fill_1  FILLER_26_104
timestamp 1677579658
transform 1 0 11136 0 1 20412
box -48 -56 144 834
use sg13g2_decap_4  FILLER_26_122
timestamp 1679577901
transform 1 0 12864 0 1 20412
box -48 -56 432 834
use sg13g2_decap_8  FILLER_26_160
timestamp 1679581782
transform 1 0 16512 0 1 20412
box -48 -56 720 834
use sg13g2_fill_1  FILLER_27_17
timestamp 1677579658
transform 1 0 2784 0 -1 21924
box -48 -56 144 834
use sg13g2_fill_1  FILLER_27_39
timestamp 1677579658
transform 1 0 4896 0 -1 21924
box -48 -56 144 834
use sg13g2_fill_1  FILLER_27_83
timestamp 1677579658
transform 1 0 9120 0 -1 21924
box -48 -56 144 834
use sg13g2_fill_1  FILLER_27_144
timestamp 1677579658
transform 1 0 14976 0 -1 21924
box -48 -56 144 834
use sg13g2_decap_4  FILLER_27_172
timestamp 1679577901
transform 1 0 17664 0 -1 21924
box -48 -56 432 834
use sg13g2_fill_1  FILLER_27_181
timestamp 1677579658
transform 1 0 18528 0 -1 21924
box -48 -56 144 834
use sg13g2_fill_1  FILLER_27_199
timestamp 1677579658
transform 1 0 20256 0 -1 21924
box -48 -56 144 834
use sg13g2_decap_8  FILLER_28_0
timestamp 1679581782
transform 1 0 1152 0 1 21924
box -48 -56 720 834
use sg13g2_decap_4  FILLER_28_7
timestamp 1679577901
transform 1 0 1824 0 1 21924
box -48 -56 432 834
use sg13g2_fill_1  FILLER_28_11
timestamp 1677579658
transform 1 0 2208 0 1 21924
box -48 -56 144 834
use sg13g2_fill_1  FILLER_28_39
timestamp 1677579658
transform 1 0 4896 0 1 21924
box -48 -56 144 834
use sg13g2_fill_2  FILLER_28_67
timestamp 1677580104
transform 1 0 7584 0 1 21924
box -48 -56 240 834
use sg13g2_fill_1  FILLER_28_69
timestamp 1677579658
transform 1 0 7776 0 1 21924
box -48 -56 144 834
use sg13g2_decap_4  FILLER_28_118
timestamp 1679577901
transform 1 0 12480 0 1 21924
box -48 -56 432 834
use sg13g2_fill_2  FILLER_28_122
timestamp 1677580104
transform 1 0 12864 0 1 21924
box -48 -56 240 834
use sg13g2_decap_8  FILLER_28_157
timestamp 1679581782
transform 1 0 16224 0 1 21924
box -48 -56 720 834
use sg13g2_fill_1  FILLER_28_164
timestamp 1677579658
transform 1 0 16896 0 1 21924
box -48 -56 144 834
use sg13g2_decap_4  FILLER_28_196
timestamp 1679577901
transform 1 0 19968 0 1 21924
box -48 -56 432 834
use sg13g2_fill_2  FILLER_29_17
timestamp 1677580104
transform 1 0 2784 0 -1 23436
box -48 -56 240 834
use sg13g2_fill_1  FILLER_29_61
timestamp 1677579658
transform 1 0 7008 0 -1 23436
box -48 -56 144 834
use sg13g2_fill_2  FILLER_29_96
timestamp 1677580104
transform 1 0 10368 0 -1 23436
box -48 -56 240 834
use sg13g2_decap_8  FILLER_29_115
timestamp 1679581782
transform 1 0 12192 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_122
timestamp 1679581782
transform 1 0 12864 0 -1 23436
box -48 -56 720 834
use sg13g2_fill_2  FILLER_29_129
timestamp 1677580104
transform 1 0 13536 0 -1 23436
box -48 -56 240 834
use sg13g2_fill_1  FILLER_29_131
timestamp 1677579658
transform 1 0 13728 0 -1 23436
box -48 -56 144 834
use sg13g2_fill_2  FILLER_29_149
timestamp 1677580104
transform 1 0 15456 0 -1 23436
box -48 -56 240 834
use sg13g2_fill_1  FILLER_29_178
timestamp 1677579658
transform 1 0 18240 0 -1 23436
box -48 -56 144 834
use sg13g2_decap_4  FILLER_29_196
timestamp 1679577901
transform 1 0 19968 0 -1 23436
box -48 -56 432 834
use sg13g2_fill_1  FILLER_30_17
timestamp 1677579658
transform 1 0 2784 0 1 23436
box -48 -56 144 834
use sg13g2_decap_8  FILLER_30_75
timestamp 1679581782
transform 1 0 8352 0 1 23436
box -48 -56 720 834
use sg13g2_fill_2  FILLER_30_82
timestamp 1677580104
transform 1 0 9024 0 1 23436
box -48 -56 240 834
use sg13g2_fill_1  FILLER_30_84
timestamp 1677579658
transform 1 0 9216 0 1 23436
box -48 -56 144 834
use sg13g2_decap_4  FILLER_30_102
timestamp 1679577901
transform 1 0 10944 0 1 23436
box -48 -56 432 834
use sg13g2_decap_4  FILLER_30_173
timestamp 1679577901
transform 1 0 17760 0 1 23436
box -48 -56 432 834
use sg13g2_fill_1  FILLER_30_177
timestamp 1677579658
transform 1 0 18144 0 1 23436
box -48 -56 144 834
use sg13g2_fill_1  FILLER_30_199
timestamp 1677579658
transform 1 0 20256 0 1 23436
box -48 -56 144 834
use sg13g2_decap_8  FILLER_31_0
timestamp 1679581782
transform 1 0 1152 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_7
timestamp 1679581782
transform 1 0 1824 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_14
timestamp 1679581782
transform 1 0 2496 0 -1 24948
box -48 -56 720 834
use sg13g2_fill_1  FILLER_31_21
timestamp 1677579658
transform 1 0 3168 0 -1 24948
box -48 -56 144 834
use sg13g2_decap_8  FILLER_31_27
timestamp 1679581782
transform 1 0 3744 0 -1 24948
box -48 -56 720 834
use sg13g2_fill_2  FILLER_31_34
timestamp 1677580104
transform 1 0 4416 0 -1 24948
box -48 -56 240 834
use sg13g2_fill_1  FILLER_31_36
timestamp 1677579658
transform 1 0 4608 0 -1 24948
box -48 -56 144 834
use sg13g2_fill_1  FILLER_31_54
timestamp 1677579658
transform 1 0 6336 0 -1 24948
box -48 -56 144 834
use sg13g2_decap_4  FILLER_31_62
timestamp 1679577901
transform 1 0 7104 0 -1 24948
box -48 -56 432 834
use sg13g2_decap_4  FILLER_31_76
timestamp 1679577901
transform 1 0 8448 0 -1 24948
box -48 -56 432 834
use sg13g2_fill_2  FILLER_31_116
timestamp 1677580104
transform 1 0 12288 0 -1 24948
box -48 -56 240 834
use sg13g2_fill_1  FILLER_31_118
timestamp 1677579658
transform 1 0 12480 0 -1 24948
box -48 -56 144 834
use sg13g2_decap_4  FILLER_31_155
timestamp 1679577901
transform 1 0 16032 0 -1 24948
box -48 -56 432 834
use sg13g2_fill_1  FILLER_31_159
timestamp 1677579658
transform 1 0 16416 0 -1 24948
box -48 -56 144 834
use sg13g2_fill_2  FILLER_31_177
timestamp 1677580104
transform 1 0 18144 0 -1 24948
box -48 -56 240 834
use sg13g2_fill_1  FILLER_31_179
timestamp 1677579658
transform 1 0 18336 0 -1 24948
box -48 -56 144 834
use sg13g2_decap_8  FILLER_32_0
timestamp 1679581782
transform 1 0 1152 0 1 24948
box -48 -56 720 834
use sg13g2_fill_2  FILLER_32_7
timestamp 1677580104
transform 1 0 1824 0 1 24948
box -48 -56 240 834
use sg13g2_fill_1  FILLER_32_9
timestamp 1677579658
transform 1 0 2016 0 1 24948
box -48 -56 144 834
use sg13g2_fill_2  FILLER_32_31
timestamp 1677580104
transform 1 0 4128 0 1 24948
box -48 -56 240 834
use sg13g2_fill_1  FILLER_32_89
timestamp 1677579658
transform 1 0 9696 0 1 24948
box -48 -56 144 834
use sg13g2_decap_4  FILLER_32_102
timestamp 1679577901
transform 1 0 10944 0 1 24948
box -48 -56 432 834
use sg13g2_fill_1  FILLER_32_106
timestamp 1677579658
transform 1 0 11328 0 1 24948
box -48 -56 144 834
use sg13g2_decap_8  FILLER_32_117
timestamp 1679581782
transform 1 0 12384 0 1 24948
box -48 -56 720 834
use sg13g2_decap_4  FILLER_32_124
timestamp 1679577901
transform 1 0 13056 0 1 24948
box -48 -56 432 834
use sg13g2_decap_8  FILLER_32_151
timestamp 1679581782
transform 1 0 15648 0 1 24948
box -48 -56 720 834
use sg13g2_decap_4  FILLER_32_158
timestamp 1679577901
transform 1 0 16320 0 1 24948
box -48 -56 432 834
use sg13g2_fill_2  FILLER_32_198
timestamp 1677580104
transform 1 0 20160 0 1 24948
box -48 -56 240 834
use sg13g2_fill_2  FILLER_33_0
timestamp 1677580104
transform 1 0 1152 0 -1 26460
box -48 -56 240 834
use sg13g2_fill_1  FILLER_33_2
timestamp 1677579658
transform 1 0 1344 0 -1 26460
box -48 -56 144 834
use sg13g2_decap_8  FILLER_33_56
timestamp 1679581782
transform 1 0 6528 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_63
timestamp 1679581782
transform 1 0 7200 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_70
timestamp 1679581782
transform 1 0 7872 0 -1 26460
box -48 -56 720 834
use sg13g2_fill_2  FILLER_33_77
timestamp 1677580104
transform 1 0 8544 0 -1 26460
box -48 -56 240 834
use sg13g2_fill_1  FILLER_33_117
timestamp 1677579658
transform 1 0 12384 0 -1 26460
box -48 -56 144 834
use sg13g2_decap_8  FILLER_34_17
timestamp 1679581782
transform 1 0 2784 0 1 26460
box -48 -56 720 834
use sg13g2_fill_1  FILLER_34_24
timestamp 1677579658
transform 1 0 3456 0 1 26460
box -48 -56 144 834
use sg13g2_fill_2  FILLER_34_59
timestamp 1677580104
transform 1 0 6816 0 1 26460
box -48 -56 240 834
use sg13g2_fill_2  FILLER_34_78
timestamp 1677580104
transform 1 0 8640 0 1 26460
box -48 -56 240 834
use sg13g2_fill_1  FILLER_34_80
timestamp 1677579658
transform 1 0 8832 0 1 26460
box -48 -56 144 834
use sg13g2_fill_2  FILLER_34_113
timestamp 1677580104
transform 1 0 12000 0 1 26460
box -48 -56 240 834
use sg13g2_fill_1  FILLER_34_115
timestamp 1677579658
transform 1 0 12192 0 1 26460
box -48 -56 144 834
use sg13g2_fill_1  FILLER_34_133
timestamp 1677579658
transform 1 0 13920 0 1 26460
box -48 -56 144 834
use sg13g2_decap_8  FILLER_34_163
timestamp 1679581782
transform 1 0 16800 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_170
timestamp 1679581782
transform 1 0 17472 0 1 26460
box -48 -56 720 834
use sg13g2_fill_2  FILLER_34_177
timestamp 1677580104
transform 1 0 18144 0 1 26460
box -48 -56 240 834
use sg13g2_fill_1  FILLER_34_188
timestamp 1677579658
transform 1 0 19200 0 1 26460
box -48 -56 144 834
use sg13g2_fill_2  FILLER_34_197
timestamp 1677580104
transform 1 0 20064 0 1 26460
box -48 -56 240 834
use sg13g2_fill_1  FILLER_34_199
timestamp 1677579658
transform 1 0 20256 0 1 26460
box -48 -56 144 834
use sg13g2_decap_4  FILLER_35_0
timestamp 1679577901
transform 1 0 1152 0 -1 27972
box -48 -56 432 834
use sg13g2_fill_1  FILLER_35_4
timestamp 1677579658
transform 1 0 1536 0 -1 27972
box -48 -56 144 834
use sg13g2_decap_4  FILLER_35_39
timestamp 1679577901
transform 1 0 4896 0 -1 27972
box -48 -56 432 834
use sg13g2_decap_4  FILLER_35_53
timestamp 1679577901
transform 1 0 6240 0 -1 27972
box -48 -56 432 834
use sg13g2_fill_2  FILLER_35_74
timestamp 1677580104
transform 1 0 8256 0 -1 27972
box -48 -56 240 834
use sg13g2_fill_1  FILLER_35_84
timestamp 1677579658
transform 1 0 9216 0 -1 27972
box -48 -56 144 834
use sg13g2_decap_4  FILLER_35_90
timestamp 1679577901
transform 1 0 9792 0 -1 27972
box -48 -56 432 834
use sg13g2_fill_2  FILLER_35_94
timestamp 1677580104
transform 1 0 10176 0 -1 27972
box -48 -56 240 834
use sg13g2_decap_8  FILLER_35_118
timestamp 1679581782
transform 1 0 12480 0 -1 27972
box -48 -56 720 834
use sg13g2_fill_2  FILLER_35_125
timestamp 1677580104
transform 1 0 13152 0 -1 27972
box -48 -56 240 834
use sg13g2_fill_1  FILLER_35_127
timestamp 1677579658
transform 1 0 13344 0 -1 27972
box -48 -56 144 834
use sg13g2_fill_1  FILLER_35_150
timestamp 1677579658
transform 1 0 15552 0 -1 27972
box -48 -56 144 834
use sg13g2_fill_2  FILLER_35_168
timestamp 1677580104
transform 1 0 17280 0 -1 27972
box -48 -56 240 834
use sg13g2_decap_4  FILLER_35_196
timestamp 1679577901
transform 1 0 19968 0 -1 27972
box -48 -56 432 834
use sg13g2_fill_1  FILLER_36_0
timestamp 1677579658
transform 1 0 1152 0 1 27972
box -48 -56 144 834
use sg13g2_decap_4  FILLER_36_43
timestamp 1679577901
transform 1 0 5280 0 1 27972
box -48 -56 432 834
use sg13g2_decap_8  FILLER_36_126
timestamp 1679581782
transform 1 0 13248 0 1 27972
box -48 -56 720 834
use sg13g2_decap_4  FILLER_36_133
timestamp 1679577901
transform 1 0 13920 0 1 27972
box -48 -56 432 834
use sg13g2_fill_1  FILLER_36_157
timestamp 1677579658
transform 1 0 16224 0 1 27972
box -48 -56 144 834
use sg13g2_fill_1  FILLER_36_179
timestamp 1677579658
transform 1 0 18336 0 1 27972
box -48 -56 144 834
use sg13g2_fill_2  FILLER_36_197
timestamp 1677580104
transform 1 0 20064 0 1 27972
box -48 -56 240 834
use sg13g2_fill_1  FILLER_36_199
timestamp 1677579658
transform 1 0 20256 0 1 27972
box -48 -56 144 834
use sg13g2_decap_8  FILLER_37_0
timestamp 1679581782
transform 1 0 1152 0 -1 29484
box -48 -56 720 834
use sg13g2_fill_2  FILLER_37_7
timestamp 1677580104
transform 1 0 1824 0 -1 29484
box -48 -56 240 834
use sg13g2_fill_2  FILLER_37_26
timestamp 1677580104
transform 1 0 3648 0 -1 29484
box -48 -56 240 834
use sg13g2_decap_8  FILLER_37_57
timestamp 1679581782
transform 1 0 6624 0 -1 29484
box -48 -56 720 834
use sg13g2_fill_2  FILLER_37_84
timestamp 1677580104
transform 1 0 9216 0 -1 29484
box -48 -56 240 834
use sg13g2_fill_1  FILLER_37_103
timestamp 1677579658
transform 1 0 11040 0 -1 29484
box -48 -56 144 834
use sg13g2_fill_1  FILLER_37_114
timestamp 1677579658
transform 1 0 12096 0 -1 29484
box -48 -56 144 834
use sg13g2_decap_8  FILLER_37_153
timestamp 1679581782
transform 1 0 15840 0 -1 29484
box -48 -56 720 834
use sg13g2_fill_1  FILLER_38_0
timestamp 1677579658
transform 1 0 1152 0 1 29484
box -48 -56 144 834
use sg13g2_decap_4  FILLER_38_18
timestamp 1679577901
transform 1 0 2880 0 1 29484
box -48 -56 432 834
use sg13g2_fill_2  FILLER_38_22
timestamp 1677580104
transform 1 0 3264 0 1 29484
box -48 -56 240 834
use sg13g2_fill_2  FILLER_38_41
timestamp 1677580104
transform 1 0 5088 0 1 29484
box -48 -56 240 834
use sg13g2_fill_1  FILLER_38_43
timestamp 1677579658
transform 1 0 5280 0 1 29484
box -48 -56 144 834
use sg13g2_fill_2  FILLER_38_54
timestamp 1677580104
transform 1 0 6336 0 1 29484
box -48 -56 240 834
use sg13g2_fill_1  FILLER_38_56
timestamp 1677579658
transform 1 0 6528 0 1 29484
box -48 -56 144 834
use sg13g2_fill_1  FILLER_38_77
timestamp 1677579658
transform 1 0 8544 0 1 29484
box -48 -56 144 834
use sg13g2_decap_4  FILLER_38_88
timestamp 1679577901
transform 1 0 9600 0 1 29484
box -48 -56 432 834
use sg13g2_fill_1  FILLER_38_168
timestamp 1677579658
transform 1 0 17280 0 1 29484
box -48 -56 144 834
use sg13g2_fill_1  FILLER_38_199
timestamp 1677579658
transform 1 0 20256 0 1 29484
box -48 -56 144 834
use sg13g2_decap_8  FILLER_39_0
timestamp 1679581782
transform 1 0 1152 0 -1 30996
box -48 -56 720 834
use sg13g2_fill_2  FILLER_39_7
timestamp 1677580104
transform 1 0 1824 0 -1 30996
box -48 -56 240 834
use sg13g2_fill_1  FILLER_39_9
timestamp 1677579658
transform 1 0 2016 0 -1 30996
box -48 -56 144 834
use sg13g2_decap_4  FILLER_39_31
timestamp 1679577901
transform 1 0 4128 0 -1 30996
box -48 -56 432 834
use sg13g2_fill_1  FILLER_39_35
timestamp 1677579658
transform 1 0 4512 0 -1 30996
box -48 -56 144 834
use sg13g2_decap_8  FILLER_39_57
timestamp 1679581782
transform 1 0 6624 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_64
timestamp 1679581782
transform 1 0 7296 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_4  FILLER_39_71
timestamp 1679577901
transform 1 0 7968 0 -1 30996
box -48 -56 432 834
use sg13g2_fill_1  FILLER_39_75
timestamp 1677579658
transform 1 0 8352 0 -1 30996
box -48 -56 144 834
use sg13g2_fill_2  FILLER_39_98
timestamp 1677580104
transform 1 0 10560 0 -1 30996
box -48 -56 240 834
use sg13g2_decap_8  FILLER_39_120
timestamp 1679581782
transform 1 0 12672 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_4  FILLER_39_127
timestamp 1679577901
transform 1 0 13344 0 -1 30996
box -48 -56 432 834
use sg13g2_fill_2  FILLER_39_131
timestamp 1677580104
transform 1 0 13728 0 -1 30996
box -48 -56 240 834
use sg13g2_fill_2  FILLER_39_155
timestamp 1677580104
transform 1 0 16032 0 -1 30996
box -48 -56 240 834
use sg13g2_decap_8  FILLER_40_0
timestamp 1679581782
transform 1 0 1152 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_7
timestamp 1679581782
transform 1 0 1824 0 1 30996
box -48 -56 720 834
use sg13g2_fill_1  FILLER_40_14
timestamp 1677579658
transform 1 0 2496 0 1 30996
box -48 -56 144 834
use sg13g2_fill_2  FILLER_40_70
timestamp 1677580104
transform 1 0 7872 0 1 30996
box -48 -56 240 834
use sg13g2_fill_1  FILLER_40_72
timestamp 1677579658
transform 1 0 8064 0 1 30996
box -48 -56 144 834
use sg13g2_fill_1  FILLER_40_94
timestamp 1677579658
transform 1 0 10176 0 1 30996
box -48 -56 144 834
use sg13g2_decap_4  FILLER_40_116
timestamp 1679577901
transform 1 0 12288 0 1 30996
box -48 -56 432 834
use sg13g2_decap_8  FILLER_40_150
timestamp 1679581782
transform 1 0 15552 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_157
timestamp 1679581782
transform 1 0 16224 0 1 30996
box -48 -56 720 834
use sg13g2_fill_2  FILLER_40_164
timestamp 1677580104
transform 1 0 16896 0 1 30996
box -48 -56 240 834
use sg13g2_decap_8  FILLER_41_0
timestamp 1679581782
transform 1 0 1152 0 -1 32508
box -48 -56 720 834
use sg13g2_fill_2  FILLER_41_7
timestamp 1677580104
transform 1 0 1824 0 -1 32508
box -48 -56 240 834
use sg13g2_decap_4  FILLER_41_26
timestamp 1679577901
transform 1 0 3648 0 -1 32508
box -48 -56 432 834
use sg13g2_fill_1  FILLER_41_30
timestamp 1677579658
transform 1 0 4032 0 -1 32508
box -48 -56 144 834
use sg13g2_fill_2  FILLER_41_75
timestamp 1677580104
transform 1 0 8352 0 -1 32508
box -48 -56 240 834
use sg13g2_fill_1  FILLER_41_77
timestamp 1677579658
transform 1 0 8544 0 -1 32508
box -48 -56 144 834
use sg13g2_decap_8  FILLER_41_95
timestamp 1679581782
transform 1 0 10272 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_102
timestamp 1679581782
transform 1 0 10944 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_109
timestamp 1679581782
transform 1 0 11616 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_4  FILLER_41_116
timestamp 1679577901
transform 1 0 12288 0 -1 32508
box -48 -56 432 834
use sg13g2_fill_2  FILLER_41_120
timestamp 1677580104
transform 1 0 12672 0 -1 32508
box -48 -56 240 834
use sg13g2_decap_8  FILLER_41_142
timestamp 1679581782
transform 1 0 14784 0 -1 32508
box -48 -56 720 834
use sg13g2_fill_2  FILLER_41_149
timestamp 1677580104
transform 1 0 15456 0 -1 32508
box -48 -56 240 834
use sg13g2_fill_1  FILLER_41_151
timestamp 1677579658
transform 1 0 15648 0 -1 32508
box -48 -56 144 834
use sg13g2_fill_2  FILLER_41_173
timestamp 1677580104
transform 1 0 17760 0 -1 32508
box -48 -56 240 834
use sg13g2_decap_8  FILLER_42_0
timestamp 1679581782
transform 1 0 1152 0 1 32508
box -48 -56 720 834
use sg13g2_fill_1  FILLER_42_7
timestamp 1677579658
transform 1 0 1824 0 1 32508
box -48 -56 144 834
use sg13g2_decap_4  FILLER_42_29
timestamp 1679577901
transform 1 0 3936 0 1 32508
box -48 -56 432 834
use sg13g2_fill_1  FILLER_42_50
timestamp 1677579658
transform 1 0 5952 0 1 32508
box -48 -56 144 834
use sg13g2_fill_1  FILLER_42_59
timestamp 1677579658
transform 1 0 6816 0 1 32508
box -48 -56 144 834
use sg13g2_fill_1  FILLER_42_77
timestamp 1677579658
transform 1 0 8544 0 1 32508
box -48 -56 144 834
use sg13g2_decap_8  FILLER_42_95
timestamp 1679581782
transform 1 0 10272 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_102
timestamp 1679581782
transform 1 0 10944 0 1 32508
box -48 -56 720 834
use sg13g2_fill_2  FILLER_42_109
timestamp 1677580104
transform 1 0 11616 0 1 32508
box -48 -56 240 834
use sg13g2_decap_4  FILLER_42_128
timestamp 1679577901
transform 1 0 13440 0 1 32508
box -48 -56 432 834
use sg13g2_fill_2  FILLER_42_132
timestamp 1677580104
transform 1 0 13824 0 1 32508
box -48 -56 240 834
use sg13g2_fill_1  FILLER_42_199
timestamp 1677579658
transform 1 0 20256 0 1 32508
box -48 -56 144 834
use sg13g2_decap_8  FILLER_43_17
timestamp 1679581782
transform 1 0 2784 0 -1 34020
box -48 -56 720 834
use sg13g2_fill_2  FILLER_43_24
timestamp 1677580104
transform 1 0 3456 0 -1 34020
box -48 -56 240 834
use sg13g2_fill_1  FILLER_43_26
timestamp 1677579658
transform 1 0 3648 0 -1 34020
box -48 -56 144 834
use sg13g2_fill_2  FILLER_43_146
timestamp 1677580104
transform 1 0 15168 0 -1 34020
box -48 -56 240 834
use sg13g2_fill_2  FILLER_43_175
timestamp 1677580104
transform 1 0 17952 0 -1 34020
box -48 -56 240 834
use sg13g2_fill_1  FILLER_43_177
timestamp 1677579658
transform 1 0 18144 0 -1 34020
box -48 -56 144 834
use sg13g2_fill_1  FILLER_43_199
timestamp 1677579658
transform 1 0 20256 0 -1 34020
box -48 -56 144 834
use sg13g2_fill_2  FILLER_44_0
timestamp 1677580104
transform 1 0 1152 0 1 34020
box -48 -56 240 834
use sg13g2_fill_1  FILLER_44_2
timestamp 1677579658
transform 1 0 1344 0 1 34020
box -48 -56 144 834
use sg13g2_fill_1  FILLER_44_49
timestamp 1677579658
transform 1 0 5856 0 1 34020
box -48 -56 144 834
use sg13g2_fill_2  FILLER_44_72
timestamp 1677580104
transform 1 0 8064 0 1 34020
box -48 -56 240 834
use sg13g2_fill_1  FILLER_44_74
timestamp 1677579658
transform 1 0 8256 0 1 34020
box -48 -56 144 834
use sg13g2_fill_1  FILLER_44_78
timestamp 1677579658
transform 1 0 8640 0 1 34020
box -48 -56 144 834
use sg13g2_fill_2  FILLER_44_147
timestamp 1677580104
transform 1 0 15264 0 1 34020
box -48 -56 240 834
use sg13g2_fill_2  FILLER_44_166
timestamp 1677580104
transform 1 0 17088 0 1 34020
box -48 -56 240 834
use sg13g2_fill_1  FILLER_44_168
timestamp 1677579658
transform 1 0 17280 0 1 34020
box -48 -56 144 834
use sg13g2_fill_1  FILLER_44_199
timestamp 1677579658
transform 1 0 20256 0 1 34020
box -48 -56 144 834
use sg13g2_fill_2  FILLER_45_0
timestamp 1677580104
transform 1 0 1152 0 -1 35532
box -48 -56 240 834
use sg13g2_fill_1  FILLER_45_2
timestamp 1677579658
transform 1 0 1344 0 -1 35532
box -48 -56 144 834
use sg13g2_fill_2  FILLER_45_24
timestamp 1677580104
transform 1 0 3456 0 -1 35532
box -48 -56 240 834
use sg13g2_fill_1  FILLER_45_26
timestamp 1677579658
transform 1 0 3648 0 -1 35532
box -48 -56 144 834
use sg13g2_fill_2  FILLER_45_31
timestamp 1677580104
transform 1 0 4128 0 -1 35532
box -48 -56 240 834
use sg13g2_fill_2  FILLER_45_67
timestamp 1677580104
transform 1 0 7584 0 -1 35532
box -48 -56 240 834
use sg13g2_fill_1  FILLER_45_69
timestamp 1677579658
transform 1 0 7776 0 -1 35532
box -48 -56 144 834
use sg13g2_fill_2  FILLER_45_109
timestamp 1677580104
transform 1 0 11616 0 -1 35532
box -48 -56 240 834
use sg13g2_fill_2  FILLER_45_128
timestamp 1677580104
transform 1 0 13440 0 -1 35532
box -48 -56 240 834
use sg13g2_fill_2  FILLER_45_168
timestamp 1677580104
transform 1 0 17280 0 -1 35532
box -48 -56 240 834
use sg13g2_fill_1  FILLER_45_170
timestamp 1677579658
transform 1 0 17472 0 -1 35532
box -48 -56 144 834
use sg13g2_fill_2  FILLER_46_0
timestamp 1677580104
transform 1 0 1152 0 1 35532
box -48 -56 240 834
use sg13g2_fill_2  FILLER_46_27
timestamp 1677580104
transform 1 0 3744 0 1 35532
box -48 -56 240 834
use sg13g2_fill_2  FILLER_46_78
timestamp 1677580104
transform 1 0 8640 0 1 35532
box -48 -56 240 834
use sg13g2_fill_1  FILLER_46_80
timestamp 1677579658
transform 1 0 8832 0 1 35532
box -48 -56 144 834
use sg13g2_decap_8  FILLER_46_125
timestamp 1679581782
transform 1 0 13152 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_132
timestamp 1679581782
transform 1 0 13824 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_139
timestamp 1679581782
transform 1 0 14496 0 1 35532
box -48 -56 720 834
use sg13g2_fill_1  FILLER_46_199
timestamp 1677579658
transform 1 0 20256 0 1 35532
box -48 -56 144 834
use sg13g2_fill_2  FILLER_47_17
timestamp 1677580104
transform 1 0 2784 0 -1 37044
box -48 -56 240 834
use sg13g2_decap_4  FILLER_47_82
timestamp 1679577901
transform 1 0 9024 0 -1 37044
box -48 -56 432 834
use sg13g2_decap_8  FILLER_47_124
timestamp 1679581782
transform 1 0 13056 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_131
timestamp 1679581782
transform 1 0 13728 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_138
timestamp 1679581782
transform 1 0 14400 0 -1 37044
box -48 -56 720 834
use sg13g2_fill_2  FILLER_47_162
timestamp 1677580104
transform 1 0 16704 0 -1 37044
box -48 -56 240 834
use sg13g2_fill_2  FILLER_47_173
timestamp 1677580104
transform 1 0 17760 0 -1 37044
box -48 -56 240 834
use sg13g2_fill_1  FILLER_47_175
timestamp 1677579658
transform 1 0 17952 0 -1 37044
box -48 -56 144 834
use sg13g2_fill_2  FILLER_48_0
timestamp 1677580104
transform 1 0 1152 0 1 37044
box -48 -56 240 834
use sg13g2_fill_2  FILLER_48_31
timestamp 1677580104
transform 1 0 4128 0 1 37044
box -48 -56 240 834
use sg13g2_decap_8  FILLER_48_95
timestamp 1679581782
transform 1 0 10272 0 1 37044
box -48 -56 720 834
use sg13g2_decap_4  FILLER_48_102
timestamp 1679577901
transform 1 0 10944 0 1 37044
box -48 -56 432 834
use sg13g2_fill_1  FILLER_48_106
timestamp 1677579658
transform 1 0 11328 0 1 37044
box -48 -56 144 834
use sg13g2_decap_8  FILLER_48_124
timestamp 1679581782
transform 1 0 13056 0 1 37044
box -48 -56 720 834
use sg13g2_fill_2  FILLER_48_131
timestamp 1677580104
transform 1 0 13728 0 1 37044
box -48 -56 240 834
use sg13g2_fill_2  FILLER_48_154
timestamp 1677580104
transform 1 0 15936 0 1 37044
box -48 -56 240 834
use sg13g2_fill_2  FILLER_48_173
timestamp 1677580104
transform 1 0 17760 0 1 37044
box -48 -56 240 834
use sg13g2_fill_1  FILLER_48_175
timestamp 1677579658
transform 1 0 17952 0 1 37044
box -48 -56 144 834
use sg13g2_fill_1  FILLER_49_17
timestamp 1677579658
transform 1 0 2784 0 -1 38556
box -48 -56 144 834
use sg13g2_fill_1  FILLER_49_26
timestamp 1677579658
transform 1 0 3648 0 -1 38556
box -48 -56 144 834
use sg13g2_fill_2  FILLER_49_48
timestamp 1677580104
transform 1 0 5760 0 -1 38556
box -48 -56 240 834
use sg13g2_fill_1  FILLER_49_53
timestamp 1677579658
transform 1 0 6240 0 -1 38556
box -48 -56 144 834
use sg13g2_decap_4  FILLER_49_94
timestamp 1679577901
transform 1 0 10176 0 -1 38556
box -48 -56 432 834
use sg13g2_decap_4  FILLER_49_115
timestamp 1679577901
transform 1 0 12192 0 -1 38556
box -48 -56 432 834
use sg13g2_fill_2  FILLER_49_119
timestamp 1677580104
transform 1 0 12576 0 -1 38556
box -48 -56 240 834
use sg13g2_fill_1  FILLER_50_0
timestamp 1677579658
transform 1 0 1152 0 1 38556
box -48 -56 144 834
use sg13g2_fill_1  FILLER_50_120
timestamp 1677579658
transform 1 0 12672 0 1 38556
box -48 -56 144 834
use sg13g2_decap_8  FILLER_50_125
timestamp 1679581782
transform 1 0 13152 0 1 38556
box -48 -56 720 834
use sg13g2_fill_1  FILLER_50_132
timestamp 1677579658
transform 1 0 13824 0 1 38556
box -48 -56 144 834
use sg13g2_fill_1  FILLER_50_179
timestamp 1677579658
transform 1 0 18336 0 1 38556
box -48 -56 144 834
use sg13g2_fill_1  FILLER_51_28
timestamp 1677579658
transform 1 0 3840 0 -1 40068
box -48 -56 144 834
use sg13g2_fill_1  FILLER_51_93
timestamp 1677579658
transform 1 0 10080 0 -1 40068
box -48 -56 144 834
use sg13g2_fill_1  FILLER_51_124
timestamp 1677579658
transform 1 0 13056 0 -1 40068
box -48 -56 144 834
use sg13g2_fill_1  FILLER_51_163
timestamp 1677579658
transform 1 0 16800 0 -1 40068
box -48 -56 144 834
use sg13g2_fill_1  FILLER_51_176
timestamp 1677579658
transform 1 0 18048 0 -1 40068
box -48 -56 144 834
use sg13g2_fill_2  FILLER_51_188
timestamp 1677580104
transform 1 0 19200 0 -1 40068
box -48 -56 240 834
use sg13g2_fill_2  FILLER_51_194
timestamp 1677580104
transform 1 0 19776 0 -1 40068
box -48 -56 240 834
use sg13g2_decap_4  FILLER_52_13
timestamp 1679577901
transform 1 0 2400 0 1 40068
box -48 -56 432 834
use sg13g2_fill_1  FILLER_52_117
timestamp 1677579658
transform 1 0 12384 0 1 40068
box -48 -56 144 834
use sg13g2_fill_1  FILLER_52_168
timestamp 1677579658
transform 1 0 17280 0 1 40068
box -48 -56 144 834
use sg13g2_fill_1  FILLER_52_188
timestamp 1677579658
transform 1 0 19200 0 1 40068
box -48 -56 144 834
use sg13g2_fill_1  FILLER_52_193
timestamp 1677579658
transform 1 0 19680 0 1 40068
box -48 -56 144 834
use sg13g2_fill_2  FILLER_52_198
timestamp 1677580104
transform 1 0 20160 0 1 40068
box -48 -56 240 834
use sg13g2_fill_1  FILLER_53_3
timestamp 1677579658
transform 1 0 1440 0 -1 41580
box -48 -56 144 834
use sg13g2_decap_8  FILLER_53_99
timestamp 1679581782
transform 1 0 10656 0 -1 41580
box -48 -56 720 834
use sg13g2_fill_2  FILLER_53_106
timestamp 1677580104
transform 1 0 11328 0 -1 41580
box -48 -56 240 834
use sg13g2_fill_2  FILLER_53_129
timestamp 1677580104
transform 1 0 13536 0 -1 41580
box -48 -56 240 834
use sg13g2_fill_2  FILLER_53_135
timestamp 1677580104
transform 1 0 14112 0 -1 41580
box -48 -56 240 834
use sg13g2_fill_2  FILLER_53_149
timestamp 1677580104
transform 1 0 15456 0 -1 41580
box -48 -56 240 834
use sg13g2_fill_1  FILLER_53_166
timestamp 1677579658
transform 1 0 17088 0 -1 41580
box -48 -56 144 834
use sg13g2_fill_1  FILLER_53_175
timestamp 1677579658
transform 1 0 17952 0 -1 41580
box -48 -56 144 834
use sg13g2_fill_1  FILLER_53_188
timestamp 1677579658
transform 1 0 19200 0 -1 41580
box -48 -56 144 834
use sg13g2_fill_2  FILLER_53_197
timestamp 1677580104
transform 1 0 20064 0 -1 41580
box -48 -56 240 834
use sg13g2_fill_1  FILLER_53_199
timestamp 1677579658
transform 1 0 20256 0 -1 41580
box -48 -56 144 834
<< labels >>
flabel metal3 s 21424 23396 21504 23476 0 FreeSans 320 0 0 0 CLK_TT_PROJECT
port 0 nsew signal output
flabel metal3 s 0 16172 80 16252 0 FreeSans 320 0 0 0 E1END[0]
port 1 nsew signal input
flabel metal3 s 0 16508 80 16588 0 FreeSans 320 0 0 0 E1END[1]
port 2 nsew signal input
flabel metal3 s 0 16844 80 16924 0 FreeSans 320 0 0 0 E1END[2]
port 3 nsew signal input
flabel metal3 s 0 17180 80 17260 0 FreeSans 320 0 0 0 E1END[3]
port 4 nsew signal input
flabel metal3 s 0 20204 80 20284 0 FreeSans 320 0 0 0 E2END[0]
port 5 nsew signal input
flabel metal3 s 0 20540 80 20620 0 FreeSans 320 0 0 0 E2END[1]
port 6 nsew signal input
flabel metal3 s 0 20876 80 20956 0 FreeSans 320 0 0 0 E2END[2]
port 7 nsew signal input
flabel metal3 s 0 21212 80 21292 0 FreeSans 320 0 0 0 E2END[3]
port 8 nsew signal input
flabel metal3 s 0 21548 80 21628 0 FreeSans 320 0 0 0 E2END[4]
port 9 nsew signal input
flabel metal3 s 0 21884 80 21964 0 FreeSans 320 0 0 0 E2END[5]
port 10 nsew signal input
flabel metal3 s 0 22220 80 22300 0 FreeSans 320 0 0 0 E2END[6]
port 11 nsew signal input
flabel metal3 s 0 22556 80 22636 0 FreeSans 320 0 0 0 E2END[7]
port 12 nsew signal input
flabel metal3 s 0 17516 80 17596 0 FreeSans 320 0 0 0 E2MID[0]
port 13 nsew signal input
flabel metal3 s 0 17852 80 17932 0 FreeSans 320 0 0 0 E2MID[1]
port 14 nsew signal input
flabel metal3 s 0 18188 80 18268 0 FreeSans 320 0 0 0 E2MID[2]
port 15 nsew signal input
flabel metal3 s 0 18524 80 18604 0 FreeSans 320 0 0 0 E2MID[3]
port 16 nsew signal input
flabel metal3 s 0 18860 80 18940 0 FreeSans 320 0 0 0 E2MID[4]
port 17 nsew signal input
flabel metal3 s 0 19196 80 19276 0 FreeSans 320 0 0 0 E2MID[5]
port 18 nsew signal input
flabel metal3 s 0 19532 80 19612 0 FreeSans 320 0 0 0 E2MID[6]
port 19 nsew signal input
flabel metal3 s 0 19868 80 19948 0 FreeSans 320 0 0 0 E2MID[7]
port 20 nsew signal input
flabel metal3 s 0 28268 80 28348 0 FreeSans 320 0 0 0 E6END[0]
port 21 nsew signal input
flabel metal3 s 0 31628 80 31708 0 FreeSans 320 0 0 0 E6END[10]
port 22 nsew signal input
flabel metal3 s 0 31964 80 32044 0 FreeSans 320 0 0 0 E6END[11]
port 23 nsew signal input
flabel metal3 s 0 28604 80 28684 0 FreeSans 320 0 0 0 E6END[1]
port 24 nsew signal input
flabel metal3 s 0 28940 80 29020 0 FreeSans 320 0 0 0 E6END[2]
port 25 nsew signal input
flabel metal3 s 0 29276 80 29356 0 FreeSans 320 0 0 0 E6END[3]
port 26 nsew signal input
flabel metal3 s 0 29612 80 29692 0 FreeSans 320 0 0 0 E6END[4]
port 27 nsew signal input
flabel metal3 s 0 29948 80 30028 0 FreeSans 320 0 0 0 E6END[5]
port 28 nsew signal input
flabel metal3 s 0 30284 80 30364 0 FreeSans 320 0 0 0 E6END[6]
port 29 nsew signal input
flabel metal3 s 0 30620 80 30700 0 FreeSans 320 0 0 0 E6END[7]
port 30 nsew signal input
flabel metal3 s 0 30956 80 31036 0 FreeSans 320 0 0 0 E6END[8]
port 31 nsew signal input
flabel metal3 s 0 31292 80 31372 0 FreeSans 320 0 0 0 E6END[9]
port 32 nsew signal input
flabel metal3 s 0 22892 80 22972 0 FreeSans 320 0 0 0 EE4END[0]
port 33 nsew signal input
flabel metal3 s 0 26252 80 26332 0 FreeSans 320 0 0 0 EE4END[10]
port 34 nsew signal input
flabel metal3 s 0 26588 80 26668 0 FreeSans 320 0 0 0 EE4END[11]
port 35 nsew signal input
flabel metal3 s 0 26924 80 27004 0 FreeSans 320 0 0 0 EE4END[12]
port 36 nsew signal input
flabel metal3 s 0 27260 80 27340 0 FreeSans 320 0 0 0 EE4END[13]
port 37 nsew signal input
flabel metal3 s 0 27596 80 27676 0 FreeSans 320 0 0 0 EE4END[14]
port 38 nsew signal input
flabel metal3 s 0 27932 80 28012 0 FreeSans 320 0 0 0 EE4END[15]
port 39 nsew signal input
flabel metal3 s 0 23228 80 23308 0 FreeSans 320 0 0 0 EE4END[1]
port 40 nsew signal input
flabel metal3 s 0 23564 80 23644 0 FreeSans 320 0 0 0 EE4END[2]
port 41 nsew signal input
flabel metal3 s 0 23900 80 23980 0 FreeSans 320 0 0 0 EE4END[3]
port 42 nsew signal input
flabel metal3 s 0 24236 80 24316 0 FreeSans 320 0 0 0 EE4END[4]
port 43 nsew signal input
flabel metal3 s 0 24572 80 24652 0 FreeSans 320 0 0 0 EE4END[5]
port 44 nsew signal input
flabel metal3 s 0 24908 80 24988 0 FreeSans 320 0 0 0 EE4END[6]
port 45 nsew signal input
flabel metal3 s 0 25244 80 25324 0 FreeSans 320 0 0 0 EE4END[7]
port 46 nsew signal input
flabel metal3 s 0 25580 80 25660 0 FreeSans 320 0 0 0 EE4END[8]
port 47 nsew signal input
flabel metal3 s 0 25916 80 25996 0 FreeSans 320 0 0 0 EE4END[9]
port 48 nsew signal input
flabel metal3 s 21424 22892 21504 22972 0 FreeSans 320 0 0 0 ENA_TT_PROJECT
port 49 nsew signal output
flabel metal3 s 0 32300 80 32380 0 FreeSans 320 0 0 0 FrameData[0]
port 50 nsew signal input
flabel metal3 s 0 35660 80 35740 0 FreeSans 320 0 0 0 FrameData[10]
port 51 nsew signal input
flabel metal3 s 0 35996 80 36076 0 FreeSans 320 0 0 0 FrameData[11]
port 52 nsew signal input
flabel metal3 s 0 36332 80 36412 0 FreeSans 320 0 0 0 FrameData[12]
port 53 nsew signal input
flabel metal3 s 0 36668 80 36748 0 FreeSans 320 0 0 0 FrameData[13]
port 54 nsew signal input
flabel metal3 s 0 37004 80 37084 0 FreeSans 320 0 0 0 FrameData[14]
port 55 nsew signal input
flabel metal3 s 0 37340 80 37420 0 FreeSans 320 0 0 0 FrameData[15]
port 56 nsew signal input
flabel metal3 s 0 37676 80 37756 0 FreeSans 320 0 0 0 FrameData[16]
port 57 nsew signal input
flabel metal3 s 0 38012 80 38092 0 FreeSans 320 0 0 0 FrameData[17]
port 58 nsew signal input
flabel metal3 s 0 38348 80 38428 0 FreeSans 320 0 0 0 FrameData[18]
port 59 nsew signal input
flabel metal3 s 0 38684 80 38764 0 FreeSans 320 0 0 0 FrameData[19]
port 60 nsew signal input
flabel metal3 s 0 32636 80 32716 0 FreeSans 320 0 0 0 FrameData[1]
port 61 nsew signal input
flabel metal3 s 0 39020 80 39100 0 FreeSans 320 0 0 0 FrameData[20]
port 62 nsew signal input
flabel metal3 s 0 39356 80 39436 0 FreeSans 320 0 0 0 FrameData[21]
port 63 nsew signal input
flabel metal3 s 0 39692 80 39772 0 FreeSans 320 0 0 0 FrameData[22]
port 64 nsew signal input
flabel metal3 s 0 40028 80 40108 0 FreeSans 320 0 0 0 FrameData[23]
port 65 nsew signal input
flabel metal3 s 0 40364 80 40444 0 FreeSans 320 0 0 0 FrameData[24]
port 66 nsew signal input
flabel metal3 s 0 40700 80 40780 0 FreeSans 320 0 0 0 FrameData[25]
port 67 nsew signal input
flabel metal3 s 0 41036 80 41116 0 FreeSans 320 0 0 0 FrameData[26]
port 68 nsew signal input
flabel metal3 s 0 41372 80 41452 0 FreeSans 320 0 0 0 FrameData[27]
port 69 nsew signal input
flabel metal3 s 0 41708 80 41788 0 FreeSans 320 0 0 0 FrameData[28]
port 70 nsew signal input
flabel metal3 s 0 42044 80 42124 0 FreeSans 320 0 0 0 FrameData[29]
port 71 nsew signal input
flabel metal3 s 0 32972 80 33052 0 FreeSans 320 0 0 0 FrameData[2]
port 72 nsew signal input
flabel metal3 s 0 42380 80 42460 0 FreeSans 320 0 0 0 FrameData[30]
port 73 nsew signal input
flabel metal3 s 0 42716 80 42796 0 FreeSans 320 0 0 0 FrameData[31]
port 74 nsew signal input
flabel metal3 s 0 33308 80 33388 0 FreeSans 320 0 0 0 FrameData[3]
port 75 nsew signal input
flabel metal3 s 0 33644 80 33724 0 FreeSans 320 0 0 0 FrameData[4]
port 76 nsew signal input
flabel metal3 s 0 33980 80 34060 0 FreeSans 320 0 0 0 FrameData[5]
port 77 nsew signal input
flabel metal3 s 0 34316 80 34396 0 FreeSans 320 0 0 0 FrameData[6]
port 78 nsew signal input
flabel metal3 s 0 34652 80 34732 0 FreeSans 320 0 0 0 FrameData[7]
port 79 nsew signal input
flabel metal3 s 0 34988 80 35068 0 FreeSans 320 0 0 0 FrameData[8]
port 80 nsew signal input
flabel metal3 s 0 35324 80 35404 0 FreeSans 320 0 0 0 FrameData[9]
port 81 nsew signal input
flabel metal3 s 21424 24404 21504 24484 0 FreeSans 320 0 0 0 FrameData_O[0]
port 82 nsew signal output
flabel metal3 s 21424 29444 21504 29524 0 FreeSans 320 0 0 0 FrameData_O[10]
port 83 nsew signal output
flabel metal3 s 21424 29948 21504 30028 0 FreeSans 320 0 0 0 FrameData_O[11]
port 84 nsew signal output
flabel metal3 s 21424 30452 21504 30532 0 FreeSans 320 0 0 0 FrameData_O[12]
port 85 nsew signal output
flabel metal3 s 21424 30956 21504 31036 0 FreeSans 320 0 0 0 FrameData_O[13]
port 86 nsew signal output
flabel metal3 s 21424 31460 21504 31540 0 FreeSans 320 0 0 0 FrameData_O[14]
port 87 nsew signal output
flabel metal3 s 21424 31964 21504 32044 0 FreeSans 320 0 0 0 FrameData_O[15]
port 88 nsew signal output
flabel metal3 s 21424 32468 21504 32548 0 FreeSans 320 0 0 0 FrameData_O[16]
port 89 nsew signal output
flabel metal3 s 21424 32972 21504 33052 0 FreeSans 320 0 0 0 FrameData_O[17]
port 90 nsew signal output
flabel metal3 s 21424 33476 21504 33556 0 FreeSans 320 0 0 0 FrameData_O[18]
port 91 nsew signal output
flabel metal3 s 21424 33980 21504 34060 0 FreeSans 320 0 0 0 FrameData_O[19]
port 92 nsew signal output
flabel metal3 s 21424 24908 21504 24988 0 FreeSans 320 0 0 0 FrameData_O[1]
port 93 nsew signal output
flabel metal3 s 21424 34484 21504 34564 0 FreeSans 320 0 0 0 FrameData_O[20]
port 94 nsew signal output
flabel metal3 s 21424 34988 21504 35068 0 FreeSans 320 0 0 0 FrameData_O[21]
port 95 nsew signal output
flabel metal3 s 21424 35492 21504 35572 0 FreeSans 320 0 0 0 FrameData_O[22]
port 96 nsew signal output
flabel metal3 s 21424 35996 21504 36076 0 FreeSans 320 0 0 0 FrameData_O[23]
port 97 nsew signal output
flabel metal3 s 21424 36500 21504 36580 0 FreeSans 320 0 0 0 FrameData_O[24]
port 98 nsew signal output
flabel metal3 s 21424 37004 21504 37084 0 FreeSans 320 0 0 0 FrameData_O[25]
port 99 nsew signal output
flabel metal3 s 21424 37508 21504 37588 0 FreeSans 320 0 0 0 FrameData_O[26]
port 100 nsew signal output
flabel metal3 s 21424 38012 21504 38092 0 FreeSans 320 0 0 0 FrameData_O[27]
port 101 nsew signal output
flabel metal3 s 21424 38516 21504 38596 0 FreeSans 320 0 0 0 FrameData_O[28]
port 102 nsew signal output
flabel metal3 s 21424 39020 21504 39100 0 FreeSans 320 0 0 0 FrameData_O[29]
port 103 nsew signal output
flabel metal3 s 21424 25412 21504 25492 0 FreeSans 320 0 0 0 FrameData_O[2]
port 104 nsew signal output
flabel metal3 s 21424 39524 21504 39604 0 FreeSans 320 0 0 0 FrameData_O[30]
port 105 nsew signal output
flabel metal3 s 21424 40028 21504 40108 0 FreeSans 320 0 0 0 FrameData_O[31]
port 106 nsew signal output
flabel metal3 s 21424 25916 21504 25996 0 FreeSans 320 0 0 0 FrameData_O[3]
port 107 nsew signal output
flabel metal3 s 21424 26420 21504 26500 0 FreeSans 320 0 0 0 FrameData_O[4]
port 108 nsew signal output
flabel metal3 s 21424 26924 21504 27004 0 FreeSans 320 0 0 0 FrameData_O[5]
port 109 nsew signal output
flabel metal3 s 21424 27428 21504 27508 0 FreeSans 320 0 0 0 FrameData_O[6]
port 110 nsew signal output
flabel metal3 s 21424 27932 21504 28012 0 FreeSans 320 0 0 0 FrameData_O[7]
port 111 nsew signal output
flabel metal3 s 21424 28436 21504 28516 0 FreeSans 320 0 0 0 FrameData_O[8]
port 112 nsew signal output
flabel metal3 s 21424 28940 21504 29020 0 FreeSans 320 0 0 0 FrameData_O[9]
port 113 nsew signal output
flabel metal2 s 15800 0 15880 80 0 FreeSans 320 0 0 0 FrameStrobe[0]
port 114 nsew signal input
flabel metal2 s 17720 0 17800 80 0 FreeSans 320 0 0 0 FrameStrobe[10]
port 115 nsew signal input
flabel metal2 s 17912 0 17992 80 0 FreeSans 320 0 0 0 FrameStrobe[11]
port 116 nsew signal input
flabel metal2 s 18104 0 18184 80 0 FreeSans 320 0 0 0 FrameStrobe[12]
port 117 nsew signal input
flabel metal2 s 18296 0 18376 80 0 FreeSans 320 0 0 0 FrameStrobe[13]
port 118 nsew signal input
flabel metal2 s 18488 0 18568 80 0 FreeSans 320 0 0 0 FrameStrobe[14]
port 119 nsew signal input
flabel metal2 s 18680 0 18760 80 0 FreeSans 320 0 0 0 FrameStrobe[15]
port 120 nsew signal input
flabel metal2 s 18872 0 18952 80 0 FreeSans 320 0 0 0 FrameStrobe[16]
port 121 nsew signal input
flabel metal2 s 19064 0 19144 80 0 FreeSans 320 0 0 0 FrameStrobe[17]
port 122 nsew signal input
flabel metal2 s 19256 0 19336 80 0 FreeSans 320 0 0 0 FrameStrobe[18]
port 123 nsew signal input
flabel metal2 s 19448 0 19528 80 0 FreeSans 320 0 0 0 FrameStrobe[19]
port 124 nsew signal input
flabel metal2 s 15992 0 16072 80 0 FreeSans 320 0 0 0 FrameStrobe[1]
port 125 nsew signal input
flabel metal2 s 16184 0 16264 80 0 FreeSans 320 0 0 0 FrameStrobe[2]
port 126 nsew signal input
flabel metal2 s 16376 0 16456 80 0 FreeSans 320 0 0 0 FrameStrobe[3]
port 127 nsew signal input
flabel metal2 s 16568 0 16648 80 0 FreeSans 320 0 0 0 FrameStrobe[4]
port 128 nsew signal input
flabel metal2 s 16760 0 16840 80 0 FreeSans 320 0 0 0 FrameStrobe[5]
port 129 nsew signal input
flabel metal2 s 16952 0 17032 80 0 FreeSans 320 0 0 0 FrameStrobe[6]
port 130 nsew signal input
flabel metal2 s 17144 0 17224 80 0 FreeSans 320 0 0 0 FrameStrobe[7]
port 131 nsew signal input
flabel metal2 s 17336 0 17416 80 0 FreeSans 320 0 0 0 FrameStrobe[8]
port 132 nsew signal input
flabel metal2 s 17528 0 17608 80 0 FreeSans 320 0 0 0 FrameStrobe[9]
port 133 nsew signal input
flabel metal2 s 15800 42928 15880 43008 0 FreeSans 320 0 0 0 FrameStrobe_O[0]
port 134 nsew signal output
flabel metal2 s 17720 42928 17800 43008 0 FreeSans 320 0 0 0 FrameStrobe_O[10]
port 135 nsew signal output
flabel metal2 s 17912 42928 17992 43008 0 FreeSans 320 0 0 0 FrameStrobe_O[11]
port 136 nsew signal output
flabel metal2 s 18104 42928 18184 43008 0 FreeSans 320 0 0 0 FrameStrobe_O[12]
port 137 nsew signal output
flabel metal2 s 18296 42928 18376 43008 0 FreeSans 320 0 0 0 FrameStrobe_O[13]
port 138 nsew signal output
flabel metal2 s 18488 42928 18568 43008 0 FreeSans 320 0 0 0 FrameStrobe_O[14]
port 139 nsew signal output
flabel metal2 s 18680 42928 18760 43008 0 FreeSans 320 0 0 0 FrameStrobe_O[15]
port 140 nsew signal output
flabel metal2 s 18872 42928 18952 43008 0 FreeSans 320 0 0 0 FrameStrobe_O[16]
port 141 nsew signal output
flabel metal2 s 19064 42928 19144 43008 0 FreeSans 320 0 0 0 FrameStrobe_O[17]
port 142 nsew signal output
flabel metal2 s 19256 42928 19336 43008 0 FreeSans 320 0 0 0 FrameStrobe_O[18]
port 143 nsew signal output
flabel metal2 s 19448 42928 19528 43008 0 FreeSans 320 0 0 0 FrameStrobe_O[19]
port 144 nsew signal output
flabel metal2 s 15992 42928 16072 43008 0 FreeSans 320 0 0 0 FrameStrobe_O[1]
port 145 nsew signal output
flabel metal2 s 16184 42928 16264 43008 0 FreeSans 320 0 0 0 FrameStrobe_O[2]
port 146 nsew signal output
flabel metal2 s 16376 42928 16456 43008 0 FreeSans 320 0 0 0 FrameStrobe_O[3]
port 147 nsew signal output
flabel metal2 s 16568 42928 16648 43008 0 FreeSans 320 0 0 0 FrameStrobe_O[4]
port 148 nsew signal output
flabel metal2 s 16760 42928 16840 43008 0 FreeSans 320 0 0 0 FrameStrobe_O[5]
port 149 nsew signal output
flabel metal2 s 16952 42928 17032 43008 0 FreeSans 320 0 0 0 FrameStrobe_O[6]
port 150 nsew signal output
flabel metal2 s 17144 42928 17224 43008 0 FreeSans 320 0 0 0 FrameStrobe_O[7]
port 151 nsew signal output
flabel metal2 s 17336 42928 17416 43008 0 FreeSans 320 0 0 0 FrameStrobe_O[8]
port 152 nsew signal output
flabel metal2 s 17528 42928 17608 43008 0 FreeSans 320 0 0 0 FrameStrobe_O[9]
port 153 nsew signal output
flabel metal2 s 1784 42928 1864 43008 0 FreeSans 320 0 0 0 N1BEG[0]
port 154 nsew signal output
flabel metal2 s 1976 42928 2056 43008 0 FreeSans 320 0 0 0 N1BEG[1]
port 155 nsew signal output
flabel metal2 s 2168 42928 2248 43008 0 FreeSans 320 0 0 0 N1BEG[2]
port 156 nsew signal output
flabel metal2 s 2360 42928 2440 43008 0 FreeSans 320 0 0 0 N1BEG[3]
port 157 nsew signal output
flabel metal2 s 1784 0 1864 80 0 FreeSans 320 0 0 0 N1END[0]
port 158 nsew signal input
flabel metal2 s 1976 0 2056 80 0 FreeSans 320 0 0 0 N1END[1]
port 159 nsew signal input
flabel metal2 s 2168 0 2248 80 0 FreeSans 320 0 0 0 N1END[2]
port 160 nsew signal input
flabel metal2 s 2360 0 2440 80 0 FreeSans 320 0 0 0 N1END[3]
port 161 nsew signal input
flabel metal2 s 2552 42928 2632 43008 0 FreeSans 320 0 0 0 N2BEG[0]
port 162 nsew signal output
flabel metal2 s 2744 42928 2824 43008 0 FreeSans 320 0 0 0 N2BEG[1]
port 163 nsew signal output
flabel metal2 s 2936 42928 3016 43008 0 FreeSans 320 0 0 0 N2BEG[2]
port 164 nsew signal output
flabel metal2 s 3128 42928 3208 43008 0 FreeSans 320 0 0 0 N2BEG[3]
port 165 nsew signal output
flabel metal2 s 3320 42928 3400 43008 0 FreeSans 320 0 0 0 N2BEG[4]
port 166 nsew signal output
flabel metal2 s 3512 42928 3592 43008 0 FreeSans 320 0 0 0 N2BEG[5]
port 167 nsew signal output
flabel metal2 s 3704 42928 3784 43008 0 FreeSans 320 0 0 0 N2BEG[6]
port 168 nsew signal output
flabel metal2 s 3896 42928 3976 43008 0 FreeSans 320 0 0 0 N2BEG[7]
port 169 nsew signal output
flabel metal2 s 4088 42928 4168 43008 0 FreeSans 320 0 0 0 N2BEGb[0]
port 170 nsew signal output
flabel metal2 s 4280 42928 4360 43008 0 FreeSans 320 0 0 0 N2BEGb[1]
port 171 nsew signal output
flabel metal2 s 4472 42928 4552 43008 0 FreeSans 320 0 0 0 N2BEGb[2]
port 172 nsew signal output
flabel metal2 s 4664 42928 4744 43008 0 FreeSans 320 0 0 0 N2BEGb[3]
port 173 nsew signal output
flabel metal2 s 4856 42928 4936 43008 0 FreeSans 320 0 0 0 N2BEGb[4]
port 174 nsew signal output
flabel metal2 s 5048 42928 5128 43008 0 FreeSans 320 0 0 0 N2BEGb[5]
port 175 nsew signal output
flabel metal2 s 5240 42928 5320 43008 0 FreeSans 320 0 0 0 N2BEGb[6]
port 176 nsew signal output
flabel metal2 s 5432 42928 5512 43008 0 FreeSans 320 0 0 0 N2BEGb[7]
port 177 nsew signal output
flabel metal2 s 4088 0 4168 80 0 FreeSans 320 0 0 0 N2END[0]
port 178 nsew signal input
flabel metal2 s 4280 0 4360 80 0 FreeSans 320 0 0 0 N2END[1]
port 179 nsew signal input
flabel metal2 s 4472 0 4552 80 0 FreeSans 320 0 0 0 N2END[2]
port 180 nsew signal input
flabel metal2 s 4664 0 4744 80 0 FreeSans 320 0 0 0 N2END[3]
port 181 nsew signal input
flabel metal2 s 4856 0 4936 80 0 FreeSans 320 0 0 0 N2END[4]
port 182 nsew signal input
flabel metal2 s 5048 0 5128 80 0 FreeSans 320 0 0 0 N2END[5]
port 183 nsew signal input
flabel metal2 s 5240 0 5320 80 0 FreeSans 320 0 0 0 N2END[6]
port 184 nsew signal input
flabel metal2 s 5432 0 5512 80 0 FreeSans 320 0 0 0 N2END[7]
port 185 nsew signal input
flabel metal2 s 2552 0 2632 80 0 FreeSans 320 0 0 0 N2MID[0]
port 186 nsew signal input
flabel metal2 s 2744 0 2824 80 0 FreeSans 320 0 0 0 N2MID[1]
port 187 nsew signal input
flabel metal2 s 2936 0 3016 80 0 FreeSans 320 0 0 0 N2MID[2]
port 188 nsew signal input
flabel metal2 s 3128 0 3208 80 0 FreeSans 320 0 0 0 N2MID[3]
port 189 nsew signal input
flabel metal2 s 3320 0 3400 80 0 FreeSans 320 0 0 0 N2MID[4]
port 190 nsew signal input
flabel metal2 s 3512 0 3592 80 0 FreeSans 320 0 0 0 N2MID[5]
port 191 nsew signal input
flabel metal2 s 3704 0 3784 80 0 FreeSans 320 0 0 0 N2MID[6]
port 192 nsew signal input
flabel metal2 s 3896 0 3976 80 0 FreeSans 320 0 0 0 N2MID[7]
port 193 nsew signal input
flabel metal2 s 5624 42928 5704 43008 0 FreeSans 320 0 0 0 N4BEG[0]
port 194 nsew signal output
flabel metal2 s 7544 42928 7624 43008 0 FreeSans 320 0 0 0 N4BEG[10]
port 195 nsew signal output
flabel metal2 s 7736 42928 7816 43008 0 FreeSans 320 0 0 0 N4BEG[11]
port 196 nsew signal output
flabel metal2 s 7928 42928 8008 43008 0 FreeSans 320 0 0 0 N4BEG[12]
port 197 nsew signal output
flabel metal2 s 8120 42928 8200 43008 0 FreeSans 320 0 0 0 N4BEG[13]
port 198 nsew signal output
flabel metal2 s 8312 42928 8392 43008 0 FreeSans 320 0 0 0 N4BEG[14]
port 199 nsew signal output
flabel metal2 s 8504 42928 8584 43008 0 FreeSans 320 0 0 0 N4BEG[15]
port 200 nsew signal output
flabel metal2 s 5816 42928 5896 43008 0 FreeSans 320 0 0 0 N4BEG[1]
port 201 nsew signal output
flabel metal2 s 6008 42928 6088 43008 0 FreeSans 320 0 0 0 N4BEG[2]
port 202 nsew signal output
flabel metal2 s 6200 42928 6280 43008 0 FreeSans 320 0 0 0 N4BEG[3]
port 203 nsew signal output
flabel metal2 s 6392 42928 6472 43008 0 FreeSans 320 0 0 0 N4BEG[4]
port 204 nsew signal output
flabel metal2 s 6584 42928 6664 43008 0 FreeSans 320 0 0 0 N4BEG[5]
port 205 nsew signal output
flabel metal2 s 6776 42928 6856 43008 0 FreeSans 320 0 0 0 N4BEG[6]
port 206 nsew signal output
flabel metal2 s 6968 42928 7048 43008 0 FreeSans 320 0 0 0 N4BEG[7]
port 207 nsew signal output
flabel metal2 s 7160 42928 7240 43008 0 FreeSans 320 0 0 0 N4BEG[8]
port 208 nsew signal output
flabel metal2 s 7352 42928 7432 43008 0 FreeSans 320 0 0 0 N4BEG[9]
port 209 nsew signal output
flabel metal2 s 5624 0 5704 80 0 FreeSans 320 0 0 0 N4END[0]
port 210 nsew signal input
flabel metal2 s 7544 0 7624 80 0 FreeSans 320 0 0 0 N4END[10]
port 211 nsew signal input
flabel metal2 s 7736 0 7816 80 0 FreeSans 320 0 0 0 N4END[11]
port 212 nsew signal input
flabel metal2 s 7928 0 8008 80 0 FreeSans 320 0 0 0 N4END[12]
port 213 nsew signal input
flabel metal2 s 8120 0 8200 80 0 FreeSans 320 0 0 0 N4END[13]
port 214 nsew signal input
flabel metal2 s 8312 0 8392 80 0 FreeSans 320 0 0 0 N4END[14]
port 215 nsew signal input
flabel metal2 s 8504 0 8584 80 0 FreeSans 320 0 0 0 N4END[15]
port 216 nsew signal input
flabel metal2 s 5816 0 5896 80 0 FreeSans 320 0 0 0 N4END[1]
port 217 nsew signal input
flabel metal2 s 6008 0 6088 80 0 FreeSans 320 0 0 0 N4END[2]
port 218 nsew signal input
flabel metal2 s 6200 0 6280 80 0 FreeSans 320 0 0 0 N4END[3]
port 219 nsew signal input
flabel metal2 s 6392 0 6472 80 0 FreeSans 320 0 0 0 N4END[4]
port 220 nsew signal input
flabel metal2 s 6584 0 6664 80 0 FreeSans 320 0 0 0 N4END[5]
port 221 nsew signal input
flabel metal2 s 6776 0 6856 80 0 FreeSans 320 0 0 0 N4END[6]
port 222 nsew signal input
flabel metal2 s 6968 0 7048 80 0 FreeSans 320 0 0 0 N4END[7]
port 223 nsew signal input
flabel metal2 s 7160 0 7240 80 0 FreeSans 320 0 0 0 N4END[8]
port 224 nsew signal input
flabel metal2 s 7352 0 7432 80 0 FreeSans 320 0 0 0 N4END[9]
port 225 nsew signal input
flabel metal3 s 21424 23900 21504 23980 0 FreeSans 320 0 0 0 RST_N_TT_PROJECT
port 226 nsew signal output
flabel metal2 s 8696 0 8776 80 0 FreeSans 320 0 0 0 S1BEG[0]
port 227 nsew signal output
flabel metal2 s 8888 0 8968 80 0 FreeSans 320 0 0 0 S1BEG[1]
port 228 nsew signal output
flabel metal2 s 9080 0 9160 80 0 FreeSans 320 0 0 0 S1BEG[2]
port 229 nsew signal output
flabel metal2 s 9272 0 9352 80 0 FreeSans 320 0 0 0 S1BEG[3]
port 230 nsew signal output
flabel metal2 s 8696 42928 8776 43008 0 FreeSans 320 0 0 0 S1END[0]
port 231 nsew signal input
flabel metal2 s 8888 42928 8968 43008 0 FreeSans 320 0 0 0 S1END[1]
port 232 nsew signal input
flabel metal2 s 9080 42928 9160 43008 0 FreeSans 320 0 0 0 S1END[2]
port 233 nsew signal input
flabel metal2 s 9272 42928 9352 43008 0 FreeSans 320 0 0 0 S1END[3]
port 234 nsew signal input
flabel metal2 s 9464 0 9544 80 0 FreeSans 320 0 0 0 S2BEG[0]
port 235 nsew signal output
flabel metal2 s 9656 0 9736 80 0 FreeSans 320 0 0 0 S2BEG[1]
port 236 nsew signal output
flabel metal2 s 9848 0 9928 80 0 FreeSans 320 0 0 0 S2BEG[2]
port 237 nsew signal output
flabel metal2 s 10040 0 10120 80 0 FreeSans 320 0 0 0 S2BEG[3]
port 238 nsew signal output
flabel metal2 s 10232 0 10312 80 0 FreeSans 320 0 0 0 S2BEG[4]
port 239 nsew signal output
flabel metal2 s 10424 0 10504 80 0 FreeSans 320 0 0 0 S2BEG[5]
port 240 nsew signal output
flabel metal2 s 10616 0 10696 80 0 FreeSans 320 0 0 0 S2BEG[6]
port 241 nsew signal output
flabel metal2 s 10808 0 10888 80 0 FreeSans 320 0 0 0 S2BEG[7]
port 242 nsew signal output
flabel metal2 s 11000 0 11080 80 0 FreeSans 320 0 0 0 S2BEGb[0]
port 243 nsew signal output
flabel metal2 s 11192 0 11272 80 0 FreeSans 320 0 0 0 S2BEGb[1]
port 244 nsew signal output
flabel metal2 s 11384 0 11464 80 0 FreeSans 320 0 0 0 S2BEGb[2]
port 245 nsew signal output
flabel metal2 s 11576 0 11656 80 0 FreeSans 320 0 0 0 S2BEGb[3]
port 246 nsew signal output
flabel metal2 s 11768 0 11848 80 0 FreeSans 320 0 0 0 S2BEGb[4]
port 247 nsew signal output
flabel metal2 s 11960 0 12040 80 0 FreeSans 320 0 0 0 S2BEGb[5]
port 248 nsew signal output
flabel metal2 s 12152 0 12232 80 0 FreeSans 320 0 0 0 S2BEGb[6]
port 249 nsew signal output
flabel metal2 s 12344 0 12424 80 0 FreeSans 320 0 0 0 S2BEGb[7]
port 250 nsew signal output
flabel metal2 s 11000 42928 11080 43008 0 FreeSans 320 0 0 0 S2END[0]
port 251 nsew signal input
flabel metal2 s 11192 42928 11272 43008 0 FreeSans 320 0 0 0 S2END[1]
port 252 nsew signal input
flabel metal2 s 11384 42928 11464 43008 0 FreeSans 320 0 0 0 S2END[2]
port 253 nsew signal input
flabel metal2 s 11576 42928 11656 43008 0 FreeSans 320 0 0 0 S2END[3]
port 254 nsew signal input
flabel metal2 s 11768 42928 11848 43008 0 FreeSans 320 0 0 0 S2END[4]
port 255 nsew signal input
flabel metal2 s 11960 42928 12040 43008 0 FreeSans 320 0 0 0 S2END[5]
port 256 nsew signal input
flabel metal2 s 12152 42928 12232 43008 0 FreeSans 320 0 0 0 S2END[6]
port 257 nsew signal input
flabel metal2 s 12344 42928 12424 43008 0 FreeSans 320 0 0 0 S2END[7]
port 258 nsew signal input
flabel metal2 s 9464 42928 9544 43008 0 FreeSans 320 0 0 0 S2MID[0]
port 259 nsew signal input
flabel metal2 s 9656 42928 9736 43008 0 FreeSans 320 0 0 0 S2MID[1]
port 260 nsew signal input
flabel metal2 s 9848 42928 9928 43008 0 FreeSans 320 0 0 0 S2MID[2]
port 261 nsew signal input
flabel metal2 s 10040 42928 10120 43008 0 FreeSans 320 0 0 0 S2MID[3]
port 262 nsew signal input
flabel metal2 s 10232 42928 10312 43008 0 FreeSans 320 0 0 0 S2MID[4]
port 263 nsew signal input
flabel metal2 s 10424 42928 10504 43008 0 FreeSans 320 0 0 0 S2MID[5]
port 264 nsew signal input
flabel metal2 s 10616 42928 10696 43008 0 FreeSans 320 0 0 0 S2MID[6]
port 265 nsew signal input
flabel metal2 s 10808 42928 10888 43008 0 FreeSans 320 0 0 0 S2MID[7]
port 266 nsew signal input
flabel metal2 s 12536 0 12616 80 0 FreeSans 320 0 0 0 S4BEG[0]
port 267 nsew signal output
flabel metal2 s 14456 0 14536 80 0 FreeSans 320 0 0 0 S4BEG[10]
port 268 nsew signal output
flabel metal2 s 14648 0 14728 80 0 FreeSans 320 0 0 0 S4BEG[11]
port 269 nsew signal output
flabel metal2 s 14840 0 14920 80 0 FreeSans 320 0 0 0 S4BEG[12]
port 270 nsew signal output
flabel metal2 s 15032 0 15112 80 0 FreeSans 320 0 0 0 S4BEG[13]
port 271 nsew signal output
flabel metal2 s 15224 0 15304 80 0 FreeSans 320 0 0 0 S4BEG[14]
port 272 nsew signal output
flabel metal2 s 15416 0 15496 80 0 FreeSans 320 0 0 0 S4BEG[15]
port 273 nsew signal output
flabel metal2 s 12728 0 12808 80 0 FreeSans 320 0 0 0 S4BEG[1]
port 274 nsew signal output
flabel metal2 s 12920 0 13000 80 0 FreeSans 320 0 0 0 S4BEG[2]
port 275 nsew signal output
flabel metal2 s 13112 0 13192 80 0 FreeSans 320 0 0 0 S4BEG[3]
port 276 nsew signal output
flabel metal2 s 13304 0 13384 80 0 FreeSans 320 0 0 0 S4BEG[4]
port 277 nsew signal output
flabel metal2 s 13496 0 13576 80 0 FreeSans 320 0 0 0 S4BEG[5]
port 278 nsew signal output
flabel metal2 s 13688 0 13768 80 0 FreeSans 320 0 0 0 S4BEG[6]
port 279 nsew signal output
flabel metal2 s 13880 0 13960 80 0 FreeSans 320 0 0 0 S4BEG[7]
port 280 nsew signal output
flabel metal2 s 14072 0 14152 80 0 FreeSans 320 0 0 0 S4BEG[8]
port 281 nsew signal output
flabel metal2 s 14264 0 14344 80 0 FreeSans 320 0 0 0 S4BEG[9]
port 282 nsew signal output
flabel metal2 s 12536 42928 12616 43008 0 FreeSans 320 0 0 0 S4END[0]
port 283 nsew signal input
flabel metal2 s 14456 42928 14536 43008 0 FreeSans 320 0 0 0 S4END[10]
port 284 nsew signal input
flabel metal2 s 14648 42928 14728 43008 0 FreeSans 320 0 0 0 S4END[11]
port 285 nsew signal input
flabel metal2 s 14840 42928 14920 43008 0 FreeSans 320 0 0 0 S4END[12]
port 286 nsew signal input
flabel metal2 s 15032 42928 15112 43008 0 FreeSans 320 0 0 0 S4END[13]
port 287 nsew signal input
flabel metal2 s 15224 42928 15304 43008 0 FreeSans 320 0 0 0 S4END[14]
port 288 nsew signal input
flabel metal2 s 15416 42928 15496 43008 0 FreeSans 320 0 0 0 S4END[15]
port 289 nsew signal input
flabel metal2 s 12728 42928 12808 43008 0 FreeSans 320 0 0 0 S4END[1]
port 290 nsew signal input
flabel metal2 s 12920 42928 13000 43008 0 FreeSans 320 0 0 0 S4END[2]
port 291 nsew signal input
flabel metal2 s 13112 42928 13192 43008 0 FreeSans 320 0 0 0 S4END[3]
port 292 nsew signal input
flabel metal2 s 13304 42928 13384 43008 0 FreeSans 320 0 0 0 S4END[4]
port 293 nsew signal input
flabel metal2 s 13496 42928 13576 43008 0 FreeSans 320 0 0 0 S4END[5]
port 294 nsew signal input
flabel metal2 s 13688 42928 13768 43008 0 FreeSans 320 0 0 0 S4END[6]
port 295 nsew signal input
flabel metal2 s 13880 42928 13960 43008 0 FreeSans 320 0 0 0 S4END[7]
port 296 nsew signal input
flabel metal2 s 14072 42928 14152 43008 0 FreeSans 320 0 0 0 S4END[8]
port 297 nsew signal input
flabel metal2 s 14264 42928 14344 43008 0 FreeSans 320 0 0 0 S4END[9]
port 298 nsew signal input
flabel metal3 s 21424 18860 21504 18940 0 FreeSans 320 0 0 0 UIO_IN_TT_PROJECT0
port 299 nsew signal output
flabel metal3 s 21424 19364 21504 19444 0 FreeSans 320 0 0 0 UIO_IN_TT_PROJECT1
port 300 nsew signal output
flabel metal3 s 21424 19868 21504 19948 0 FreeSans 320 0 0 0 UIO_IN_TT_PROJECT2
port 301 nsew signal output
flabel metal3 s 21424 20372 21504 20452 0 FreeSans 320 0 0 0 UIO_IN_TT_PROJECT3
port 302 nsew signal output
flabel metal3 s 21424 20876 21504 20956 0 FreeSans 320 0 0 0 UIO_IN_TT_PROJECT4
port 303 nsew signal output
flabel metal3 s 21424 21380 21504 21460 0 FreeSans 320 0 0 0 UIO_IN_TT_PROJECT5
port 304 nsew signal output
flabel metal3 s 21424 21884 21504 21964 0 FreeSans 320 0 0 0 UIO_IN_TT_PROJECT6
port 305 nsew signal output
flabel metal3 s 21424 22388 21504 22468 0 FreeSans 320 0 0 0 UIO_IN_TT_PROJECT7
port 306 nsew signal output
flabel metal3 s 21424 10796 21504 10876 0 FreeSans 320 0 0 0 UIO_OE_TT_PROJECT0
port 307 nsew signal input
flabel metal3 s 21424 11300 21504 11380 0 FreeSans 320 0 0 0 UIO_OE_TT_PROJECT1
port 308 nsew signal input
flabel metal3 s 21424 11804 21504 11884 0 FreeSans 320 0 0 0 UIO_OE_TT_PROJECT2
port 309 nsew signal input
flabel metal3 s 21424 12308 21504 12388 0 FreeSans 320 0 0 0 UIO_OE_TT_PROJECT3
port 310 nsew signal input
flabel metal3 s 21424 12812 21504 12892 0 FreeSans 320 0 0 0 UIO_OE_TT_PROJECT4
port 311 nsew signal input
flabel metal3 s 21424 13316 21504 13396 0 FreeSans 320 0 0 0 UIO_OE_TT_PROJECT5
port 312 nsew signal input
flabel metal3 s 21424 13820 21504 13900 0 FreeSans 320 0 0 0 UIO_OE_TT_PROJECT6
port 313 nsew signal input
flabel metal3 s 21424 14324 21504 14404 0 FreeSans 320 0 0 0 UIO_OE_TT_PROJECT7
port 314 nsew signal input
flabel metal3 s 21424 6764 21504 6844 0 FreeSans 320 0 0 0 UIO_OUT_TT_PROJECT0
port 315 nsew signal input
flabel metal3 s 21424 7268 21504 7348 0 FreeSans 320 0 0 0 UIO_OUT_TT_PROJECT1
port 316 nsew signal input
flabel metal3 s 21424 7772 21504 7852 0 FreeSans 320 0 0 0 UIO_OUT_TT_PROJECT2
port 317 nsew signal input
flabel metal3 s 21424 8276 21504 8356 0 FreeSans 320 0 0 0 UIO_OUT_TT_PROJECT3
port 318 nsew signal input
flabel metal3 s 21424 8780 21504 8860 0 FreeSans 320 0 0 0 UIO_OUT_TT_PROJECT4
port 319 nsew signal input
flabel metal3 s 21424 9284 21504 9364 0 FreeSans 320 0 0 0 UIO_OUT_TT_PROJECT5
port 320 nsew signal input
flabel metal3 s 21424 9788 21504 9868 0 FreeSans 320 0 0 0 UIO_OUT_TT_PROJECT6
port 321 nsew signal input
flabel metal3 s 21424 10292 21504 10372 0 FreeSans 320 0 0 0 UIO_OUT_TT_PROJECT7
port 322 nsew signal input
flabel metal3 s 21424 14828 21504 14908 0 FreeSans 320 0 0 0 UI_IN_TT_PROJECT0
port 323 nsew signal output
flabel metal3 s 21424 15332 21504 15412 0 FreeSans 320 0 0 0 UI_IN_TT_PROJECT1
port 324 nsew signal output
flabel metal3 s 21424 15836 21504 15916 0 FreeSans 320 0 0 0 UI_IN_TT_PROJECT2
port 325 nsew signal output
flabel metal3 s 21424 16340 21504 16420 0 FreeSans 320 0 0 0 UI_IN_TT_PROJECT3
port 326 nsew signal output
flabel metal3 s 21424 16844 21504 16924 0 FreeSans 320 0 0 0 UI_IN_TT_PROJECT4
port 327 nsew signal output
flabel metal3 s 21424 17348 21504 17428 0 FreeSans 320 0 0 0 UI_IN_TT_PROJECT5
port 328 nsew signal output
flabel metal3 s 21424 17852 21504 17932 0 FreeSans 320 0 0 0 UI_IN_TT_PROJECT6
port 329 nsew signal output
flabel metal3 s 21424 18356 21504 18436 0 FreeSans 320 0 0 0 UI_IN_TT_PROJECT7
port 330 nsew signal output
flabel metal3 s 21424 2732 21504 2812 0 FreeSans 320 0 0 0 UO_OUT_TT_PROJECT0
port 331 nsew signal input
flabel metal3 s 21424 3236 21504 3316 0 FreeSans 320 0 0 0 UO_OUT_TT_PROJECT1
port 332 nsew signal input
flabel metal3 s 21424 3740 21504 3820 0 FreeSans 320 0 0 0 UO_OUT_TT_PROJECT2
port 333 nsew signal input
flabel metal3 s 21424 4244 21504 4324 0 FreeSans 320 0 0 0 UO_OUT_TT_PROJECT3
port 334 nsew signal input
flabel metal3 s 21424 4748 21504 4828 0 FreeSans 320 0 0 0 UO_OUT_TT_PROJECT4
port 335 nsew signal input
flabel metal3 s 21424 5252 21504 5332 0 FreeSans 320 0 0 0 UO_OUT_TT_PROJECT5
port 336 nsew signal input
flabel metal3 s 21424 5756 21504 5836 0 FreeSans 320 0 0 0 UO_OUT_TT_PROJECT6
port 337 nsew signal input
flabel metal3 s 21424 6260 21504 6340 0 FreeSans 320 0 0 0 UO_OUT_TT_PROJECT7
port 338 nsew signal input
flabel metal2 s 15608 0 15688 80 0 FreeSans 320 0 0 0 UserCLK
port 339 nsew signal input
flabel metal2 s 15608 42928 15688 43008 0 FreeSans 320 0 0 0 UserCLKo
port 340 nsew signal output
flabel metal6 s 4892 0 5332 43008 0 FreeSans 2624 90 0 0 VGND
port 341 nsew ground bidirectional
flabel metal6 s 4892 0 5332 328 0 FreeSans 2624 0 0 0 VGND
port 341 nsew ground bidirectional
flabel metal6 s 4892 42680 5332 43008 0 FreeSans 2624 0 0 0 VGND
port 341 nsew ground bidirectional
flabel metal6 s 20012 0 20452 43008 0 FreeSans 2624 90 0 0 VGND
port 341 nsew ground bidirectional
flabel metal6 s 20012 0 20452 328 0 FreeSans 2624 0 0 0 VGND
port 341 nsew ground bidirectional
flabel metal6 s 20012 42680 20452 43008 0 FreeSans 2624 0 0 0 VGND
port 341 nsew ground bidirectional
flabel metal6 s 3652 0 4092 43008 0 FreeSans 2624 90 0 0 VPWR
port 342 nsew power bidirectional
flabel metal6 s 3652 0 4092 328 0 FreeSans 2624 0 0 0 VPWR
port 342 nsew power bidirectional
flabel metal6 s 3652 42680 4092 43008 0 FreeSans 2624 0 0 0 VPWR
port 342 nsew power bidirectional
flabel metal6 s 18772 0 19212 43008 0 FreeSans 2624 90 0 0 VPWR
port 342 nsew power bidirectional
flabel metal6 s 18772 0 19212 328 0 FreeSans 2624 0 0 0 VPWR
port 342 nsew power bidirectional
flabel metal6 s 18772 42680 19212 43008 0 FreeSans 2624 0 0 0 VPWR
port 342 nsew power bidirectional
flabel metal3 s 0 44 80 124 0 FreeSans 320 0 0 0 W1BEG[0]
port 343 nsew signal output
flabel metal3 s 0 380 80 460 0 FreeSans 320 0 0 0 W1BEG[1]
port 344 nsew signal output
flabel metal3 s 0 716 80 796 0 FreeSans 320 0 0 0 W1BEG[2]
port 345 nsew signal output
flabel metal3 s 0 1052 80 1132 0 FreeSans 320 0 0 0 W1BEG[3]
port 346 nsew signal output
flabel metal3 s 0 1388 80 1468 0 FreeSans 320 0 0 0 W2BEG[0]
port 347 nsew signal output
flabel metal3 s 0 1724 80 1804 0 FreeSans 320 0 0 0 W2BEG[1]
port 348 nsew signal output
flabel metal3 s 0 2060 80 2140 0 FreeSans 320 0 0 0 W2BEG[2]
port 349 nsew signal output
flabel metal3 s 0 2396 80 2476 0 FreeSans 320 0 0 0 W2BEG[3]
port 350 nsew signal output
flabel metal3 s 0 2732 80 2812 0 FreeSans 320 0 0 0 W2BEG[4]
port 351 nsew signal output
flabel metal3 s 0 3068 80 3148 0 FreeSans 320 0 0 0 W2BEG[5]
port 352 nsew signal output
flabel metal3 s 0 3404 80 3484 0 FreeSans 320 0 0 0 W2BEG[6]
port 353 nsew signal output
flabel metal3 s 0 3740 80 3820 0 FreeSans 320 0 0 0 W2BEG[7]
port 354 nsew signal output
flabel metal3 s 0 4076 80 4156 0 FreeSans 320 0 0 0 W2BEGb[0]
port 355 nsew signal output
flabel metal3 s 0 4412 80 4492 0 FreeSans 320 0 0 0 W2BEGb[1]
port 356 nsew signal output
flabel metal3 s 0 4748 80 4828 0 FreeSans 320 0 0 0 W2BEGb[2]
port 357 nsew signal output
flabel metal3 s 0 5084 80 5164 0 FreeSans 320 0 0 0 W2BEGb[3]
port 358 nsew signal output
flabel metal3 s 0 5420 80 5500 0 FreeSans 320 0 0 0 W2BEGb[4]
port 359 nsew signal output
flabel metal3 s 0 5756 80 5836 0 FreeSans 320 0 0 0 W2BEGb[5]
port 360 nsew signal output
flabel metal3 s 0 6092 80 6172 0 FreeSans 320 0 0 0 W2BEGb[6]
port 361 nsew signal output
flabel metal3 s 0 6428 80 6508 0 FreeSans 320 0 0 0 W2BEGb[7]
port 362 nsew signal output
flabel metal3 s 0 12140 80 12220 0 FreeSans 320 0 0 0 W6BEG[0]
port 363 nsew signal output
flabel metal3 s 0 15500 80 15580 0 FreeSans 320 0 0 0 W6BEG[10]
port 364 nsew signal output
flabel metal3 s 0 15836 80 15916 0 FreeSans 320 0 0 0 W6BEG[11]
port 365 nsew signal output
flabel metal3 s 0 12476 80 12556 0 FreeSans 320 0 0 0 W6BEG[1]
port 366 nsew signal output
flabel metal3 s 0 12812 80 12892 0 FreeSans 320 0 0 0 W6BEG[2]
port 367 nsew signal output
flabel metal3 s 0 13148 80 13228 0 FreeSans 320 0 0 0 W6BEG[3]
port 368 nsew signal output
flabel metal3 s 0 13484 80 13564 0 FreeSans 320 0 0 0 W6BEG[4]
port 369 nsew signal output
flabel metal3 s 0 13820 80 13900 0 FreeSans 320 0 0 0 W6BEG[5]
port 370 nsew signal output
flabel metal3 s 0 14156 80 14236 0 FreeSans 320 0 0 0 W6BEG[6]
port 371 nsew signal output
flabel metal3 s 0 14492 80 14572 0 FreeSans 320 0 0 0 W6BEG[7]
port 372 nsew signal output
flabel metal3 s 0 14828 80 14908 0 FreeSans 320 0 0 0 W6BEG[8]
port 373 nsew signal output
flabel metal3 s 0 15164 80 15244 0 FreeSans 320 0 0 0 W6BEG[9]
port 374 nsew signal output
flabel metal3 s 0 6764 80 6844 0 FreeSans 320 0 0 0 WW4BEG[0]
port 375 nsew signal output
flabel metal3 s 0 10124 80 10204 0 FreeSans 320 0 0 0 WW4BEG[10]
port 376 nsew signal output
flabel metal3 s 0 10460 80 10540 0 FreeSans 320 0 0 0 WW4BEG[11]
port 377 nsew signal output
flabel metal3 s 0 10796 80 10876 0 FreeSans 320 0 0 0 WW4BEG[12]
port 378 nsew signal output
flabel metal3 s 0 11132 80 11212 0 FreeSans 320 0 0 0 WW4BEG[13]
port 379 nsew signal output
flabel metal3 s 0 11468 80 11548 0 FreeSans 320 0 0 0 WW4BEG[14]
port 380 nsew signal output
flabel metal3 s 0 11804 80 11884 0 FreeSans 320 0 0 0 WW4BEG[15]
port 381 nsew signal output
flabel metal3 s 0 7100 80 7180 0 FreeSans 320 0 0 0 WW4BEG[1]
port 382 nsew signal output
flabel metal3 s 0 7436 80 7516 0 FreeSans 320 0 0 0 WW4BEG[2]
port 383 nsew signal output
flabel metal3 s 0 7772 80 7852 0 FreeSans 320 0 0 0 WW4BEG[3]
port 384 nsew signal output
flabel metal3 s 0 8108 80 8188 0 FreeSans 320 0 0 0 WW4BEG[4]
port 385 nsew signal output
flabel metal3 s 0 8444 80 8524 0 FreeSans 320 0 0 0 WW4BEG[5]
port 386 nsew signal output
flabel metal3 s 0 8780 80 8860 0 FreeSans 320 0 0 0 WW4BEG[6]
port 387 nsew signal output
flabel metal3 s 0 9116 80 9196 0 FreeSans 320 0 0 0 WW4BEG[7]
port 388 nsew signal output
flabel metal3 s 0 9452 80 9532 0 FreeSans 320 0 0 0 WW4BEG[8]
port 389 nsew signal output
flabel metal3 s 0 9788 80 9868 0 FreeSans 320 0 0 0 WW4BEG[9]
port 390 nsew signal output
rlabel metal1 10802 41580 10802 41580 0 VGND
rlabel metal1 10752 40824 10752 40824 0 VPWR
rlabel metal3 21378 23436 21378 23436 0 CLK_TT_PROJECT
rlabel metal3 1440 16296 1440 16296 0 E1END[0]
rlabel metal3 11616 18816 11616 18816 0 E1END[1]
rlabel metal2 15456 35658 15456 35658 0 E1END[2]
rlabel metal2 7296 17472 7296 17472 0 E1END[3]
rlabel metal2 2208 18690 2208 18690 0 E2END[0]
rlabel metal2 12288 33180 12288 33180 0 E2END[1]
rlabel metal2 18624 34986 18624 34986 0 E2END[2]
rlabel metal2 9024 35784 9024 35784 0 E2END[3]
rlabel metal2 8160 33852 8160 33852 0 E2END[4]
rlabel metal3 1182 21924 1182 21924 0 E2END[5]
rlabel metal3 1230 22260 1230 22260 0 E2END[6]
rlabel metal3 1230 22596 1230 22596 0 E2END[7]
rlabel metal2 2496 18480 2496 18480 0 E2MID[0]
rlabel metal2 11520 19950 11520 19950 0 E2MID[1]
rlabel metal3 654 18228 654 18228 0 E2MID[2]
rlabel metal2 2400 37170 2400 37170 0 E2MID[3]
rlabel metal3 1344 18984 1344 18984 0 E2MID[4]
rlabel metal2 17472 20580 17472 20580 0 E2MID[5]
rlabel metal2 17856 23226 17856 23226 0 E2MID[6]
rlabel metal3 942 19908 942 19908 0 E2MID[7]
rlabel metal2 2064 19404 2064 19404 0 E6END[0]
rlabel metal2 11808 35154 11808 35154 0 E6END[10]
rlabel metal2 6528 31710 6528 31710 0 E6END[11]
rlabel metal2 15264 31374 15264 31374 0 E6END[1]
rlabel metal2 2496 39438 2496 39438 0 E6END[2]
rlabel metal2 5952 32382 5952 32382 0 E6END[3]
rlabel metal3 126 29652 126 29652 0 E6END[4]
rlabel metal3 17424 20076 17424 20076 0 E6END[5]
rlabel metal2 1920 35448 1920 35448 0 E6END[6]
rlabel metal3 1872 28392 1872 28392 0 E6END[7]
rlabel metal3 1374 30996 1374 30996 0 E6END[8]
rlabel metal2 14832 29064 14832 29064 0 E6END[9]
rlabel metal2 1152 21882 1152 21882 0 EE4END[0]
rlabel metal3 558 26292 558 26292 0 EE4END[10]
rlabel metal3 1290 26628 1290 26628 0 EE4END[11]
rlabel metal3 3534 26964 3534 26964 0 EE4END[12]
rlabel metal2 17376 25494 17376 25494 0 EE4END[13]
rlabel metal3 702 27636 702 27636 0 EE4END[14]
rlabel metal2 4512 28224 4512 28224 0 EE4END[15]
rlabel metal3 7680 23394 7680 23394 0 EE4END[1]
rlabel via2 78 23604 78 23604 0 EE4END[2]
rlabel metal3 480 23898 480 23898 0 EE4END[3]
rlabel metal2 6528 24066 6528 24066 0 EE4END[4]
rlabel metal3 1038 24612 1038 24612 0 EE4END[5]
rlabel metal3 126 24948 126 24948 0 EE4END[6]
rlabel metal3 2208 25326 2208 25326 0 EE4END[7]
rlabel metal3 558 25620 558 25620 0 EE4END[8]
rlabel metal3 990 25956 990 25956 0 EE4END[9]
rlabel metal2 18816 23268 18816 23268 0 ENA_TT_PROJECT
rlabel metal2 2208 7854 2208 7854 0 FrameData[0]
rlabel metal2 15168 36750 15168 36750 0 FrameData[10]
rlabel metal2 17376 19194 17376 19194 0 FrameData[11]
rlabel metal2 17184 19068 17184 19068 0 FrameData[12]
rlabel metal2 20256 17850 20256 17850 0 FrameData[13]
rlabel metal3 606 37044 606 37044 0 FrameData[14]
rlabel metal3 12624 19992 12624 19992 0 FrameData[15]
rlabel metal2 1536 10752 1536 10752 0 FrameData[16]
rlabel metal2 1344 15540 1344 15540 0 FrameData[17]
rlabel metal2 1344 17976 1344 17976 0 FrameData[18]
rlabel metal2 2400 16254 2400 16254 0 FrameData[19]
rlabel metal2 1296 5628 1296 5628 0 FrameData[1]
rlabel metal2 1152 39270 1152 39270 0 FrameData[20]
rlabel metal3 1086 39396 1086 39396 0 FrameData[21]
rlabel metal2 12480 2100 12480 2100 0 FrameData[22]
rlabel metal3 1182 40068 1182 40068 0 FrameData[23]
rlabel metal3 2112 4914 2112 4914 0 FrameData[24]
rlabel metal2 1344 4368 1344 4368 0 FrameData[25]
rlabel metal3 12576 31332 12576 31332 0 FrameData[26]
rlabel metal2 11952 17052 11952 17052 0 FrameData[27]
rlabel metal2 12192 15330 12192 15330 0 FrameData[28]
rlabel metal3 13440 14028 13440 14028 0 FrameData[29]
rlabel metal3 510 33012 510 33012 0 FrameData[2]
rlabel metal2 11616 12390 11616 12390 0 FrameData[30]
rlabel metal3 846 42756 846 42756 0 FrameData[31]
rlabel metal2 1296 23772 1296 23772 0 FrameData[3]
rlabel metal2 1632 18186 1632 18186 0 FrameData[4]
rlabel metal3 126 34020 126 34020 0 FrameData[5]
rlabel metal2 18768 29988 18768 29988 0 FrameData[6]
rlabel metal2 2496 32592 2496 32592 0 FrameData[7]
rlabel metal2 1920 9786 1920 9786 0 FrameData[8]
rlabel metal2 1440 1764 1440 1764 0 FrameData[9]
rlabel metal3 20658 24444 20658 24444 0 FrameData_O[0]
rlabel metal2 19872 30366 19872 30366 0 FrameData_O[10]
rlabel metal2 17856 30576 17856 30576 0 FrameData_O[11]
rlabel metal3 21042 30492 21042 30492 0 FrameData_O[12]
rlabel metal3 21090 30996 21090 30996 0 FrameData_O[13]
rlabel metal3 20850 31500 20850 31500 0 FrameData_O[14]
rlabel metal3 20658 32004 20658 32004 0 FrameData_O[15]
rlabel metal3 20994 32508 20994 32508 0 FrameData_O[16]
rlabel metal2 19488 32088 19488 32088 0 FrameData_O[17]
rlabel metal3 21042 33516 21042 33516 0 FrameData_O[18]
rlabel metal3 20832 38892 20832 38892 0 FrameData_O[19]
rlabel metal3 20544 24780 20544 24780 0 FrameData_O[1]
rlabel metal3 19554 34524 19554 34524 0 FrameData_O[20]
rlabel metal3 20832 38976 20832 38976 0 FrameData_O[21]
rlabel metal2 19776 38724 19776 38724 0 FrameData_O[22]
rlabel metal3 20496 38808 20496 38808 0 FrameData_O[23]
rlabel metal3 17760 36498 17760 36498 0 FrameData_O[24]
rlabel metal2 20016 40236 20016 40236 0 FrameData_O[25]
rlabel metal2 17952 40488 17952 40488 0 FrameData_O[26]
rlabel metal3 20994 38052 20994 38052 0 FrameData_O[27]
rlabel metal3 21042 38556 21042 38556 0 FrameData_O[28]
rlabel metal3 20802 39060 20802 39060 0 FrameData_O[29]
rlabel metal2 19872 25788 19872 25788 0 FrameData_O[2]
rlabel metal2 19824 39564 19824 39564 0 FrameData_O[30]
rlabel metal3 20544 40026 20544 40026 0 FrameData_O[31]
rlabel metal3 20850 25956 20850 25956 0 FrameData_O[3]
rlabel metal3 21378 26460 21378 26460 0 FrameData_O[4]
rlabel metal3 20706 26964 20706 26964 0 FrameData_O[5]
rlabel metal3 20178 27468 20178 27468 0 FrameData_O[6]
rlabel metal3 19776 29316 19776 29316 0 FrameData_O[7]
rlabel metal3 20850 28476 20850 28476 0 FrameData_O[8]
rlabel metal3 20976 29232 20976 29232 0 FrameData_O[9]
rlabel metal2 15840 324 15840 324 0 FrameStrobe[0]
rlabel metal2 17760 618 17760 618 0 FrameStrobe[10]
rlabel metal2 17952 366 17952 366 0 FrameStrobe[11]
rlabel metal2 18144 366 18144 366 0 FrameStrobe[12]
rlabel metal2 18336 366 18336 366 0 FrameStrobe[13]
rlabel metal2 18528 366 18528 366 0 FrameStrobe[14]
rlabel metal2 18720 282 18720 282 0 FrameStrobe[15]
rlabel metal2 18912 702 18912 702 0 FrameStrobe[16]
rlabel metal2 19104 660 19104 660 0 FrameStrobe[17]
rlabel metal2 19296 324 19296 324 0 FrameStrobe[18]
rlabel metal2 19488 366 19488 366 0 FrameStrobe[19]
rlabel metal2 16032 744 16032 744 0 FrameStrobe[1]
rlabel metal2 2496 20034 2496 20034 0 FrameStrobe[2]
rlabel metal2 16416 912 16416 912 0 FrameStrobe[3]
rlabel metal2 17856 13986 17856 13986 0 FrameStrobe[4]
rlabel metal2 2496 5334 2496 5334 0 FrameStrobe[5]
rlabel metal3 17136 35700 17136 35700 0 FrameStrobe[6]
rlabel metal2 2448 20748 2448 20748 0 FrameStrobe[7]
rlabel metal2 2448 38220 2448 38220 0 FrameStrobe[8]
rlabel metal2 17568 450 17568 450 0 FrameStrobe[9]
rlabel metal2 16128 40656 16128 40656 0 FrameStrobe_O[0]
rlabel metal2 17808 41412 17808 41412 0 FrameStrobe_O[10]
rlabel metal2 18528 40698 18528 40698 0 FrameStrobe_O[11]
rlabel metal2 18144 42180 18144 42180 0 FrameStrobe_O[12]
rlabel metal2 19776 41454 19776 41454 0 FrameStrobe_O[13]
rlabel metal2 18480 39900 18480 39900 0 FrameStrobe_O[14]
rlabel metal2 17856 36582 17856 36582 0 FrameStrobe_O[15]
rlabel metal2 18960 39900 18960 39900 0 FrameStrobe_O[16]
rlabel metal2 18288 37632 18288 37632 0 FrameStrobe_O[17]
rlabel metal2 11808 41160 11808 41160 0 FrameStrobe_O[18]
rlabel metal3 19104 41412 19104 41412 0 FrameStrobe_O[19]
rlabel metal2 16560 40656 16560 40656 0 FrameStrobe_O[1]
rlabel metal2 16176 41412 16176 41412 0 FrameStrobe_O[2]
rlabel metal3 16704 40656 16704 40656 0 FrameStrobe_O[3]
rlabel metal3 16608 18732 16608 18732 0 FrameStrobe_O[4]
rlabel metal2 16800 42096 16800 42096 0 FrameStrobe_O[5]
rlabel metal2 17136 41412 17136 41412 0 FrameStrobe_O[6]
rlabel metal3 18816 40656 18816 40656 0 FrameStrobe_O[7]
rlabel metal2 18912 41160 18912 41160 0 FrameStrobe_O[8]
rlabel metal3 17856 40656 17856 40656 0 FrameStrobe_O[9]
rlabel metal2 6192 6636 6192 6636 0 Inst_E_TT_IF_ConfigMem.Inst_frame0_bit0.Q
rlabel metal2 7776 6890 7776 6890 0 Inst_E_TT_IF_ConfigMem.Inst_frame0_bit1.Q
rlabel metal2 4416 36162 4416 36162 0 Inst_E_TT_IF_ConfigMem.Inst_frame0_bit10.Q
rlabel metal2 5904 35364 5904 35364 0 Inst_E_TT_IF_ConfigMem.Inst_frame0_bit11.Q
rlabel metal2 9984 37681 9984 37681 0 Inst_E_TT_IF_ConfigMem.Inst_frame0_bit12.Q
rlabel metal3 8160 37380 8160 37380 0 Inst_E_TT_IF_ConfigMem.Inst_frame0_bit13.Q
rlabel metal2 8160 36120 8160 36120 0 Inst_E_TT_IF_ConfigMem.Inst_frame0_bit14.Q
rlabel metal2 6432 36750 6432 36750 0 Inst_E_TT_IF_ConfigMem.Inst_frame0_bit15.Q
rlabel metal2 5088 37590 5088 37590 0 Inst_E_TT_IF_ConfigMem.Inst_frame0_bit16.Q
rlabel metal3 6144 38724 6144 38724 0 Inst_E_TT_IF_ConfigMem.Inst_frame0_bit17.Q
rlabel metal3 3408 38724 3408 38724 0 Inst_E_TT_IF_ConfigMem.Inst_frame0_bit18.Q
rlabel metal2 7872 40023 7872 40023 0 Inst_E_TT_IF_ConfigMem.Inst_frame0_bit19.Q
rlabel metal2 13824 18606 13824 18606 0 Inst_E_TT_IF_ConfigMem.Inst_frame0_bit2.Q
rlabel metal2 10560 38850 10560 38850 0 Inst_E_TT_IF_ConfigMem.Inst_frame0_bit20.Q
rlabel metal2 12096 38642 12096 38642 0 Inst_E_TT_IF_ConfigMem.Inst_frame0_bit21.Q
rlabel metal2 8544 39060 8544 39060 0 Inst_E_TT_IF_ConfigMem.Inst_frame0_bit22.Q
rlabel metal2 9984 40154 9984 40154 0 Inst_E_TT_IF_ConfigMem.Inst_frame0_bit23.Q
rlabel metal2 5664 15414 5664 15414 0 Inst_E_TT_IF_ConfigMem.Inst_frame0_bit24.Q
rlabel metal3 5616 15708 5616 15708 0 Inst_E_TT_IF_ConfigMem.Inst_frame0_bit25.Q
rlabel via1 14496 31330 14496 31330 0 Inst_E_TT_IF_ConfigMem.Inst_frame0_bit26.Q
rlabel metal3 14738 31332 14738 31332 0 Inst_E_TT_IF_ConfigMem.Inst_frame0_bit27.Q
rlabel metal2 12000 39900 12000 39900 0 Inst_E_TT_IF_ConfigMem.Inst_frame0_bit28.Q
rlabel metal2 12000 40362 12000 40362 0 Inst_E_TT_IF_ConfigMem.Inst_frame0_bit29.Q
rlabel metal2 15648 18186 15648 18186 0 Inst_E_TT_IF_ConfigMem.Inst_frame0_bit3.Q
rlabel metal2 5856 33390 5856 33390 0 Inst_E_TT_IF_ConfigMem.Inst_frame0_bit30.Q
rlabel metal3 4944 33852 4944 33852 0 Inst_E_TT_IF_ConfigMem.Inst_frame0_bit31.Q
rlabel metal2 13440 34272 13440 34272 0 Inst_E_TT_IF_ConfigMem.Inst_frame0_bit4.Q
rlabel metal2 15072 34104 15072 34104 0 Inst_E_TT_IF_ConfigMem.Inst_frame0_bit5.Q
rlabel metal2 10128 11928 10128 11928 0 Inst_E_TT_IF_ConfigMem.Inst_frame0_bit6.Q
rlabel metal2 12384 13734 12384 13734 0 Inst_E_TT_IF_ConfigMem.Inst_frame0_bit7.Q
rlabel metal2 8160 1974 8160 1974 0 Inst_E_TT_IF_ConfigMem.Inst_frame0_bit8.Q
rlabel metal2 9696 1631 9696 1631 0 Inst_E_TT_IF_ConfigMem.Inst_frame0_bit9.Q
rlabel metal2 5568 26502 5568 26502 0 Inst_E_TT_IF_ConfigMem.Inst_frame1_bit0.Q
rlabel metal2 5808 25536 5808 25536 0 Inst_E_TT_IF_ConfigMem.Inst_frame1_bit1.Q
rlabel metal2 14016 19488 14016 19488 0 Inst_E_TT_IF_ConfigMem.Inst_frame1_bit10.Q
rlabel via2 15552 19238 15552 19238 0 Inst_E_TT_IF_ConfigMem.Inst_frame1_bit11.Q
rlabel metal2 14208 37968 14208 37968 0 Inst_E_TT_IF_ConfigMem.Inst_frame1_bit12.Q
rlabel metal2 15720 37464 15720 37464 0 Inst_E_TT_IF_ConfigMem.Inst_frame1_bit13.Q
rlabel metal2 10176 13650 10176 13650 0 Inst_E_TT_IF_ConfigMem.Inst_frame1_bit14.Q
rlabel metal2 11712 15001 11712 15001 0 Inst_E_TT_IF_ConfigMem.Inst_frame1_bit15.Q
rlabel metal2 5664 11046 5664 11046 0 Inst_E_TT_IF_ConfigMem.Inst_frame1_bit16.Q
rlabel metal3 7104 10332 7104 10332 0 Inst_E_TT_IF_ConfigMem.Inst_frame1_bit17.Q
rlabel metal2 13632 16254 13632 16254 0 Inst_E_TT_IF_ConfigMem.Inst_frame1_bit18.Q
rlabel metal2 15312 15708 15312 15708 0 Inst_E_TT_IF_ConfigMem.Inst_frame1_bit19.Q
rlabel metal3 17424 23100 17424 23100 0 Inst_E_TT_IF_ConfigMem.Inst_frame1_bit2.Q
rlabel metal2 14064 38892 14064 38892 0 Inst_E_TT_IF_ConfigMem.Inst_frame1_bit20.Q
rlabel metal2 15648 39193 15648 39193 0 Inst_E_TT_IF_ConfigMem.Inst_frame1_bit21.Q
rlabel metal2 7200 15592 7200 15592 0 Inst_E_TT_IF_ConfigMem.Inst_frame1_bit22.Q
rlabel metal3 8352 14952 8352 14952 0 Inst_E_TT_IF_ConfigMem.Inst_frame1_bit23.Q
rlabel metal2 6096 3696 6096 3696 0 Inst_E_TT_IF_ConfigMem.Inst_frame1_bit24.Q
rlabel metal3 7344 4368 7344 4368 0 Inst_E_TT_IF_ConfigMem.Inst_frame1_bit25.Q
rlabel metal2 11904 17262 11904 17262 0 Inst_E_TT_IF_ConfigMem.Inst_frame1_bit26.Q
rlabel metal2 13584 17220 13584 17220 0 Inst_E_TT_IF_ConfigMem.Inst_frame1_bit27.Q
rlabel metal2 13344 40362 13344 40362 0 Inst_E_TT_IF_ConfigMem.Inst_frame1_bit28.Q
rlabel metal2 14880 39981 14880 39981 0 Inst_E_TT_IF_ConfigMem.Inst_frame1_bit29.Q
rlabel metal2 17328 23772 17328 23772 0 Inst_E_TT_IF_ConfigMem.Inst_frame1_bit3.Q
rlabel metal2 9600 15582 9600 15582 0 Inst_E_TT_IF_ConfigMem.Inst_frame1_bit30.Q
rlabel metal2 11232 15960 11232 15960 0 Inst_E_TT_IF_ConfigMem.Inst_frame1_bit31.Q
rlabel metal2 6624 35910 6624 35910 0 Inst_E_TT_IF_ConfigMem.Inst_frame1_bit4.Q
rlabel metal2 8640 36792 8640 36792 0 Inst_E_TT_IF_ConfigMem.Inst_frame1_bit5.Q
rlabel metal3 8304 36708 8304 36708 0 Inst_E_TT_IF_ConfigMem.Inst_frame1_bit6.Q
rlabel metal2 10032 35196 10032 35196 0 Inst_E_TT_IF_ConfigMem.Inst_frame1_bit7.Q
rlabel metal3 4992 2604 4992 2604 0 Inst_E_TT_IF_ConfigMem.Inst_frame1_bit8.Q
rlabel metal2 6816 1470 6816 1470 0 Inst_E_TT_IF_ConfigMem.Inst_frame1_bit9.Q
rlabel metal2 7680 24864 7680 24864 0 Inst_E_TT_IF_ConfigMem.Inst_frame2_bit0.Q
rlabel metal2 19344 19488 19344 19488 0 Inst_E_TT_IF_ConfigMem.Inst_frame2_bit1.Q
rlabel metal2 4128 20496 4128 20496 0 Inst_E_TT_IF_ConfigMem.Inst_frame2_bit10.Q
rlabel metal2 4272 18564 4272 18564 0 Inst_E_TT_IF_ConfigMem.Inst_frame2_bit11.Q
rlabel metal2 4416 19530 4416 19530 0 Inst_E_TT_IF_ConfigMem.Inst_frame2_bit12.Q
rlabel metal3 14976 20580 14976 20580 0 Inst_E_TT_IF_ConfigMem.Inst_frame2_bit13.Q
rlabel metal2 14400 22008 14400 22008 0 Inst_E_TT_IF_ConfigMem.Inst_frame2_bit14.Q
rlabel metal2 14976 21084 14976 21084 0 Inst_E_TT_IF_ConfigMem.Inst_frame2_bit15.Q
rlabel metal2 19488 36456 19488 36456 0 Inst_E_TT_IF_ConfigMem.Inst_frame2_bit16.Q
rlabel metal3 19008 35196 19008 35196 0 Inst_E_TT_IF_ConfigMem.Inst_frame2_bit17.Q
rlabel metal2 19536 32844 19536 32844 0 Inst_E_TT_IF_ConfigMem.Inst_frame2_bit18.Q
rlabel metal2 9072 25116 9072 25116 0 Inst_E_TT_IF_ConfigMem.Inst_frame2_bit19.Q
rlabel metal2 17952 19950 17952 19950 0 Inst_E_TT_IF_ConfigMem.Inst_frame2_bit2.Q
rlabel metal2 10944 24295 10944 24295 0 Inst_E_TT_IF_ConfigMem.Inst_frame2_bit20.Q
rlabel metal3 11808 23268 11808 23268 0 Inst_E_TT_IF_ConfigMem.Inst_frame2_bit21.Q
rlabel metal3 9024 23100 9024 23100 0 Inst_E_TT_IF_ConfigMem.Inst_frame2_bit22.Q
rlabel via1 9600 22262 9600 22262 0 Inst_E_TT_IF_ConfigMem.Inst_frame2_bit23.Q
rlabel metal2 11712 22302 11712 22302 0 Inst_E_TT_IF_ConfigMem.Inst_frame2_bit24.Q
rlabel metal3 18720 23772 18720 23772 0 Inst_E_TT_IF_ConfigMem.Inst_frame2_bit25.Q
rlabel metal2 19296 23772 19296 23772 0 Inst_E_TT_IF_ConfigMem.Inst_frame2_bit26.Q
rlabel metal2 19968 22008 19968 22008 0 Inst_E_TT_IF_ConfigMem.Inst_frame2_bit27.Q
rlabel metal2 18432 29358 18432 29358 0 Inst_E_TT_IF_ConfigMem.Inst_frame2_bit28.Q
rlabel metal3 18480 29316 18480 29316 0 Inst_E_TT_IF_ConfigMem.Inst_frame2_bit29.Q
rlabel metal2 19584 19404 19584 19404 0 Inst_E_TT_IF_ConfigMem.Inst_frame2_bit3.Q
rlabel metal3 19584 27636 19584 27636 0 Inst_E_TT_IF_ConfigMem.Inst_frame2_bit30.Q
rlabel metal3 3552 26796 3552 26796 0 Inst_E_TT_IF_ConfigMem.Inst_frame2_bit31.Q
rlabel metal3 17760 31332 17760 31332 0 Inst_E_TT_IF_ConfigMem.Inst_frame2_bit4.Q
rlabel metal2 18432 30359 18432 30359 0 Inst_E_TT_IF_ConfigMem.Inst_frame2_bit5.Q
rlabel metal2 19200 29442 19200 29442 0 Inst_E_TT_IF_ConfigMem.Inst_frame2_bit6.Q
rlabel metal2 3504 28896 3504 28896 0 Inst_E_TT_IF_ConfigMem.Inst_frame2_bit7.Q
rlabel metal2 4896 29652 4896 29652 0 Inst_E_TT_IF_ConfigMem.Inst_frame2_bit8.Q
rlabel metal2 5472 28266 5472 28266 0 Inst_E_TT_IF_ConfigMem.Inst_frame2_bit9.Q
rlabel via1 6816 14025 6816 14025 0 Inst_E_TT_IF_ConfigMem.Inst_frame3_bit0.Q
rlabel metal2 8448 13692 8448 13692 0 Inst_E_TT_IF_ConfigMem.Inst_frame3_bit1.Q
rlabel metal2 11040 11839 11040 11839 0 Inst_E_TT_IF_ConfigMem.Inst_frame3_bit10.Q
rlabel metal2 9216 12558 9216 12558 0 Inst_E_TT_IF_ConfigMem.Inst_frame3_bit11.Q
rlabel metal2 18480 17787 18480 17787 0 Inst_E_TT_IF_ConfigMem.Inst_frame3_bit12.Q
rlabel metal2 16944 17220 16944 17220 0 Inst_E_TT_IF_ConfigMem.Inst_frame3_bit13.Q
rlabel metal2 17280 11970 17280 11970 0 Inst_E_TT_IF_ConfigMem.Inst_frame3_bit14.Q
rlabel metal2 15360 12222 15360 12222 0 Inst_E_TT_IF_ConfigMem.Inst_frame3_bit15.Q
rlabel metal2 4176 14196 4176 14196 0 Inst_E_TT_IF_ConfigMem.Inst_frame3_bit16.Q
rlabel metal2 2688 14994 2688 14994 0 Inst_E_TT_IF_ConfigMem.Inst_frame3_bit17.Q
rlabel metal2 1728 18144 1728 18144 0 Inst_E_TT_IF_ConfigMem.Inst_frame3_bit18.Q
rlabel metal2 2736 16800 2736 16800 0 Inst_E_TT_IF_ConfigMem.Inst_frame3_bit19.Q
rlabel metal2 7344 8904 7344 8904 0 Inst_E_TT_IF_ConfigMem.Inst_frame3_bit2.Q
rlabel metal2 3264 16296 3264 16296 0 Inst_E_TT_IF_ConfigMem.Inst_frame3_bit20.Q
rlabel via2 14688 23774 14688 23774 0 Inst_E_TT_IF_ConfigMem.Inst_frame3_bit21.Q
rlabel metal2 15264 23940 15264 23940 0 Inst_E_TT_IF_ConfigMem.Inst_frame3_bit22.Q
rlabel metal2 15360 23310 15360 23310 0 Inst_E_TT_IF_ConfigMem.Inst_frame3_bit23.Q
rlabel metal2 17952 38640 17952 38640 0 Inst_E_TT_IF_ConfigMem.Inst_frame3_bit24.Q
rlabel metal3 17136 38052 17136 38052 0 Inst_E_TT_IF_ConfigMem.Inst_frame3_bit25.Q
rlabel metal2 18528 36876 18528 36876 0 Inst_E_TT_IF_ConfigMem.Inst_frame3_bit26.Q
rlabel metal2 9600 27216 9600 27216 0 Inst_E_TT_IF_ConfigMem.Inst_frame3_bit27.Q
rlabel metal2 10464 26373 10464 26373 0 Inst_E_TT_IF_ConfigMem.Inst_frame3_bit28.Q
rlabel metal2 11616 25452 11616 25452 0 Inst_E_TT_IF_ConfigMem.Inst_frame3_bit29.Q
rlabel metal3 8016 8820 8016 8820 0 Inst_E_TT_IF_ConfigMem.Inst_frame3_bit3.Q
rlabel metal2 6432 23310 6432 23310 0 Inst_E_TT_IF_ConfigMem.Inst_frame3_bit30.Q
rlabel metal2 6816 24528 6816 24528 0 Inst_E_TT_IF_ConfigMem.Inst_frame3_bit31.Q
rlabel metal2 15840 14277 15840 14277 0 Inst_E_TT_IF_ConfigMem.Inst_frame3_bit4.Q
rlabel metal3 16896 13440 16896 13440 0 Inst_E_TT_IF_ConfigMem.Inst_frame3_bit5.Q
rlabel metal3 17328 9660 17328 9660 0 Inst_E_TT_IF_ConfigMem.Inst_frame3_bit6.Q
rlabel metal3 15168 8820 15168 8820 0 Inst_E_TT_IF_ConfigMem.Inst_frame3_bit7.Q
rlabel metal2 5520 12684 5520 12684 0 Inst_E_TT_IF_ConfigMem.Inst_frame3_bit8.Q
rlabel metal2 3840 13146 3840 13146 0 Inst_E_TT_IF_ConfigMem.Inst_frame3_bit9.Q
rlabel metal3 3744 7140 3744 7140 0 Inst_E_TT_IF_ConfigMem.Inst_frame4_bit0.Q
rlabel metal3 5760 5880 5760 5880 0 Inst_E_TT_IF_ConfigMem.Inst_frame4_bit1.Q
rlabel metal2 10608 9660 10608 9660 0 Inst_E_TT_IF_ConfigMem.Inst_frame4_bit10.Q
rlabel metal2 8928 10248 8928 10248 0 Inst_E_TT_IF_ConfigMem.Inst_frame4_bit11.Q
rlabel via2 17856 15537 17856 15537 0 Inst_E_TT_IF_ConfigMem.Inst_frame4_bit12.Q
rlabel metal3 16656 15540 16656 15540 0 Inst_E_TT_IF_ConfigMem.Inst_frame4_bit13.Q
rlabel metal2 15792 9660 15792 9660 0 Inst_E_TT_IF_ConfigMem.Inst_frame4_bit14.Q
rlabel metal2 14640 10080 14640 10080 0 Inst_E_TT_IF_ConfigMem.Inst_frame4_bit15.Q
rlabel metal2 4224 11977 4224 11977 0 Inst_E_TT_IF_ConfigMem.Inst_frame4_bit16.Q
rlabel metal2 2688 11424 2688 11424 0 Inst_E_TT_IF_ConfigMem.Inst_frame4_bit17.Q
rlabel metal2 13056 7644 13056 7644 0 Inst_E_TT_IF_ConfigMem.Inst_frame4_bit18.Q
rlabel metal2 11136 8022 11136 8022 0 Inst_E_TT_IF_ConfigMem.Inst_frame4_bit19.Q
rlabel metal2 11136 8904 11136 8904 0 Inst_E_TT_IF_ConfigMem.Inst_frame4_bit2.Q
rlabel metal2 17280 6678 17280 6678 0 Inst_E_TT_IF_ConfigMem.Inst_frame4_bit20.Q
rlabel metal2 15456 6510 15456 6510 0 Inst_E_TT_IF_ConfigMem.Inst_frame4_bit21.Q
rlabel metal2 16704 8701 16704 8701 0 Inst_E_TT_IF_ConfigMem.Inst_frame4_bit22.Q
rlabel metal2 15120 8148 15120 8148 0 Inst_E_TT_IF_ConfigMem.Inst_frame4_bit23.Q
rlabel metal2 2736 3612 2736 3612 0 Inst_E_TT_IF_ConfigMem.Inst_frame4_bit24.Q
rlabel metal2 4608 4074 4608 4074 0 Inst_E_TT_IF_ConfigMem.Inst_frame4_bit25.Q
rlabel metal2 6816 11634 6816 11634 0 Inst_E_TT_IF_ConfigMem.Inst_frame4_bit26.Q
rlabel metal3 8688 11172 8688 11172 0 Inst_E_TT_IF_ConfigMem.Inst_frame4_bit27.Q
rlabel metal2 13632 14448 13632 14448 0 Inst_E_TT_IF_ConfigMem.Inst_frame4_bit28.Q
rlabel metal2 15264 14448 15264 14448 0 Inst_E_TT_IF_ConfigMem.Inst_frame4_bit29.Q
rlabel metal3 12816 8820 12816 8820 0 Inst_E_TT_IF_ConfigMem.Inst_frame4_bit3.Q
rlabel metal2 13056 12936 13056 12936 0 Inst_E_TT_IF_ConfigMem.Inst_frame4_bit30.Q
rlabel metal2 14688 12936 14688 12936 0 Inst_E_TT_IF_ConfigMem.Inst_frame4_bit31.Q
rlabel metal3 18000 14196 18000 14196 0 Inst_E_TT_IF_ConfigMem.Inst_frame4_bit4.Q
rlabel metal2 19872 15001 19872 15001 0 Inst_E_TT_IF_ConfigMem.Inst_frame4_bit5.Q
rlabel metal3 19440 9660 19440 9660 0 Inst_E_TT_IF_ConfigMem.Inst_frame4_bit6.Q
rlabel metal2 20064 8904 20064 8904 0 Inst_E_TT_IF_ConfigMem.Inst_frame4_bit7.Q
rlabel metal3 3600 9492 3600 9492 0 Inst_E_TT_IF_ConfigMem.Inst_frame4_bit8.Q
rlabel metal2 5616 8148 5616 8148 0 Inst_E_TT_IF_ConfigMem.Inst_frame4_bit9.Q
rlabel metal2 2880 6717 2880 6717 0 Inst_E_TT_IF_ConfigMem.Inst_frame5_bit0.Q
rlabel metal2 2736 5880 2736 5880 0 Inst_E_TT_IF_ConfigMem.Inst_frame5_bit1.Q
rlabel metal2 11808 11172 11808 11172 0 Inst_E_TT_IF_ConfigMem.Inst_frame5_bit10.Q
rlabel metal2 12816 10227 12816 10227 0 Inst_E_TT_IF_ConfigMem.Inst_frame5_bit11.Q
rlabel metal2 20208 16464 20208 16464 0 Inst_E_TT_IF_ConfigMem.Inst_frame5_bit12.Q
rlabel metal2 18624 17175 18624 17175 0 Inst_E_TT_IF_ConfigMem.Inst_frame5_bit13.Q
rlabel metal2 18480 11172 18480 11172 0 Inst_E_TT_IF_ConfigMem.Inst_frame5_bit14.Q
rlabel metal2 20064 11172 20064 11172 0 Inst_E_TT_IF_ConfigMem.Inst_frame5_bit15.Q
rlabel metal2 3264 10122 3264 10122 0 Inst_E_TT_IF_ConfigMem.Inst_frame5_bit16.Q
rlabel metal2 4944 8820 4944 8820 0 Inst_E_TT_IF_ConfigMem.Inst_frame5_bit17.Q
rlabel metal3 9168 5880 9168 5880 0 Inst_E_TT_IF_ConfigMem.Inst_frame5_bit18.Q
rlabel metal2 8352 6132 8352 6132 0 Inst_E_TT_IF_ConfigMem.Inst_frame5_bit19.Q
rlabel metal2 8448 7189 8448 7189 0 Inst_E_TT_IF_ConfigMem.Inst_frame5_bit2.Q
rlabel metal2 17760 6174 17760 6174 0 Inst_E_TT_IF_ConfigMem.Inst_frame5_bit20.Q
rlabel metal3 19776 3612 19776 3612 0 Inst_E_TT_IF_ConfigMem.Inst_frame5_bit21.Q
rlabel metal2 18192 2100 18192 2100 0 Inst_E_TT_IF_ConfigMem.Inst_frame5_bit22.Q
rlabel metal3 19872 3360 19872 3360 0 Inst_E_TT_IF_ConfigMem.Inst_frame5_bit23.Q
rlabel metal2 3936 4998 3936 4998 0 Inst_E_TT_IF_ConfigMem.Inst_frame5_bit24.Q
rlabel metal2 5760 3654 5760 3654 0 Inst_E_TT_IF_ConfigMem.Inst_frame5_bit25.Q
rlabel metal2 11328 6174 11328 6174 0 Inst_E_TT_IF_ConfigMem.Inst_frame5_bit26.Q
rlabel metal2 13152 6132 13152 6132 0 Inst_E_TT_IF_ConfigMem.Inst_frame5_bit27.Q
rlabel metal2 18336 5166 18336 5166 0 Inst_E_TT_IF_ConfigMem.Inst_frame5_bit28.Q
rlabel metal3 19824 2856 19824 2856 0 Inst_E_TT_IF_ConfigMem.Inst_frame5_bit29.Q
rlabel metal2 9984 7434 9984 7434 0 Inst_E_TT_IF_ConfigMem.Inst_frame5_bit3.Q
rlabel metal2 17952 7434 17952 7434 0 Inst_E_TT_IF_ConfigMem.Inst_frame5_bit30.Q
rlabel metal2 20016 5040 20016 5040 0 Inst_E_TT_IF_ConfigMem.Inst_frame5_bit31.Q
rlabel metal2 20064 12684 20064 12684 0 Inst_E_TT_IF_ConfigMem.Inst_frame5_bit4.Q
rlabel metal2 18432 13146 18432 13146 0 Inst_E_TT_IF_ConfigMem.Inst_frame5_bit5.Q
rlabel metal2 16512 4165 16512 4165 0 Inst_E_TT_IF_ConfigMem.Inst_frame5_bit6.Q
rlabel metal2 14976 3864 14976 3864 0 Inst_E_TT_IF_ConfigMem.Inst_frame5_bit7.Q
rlabel metal2 4656 1260 4656 1260 0 Inst_E_TT_IF_ConfigMem.Inst_frame5_bit8.Q
rlabel metal2 2976 2100 2976 2100 0 Inst_E_TT_IF_ConfigMem.Inst_frame5_bit9.Q
rlabel metal2 9744 17220 9744 17220 0 Inst_E_TT_IF_ConfigMem.Inst_frame6_bit0.Q
rlabel metal2 11280 17787 11280 17787 0 Inst_E_TT_IF_ConfigMem.Inst_frame6_bit1.Q
rlabel metal2 18432 25795 18432 25795 0 Inst_E_TT_IF_ConfigMem.Inst_frame6_bit10.Q
rlabel metal2 19008 26544 19008 26544 0 Inst_E_TT_IF_ConfigMem.Inst_frame6_bit11.Q
rlabel metal2 15840 32802 15840 32802 0 Inst_E_TT_IF_ConfigMem.Inst_frame6_bit12.Q
rlabel metal2 17376 32804 17376 32804 0 Inst_E_TT_IF_ConfigMem.Inst_frame6_bit13.Q
rlabel metal2 17184 33726 17184 33726 0 Inst_E_TT_IF_ConfigMem.Inst_frame6_bit14.Q
rlabel metal2 12384 27636 12384 27636 0 Inst_E_TT_IF_ConfigMem.Inst_frame6_bit15.Q
rlabel metal3 12192 30072 12192 30072 0 Inst_E_TT_IF_ConfigMem.Inst_frame6_bit16.Q
rlabel metal2 11808 28350 11808 28350 0 Inst_E_TT_IF_ConfigMem.Inst_frame6_bit17.Q
rlabel metal2 7440 3612 7440 3612 0 Inst_E_TT_IF_ConfigMem.Inst_frame6_bit18.Q
rlabel metal2 9216 3864 9216 3864 0 Inst_E_TT_IF_ConfigMem.Inst_frame6_bit19.Q
rlabel metal2 11040 20118 11040 20118 0 Inst_E_TT_IF_ConfigMem.Inst_frame6_bit2.Q
rlabel via1 13344 4946 13344 4946 0 Inst_E_TT_IF_ConfigMem.Inst_frame6_bit20.Q
rlabel metal2 14688 4494 14688 4494 0 Inst_E_TT_IF_ConfigMem.Inst_frame6_bit21.Q
rlabel metal2 14880 1848 14880 1848 0 Inst_E_TT_IF_ConfigMem.Inst_frame6_bit22.Q
rlabel metal2 16896 1596 16896 1596 0 Inst_E_TT_IF_ConfigMem.Inst_frame6_bit23.Q
rlabel metal3 9984 4116 9984 4116 0 Inst_E_TT_IF_ConfigMem.Inst_frame6_bit24.Q
rlabel metal2 11712 4249 11712 4249 0 Inst_E_TT_IF_ConfigMem.Inst_frame6_bit25.Q
rlabel metal2 13344 3276 13344 3276 0 Inst_E_TT_IF_ConfigMem.Inst_frame6_bit26.Q
rlabel metal2 11328 3486 11328 3486 0 Inst_E_TT_IF_ConfigMem.Inst_frame6_bit27.Q
rlabel metal2 18432 3108 18432 3108 0 Inst_E_TT_IF_ConfigMem.Inst_frame6_bit28.Q
rlabel metal2 16800 2898 16800 2898 0 Inst_E_TT_IF_ConfigMem.Inst_frame6_bit29.Q
rlabel metal2 12576 19775 12576 19775 0 Inst_E_TT_IF_ConfigMem.Inst_frame6_bit3.Q
rlabel metal2 14112 7441 14112 7441 0 Inst_E_TT_IF_ConfigMem.Inst_frame6_bit30.Q
rlabel metal3 15168 6636 15168 6636 0 Inst_E_TT_IF_ConfigMem.Inst_frame6_bit31.Q
rlabel metal2 8784 16464 8784 16464 0 Inst_E_TT_IF_ConfigMem.Inst_frame6_bit4.Q
rlabel metal2 7200 17682 7200 17682 0 Inst_E_TT_IF_ConfigMem.Inst_frame6_bit5.Q
rlabel metal2 6528 21462 6528 21462 0 Inst_E_TT_IF_ConfigMem.Inst_frame6_bit6.Q
rlabel metal2 7344 20076 7344 20076 0 Inst_E_TT_IF_ConfigMem.Inst_frame6_bit7.Q
rlabel metal2 6816 22680 6816 22680 0 Inst_E_TT_IF_ConfigMem.Inst_frame6_bit8.Q
rlabel metal2 18912 25326 18912 25326 0 Inst_E_TT_IF_ConfigMem.Inst_frame6_bit9.Q
rlabel metal2 2304 31164 2304 31164 0 Inst_E_TT_IF_ConfigMem.Inst_frame7_bit0.Q
rlabel metal2 3840 31119 3840 31119 0 Inst_E_TT_IF_ConfigMem.Inst_frame7_bit1.Q
rlabel metal2 16608 37128 16608 37128 0 Inst_E_TT_IF_ConfigMem.Inst_frame7_bit10.Q
rlabel metal2 8832 29778 8832 29778 0 Inst_E_TT_IF_ConfigMem.Inst_frame7_bit11.Q
rlabel metal3 9216 29736 9216 29736 0 Inst_E_TT_IF_ConfigMem.Inst_frame7_bit12.Q
rlabel metal2 8352 29778 8352 29778 0 Inst_E_TT_IF_ConfigMem.Inst_frame7_bit13.Q
rlabel metal2 4896 17094 4896 17094 0 Inst_E_TT_IF_ConfigMem.Inst_frame7_bit14.Q
rlabel metal2 6432 17343 6432 17343 0 Inst_E_TT_IF_ConfigMem.Inst_frame7_bit15.Q
rlabel metal2 14016 29200 14016 29200 0 Inst_E_TT_IF_ConfigMem.Inst_frame7_bit16.Q
rlabel metal3 15840 28560 15840 28560 0 Inst_E_TT_IF_ConfigMem.Inst_frame7_bit17.Q
rlabel metal2 11328 35994 11328 35994 0 Inst_E_TT_IF_ConfigMem.Inst_frame7_bit18.Q
rlabel metal2 13344 35616 13344 35616 0 Inst_E_TT_IF_ConfigMem.Inst_frame7_bit19.Q
rlabel metal3 3792 21588 3792 21588 0 Inst_E_TT_IF_ConfigMem.Inst_frame7_bit2.Q
rlabel metal2 6048 31626 6048 31626 0 Inst_E_TT_IF_ConfigMem.Inst_frame7_bit20.Q
rlabel via1 7584 31334 7584 31334 0 Inst_E_TT_IF_ConfigMem.Inst_frame7_bit21.Q
rlabel metal2 2688 25956 2688 25956 0 Inst_E_TT_IF_ConfigMem.Inst_frame7_bit22.Q
rlabel metal2 3840 25333 3840 25333 0 Inst_E_TT_IF_ConfigMem.Inst_frame7_bit23.Q
rlabel metal2 11040 21630 11040 21630 0 Inst_E_TT_IF_ConfigMem.Inst_frame7_bit24.Q
rlabel metal2 12720 21000 12720 21000 0 Inst_E_TT_IF_ConfigMem.Inst_frame7_bit25.Q
rlabel metal2 12288 31080 12288 31080 0 Inst_E_TT_IF_ConfigMem.Inst_frame7_bit26.Q
rlabel metal2 10464 31080 10464 31080 0 Inst_E_TT_IF_ConfigMem.Inst_frame7_bit27.Q
rlabel metal2 9936 31395 9936 31395 0 Inst_E_TT_IF_ConfigMem.Inst_frame7_bit28.Q
rlabel metal2 8352 32004 8352 32004 0 Inst_E_TT_IF_ConfigMem.Inst_frame7_bit29.Q
rlabel metal3 3696 23604 3696 23604 0 Inst_E_TT_IF_ConfigMem.Inst_frame7_bit3.Q
rlabel metal2 9888 18984 9888 18984 0 Inst_E_TT_IF_ConfigMem.Inst_frame7_bit30.Q
rlabel via1 8256 19235 8256 19235 0 Inst_E_TT_IF_ConfigMem.Inst_frame7_bit31.Q
rlabel metal2 2640 21000 2640 21000 0 Inst_E_TT_IF_ConfigMem.Inst_frame7_bit4.Q
rlabel metal2 14496 28014 14496 28014 0 Inst_E_TT_IF_ConfigMem.Inst_frame7_bit5.Q
rlabel metal2 15648 26082 15648 26082 0 Inst_E_TT_IF_ConfigMem.Inst_frame7_bit6.Q
rlabel metal2 14736 26124 14736 26124 0 Inst_E_TT_IF_ConfigMem.Inst_frame7_bit7.Q
rlabel metal2 15264 35364 15264 35364 0 Inst_E_TT_IF_ConfigMem.Inst_frame7_bit8.Q
rlabel metal2 16992 34895 16992 34895 0 Inst_E_TT_IF_ConfigMem.Inst_frame7_bit9.Q
rlabel metal2 2688 23310 2688 23310 0 Inst_E_TT_IF_ConfigMem.Inst_frame8_bit10.Q
rlabel metal2 4560 23268 4560 23268 0 Inst_E_TT_IF_ConfigMem.Inst_frame8_bit11.Q
rlabel metal2 13824 29904 13824 29904 0 Inst_E_TT_IF_ConfigMem.Inst_frame8_bit12.Q
rlabel metal2 15360 29869 15360 29869 0 Inst_E_TT_IF_ConfigMem.Inst_frame8_bit13.Q
rlabel metal2 11040 36414 11040 36414 0 Inst_E_TT_IF_ConfigMem.Inst_frame8_bit14.Q
rlabel via1 12816 36703 12816 36703 0 Inst_E_TT_IF_ConfigMem.Inst_frame8_bit15.Q
rlabel metal2 4800 30912 4800 30912 0 Inst_E_TT_IF_ConfigMem.Inst_frame8_bit16.Q
rlabel metal2 6336 30909 6336 30909 0 Inst_E_TT_IF_ConfigMem.Inst_frame8_bit17.Q
rlabel metal2 3360 27846 3360 27846 0 Inst_E_TT_IF_ConfigMem.Inst_frame8_bit18.Q
rlabel metal2 2976 28987 2976 28987 0 Inst_E_TT_IF_ConfigMem.Inst_frame8_bit19.Q
rlabel metal2 2016 36540 2016 36540 0 Inst_E_TT_IF_ConfigMem.Inst_frame8_bit20.Q
rlabel metal2 3456 36841 3456 36841 0 Inst_E_TT_IF_ConfigMem.Inst_frame8_bit21.Q
rlabel via1 2160 32848 2160 32848 0 Inst_E_TT_IF_ConfigMem.Inst_frame8_bit22.Q
rlabel metal3 3264 32844 3264 32844 0 Inst_E_TT_IF_ConfigMem.Inst_frame8_bit23.Q
rlabel via1 3984 34360 3984 34360 0 Inst_E_TT_IF_ConfigMem.Inst_frame8_bit24.Q
rlabel metal2 2400 34818 2400 34818 0 Inst_E_TT_IF_ConfigMem.Inst_frame8_bit25.Q
rlabel metal2 2304 38640 2304 38640 0 Inst_E_TT_IF_ConfigMem.Inst_frame8_bit26.Q
rlabel metal3 5808 37632 5808 37632 0 Inst_E_TT_IF_ConfigMem.Inst_frame8_bit27.Q
rlabel via1 3600 39727 3600 39727 0 Inst_E_TT_IF_ConfigMem.Inst_frame8_bit28.Q
rlabel metal2 2016 39774 2016 39774 0 Inst_E_TT_IF_ConfigMem.Inst_frame8_bit29.Q
rlabel metal2 13344 33348 13344 33348 0 Inst_E_TT_IF_ConfigMem.Inst_frame8_bit30.Q
rlabel metal2 11712 33726 11712 33726 0 Inst_E_TT_IF_ConfigMem.Inst_frame8_bit31.Q
rlabel metal2 1536 31458 1536 31458 0 Inst_E_TT_IF_switch_matrix.N1BEG0
rlabel metal2 2304 32676 2304 32676 0 Inst_E_TT_IF_switch_matrix.N1BEG1
rlabel metal2 1536 34902 1536 34902 0 Inst_E_TT_IF_switch_matrix.N1BEG2
rlabel metal2 1440 35700 1440 35700 0 Inst_E_TT_IF_switch_matrix.N1BEG3
rlabel metal4 8208 32676 8208 32676 0 Inst_E_TT_IF_switch_matrix.N2BEG0
rlabel metal2 4032 35196 4032 35196 0 Inst_E_TT_IF_switch_matrix.N2BEG1
rlabel metal2 1392 37464 1392 37464 0 Inst_E_TT_IF_switch_matrix.N2BEG2
rlabel metal2 1824 37296 1824 37296 0 Inst_E_TT_IF_switch_matrix.N2BEG3
rlabel metal2 4080 37296 4080 37296 0 Inst_E_TT_IF_switch_matrix.N2BEG4
rlabel metal2 3408 38136 3408 38136 0 Inst_E_TT_IF_switch_matrix.N2BEG5
rlabel metal2 13440 33957 13440 33957 0 Inst_E_TT_IF_switch_matrix.N2BEG6
rlabel metal3 1680 38976 1680 38976 0 Inst_E_TT_IF_switch_matrix.N2BEG7
rlabel metal2 5808 35196 5808 35196 0 Inst_E_TT_IF_switch_matrix.N4BEG0
rlabel metal3 14640 34776 14640 34776 0 Inst_E_TT_IF_switch_matrix.N4BEG1
rlabel metal2 16944 41160 16944 41160 0 Inst_E_TT_IF_switch_matrix.N4BEG2
rlabel metal3 7680 30240 7680 30240 0 Inst_E_TT_IF_switch_matrix.N4BEG3
rlabel metal3 6960 3444 6960 3444 0 Inst_E_TT_IF_switch_matrix.S1BEG0
rlabel metal3 15600 29232 15600 29232 0 Inst_E_TT_IF_switch_matrix.S1BEG1
rlabel metal4 13056 18438 13056 18438 0 Inst_E_TT_IF_switch_matrix.S1BEG2
rlabel metal2 8592 14280 8592 14280 0 Inst_E_TT_IF_switch_matrix.S1BEG3
rlabel metal4 2400 4158 2400 4158 0 Inst_E_TT_IF_switch_matrix.S2BEG0
rlabel metal3 12720 21672 12720 21672 0 Inst_E_TT_IF_switch_matrix.S2BEG1
rlabel metal4 12192 16884 12192 16884 0 Inst_E_TT_IF_switch_matrix.S2BEG2
rlabel metal3 10032 20076 10032 20076 0 Inst_E_TT_IF_switch_matrix.S2BEG3
rlabel metal3 10416 1596 10416 1596 0 Inst_E_TT_IF_switch_matrix.S2BEG4
rlabel metal4 11424 10164 11424 10164 0 Inst_E_TT_IF_switch_matrix.S2BEG5
rlabel metal3 12336 20076 12336 20076 0 Inst_E_TT_IF_switch_matrix.S2BEG6
rlabel metal3 9120 10164 9120 10164 0 Inst_E_TT_IF_switch_matrix.S2BEG7
rlabel metal3 14928 1176 14928 1176 0 Inst_E_TT_IF_switch_matrix.S4BEG0
rlabel metal2 18432 1848 18432 1848 0 Inst_E_TT_IF_switch_matrix.S4BEG1
rlabel metal3 17328 1176 17328 1176 0 Inst_E_TT_IF_switch_matrix.S4BEG2
rlabel metal3 13536 1680 13536 1680 0 Inst_E_TT_IF_switch_matrix.S4BEG3
rlabel metal3 6000 1680 6000 1680 0 Inst_E_TT_IF_switch_matrix.W1BEG0
rlabel metal2 14400 3570 14400 3570 0 Inst_E_TT_IF_switch_matrix.W1BEG1
rlabel metal3 5136 1764 5136 1764 0 Inst_E_TT_IF_switch_matrix.W1BEG2
rlabel metal2 11904 4116 11904 4116 0 Inst_E_TT_IF_switch_matrix.W1BEG3
rlabel metal2 2496 1638 2496 1638 0 Inst_E_TT_IF_switch_matrix.W2BEG0
rlabel metal2 1728 1092 1728 1092 0 Inst_E_TT_IF_switch_matrix.W2BEG1
rlabel metal2 1440 4032 1440 4032 0 Inst_E_TT_IF_switch_matrix.W2BEG2
rlabel metal2 1776 2688 1776 2688 0 Inst_E_TT_IF_switch_matrix.W2BEG3
rlabel metal2 2016 4032 2016 4032 0 Inst_E_TT_IF_switch_matrix.W2BEG4
rlabel metal2 1680 3360 1680 3360 0 Inst_E_TT_IF_switch_matrix.W2BEG5
rlabel metal2 2496 3486 2496 3486 0 Inst_E_TT_IF_switch_matrix.W2BEG6
rlabel metal3 3648 2688 3648 2688 0 Inst_E_TT_IF_switch_matrix.W2BEG7
rlabel metal2 2208 5334 2208 5334 0 Inst_E_TT_IF_switch_matrix.W2BEGb0
rlabel metal2 18528 14868 18528 14868 0 Inst_E_TT_IF_switch_matrix.W2BEGb1
rlabel metal2 20256 6258 20256 6258 0 Inst_E_TT_IF_switch_matrix.W2BEGb2
rlabel metal2 2496 6336 2496 6336 0 Inst_E_TT_IF_switch_matrix.W2BEGb3
rlabel metal2 1920 5586 1920 5586 0 Inst_E_TT_IF_switch_matrix.W2BEGb4
rlabel metal2 19776 6930 19776 6930 0 Inst_E_TT_IF_switch_matrix.W2BEGb5
rlabel metal3 18768 4200 18768 4200 0 Inst_E_TT_IF_switch_matrix.W2BEGb6
rlabel metal2 5664 4998 5664 4998 0 Inst_E_TT_IF_switch_matrix.W2BEGb7
rlabel metal2 8544 11676 8544 11676 0 Inst_E_TT_IF_switch_matrix.W6BEG0
rlabel metal2 2016 13860 2016 13860 0 Inst_E_TT_IF_switch_matrix.W6BEG1
rlabel metal2 1632 13566 1632 13566 0 Inst_E_TT_IF_switch_matrix.W6BEG10
rlabel metal2 4416 14700 4416 14700 0 Inst_E_TT_IF_switch_matrix.W6BEG11
rlabel metal2 1728 12348 1728 12348 0 Inst_E_TT_IF_switch_matrix.W6BEG2
rlabel metal2 8544 13272 8544 13272 0 Inst_E_TT_IF_switch_matrix.W6BEG3
rlabel metal2 2112 10752 2112 10752 0 Inst_E_TT_IF_switch_matrix.W6BEG4
rlabel metal3 2112 13902 2112 13902 0 Inst_E_TT_IF_switch_matrix.W6BEG5
rlabel metal3 17376 13314 17376 13314 0 Inst_E_TT_IF_switch_matrix.W6BEG6
rlabel metal2 1728 13986 1728 13986 0 Inst_E_TT_IF_switch_matrix.W6BEG7
rlabel metal2 2496 13314 2496 13314 0 Inst_E_TT_IF_switch_matrix.W6BEG8
rlabel metal2 18240 17262 18240 17262 0 Inst_E_TT_IF_switch_matrix.W6BEG9
rlabel metal3 1728 6300 1728 6300 0 Inst_E_TT_IF_switch_matrix.WW4BEG0
rlabel metal2 20141 6340 20141 6340 0 Inst_E_TT_IF_switch_matrix.WW4BEG1
rlabel metal2 1728 10332 1728 10332 0 Inst_E_TT_IF_switch_matrix.WW4BEG10
rlabel metal2 3120 11424 3120 11424 0 Inst_E_TT_IF_switch_matrix.WW4BEG11
rlabel metal3 12864 7980 12864 7980 0 Inst_E_TT_IF_switch_matrix.WW4BEG12
rlabel metal2 2112 6510 2112 6510 0 Inst_E_TT_IF_switch_matrix.WW4BEG13
rlabel metal2 2112 8652 2112 8652 0 Inst_E_TT_IF_switch_matrix.WW4BEG14
rlabel metal2 1536 4410 1536 4410 0 Inst_E_TT_IF_switch_matrix.WW4BEG15
rlabel metal2 2016 7308 2016 7308 0 Inst_E_TT_IF_switch_matrix.WW4BEG2
rlabel metal3 4128 7182 4128 7182 0 Inst_E_TT_IF_switch_matrix.WW4BEG3
rlabel metal2 2016 8316 2016 8316 0 Inst_E_TT_IF_switch_matrix.WW4BEG4
rlabel metal2 19968 14532 19968 14532 0 Inst_E_TT_IF_switch_matrix.WW4BEG5
rlabel metal2 1632 9366 1632 9366 0 Inst_E_TT_IF_switch_matrix.WW4BEG6
rlabel metal2 2880 9156 2880 9156 0 Inst_E_TT_IF_switch_matrix.WW4BEG7
rlabel metal2 2496 9324 2496 9324 0 Inst_E_TT_IF_switch_matrix.WW4BEG8
rlabel metal3 17856 13440 17856 13440 0 Inst_E_TT_IF_switch_matrix.WW4BEG9
rlabel metal2 1488 37884 1488 37884 0 N1BEG[0]
rlabel metal2 1968 39900 1968 39900 0 N1BEG[1]
rlabel metal2 1776 38220 1776 38220 0 N1BEG[2]
rlabel metal3 2352 38556 2352 38556 0 N1BEG[3]
rlabel metal2 1824 1248 1824 1248 0 N1END[0]
rlabel metal2 2016 1290 2016 1290 0 N1END[1]
rlabel metal2 2208 702 2208 702 0 N1END[2]
rlabel metal2 2400 366 2400 366 0 N1END[3]
rlabel metal2 10368 41622 10368 41622 0 N2BEG[0]
rlabel metal3 3456 35028 3456 35028 0 N2BEG[1]
rlabel metal2 1632 37674 1632 37674 0 N2BEG[2]
rlabel metal3 2400 37632 2400 37632 0 N2BEG[3]
rlabel metal2 3120 38388 3120 38388 0 N2BEG[4]
rlabel metal2 3552 38976 3552 38976 0 N2BEG[5]
rlabel metal2 12864 39102 12864 39102 0 N2BEG[6]
rlabel metal3 2028 39060 2028 39060 0 N2BEG[7]
rlabel metal2 6816 38976 6816 38976 0 N2BEGb[0]
rlabel metal2 1680 39900 1680 39900 0 N2BEGb[1]
rlabel metal2 1776 40656 1776 40656 0 N2BEGb[2]
rlabel metal2 7056 37632 7056 37632 0 N2BEGb[3]
rlabel metal2 9600 41118 9600 41118 0 N2BEGb[4]
rlabel metal2 2112 41370 2112 41370 0 N2BEGb[5]
rlabel metal2 4128 38388 4128 38388 0 N2BEGb[6]
rlabel metal2 5376 39942 5376 39942 0 N2BEGb[7]
rlabel metal2 4128 450 4128 450 0 N2END[0]
rlabel metal4 1152 18480 1152 18480 0 N2END[1]
rlabel metal2 4512 492 4512 492 0 N2END[2]
rlabel metal2 4704 240 4704 240 0 N2END[3]
rlabel metal4 1248 18396 1248 18396 0 N2END[4]
rlabel metal2 5088 324 5088 324 0 N2END[5]
rlabel metal2 5280 156 5280 156 0 N2END[6]
rlabel metal2 5472 366 5472 366 0 N2END[7]
rlabel metal3 4752 2184 4752 2184 0 N2MID[0]
rlabel metal2 1536 39606 1536 39606 0 N2MID[1]
rlabel metal2 1344 41034 1344 41034 0 N2MID[2]
rlabel metal4 2160 15120 2160 15120 0 N2MID[3]
rlabel metal4 1056 17220 1056 17220 0 N2MID[4]
rlabel metal3 2064 40320 2064 40320 0 N2MID[5]
rlabel metal2 17568 22974 17568 22974 0 N2MID[6]
rlabel metal4 2304 17388 2304 17388 0 N2MID[7]
rlabel metal2 3072 41538 3072 41538 0 N4BEG[0]
rlabel metal2 7584 42306 7584 42306 0 N4BEG[10]
rlabel metal2 7776 42348 7776 42348 0 N4BEG[11]
rlabel metal2 5856 40908 5856 40908 0 N4BEG[12]
rlabel metal3 12582 41412 12582 41412 0 N4BEG[13]
rlabel metal2 8352 42012 8352 42012 0 N4BEG[14]
rlabel metal2 6144 41454 6144 41454 0 N4BEG[15]
rlabel metal2 5328 38724 5328 38724 0 N4BEG[1]
rlabel metal2 3456 41412 3456 41412 0 N4BEG[2]
rlabel metal2 5760 41706 5760 41706 0 N4BEG[3]
rlabel metal2 6240 40320 6240 40320 0 N4BEG[4]
rlabel metal3 6000 40656 6000 40656 0 N4BEG[5]
rlabel metal2 6624 39858 6624 39858 0 N4BEG[6]
rlabel metal2 9984 41664 9984 41664 0 N4BEG[7]
rlabel metal3 7584 40656 7584 40656 0 N4BEG[8]
rlabel metal4 7536 35280 7536 35280 0 N4BEG[9]
rlabel metal2 6864 11508 6864 11508 0 N4END[0]
rlabel metal3 7248 13776 7248 13776 0 N4END[10]
rlabel metal2 7776 366 7776 366 0 N4END[11]
rlabel metal2 7968 618 7968 618 0 N4END[12]
rlabel metal2 8160 744 8160 744 0 N4END[13]
rlabel metal2 8352 324 8352 324 0 N4END[14]
rlabel metal2 8544 534 8544 534 0 N4END[15]
rlabel metal2 13728 13440 13728 13440 0 N4END[1]
rlabel metal2 13200 13188 13200 13188 0 N4END[2]
rlabel metal3 6432 14028 6432 14028 0 N4END[3]
rlabel metal2 6432 660 6432 660 0 N4END[4]
rlabel metal2 6624 492 6624 492 0 N4END[5]
rlabel metal2 6816 408 6816 408 0 N4END[6]
rlabel metal2 7008 660 7008 660 0 N4END[7]
rlabel metal2 7200 660 7200 660 0 N4END[8]
rlabel metal2 7392 618 7392 618 0 N4END[9]
rlabel metal3 13488 24192 13488 24192 0 RST_N_TT_PROJECT
rlabel metal2 8736 492 8736 492 0 S1BEG[0]
rlabel metal2 15264 1974 15264 1974 0 S1BEG[1]
rlabel metal2 12864 756 12864 756 0 S1BEG[2]
rlabel metal3 8976 2436 8976 2436 0 S1BEG[3]
rlabel metal2 6528 17472 6528 17472 0 S1END[0]
rlabel metal2 12720 17724 12720 17724 0 S1END[1]
rlabel metal2 12576 38514 12576 38514 0 S1END[2]
rlabel metal3 7872 15540 7872 15540 0 S1END[3]
rlabel metal2 9504 282 9504 282 0 S2BEG[0]
rlabel metal2 12480 672 12480 672 0 S2BEG[1]
rlabel metal2 9888 870 9888 870 0 S2BEG[2]
rlabel metal2 9984 1722 9984 1722 0 S2BEG[3]
rlabel metal2 10272 492 10272 492 0 S2BEG[4]
rlabel metal2 10944 1638 10944 1638 0 S2BEG[5]
rlabel metal2 12096 1512 12096 1512 0 S2BEG[6]
rlabel metal2 9600 2352 9600 2352 0 S2BEG[7]
rlabel metal2 10368 1386 10368 1386 0 S2BEGb[0]
rlabel metal2 11232 492 11232 492 0 S2BEGb[1]
rlabel metal2 11424 366 11424 366 0 S2BEGb[2]
rlabel metal2 11616 282 11616 282 0 S2BEGb[3]
rlabel metal2 11808 660 11808 660 0 S2BEGb[4]
rlabel metal2 12000 492 12000 492 0 S2BEGb[5]
rlabel metal2 12192 450 12192 450 0 S2BEGb[6]
rlabel metal2 12384 576 12384 576 0 S2BEGb[7]
rlabel metal2 11040 41634 11040 41634 0 S2END[0]
rlabel metal2 10944 37128 10944 37128 0 S2END[1]
rlabel metal2 11424 42516 11424 42516 0 S2END[2]
rlabel metal2 11616 42306 11616 42306 0 S2END[3]
rlabel metal2 6144 37464 6144 37464 0 S2END[4]
rlabel metal2 12000 42432 12000 42432 0 S2END[5]
rlabel metal2 12192 41508 12192 41508 0 S2END[6]
rlabel metal2 12384 42768 12384 42768 0 S2END[7]
rlabel metal3 9456 2352 9456 2352 0 S2MID[0]
rlabel metal2 10512 1176 10512 1176 0 S2MID[1]
rlabel metal2 8880 37380 8880 37380 0 S2MID[2]
rlabel metal3 10896 37296 10896 37296 0 S2MID[3]
rlabel metal3 10416 36624 10416 36624 0 S2MID[4]
rlabel metal2 10464 42264 10464 42264 0 S2MID[5]
rlabel metal3 11280 1848 11280 1848 0 S2MID[6]
rlabel metal4 11616 20034 11616 20034 0 S2MID[7]
rlabel metal2 12576 492 12576 492 0 S4BEG[0]
rlabel metal2 14496 156 14496 156 0 S4BEG[10]
rlabel metal2 14688 450 14688 450 0 S4BEG[11]
rlabel metal2 14880 492 14880 492 0 S4BEG[12]
rlabel metal2 18240 630 18240 630 0 S4BEG[13]
rlabel metal2 15264 282 15264 282 0 S4BEG[14]
rlabel metal2 15456 366 15456 366 0 S4BEG[15]
rlabel metal2 12768 282 12768 282 0 S4BEG[1]
rlabel metal2 12960 1248 12960 1248 0 S4BEG[2]
rlabel metal2 13152 240 13152 240 0 S4BEG[3]
rlabel metal2 13344 1122 13344 1122 0 S4BEG[4]
rlabel metal2 13536 492 13536 492 0 S4BEG[5]
rlabel metal2 13728 702 13728 702 0 S4BEG[6]
rlabel metal2 13920 660 13920 660 0 S4BEG[7]
rlabel metal2 14112 366 14112 366 0 S4BEG[8]
rlabel metal2 14304 198 14304 198 0 S4BEG[9]
rlabel metal2 12576 42264 12576 42264 0 S4END[0]
rlabel metal2 14496 42264 14496 42264 0 S4END[10]
rlabel metal2 14688 42264 14688 42264 0 S4END[11]
rlabel metal2 14880 42054 14880 42054 0 S4END[12]
rlabel metal2 15072 42054 15072 42054 0 S4END[13]
rlabel metal2 15264 41718 15264 41718 0 S4END[14]
rlabel metal2 15456 42054 15456 42054 0 S4END[15]
rlabel metal2 14688 16128 14688 16128 0 S4END[1]
rlabel metal2 13488 18816 13488 18816 0 S4END[2]
rlabel metal2 13152 42810 13152 42810 0 S4END[3]
rlabel metal2 13344 42264 13344 42264 0 S4END[4]
rlabel metal2 13536 42306 13536 42306 0 S4END[5]
rlabel metal2 13728 42264 13728 42264 0 S4END[6]
rlabel metal2 14640 2268 14640 2268 0 S4END[7]
rlabel metal3 14064 2688 14064 2688 0 S4END[8]
rlabel metal3 14592 1848 14592 1848 0 S4END[9]
rlabel metal3 20994 18900 20994 18900 0 UIO_IN_TT_PROJECT0
rlabel metal3 21090 19404 21090 19404 0 UIO_IN_TT_PROJECT1
rlabel metal3 21378 19908 21378 19908 0 UIO_IN_TT_PROJECT2
rlabel metal2 12192 22428 12192 22428 0 UIO_IN_TT_PROJECT3
rlabel metal2 12384 21672 12384 21672 0 UIO_IN_TT_PROJECT4
rlabel metal2 19872 21924 19872 21924 0 UIO_IN_TT_PROJECT5
rlabel metal3 21138 21924 21138 21924 0 UIO_IN_TT_PROJECT6
rlabel metal4 16416 23772 16416 23772 0 UIO_IN_TT_PROJECT7
rlabel metal3 20802 10836 20802 10836 0 UIO_OE_TT_PROJECT0
rlabel metal3 20544 11382 20544 11382 0 UIO_OE_TT_PROJECT1
rlabel metal2 18912 11802 18912 11802 0 UIO_OE_TT_PROJECT2
rlabel metal3 21234 12348 21234 12348 0 UIO_OE_TT_PROJECT3
rlabel metal3 20994 12852 20994 12852 0 UIO_OE_TT_PROJECT4
rlabel metal2 20736 11886 20736 11886 0 UIO_OE_TT_PROJECT5
rlabel metal4 20736 11970 20736 11970 0 UIO_OE_TT_PROJECT6
rlabel metal3 20994 14364 20994 14364 0 UIO_OE_TT_PROJECT7
rlabel metal3 20994 6804 20994 6804 0 UIO_OUT_TT_PROJECT0
rlabel metal2 20064 16716 20064 16716 0 UIO_OUT_TT_PROJECT1
rlabel metal3 21464 8064 21464 8064 0 UIO_OUT_TT_PROJECT2
rlabel metal3 20994 8316 20994 8316 0 UIO_OUT_TT_PROJECT3
rlabel metal3 20802 8820 20802 8820 0 UIO_OUT_TT_PROJECT4
rlabel metal2 19008 13314 19008 13314 0 UIO_OUT_TT_PROJECT5
rlabel metal3 20544 9786 20544 9786 0 UIO_OUT_TT_PROJECT6
rlabel metal3 4224 12516 4224 12516 0 UIO_OUT_TT_PROJECT7
rlabel metal2 4128 15624 4128 15624 0 UI_IN_TT_PROJECT0
rlabel metal3 18834 15372 18834 15372 0 UI_IN_TT_PROJECT1
rlabel metal3 21282 15876 21282 15876 0 UI_IN_TT_PROJECT2
rlabel metal3 21090 16380 21090 16380 0 UI_IN_TT_PROJECT3
rlabel metal3 21186 16884 21186 16884 0 UI_IN_TT_PROJECT4
rlabel metal3 21042 17388 21042 17388 0 UI_IN_TT_PROJECT5
rlabel metal3 20658 17892 20658 17892 0 UI_IN_TT_PROJECT6
rlabel metal3 21330 18396 21330 18396 0 UI_IN_TT_PROJECT7
rlabel metal2 11424 3276 11424 3276 0 UO_OUT_TT_PROJECT0
rlabel metal2 16128 7056 16128 7056 0 UO_OUT_TT_PROJECT1
rlabel metal3 20544 3822 20544 3822 0 UO_OUT_TT_PROJECT2
rlabel metal3 20994 4284 20994 4284 0 UO_OUT_TT_PROJECT3
rlabel via2 21426 4788 21426 4788 0 UO_OUT_TT_PROJECT4
rlabel metal3 21426 5292 21426 5292 0 UO_OUT_TT_PROJECT5
rlabel metal2 19680 10416 19680 10416 0 UO_OUT_TT_PROJECT6
rlabel metal3 21426 6300 21426 6300 0 UO_OUT_TT_PROJECT7
rlabel metal2 15648 366 15648 366 0 UserCLK
rlabel metal2 15696 41412 15696 41412 0 UserCLKo
rlabel metal3 1290 84 1290 84 0 W1BEG[0]
rlabel metal3 2142 420 2142 420 0 W1BEG[1]
rlabel metal3 1710 756 1710 756 0 W1BEG[2]
rlabel metal3 222 1092 222 1092 0 W1BEG[3]
rlabel metal2 2304 1344 2304 1344 0 W2BEG[0]
rlabel metal2 1536 1512 1536 1512 0 W2BEG[1]
rlabel metal2 1920 1680 1920 1680 0 W2BEG[2]
rlabel metal3 798 2436 798 2436 0 W2BEG[3]
rlabel metal3 990 2772 990 2772 0 W2BEG[4]
rlabel metal3 798 3108 798 3108 0 W2BEG[5]
rlabel metal3 1182 3444 1182 3444 0 W2BEG[6]
rlabel metal2 2256 2856 2256 2856 0 W2BEG[7]
rlabel metal2 1920 3864 1920 3864 0 W2BEGb[0]
rlabel metal2 17760 4410 17760 4410 0 W2BEGb[1]
rlabel metal3 1278 4788 1278 4788 0 W2BEGb[2]
rlabel metal3 1182 5124 1182 5124 0 W2BEGb[3]
rlabel metal2 1728 5124 1728 5124 0 W2BEGb[4]
rlabel metal2 8832 6384 8832 6384 0 W2BEGb[5]
rlabel metal2 17376 5250 17376 5250 0 W2BEGb[6]
rlabel metal3 78 6468 78 6468 0 W2BEGb[7]
rlabel metal2 1536 12054 1536 12054 0 W6BEG[0]
rlabel metal3 798 15540 798 15540 0 W6BEG[10]
rlabel metal3 990 15876 990 15876 0 W6BEG[11]
rlabel metal3 894 12516 894 12516 0 W6BEG[1]
rlabel metal2 1536 12600 1536 12600 0 W6BEG[2]
rlabel metal2 1920 12726 1920 12726 0 W6BEG[3]
rlabel metal2 1872 11928 1872 11928 0 W6BEG[4]
rlabel metal3 990 13860 990 13860 0 W6BEG[5]
rlabel metal2 1344 13818 1344 13818 0 W6BEG[6]
rlabel metal2 1536 14364 1536 14364 0 W6BEG[7]
rlabel metal2 2304 14532 2304 14532 0 W6BEG[8]
rlabel metal2 17952 15498 17952 15498 0 W6BEG[9]
rlabel metal2 1536 6720 1536 6720 0 WW4BEG[0]
rlabel metal2 1488 9660 1488 9660 0 WW4BEG[10]
rlabel metal2 2880 10626 2880 10626 0 WW4BEG[11]
rlabel metal2 1392 8148 1392 8148 0 WW4BEG[12]
rlabel metal2 1920 7182 1920 7182 0 WW4BEG[13]
rlabel metal2 1872 8820 1872 8820 0 WW4BEG[14]
rlabel metal2 1344 4872 1344 4872 0 WW4BEG[15]
rlabel metal3 1086 7140 1086 7140 0 WW4BEG[1]
rlabel metal2 1824 7434 1824 7434 0 WW4BEG[2]
rlabel metal2 1392 7392 1392 7392 0 WW4BEG[3]
rlabel metal3 942 8148 942 8148 0 WW4BEG[4]
rlabel metal3 318 8484 318 8484 0 WW4BEG[5]
rlabel metal3 798 8820 798 8820 0 WW4BEG[6]
rlabel metal2 2688 8988 2688 8988 0 WW4BEG[7]
rlabel metal2 2304 9156 2304 9156 0 WW4BEG[8]
rlabel metal2 14208 9576 14208 9576 0 WW4BEG[9]
rlabel metal2 8160 34902 8160 34902 0 _000_
rlabel metal3 9168 32844 9168 32844 0 _001_
rlabel metal3 7056 32844 7056 32844 0 _002_
rlabel metal3 12384 39144 12384 39144 0 _003_
rlabel metal2 14784 31626 14784 31626 0 _004_
rlabel metal3 6192 14700 6192 14700 0 _005_
rlabel metal2 13920 25221 13920 25221 0 _006_
rlabel metal3 4608 19320 4608 19320 0 _007_
rlabel metal2 3600 17976 3600 17976 0 _008_
rlabel metal2 11952 26880 11952 26880 0 _009_
rlabel metal3 12768 30408 12768 30408 0 _010_
rlabel metal2 7680 21042 7680 21042 0 _011_
rlabel metal2 7872 20496 7872 20496 0 _012_
rlabel metal2 9168 29820 9168 29820 0 _013_
rlabel metal2 8544 29400 8544 29400 0 _014_
rlabel metal2 14112 25326 14112 25326 0 _015_
rlabel metal3 16080 26292 16080 26292 0 _016_
rlabel metal2 14208 27342 14208 27342 0 _017_
rlabel metal2 3072 22008 3072 22008 0 _018_
rlabel metal3 4032 20748 4032 20748 0 _019_
rlabel metal2 9984 33138 9984 33138 0 _020_
rlabel metal2 10080 33390 10080 33390 0 _021_
rlabel metal2 9840 32844 9840 32844 0 _022_
rlabel metal3 9312 33012 9312 33012 0 _023_
rlabel metal2 8256 35112 8256 35112 0 _024_
rlabel metal3 7296 34356 7296 34356 0 _025_
rlabel metal2 6336 35028 6336 35028 0 _026_
rlabel metal2 6048 34482 6048 34482 0 _027_
rlabel metal2 9888 35238 9888 35238 0 _028_
rlabel metal2 10368 35070 10368 35070 0 _029_
rlabel metal3 11382 35112 11382 35112 0 _030_
rlabel metal2 8880 34860 8880 34860 0 _031_
rlabel metal2 9120 36582 9120 36582 0 _032_
rlabel metal2 9120 34608 9120 34608 0 _033_
rlabel metal2 9360 33096 9360 33096 0 _034_
rlabel metal2 7968 37170 7968 37170 0 _035_
rlabel metal2 9696 33558 9696 33558 0 _036_
rlabel metal2 7872 35364 7872 35364 0 _037_
rlabel metal2 10176 34316 10176 34316 0 _038_
rlabel metal2 12288 10332 12288 10332 0 _039_
rlabel via2 11712 28138 11712 28138 0 _040_
rlabel metal3 12432 17892 12432 17892 0 _041_
rlabel metal2 5184 26208 5184 26208 0 _042_
rlabel metal3 5856 25956 5856 25956 0 _043_
rlabel metal3 6432 26796 6432 26796 0 _044_
rlabel metal3 6432 26208 6432 26208 0 _045_
rlabel metal2 6048 26208 6048 26208 0 _046_
rlabel metal3 15168 19824 15168 19824 0 _047_
rlabel metal2 18096 13272 18096 13272 0 _048_
rlabel metal2 17904 27468 17904 27468 0 _049_
rlabel metal2 18336 30072 18336 30072 0 _050_
rlabel metal3 18576 27804 18576 27804 0 _051_
rlabel metal3 19536 27720 19536 27720 0 _052_
rlabel metal2 19488 27888 19488 27888 0 _053_
rlabel metal2 14112 13314 14112 13314 0 _054_
rlabel metal2 17952 17934 17952 17934 0 _055_
rlabel metal2 18912 22302 18912 22302 0 _056_
rlabel metal2 19680 23856 19680 23856 0 _057_
rlabel metal2 18336 22764 18336 22764 0 _058_
rlabel metal3 19584 23730 19584 23730 0 _059_
rlabel metal2 19584 22932 19584 22932 0 _060_
rlabel metal2 4512 7266 4512 7266 0 _061_
rlabel metal3 10080 12516 10080 12516 0 _062_
rlabel metal2 6528 20160 6528 20160 0 _063_
rlabel metal2 7632 23100 7632 23100 0 _064_
rlabel metal2 9504 21126 9504 21126 0 _065_
rlabel metal2 9648 20748 9648 20748 0 _066_
rlabel metal2 12000 21168 12000 21168 0 _067_
rlabel metal3 10560 22344 10560 22344 0 _068_
rlabel metal2 11520 16170 11520 16170 0 _069_
rlabel metal2 11808 8316 11808 8316 0 _070_
rlabel metal2 11136 24864 11136 24864 0 _071_
rlabel metal2 9888 25368 9888 25368 0 _072_
rlabel metal2 11040 24664 11040 24664 0 _073_
rlabel metal3 11568 24612 11568 24612 0 _074_
rlabel metal2 11760 24696 11760 24696 0 _075_
rlabel metal2 16896 13902 16896 13902 0 _076_
rlabel metal2 18912 13356 18912 13356 0 _077_
rlabel metal2 19776 33054 19776 33054 0 _078_
rlabel metal3 20064 35364 20064 35364 0 _079_
rlabel metal2 18000 34356 18000 34356 0 _080_
rlabel metal2 20064 35238 20064 35238 0 _081_
rlabel metal2 19872 33012 19872 33012 0 _082_
rlabel metal3 14448 13188 14448 13188 0 _083_
rlabel metal2 16320 14532 16320 14532 0 _084_
rlabel metal2 14928 20328 14928 20328 0 _085_
rlabel metal3 15504 20160 15504 20160 0 _086_
rlabel metal2 16032 22176 16032 22176 0 _087_
rlabel metal2 15648 21756 15648 21756 0 _088_
rlabel metal3 15264 21588 15264 21588 0 _089_
rlabel metal2 11808 9912 11808 9912 0 _090_
rlabel metal2 4992 21378 4992 21378 0 _091_
rlabel metal2 7392 14070 7392 14070 0 _092_
rlabel metal2 5952 20788 5952 20788 0 _093_
rlabel metal3 4416 18312 4416 18312 0 _094_
rlabel metal2 4608 20832 4608 20832 0 _095_
rlabel metal2 4704 19278 4704 19278 0 _096_
rlabel metal3 5136 18732 5136 18732 0 _097_
rlabel metal3 4752 20076 4752 20076 0 _098_
rlabel metal2 8928 15750 8928 15750 0 _099_
rlabel metal2 5712 27636 5712 27636 0 _100_
rlabel metal3 6240 29148 6240 29148 0 _101_
rlabel metal2 5760 29904 5760 29904 0 _102_
rlabel metal2 6336 29400 6336 29400 0 _103_
rlabel metal3 6192 29064 6192 29064 0 _104_
rlabel metal2 17376 17766 17376 17766 0 _105_
rlabel metal3 19056 29148 19056 29148 0 _106_
rlabel metal3 18960 31332 18960 31332 0 _107_
rlabel metal2 16512 31080 16512 31080 0 _108_
rlabel metal2 19296 31416 19296 31416 0 _109_
rlabel metal2 19584 29526 19584 29526 0 _110_
rlabel metal2 19104 18732 19104 18732 0 _111_
rlabel metal2 18672 18564 18672 18564 0 _112_
rlabel metal3 19344 18732 19344 18732 0 _113_
rlabel metal3 19968 20580 19968 20580 0 _114_
rlabel metal2 20016 19236 20016 19236 0 _115_
rlabel metal2 19200 19824 19200 19824 0 _116_
rlabel metal3 5280 13188 5280 13188 0 _117_
rlabel metal2 5472 23856 5472 23856 0 _118_
rlabel metal2 8064 23730 8064 23730 0 _119_
rlabel metal3 7584 23772 7584 23772 0 _120_
rlabel metal2 8256 23898 8256 23898 0 _121_
rlabel metal2 7920 24612 7920 24612 0 _122_
rlabel metal2 11904 14994 11904 14994 0 _123_
rlabel metal2 11904 25368 11904 25368 0 _124_
rlabel metal2 11136 26712 11136 26712 0 _125_
rlabel metal2 9408 27588 9408 27588 0 _126_
rlabel metal2 11424 27090 11424 27090 0 _127_
rlabel metal2 12000 25620 12000 25620 0 _128_
rlabel metal2 17472 16128 17472 16128 0 _129_
rlabel metal2 18912 38262 18912 38262 0 _130_
rlabel metal3 18480 38892 18480 38892 0 _131_
rlabel metal2 16320 39396 16320 39396 0 _132_
rlabel metal2 18912 38934 18912 38934 0 _133_
rlabel metal2 19056 38304 19056 38304 0 _134_
rlabel metal2 15744 19047 15744 19047 0 _135_
rlabel metal2 14352 24780 14352 24780 0 _136_
rlabel metal2 14880 25242 14880 25242 0 _137_
rlabel metal2 15072 24360 15072 24360 0 _138_
rlabel metal2 15648 24906 15648 24906 0 _139_
rlabel metal2 15552 24150 15552 24150 0 _140_
rlabel metal2 3312 18060 3312 18060 0 _141_
rlabel metal2 3360 15582 3360 15582 0 _142_
rlabel metal2 3168 18396 3168 18396 0 _143_
rlabel metal2 3264 15792 3264 15792 0 _144_
rlabel metal2 3552 15708 3552 15708 0 _145_
rlabel metal2 3504 16212 3504 16212 0 _146_
rlabel metal2 12288 27804 12288 27804 0 _147_
rlabel metal2 12576 28392 12576 28392 0 _148_
rlabel metal2 13152 28602 13152 28602 0 _149_
rlabel metal2 12672 28224 12672 28224 0 _150_
rlabel metal2 10272 29400 10272 29400 0 _151_
rlabel metal2 10224 28644 10224 28644 0 _152_
rlabel metal2 17472 33222 17472 33222 0 _153_
rlabel metal2 17664 32592 17664 32592 0 _154_
rlabel metal2 18912 26628 18912 26628 0 _155_
rlabel metal2 19104 26250 19104 26250 0 _156_
rlabel metal2 19296 26208 19296 26208 0 _157_
rlabel metal2 18672 24612 18672 24612 0 _158_
rlabel metal2 18816 24864 18816 24864 0 _159_
rlabel metal2 19488 24528 19488 24528 0 _160_
rlabel metal2 19392 24990 19392 24990 0 _161_
rlabel metal3 6192 20076 6192 20076 0 _162_
rlabel metal2 7008 20496 7008 20496 0 _163_
rlabel metal2 7584 20958 7584 20958 0 _164_
rlabel metal2 7872 21294 7872 21294 0 _165_
rlabel metal2 6144 21084 6144 21084 0 _166_
rlabel metal2 6816 21252 6816 21252 0 _167_
rlabel metal2 7584 20328 7584 20328 0 _168_
rlabel metal2 7248 19908 7248 19908 0 _169_
rlabel metal3 8784 28224 8784 28224 0 _170_
rlabel metal2 8928 29190 8928 29190 0 _171_
rlabel via1 9026 29148 9026 29148 0 _172_
rlabel metal2 8784 30828 8784 30828 0 _173_
rlabel metal2 9312 29400 9312 29400 0 _174_
rlabel metal2 8160 29232 8160 29232 0 _175_
rlabel metal2 19920 36876 19920 36876 0 _176_
rlabel metal2 17184 35784 17184 35784 0 _177_
rlabel metal3 15456 24528 15456 24528 0 _178_
rlabel metal2 16128 27300 16128 27300 0 _179_
rlabel metal2 15360 26754 15360 26754 0 _180_
rlabel metal3 15936 26796 15936 26796 0 _181_
rlabel metal2 15744 26901 15744 26901 0 _182_
rlabel metal2 14256 25536 14256 25536 0 _183_
rlabel metal3 14880 26292 14880 26292 0 _184_
rlabel metal2 15264 25578 15264 25578 0 _185_
rlabel metal2 15600 26544 15600 26544 0 _186_
rlabel metal2 4560 21756 4560 21756 0 _187_
rlabel metal2 4320 22008 4320 22008 0 _188_
rlabel metal2 3552 20790 3552 20790 0 _189_
rlabel metal2 3744 20832 3744 20832 0 _190_
rlabel metal2 3312 24612 3312 24612 0 _191_
rlabel metal2 3360 20748 3360 20748 0 _192_
rlabel metal2 4224 21462 4224 21462 0 _193_
rlabel metal2 4032 21798 4032 21798 0 _194_
rlabel metal3 17856 23268 17856 23268 0 _195_
rlabel metal2 17424 23268 17424 23268 0 _196_
rlabel metal3 5136 32844 5136 32844 0 _197_
rlabel metal2 6432 32676 6432 32676 0 _198_
rlabel via1 7104 31336 7104 31336 0 _199_
rlabel metal2 11904 40152 11904 40152 0 _200_
rlabel metal3 12576 39900 12576 39900 0 _201_
rlabel metal2 12240 36708 12240 36708 0 _202_
rlabel metal2 14352 30492 14352 30492 0 _203_
rlabel metal2 15456 31332 15456 31332 0 _204_
rlabel metal2 14880 30492 14880 30492 0 _205_
rlabel metal2 5568 14784 5568 14784 0 _206_
rlabel metal3 6048 16044 6048 16044 0 _207_
rlabel metal2 5856 17052 5856 17052 0 _208_
rlabel metal2 19104 32214 19104 32214 0 clknet_0_UserCLK
rlabel metal2 19824 26376 19824 26376 0 clknet_1_0__leaf_UserCLK
rlabel metal3 17616 37632 17616 37632 0 clknet_1_1__leaf_UserCLK
<< properties >>
string FIXED_BBOX 0 0 21504 43008
<< end >>
