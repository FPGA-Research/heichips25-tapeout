magic
tech ihp-sg13g2
magscale 1 2
timestamp 1752747676
<< metal1 >>
rect 1152 9848 41856 9872
rect 1152 9808 4928 9848
rect 4968 9808 5010 9848
rect 5050 9808 5092 9848
rect 5132 9808 5174 9848
rect 5214 9808 5256 9848
rect 5296 9808 20048 9848
rect 20088 9808 20130 9848
rect 20170 9808 20212 9848
rect 20252 9808 20294 9848
rect 20334 9808 20376 9848
rect 20416 9808 35168 9848
rect 35208 9808 35250 9848
rect 35290 9808 35332 9848
rect 35372 9808 35414 9848
rect 35454 9808 35496 9848
rect 35536 9808 41856 9848
rect 1152 9784 41856 9808
rect 4099 9680 4157 9681
rect 4099 9640 4108 9680
rect 4148 9640 4157 9680
rect 4099 9639 4157 9640
rect 4579 9680 4637 9681
rect 4579 9640 4588 9680
rect 4628 9640 4637 9680
rect 4579 9639 4637 9640
rect 9195 9680 9237 9689
rect 9195 9640 9196 9680
rect 9236 9640 9237 9680
rect 9195 9631 9237 9640
rect 11691 9680 11733 9689
rect 11691 9640 11692 9680
rect 11732 9640 11733 9680
rect 11691 9631 11733 9640
rect 13323 9680 13365 9689
rect 13323 9640 13324 9680
rect 13364 9640 13365 9680
rect 13323 9631 13365 9640
rect 16683 9680 16725 9689
rect 16683 9640 16684 9680
rect 16724 9640 16725 9680
rect 16683 9631 16725 9640
rect 19467 9680 19509 9689
rect 19467 9640 19468 9680
rect 19508 9640 19509 9680
rect 19467 9631 19509 9640
rect 21387 9680 21429 9689
rect 21387 9640 21388 9680
rect 21428 9640 21429 9680
rect 21387 9631 21429 9640
rect 32043 9680 32085 9689
rect 32043 9640 32044 9680
rect 32084 9640 32085 9680
rect 32043 9631 32085 9640
rect 32427 9680 32469 9689
rect 32427 9640 32428 9680
rect 32468 9640 32469 9680
rect 32427 9631 32469 9640
rect 32811 9680 32853 9689
rect 32811 9640 32812 9680
rect 32852 9640 32853 9680
rect 32811 9631 32853 9640
rect 37707 9680 37749 9689
rect 37707 9640 37708 9680
rect 37748 9640 37749 9680
rect 37707 9631 37749 9640
rect 40683 9680 40725 9689
rect 40683 9640 40684 9680
rect 40724 9640 40725 9680
rect 40683 9631 40725 9640
rect 41451 9680 41493 9689
rect 41451 9640 41452 9680
rect 41492 9640 41493 9680
rect 41451 9631 41493 9640
rect 2955 9596 2997 9605
rect 2955 9556 2956 9596
rect 2996 9556 2997 9596
rect 2955 9547 2997 9556
rect 1507 9512 1565 9513
rect 1507 9472 1516 9512
rect 1556 9472 1565 9512
rect 1507 9471 1565 9472
rect 2755 9512 2813 9513
rect 2755 9472 2764 9512
rect 2804 9472 2813 9512
rect 2755 9471 2813 9472
rect 3339 9512 3381 9521
rect 3339 9472 3340 9512
rect 3380 9472 3381 9512
rect 3339 9463 3381 9472
rect 3435 9512 3477 9521
rect 3435 9472 3436 9512
rect 3476 9472 3477 9512
rect 3435 9463 3477 9472
rect 3531 9512 3573 9521
rect 3531 9472 3532 9512
rect 3572 9472 3573 9512
rect 3531 9463 3573 9472
rect 3627 9512 3669 9521
rect 3627 9472 3628 9512
rect 3668 9472 3669 9512
rect 3627 9463 3669 9472
rect 3819 9512 3861 9521
rect 3819 9472 3820 9512
rect 3860 9472 3861 9512
rect 3819 9463 3861 9472
rect 3915 9512 3957 9521
rect 3915 9472 3916 9512
rect 3956 9472 3957 9512
rect 3915 9463 3957 9472
rect 4299 9512 4341 9521
rect 4299 9472 4300 9512
rect 4340 9472 4341 9512
rect 4299 9463 4341 9472
rect 4395 9512 4437 9521
rect 4395 9472 4396 9512
rect 4436 9472 4437 9512
rect 4395 9463 4437 9472
rect 4491 9512 4533 9521
rect 4491 9472 4492 9512
rect 4532 9472 4533 9512
rect 4491 9463 4533 9472
rect 7747 9512 7805 9513
rect 7747 9472 7756 9512
rect 7796 9472 7805 9512
rect 7747 9471 7805 9472
rect 8995 9512 9053 9513
rect 8995 9472 9004 9512
rect 9044 9472 9053 9512
rect 8995 9471 9053 9472
rect 10243 9512 10301 9513
rect 10243 9472 10252 9512
rect 10292 9472 10301 9512
rect 10243 9471 10301 9472
rect 11491 9512 11549 9513
rect 11491 9472 11500 9512
rect 11540 9472 11549 9512
rect 11491 9471 11549 9472
rect 11875 9512 11933 9513
rect 11875 9472 11884 9512
rect 11924 9472 11933 9512
rect 11875 9471 11933 9472
rect 13123 9512 13181 9513
rect 13123 9472 13132 9512
rect 13172 9472 13181 9512
rect 13123 9471 13181 9472
rect 15235 9512 15293 9513
rect 15235 9472 15244 9512
rect 15284 9472 15293 9512
rect 15235 9471 15293 9472
rect 16483 9512 16541 9513
rect 16483 9472 16492 9512
rect 16532 9472 16541 9512
rect 16483 9471 16541 9472
rect 17827 9512 17885 9513
rect 17827 9472 17836 9512
rect 17876 9472 17885 9512
rect 17827 9471 17885 9472
rect 19075 9512 19133 9513
rect 19075 9472 19084 9512
rect 19124 9472 19133 9512
rect 19075 9471 19133 9472
rect 22435 9512 22493 9513
rect 22435 9472 22444 9512
rect 22484 9472 22493 9512
rect 22435 9471 22493 9472
rect 23683 9512 23741 9513
rect 23683 9472 23692 9512
rect 23732 9472 23741 9512
rect 23683 9471 23741 9472
rect 24259 9512 24317 9513
rect 24259 9472 24268 9512
rect 24308 9472 24317 9512
rect 24259 9471 24317 9472
rect 25507 9512 25565 9513
rect 25507 9472 25516 9512
rect 25556 9472 25565 9512
rect 25507 9471 25565 9472
rect 27715 9512 27773 9513
rect 27715 9472 27724 9512
rect 27764 9472 27773 9512
rect 27715 9471 27773 9472
rect 28963 9512 29021 9513
rect 28963 9472 28972 9512
rect 29012 9472 29021 9512
rect 28963 9471 29021 9472
rect 29539 9512 29597 9513
rect 29539 9472 29548 9512
rect 29588 9472 29597 9512
rect 29539 9471 29597 9472
rect 30499 9512 30557 9513
rect 30499 9472 30508 9512
rect 30548 9472 30557 9512
rect 30499 9471 30557 9472
rect 30787 9512 30845 9513
rect 30787 9472 30796 9512
rect 30836 9472 30845 9512
rect 30787 9471 30845 9472
rect 31659 9512 31701 9521
rect 31659 9472 31660 9512
rect 31700 9472 31701 9512
rect 31659 9463 31701 9472
rect 34531 9512 34589 9513
rect 34531 9472 34540 9512
rect 34580 9472 34589 9512
rect 34531 9471 34589 9472
rect 35203 9512 35261 9513
rect 35203 9472 35212 9512
rect 35252 9472 35261 9512
rect 35203 9471 35261 9472
rect 36163 9512 36221 9513
rect 36163 9472 36172 9512
rect 36212 9472 36221 9512
rect 36163 9471 36221 9472
rect 36547 9512 36605 9513
rect 36547 9472 36556 9512
rect 36596 9472 36605 9512
rect 36547 9471 36605 9472
rect 19651 9428 19709 9429
rect 19651 9388 19660 9428
rect 19700 9388 19709 9428
rect 19651 9387 19709 9388
rect 21187 9428 21245 9429
rect 21187 9388 21196 9428
rect 21236 9388 21245 9428
rect 21187 9387 21245 9388
rect 32227 9428 32285 9429
rect 32227 9388 32236 9428
rect 32276 9388 32285 9428
rect 32227 9387 32285 9388
rect 32611 9428 32669 9429
rect 32611 9388 32620 9428
rect 32660 9388 32669 9428
rect 32611 9387 32669 9388
rect 32995 9428 33053 9429
rect 32995 9388 33004 9428
rect 33044 9388 33053 9428
rect 32995 9387 33053 9388
rect 37891 9428 37949 9429
rect 37891 9388 37900 9428
rect 37940 9388 37949 9428
rect 37891 9387 37949 9388
rect 40483 9428 40541 9429
rect 40483 9388 40492 9428
rect 40532 9388 40541 9428
rect 40483 9387 40541 9388
rect 40867 9428 40925 9429
rect 40867 9388 40876 9428
rect 40916 9388 40925 9428
rect 40867 9387 40925 9388
rect 41251 9428 41309 9429
rect 41251 9388 41260 9428
rect 41300 9388 41309 9428
rect 41251 9387 41309 9388
rect 33387 9344 33429 9353
rect 33387 9304 33388 9344
rect 33428 9304 33429 9344
rect 33387 9295 33429 9304
rect 34827 9344 34869 9353
rect 34827 9304 34828 9344
rect 34868 9304 34869 9344
rect 34827 9295 34869 9304
rect 36843 9344 36885 9353
rect 36843 9304 36844 9344
rect 36884 9304 36885 9344
rect 36843 9295 36885 9304
rect 41067 9344 41109 9353
rect 41067 9304 41068 9344
rect 41108 9304 41109 9344
rect 41067 9295 41109 9304
rect 19275 9260 19317 9269
rect 19275 9220 19276 9260
rect 19316 9220 19317 9260
rect 19275 9211 19317 9220
rect 23883 9260 23925 9269
rect 23883 9220 23884 9260
rect 23924 9220 23925 9260
rect 23883 9211 23925 9220
rect 25707 9260 25749 9269
rect 25707 9220 25708 9260
rect 25748 9220 25749 9260
rect 25707 9211 25749 9220
rect 29163 9260 29205 9269
rect 29163 9220 29164 9260
rect 29204 9220 29205 9260
rect 29163 9211 29205 9220
rect 34251 9260 34293 9269
rect 34251 9220 34252 9260
rect 34292 9220 34293 9260
rect 34251 9211 34293 9220
rect 35883 9260 35925 9269
rect 35883 9220 35884 9260
rect 35924 9220 35925 9260
rect 35883 9211 35925 9220
rect 1152 9092 41856 9116
rect 1152 9052 3688 9092
rect 3728 9052 3770 9092
rect 3810 9052 3852 9092
rect 3892 9052 3934 9092
rect 3974 9052 4016 9092
rect 4056 9052 18808 9092
rect 18848 9052 18890 9092
rect 18930 9052 18972 9092
rect 19012 9052 19054 9092
rect 19094 9052 19136 9092
rect 19176 9052 33928 9092
rect 33968 9052 34010 9092
rect 34050 9052 34092 9092
rect 34132 9052 34174 9092
rect 34214 9052 34256 9092
rect 34296 9052 41856 9092
rect 1152 9028 41856 9052
rect 3627 8924 3669 8933
rect 3627 8884 3628 8924
rect 3668 8884 3669 8924
rect 3627 8875 3669 8884
rect 9483 8840 9525 8849
rect 9483 8800 9484 8840
rect 9524 8800 9525 8840
rect 9483 8791 9525 8800
rect 13899 8840 13941 8849
rect 13899 8800 13900 8840
rect 13940 8800 13941 8840
rect 13899 8791 13941 8800
rect 15531 8840 15573 8849
rect 15531 8800 15532 8840
rect 15572 8800 15573 8840
rect 15531 8791 15573 8800
rect 20043 8840 20085 8849
rect 20043 8800 20044 8840
rect 20084 8800 20085 8840
rect 20043 8791 20085 8800
rect 29259 8840 29301 8849
rect 29259 8800 29260 8840
rect 29300 8800 29301 8840
rect 29259 8791 29301 8800
rect 29739 8840 29781 8849
rect 29739 8800 29740 8840
rect 29780 8800 29781 8840
rect 29739 8791 29781 8800
rect 31755 8840 31797 8849
rect 31755 8800 31756 8840
rect 31796 8800 31797 8840
rect 31755 8791 31797 8800
rect 32139 8840 32181 8849
rect 32139 8800 32140 8840
rect 32180 8800 32181 8840
rect 32139 8791 32181 8800
rect 32523 8840 32565 8849
rect 32523 8800 32524 8840
rect 32564 8800 32565 8840
rect 32523 8791 32565 8800
rect 32907 8840 32949 8849
rect 32907 8800 32908 8840
rect 32948 8800 32949 8840
rect 32907 8791 32949 8800
rect 36171 8840 36213 8849
rect 36171 8800 36172 8840
rect 36212 8800 36213 8840
rect 36171 8791 36213 8800
rect 36555 8840 36597 8849
rect 36555 8800 36556 8840
rect 36596 8800 36597 8840
rect 36555 8791 36597 8800
rect 38763 8840 38805 8849
rect 38763 8800 38764 8840
rect 38804 8800 38805 8840
rect 38763 8791 38805 8800
rect 39147 8840 39189 8849
rect 39147 8800 39148 8840
rect 39188 8800 39189 8840
rect 39147 8791 39189 8800
rect 40011 8840 40053 8849
rect 40011 8800 40012 8840
rect 40052 8800 40053 8840
rect 40011 8791 40053 8800
rect 40395 8840 40437 8849
rect 40395 8800 40396 8840
rect 40436 8800 40437 8840
rect 40395 8791 40437 8800
rect 41067 8840 41109 8849
rect 41067 8800 41068 8840
rect 41108 8800 41109 8840
rect 41067 8791 41109 8800
rect 41451 8840 41493 8849
rect 41451 8800 41452 8840
rect 41492 8800 41493 8840
rect 41451 8791 41493 8800
rect 19843 8756 19901 8757
rect 19227 8714 19269 8723
rect 19843 8716 19852 8756
rect 19892 8716 19901 8756
rect 19843 8715 19901 8716
rect 22443 8756 22485 8765
rect 22443 8716 22444 8756
rect 22484 8716 22485 8756
rect 1603 8672 1661 8673
rect 1603 8632 1612 8672
rect 1652 8632 1661 8672
rect 1603 8631 1661 8632
rect 2851 8672 2909 8673
rect 2851 8632 2860 8672
rect 2900 8632 2909 8672
rect 2851 8631 2909 8632
rect 3523 8672 3581 8673
rect 3523 8632 3532 8672
rect 3572 8632 3581 8672
rect 3523 8631 3581 8632
rect 3627 8672 3669 8681
rect 3627 8632 3628 8672
rect 3668 8632 3669 8672
rect 3627 8623 3669 8632
rect 3811 8672 3869 8673
rect 3811 8632 3820 8672
rect 3860 8632 3869 8672
rect 3811 8631 3869 8632
rect 4011 8672 4053 8681
rect 4011 8632 4012 8672
rect 4052 8632 4053 8672
rect 4011 8623 4053 8632
rect 4107 8672 4149 8681
rect 4107 8632 4108 8672
rect 4148 8632 4149 8672
rect 4107 8623 4149 8632
rect 4203 8672 4245 8681
rect 4203 8632 4204 8672
rect 4244 8632 4245 8672
rect 4203 8623 4245 8632
rect 4299 8672 4341 8681
rect 4299 8632 4300 8672
rect 4340 8632 4341 8672
rect 4299 8623 4341 8632
rect 4771 8672 4829 8673
rect 4771 8632 4780 8672
rect 4820 8632 4829 8672
rect 4771 8631 4829 8632
rect 6019 8672 6077 8673
rect 6019 8632 6028 8672
rect 6068 8632 6077 8672
rect 6019 8631 6077 8632
rect 6403 8672 6461 8673
rect 6403 8632 6412 8672
rect 6452 8632 6461 8672
rect 6403 8631 6461 8632
rect 7651 8672 7709 8673
rect 7651 8632 7660 8672
rect 7700 8632 7709 8672
rect 7651 8631 7709 8632
rect 8035 8672 8093 8673
rect 8035 8632 8044 8672
rect 8084 8632 8093 8672
rect 8035 8631 8093 8632
rect 9283 8672 9341 8673
rect 9283 8632 9292 8672
rect 9332 8632 9341 8672
rect 9283 8631 9341 8632
rect 9667 8672 9725 8673
rect 9667 8632 9676 8672
rect 9716 8632 9725 8672
rect 9667 8631 9725 8632
rect 10915 8672 10973 8673
rect 10915 8632 10924 8672
rect 10964 8632 10973 8672
rect 10915 8631 10973 8632
rect 12451 8672 12509 8673
rect 12451 8632 12460 8672
rect 12500 8632 12509 8672
rect 12451 8631 12509 8632
rect 13699 8672 13757 8673
rect 13699 8632 13708 8672
rect 13748 8632 13757 8672
rect 13699 8631 13757 8632
rect 14083 8672 14141 8673
rect 14083 8632 14092 8672
rect 14132 8632 14141 8672
rect 14083 8631 14141 8632
rect 15331 8672 15389 8673
rect 15331 8632 15340 8672
rect 15380 8632 15389 8672
rect 15331 8631 15389 8632
rect 15907 8672 15965 8673
rect 15907 8632 15916 8672
rect 15956 8632 15965 8672
rect 15907 8631 15965 8632
rect 17155 8672 17213 8673
rect 17155 8632 17164 8672
rect 17204 8632 17213 8672
rect 17155 8631 17213 8632
rect 17643 8672 17685 8681
rect 17643 8632 17644 8672
rect 17684 8632 17685 8672
rect 17643 8623 17685 8632
rect 17739 8672 17781 8681
rect 17739 8632 17740 8672
rect 17780 8632 17781 8672
rect 17739 8623 17781 8632
rect 18123 8672 18165 8681
rect 18123 8632 18124 8672
rect 18164 8632 18165 8672
rect 18123 8623 18165 8632
rect 18219 8672 18261 8681
rect 19227 8674 19228 8714
rect 19268 8674 19269 8714
rect 22443 8707 22485 8716
rect 29443 8756 29501 8757
rect 29443 8716 29452 8756
rect 29492 8716 29501 8756
rect 29443 8715 29501 8716
rect 29923 8756 29981 8757
rect 29923 8716 29932 8756
rect 29972 8716 29981 8756
rect 29923 8715 29981 8716
rect 31939 8756 31997 8757
rect 31939 8716 31948 8756
rect 31988 8716 31997 8756
rect 31939 8715 31997 8716
rect 32323 8756 32381 8757
rect 32323 8716 32332 8756
rect 32372 8716 32381 8756
rect 32323 8715 32381 8716
rect 32707 8756 32765 8757
rect 32707 8716 32716 8756
rect 32756 8716 32765 8756
rect 32707 8715 32765 8716
rect 33091 8756 33149 8757
rect 33091 8716 33100 8756
rect 33140 8716 33149 8756
rect 33091 8715 33149 8716
rect 36355 8756 36413 8757
rect 36355 8716 36364 8756
rect 36404 8716 36413 8756
rect 36355 8715 36413 8716
rect 36739 8756 36797 8757
rect 36739 8716 36748 8756
rect 36788 8716 36797 8756
rect 36739 8715 36797 8716
rect 38563 8756 38621 8757
rect 38563 8716 38572 8756
rect 38612 8716 38621 8756
rect 38563 8715 38621 8716
rect 38947 8756 39005 8757
rect 38947 8716 38956 8756
rect 38996 8716 39005 8756
rect 38947 8715 39005 8716
rect 39811 8756 39869 8757
rect 39811 8716 39820 8756
rect 39860 8716 39869 8756
rect 39811 8715 39869 8716
rect 40195 8756 40253 8757
rect 40195 8716 40204 8756
rect 40244 8716 40253 8756
rect 40195 8715 40253 8716
rect 40867 8756 40925 8757
rect 40867 8716 40876 8756
rect 40916 8716 40925 8756
rect 40867 8715 40925 8716
rect 41251 8756 41309 8757
rect 41251 8716 41260 8756
rect 41300 8716 41309 8756
rect 41251 8715 41309 8716
rect 23547 8681 23589 8690
rect 27003 8681 27045 8690
rect 18219 8632 18220 8672
rect 18260 8632 18261 8672
rect 18219 8623 18261 8632
rect 18691 8672 18749 8673
rect 18691 8632 18700 8672
rect 18740 8632 18749 8672
rect 19227 8665 19269 8674
rect 20227 8672 20285 8673
rect 18691 8631 18749 8632
rect 20227 8632 20236 8672
rect 20276 8632 20285 8672
rect 20227 8631 20285 8632
rect 21475 8672 21533 8673
rect 21475 8632 21484 8672
rect 21524 8632 21533 8672
rect 21475 8631 21533 8632
rect 21963 8672 22005 8681
rect 21963 8632 21964 8672
rect 22004 8632 22005 8672
rect 21963 8623 22005 8632
rect 22059 8672 22101 8681
rect 22059 8632 22060 8672
rect 22100 8632 22101 8672
rect 22059 8623 22101 8632
rect 22539 8672 22581 8681
rect 22539 8632 22540 8672
rect 22580 8632 22581 8672
rect 22539 8623 22581 8632
rect 23011 8672 23069 8673
rect 23011 8632 23020 8672
rect 23060 8632 23069 8672
rect 23547 8641 23548 8681
rect 23588 8641 23589 8681
rect 23547 8632 23589 8641
rect 25419 8672 25461 8681
rect 25419 8632 25420 8672
rect 25460 8632 25461 8672
rect 23011 8631 23069 8632
rect 25419 8623 25461 8632
rect 25515 8672 25557 8681
rect 25515 8632 25516 8672
rect 25556 8632 25557 8672
rect 25515 8623 25557 8632
rect 25899 8672 25941 8681
rect 25899 8632 25900 8672
rect 25940 8632 25941 8672
rect 25899 8623 25941 8632
rect 25995 8672 26037 8681
rect 25995 8632 25996 8672
rect 26036 8632 26037 8672
rect 25995 8623 26037 8632
rect 26467 8672 26525 8673
rect 26467 8632 26476 8672
rect 26516 8632 26525 8672
rect 27003 8641 27004 8681
rect 27044 8641 27045 8681
rect 27003 8632 27045 8641
rect 27523 8672 27581 8673
rect 27523 8632 27532 8672
rect 27572 8632 27581 8672
rect 26467 8631 26525 8632
rect 27523 8631 27581 8632
rect 28771 8672 28829 8673
rect 28771 8632 28780 8672
rect 28820 8632 28829 8672
rect 28771 8631 28829 8632
rect 30115 8672 30173 8673
rect 30115 8632 30124 8672
rect 30164 8632 30173 8672
rect 30115 8631 30173 8632
rect 31363 8672 31421 8673
rect 31363 8632 31372 8672
rect 31412 8632 31421 8672
rect 31363 8631 31421 8632
rect 33955 8672 34013 8673
rect 33955 8632 33964 8672
rect 34004 8632 34013 8672
rect 33955 8631 34013 8632
rect 34819 8672 34877 8673
rect 34819 8632 34828 8672
rect 34868 8632 34877 8672
rect 34819 8631 34877 8632
rect 36931 8672 36989 8673
rect 36931 8632 36940 8672
rect 36980 8632 36989 8672
rect 36931 8631 36989 8632
rect 38179 8672 38237 8673
rect 38179 8632 38188 8672
rect 38228 8632 38237 8672
rect 38179 8631 38237 8632
rect 3051 8588 3093 8597
rect 3051 8548 3052 8588
rect 3092 8548 3093 8588
rect 3051 8539 3093 8548
rect 17355 8588 17397 8597
rect 17355 8548 17356 8588
rect 17396 8548 17397 8588
rect 17355 8539 17397 8548
rect 21675 8588 21717 8597
rect 21675 8548 21676 8588
rect 21716 8548 21717 8588
rect 21675 8539 21717 8548
rect 27339 8588 27381 8597
rect 27339 8548 27340 8588
rect 27380 8548 27381 8588
rect 27339 8539 27381 8548
rect 33579 8588 33621 8597
rect 33579 8548 33580 8588
rect 33620 8548 33621 8588
rect 33579 8539 33621 8548
rect 6219 8504 6261 8513
rect 6219 8464 6220 8504
rect 6260 8464 6261 8504
rect 6219 8455 6261 8464
rect 7851 8504 7893 8513
rect 7851 8464 7852 8504
rect 7892 8464 7893 8504
rect 7851 8455 7893 8464
rect 11115 8504 11157 8513
rect 11115 8464 11116 8504
rect 11156 8464 11157 8504
rect 11115 8455 11157 8464
rect 19371 8504 19413 8513
rect 19371 8464 19372 8504
rect 19412 8464 19413 8504
rect 19371 8455 19413 8464
rect 23691 8504 23733 8513
rect 23691 8464 23692 8504
rect 23732 8464 23733 8504
rect 23691 8455 23733 8464
rect 27147 8504 27189 8513
rect 27147 8464 27148 8504
rect 27188 8464 27189 8504
rect 27147 8455 27189 8464
rect 31563 8504 31605 8513
rect 31563 8464 31564 8504
rect 31604 8464 31605 8504
rect 31563 8455 31605 8464
rect 35971 8504 36029 8505
rect 35971 8464 35980 8504
rect 36020 8464 36029 8504
rect 35971 8463 36029 8464
rect 38379 8504 38421 8513
rect 38379 8464 38380 8504
rect 38420 8464 38421 8504
rect 38379 8455 38421 8464
rect 1152 8336 41856 8360
rect 1152 8296 4928 8336
rect 4968 8296 5010 8336
rect 5050 8296 5092 8336
rect 5132 8296 5174 8336
rect 5214 8296 5256 8336
rect 5296 8296 20048 8336
rect 20088 8296 20130 8336
rect 20170 8296 20212 8336
rect 20252 8296 20294 8336
rect 20334 8296 20376 8336
rect 20416 8296 35168 8336
rect 35208 8296 35250 8336
rect 35290 8296 35332 8336
rect 35372 8296 35414 8336
rect 35454 8296 35496 8336
rect 35536 8296 41856 8336
rect 1152 8272 41856 8296
rect 2859 8168 2901 8177
rect 2859 8128 2860 8168
rect 2900 8128 2901 8168
rect 2859 8119 2901 8128
rect 8323 8168 8381 8169
rect 8323 8128 8332 8168
rect 8372 8128 8381 8168
rect 8323 8127 8381 8128
rect 10347 8168 10389 8177
rect 10347 8128 10348 8168
rect 10388 8128 10389 8168
rect 10347 8119 10389 8128
rect 22539 8168 22581 8177
rect 22539 8128 22540 8168
rect 22580 8128 22581 8168
rect 22539 8119 22581 8128
rect 33291 8168 33333 8177
rect 33291 8128 33292 8168
rect 33332 8128 33333 8168
rect 33291 8119 33333 8128
rect 40683 8168 40725 8177
rect 40683 8128 40684 8168
rect 40724 8128 40725 8168
rect 40683 8119 40725 8128
rect 41451 8168 41493 8177
rect 41451 8128 41452 8168
rect 41492 8128 41493 8168
rect 41451 8119 41493 8128
rect 7371 8084 7413 8093
rect 7371 8044 7372 8084
rect 7412 8044 7413 8084
rect 7371 8035 7413 8044
rect 27051 8084 27093 8093
rect 27051 8044 27052 8084
rect 27092 8044 27093 8084
rect 27051 8035 27093 8044
rect 30411 8084 30453 8093
rect 30411 8044 30412 8084
rect 30452 8044 30453 8084
rect 30411 8035 30453 8044
rect 32811 8084 32853 8093
rect 32811 8044 32812 8084
rect 32852 8044 32853 8084
rect 32811 8035 32853 8044
rect 1411 8000 1469 8001
rect 1411 7960 1420 8000
rect 1460 7960 1469 8000
rect 1411 7959 1469 7960
rect 2659 8000 2717 8001
rect 2659 7960 2668 8000
rect 2708 7960 2717 8000
rect 2659 7959 2717 7960
rect 3043 8000 3101 8001
rect 3043 7960 3052 8000
rect 3092 7960 3101 8000
rect 3043 7959 3101 7960
rect 3435 8000 3477 8009
rect 3435 7960 3436 8000
rect 3476 7960 3477 8000
rect 3435 7951 3477 7960
rect 3531 8000 3573 8009
rect 3531 7960 3532 8000
rect 3572 7960 3573 8000
rect 3531 7951 3573 7960
rect 3627 8000 3669 8009
rect 3627 7960 3628 8000
rect 3668 7960 3669 8000
rect 3627 7951 3669 7960
rect 4003 8000 4061 8001
rect 4003 7960 4012 8000
rect 4052 7960 4061 8000
rect 4003 7959 4061 7960
rect 5251 8000 5309 8001
rect 5251 7960 5260 8000
rect 5300 7960 5309 8000
rect 5251 7959 5309 7960
rect 5923 8000 5981 8001
rect 5923 7960 5932 8000
rect 5972 7960 5981 8000
rect 5923 7959 5981 7960
rect 7171 8000 7229 8001
rect 7171 7960 7180 8000
rect 7220 7960 7229 8000
rect 7171 7959 7229 7960
rect 7851 8000 7893 8009
rect 7851 7960 7852 8000
rect 7892 7960 7893 8000
rect 7851 7951 7893 7960
rect 7947 8000 7989 8009
rect 7947 7960 7948 8000
rect 7988 7960 7989 8000
rect 7947 7951 7989 7960
rect 8043 8000 8085 8009
rect 8043 7960 8044 8000
rect 8084 7960 8085 8000
rect 8043 7951 8085 7960
rect 8139 8000 8181 8009
rect 8139 7960 8140 8000
rect 8180 7960 8181 8000
rect 8139 7951 8181 7960
rect 8523 8000 8565 8009
rect 8523 7960 8524 8000
rect 8564 7960 8565 8000
rect 8523 7951 8565 7960
rect 8619 8000 8661 8009
rect 8619 7960 8620 8000
rect 8660 7960 8661 8000
rect 8619 7951 8661 7960
rect 8899 8000 8957 8001
rect 8899 7960 8908 8000
rect 8948 7960 8957 8000
rect 8899 7959 8957 7960
rect 10147 8000 10205 8001
rect 10147 7960 10156 8000
rect 10196 7960 10205 8000
rect 10147 7959 10205 7960
rect 10531 8000 10589 8001
rect 10531 7960 10540 8000
rect 10580 7960 10589 8000
rect 10531 7959 10589 7960
rect 11779 8000 11837 8001
rect 11779 7960 11788 8000
rect 11828 7960 11837 8000
rect 11779 7959 11837 7960
rect 12163 8000 12221 8001
rect 12163 7960 12172 8000
rect 12212 7960 12221 8000
rect 12163 7959 12221 7960
rect 13411 8000 13469 8001
rect 13411 7960 13420 8000
rect 13460 7960 13469 8000
rect 13411 7959 13469 7960
rect 13795 8000 13853 8001
rect 13795 7960 13804 8000
rect 13844 7960 13853 8000
rect 13795 7959 13853 7960
rect 15043 8000 15101 8001
rect 15043 7960 15052 8000
rect 15092 7960 15101 8000
rect 15043 7959 15101 7960
rect 16099 8000 16157 8001
rect 16099 7960 16108 8000
rect 16148 7960 16157 8000
rect 16099 7959 16157 7960
rect 17347 8000 17405 8001
rect 17347 7960 17356 8000
rect 17396 7960 17405 8000
rect 17347 7959 17405 7960
rect 17827 8000 17885 8001
rect 17827 7960 17836 8000
rect 17876 7960 17885 8000
rect 17827 7959 17885 7960
rect 19075 8000 19133 8001
rect 19075 7960 19084 8000
rect 19124 7960 19133 8000
rect 19075 7959 19133 7960
rect 19747 8000 19805 8001
rect 19747 7960 19756 8000
rect 19796 7960 19805 8000
rect 19747 7959 19805 7960
rect 20995 8000 21053 8001
rect 20995 7960 21004 8000
rect 21044 7960 21053 8000
rect 20995 7959 21053 7960
rect 22819 8000 22877 8001
rect 22819 7960 22828 8000
rect 22868 7960 22877 8000
rect 22819 7959 22877 7960
rect 24067 8000 24125 8001
rect 24067 7960 24076 8000
rect 24116 7960 24125 8000
rect 24067 7959 24125 7960
rect 25323 8000 25365 8009
rect 25323 7960 25324 8000
rect 25364 7960 25365 8000
rect 25323 7951 25365 7960
rect 25419 8000 25461 8009
rect 25419 7960 25420 8000
rect 25460 7960 25461 8000
rect 25419 7951 25461 7960
rect 25899 8000 25941 8009
rect 25899 7960 25900 8000
rect 25940 7960 25941 8000
rect 25899 7951 25941 7960
rect 26371 8000 26429 8001
rect 26371 7960 26380 8000
rect 26420 7960 26429 8000
rect 28683 8000 28725 8009
rect 26371 7959 26429 7960
rect 26859 7986 26901 7995
rect 26859 7946 26860 7986
rect 26900 7946 26901 7986
rect 28683 7960 28684 8000
rect 28724 7960 28725 8000
rect 28683 7951 28725 7960
rect 28779 8000 28821 8009
rect 28779 7960 28780 8000
rect 28820 7960 28821 8000
rect 28779 7951 28821 7960
rect 29731 8000 29789 8001
rect 29731 7960 29740 8000
rect 29780 7960 29789 8000
rect 31083 8000 31125 8009
rect 29731 7959 29789 7960
rect 30267 7958 30309 7967
rect 26859 7937 26901 7946
rect 3147 7916 3189 7925
rect 3147 7876 3148 7916
rect 3188 7876 3189 7916
rect 3147 7867 3189 7876
rect 21571 7916 21629 7917
rect 21571 7876 21580 7916
rect 21620 7876 21629 7916
rect 21571 7875 21629 7876
rect 22339 7916 22397 7917
rect 22339 7876 22348 7916
rect 22388 7876 22397 7916
rect 22339 7875 22397 7876
rect 25803 7916 25845 7925
rect 25803 7876 25804 7916
rect 25844 7876 25845 7916
rect 25803 7867 25845 7876
rect 27427 7916 27485 7917
rect 27427 7876 27436 7916
rect 27476 7876 27485 7916
rect 27427 7875 27485 7876
rect 29163 7916 29205 7925
rect 29163 7876 29164 7916
rect 29204 7876 29205 7916
rect 29163 7867 29205 7876
rect 29259 7916 29301 7925
rect 29259 7876 29260 7916
rect 29300 7876 29301 7916
rect 30267 7918 30268 7958
rect 30308 7918 30309 7958
rect 31083 7960 31084 8000
rect 31124 7960 31125 8000
rect 31083 7951 31125 7960
rect 31179 8000 31221 8009
rect 31179 7960 31180 8000
rect 31220 7960 31221 8000
rect 31179 7951 31221 7960
rect 32131 8000 32189 8001
rect 32131 7960 32140 8000
rect 32180 7960 32189 8000
rect 34059 8000 34101 8009
rect 32131 7959 32189 7960
rect 32619 7986 32661 7995
rect 32619 7946 32620 7986
rect 32660 7946 32661 7986
rect 34059 7960 34060 8000
rect 34100 7960 34101 8000
rect 34059 7951 34101 7960
rect 34435 8000 34493 8001
rect 34435 7960 34444 8000
rect 34484 7960 34493 8000
rect 34435 7959 34493 7960
rect 35299 8000 35357 8001
rect 35299 7960 35308 8000
rect 35348 7960 35357 8000
rect 35299 7959 35357 7960
rect 36835 8000 36893 8001
rect 36835 7960 36844 8000
rect 36884 7960 36893 8000
rect 36835 7959 36893 7960
rect 38083 8000 38141 8001
rect 38083 7960 38092 8000
rect 38132 7960 38141 8000
rect 38083 7959 38141 7960
rect 32619 7937 32661 7946
rect 30267 7909 30309 7918
rect 30787 7916 30845 7917
rect 29259 7867 29301 7876
rect 30787 7876 30796 7916
rect 30836 7876 30845 7916
rect 30787 7875 30845 7876
rect 31563 7916 31605 7925
rect 31563 7876 31564 7916
rect 31604 7876 31605 7916
rect 31563 7867 31605 7876
rect 31659 7916 31701 7925
rect 31659 7876 31660 7916
rect 31700 7876 31701 7916
rect 31659 7867 31701 7876
rect 33091 7916 33149 7917
rect 33091 7876 33100 7916
rect 33140 7876 33149 7916
rect 33091 7875 33149 7876
rect 40483 7916 40541 7917
rect 40483 7876 40492 7916
rect 40532 7876 40541 7916
rect 40483 7875 40541 7876
rect 40867 7916 40925 7917
rect 40867 7876 40876 7916
rect 40916 7876 40925 7916
rect 40867 7875 40925 7876
rect 41251 7916 41309 7917
rect 41251 7876 41260 7916
rect 41300 7876 41309 7916
rect 41251 7875 41309 7876
rect 30603 7832 30645 7841
rect 30603 7792 30604 7832
rect 30644 7792 30645 7832
rect 30603 7783 30645 7792
rect 41067 7832 41109 7841
rect 41067 7792 41068 7832
rect 41108 7792 41109 7832
rect 41067 7783 41109 7792
rect 2859 7748 2901 7757
rect 2859 7708 2860 7748
rect 2900 7708 2901 7748
rect 2859 7699 2901 7708
rect 3811 7748 3869 7749
rect 3811 7708 3820 7748
rect 3860 7708 3869 7748
rect 3811 7707 3869 7708
rect 5451 7748 5493 7757
rect 5451 7708 5452 7748
rect 5492 7708 5493 7748
rect 5451 7699 5493 7708
rect 11979 7748 12021 7757
rect 11979 7708 11980 7748
rect 12020 7708 12021 7748
rect 11979 7699 12021 7708
rect 13611 7748 13653 7757
rect 13611 7708 13612 7748
rect 13652 7708 13653 7748
rect 13611 7699 13653 7708
rect 15243 7748 15285 7757
rect 15243 7708 15244 7748
rect 15284 7708 15285 7748
rect 15243 7699 15285 7708
rect 17547 7748 17589 7757
rect 17547 7708 17548 7748
rect 17588 7708 17589 7748
rect 17547 7699 17589 7708
rect 19275 7748 19317 7757
rect 19275 7708 19276 7748
rect 19316 7708 19317 7748
rect 19275 7699 19317 7708
rect 21195 7748 21237 7757
rect 21195 7708 21196 7748
rect 21236 7708 21237 7748
rect 21195 7699 21237 7708
rect 21387 7748 21429 7757
rect 21387 7708 21388 7748
rect 21428 7708 21429 7748
rect 21387 7699 21429 7708
rect 24267 7748 24309 7757
rect 24267 7708 24268 7748
rect 24308 7708 24309 7748
rect 24267 7699 24309 7708
rect 27243 7748 27285 7757
rect 27243 7708 27244 7748
rect 27284 7708 27285 7748
rect 27243 7699 27285 7708
rect 36451 7748 36509 7749
rect 36451 7708 36460 7748
rect 36500 7708 36509 7748
rect 36451 7707 36509 7708
rect 36651 7748 36693 7757
rect 36651 7708 36652 7748
rect 36692 7708 36693 7748
rect 36651 7699 36693 7708
rect 1152 7580 41856 7604
rect 1152 7540 3688 7580
rect 3728 7540 3770 7580
rect 3810 7540 3852 7580
rect 3892 7540 3934 7580
rect 3974 7540 4016 7580
rect 4056 7540 18808 7580
rect 18848 7540 18890 7580
rect 18930 7540 18972 7580
rect 19012 7540 19054 7580
rect 19094 7540 19136 7580
rect 19176 7540 33928 7580
rect 33968 7540 34010 7580
rect 34050 7540 34092 7580
rect 34132 7540 34174 7580
rect 34214 7540 34256 7580
rect 34296 7540 41856 7580
rect 1152 7516 41856 7540
rect 3723 7412 3765 7421
rect 3723 7372 3724 7412
rect 3764 7372 3765 7412
rect 3723 7363 3765 7372
rect 25611 7412 25653 7421
rect 25611 7372 25612 7412
rect 25652 7372 25653 7412
rect 25611 7363 25653 7372
rect 26283 7412 26325 7421
rect 26283 7372 26284 7412
rect 26324 7372 26325 7412
rect 26283 7363 26325 7372
rect 30315 7412 30357 7421
rect 30315 7372 30316 7412
rect 30356 7372 30357 7412
rect 30315 7363 30357 7372
rect 33099 7412 33141 7421
rect 33099 7372 33100 7412
rect 33140 7372 33141 7412
rect 33099 7363 33141 7372
rect 40683 7412 40725 7421
rect 40683 7372 40684 7412
rect 40724 7372 40725 7412
rect 40683 7363 40725 7372
rect 4395 7328 4437 7337
rect 4395 7288 4396 7328
rect 4436 7288 4437 7328
rect 4395 7279 4437 7288
rect 7755 7244 7797 7253
rect 7755 7204 7756 7244
rect 7796 7204 7797 7244
rect 7755 7195 7797 7204
rect 14283 7244 14325 7253
rect 14283 7204 14284 7244
rect 14324 7204 14325 7244
rect 14283 7195 14325 7204
rect 14379 7244 14421 7253
rect 14379 7204 14380 7244
rect 14420 7204 14421 7244
rect 21379 7244 21437 7245
rect 14379 7195 14421 7204
rect 20859 7202 20901 7211
rect 21379 7204 21388 7244
rect 21428 7204 21437 7244
rect 21379 7203 21437 7204
rect 23395 7244 23453 7245
rect 23395 7204 23404 7244
rect 23444 7204 23453 7244
rect 23395 7203 23453 7204
rect 25891 7244 25949 7245
rect 25891 7204 25900 7244
rect 25940 7204 25949 7244
rect 25891 7203 25949 7204
rect 30691 7244 30749 7245
rect 30691 7204 30700 7244
rect 30740 7204 30749 7244
rect 30691 7203 30749 7204
rect 38475 7244 38517 7253
rect 38475 7204 38476 7244
rect 38516 7204 38517 7244
rect 8859 7169 8901 7178
rect 12843 7174 12885 7183
rect 2955 7160 2997 7169
rect 2955 7120 2956 7160
rect 2996 7120 2997 7160
rect 2955 7111 2997 7120
rect 3051 7160 3093 7169
rect 3051 7120 3052 7160
rect 3092 7120 3093 7160
rect 3051 7111 3093 7120
rect 3147 7160 3189 7169
rect 3147 7120 3148 7160
rect 3188 7120 3189 7160
rect 3147 7111 3189 7120
rect 3243 7160 3285 7169
rect 3243 7120 3244 7160
rect 3284 7120 3285 7160
rect 3243 7111 3285 7120
rect 3435 7160 3477 7169
rect 3435 7120 3436 7160
rect 3476 7120 3477 7160
rect 3435 7111 3477 7120
rect 3531 7160 3573 7169
rect 3531 7120 3532 7160
rect 3572 7120 3573 7160
rect 3531 7111 3573 7120
rect 4395 7152 4437 7161
rect 4395 7112 4396 7152
rect 4436 7112 4437 7152
rect 4395 7103 4437 7112
rect 4779 7160 4821 7169
rect 4779 7120 4780 7160
rect 4820 7120 4821 7160
rect 4779 7111 4821 7120
rect 4875 7160 4917 7169
rect 4875 7120 4876 7160
rect 4916 7120 4917 7160
rect 4875 7111 4917 7120
rect 5259 7160 5301 7169
rect 5259 7120 5260 7160
rect 5300 7120 5301 7160
rect 5259 7111 5301 7120
rect 5355 7160 5397 7169
rect 5355 7120 5356 7160
rect 5396 7120 5397 7160
rect 5355 7111 5397 7120
rect 5451 7160 5493 7169
rect 5451 7120 5452 7160
rect 5492 7120 5493 7160
rect 5451 7111 5493 7120
rect 5547 7160 5589 7169
rect 5547 7120 5548 7160
rect 5588 7120 5589 7160
rect 5547 7111 5589 7120
rect 5739 7160 5781 7169
rect 5739 7120 5740 7160
rect 5780 7120 5781 7160
rect 5739 7111 5781 7120
rect 5835 7160 5877 7169
rect 5835 7120 5836 7160
rect 5876 7120 5877 7160
rect 5835 7111 5877 7120
rect 5931 7160 5973 7169
rect 5931 7120 5932 7160
rect 5972 7120 5973 7160
rect 5931 7111 5973 7120
rect 6027 7160 6069 7169
rect 6027 7120 6028 7160
rect 6068 7120 6069 7160
rect 6027 7111 6069 7120
rect 6219 7160 6261 7169
rect 6219 7120 6220 7160
rect 6260 7120 6261 7160
rect 6219 7111 6261 7120
rect 6315 7160 6357 7169
rect 6315 7120 6316 7160
rect 6356 7120 6357 7160
rect 6315 7111 6357 7120
rect 6795 7160 6837 7169
rect 6795 7120 6796 7160
rect 6836 7120 6837 7160
rect 6795 7111 6837 7120
rect 6891 7160 6933 7169
rect 6891 7120 6892 7160
rect 6932 7120 6933 7160
rect 6891 7111 6933 7120
rect 6987 7160 7029 7169
rect 6987 7120 6988 7160
rect 7028 7120 7029 7160
rect 6987 7111 7029 7120
rect 7275 7160 7317 7169
rect 7275 7120 7276 7160
rect 7316 7120 7317 7160
rect 7275 7111 7317 7120
rect 7371 7160 7413 7169
rect 7371 7120 7372 7160
rect 7412 7120 7413 7160
rect 7371 7111 7413 7120
rect 7851 7160 7893 7169
rect 7851 7120 7852 7160
rect 7892 7120 7893 7160
rect 7851 7111 7893 7120
rect 8323 7160 8381 7161
rect 8323 7120 8332 7160
rect 8372 7120 8381 7160
rect 8859 7129 8860 7169
rect 8900 7129 8901 7169
rect 8859 7120 8901 7129
rect 9195 7160 9237 7169
rect 9195 7120 9196 7160
rect 9236 7120 9237 7160
rect 8323 7119 8381 7120
rect 9195 7111 9237 7120
rect 9291 7160 9333 7169
rect 9291 7120 9292 7160
rect 9332 7120 9333 7160
rect 9291 7111 9333 7120
rect 9675 7160 9717 7169
rect 9675 7120 9676 7160
rect 9716 7120 9717 7160
rect 9675 7111 9717 7120
rect 9771 7160 9813 7169
rect 9771 7120 9772 7160
rect 9812 7120 9813 7160
rect 9771 7111 9813 7120
rect 9867 7160 9909 7169
rect 9867 7120 9868 7160
rect 9908 7120 9909 7160
rect 9867 7111 9909 7120
rect 9963 7160 10005 7169
rect 9963 7120 9964 7160
rect 10004 7120 10005 7160
rect 9963 7111 10005 7120
rect 11307 7160 11349 7169
rect 11307 7120 11308 7160
rect 11348 7120 11349 7160
rect 11307 7111 11349 7120
rect 11403 7160 11445 7169
rect 11403 7120 11404 7160
rect 11444 7120 11445 7160
rect 11403 7111 11445 7120
rect 11787 7160 11829 7169
rect 11787 7120 11788 7160
rect 11828 7120 11829 7160
rect 11787 7111 11829 7120
rect 11883 7160 11925 7169
rect 11883 7120 11884 7160
rect 11924 7120 11925 7160
rect 11883 7111 11925 7120
rect 12355 7160 12413 7161
rect 12355 7120 12364 7160
rect 12404 7120 12413 7160
rect 12843 7134 12844 7174
rect 12884 7134 12885 7174
rect 15339 7174 15381 7183
rect 12843 7125 12885 7134
rect 13803 7160 13845 7169
rect 12355 7119 12413 7120
rect 13803 7120 13804 7160
rect 13844 7120 13845 7160
rect 13803 7111 13845 7120
rect 13899 7160 13941 7169
rect 13899 7120 13900 7160
rect 13940 7120 13941 7160
rect 13899 7111 13941 7120
rect 14851 7160 14909 7161
rect 14851 7120 14860 7160
rect 14900 7120 14909 7160
rect 15339 7134 15340 7174
rect 15380 7134 15381 7174
rect 15339 7125 15381 7134
rect 16291 7160 16349 7161
rect 14851 7119 14909 7120
rect 16291 7120 16300 7160
rect 16340 7120 16349 7160
rect 16291 7119 16349 7120
rect 17539 7160 17597 7161
rect 17539 7120 17548 7160
rect 17588 7120 17597 7160
rect 17539 7119 17597 7120
rect 19275 7160 19317 7169
rect 19275 7120 19276 7160
rect 19316 7120 19317 7160
rect 19275 7111 19317 7120
rect 19371 7160 19413 7169
rect 19371 7120 19372 7160
rect 19412 7120 19413 7160
rect 19371 7111 19413 7120
rect 19755 7160 19797 7169
rect 19755 7120 19756 7160
rect 19796 7120 19797 7160
rect 19755 7111 19797 7120
rect 19851 7160 19893 7169
rect 20859 7162 20860 7202
rect 20900 7162 20901 7202
rect 38475 7195 38517 7204
rect 40483 7244 40541 7245
rect 40483 7204 40492 7244
rect 40532 7204 40541 7244
rect 40483 7203 40541 7204
rect 40867 7244 40925 7245
rect 40867 7204 40876 7244
rect 40916 7204 40925 7244
rect 40867 7203 40925 7204
rect 36651 7174 36693 7183
rect 19851 7120 19852 7160
rect 19892 7120 19893 7160
rect 19851 7111 19893 7120
rect 20323 7160 20381 7161
rect 20323 7120 20332 7160
rect 20372 7120 20381 7160
rect 20859 7153 20901 7162
rect 24163 7160 24221 7161
rect 20323 7119 20381 7120
rect 24163 7120 24172 7160
rect 24212 7120 24221 7160
rect 24163 7119 24221 7120
rect 25411 7160 25469 7161
rect 25411 7120 25420 7160
rect 25460 7120 25469 7160
rect 25411 7119 25469 7120
rect 26467 7160 26525 7161
rect 26467 7120 26476 7160
rect 26516 7120 26525 7160
rect 26467 7119 26525 7120
rect 27715 7160 27773 7161
rect 27715 7120 27724 7160
rect 27764 7120 27773 7160
rect 27715 7119 27773 7120
rect 28867 7160 28925 7161
rect 28867 7120 28876 7160
rect 28916 7120 28925 7160
rect 28867 7119 28925 7120
rect 30115 7160 30173 7161
rect 30115 7120 30124 7160
rect 30164 7120 30173 7160
rect 30115 7119 30173 7120
rect 31651 7160 31709 7161
rect 31651 7120 31660 7160
rect 31700 7120 31709 7160
rect 31651 7119 31709 7120
rect 32899 7160 32957 7161
rect 32899 7120 32908 7160
rect 32948 7120 32957 7160
rect 32899 7119 32957 7120
rect 33379 7160 33437 7161
rect 33379 7120 33388 7160
rect 33428 7120 33437 7160
rect 33379 7119 33437 7120
rect 34627 7160 34685 7161
rect 34627 7120 34636 7160
rect 34676 7120 34685 7160
rect 34627 7119 34685 7120
rect 35115 7160 35157 7169
rect 35115 7120 35116 7160
rect 35156 7120 35157 7160
rect 35115 7111 35157 7120
rect 35211 7160 35253 7169
rect 35211 7120 35212 7160
rect 35252 7120 35253 7160
rect 35211 7111 35253 7120
rect 35595 7160 35637 7169
rect 35595 7120 35596 7160
rect 35636 7120 35637 7160
rect 35595 7111 35637 7120
rect 35691 7160 35733 7169
rect 35691 7120 35692 7160
rect 35732 7120 35733 7160
rect 35691 7111 35733 7120
rect 36163 7160 36221 7161
rect 36163 7120 36172 7160
rect 36212 7120 36221 7160
rect 36651 7134 36652 7174
rect 36692 7134 36693 7174
rect 36651 7125 36693 7134
rect 37995 7160 38037 7169
rect 36163 7119 36221 7120
rect 37995 7120 37996 7160
rect 38036 7120 38037 7160
rect 37995 7111 38037 7120
rect 38091 7160 38133 7169
rect 38091 7120 38092 7160
rect 38132 7120 38133 7160
rect 38091 7111 38133 7120
rect 38571 7160 38613 7169
rect 39531 7165 39573 7174
rect 38571 7120 38572 7160
rect 38612 7120 38613 7160
rect 38571 7111 38613 7120
rect 39043 7160 39101 7161
rect 39043 7120 39052 7160
rect 39092 7120 39101 7160
rect 39043 7119 39101 7120
rect 39531 7125 39532 7165
rect 39572 7125 39573 7165
rect 39531 7116 39573 7125
rect 3619 7076 3677 7077
rect 3619 7036 3628 7076
rect 3668 7036 3677 7076
rect 3619 7035 3677 7036
rect 9003 7076 9045 7085
rect 9003 7036 9004 7076
rect 9044 7036 9045 7076
rect 9003 7027 9045 7036
rect 21003 7076 21045 7085
rect 21003 7036 21004 7076
rect 21044 7036 21045 7076
rect 21003 7027 21045 7036
rect 34827 7076 34869 7085
rect 34827 7036 34828 7076
rect 34868 7036 34869 7076
rect 34827 7027 34869 7036
rect 3715 6992 3773 6993
rect 3715 6952 3724 6992
rect 3764 6952 3773 6992
rect 3715 6951 3773 6952
rect 4587 6992 4629 7001
rect 4587 6952 4588 6992
rect 4628 6952 4629 6992
rect 4587 6943 4629 6952
rect 5059 6992 5117 6993
rect 5059 6952 5068 6992
rect 5108 6952 5117 6992
rect 5059 6951 5117 6952
rect 6499 6992 6557 6993
rect 6499 6952 6508 6992
rect 6548 6952 6557 6992
rect 6499 6951 6557 6952
rect 6691 6992 6749 6993
rect 6691 6952 6700 6992
rect 6740 6952 6749 6992
rect 6691 6951 6749 6952
rect 9475 6992 9533 6993
rect 9475 6952 9484 6992
rect 9524 6952 9533 6992
rect 9475 6951 9533 6952
rect 13035 6992 13077 7001
rect 13035 6952 13036 6992
rect 13076 6952 13077 6992
rect 13035 6943 13077 6952
rect 15531 6992 15573 7001
rect 15531 6952 15532 6992
rect 15572 6952 15573 6992
rect 15531 6943 15573 6952
rect 17739 6992 17781 7001
rect 17739 6952 17740 6992
rect 17780 6952 17781 6992
rect 17739 6943 17781 6952
rect 21195 6992 21237 7001
rect 21195 6952 21196 6992
rect 21236 6952 21237 6992
rect 21195 6943 21237 6952
rect 23211 6992 23253 7001
rect 23211 6952 23212 6992
rect 23252 6952 23253 6992
rect 23211 6943 23253 6952
rect 26091 6992 26133 7001
rect 26091 6952 26092 6992
rect 26132 6952 26133 6992
rect 26091 6943 26133 6952
rect 30507 6992 30549 7001
rect 30507 6952 30508 6992
rect 30548 6952 30549 6992
rect 30507 6943 30549 6952
rect 36843 6992 36885 7001
rect 36843 6952 36844 6992
rect 36884 6952 36885 6992
rect 36843 6943 36885 6952
rect 39723 6992 39765 7001
rect 39723 6952 39724 6992
rect 39764 6952 39765 6992
rect 39723 6943 39765 6952
rect 41067 6992 41109 7001
rect 41067 6952 41068 6992
rect 41108 6952 41109 6992
rect 41067 6943 41109 6952
rect 1152 6824 41856 6848
rect 1152 6784 4928 6824
rect 4968 6784 5010 6824
rect 5050 6784 5092 6824
rect 5132 6784 5174 6824
rect 5214 6784 5256 6824
rect 5296 6784 20048 6824
rect 20088 6784 20130 6824
rect 20170 6784 20212 6824
rect 20252 6784 20294 6824
rect 20334 6784 20376 6824
rect 20416 6784 35168 6824
rect 35208 6784 35250 6824
rect 35290 6784 35332 6824
rect 35372 6784 35414 6824
rect 35454 6784 35496 6824
rect 35536 6784 41856 6824
rect 1152 6760 41856 6784
rect 5827 6656 5885 6657
rect 5827 6616 5836 6656
rect 5876 6616 5885 6656
rect 5827 6615 5885 6616
rect 6307 6656 6365 6657
rect 6307 6616 6316 6656
rect 6356 6616 6365 6656
rect 6307 6615 6365 6616
rect 9003 6656 9045 6665
rect 9003 6616 9004 6656
rect 9044 6616 9045 6656
rect 9003 6607 9045 6616
rect 21291 6656 21333 6665
rect 21291 6616 21292 6656
rect 21332 6616 21333 6656
rect 21291 6607 21333 6616
rect 37323 6656 37365 6665
rect 37323 6616 37324 6656
rect 37364 6616 37365 6656
rect 37323 6607 37365 6616
rect 39435 6656 39477 6665
rect 39435 6616 39436 6656
rect 39476 6616 39477 6656
rect 39435 6607 39477 6616
rect 40683 6656 40725 6665
rect 40683 6616 40684 6656
rect 40724 6616 40725 6656
rect 40683 6607 40725 6616
rect 3531 6572 3573 6581
rect 3531 6532 3532 6572
rect 3572 6532 3573 6572
rect 3531 6523 3573 6532
rect 6795 6572 6837 6581
rect 6795 6532 6796 6572
rect 6836 6532 6837 6572
rect 6795 6523 6837 6532
rect 19659 6572 19701 6581
rect 19659 6532 19660 6572
rect 19700 6532 19701 6572
rect 19659 6523 19701 6532
rect 23307 6572 23349 6581
rect 23307 6532 23308 6572
rect 23348 6532 23349 6572
rect 23307 6523 23349 6532
rect 1699 6488 1757 6489
rect 1699 6448 1708 6488
rect 1748 6448 1757 6488
rect 1699 6447 1757 6448
rect 2947 6488 3005 6489
rect 2947 6448 2956 6488
rect 2996 6448 3005 6488
rect 2947 6447 3005 6448
rect 3435 6488 3477 6497
rect 3435 6448 3436 6488
rect 3476 6448 3477 6488
rect 3435 6439 3477 6448
rect 3619 6488 3677 6489
rect 3619 6448 3628 6488
rect 3668 6448 3677 6488
rect 3619 6447 3677 6448
rect 3907 6488 3965 6489
rect 3907 6448 3916 6488
rect 3956 6448 3965 6488
rect 3907 6447 3965 6448
rect 4203 6488 4245 6497
rect 4203 6448 4204 6488
rect 4244 6448 4245 6488
rect 4203 6439 4245 6448
rect 4299 6488 4341 6497
rect 4299 6448 4300 6488
rect 4340 6448 4341 6488
rect 4299 6439 4341 6448
rect 4862 6488 4920 6489
rect 4862 6448 4871 6488
rect 4911 6448 4920 6488
rect 4862 6447 4920 6448
rect 4971 6488 5013 6497
rect 4971 6448 4972 6488
rect 5012 6448 5013 6488
rect 4971 6439 5013 6448
rect 5067 6488 5109 6497
rect 5067 6448 5068 6488
rect 5108 6448 5109 6488
rect 5067 6439 5109 6448
rect 5251 6488 5309 6489
rect 5251 6448 5260 6488
rect 5300 6448 5309 6488
rect 5251 6447 5309 6448
rect 5347 6488 5405 6489
rect 5347 6448 5356 6488
rect 5396 6448 5405 6488
rect 5347 6447 5405 6448
rect 5547 6488 5589 6497
rect 5547 6448 5548 6488
rect 5588 6448 5589 6488
rect 5547 6439 5589 6448
rect 5643 6488 5685 6497
rect 5643 6448 5644 6488
rect 5684 6448 5685 6488
rect 5643 6439 5685 6448
rect 5739 6488 5781 6497
rect 5739 6448 5740 6488
rect 5780 6448 5781 6488
rect 5739 6439 5781 6448
rect 6027 6488 6069 6497
rect 6027 6448 6028 6488
rect 6068 6448 6069 6488
rect 6027 6439 6069 6448
rect 6123 6488 6165 6497
rect 6123 6448 6124 6488
rect 6164 6448 6165 6488
rect 6123 6439 6165 6448
rect 6219 6488 6261 6497
rect 6219 6448 6220 6488
rect 6260 6448 6261 6488
rect 6219 6439 6261 6448
rect 6891 6488 6933 6497
rect 6891 6448 6892 6488
rect 6932 6448 6933 6488
rect 6891 6439 6933 6448
rect 7171 6488 7229 6489
rect 7171 6448 7180 6488
rect 7220 6448 7229 6488
rect 7171 6447 7229 6448
rect 7555 6488 7613 6489
rect 7555 6448 7564 6488
rect 7604 6448 7613 6488
rect 7555 6447 7613 6448
rect 8803 6488 8861 6489
rect 8803 6448 8812 6488
rect 8852 6448 8861 6488
rect 8803 6447 8861 6448
rect 9859 6488 9917 6489
rect 9859 6448 9868 6488
rect 9908 6448 9917 6488
rect 9859 6447 9917 6448
rect 11107 6488 11165 6489
rect 11107 6448 11116 6488
rect 11156 6448 11165 6488
rect 11107 6447 11165 6448
rect 12259 6488 12317 6489
rect 12259 6448 12268 6488
rect 12308 6448 12317 6488
rect 12259 6447 12317 6448
rect 13507 6488 13565 6489
rect 13507 6448 13516 6488
rect 13556 6448 13565 6488
rect 13507 6447 13565 6448
rect 14755 6488 14813 6489
rect 14755 6448 14764 6488
rect 14804 6448 14813 6488
rect 14755 6447 14813 6448
rect 16003 6488 16061 6489
rect 16003 6448 16012 6488
rect 16052 6448 16061 6488
rect 16003 6447 16061 6448
rect 17931 6488 17973 6497
rect 17931 6448 17932 6488
rect 17972 6448 17973 6488
rect 17931 6439 17973 6448
rect 18027 6488 18069 6497
rect 18027 6448 18028 6488
rect 18068 6448 18069 6488
rect 18027 6439 18069 6448
rect 18411 6488 18453 6497
rect 18411 6448 18412 6488
rect 18452 6448 18453 6488
rect 18411 6439 18453 6448
rect 18979 6488 19037 6489
rect 18979 6448 18988 6488
rect 19028 6448 19037 6488
rect 19843 6488 19901 6489
rect 18979 6447 19037 6448
rect 19467 6474 19509 6483
rect 19467 6434 19468 6474
rect 19508 6434 19509 6474
rect 19843 6448 19852 6488
rect 19892 6448 19901 6488
rect 19843 6447 19901 6448
rect 21091 6488 21149 6489
rect 21091 6448 21100 6488
rect 21140 6448 21149 6488
rect 21091 6447 21149 6448
rect 21579 6488 21621 6497
rect 21579 6448 21580 6488
rect 21620 6448 21621 6488
rect 21579 6439 21621 6448
rect 21675 6488 21717 6497
rect 21675 6448 21676 6488
rect 21716 6448 21717 6488
rect 21675 6439 21717 6448
rect 22059 6488 22101 6497
rect 22059 6448 22060 6488
rect 22100 6448 22101 6488
rect 22059 6439 22101 6448
rect 22627 6488 22685 6489
rect 22627 6448 22636 6488
rect 22676 6448 22685 6488
rect 24355 6488 24413 6489
rect 22627 6447 22685 6448
rect 23163 6446 23205 6455
rect 24355 6448 24364 6488
rect 24404 6448 24413 6488
rect 24355 6447 24413 6448
rect 25603 6488 25661 6489
rect 25603 6448 25612 6488
rect 25652 6448 25661 6488
rect 25603 6447 25661 6448
rect 26467 6488 26525 6489
rect 26467 6448 26476 6488
rect 26516 6448 26525 6488
rect 26467 6447 26525 6448
rect 27715 6488 27773 6489
rect 27715 6448 27724 6488
rect 27764 6448 27773 6488
rect 27715 6447 27773 6448
rect 28291 6488 28349 6489
rect 28291 6448 28300 6488
rect 28340 6448 28349 6488
rect 28291 6447 28349 6448
rect 29539 6488 29597 6489
rect 29539 6448 29548 6488
rect 29588 6448 29597 6488
rect 29539 6447 29597 6448
rect 30499 6488 30557 6489
rect 30499 6448 30508 6488
rect 30548 6448 30557 6488
rect 30499 6447 30557 6448
rect 32515 6488 32573 6489
rect 32515 6448 32524 6488
rect 32564 6448 32573 6488
rect 32515 6447 32573 6448
rect 33763 6488 33821 6489
rect 33763 6448 33772 6488
rect 33812 6448 33821 6488
rect 33763 6447 33821 6448
rect 36939 6488 36981 6497
rect 36939 6448 36940 6488
rect 36980 6448 36981 6488
rect 19467 6425 19509 6434
rect 18507 6404 18549 6413
rect 18507 6364 18508 6404
rect 18548 6364 18549 6404
rect 18507 6355 18549 6364
rect 22155 6404 22197 6413
rect 22155 6364 22156 6404
rect 22196 6364 22197 6404
rect 23163 6406 23164 6446
rect 23204 6406 23205 6446
rect 23163 6397 23205 6406
rect 31747 6446 31805 6447
rect 31747 6406 31756 6446
rect 31796 6406 31805 6446
rect 36939 6439 36981 6448
rect 37987 6488 38045 6489
rect 37987 6448 37996 6488
rect 38036 6448 38045 6488
rect 37987 6447 38045 6448
rect 39235 6488 39293 6489
rect 39235 6448 39244 6488
rect 39284 6448 39293 6488
rect 39235 6447 39293 6448
rect 31747 6405 31805 6406
rect 23683 6404 23741 6405
rect 22155 6355 22197 6364
rect 23683 6364 23692 6404
rect 23732 6364 23741 6404
rect 23683 6363 23741 6364
rect 26275 6404 26333 6405
rect 26275 6364 26284 6404
rect 26324 6364 26333 6404
rect 26275 6363 26333 6364
rect 32323 6404 32381 6405
rect 32323 6364 32332 6404
rect 32372 6364 32381 6404
rect 32323 6363 32381 6364
rect 36547 6404 36605 6405
rect 36547 6364 36556 6404
rect 36596 6364 36605 6404
rect 36547 6363 36605 6364
rect 39811 6404 39869 6405
rect 39811 6364 39820 6404
rect 39860 6364 39869 6404
rect 39811 6363 39869 6364
rect 40483 6404 40541 6405
rect 40483 6364 40492 6404
rect 40532 6364 40541 6404
rect 40483 6363 40541 6364
rect 40867 6404 40925 6405
rect 40867 6364 40876 6404
rect 40916 6364 40925 6404
rect 40867 6363 40925 6364
rect 3147 6320 3189 6329
rect 3147 6280 3148 6320
rect 3188 6280 3189 6320
rect 3147 6271 3189 6280
rect 4579 6320 4637 6321
rect 4579 6280 4588 6320
rect 4628 6280 4637 6320
rect 4579 6279 4637 6280
rect 6499 6320 6557 6321
rect 6499 6280 6508 6320
rect 6548 6280 6557 6320
rect 6499 6279 6557 6280
rect 27915 6320 27957 6329
rect 27915 6280 27916 6320
rect 27956 6280 27957 6320
rect 27915 6271 27957 6280
rect 36363 6320 36405 6329
rect 36363 6280 36364 6320
rect 36404 6280 36405 6320
rect 36363 6271 36405 6280
rect 39627 6320 39669 6329
rect 39627 6280 39628 6320
rect 39668 6280 39669 6320
rect 39627 6271 39669 6280
rect 41067 6320 41109 6329
rect 41067 6280 41068 6320
rect 41108 6280 41109 6320
rect 41067 6271 41109 6280
rect 5355 6236 5397 6245
rect 5355 6196 5356 6236
rect 5396 6196 5397 6236
rect 5355 6187 5397 6196
rect 11307 6236 11349 6245
rect 11307 6196 11308 6236
rect 11348 6196 11349 6236
rect 11307 6187 11349 6196
rect 13707 6236 13749 6245
rect 13707 6196 13708 6236
rect 13748 6196 13749 6236
rect 13707 6187 13749 6196
rect 16203 6236 16245 6245
rect 16203 6196 16204 6236
rect 16244 6196 16245 6236
rect 16203 6187 16245 6196
rect 23499 6236 23541 6245
rect 23499 6196 23500 6236
rect 23540 6196 23541 6236
rect 23499 6187 23541 6196
rect 25803 6236 25845 6245
rect 25803 6196 25804 6236
rect 25844 6196 25845 6236
rect 25803 6187 25845 6196
rect 26091 6236 26133 6245
rect 26091 6196 26092 6236
rect 26132 6196 26133 6236
rect 26091 6187 26133 6196
rect 29739 6236 29781 6245
rect 29739 6196 29740 6236
rect 29780 6196 29781 6236
rect 29739 6187 29781 6196
rect 31947 6236 31989 6245
rect 31947 6196 31948 6236
rect 31988 6196 31989 6236
rect 31947 6187 31989 6196
rect 32139 6236 32181 6245
rect 32139 6196 32140 6236
rect 32180 6196 32181 6236
rect 32139 6187 32181 6196
rect 33963 6236 34005 6245
rect 33963 6196 33964 6236
rect 34004 6196 34005 6236
rect 33963 6187 34005 6196
rect 1152 6068 41856 6092
rect 1152 6028 3688 6068
rect 3728 6028 3770 6068
rect 3810 6028 3852 6068
rect 3892 6028 3934 6068
rect 3974 6028 4016 6068
rect 4056 6028 18808 6068
rect 18848 6028 18890 6068
rect 18930 6028 18972 6068
rect 19012 6028 19054 6068
rect 19094 6028 19136 6068
rect 19176 6028 33928 6068
rect 33968 6028 34010 6068
rect 34050 6028 34092 6068
rect 34132 6028 34174 6068
rect 34214 6028 34256 6068
rect 34296 6028 41856 6068
rect 1152 6004 41856 6028
rect 4107 5900 4149 5909
rect 4107 5860 4108 5900
rect 4148 5860 4149 5900
rect 4107 5851 4149 5860
rect 4875 5900 4917 5909
rect 4875 5860 4876 5900
rect 4916 5860 4917 5900
rect 4875 5851 4917 5860
rect 19467 5900 19509 5909
rect 19467 5860 19468 5900
rect 19508 5860 19509 5900
rect 19467 5851 19509 5860
rect 23499 5900 23541 5909
rect 23499 5860 23500 5900
rect 23540 5860 23541 5900
rect 23499 5851 23541 5860
rect 41067 5900 41109 5909
rect 41067 5860 41068 5900
rect 41108 5860 41109 5900
rect 41067 5851 41109 5860
rect 5355 5816 5397 5825
rect 5355 5776 5356 5816
rect 5396 5776 5397 5816
rect 5355 5767 5397 5776
rect 40683 5816 40725 5825
rect 40683 5776 40684 5816
rect 40724 5776 40725 5816
rect 40683 5767 40725 5776
rect 10539 5732 10581 5741
rect 10539 5692 10540 5732
rect 10580 5692 10581 5732
rect 10539 5683 10581 5692
rect 20227 5732 20285 5733
rect 20227 5692 20236 5732
rect 20276 5692 20285 5732
rect 20227 5691 20285 5692
rect 24459 5732 24501 5741
rect 24459 5692 24460 5732
rect 24500 5692 24501 5732
rect 26851 5732 26909 5733
rect 24459 5683 24501 5692
rect 25467 5690 25509 5699
rect 26851 5692 26860 5732
rect 26900 5692 26909 5732
rect 29731 5732 29789 5733
rect 26851 5691 26909 5692
rect 11595 5662 11637 5671
rect 1603 5648 1661 5649
rect 1603 5608 1612 5648
rect 1652 5608 1661 5648
rect 1603 5607 1661 5608
rect 2851 5648 2909 5649
rect 2851 5608 2860 5648
rect 2900 5608 2909 5648
rect 2851 5607 2909 5608
rect 4107 5648 4149 5657
rect 4107 5608 4108 5648
rect 4148 5608 4149 5648
rect 4107 5599 4149 5608
rect 4299 5648 4341 5657
rect 4299 5608 4300 5648
rect 4340 5608 4341 5648
rect 4299 5599 4341 5608
rect 4387 5648 4445 5649
rect 4387 5608 4396 5648
rect 4436 5608 4445 5648
rect 4387 5607 4445 5608
rect 4587 5648 4629 5657
rect 4587 5608 4588 5648
rect 4628 5608 4629 5648
rect 4587 5599 4629 5608
rect 4875 5648 4917 5657
rect 4875 5608 4876 5648
rect 4916 5608 4917 5648
rect 4875 5599 4917 5608
rect 5059 5648 5117 5649
rect 5059 5608 5068 5648
rect 5108 5608 5117 5648
rect 5059 5607 5117 5608
rect 5163 5648 5205 5657
rect 5163 5608 5164 5648
rect 5204 5608 5205 5648
rect 5163 5599 5205 5608
rect 5355 5648 5397 5657
rect 5355 5608 5356 5648
rect 5396 5608 5397 5648
rect 5355 5599 5397 5608
rect 5643 5648 5685 5657
rect 5643 5608 5644 5648
rect 5684 5608 5685 5648
rect 5643 5599 5685 5608
rect 5739 5648 5781 5657
rect 5739 5608 5740 5648
rect 5780 5608 5781 5648
rect 5739 5599 5781 5608
rect 6123 5648 6165 5657
rect 6123 5608 6124 5648
rect 6164 5608 6165 5648
rect 6123 5599 6165 5608
rect 6219 5648 6261 5657
rect 7179 5653 7221 5662
rect 6219 5608 6220 5648
rect 6260 5608 6261 5648
rect 6219 5599 6261 5608
rect 6691 5648 6749 5649
rect 6691 5608 6700 5648
rect 6740 5608 6749 5648
rect 6691 5607 6749 5608
rect 7179 5613 7180 5653
rect 7220 5613 7221 5653
rect 7179 5604 7221 5613
rect 8323 5648 8381 5649
rect 8323 5608 8332 5648
rect 8372 5608 8381 5648
rect 8323 5607 8381 5608
rect 9571 5648 9629 5649
rect 9571 5608 9580 5648
rect 9620 5608 9629 5648
rect 9571 5607 9629 5608
rect 10059 5648 10101 5657
rect 10059 5608 10060 5648
rect 10100 5608 10101 5648
rect 10059 5599 10101 5608
rect 10155 5648 10197 5657
rect 10155 5608 10156 5648
rect 10196 5608 10197 5648
rect 10155 5599 10197 5608
rect 10635 5648 10677 5657
rect 10635 5608 10636 5648
rect 10676 5608 10677 5648
rect 10635 5599 10677 5608
rect 11107 5648 11165 5649
rect 11107 5608 11116 5648
rect 11156 5608 11165 5648
rect 11595 5622 11596 5662
rect 11636 5622 11637 5662
rect 11595 5613 11637 5622
rect 13123 5648 13181 5649
rect 11107 5607 11165 5608
rect 13123 5608 13132 5648
rect 13172 5608 13181 5648
rect 13123 5607 13181 5608
rect 14371 5648 14429 5649
rect 14371 5608 14380 5648
rect 14420 5608 14429 5648
rect 14371 5607 14429 5608
rect 14755 5648 14813 5649
rect 14755 5608 14764 5648
rect 14804 5608 14813 5648
rect 14755 5607 14813 5608
rect 16003 5648 16061 5649
rect 16003 5608 16012 5648
rect 16052 5608 16061 5648
rect 16003 5607 16061 5608
rect 16387 5648 16445 5649
rect 16387 5608 16396 5648
rect 16436 5608 16445 5648
rect 16387 5607 16445 5608
rect 17635 5648 17693 5649
rect 17635 5608 17644 5648
rect 17684 5608 17693 5648
rect 17635 5607 17693 5608
rect 18019 5648 18077 5649
rect 18019 5608 18028 5648
rect 18068 5608 18077 5648
rect 18019 5607 18077 5608
rect 19267 5648 19325 5649
rect 19267 5608 19276 5648
rect 19316 5608 19325 5648
rect 19267 5607 19325 5608
rect 22051 5648 22109 5649
rect 22051 5608 22060 5648
rect 22100 5608 22109 5648
rect 22051 5607 22109 5608
rect 23299 5648 23357 5649
rect 23299 5608 23308 5648
rect 23348 5608 23357 5648
rect 23299 5607 23357 5608
rect 23883 5648 23925 5657
rect 23883 5608 23884 5648
rect 23924 5608 23925 5648
rect 23883 5599 23925 5608
rect 23979 5648 24021 5657
rect 23979 5608 23980 5648
rect 24020 5608 24021 5648
rect 23979 5599 24021 5608
rect 24363 5648 24405 5657
rect 25467 5650 25468 5690
rect 25508 5650 25509 5690
rect 29211 5690 29253 5699
rect 29731 5692 29740 5732
rect 29780 5692 29789 5732
rect 29731 5691 29789 5692
rect 35883 5732 35925 5741
rect 35883 5692 35884 5732
rect 35924 5692 35925 5732
rect 28694 5661 28736 5670
rect 24363 5608 24364 5648
rect 24404 5608 24405 5648
rect 24363 5599 24405 5608
rect 24931 5648 24989 5649
rect 24931 5608 24940 5648
rect 24980 5608 24989 5648
rect 25467 5641 25509 5650
rect 27627 5648 27669 5657
rect 24931 5607 24989 5608
rect 27627 5608 27628 5648
rect 27668 5608 27669 5648
rect 27627 5599 27669 5608
rect 27723 5648 27765 5657
rect 27723 5608 27724 5648
rect 27764 5608 27765 5648
rect 27723 5599 27765 5608
rect 28107 5648 28149 5657
rect 28107 5608 28108 5648
rect 28148 5608 28149 5648
rect 28107 5599 28149 5608
rect 28203 5648 28245 5657
rect 28203 5608 28204 5648
rect 28244 5608 28245 5648
rect 28694 5621 28695 5661
rect 28735 5621 28736 5661
rect 29211 5650 29212 5690
rect 29252 5650 29253 5690
rect 35883 5683 35925 5692
rect 40483 5732 40541 5733
rect 40483 5692 40492 5732
rect 40532 5692 40541 5732
rect 40483 5691 40541 5692
rect 40867 5732 40925 5733
rect 40867 5692 40876 5732
rect 40916 5692 40925 5732
rect 40867 5691 40925 5692
rect 33387 5662 33429 5671
rect 29211 5641 29253 5650
rect 30115 5648 30173 5649
rect 28694 5612 28736 5621
rect 28203 5599 28245 5608
rect 30115 5608 30124 5648
rect 30164 5608 30173 5648
rect 30115 5607 30173 5608
rect 31363 5648 31421 5649
rect 31363 5608 31372 5648
rect 31412 5608 31421 5648
rect 31363 5607 31421 5608
rect 31851 5648 31893 5657
rect 31851 5608 31852 5648
rect 31892 5608 31893 5648
rect 31851 5599 31893 5608
rect 31947 5648 31989 5657
rect 31947 5608 31948 5648
rect 31988 5608 31989 5648
rect 31947 5599 31989 5608
rect 32331 5648 32373 5657
rect 32331 5608 32332 5648
rect 32372 5608 32373 5648
rect 32331 5599 32373 5608
rect 32427 5648 32469 5657
rect 32427 5608 32428 5648
rect 32468 5608 32469 5648
rect 32427 5599 32469 5608
rect 32899 5648 32957 5649
rect 32899 5608 32908 5648
rect 32948 5608 32957 5648
rect 33387 5622 33388 5662
rect 33428 5622 33429 5662
rect 36891 5657 36933 5666
rect 33387 5613 33429 5622
rect 35307 5648 35349 5657
rect 32899 5607 32957 5608
rect 35307 5608 35308 5648
rect 35348 5608 35349 5648
rect 35307 5599 35349 5608
rect 35403 5648 35445 5657
rect 35403 5608 35404 5648
rect 35444 5608 35445 5648
rect 35403 5599 35445 5608
rect 35787 5648 35829 5657
rect 35787 5608 35788 5648
rect 35828 5608 35829 5648
rect 35787 5599 35829 5608
rect 36355 5648 36413 5649
rect 36355 5608 36364 5648
rect 36404 5608 36413 5648
rect 36891 5617 36892 5657
rect 36932 5617 36933 5657
rect 36891 5608 36933 5617
rect 36355 5607 36413 5608
rect 3051 5564 3093 5573
rect 3051 5524 3052 5564
rect 3092 5524 3093 5564
rect 3051 5515 3093 5524
rect 7371 5564 7413 5573
rect 7371 5524 7372 5564
rect 7412 5524 7413 5564
rect 7371 5515 7413 5524
rect 9771 5564 9813 5573
rect 9771 5524 9772 5564
rect 9812 5524 9813 5564
rect 9771 5515 9813 5524
rect 29355 5564 29397 5573
rect 29355 5524 29356 5564
rect 29396 5524 29397 5564
rect 29355 5515 29397 5524
rect 31563 5564 31605 5573
rect 31563 5524 31564 5564
rect 31604 5524 31605 5564
rect 31563 5515 31605 5524
rect 11787 5480 11829 5489
rect 11787 5440 11788 5480
rect 11828 5440 11829 5480
rect 11787 5431 11829 5440
rect 14571 5480 14613 5489
rect 14571 5440 14572 5480
rect 14612 5440 14613 5480
rect 14571 5431 14613 5440
rect 16203 5480 16245 5489
rect 16203 5440 16204 5480
rect 16244 5440 16245 5480
rect 16203 5431 16245 5440
rect 17835 5480 17877 5489
rect 17835 5440 17836 5480
rect 17876 5440 17877 5480
rect 17835 5431 17877 5440
rect 20427 5480 20469 5489
rect 20427 5440 20428 5480
rect 20468 5440 20469 5480
rect 20427 5431 20469 5440
rect 25611 5480 25653 5489
rect 25611 5440 25612 5480
rect 25652 5440 25653 5480
rect 25611 5431 25653 5440
rect 27051 5480 27093 5489
rect 27051 5440 27052 5480
rect 27092 5440 27093 5480
rect 27051 5431 27093 5440
rect 29547 5480 29589 5489
rect 29547 5440 29548 5480
rect 29588 5440 29589 5480
rect 29547 5431 29589 5440
rect 33579 5480 33621 5489
rect 33579 5440 33580 5480
rect 33620 5440 33621 5480
rect 33579 5431 33621 5440
rect 37035 5480 37077 5489
rect 37035 5440 37036 5480
rect 37076 5440 37077 5480
rect 37035 5431 37077 5440
rect 1152 5312 41856 5336
rect 1152 5272 4928 5312
rect 4968 5272 5010 5312
rect 5050 5272 5092 5312
rect 5132 5272 5174 5312
rect 5214 5272 5256 5312
rect 5296 5272 20048 5312
rect 20088 5272 20130 5312
rect 20170 5272 20212 5312
rect 20252 5272 20294 5312
rect 20334 5272 20376 5312
rect 20416 5272 35168 5312
rect 35208 5272 35250 5312
rect 35290 5272 35332 5312
rect 35372 5272 35414 5312
rect 35454 5272 35496 5312
rect 35536 5272 41856 5312
rect 1152 5248 41856 5272
rect 4195 5144 4253 5145
rect 4195 5104 4204 5144
rect 4244 5104 4253 5144
rect 4195 5103 4253 5104
rect 4587 5144 4629 5153
rect 4587 5104 4588 5144
rect 4628 5104 4629 5144
rect 4587 5095 4629 5104
rect 20523 5144 20565 5153
rect 20523 5104 20524 5144
rect 20564 5104 20565 5144
rect 20523 5095 20565 5104
rect 35595 5144 35637 5153
rect 35595 5104 35596 5144
rect 35636 5104 35637 5144
rect 35595 5095 35637 5104
rect 37323 5144 37365 5153
rect 37323 5104 37324 5144
rect 37364 5104 37365 5144
rect 37323 5095 37365 5104
rect 3627 5060 3669 5069
rect 3627 5020 3628 5060
rect 3668 5020 3669 5060
rect 3627 5011 3669 5020
rect 7275 5060 7317 5069
rect 7275 5020 7276 5060
rect 7316 5020 7317 5060
rect 7275 5011 7317 5020
rect 15627 5060 15669 5069
rect 15627 5020 15628 5060
rect 15668 5020 15669 5060
rect 15627 5011 15669 5020
rect 18507 5060 18549 5069
rect 18507 5020 18508 5060
rect 18548 5020 18549 5060
rect 18507 5011 18549 5020
rect 23115 5060 23157 5069
rect 23115 5020 23116 5060
rect 23156 5020 23157 5060
rect 23115 5011 23157 5020
rect 25131 5060 25173 5069
rect 25131 5020 25132 5060
rect 25172 5020 25173 5060
rect 25131 5011 25173 5020
rect 33675 5060 33717 5069
rect 33675 5020 33676 5060
rect 33716 5020 33717 5060
rect 33675 5011 33717 5020
rect 40011 5060 40053 5069
rect 40011 5020 40012 5060
rect 40052 5020 40053 5060
rect 40011 5011 40053 5020
rect 1603 4976 1661 4977
rect 1603 4936 1612 4976
rect 1652 4936 1661 4976
rect 1603 4935 1661 4936
rect 2851 4976 2909 4977
rect 2851 4936 2860 4976
rect 2900 4936 2909 4976
rect 2851 4935 2909 4936
rect 3723 4976 3765 4985
rect 3723 4936 3724 4976
rect 3764 4936 3765 4976
rect 3723 4927 3765 4936
rect 3819 4976 3861 4985
rect 3819 4936 3820 4976
rect 3860 4936 3861 4976
rect 3819 4927 3861 4936
rect 3915 4976 3957 4985
rect 3915 4936 3916 4976
rect 3956 4936 3957 4976
rect 3915 4927 3957 4936
rect 4107 4976 4149 4985
rect 4107 4936 4108 4976
rect 4148 4936 4149 4976
rect 4107 4927 4149 4936
rect 4299 4976 4341 4985
rect 4299 4936 4300 4976
rect 4340 4936 4341 4976
rect 4299 4927 4341 4936
rect 4387 4976 4445 4977
rect 4387 4936 4396 4976
rect 4436 4936 4445 4976
rect 4387 4935 4445 4936
rect 4675 4976 4733 4977
rect 4675 4936 4684 4976
rect 4724 4936 4733 4976
rect 4675 4935 4733 4936
rect 5067 4976 5109 4985
rect 5067 4936 5068 4976
rect 5108 4936 5109 4976
rect 5067 4927 5109 4936
rect 5251 4976 5309 4977
rect 5251 4936 5260 4976
rect 5300 4936 5309 4976
rect 5251 4935 5309 4936
rect 5547 4976 5589 4985
rect 5547 4936 5548 4976
rect 5588 4936 5589 4976
rect 5547 4927 5589 4936
rect 5643 4976 5685 4985
rect 5643 4936 5644 4976
rect 5684 4936 5685 4976
rect 5643 4927 5685 4936
rect 6123 4976 6165 4985
rect 6123 4936 6124 4976
rect 6164 4936 6165 4976
rect 6123 4927 6165 4936
rect 6595 4976 6653 4977
rect 6595 4936 6604 4976
rect 6644 4936 6653 4976
rect 8419 4976 8477 4977
rect 6595 4935 6653 4936
rect 7083 4966 7125 4975
rect 7083 4926 7084 4966
rect 7124 4926 7125 4966
rect 8419 4936 8428 4976
rect 8468 4936 8477 4976
rect 8419 4935 8477 4936
rect 8715 4976 8757 4985
rect 8715 4936 8716 4976
rect 8756 4936 8757 4976
rect 8715 4927 8757 4936
rect 8811 4976 8853 4985
rect 8811 4936 8812 4976
rect 8852 4936 8853 4976
rect 8811 4927 8853 4936
rect 9283 4976 9341 4977
rect 9283 4936 9292 4976
rect 9332 4936 9341 4976
rect 9283 4935 9341 4936
rect 10531 4976 10589 4977
rect 10531 4936 10540 4976
rect 10580 4936 10589 4976
rect 10531 4935 10589 4936
rect 11107 4976 11165 4977
rect 11107 4936 11116 4976
rect 11156 4936 11165 4976
rect 11107 4935 11165 4936
rect 12355 4976 12413 4977
rect 12355 4936 12364 4976
rect 12404 4936 12413 4976
rect 12355 4935 12413 4936
rect 13899 4976 13941 4985
rect 13899 4936 13900 4976
rect 13940 4936 13941 4976
rect 13899 4927 13941 4936
rect 13995 4976 14037 4985
rect 13995 4936 13996 4976
rect 14036 4936 14037 4976
rect 13995 4927 14037 4936
rect 14947 4976 15005 4977
rect 14947 4936 14956 4976
rect 14996 4936 15005 4976
rect 14947 4935 15005 4936
rect 15435 4971 15477 4980
rect 15435 4931 15436 4971
rect 15476 4931 15477 4971
rect 7083 4917 7125 4926
rect 15435 4922 15477 4931
rect 16779 4976 16821 4985
rect 16779 4936 16780 4976
rect 16820 4936 16821 4976
rect 16779 4927 16821 4936
rect 16875 4976 16917 4985
rect 16875 4936 16876 4976
rect 16916 4936 16917 4976
rect 16875 4927 16917 4936
rect 17827 4976 17885 4977
rect 17827 4936 17836 4976
rect 17876 4936 17885 4976
rect 17827 4935 17885 4936
rect 18315 4971 18357 4980
rect 18315 4931 18316 4971
rect 18356 4931 18357 4971
rect 18315 4922 18357 4931
rect 18795 4976 18837 4985
rect 18795 4936 18796 4976
rect 18836 4936 18837 4976
rect 18795 4927 18837 4936
rect 18891 4976 18933 4985
rect 18891 4936 18892 4976
rect 18932 4936 18933 4976
rect 18891 4927 18933 4936
rect 19843 4976 19901 4977
rect 19843 4936 19852 4976
rect 19892 4936 19901 4976
rect 21667 4976 21725 4977
rect 19843 4935 19901 4936
rect 20379 4934 20421 4943
rect 21667 4936 21676 4976
rect 21716 4936 21725 4976
rect 21667 4935 21725 4936
rect 22915 4976 22973 4977
rect 22915 4936 22924 4976
rect 22964 4936 22973 4976
rect 22915 4935 22973 4936
rect 23403 4976 23445 4985
rect 23403 4936 23404 4976
rect 23444 4936 23445 4976
rect 6027 4892 6069 4901
rect 6027 4852 6028 4892
rect 6068 4852 6069 4892
rect 6027 4843 6069 4852
rect 14379 4892 14421 4901
rect 14379 4852 14380 4892
rect 14420 4852 14421 4892
rect 14379 4843 14421 4852
rect 14475 4892 14517 4901
rect 14475 4852 14476 4892
rect 14516 4852 14517 4892
rect 14475 4843 14517 4852
rect 17259 4892 17301 4901
rect 17259 4852 17260 4892
rect 17300 4852 17301 4892
rect 17259 4843 17301 4852
rect 17355 4892 17397 4901
rect 17355 4852 17356 4892
rect 17396 4852 17397 4892
rect 17355 4843 17397 4852
rect 19275 4892 19317 4901
rect 19275 4852 19276 4892
rect 19316 4852 19317 4892
rect 19275 4843 19317 4852
rect 19371 4892 19413 4901
rect 19371 4852 19372 4892
rect 19412 4852 19413 4892
rect 20379 4894 20380 4934
rect 20420 4894 20421 4934
rect 23403 4927 23445 4936
rect 23499 4976 23541 4985
rect 23499 4936 23500 4976
rect 23540 4936 23541 4976
rect 23499 4927 23541 4936
rect 24451 4976 24509 4977
rect 24451 4936 24460 4976
rect 24500 4936 24509 4976
rect 26371 4976 26429 4977
rect 24451 4935 24509 4936
rect 24939 4962 24981 4971
rect 24939 4922 24940 4962
rect 24980 4922 24981 4962
rect 26371 4936 26380 4976
rect 26420 4936 26429 4976
rect 26371 4935 26429 4936
rect 27619 4976 27677 4977
rect 27619 4936 27628 4976
rect 27668 4936 27677 4976
rect 27619 4935 27677 4936
rect 29059 4976 29117 4977
rect 29059 4936 29068 4976
rect 29108 4936 29117 4976
rect 29059 4935 29117 4936
rect 30307 4976 30365 4977
rect 30307 4936 30316 4976
rect 30356 4936 30365 4976
rect 30307 4935 30365 4936
rect 31947 4976 31989 4985
rect 31947 4936 31948 4976
rect 31988 4936 31989 4976
rect 31947 4927 31989 4936
rect 32043 4976 32085 4985
rect 32043 4936 32044 4976
rect 32084 4936 32085 4976
rect 32043 4927 32085 4936
rect 32995 4976 33053 4977
rect 32995 4936 33004 4976
rect 33044 4936 33053 4976
rect 34147 4976 34205 4977
rect 32995 4935 33053 4936
rect 33483 4962 33525 4971
rect 24939 4913 24981 4922
rect 33483 4922 33484 4962
rect 33524 4922 33525 4962
rect 34147 4936 34156 4976
rect 34196 4936 34205 4976
rect 34147 4935 34205 4936
rect 35395 4976 35453 4977
rect 35395 4936 35404 4976
rect 35444 4936 35453 4976
rect 35395 4935 35453 4936
rect 35875 4976 35933 4977
rect 35875 4936 35884 4976
rect 35924 4936 35933 4976
rect 35875 4935 35933 4936
rect 37123 4976 37181 4977
rect 37123 4936 37132 4976
rect 37172 4936 37181 4976
rect 37123 4935 37181 4936
rect 38283 4976 38325 4985
rect 38283 4936 38284 4976
rect 38324 4936 38325 4976
rect 38283 4927 38325 4936
rect 38379 4976 38421 4985
rect 38379 4936 38380 4976
rect 38420 4936 38421 4976
rect 38379 4927 38421 4936
rect 38763 4976 38805 4985
rect 38763 4936 38764 4976
rect 38804 4936 38805 4976
rect 38763 4927 38805 4936
rect 39331 4976 39389 4977
rect 39331 4936 39340 4976
rect 39380 4936 39389 4976
rect 39331 4935 39389 4936
rect 39819 4962 39861 4971
rect 33483 4913 33525 4922
rect 39819 4922 39820 4962
rect 39860 4922 39861 4962
rect 39819 4913 39861 4922
rect 20379 4885 20421 4894
rect 20707 4892 20765 4893
rect 19371 4843 19413 4852
rect 20707 4852 20716 4892
rect 20756 4852 20765 4892
rect 20707 4851 20765 4852
rect 21091 4892 21149 4893
rect 21091 4852 21100 4892
rect 21140 4852 21149 4892
rect 21091 4851 21149 4852
rect 23883 4892 23925 4901
rect 23883 4852 23884 4892
rect 23924 4852 23925 4892
rect 23883 4843 23925 4852
rect 23979 4892 24021 4901
rect 23979 4852 23980 4892
rect 24020 4852 24021 4892
rect 23979 4843 24021 4852
rect 25507 4892 25565 4893
rect 25507 4852 25516 4892
rect 25556 4852 25565 4892
rect 25507 4851 25565 4852
rect 32427 4892 32469 4901
rect 32427 4852 32428 4892
rect 32468 4852 32469 4892
rect 32427 4843 32469 4852
rect 32523 4892 32565 4901
rect 32523 4852 32524 4892
rect 32564 4852 32565 4892
rect 32523 4843 32565 4852
rect 38859 4892 38901 4901
rect 38859 4852 38860 4892
rect 38900 4852 38901 4892
rect 38859 4843 38901 4852
rect 40483 4892 40541 4893
rect 40483 4852 40492 4892
rect 40532 4852 40541 4892
rect 40483 4851 40541 4852
rect 40867 4892 40925 4893
rect 40867 4852 40876 4892
rect 40916 4852 40925 4892
rect 40867 4851 40925 4852
rect 41251 4892 41309 4893
rect 41251 4852 41260 4892
rect 41300 4852 41309 4892
rect 41251 4851 41309 4852
rect 3051 4808 3093 4817
rect 3051 4768 3052 4808
rect 3092 4768 3093 4808
rect 3051 4759 3093 4768
rect 21291 4808 21333 4817
rect 21291 4768 21292 4808
rect 21332 4768 21333 4808
rect 21291 4759 21333 4768
rect 40683 4808 40725 4817
rect 40683 4768 40684 4808
rect 40724 4768 40725 4808
rect 40683 4759 40725 4768
rect 41067 4808 41109 4817
rect 41067 4768 41068 4808
rect 41108 4768 41109 4808
rect 41067 4759 41109 4768
rect 41451 4808 41493 4817
rect 41451 4768 41452 4808
rect 41492 4768 41493 4808
rect 41451 4759 41493 4768
rect 4587 4724 4629 4733
rect 4587 4684 4588 4724
rect 4628 4684 4629 4724
rect 4587 4675 4629 4684
rect 5163 4724 5205 4733
rect 5163 4684 5164 4724
rect 5204 4684 5205 4724
rect 5163 4675 5205 4684
rect 9091 4724 9149 4725
rect 9091 4684 9100 4724
rect 9140 4684 9149 4724
rect 9091 4683 9149 4684
rect 10731 4724 10773 4733
rect 10731 4684 10732 4724
rect 10772 4684 10773 4724
rect 10731 4675 10773 4684
rect 12555 4724 12597 4733
rect 12555 4684 12556 4724
rect 12596 4684 12597 4724
rect 12555 4675 12597 4684
rect 20907 4724 20949 4733
rect 20907 4684 20908 4724
rect 20948 4684 20949 4724
rect 20907 4675 20949 4684
rect 25323 4724 25365 4733
rect 25323 4684 25324 4724
rect 25364 4684 25365 4724
rect 25323 4675 25365 4684
rect 27819 4724 27861 4733
rect 27819 4684 27820 4724
rect 27860 4684 27861 4724
rect 27819 4675 27861 4684
rect 30507 4724 30549 4733
rect 30507 4684 30508 4724
rect 30548 4684 30549 4724
rect 30507 4675 30549 4684
rect 1152 4556 41856 4580
rect 1152 4516 3688 4556
rect 3728 4516 3770 4556
rect 3810 4516 3852 4556
rect 3892 4516 3934 4556
rect 3974 4516 4016 4556
rect 4056 4516 18808 4556
rect 18848 4516 18890 4556
rect 18930 4516 18972 4556
rect 19012 4516 19054 4556
rect 19094 4516 19136 4556
rect 19176 4516 33928 4556
rect 33968 4516 34010 4556
rect 34050 4516 34092 4556
rect 34132 4516 34174 4556
rect 34214 4516 34256 4556
rect 34296 4516 41856 4556
rect 1152 4492 41856 4516
rect 9483 4388 9525 4397
rect 9483 4348 9484 4388
rect 9524 4348 9525 4388
rect 9483 4339 9525 4348
rect 18795 4388 18837 4397
rect 18795 4348 18796 4388
rect 18836 4348 18837 4388
rect 18795 4339 18837 4348
rect 20715 4388 20757 4397
rect 20715 4348 20716 4388
rect 20756 4348 20757 4388
rect 20715 4339 20757 4348
rect 24267 4388 24309 4397
rect 24267 4348 24268 4388
rect 24308 4348 24309 4388
rect 24267 4339 24309 4348
rect 33387 4388 33429 4397
rect 33387 4348 33388 4388
rect 33428 4348 33429 4388
rect 33387 4339 33429 4348
rect 40299 4388 40341 4397
rect 40299 4348 40300 4388
rect 40340 4348 40341 4388
rect 40299 4339 40341 4348
rect 41067 4388 41109 4397
rect 41067 4348 41068 4388
rect 41108 4348 41109 4388
rect 41067 4339 41109 4348
rect 4195 4304 4253 4305
rect 4195 4264 4204 4304
rect 4244 4264 4253 4304
rect 4195 4263 4253 4264
rect 5067 4304 5109 4313
rect 5067 4264 5068 4304
rect 5108 4264 5109 4304
rect 5067 4255 5109 4264
rect 31267 4304 31325 4305
rect 31267 4264 31276 4304
rect 31316 4264 31325 4304
rect 31267 4263 31325 4264
rect 6219 4220 6261 4229
rect 6219 4180 6220 4220
rect 6260 4180 6261 4220
rect 6219 4171 6261 4180
rect 23203 4220 23261 4221
rect 23203 4180 23212 4220
rect 23252 4180 23261 4220
rect 23203 4179 23261 4180
rect 23491 4220 23549 4221
rect 23491 4180 23500 4220
rect 23540 4180 23549 4220
rect 23491 4179 23549 4180
rect 24067 4220 24125 4221
rect 24067 4180 24076 4220
rect 24116 4180 24125 4220
rect 24067 4179 24125 4180
rect 27043 4220 27101 4221
rect 27043 4180 27052 4220
rect 27092 4180 27101 4220
rect 27043 4179 27101 4180
rect 29635 4220 29693 4221
rect 29635 4180 29644 4220
rect 29684 4180 29693 4220
rect 29635 4179 29693 4180
rect 32803 4220 32861 4221
rect 32803 4180 32812 4220
rect 32852 4180 32861 4220
rect 32803 4179 32861 4180
rect 33187 4220 33245 4221
rect 33187 4180 33196 4220
rect 33236 4180 33245 4220
rect 33187 4179 33245 4180
rect 36835 4220 36893 4221
rect 36835 4180 36844 4220
rect 36884 4180 36893 4220
rect 36835 4179 36893 4180
rect 40483 4220 40541 4221
rect 40483 4180 40492 4220
rect 40532 4180 40541 4220
rect 40483 4179 40541 4180
rect 40867 4220 40925 4221
rect 40867 4180 40876 4220
rect 40916 4180 40925 4220
rect 40867 4179 40925 4180
rect 41251 4220 41309 4221
rect 41251 4180 41260 4220
rect 41300 4180 41309 4220
rect 41251 4179 41309 4180
rect 1507 4136 1565 4137
rect 1507 4096 1516 4136
rect 1556 4096 1565 4136
rect 1507 4095 1565 4096
rect 2755 4136 2813 4137
rect 2755 4096 2764 4136
rect 2804 4096 2813 4136
rect 2755 4095 2813 4096
rect 3523 4136 3581 4137
rect 3523 4096 3532 4136
rect 3572 4096 3581 4136
rect 3523 4095 3581 4096
rect 3819 4136 3861 4145
rect 3819 4096 3820 4136
rect 3860 4096 3861 4136
rect 3819 4087 3861 4096
rect 3915 4136 3957 4145
rect 3915 4096 3916 4136
rect 3956 4096 3957 4136
rect 3915 4087 3957 4096
rect 4395 4136 4437 4145
rect 4395 4096 4396 4136
rect 4436 4096 4437 4136
rect 4395 4087 4437 4096
rect 4587 4136 4629 4145
rect 4587 4096 4588 4136
rect 4628 4096 4629 4136
rect 4587 4087 4629 4096
rect 4675 4136 4733 4137
rect 4675 4096 4684 4136
rect 4724 4096 4733 4136
rect 4675 4095 4733 4096
rect 5067 4136 5109 4145
rect 5067 4096 5068 4136
rect 5108 4096 5109 4136
rect 5067 4087 5109 4096
rect 5643 4136 5685 4145
rect 5643 4096 5644 4136
rect 5684 4096 5685 4136
rect 5643 4087 5685 4096
rect 5739 4136 5781 4145
rect 5739 4096 5740 4136
rect 5780 4096 5781 4136
rect 5739 4087 5781 4096
rect 6123 4136 6165 4145
rect 7179 4141 7221 4150
rect 15579 4145 15621 4154
rect 6123 4096 6124 4136
rect 6164 4096 6165 4136
rect 6123 4087 6165 4096
rect 6691 4136 6749 4137
rect 6691 4096 6700 4136
rect 6740 4096 6749 4136
rect 6691 4095 6749 4096
rect 7179 4101 7180 4141
rect 7220 4101 7221 4141
rect 7179 4092 7221 4101
rect 8035 4136 8093 4137
rect 8035 4096 8044 4136
rect 8084 4096 8093 4136
rect 8035 4095 8093 4096
rect 9283 4136 9341 4137
rect 9283 4096 9292 4136
rect 9332 4096 9341 4136
rect 9283 4095 9341 4096
rect 10435 4136 10493 4137
rect 10435 4096 10444 4136
rect 10484 4096 10493 4136
rect 10435 4095 10493 4096
rect 11683 4136 11741 4137
rect 11683 4096 11692 4136
rect 11732 4096 11741 4136
rect 11683 4095 11741 4096
rect 12067 4136 12125 4137
rect 12067 4096 12076 4136
rect 12116 4096 12125 4136
rect 12067 4095 12125 4096
rect 13315 4136 13373 4137
rect 13315 4096 13324 4136
rect 13364 4096 13373 4136
rect 13315 4095 13373 4096
rect 13995 4136 14037 4145
rect 13995 4096 13996 4136
rect 14036 4096 14037 4136
rect 13995 4087 14037 4096
rect 14091 4136 14133 4145
rect 14091 4096 14092 4136
rect 14132 4096 14133 4136
rect 14091 4087 14133 4096
rect 14475 4136 14517 4145
rect 14475 4096 14476 4136
rect 14516 4096 14517 4136
rect 14475 4087 14517 4096
rect 14571 4136 14613 4145
rect 14571 4096 14572 4136
rect 14612 4096 14613 4136
rect 14571 4087 14613 4096
rect 15043 4136 15101 4137
rect 15043 4096 15052 4136
rect 15092 4096 15101 4136
rect 15579 4105 15580 4145
rect 15620 4105 15621 4145
rect 15579 4096 15621 4105
rect 17347 4136 17405 4137
rect 17347 4096 17356 4136
rect 17396 4096 17405 4136
rect 15043 4095 15101 4096
rect 17347 4095 17405 4096
rect 18595 4136 18653 4137
rect 18595 4096 18604 4136
rect 18644 4096 18653 4136
rect 18595 4095 18653 4096
rect 19267 4136 19325 4137
rect 19267 4096 19276 4136
rect 19316 4096 19325 4136
rect 19267 4095 19325 4096
rect 20515 4136 20573 4137
rect 20515 4096 20524 4136
rect 20564 4096 20573 4136
rect 20515 4095 20573 4096
rect 21099 4136 21141 4145
rect 21099 4096 21100 4136
rect 21140 4096 21141 4136
rect 21099 4087 21141 4096
rect 21195 4136 21237 4145
rect 21195 4096 21196 4136
rect 21236 4096 21237 4136
rect 21195 4087 21237 4096
rect 21579 4136 21621 4145
rect 21579 4096 21580 4136
rect 21620 4096 21621 4136
rect 21579 4087 21621 4096
rect 21675 4136 21717 4145
rect 22635 4141 22677 4150
rect 29115 4145 29157 4154
rect 21675 4096 21676 4136
rect 21716 4096 21717 4136
rect 21675 4087 21717 4096
rect 22147 4136 22205 4137
rect 22147 4096 22156 4136
rect 22196 4096 22205 4136
rect 22147 4095 22205 4096
rect 22635 4101 22636 4141
rect 22676 4101 22677 4141
rect 22635 4092 22677 4101
rect 24451 4136 24509 4137
rect 24451 4096 24460 4136
rect 24500 4096 24509 4136
rect 24451 4095 24509 4096
rect 25699 4136 25757 4137
rect 25699 4096 25708 4136
rect 25748 4096 25757 4136
rect 25699 4095 25757 4096
rect 27531 4136 27573 4145
rect 27531 4096 27532 4136
rect 27572 4096 27573 4136
rect 27531 4087 27573 4096
rect 27627 4136 27669 4145
rect 27627 4096 27628 4136
rect 27668 4096 27669 4136
rect 27627 4087 27669 4096
rect 28011 4136 28053 4145
rect 28011 4096 28012 4136
rect 28052 4096 28053 4136
rect 28011 4087 28053 4096
rect 28107 4136 28149 4145
rect 28107 4096 28108 4136
rect 28148 4096 28149 4136
rect 28107 4087 28149 4096
rect 28579 4136 28637 4137
rect 28579 4096 28588 4136
rect 28628 4096 28637 4136
rect 29115 4105 29116 4145
rect 29156 4105 29157 4145
rect 29115 4096 29157 4105
rect 30595 4136 30653 4137
rect 30595 4096 30604 4136
rect 30644 4096 30653 4136
rect 28579 4095 28637 4096
rect 30595 4095 30653 4096
rect 30891 4136 30933 4145
rect 30891 4096 30892 4136
rect 30932 4096 30933 4136
rect 30891 4087 30933 4096
rect 33571 4136 33629 4137
rect 33571 4096 33580 4136
rect 33620 4096 33629 4136
rect 33571 4095 33629 4096
rect 34819 4136 34877 4137
rect 34819 4096 34828 4136
rect 34868 4096 34877 4136
rect 34819 4095 34877 4096
rect 35011 4136 35069 4137
rect 35011 4096 35020 4136
rect 35060 4096 35069 4136
rect 35011 4095 35069 4096
rect 36259 4136 36317 4137
rect 36259 4096 36268 4136
rect 36308 4096 36317 4136
rect 36259 4095 36317 4096
rect 37219 4136 37277 4137
rect 37219 4096 37228 4136
rect 37268 4096 37277 4136
rect 37219 4095 37277 4096
rect 38467 4136 38525 4137
rect 38467 4096 38476 4136
rect 38516 4096 38525 4136
rect 38467 4095 38525 4096
rect 38851 4136 38909 4137
rect 38851 4096 38860 4136
rect 38900 4096 38909 4136
rect 38851 4095 38909 4096
rect 40099 4136 40157 4137
rect 40099 4096 40108 4136
rect 40148 4096 40157 4136
rect 40099 4095 40157 4096
rect 2955 4052 2997 4061
rect 2955 4012 2956 4052
rect 2996 4012 2997 4052
rect 2955 4003 2997 4012
rect 13515 4052 13557 4061
rect 13515 4012 13516 4052
rect 13556 4012 13557 4052
rect 13515 4003 13557 4012
rect 15723 4052 15765 4061
rect 15723 4012 15724 4052
rect 15764 4012 15765 4052
rect 15723 4003 15765 4012
rect 29259 4052 29301 4061
rect 29259 4012 29260 4052
rect 29300 4012 29301 4052
rect 29259 4003 29301 4012
rect 30987 4052 31029 4061
rect 30987 4012 30988 4052
rect 31028 4012 31029 4052
rect 30987 4003 31029 4012
rect 4483 3968 4541 3969
rect 4483 3928 4492 3968
rect 4532 3928 4541 3968
rect 4483 3927 4541 3928
rect 4875 3968 4917 3977
rect 4875 3928 4876 3968
rect 4916 3928 4917 3968
rect 4875 3919 4917 3928
rect 7371 3968 7413 3977
rect 7371 3928 7372 3968
rect 7412 3928 7413 3968
rect 7371 3919 7413 3928
rect 11883 3968 11925 3977
rect 11883 3928 11884 3968
rect 11924 3928 11925 3968
rect 11883 3919 11925 3928
rect 22827 3968 22869 3977
rect 22827 3928 22828 3968
rect 22868 3928 22869 3968
rect 22827 3919 22869 3928
rect 23019 3968 23061 3977
rect 23019 3928 23020 3968
rect 23060 3928 23061 3968
rect 23019 3919 23061 3928
rect 23691 3968 23733 3977
rect 23691 3928 23692 3968
rect 23732 3928 23733 3968
rect 23691 3919 23733 3928
rect 23883 3968 23925 3977
rect 23883 3928 23884 3968
rect 23924 3928 23925 3968
rect 23883 3919 23925 3928
rect 27243 3968 27285 3977
rect 27243 3928 27244 3968
rect 27284 3928 27285 3968
rect 27243 3919 27285 3928
rect 29451 3968 29493 3977
rect 29451 3928 29452 3968
rect 29492 3928 29493 3968
rect 29451 3919 29493 3928
rect 32619 3968 32661 3977
rect 32619 3928 32620 3968
rect 32660 3928 32661 3968
rect 32619 3919 32661 3928
rect 33003 3968 33045 3977
rect 33003 3928 33004 3968
rect 33044 3928 33045 3968
rect 33003 3919 33045 3928
rect 36459 3968 36501 3977
rect 36459 3928 36460 3968
rect 36500 3928 36501 3968
rect 36459 3919 36501 3928
rect 36651 3968 36693 3977
rect 36651 3928 36652 3968
rect 36692 3928 36693 3968
rect 36651 3919 36693 3928
rect 38667 3968 38709 3977
rect 38667 3928 38668 3968
rect 38708 3928 38709 3968
rect 38667 3919 38709 3928
rect 40683 3968 40725 3977
rect 40683 3928 40684 3968
rect 40724 3928 40725 3968
rect 40683 3919 40725 3928
rect 41451 3968 41493 3977
rect 41451 3928 41452 3968
rect 41492 3928 41493 3968
rect 41451 3919 41493 3928
rect 1152 3800 41856 3824
rect 1152 3760 4928 3800
rect 4968 3760 5010 3800
rect 5050 3760 5092 3800
rect 5132 3760 5174 3800
rect 5214 3760 5256 3800
rect 5296 3760 20048 3800
rect 20088 3760 20130 3800
rect 20170 3760 20212 3800
rect 20252 3760 20294 3800
rect 20334 3760 20376 3800
rect 20416 3760 35168 3800
rect 35208 3760 35250 3800
rect 35290 3760 35332 3800
rect 35372 3760 35414 3800
rect 35454 3760 35496 3800
rect 35536 3760 41856 3800
rect 1152 3736 41856 3760
rect 4003 3632 4061 3633
rect 4003 3592 4012 3632
rect 4052 3592 4061 3632
rect 4003 3591 4061 3592
rect 10155 3632 10197 3641
rect 10155 3592 10156 3632
rect 10196 3592 10197 3632
rect 10155 3583 10197 3592
rect 12843 3632 12885 3641
rect 12843 3592 12844 3632
rect 12884 3592 12885 3632
rect 12843 3583 12885 3592
rect 15627 3632 15669 3641
rect 15627 3592 15628 3632
rect 15668 3592 15669 3632
rect 15627 3583 15669 3592
rect 21099 3632 21141 3641
rect 21099 3592 21100 3632
rect 21140 3592 21141 3632
rect 21099 3583 21141 3592
rect 22827 3632 22869 3641
rect 22827 3592 22828 3632
rect 22868 3592 22869 3632
rect 22827 3583 22869 3592
rect 29547 3632 29589 3641
rect 29547 3592 29548 3632
rect 29588 3592 29589 3632
rect 29547 3583 29589 3592
rect 3339 3548 3381 3557
rect 3339 3508 3340 3548
rect 3380 3508 3381 3548
rect 3339 3499 3381 3508
rect 7275 3548 7317 3557
rect 7275 3508 7276 3548
rect 7316 3508 7317 3548
rect 7275 3499 7317 3508
rect 7755 3548 7797 3557
rect 7755 3508 7756 3548
rect 7796 3508 7797 3548
rect 7755 3499 7797 3508
rect 18027 3548 18069 3557
rect 18027 3508 18028 3548
rect 18068 3508 18069 3548
rect 18027 3499 18069 3508
rect 24651 3548 24693 3557
rect 24651 3508 24652 3548
rect 24692 3508 24693 3548
rect 24651 3499 24693 3508
rect 26667 3548 26709 3557
rect 26667 3508 26668 3548
rect 26708 3508 26709 3548
rect 26667 3499 26709 3508
rect 31467 3548 31509 3557
rect 31467 3508 31468 3548
rect 31508 3508 31509 3548
rect 31467 3499 31509 3508
rect 33483 3548 33525 3557
rect 33483 3508 33484 3548
rect 33524 3508 33525 3548
rect 33483 3499 33525 3508
rect 35883 3548 35925 3557
rect 35883 3508 35884 3548
rect 35924 3508 35925 3548
rect 35883 3499 35925 3508
rect 37899 3548 37941 3557
rect 37899 3508 37900 3548
rect 37940 3508 37941 3548
rect 37899 3499 37941 3508
rect 1603 3464 1661 3465
rect 1603 3424 1612 3464
rect 1652 3424 1661 3464
rect 1603 3423 1661 3424
rect 2851 3464 2909 3465
rect 2851 3424 2860 3464
rect 2900 3424 2909 3464
rect 3427 3464 3485 3465
rect 2851 3423 2909 3424
rect 3243 3449 3285 3458
rect 3243 3409 3244 3449
rect 3284 3409 3285 3449
rect 3427 3424 3436 3464
rect 3476 3424 3485 3464
rect 3427 3423 3485 3424
rect 3619 3464 3677 3465
rect 3619 3424 3628 3464
rect 3668 3424 3677 3464
rect 3619 3423 3677 3424
rect 3715 3464 3773 3465
rect 3715 3424 3724 3464
rect 3764 3424 3773 3464
rect 3715 3423 3773 3424
rect 3915 3464 3957 3473
rect 3915 3424 3916 3464
rect 3956 3424 3957 3464
rect 3915 3415 3957 3424
rect 4011 3464 4053 3473
rect 4011 3424 4012 3464
rect 4052 3424 4053 3464
rect 4011 3415 4053 3424
rect 4147 3464 4205 3465
rect 4147 3424 4156 3464
rect 4196 3424 4205 3464
rect 4147 3423 4205 3424
rect 4491 3464 4533 3473
rect 4491 3424 4492 3464
rect 4532 3424 4533 3464
rect 4491 3415 4533 3424
rect 4587 3464 4629 3473
rect 4587 3424 4588 3464
rect 4628 3424 4629 3464
rect 4587 3415 4629 3424
rect 4683 3464 4725 3473
rect 4683 3424 4684 3464
rect 4724 3424 4725 3464
rect 4683 3415 4725 3424
rect 4779 3464 4821 3473
rect 4779 3424 4780 3464
rect 4820 3424 4821 3464
rect 4779 3415 4821 3424
rect 4971 3464 5013 3473
rect 4971 3424 4972 3464
rect 5012 3424 5013 3464
rect 4971 3415 5013 3424
rect 5067 3464 5109 3473
rect 5067 3424 5068 3464
rect 5108 3424 5109 3464
rect 5067 3415 5109 3424
rect 5163 3464 5205 3473
rect 5163 3424 5164 3464
rect 5204 3424 5205 3464
rect 5163 3415 5205 3424
rect 5259 3464 5301 3473
rect 5259 3424 5260 3464
rect 5300 3424 5301 3464
rect 5259 3415 5301 3424
rect 5547 3464 5589 3473
rect 5547 3424 5548 3464
rect 5588 3424 5589 3464
rect 5547 3415 5589 3424
rect 5643 3464 5685 3473
rect 5643 3424 5644 3464
rect 5684 3424 5685 3464
rect 5643 3415 5685 3424
rect 6027 3464 6069 3473
rect 6027 3424 6028 3464
rect 6068 3424 6069 3464
rect 6027 3415 6069 3424
rect 6123 3464 6165 3473
rect 6123 3424 6124 3464
rect 6164 3424 6165 3464
rect 6123 3415 6165 3424
rect 6595 3464 6653 3465
rect 6595 3424 6604 3464
rect 6644 3424 6653 3464
rect 6595 3423 6653 3424
rect 7083 3459 7125 3468
rect 7083 3419 7084 3459
rect 7124 3419 7125 3459
rect 7083 3410 7125 3419
rect 7851 3464 7893 3473
rect 7851 3424 7852 3464
rect 7892 3424 7893 3464
rect 7851 3415 7893 3424
rect 8131 3464 8189 3465
rect 8131 3424 8140 3464
rect 8180 3424 8189 3464
rect 8131 3423 8189 3424
rect 8707 3464 8765 3465
rect 8707 3424 8716 3464
rect 8756 3424 8765 3464
rect 8707 3423 8765 3424
rect 9955 3464 10013 3465
rect 9955 3424 9964 3464
rect 10004 3424 10013 3464
rect 9955 3423 10013 3424
rect 11115 3464 11157 3473
rect 11115 3424 11116 3464
rect 11156 3424 11157 3464
rect 11115 3415 11157 3424
rect 11211 3464 11253 3473
rect 11211 3424 11212 3464
rect 11252 3424 11253 3464
rect 11211 3415 11253 3424
rect 12163 3464 12221 3465
rect 12163 3424 12172 3464
rect 12212 3424 12221 3464
rect 12163 3423 12221 3424
rect 12651 3459 12693 3468
rect 12651 3419 12652 3459
rect 12692 3419 12693 3459
rect 14179 3464 14237 3465
rect 14179 3424 14188 3464
rect 14228 3424 14237 3464
rect 14179 3423 14237 3424
rect 15427 3464 15485 3465
rect 15427 3424 15436 3464
rect 15476 3424 15485 3464
rect 15427 3423 15485 3424
rect 16299 3464 16341 3473
rect 16299 3424 16300 3464
rect 16340 3424 16341 3464
rect 12651 3410 12693 3419
rect 16299 3415 16341 3424
rect 16395 3464 16437 3473
rect 16395 3424 16396 3464
rect 16436 3424 16437 3464
rect 16395 3415 16437 3424
rect 16875 3464 16917 3473
rect 16875 3424 16876 3464
rect 16916 3424 16917 3464
rect 16875 3415 16917 3424
rect 17347 3464 17405 3465
rect 17347 3424 17356 3464
rect 17396 3424 17405 3464
rect 17347 3423 17405 3424
rect 17835 3459 17877 3468
rect 17835 3419 17836 3459
rect 17876 3419 17877 3459
rect 19651 3464 19709 3465
rect 19651 3424 19660 3464
rect 19700 3424 19709 3464
rect 19651 3423 19709 3424
rect 20899 3464 20957 3465
rect 20899 3424 20908 3464
rect 20948 3424 20957 3464
rect 20899 3423 20957 3424
rect 21379 3464 21437 3465
rect 21379 3424 21388 3464
rect 21428 3424 21437 3464
rect 21379 3423 21437 3424
rect 22627 3464 22685 3465
rect 22627 3424 22636 3464
rect 22676 3424 22685 3464
rect 22627 3423 22685 3424
rect 23203 3464 23261 3465
rect 23203 3424 23212 3464
rect 23252 3424 23261 3464
rect 23203 3423 23261 3424
rect 24451 3464 24509 3465
rect 24451 3424 24460 3464
rect 24500 3424 24509 3464
rect 24451 3423 24509 3424
rect 24939 3464 24981 3473
rect 24939 3424 24940 3464
rect 24980 3424 24981 3464
rect 17835 3410 17877 3419
rect 24939 3415 24981 3424
rect 25035 3464 25077 3473
rect 25035 3424 25036 3464
rect 25076 3424 25077 3464
rect 25035 3415 25077 3424
rect 25419 3464 25461 3473
rect 25419 3424 25420 3464
rect 25460 3424 25461 3464
rect 25419 3415 25461 3424
rect 25515 3464 25557 3473
rect 25515 3424 25516 3464
rect 25556 3424 25557 3464
rect 25515 3415 25557 3424
rect 25987 3464 26045 3465
rect 25987 3424 25996 3464
rect 26036 3424 26045 3464
rect 28099 3464 28157 3465
rect 25987 3423 26045 3424
rect 26475 3450 26517 3459
rect 26475 3410 26476 3450
rect 26516 3410 26517 3450
rect 28099 3424 28108 3464
rect 28148 3424 28157 3464
rect 28099 3423 28157 3424
rect 29347 3464 29405 3465
rect 29347 3424 29356 3464
rect 29396 3424 29405 3464
rect 29347 3423 29405 3424
rect 30019 3464 30077 3465
rect 30019 3424 30028 3464
rect 30068 3424 30077 3464
rect 30019 3423 30077 3424
rect 31267 3464 31325 3465
rect 31267 3424 31276 3464
rect 31316 3424 31325 3464
rect 31267 3423 31325 3424
rect 31755 3464 31797 3473
rect 31755 3424 31756 3464
rect 31796 3424 31797 3464
rect 31755 3415 31797 3424
rect 31851 3464 31893 3473
rect 31851 3424 31852 3464
rect 31892 3424 31893 3464
rect 31851 3415 31893 3424
rect 32803 3464 32861 3465
rect 32803 3424 32812 3464
rect 32852 3424 32861 3464
rect 34435 3464 34493 3465
rect 32803 3423 32861 3424
rect 33291 3450 33333 3459
rect 3243 3400 3285 3409
rect 26475 3401 26517 3410
rect 33291 3410 33292 3450
rect 33332 3410 33333 3450
rect 34435 3424 34444 3464
rect 34484 3424 34493 3464
rect 34435 3423 34493 3424
rect 35683 3464 35741 3465
rect 35683 3424 35692 3464
rect 35732 3424 35741 3464
rect 35683 3423 35741 3424
rect 36171 3464 36213 3473
rect 36171 3424 36172 3464
rect 36212 3424 36213 3464
rect 36171 3415 36213 3424
rect 36267 3464 36309 3473
rect 36267 3424 36268 3464
rect 36308 3424 36309 3464
rect 36267 3415 36309 3424
rect 36747 3464 36789 3473
rect 36747 3424 36748 3464
rect 36788 3424 36789 3464
rect 36747 3415 36789 3424
rect 37219 3464 37277 3465
rect 37219 3424 37228 3464
rect 37268 3424 37277 3464
rect 37219 3423 37277 3424
rect 37707 3459 37749 3468
rect 37707 3419 37708 3459
rect 37748 3419 37749 3459
rect 38275 3464 38333 3465
rect 38275 3424 38284 3464
rect 38324 3424 38333 3464
rect 38275 3423 38333 3424
rect 39523 3464 39581 3465
rect 39523 3424 39532 3464
rect 39572 3424 39581 3464
rect 39523 3423 39581 3424
rect 37707 3410 37749 3419
rect 33291 3401 33333 3410
rect 11595 3380 11637 3389
rect 11595 3340 11596 3380
rect 11636 3340 11637 3380
rect 11595 3331 11637 3340
rect 11691 3380 11733 3389
rect 11691 3340 11692 3380
rect 11732 3340 11733 3380
rect 11691 3331 11733 3340
rect 16779 3380 16821 3389
rect 16779 3340 16780 3380
rect 16820 3340 16821 3380
rect 16779 3331 16821 3340
rect 32235 3380 32277 3389
rect 32235 3340 32236 3380
rect 32276 3340 32277 3380
rect 32235 3331 32277 3340
rect 32331 3380 32373 3389
rect 32331 3340 32332 3380
rect 32372 3340 32373 3380
rect 32331 3331 32373 3340
rect 36651 3380 36693 3389
rect 36651 3340 36652 3380
rect 36692 3340 36693 3380
rect 36651 3331 36693 3340
rect 39907 3380 39965 3381
rect 39907 3340 39916 3380
rect 39956 3340 39965 3380
rect 39907 3339 39965 3340
rect 40099 3380 40157 3381
rect 40099 3340 40108 3380
rect 40148 3340 40157 3380
rect 40099 3339 40157 3340
rect 40483 3380 40541 3381
rect 40483 3340 40492 3380
rect 40532 3340 40541 3380
rect 40483 3339 40541 3340
rect 40867 3380 40925 3381
rect 40867 3340 40876 3380
rect 40916 3340 40925 3380
rect 40867 3339 40925 3340
rect 41251 3380 41309 3381
rect 41251 3340 41260 3380
rect 41300 3340 41309 3380
rect 41251 3339 41309 3340
rect 3051 3296 3093 3305
rect 3051 3256 3052 3296
rect 3092 3256 3093 3296
rect 3051 3247 3093 3256
rect 38091 3296 38133 3305
rect 38091 3256 38092 3296
rect 38132 3256 38133 3296
rect 38091 3247 38133 3256
rect 41067 3296 41109 3305
rect 41067 3256 41068 3296
rect 41108 3256 41109 3296
rect 41067 3247 41109 3256
rect 7459 3212 7517 3213
rect 7459 3172 7468 3212
rect 7508 3172 7517 3212
rect 7459 3171 7517 3172
rect 39723 3212 39765 3221
rect 39723 3172 39724 3212
rect 39764 3172 39765 3212
rect 39723 3163 39765 3172
rect 40299 3212 40341 3221
rect 40299 3172 40300 3212
rect 40340 3172 40341 3212
rect 40299 3163 40341 3172
rect 40683 3212 40725 3221
rect 40683 3172 40684 3212
rect 40724 3172 40725 3212
rect 40683 3163 40725 3172
rect 41451 3212 41493 3221
rect 41451 3172 41452 3212
rect 41492 3172 41493 3212
rect 41451 3163 41493 3172
rect 1152 3044 41856 3068
rect 1152 3004 3688 3044
rect 3728 3004 3770 3044
rect 3810 3004 3852 3044
rect 3892 3004 3934 3044
rect 3974 3004 4016 3044
rect 4056 3004 18808 3044
rect 18848 3004 18890 3044
rect 18930 3004 18972 3044
rect 19012 3004 19054 3044
rect 19094 3004 19136 3044
rect 19176 3004 33928 3044
rect 33968 3004 34010 3044
rect 34050 3004 34092 3044
rect 34132 3004 34174 3044
rect 34214 3004 34256 3044
rect 34296 3004 41856 3044
rect 1152 2980 41856 3004
rect 2955 2876 2997 2885
rect 2955 2836 2956 2876
rect 2996 2836 2997 2876
rect 2955 2827 2997 2836
rect 4875 2876 4917 2885
rect 4875 2836 4876 2876
rect 4916 2836 4917 2876
rect 4875 2827 4917 2836
rect 27147 2876 27189 2885
rect 27147 2836 27148 2876
rect 27188 2836 27189 2876
rect 27147 2827 27189 2836
rect 20323 2792 20381 2793
rect 20323 2752 20332 2792
rect 20372 2752 20381 2792
rect 20323 2751 20381 2752
rect 24451 2792 24509 2793
rect 24451 2752 24460 2792
rect 24500 2752 24509 2792
rect 24451 2751 24509 2752
rect 32907 2792 32949 2801
rect 32907 2752 32908 2792
rect 32948 2752 32949 2792
rect 32907 2743 32949 2752
rect 41067 2792 41109 2801
rect 41067 2752 41068 2792
rect 41108 2752 41109 2792
rect 41067 2743 41109 2752
rect 11499 2708 11541 2717
rect 11499 2668 11500 2708
rect 11540 2668 11541 2708
rect 11499 2659 11541 2668
rect 14475 2708 14517 2717
rect 14475 2668 14476 2708
rect 14516 2668 14517 2708
rect 14475 2659 14517 2668
rect 20707 2708 20765 2709
rect 20707 2668 20716 2708
rect 20756 2668 20765 2708
rect 20707 2667 20765 2668
rect 20899 2708 20957 2709
rect 20899 2668 20908 2708
rect 20948 2668 20957 2708
rect 20899 2667 20957 2668
rect 21475 2708 21533 2709
rect 21475 2668 21484 2708
rect 21524 2668 21533 2708
rect 21475 2667 21533 2668
rect 22147 2708 22205 2709
rect 22147 2668 22156 2708
rect 22196 2668 22205 2708
rect 22147 2667 22205 2668
rect 22915 2708 22973 2709
rect 22915 2668 22924 2708
rect 22964 2668 22973 2708
rect 22915 2667 22973 2668
rect 23299 2708 23357 2709
rect 23299 2668 23308 2708
rect 23348 2668 23357 2708
rect 23299 2667 23357 2668
rect 24643 2708 24701 2709
rect 24643 2668 24652 2708
rect 24692 2668 24701 2708
rect 24643 2667 24701 2668
rect 25315 2708 25373 2709
rect 25315 2668 25324 2708
rect 25364 2668 25373 2708
rect 25315 2667 25373 2668
rect 32707 2708 32765 2709
rect 32707 2668 32716 2708
rect 32756 2668 32765 2708
rect 32707 2667 32765 2668
rect 35779 2708 35837 2709
rect 35779 2668 35788 2708
rect 35828 2668 35837 2708
rect 35779 2667 35837 2668
rect 36555 2708 36597 2717
rect 36555 2668 36556 2708
rect 36596 2668 36597 2708
rect 36555 2659 36597 2668
rect 38179 2708 38237 2709
rect 38179 2668 38188 2708
rect 38228 2668 38237 2708
rect 38179 2667 38237 2668
rect 38563 2708 38621 2709
rect 38563 2668 38572 2708
rect 38612 2668 38621 2708
rect 38563 2667 38621 2668
rect 40867 2708 40925 2709
rect 40867 2668 40876 2708
rect 40916 2668 40925 2708
rect 40867 2667 40925 2668
rect 41251 2708 41309 2709
rect 41251 2668 41260 2708
rect 41300 2668 41309 2708
rect 41251 2667 41309 2668
rect 2755 2645 2813 2646
rect 1507 2624 1565 2625
rect 1507 2584 1516 2624
rect 1556 2584 1565 2624
rect 2755 2605 2764 2645
rect 2804 2605 2813 2645
rect 12459 2638 12501 2647
rect 2755 2604 2813 2605
rect 3243 2624 3285 2633
rect 1507 2583 1565 2584
rect 3243 2584 3244 2624
rect 3284 2584 3285 2624
rect 3243 2575 3285 2584
rect 3339 2624 3381 2633
rect 3339 2584 3340 2624
rect 3380 2584 3381 2624
rect 3339 2575 3381 2584
rect 3435 2624 3477 2633
rect 3435 2584 3436 2624
rect 3476 2584 3477 2624
rect 3435 2575 3477 2584
rect 3531 2624 3573 2633
rect 3531 2584 3532 2624
rect 3572 2584 3573 2624
rect 3531 2575 3573 2584
rect 3723 2624 3765 2633
rect 3723 2584 3724 2624
rect 3764 2584 3765 2624
rect 3723 2575 3765 2584
rect 3819 2624 3861 2633
rect 3819 2584 3820 2624
rect 3860 2584 3861 2624
rect 3819 2575 3861 2584
rect 4203 2624 4245 2633
rect 4203 2584 4204 2624
rect 4244 2584 4245 2624
rect 4203 2575 4245 2584
rect 4299 2624 4341 2633
rect 4299 2584 4300 2624
rect 4340 2584 4341 2624
rect 4299 2575 4341 2584
rect 4875 2624 4917 2633
rect 4875 2584 4876 2624
rect 4916 2584 4917 2624
rect 4875 2575 4917 2584
rect 5163 2624 5205 2633
rect 5163 2584 5164 2624
rect 5204 2584 5205 2624
rect 5163 2575 5205 2584
rect 5923 2624 5981 2625
rect 5923 2584 5932 2624
rect 5972 2584 5981 2624
rect 5923 2583 5981 2584
rect 7171 2624 7229 2625
rect 7171 2584 7180 2624
rect 7220 2584 7229 2624
rect 7171 2583 7229 2584
rect 7555 2624 7613 2625
rect 7555 2584 7564 2624
rect 7604 2584 7613 2624
rect 7555 2583 7613 2584
rect 8803 2624 8861 2625
rect 8803 2584 8812 2624
rect 8852 2584 8861 2624
rect 8803 2583 8861 2584
rect 9187 2624 9245 2625
rect 9187 2584 9196 2624
rect 9236 2584 9245 2624
rect 9187 2583 9245 2584
rect 10435 2624 10493 2625
rect 10435 2584 10444 2624
rect 10484 2584 10493 2624
rect 10435 2583 10493 2584
rect 10923 2624 10965 2633
rect 10923 2584 10924 2624
rect 10964 2584 10965 2624
rect 10923 2575 10965 2584
rect 11019 2624 11061 2633
rect 11019 2584 11020 2624
rect 11060 2584 11061 2624
rect 11019 2575 11061 2584
rect 11403 2624 11445 2633
rect 11403 2584 11404 2624
rect 11444 2584 11445 2624
rect 11403 2575 11445 2584
rect 11971 2624 12029 2625
rect 11971 2584 11980 2624
rect 12020 2584 12029 2624
rect 12459 2598 12460 2638
rect 12500 2598 12501 2638
rect 12459 2589 12501 2598
rect 13899 2624 13941 2633
rect 11971 2583 12029 2584
rect 13899 2584 13900 2624
rect 13940 2584 13941 2624
rect 13899 2575 13941 2584
rect 13995 2624 14037 2633
rect 13995 2584 13996 2624
rect 14036 2584 14037 2624
rect 13995 2575 14037 2584
rect 14379 2624 14421 2633
rect 15435 2629 15477 2638
rect 14379 2584 14380 2624
rect 14420 2584 14421 2624
rect 14379 2575 14421 2584
rect 14947 2624 15005 2625
rect 14947 2584 14956 2624
rect 14996 2584 15005 2624
rect 14947 2583 15005 2584
rect 15435 2589 15436 2629
rect 15476 2589 15477 2629
rect 15435 2580 15477 2589
rect 15907 2624 15965 2625
rect 15907 2584 15916 2624
rect 15956 2584 15965 2624
rect 15907 2583 15965 2584
rect 17155 2624 17213 2625
rect 17155 2584 17164 2624
rect 17204 2584 17213 2624
rect 17155 2583 17213 2584
rect 17923 2624 17981 2625
rect 17923 2584 17932 2624
rect 17972 2584 17981 2624
rect 17923 2583 17981 2584
rect 19171 2624 19229 2625
rect 19171 2584 19180 2624
rect 19220 2584 19229 2624
rect 19171 2583 19229 2584
rect 19651 2624 19709 2625
rect 19651 2584 19660 2624
rect 19700 2584 19709 2624
rect 19651 2583 19709 2584
rect 19947 2624 19989 2633
rect 19947 2584 19948 2624
rect 19988 2584 19989 2624
rect 19947 2575 19989 2584
rect 23779 2624 23837 2625
rect 23779 2584 23788 2624
rect 23828 2584 23837 2624
rect 23779 2583 23837 2584
rect 24075 2624 24117 2633
rect 24075 2584 24076 2624
rect 24116 2584 24117 2624
rect 24075 2575 24117 2584
rect 24171 2624 24213 2633
rect 24171 2584 24172 2624
rect 24212 2584 24213 2624
rect 24171 2575 24213 2584
rect 25699 2624 25757 2625
rect 25699 2584 25708 2624
rect 25748 2584 25757 2624
rect 25699 2583 25757 2584
rect 26947 2624 27005 2625
rect 26947 2584 26956 2624
rect 26996 2584 27005 2624
rect 26947 2583 27005 2584
rect 27523 2624 27581 2625
rect 27523 2584 27532 2624
rect 27572 2584 27581 2624
rect 27523 2583 27581 2584
rect 28771 2624 28829 2625
rect 28771 2584 28780 2624
rect 28820 2584 28829 2624
rect 28771 2583 28829 2584
rect 29155 2624 29213 2625
rect 29155 2584 29164 2624
rect 29204 2584 29213 2624
rect 29155 2583 29213 2584
rect 30403 2624 30461 2625
rect 30403 2584 30412 2624
rect 30452 2584 30461 2624
rect 30403 2583 30461 2584
rect 30787 2624 30845 2625
rect 30787 2584 30796 2624
rect 30836 2584 30845 2624
rect 30787 2583 30845 2584
rect 32035 2624 32093 2625
rect 32035 2584 32044 2624
rect 32084 2584 32093 2624
rect 32035 2583 32093 2584
rect 33091 2624 33149 2625
rect 33091 2584 33100 2624
rect 33140 2584 33149 2624
rect 33091 2583 33149 2584
rect 34339 2624 34397 2625
rect 34339 2584 34348 2624
rect 34388 2584 34397 2624
rect 34339 2583 34397 2584
rect 36075 2624 36117 2633
rect 36075 2584 36076 2624
rect 36116 2584 36117 2624
rect 36075 2575 36117 2584
rect 36171 2624 36213 2633
rect 36171 2584 36172 2624
rect 36212 2584 36213 2624
rect 36171 2575 36213 2584
rect 36651 2624 36693 2633
rect 37611 2629 37653 2638
rect 36651 2584 36652 2624
rect 36692 2584 36693 2624
rect 36651 2575 36693 2584
rect 37123 2624 37181 2625
rect 37123 2584 37132 2624
rect 37172 2584 37181 2624
rect 37123 2583 37181 2584
rect 37611 2589 37612 2629
rect 37652 2589 37653 2629
rect 37611 2580 37653 2589
rect 39139 2624 39197 2625
rect 39139 2584 39148 2624
rect 39188 2584 39197 2624
rect 39139 2583 39197 2584
rect 40387 2624 40445 2625
rect 40387 2584 40396 2624
rect 40436 2584 40445 2624
rect 40387 2583 40445 2584
rect 15627 2540 15669 2549
rect 15627 2500 15628 2540
rect 15668 2500 15669 2540
rect 15627 2491 15669 2500
rect 19371 2540 19413 2549
rect 19371 2500 19372 2540
rect 19412 2500 19413 2540
rect 19371 2491 19413 2500
rect 20043 2540 20085 2549
rect 20043 2500 20044 2540
rect 20084 2500 20085 2540
rect 20043 2491 20085 2500
rect 37803 2540 37845 2549
rect 37803 2500 37804 2540
rect 37844 2500 37845 2540
rect 37803 2491 37845 2500
rect 38955 2540 38997 2549
rect 38955 2500 38956 2540
rect 38996 2500 38997 2540
rect 38955 2491 38997 2500
rect 4003 2456 4061 2457
rect 4003 2416 4012 2456
rect 4052 2416 4061 2456
rect 4003 2415 4061 2416
rect 4483 2456 4541 2457
rect 4483 2416 4492 2456
rect 4532 2416 4541 2456
rect 4483 2415 4541 2416
rect 7371 2456 7413 2465
rect 7371 2416 7372 2456
rect 7412 2416 7413 2456
rect 7371 2407 7413 2416
rect 9003 2456 9045 2465
rect 9003 2416 9004 2456
rect 9044 2416 9045 2456
rect 9003 2407 9045 2416
rect 10635 2456 10677 2465
rect 10635 2416 10636 2456
rect 10676 2416 10677 2456
rect 10635 2407 10677 2416
rect 12651 2456 12693 2465
rect 12651 2416 12652 2456
rect 12692 2416 12693 2456
rect 12651 2407 12693 2416
rect 17355 2456 17397 2465
rect 17355 2416 17356 2456
rect 17396 2416 17397 2456
rect 17355 2407 17397 2416
rect 20523 2456 20565 2465
rect 20523 2416 20524 2456
rect 20564 2416 20565 2456
rect 20523 2407 20565 2416
rect 21099 2456 21141 2465
rect 21099 2416 21100 2456
rect 21140 2416 21141 2456
rect 21099 2407 21141 2416
rect 21675 2456 21717 2465
rect 21675 2416 21676 2456
rect 21716 2416 21717 2456
rect 21675 2407 21717 2416
rect 21963 2456 22005 2465
rect 21963 2416 21964 2456
rect 22004 2416 22005 2456
rect 21963 2407 22005 2416
rect 23115 2456 23157 2465
rect 23115 2416 23116 2456
rect 23156 2416 23157 2456
rect 23115 2407 23157 2416
rect 23499 2456 23541 2465
rect 23499 2416 23500 2456
rect 23540 2416 23541 2456
rect 23499 2407 23541 2416
rect 24843 2456 24885 2465
rect 24843 2416 24844 2456
rect 24884 2416 24885 2456
rect 24843 2407 24885 2416
rect 25515 2456 25557 2465
rect 25515 2416 25516 2456
rect 25556 2416 25557 2456
rect 25515 2407 25557 2416
rect 27339 2456 27381 2465
rect 27339 2416 27340 2456
rect 27380 2416 27381 2456
rect 27339 2407 27381 2416
rect 28971 2456 29013 2465
rect 28971 2416 28972 2456
rect 29012 2416 29013 2456
rect 28971 2407 29013 2416
rect 30603 2456 30645 2465
rect 30603 2416 30604 2456
rect 30644 2416 30645 2456
rect 30603 2407 30645 2416
rect 32523 2456 32565 2465
rect 32523 2416 32524 2456
rect 32564 2416 32565 2456
rect 32523 2407 32565 2416
rect 35595 2456 35637 2465
rect 35595 2416 35596 2456
rect 35636 2416 35637 2456
rect 35595 2407 35637 2416
rect 37995 2456 38037 2465
rect 37995 2416 37996 2456
rect 38036 2416 38037 2456
rect 37995 2407 38037 2416
rect 38763 2456 38805 2465
rect 38763 2416 38764 2456
rect 38804 2416 38805 2456
rect 38763 2407 38805 2416
rect 41451 2456 41493 2465
rect 41451 2416 41452 2456
rect 41492 2416 41493 2456
rect 41451 2407 41493 2416
rect 1152 2288 41856 2312
rect 1152 2248 4928 2288
rect 4968 2248 5010 2288
rect 5050 2248 5092 2288
rect 5132 2248 5174 2288
rect 5214 2248 5256 2288
rect 5296 2248 20048 2288
rect 20088 2248 20130 2288
rect 20170 2248 20212 2288
rect 20252 2248 20294 2288
rect 20334 2248 20376 2288
rect 20416 2248 35168 2288
rect 35208 2248 35250 2288
rect 35290 2248 35332 2288
rect 35372 2248 35414 2288
rect 35454 2248 35496 2288
rect 35536 2248 41856 2288
rect 1152 2224 41856 2248
rect 14859 2120 14901 2129
rect 14859 2080 14860 2120
rect 14900 2080 14901 2120
rect 14859 2071 14901 2080
rect 16875 2120 16917 2129
rect 16875 2080 16876 2120
rect 16916 2080 16917 2120
rect 16875 2071 16917 2080
rect 19179 2120 19221 2129
rect 19179 2080 19180 2120
rect 19220 2080 19221 2120
rect 19179 2071 19221 2080
rect 22059 2120 22101 2129
rect 22059 2080 22060 2120
rect 22100 2080 22101 2120
rect 22059 2071 22101 2080
rect 37035 2120 37077 2129
rect 37035 2080 37036 2120
rect 37076 2080 37077 2120
rect 37035 2071 37077 2080
rect 40203 2120 40245 2129
rect 40203 2080 40204 2120
rect 40244 2080 40245 2120
rect 40203 2071 40245 2080
rect 5259 2036 5301 2045
rect 5259 1996 5260 2036
rect 5300 1996 5301 2036
rect 5259 1987 5301 1996
rect 7275 2036 7317 2045
rect 7275 1996 7276 2036
rect 7316 1996 7317 2036
rect 7275 1987 7317 1996
rect 9579 2036 9621 2045
rect 9579 1996 9580 2036
rect 9620 1996 9621 2036
rect 9579 1987 9621 1996
rect 12843 2036 12885 2045
rect 12843 1996 12844 2036
rect 12884 1996 12885 2036
rect 12843 1987 12885 1996
rect 23883 2036 23925 2045
rect 23883 1996 23884 2036
rect 23924 1996 23925 2036
rect 23883 1987 23925 1996
rect 26475 2036 26517 2045
rect 26475 1996 26476 2036
rect 26516 1996 26517 2036
rect 26475 1987 26517 1996
rect 29451 2036 29493 2045
rect 29451 1996 29452 2036
rect 29492 1996 29493 2036
rect 29451 1987 29493 1996
rect 32235 2036 32277 2045
rect 32235 1996 32236 2036
rect 32276 1996 32277 2036
rect 32235 1987 32277 1996
rect 40011 2036 40053 2045
rect 40011 1996 40012 2036
rect 40052 1996 40053 2036
rect 40011 1987 40053 1996
rect 2179 1952 2237 1953
rect 2179 1912 2188 1952
rect 2228 1912 2237 1952
rect 2179 1911 2237 1912
rect 3427 1952 3485 1953
rect 3427 1912 3436 1952
rect 3476 1912 3485 1952
rect 3427 1911 3485 1912
rect 3811 1952 3869 1953
rect 3811 1912 3820 1952
rect 3860 1912 3869 1952
rect 3811 1911 3869 1912
rect 5059 1952 5117 1953
rect 5059 1912 5068 1952
rect 5108 1912 5117 1952
rect 5059 1911 5117 1912
rect 5547 1952 5589 1961
rect 5547 1912 5548 1952
rect 5588 1912 5589 1952
rect 5547 1903 5589 1912
rect 5643 1952 5685 1961
rect 5643 1912 5644 1952
rect 5684 1912 5685 1952
rect 5643 1903 5685 1912
rect 6027 1952 6069 1961
rect 6027 1912 6028 1952
rect 6068 1912 6069 1952
rect 6027 1903 6069 1912
rect 6595 1952 6653 1953
rect 6595 1912 6604 1952
rect 6644 1912 6653 1952
rect 6595 1911 6653 1912
rect 7083 1947 7125 1956
rect 7083 1907 7084 1947
rect 7124 1907 7125 1947
rect 7083 1898 7125 1907
rect 7851 1952 7893 1961
rect 7851 1912 7852 1952
rect 7892 1912 7893 1952
rect 7851 1903 7893 1912
rect 7947 1952 7989 1961
rect 7947 1912 7948 1952
rect 7988 1912 7989 1952
rect 7947 1903 7989 1912
rect 8331 1952 8373 1961
rect 8331 1912 8332 1952
rect 8372 1912 8373 1952
rect 8331 1903 8373 1912
rect 8899 1952 8957 1953
rect 8899 1912 8908 1952
rect 8948 1912 8957 1952
rect 8899 1911 8957 1912
rect 9387 1947 9429 1956
rect 9387 1907 9388 1947
rect 9428 1907 9429 1947
rect 9387 1898 9429 1907
rect 11115 1952 11157 1961
rect 11115 1912 11116 1952
rect 11156 1912 11157 1952
rect 11115 1903 11157 1912
rect 11211 1952 11253 1961
rect 11211 1912 11212 1952
rect 11252 1912 11253 1952
rect 11211 1903 11253 1912
rect 12163 1952 12221 1953
rect 12163 1912 12172 1952
rect 12212 1912 12221 1952
rect 12163 1911 12221 1912
rect 12651 1947 12693 1956
rect 12651 1907 12652 1947
rect 12692 1907 12693 1947
rect 13411 1952 13469 1953
rect 13411 1912 13420 1952
rect 13460 1912 13469 1952
rect 13411 1911 13469 1912
rect 14659 1952 14717 1953
rect 14659 1912 14668 1952
rect 14708 1912 14717 1952
rect 14659 1911 14717 1912
rect 15147 1952 15189 1961
rect 15147 1912 15148 1952
rect 15188 1912 15189 1952
rect 12651 1898 12693 1907
rect 15147 1903 15189 1912
rect 15243 1952 15285 1961
rect 15243 1912 15244 1952
rect 15284 1912 15285 1952
rect 15243 1903 15285 1912
rect 16195 1952 16253 1953
rect 16195 1912 16204 1952
rect 16244 1912 16253 1952
rect 17451 1952 17493 1961
rect 16195 1911 16253 1912
rect 16683 1938 16725 1947
rect 16683 1898 16684 1938
rect 16724 1898 16725 1938
rect 17451 1912 17452 1952
rect 17492 1912 17493 1952
rect 17451 1903 17493 1912
rect 17547 1952 17589 1961
rect 17547 1912 17548 1952
rect 17588 1912 17589 1952
rect 17547 1903 17589 1912
rect 18499 1952 18557 1953
rect 18499 1912 18508 1952
rect 18548 1912 18557 1952
rect 20331 1952 20373 1961
rect 18499 1911 18557 1912
rect 18987 1938 19029 1947
rect 16683 1889 16725 1898
rect 18987 1898 18988 1938
rect 19028 1898 19029 1938
rect 20331 1912 20332 1952
rect 20372 1912 20373 1952
rect 20331 1903 20373 1912
rect 20427 1952 20469 1961
rect 20427 1912 20428 1952
rect 20468 1912 20469 1952
rect 20427 1903 20469 1912
rect 21379 1952 21437 1953
rect 21379 1912 21388 1952
rect 21428 1912 21437 1952
rect 22435 1952 22493 1953
rect 21379 1911 21437 1912
rect 21867 1938 21909 1947
rect 18987 1889 19029 1898
rect 21867 1898 21868 1938
rect 21908 1898 21909 1938
rect 22435 1912 22444 1952
rect 22484 1912 22493 1952
rect 22435 1911 22493 1912
rect 23683 1952 23741 1953
rect 23683 1912 23692 1952
rect 23732 1912 23741 1952
rect 23683 1911 23741 1912
rect 24747 1952 24789 1961
rect 24747 1912 24748 1952
rect 24788 1912 24789 1952
rect 24747 1903 24789 1912
rect 24843 1952 24885 1961
rect 24843 1912 24844 1952
rect 24884 1912 24885 1952
rect 24843 1903 24885 1912
rect 25323 1952 25365 1961
rect 25323 1912 25324 1952
rect 25364 1912 25365 1952
rect 25323 1903 25365 1912
rect 25795 1952 25853 1953
rect 25795 1912 25804 1952
rect 25844 1912 25853 1952
rect 27723 1952 27765 1961
rect 25795 1911 25853 1912
rect 26283 1938 26325 1947
rect 21867 1889 21909 1898
rect 26283 1898 26284 1938
rect 26324 1898 26325 1938
rect 27723 1912 27724 1952
rect 27764 1912 27765 1952
rect 27723 1903 27765 1912
rect 27819 1952 27861 1961
rect 27819 1912 27820 1952
rect 27860 1912 27861 1952
rect 27819 1903 27861 1912
rect 28771 1952 28829 1953
rect 28771 1912 28780 1952
rect 28820 1912 28829 1952
rect 28771 1911 28829 1912
rect 29259 1947 29301 1956
rect 29259 1907 29260 1947
rect 29300 1907 29301 1947
rect 31083 1952 31125 1961
rect 29259 1898 29301 1907
rect 30507 1933 30549 1942
rect 26283 1889 26325 1898
rect 30507 1893 30508 1933
rect 30548 1893 30549 1933
rect 30507 1884 30549 1893
rect 30603 1933 30645 1942
rect 30603 1893 30604 1933
rect 30644 1893 30645 1933
rect 31083 1912 31084 1952
rect 31124 1912 31125 1952
rect 31083 1903 31125 1912
rect 31555 1952 31613 1953
rect 31555 1912 31564 1952
rect 31604 1912 31613 1952
rect 32995 1952 33053 1953
rect 31555 1911 31613 1912
rect 32043 1938 32085 1947
rect 30603 1884 30645 1893
rect 32043 1898 32044 1938
rect 32084 1898 32085 1938
rect 32995 1912 33004 1952
rect 33044 1912 33053 1952
rect 32995 1911 33053 1912
rect 34243 1952 34301 1953
rect 34243 1912 34252 1952
rect 34292 1912 34301 1952
rect 34243 1911 34301 1912
rect 35307 1952 35349 1961
rect 35307 1912 35308 1952
rect 35348 1912 35349 1952
rect 35307 1903 35349 1912
rect 35403 1952 35445 1961
rect 35403 1912 35404 1952
rect 35444 1912 35445 1952
rect 35403 1903 35445 1912
rect 35787 1952 35829 1961
rect 35787 1912 35788 1952
rect 35828 1912 35829 1952
rect 35787 1903 35829 1912
rect 36355 1952 36413 1953
rect 36355 1912 36364 1952
rect 36404 1912 36413 1952
rect 38283 1952 38325 1961
rect 36355 1911 36413 1912
rect 36843 1938 36885 1947
rect 32043 1889 32085 1898
rect 36843 1898 36844 1938
rect 36884 1898 36885 1938
rect 38283 1912 38284 1952
rect 38324 1912 38325 1952
rect 38283 1903 38325 1912
rect 38379 1952 38421 1961
rect 38379 1912 38380 1952
rect 38420 1912 38421 1952
rect 38379 1903 38421 1912
rect 38763 1952 38805 1961
rect 38763 1912 38764 1952
rect 38804 1912 38805 1952
rect 38763 1903 38805 1912
rect 38859 1952 38901 1961
rect 38859 1912 38860 1952
rect 38900 1912 38901 1952
rect 38859 1903 38901 1912
rect 39331 1952 39389 1953
rect 39331 1912 39340 1952
rect 39380 1912 39389 1952
rect 40387 1952 40445 1953
rect 39331 1911 39389 1912
rect 39819 1942 39861 1951
rect 36843 1889 36885 1898
rect 39819 1902 39820 1942
rect 39860 1902 39861 1942
rect 40387 1912 40396 1952
rect 40436 1912 40445 1952
rect 40387 1911 40445 1912
rect 41635 1952 41693 1953
rect 41635 1912 41644 1952
rect 41684 1912 41693 1952
rect 41635 1911 41693 1912
rect 39819 1893 39861 1902
rect 29827 1881 29885 1882
rect 6123 1868 6165 1877
rect 6123 1828 6124 1868
rect 6164 1828 6165 1868
rect 6123 1819 6165 1828
rect 8427 1868 8469 1877
rect 8427 1828 8428 1868
rect 8468 1828 8469 1868
rect 8427 1819 8469 1828
rect 10627 1868 10685 1869
rect 10627 1828 10636 1868
rect 10676 1828 10685 1868
rect 10627 1827 10685 1828
rect 11595 1868 11637 1877
rect 11595 1828 11596 1868
rect 11636 1828 11637 1868
rect 11595 1819 11637 1828
rect 11691 1868 11733 1877
rect 11691 1828 11692 1868
rect 11732 1828 11733 1868
rect 11691 1819 11733 1828
rect 13027 1868 13085 1869
rect 13027 1828 13036 1868
rect 13076 1828 13085 1868
rect 13027 1827 13085 1828
rect 15627 1868 15669 1877
rect 15627 1828 15628 1868
rect 15668 1828 15669 1868
rect 15627 1819 15669 1828
rect 15723 1868 15765 1877
rect 15723 1828 15724 1868
rect 15764 1828 15765 1868
rect 15723 1819 15765 1828
rect 17931 1868 17973 1877
rect 17931 1828 17932 1868
rect 17972 1828 17973 1868
rect 17931 1819 17973 1828
rect 18027 1868 18069 1877
rect 18027 1828 18028 1868
rect 18068 1828 18069 1868
rect 18027 1819 18069 1828
rect 19843 1868 19901 1869
rect 19843 1828 19852 1868
rect 19892 1828 19901 1868
rect 19843 1827 19901 1828
rect 20811 1868 20853 1877
rect 20811 1828 20812 1868
rect 20852 1828 20853 1868
rect 20811 1819 20853 1828
rect 20907 1868 20949 1877
rect 20907 1828 20908 1868
rect 20948 1828 20949 1868
rect 20907 1819 20949 1828
rect 24259 1868 24317 1869
rect 24259 1828 24268 1868
rect 24308 1828 24317 1868
rect 24259 1827 24317 1828
rect 25227 1868 25269 1877
rect 25227 1828 25228 1868
rect 25268 1828 25269 1868
rect 25227 1819 25269 1828
rect 26851 1868 26909 1869
rect 26851 1828 26860 1868
rect 26900 1828 26909 1868
rect 26851 1827 26909 1828
rect 27235 1868 27293 1869
rect 27235 1828 27244 1868
rect 27284 1828 27293 1868
rect 27235 1827 27293 1828
rect 28203 1868 28245 1877
rect 28203 1828 28204 1868
rect 28244 1828 28245 1868
rect 28203 1819 28245 1828
rect 28299 1868 28341 1877
rect 28299 1828 28300 1868
rect 28340 1828 28341 1868
rect 29827 1841 29836 1881
rect 29876 1841 29885 1881
rect 29827 1840 29885 1841
rect 30211 1868 30269 1869
rect 28299 1819 28341 1828
rect 30211 1828 30220 1868
rect 30260 1828 30269 1868
rect 30211 1827 30269 1828
rect 30987 1868 31029 1877
rect 30987 1828 30988 1868
rect 31028 1828 31029 1868
rect 30987 1819 31029 1828
rect 32611 1868 32669 1869
rect 32611 1828 32620 1868
rect 32660 1828 32669 1868
rect 32611 1827 32669 1828
rect 34627 1868 34685 1869
rect 34627 1828 34636 1868
rect 34676 1828 34685 1868
rect 34627 1827 34685 1828
rect 35883 1868 35925 1877
rect 35883 1828 35884 1868
rect 35924 1828 35925 1868
rect 35883 1819 35925 1828
rect 37699 1868 37757 1869
rect 37699 1828 37708 1868
rect 37748 1828 37757 1868
rect 37699 1827 37757 1828
rect 3627 1700 3669 1709
rect 3627 1660 3628 1700
rect 3668 1660 3669 1700
rect 3627 1651 3669 1660
rect 10827 1700 10869 1709
rect 10827 1660 10828 1700
rect 10868 1660 10869 1700
rect 10827 1651 10869 1660
rect 13227 1700 13269 1709
rect 13227 1660 13228 1700
rect 13268 1660 13269 1700
rect 13227 1651 13269 1660
rect 20043 1700 20085 1709
rect 20043 1660 20044 1700
rect 20084 1660 20085 1700
rect 20043 1651 20085 1660
rect 24075 1700 24117 1709
rect 24075 1660 24076 1700
rect 24116 1660 24117 1700
rect 24075 1651 24117 1660
rect 26667 1700 26709 1709
rect 26667 1660 26668 1700
rect 26708 1660 26709 1700
rect 26667 1651 26709 1660
rect 27435 1700 27477 1709
rect 27435 1660 27436 1700
rect 27476 1660 27477 1700
rect 27435 1651 27477 1660
rect 29643 1700 29685 1709
rect 29643 1660 29644 1700
rect 29684 1660 29685 1700
rect 29643 1651 29685 1660
rect 30027 1700 30069 1709
rect 30027 1660 30028 1700
rect 30068 1660 30069 1700
rect 30027 1651 30069 1660
rect 32427 1700 32469 1709
rect 32427 1660 32428 1700
rect 32468 1660 32469 1700
rect 32427 1651 32469 1660
rect 32811 1700 32853 1709
rect 32811 1660 32812 1700
rect 32852 1660 32853 1700
rect 32811 1651 32853 1660
rect 34443 1700 34485 1709
rect 34443 1660 34444 1700
rect 34484 1660 34485 1700
rect 34443 1651 34485 1660
rect 37515 1700 37557 1709
rect 37515 1660 37516 1700
rect 37556 1660 37557 1700
rect 37515 1651 37557 1660
rect 1152 1532 41856 1556
rect 1152 1492 3688 1532
rect 3728 1492 3770 1532
rect 3810 1492 3852 1532
rect 3892 1492 3934 1532
rect 3974 1492 4016 1532
rect 4056 1492 18808 1532
rect 18848 1492 18890 1532
rect 18930 1492 18972 1532
rect 19012 1492 19054 1532
rect 19094 1492 19136 1532
rect 19176 1492 33928 1532
rect 33968 1492 34010 1532
rect 34050 1492 34092 1532
rect 34132 1492 34174 1532
rect 34214 1492 34256 1532
rect 34296 1492 41856 1532
rect 1152 1468 41856 1492
rect 10539 1364 10581 1373
rect 10539 1324 10540 1364
rect 10580 1324 10581 1364
rect 10539 1315 10581 1324
rect 16683 1364 16725 1373
rect 16683 1324 16684 1364
rect 16724 1324 16725 1364
rect 16683 1315 16725 1324
rect 20427 1364 20469 1373
rect 20427 1324 20428 1364
rect 20468 1324 20469 1364
rect 20427 1315 20469 1324
rect 22155 1364 22197 1373
rect 22155 1324 22156 1364
rect 22196 1324 22197 1364
rect 22155 1315 22197 1324
rect 24939 1364 24981 1373
rect 24939 1324 24940 1364
rect 24980 1324 24981 1364
rect 24939 1315 24981 1324
rect 25611 1364 25653 1373
rect 25611 1324 25612 1364
rect 25652 1324 25653 1364
rect 25611 1315 25653 1324
rect 30603 1364 30645 1373
rect 30603 1324 30604 1364
rect 30644 1324 30645 1364
rect 30603 1315 30645 1324
rect 38091 1364 38133 1373
rect 38091 1324 38092 1364
rect 38132 1324 38133 1364
rect 38091 1315 38133 1324
rect 12171 1280 12213 1289
rect 12171 1240 12172 1280
rect 12212 1240 12213 1280
rect 12171 1231 12213 1240
rect 13803 1280 13845 1289
rect 13803 1240 13804 1280
rect 13844 1240 13845 1280
rect 13803 1231 13845 1240
rect 18795 1280 18837 1289
rect 18795 1240 18796 1280
rect 18836 1240 18837 1280
rect 18795 1231 18837 1240
rect 33195 1280 33237 1289
rect 33195 1240 33196 1280
rect 33236 1240 33237 1280
rect 33195 1231 33237 1240
rect 34827 1280 34869 1289
rect 34827 1240 34828 1280
rect 34868 1240 34869 1280
rect 34827 1231 34869 1240
rect 36459 1280 36501 1289
rect 36459 1240 36460 1280
rect 36500 1240 36501 1280
rect 36459 1231 36501 1240
rect 41067 1280 41109 1289
rect 41067 1240 41068 1280
rect 41108 1240 41109 1280
rect 41067 1231 41109 1240
rect 5739 1196 5781 1205
rect 5739 1156 5740 1196
rect 5780 1156 5781 1196
rect 5739 1147 5781 1156
rect 5835 1196 5877 1205
rect 5835 1156 5836 1196
rect 5876 1156 5877 1196
rect 5835 1147 5877 1156
rect 22915 1196 22973 1197
rect 22915 1156 22924 1196
rect 22964 1156 22973 1196
rect 22915 1155 22973 1156
rect 28483 1196 28541 1197
rect 28483 1156 28492 1196
rect 28532 1156 28541 1196
rect 28483 1155 28541 1156
rect 30979 1196 31037 1197
rect 30979 1156 30988 1196
rect 31028 1156 31037 1196
rect 30979 1155 31037 1156
rect 31755 1196 31797 1205
rect 31755 1156 31756 1196
rect 31796 1156 31797 1196
rect 25795 1154 25853 1155
rect 6795 1126 6837 1135
rect 1315 1112 1373 1113
rect 1315 1072 1324 1112
rect 1364 1072 1373 1112
rect 1315 1071 1373 1072
rect 2563 1112 2621 1113
rect 2563 1072 2572 1112
rect 2612 1072 2621 1112
rect 2563 1071 2621 1072
rect 3043 1112 3101 1113
rect 3043 1072 3052 1112
rect 3092 1072 3101 1112
rect 3043 1071 3101 1072
rect 4291 1112 4349 1113
rect 4291 1072 4300 1112
rect 4340 1072 4349 1112
rect 4291 1071 4349 1072
rect 5259 1112 5301 1121
rect 5259 1072 5260 1112
rect 5300 1072 5301 1112
rect 5259 1063 5301 1072
rect 5355 1112 5397 1121
rect 5355 1072 5356 1112
rect 5396 1072 5397 1112
rect 5355 1063 5397 1072
rect 6307 1112 6365 1113
rect 6307 1072 6316 1112
rect 6356 1072 6365 1112
rect 6795 1086 6796 1126
rect 6836 1086 6837 1126
rect 25795 1114 25804 1154
rect 25844 1114 25853 1154
rect 31755 1147 31797 1156
rect 31851 1196 31893 1205
rect 31851 1156 31852 1196
rect 31892 1156 31893 1196
rect 31851 1147 31893 1156
rect 39907 1196 39965 1197
rect 39907 1156 39916 1196
rect 39956 1156 39965 1196
rect 39907 1155 39965 1156
rect 40099 1196 40157 1197
rect 40099 1156 40108 1196
rect 40148 1156 40157 1196
rect 40099 1155 40157 1156
rect 40483 1196 40541 1197
rect 40483 1156 40492 1196
rect 40532 1156 40541 1196
rect 40483 1155 40541 1156
rect 40867 1196 40925 1197
rect 40867 1156 40876 1196
rect 40916 1156 40925 1196
rect 40867 1155 40925 1156
rect 41251 1196 41309 1197
rect 41251 1156 41260 1196
rect 41300 1156 41309 1196
rect 41251 1155 41309 1156
rect 32811 1126 32853 1135
rect 25795 1113 25853 1114
rect 6795 1077 6837 1086
rect 9091 1112 9149 1113
rect 6307 1071 6365 1072
rect 9091 1072 9100 1112
rect 9140 1072 9149 1112
rect 9091 1071 9149 1072
rect 10339 1112 10397 1113
rect 10339 1072 10348 1112
rect 10388 1072 10397 1112
rect 10339 1071 10397 1072
rect 10723 1112 10781 1113
rect 10723 1072 10732 1112
rect 10772 1072 10781 1112
rect 10723 1071 10781 1072
rect 11971 1112 12029 1113
rect 11971 1072 11980 1112
rect 12020 1072 12029 1112
rect 11971 1071 12029 1072
rect 12355 1112 12413 1113
rect 12355 1072 12364 1112
rect 12404 1072 12413 1112
rect 12355 1071 12413 1072
rect 13603 1112 13661 1113
rect 13603 1072 13612 1112
rect 13652 1072 13661 1112
rect 13603 1071 13661 1072
rect 15235 1112 15293 1113
rect 15235 1072 15244 1112
rect 15284 1072 15293 1112
rect 15235 1071 15293 1072
rect 16483 1112 16541 1113
rect 16483 1072 16492 1112
rect 16532 1072 16541 1112
rect 16483 1071 16541 1072
rect 17347 1112 17405 1113
rect 17347 1072 17356 1112
rect 17396 1072 17405 1112
rect 17347 1071 17405 1072
rect 18595 1112 18653 1113
rect 18595 1072 18604 1112
rect 18644 1072 18653 1112
rect 18595 1071 18653 1072
rect 18979 1112 19037 1113
rect 18979 1072 18988 1112
rect 19028 1072 19037 1112
rect 18979 1071 19037 1072
rect 20227 1112 20285 1113
rect 20227 1072 20236 1112
rect 20276 1072 20285 1112
rect 20227 1071 20285 1072
rect 20707 1112 20765 1113
rect 20707 1072 20716 1112
rect 20756 1072 20765 1112
rect 20707 1071 20765 1072
rect 21955 1112 22013 1113
rect 21955 1072 21964 1112
rect 22004 1072 22013 1112
rect 21955 1071 22013 1072
rect 24739 1112 24797 1113
rect 24739 1072 24748 1112
rect 24788 1072 24797 1112
rect 24739 1071 24797 1072
rect 27043 1112 27101 1113
rect 27043 1072 27052 1112
rect 27092 1072 27101 1112
rect 27043 1071 27101 1072
rect 29155 1112 29213 1113
rect 29155 1072 29164 1112
rect 29204 1072 29213 1112
rect 29155 1071 29213 1072
rect 30403 1112 30461 1113
rect 30403 1072 30412 1112
rect 30452 1072 30461 1112
rect 30403 1071 30461 1072
rect 31275 1112 31317 1121
rect 31275 1072 31276 1112
rect 31316 1072 31317 1112
rect 23491 1070 23549 1071
rect 4491 1028 4533 1037
rect 23491 1030 23500 1070
rect 23540 1030 23549 1070
rect 31275 1063 31317 1072
rect 31371 1112 31413 1121
rect 31371 1072 31372 1112
rect 31412 1072 31413 1112
rect 31371 1063 31413 1072
rect 32323 1112 32381 1113
rect 32323 1072 32332 1112
rect 32372 1072 32381 1112
rect 32811 1086 32812 1126
rect 32852 1086 32853 1126
rect 32811 1077 32853 1086
rect 33379 1112 33437 1113
rect 32323 1071 32381 1072
rect 33379 1072 33388 1112
rect 33428 1072 33437 1112
rect 33379 1071 33437 1072
rect 34627 1112 34685 1113
rect 34627 1072 34636 1112
rect 34676 1072 34685 1112
rect 34627 1071 34685 1072
rect 35011 1112 35069 1113
rect 35011 1072 35020 1112
rect 35060 1072 35069 1112
rect 35011 1071 35069 1072
rect 36259 1112 36317 1113
rect 36259 1072 36268 1112
rect 36308 1072 36317 1112
rect 36259 1071 36317 1072
rect 36643 1112 36701 1113
rect 36643 1072 36652 1112
rect 36692 1072 36701 1112
rect 36643 1071 36701 1072
rect 37891 1112 37949 1113
rect 37891 1072 37900 1112
rect 37940 1072 37949 1112
rect 37891 1071 37949 1072
rect 38275 1112 38333 1113
rect 38275 1072 38284 1112
rect 38324 1072 38333 1112
rect 38275 1071 38333 1072
rect 39523 1112 39581 1113
rect 39523 1072 39532 1112
rect 39572 1072 39581 1112
rect 39523 1071 39581 1072
rect 23491 1029 23549 1030
rect 4491 988 4492 1028
rect 4532 988 4533 1028
rect 4491 979 4533 988
rect 33003 1028 33045 1037
rect 33003 988 33004 1028
rect 33044 988 33045 1028
rect 33003 979 33045 988
rect 2763 944 2805 953
rect 2763 904 2764 944
rect 2804 904 2805 944
rect 2763 895 2805 904
rect 6987 944 7029 953
rect 6987 904 6988 944
rect 7028 904 7029 944
rect 6987 895 7029 904
rect 23115 944 23157 953
rect 23115 904 23116 944
rect 23156 904 23157 944
rect 23115 895 23157 904
rect 28683 944 28725 953
rect 28683 904 28684 944
rect 28724 904 28725 944
rect 28683 895 28725 904
rect 30795 944 30837 953
rect 30795 904 30796 944
rect 30836 904 30837 944
rect 30795 895 30837 904
rect 39723 944 39765 953
rect 39723 904 39724 944
rect 39764 904 39765 944
rect 39723 895 39765 904
rect 40299 944 40341 953
rect 40299 904 40300 944
rect 40340 904 40341 944
rect 40299 895 40341 904
rect 40683 944 40725 953
rect 40683 904 40684 944
rect 40724 904 40725 944
rect 40683 895 40725 904
rect 41451 944 41493 953
rect 41451 904 41452 944
rect 41492 904 41493 944
rect 41451 895 41493 904
rect 1152 776 41856 800
rect 1152 736 4928 776
rect 4968 736 5010 776
rect 5050 736 5092 776
rect 5132 736 5174 776
rect 5214 736 5256 776
rect 5296 736 20048 776
rect 20088 736 20130 776
rect 20170 736 20212 776
rect 20252 736 20294 776
rect 20334 736 20376 776
rect 20416 736 35168 776
rect 35208 736 35250 776
rect 35290 736 35332 776
rect 35372 736 35414 776
rect 35454 736 35496 776
rect 35536 736 41856 776
rect 1152 712 41856 736
<< via1 >>
rect 4928 9808 4968 9848
rect 5010 9808 5050 9848
rect 5092 9808 5132 9848
rect 5174 9808 5214 9848
rect 5256 9808 5296 9848
rect 20048 9808 20088 9848
rect 20130 9808 20170 9848
rect 20212 9808 20252 9848
rect 20294 9808 20334 9848
rect 20376 9808 20416 9848
rect 35168 9808 35208 9848
rect 35250 9808 35290 9848
rect 35332 9808 35372 9848
rect 35414 9808 35454 9848
rect 35496 9808 35536 9848
rect 4108 9640 4148 9680
rect 4588 9640 4628 9680
rect 9196 9640 9236 9680
rect 11692 9640 11732 9680
rect 13324 9640 13364 9680
rect 16684 9640 16724 9680
rect 19468 9640 19508 9680
rect 21388 9640 21428 9680
rect 32044 9640 32084 9680
rect 32428 9640 32468 9680
rect 32812 9640 32852 9680
rect 37708 9640 37748 9680
rect 40684 9640 40724 9680
rect 41452 9640 41492 9680
rect 2956 9556 2996 9596
rect 1516 9472 1556 9512
rect 2764 9472 2804 9512
rect 3340 9472 3380 9512
rect 3436 9472 3476 9512
rect 3532 9472 3572 9512
rect 3628 9472 3668 9512
rect 3820 9472 3860 9512
rect 3916 9472 3956 9512
rect 4300 9472 4340 9512
rect 4396 9472 4436 9512
rect 4492 9472 4532 9512
rect 7756 9472 7796 9512
rect 9004 9472 9044 9512
rect 10252 9472 10292 9512
rect 11500 9472 11540 9512
rect 11884 9472 11924 9512
rect 13132 9472 13172 9512
rect 15244 9472 15284 9512
rect 16492 9472 16532 9512
rect 17836 9472 17876 9512
rect 19084 9472 19124 9512
rect 22444 9472 22484 9512
rect 23692 9472 23732 9512
rect 24268 9472 24308 9512
rect 25516 9472 25556 9512
rect 27724 9472 27764 9512
rect 28972 9472 29012 9512
rect 29548 9472 29588 9512
rect 30508 9472 30548 9512
rect 30796 9472 30836 9512
rect 31660 9472 31700 9512
rect 34540 9472 34580 9512
rect 35212 9472 35252 9512
rect 36172 9472 36212 9512
rect 36556 9472 36596 9512
rect 19660 9388 19700 9428
rect 21196 9388 21236 9428
rect 32236 9388 32276 9428
rect 32620 9388 32660 9428
rect 33004 9388 33044 9428
rect 37900 9388 37940 9428
rect 40492 9388 40532 9428
rect 40876 9388 40916 9428
rect 41260 9388 41300 9428
rect 33388 9304 33428 9344
rect 34828 9304 34868 9344
rect 36844 9304 36884 9344
rect 41068 9304 41108 9344
rect 19276 9220 19316 9260
rect 23884 9220 23924 9260
rect 25708 9220 25748 9260
rect 29164 9220 29204 9260
rect 34252 9220 34292 9260
rect 35884 9220 35924 9260
rect 3688 9052 3728 9092
rect 3770 9052 3810 9092
rect 3852 9052 3892 9092
rect 3934 9052 3974 9092
rect 4016 9052 4056 9092
rect 18808 9052 18848 9092
rect 18890 9052 18930 9092
rect 18972 9052 19012 9092
rect 19054 9052 19094 9092
rect 19136 9052 19176 9092
rect 33928 9052 33968 9092
rect 34010 9052 34050 9092
rect 34092 9052 34132 9092
rect 34174 9052 34214 9092
rect 34256 9052 34296 9092
rect 3628 8884 3668 8924
rect 9484 8800 9524 8840
rect 13900 8800 13940 8840
rect 15532 8800 15572 8840
rect 20044 8800 20084 8840
rect 29260 8800 29300 8840
rect 29740 8800 29780 8840
rect 31756 8800 31796 8840
rect 32140 8800 32180 8840
rect 32524 8800 32564 8840
rect 32908 8800 32948 8840
rect 36172 8800 36212 8840
rect 36556 8800 36596 8840
rect 38764 8800 38804 8840
rect 39148 8800 39188 8840
rect 40012 8800 40052 8840
rect 40396 8800 40436 8840
rect 41068 8800 41108 8840
rect 41452 8800 41492 8840
rect 19852 8716 19892 8756
rect 22444 8716 22484 8756
rect 1612 8632 1652 8672
rect 2860 8632 2900 8672
rect 3532 8632 3572 8672
rect 3628 8632 3668 8672
rect 3820 8632 3860 8672
rect 4012 8632 4052 8672
rect 4108 8632 4148 8672
rect 4204 8632 4244 8672
rect 4300 8632 4340 8672
rect 4780 8632 4820 8672
rect 6028 8632 6068 8672
rect 6412 8632 6452 8672
rect 7660 8632 7700 8672
rect 8044 8632 8084 8672
rect 9292 8632 9332 8672
rect 9676 8632 9716 8672
rect 10924 8632 10964 8672
rect 12460 8632 12500 8672
rect 13708 8632 13748 8672
rect 14092 8632 14132 8672
rect 15340 8632 15380 8672
rect 15916 8632 15956 8672
rect 17164 8632 17204 8672
rect 17644 8632 17684 8672
rect 17740 8632 17780 8672
rect 18124 8632 18164 8672
rect 19228 8674 19268 8714
rect 29452 8716 29492 8756
rect 29932 8716 29972 8756
rect 31948 8716 31988 8756
rect 32332 8716 32372 8756
rect 32716 8716 32756 8756
rect 33100 8716 33140 8756
rect 36364 8716 36404 8756
rect 36748 8716 36788 8756
rect 38572 8716 38612 8756
rect 38956 8716 38996 8756
rect 39820 8716 39860 8756
rect 40204 8716 40244 8756
rect 40876 8716 40916 8756
rect 41260 8716 41300 8756
rect 18220 8632 18260 8672
rect 18700 8632 18740 8672
rect 20236 8632 20276 8672
rect 21484 8632 21524 8672
rect 21964 8632 22004 8672
rect 22060 8632 22100 8672
rect 22540 8632 22580 8672
rect 23020 8632 23060 8672
rect 23548 8641 23588 8681
rect 25420 8632 25460 8672
rect 25516 8632 25556 8672
rect 25900 8632 25940 8672
rect 25996 8632 26036 8672
rect 26476 8632 26516 8672
rect 27004 8641 27044 8681
rect 27532 8632 27572 8672
rect 28780 8632 28820 8672
rect 30124 8632 30164 8672
rect 31372 8632 31412 8672
rect 33964 8632 34004 8672
rect 34828 8632 34868 8672
rect 36940 8632 36980 8672
rect 38188 8632 38228 8672
rect 3052 8548 3092 8588
rect 17356 8548 17396 8588
rect 21676 8548 21716 8588
rect 27340 8548 27380 8588
rect 33580 8548 33620 8588
rect 6220 8464 6260 8504
rect 7852 8464 7892 8504
rect 11116 8464 11156 8504
rect 19372 8464 19412 8504
rect 23692 8464 23732 8504
rect 27148 8464 27188 8504
rect 31564 8464 31604 8504
rect 35980 8464 36020 8504
rect 38380 8464 38420 8504
rect 4928 8296 4968 8336
rect 5010 8296 5050 8336
rect 5092 8296 5132 8336
rect 5174 8296 5214 8336
rect 5256 8296 5296 8336
rect 20048 8296 20088 8336
rect 20130 8296 20170 8336
rect 20212 8296 20252 8336
rect 20294 8296 20334 8336
rect 20376 8296 20416 8336
rect 35168 8296 35208 8336
rect 35250 8296 35290 8336
rect 35332 8296 35372 8336
rect 35414 8296 35454 8336
rect 35496 8296 35536 8336
rect 2860 8128 2900 8168
rect 8332 8128 8372 8168
rect 10348 8128 10388 8168
rect 22540 8128 22580 8168
rect 33292 8128 33332 8168
rect 40684 8128 40724 8168
rect 41452 8128 41492 8168
rect 7372 8044 7412 8084
rect 27052 8044 27092 8084
rect 30412 8044 30452 8084
rect 32812 8044 32852 8084
rect 1420 7960 1460 8000
rect 2668 7960 2708 8000
rect 3052 7960 3092 8000
rect 3436 7960 3476 8000
rect 3532 7960 3572 8000
rect 3628 7960 3668 8000
rect 4012 7960 4052 8000
rect 5260 7960 5300 8000
rect 5932 7960 5972 8000
rect 7180 7960 7220 8000
rect 7852 7960 7892 8000
rect 7948 7960 7988 8000
rect 8044 7960 8084 8000
rect 8140 7960 8180 8000
rect 8524 7960 8564 8000
rect 8620 7960 8660 8000
rect 8908 7960 8948 8000
rect 10156 7960 10196 8000
rect 10540 7960 10580 8000
rect 11788 7960 11828 8000
rect 12172 7960 12212 8000
rect 13420 7960 13460 8000
rect 13804 7960 13844 8000
rect 15052 7960 15092 8000
rect 16108 7960 16148 8000
rect 17356 7960 17396 8000
rect 17836 7960 17876 8000
rect 19084 7960 19124 8000
rect 19756 7960 19796 8000
rect 21004 7960 21044 8000
rect 22828 7960 22868 8000
rect 24076 7960 24116 8000
rect 25324 7960 25364 8000
rect 25420 7960 25460 8000
rect 25900 7960 25940 8000
rect 26380 7960 26420 8000
rect 26860 7946 26900 7986
rect 28684 7960 28724 8000
rect 28780 7960 28820 8000
rect 29740 7960 29780 8000
rect 3148 7876 3188 7916
rect 21580 7876 21620 7916
rect 22348 7876 22388 7916
rect 25804 7876 25844 7916
rect 27436 7876 27476 7916
rect 29164 7876 29204 7916
rect 29260 7876 29300 7916
rect 30268 7918 30308 7958
rect 31084 7960 31124 8000
rect 31180 7960 31220 8000
rect 32140 7960 32180 8000
rect 32620 7946 32660 7986
rect 34060 7960 34100 8000
rect 34444 7960 34484 8000
rect 35308 7960 35348 8000
rect 36844 7960 36884 8000
rect 38092 7960 38132 8000
rect 30796 7876 30836 7916
rect 31564 7876 31604 7916
rect 31660 7876 31700 7916
rect 33100 7876 33140 7916
rect 40492 7876 40532 7916
rect 40876 7876 40916 7916
rect 41260 7876 41300 7916
rect 30604 7792 30644 7832
rect 41068 7792 41108 7832
rect 2860 7708 2900 7748
rect 3820 7708 3860 7748
rect 5452 7708 5492 7748
rect 11980 7708 12020 7748
rect 13612 7708 13652 7748
rect 15244 7708 15284 7748
rect 17548 7708 17588 7748
rect 19276 7708 19316 7748
rect 21196 7708 21236 7748
rect 21388 7708 21428 7748
rect 24268 7708 24308 7748
rect 27244 7708 27284 7748
rect 36460 7708 36500 7748
rect 36652 7708 36692 7748
rect 3688 7540 3728 7580
rect 3770 7540 3810 7580
rect 3852 7540 3892 7580
rect 3934 7540 3974 7580
rect 4016 7540 4056 7580
rect 18808 7540 18848 7580
rect 18890 7540 18930 7580
rect 18972 7540 19012 7580
rect 19054 7540 19094 7580
rect 19136 7540 19176 7580
rect 33928 7540 33968 7580
rect 34010 7540 34050 7580
rect 34092 7540 34132 7580
rect 34174 7540 34214 7580
rect 34256 7540 34296 7580
rect 3724 7372 3764 7412
rect 25612 7372 25652 7412
rect 26284 7372 26324 7412
rect 30316 7372 30356 7412
rect 33100 7372 33140 7412
rect 40684 7372 40724 7412
rect 4396 7288 4436 7328
rect 7756 7204 7796 7244
rect 14284 7204 14324 7244
rect 14380 7204 14420 7244
rect 21388 7204 21428 7244
rect 23404 7204 23444 7244
rect 25900 7204 25940 7244
rect 30700 7204 30740 7244
rect 38476 7204 38516 7244
rect 2956 7120 2996 7160
rect 3052 7120 3092 7160
rect 3148 7120 3188 7160
rect 3244 7120 3284 7160
rect 3436 7120 3476 7160
rect 3532 7120 3572 7160
rect 4396 7112 4436 7152
rect 4780 7120 4820 7160
rect 4876 7120 4916 7160
rect 5260 7120 5300 7160
rect 5356 7120 5396 7160
rect 5452 7120 5492 7160
rect 5548 7120 5588 7160
rect 5740 7120 5780 7160
rect 5836 7120 5876 7160
rect 5932 7120 5972 7160
rect 6028 7120 6068 7160
rect 6220 7120 6260 7160
rect 6316 7120 6356 7160
rect 6796 7120 6836 7160
rect 6892 7120 6932 7160
rect 6988 7120 7028 7160
rect 7276 7120 7316 7160
rect 7372 7120 7412 7160
rect 7852 7120 7892 7160
rect 8332 7120 8372 7160
rect 8860 7129 8900 7169
rect 9196 7120 9236 7160
rect 9292 7120 9332 7160
rect 9676 7120 9716 7160
rect 9772 7120 9812 7160
rect 9868 7120 9908 7160
rect 9964 7120 10004 7160
rect 11308 7120 11348 7160
rect 11404 7120 11444 7160
rect 11788 7120 11828 7160
rect 11884 7120 11924 7160
rect 12364 7120 12404 7160
rect 12844 7134 12884 7174
rect 13804 7120 13844 7160
rect 13900 7120 13940 7160
rect 14860 7120 14900 7160
rect 15340 7134 15380 7174
rect 16300 7120 16340 7160
rect 17548 7120 17588 7160
rect 19276 7120 19316 7160
rect 19372 7120 19412 7160
rect 19756 7120 19796 7160
rect 20860 7162 20900 7202
rect 40492 7204 40532 7244
rect 40876 7204 40916 7244
rect 19852 7120 19892 7160
rect 20332 7120 20372 7160
rect 24172 7120 24212 7160
rect 25420 7120 25460 7160
rect 26476 7120 26516 7160
rect 27724 7120 27764 7160
rect 28876 7120 28916 7160
rect 30124 7120 30164 7160
rect 31660 7120 31700 7160
rect 32908 7120 32948 7160
rect 33388 7120 33428 7160
rect 34636 7120 34676 7160
rect 35116 7120 35156 7160
rect 35212 7120 35252 7160
rect 35596 7120 35636 7160
rect 35692 7120 35732 7160
rect 36172 7120 36212 7160
rect 36652 7134 36692 7174
rect 37996 7120 38036 7160
rect 38092 7120 38132 7160
rect 38572 7120 38612 7160
rect 39052 7120 39092 7160
rect 39532 7125 39572 7165
rect 3628 7036 3668 7076
rect 9004 7036 9044 7076
rect 21004 7036 21044 7076
rect 34828 7036 34868 7076
rect 3724 6952 3764 6992
rect 4588 6952 4628 6992
rect 5068 6952 5108 6992
rect 6508 6952 6548 6992
rect 6700 6952 6740 6992
rect 9484 6952 9524 6992
rect 13036 6952 13076 6992
rect 15532 6952 15572 6992
rect 17740 6952 17780 6992
rect 21196 6952 21236 6992
rect 23212 6952 23252 6992
rect 26092 6952 26132 6992
rect 30508 6952 30548 6992
rect 36844 6952 36884 6992
rect 39724 6952 39764 6992
rect 41068 6952 41108 6992
rect 4928 6784 4968 6824
rect 5010 6784 5050 6824
rect 5092 6784 5132 6824
rect 5174 6784 5214 6824
rect 5256 6784 5296 6824
rect 20048 6784 20088 6824
rect 20130 6784 20170 6824
rect 20212 6784 20252 6824
rect 20294 6784 20334 6824
rect 20376 6784 20416 6824
rect 35168 6784 35208 6824
rect 35250 6784 35290 6824
rect 35332 6784 35372 6824
rect 35414 6784 35454 6824
rect 35496 6784 35536 6824
rect 5836 6616 5876 6656
rect 6316 6616 6356 6656
rect 9004 6616 9044 6656
rect 21292 6616 21332 6656
rect 37324 6616 37364 6656
rect 39436 6616 39476 6656
rect 40684 6616 40724 6656
rect 3532 6532 3572 6572
rect 6796 6532 6836 6572
rect 19660 6532 19700 6572
rect 23308 6532 23348 6572
rect 1708 6448 1748 6488
rect 2956 6448 2996 6488
rect 3436 6448 3476 6488
rect 3628 6448 3668 6488
rect 3916 6448 3956 6488
rect 4204 6448 4244 6488
rect 4300 6448 4340 6488
rect 4871 6448 4911 6488
rect 4972 6448 5012 6488
rect 5068 6448 5108 6488
rect 5260 6448 5300 6488
rect 5356 6448 5396 6488
rect 5548 6448 5588 6488
rect 5644 6448 5684 6488
rect 5740 6448 5780 6488
rect 6028 6448 6068 6488
rect 6124 6448 6164 6488
rect 6220 6448 6260 6488
rect 6892 6448 6932 6488
rect 7180 6448 7220 6488
rect 7564 6448 7604 6488
rect 8812 6448 8852 6488
rect 9868 6448 9908 6488
rect 11116 6448 11156 6488
rect 12268 6448 12308 6488
rect 13516 6448 13556 6488
rect 14764 6448 14804 6488
rect 16012 6448 16052 6488
rect 17932 6448 17972 6488
rect 18028 6448 18068 6488
rect 18412 6448 18452 6488
rect 18988 6448 19028 6488
rect 19468 6434 19508 6474
rect 19852 6448 19892 6488
rect 21100 6448 21140 6488
rect 21580 6448 21620 6488
rect 21676 6448 21716 6488
rect 22060 6448 22100 6488
rect 22636 6448 22676 6488
rect 24364 6448 24404 6488
rect 25612 6448 25652 6488
rect 26476 6448 26516 6488
rect 27724 6448 27764 6488
rect 28300 6448 28340 6488
rect 29548 6448 29588 6488
rect 30508 6448 30548 6488
rect 32524 6448 32564 6488
rect 33772 6448 33812 6488
rect 36940 6448 36980 6488
rect 18508 6364 18548 6404
rect 22156 6364 22196 6404
rect 23164 6406 23204 6446
rect 31756 6406 31796 6446
rect 37996 6448 38036 6488
rect 39244 6448 39284 6488
rect 23692 6364 23732 6404
rect 26284 6364 26324 6404
rect 32332 6364 32372 6404
rect 36556 6364 36596 6404
rect 39820 6364 39860 6404
rect 40492 6364 40532 6404
rect 40876 6364 40916 6404
rect 3148 6280 3188 6320
rect 4588 6280 4628 6320
rect 6508 6280 6548 6320
rect 27916 6280 27956 6320
rect 36364 6280 36404 6320
rect 39628 6280 39668 6320
rect 41068 6280 41108 6320
rect 5356 6196 5396 6236
rect 11308 6196 11348 6236
rect 13708 6196 13748 6236
rect 16204 6196 16244 6236
rect 23500 6196 23540 6236
rect 25804 6196 25844 6236
rect 26092 6196 26132 6236
rect 29740 6196 29780 6236
rect 31948 6196 31988 6236
rect 32140 6196 32180 6236
rect 33964 6196 34004 6236
rect 3688 6028 3728 6068
rect 3770 6028 3810 6068
rect 3852 6028 3892 6068
rect 3934 6028 3974 6068
rect 4016 6028 4056 6068
rect 18808 6028 18848 6068
rect 18890 6028 18930 6068
rect 18972 6028 19012 6068
rect 19054 6028 19094 6068
rect 19136 6028 19176 6068
rect 33928 6028 33968 6068
rect 34010 6028 34050 6068
rect 34092 6028 34132 6068
rect 34174 6028 34214 6068
rect 34256 6028 34296 6068
rect 4108 5860 4148 5900
rect 4876 5860 4916 5900
rect 19468 5860 19508 5900
rect 23500 5860 23540 5900
rect 41068 5860 41108 5900
rect 5356 5776 5396 5816
rect 40684 5776 40724 5816
rect 10540 5692 10580 5732
rect 20236 5692 20276 5732
rect 24460 5692 24500 5732
rect 26860 5692 26900 5732
rect 1612 5608 1652 5648
rect 2860 5608 2900 5648
rect 4108 5608 4148 5648
rect 4300 5608 4340 5648
rect 4396 5608 4436 5648
rect 4588 5608 4628 5648
rect 4876 5608 4916 5648
rect 5068 5608 5108 5648
rect 5164 5608 5204 5648
rect 5356 5608 5396 5648
rect 5644 5608 5684 5648
rect 5740 5608 5780 5648
rect 6124 5608 6164 5648
rect 6220 5608 6260 5648
rect 6700 5608 6740 5648
rect 7180 5613 7220 5653
rect 8332 5608 8372 5648
rect 9580 5608 9620 5648
rect 10060 5608 10100 5648
rect 10156 5608 10196 5648
rect 10636 5608 10676 5648
rect 11116 5608 11156 5648
rect 11596 5622 11636 5662
rect 13132 5608 13172 5648
rect 14380 5608 14420 5648
rect 14764 5608 14804 5648
rect 16012 5608 16052 5648
rect 16396 5608 16436 5648
rect 17644 5608 17684 5648
rect 18028 5608 18068 5648
rect 19276 5608 19316 5648
rect 22060 5608 22100 5648
rect 23308 5608 23348 5648
rect 23884 5608 23924 5648
rect 23980 5608 24020 5648
rect 25468 5650 25508 5690
rect 29740 5692 29780 5732
rect 35884 5692 35924 5732
rect 24364 5608 24404 5648
rect 24940 5608 24980 5648
rect 27628 5608 27668 5648
rect 27724 5608 27764 5648
rect 28108 5608 28148 5648
rect 28204 5608 28244 5648
rect 28695 5621 28735 5661
rect 29212 5650 29252 5690
rect 40492 5692 40532 5732
rect 40876 5692 40916 5732
rect 30124 5608 30164 5648
rect 31372 5608 31412 5648
rect 31852 5608 31892 5648
rect 31948 5608 31988 5648
rect 32332 5608 32372 5648
rect 32428 5608 32468 5648
rect 32908 5608 32948 5648
rect 33388 5622 33428 5662
rect 35308 5608 35348 5648
rect 35404 5608 35444 5648
rect 35788 5608 35828 5648
rect 36364 5608 36404 5648
rect 36892 5617 36932 5657
rect 3052 5524 3092 5564
rect 7372 5524 7412 5564
rect 9772 5524 9812 5564
rect 29356 5524 29396 5564
rect 31564 5524 31604 5564
rect 11788 5440 11828 5480
rect 14572 5440 14612 5480
rect 16204 5440 16244 5480
rect 17836 5440 17876 5480
rect 20428 5440 20468 5480
rect 25612 5440 25652 5480
rect 27052 5440 27092 5480
rect 29548 5440 29588 5480
rect 33580 5440 33620 5480
rect 37036 5440 37076 5480
rect 4928 5272 4968 5312
rect 5010 5272 5050 5312
rect 5092 5272 5132 5312
rect 5174 5272 5214 5312
rect 5256 5272 5296 5312
rect 20048 5272 20088 5312
rect 20130 5272 20170 5312
rect 20212 5272 20252 5312
rect 20294 5272 20334 5312
rect 20376 5272 20416 5312
rect 35168 5272 35208 5312
rect 35250 5272 35290 5312
rect 35332 5272 35372 5312
rect 35414 5272 35454 5312
rect 35496 5272 35536 5312
rect 4204 5104 4244 5144
rect 4588 5104 4628 5144
rect 20524 5104 20564 5144
rect 35596 5104 35636 5144
rect 37324 5104 37364 5144
rect 3628 5020 3668 5060
rect 7276 5020 7316 5060
rect 15628 5020 15668 5060
rect 18508 5020 18548 5060
rect 23116 5020 23156 5060
rect 25132 5020 25172 5060
rect 33676 5020 33716 5060
rect 40012 5020 40052 5060
rect 1612 4936 1652 4976
rect 2860 4936 2900 4976
rect 3724 4936 3764 4976
rect 3820 4936 3860 4976
rect 3916 4936 3956 4976
rect 4108 4936 4148 4976
rect 4300 4936 4340 4976
rect 4396 4936 4436 4976
rect 4684 4936 4724 4976
rect 5068 4936 5108 4976
rect 5260 4936 5300 4976
rect 5548 4936 5588 4976
rect 5644 4936 5684 4976
rect 6124 4936 6164 4976
rect 6604 4936 6644 4976
rect 7084 4926 7124 4966
rect 8428 4936 8468 4976
rect 8716 4936 8756 4976
rect 8812 4936 8852 4976
rect 9292 4936 9332 4976
rect 10540 4936 10580 4976
rect 11116 4936 11156 4976
rect 12364 4936 12404 4976
rect 13900 4936 13940 4976
rect 13996 4936 14036 4976
rect 14956 4936 14996 4976
rect 15436 4931 15476 4971
rect 16780 4936 16820 4976
rect 16876 4936 16916 4976
rect 17836 4936 17876 4976
rect 18316 4931 18356 4971
rect 18796 4936 18836 4976
rect 18892 4936 18932 4976
rect 19852 4936 19892 4976
rect 21676 4936 21716 4976
rect 22924 4936 22964 4976
rect 23404 4936 23444 4976
rect 6028 4852 6068 4892
rect 14380 4852 14420 4892
rect 14476 4852 14516 4892
rect 17260 4852 17300 4892
rect 17356 4852 17396 4892
rect 19276 4852 19316 4892
rect 19372 4852 19412 4892
rect 20380 4894 20420 4934
rect 23500 4936 23540 4976
rect 24460 4936 24500 4976
rect 24940 4922 24980 4962
rect 26380 4936 26420 4976
rect 27628 4936 27668 4976
rect 29068 4936 29108 4976
rect 30316 4936 30356 4976
rect 31948 4936 31988 4976
rect 32044 4936 32084 4976
rect 33004 4936 33044 4976
rect 33484 4922 33524 4962
rect 34156 4936 34196 4976
rect 35404 4936 35444 4976
rect 35884 4936 35924 4976
rect 37132 4936 37172 4976
rect 38284 4936 38324 4976
rect 38380 4936 38420 4976
rect 38764 4936 38804 4976
rect 39340 4936 39380 4976
rect 39820 4922 39860 4962
rect 20716 4852 20756 4892
rect 21100 4852 21140 4892
rect 23884 4852 23924 4892
rect 23980 4852 24020 4892
rect 25516 4852 25556 4892
rect 32428 4852 32468 4892
rect 32524 4852 32564 4892
rect 38860 4852 38900 4892
rect 40492 4852 40532 4892
rect 40876 4852 40916 4892
rect 41260 4852 41300 4892
rect 3052 4768 3092 4808
rect 21292 4768 21332 4808
rect 40684 4768 40724 4808
rect 41068 4768 41108 4808
rect 41452 4768 41492 4808
rect 4588 4684 4628 4724
rect 5164 4684 5204 4724
rect 9100 4684 9140 4724
rect 10732 4684 10772 4724
rect 12556 4684 12596 4724
rect 20908 4684 20948 4724
rect 25324 4684 25364 4724
rect 27820 4684 27860 4724
rect 30508 4684 30548 4724
rect 3688 4516 3728 4556
rect 3770 4516 3810 4556
rect 3852 4516 3892 4556
rect 3934 4516 3974 4556
rect 4016 4516 4056 4556
rect 18808 4516 18848 4556
rect 18890 4516 18930 4556
rect 18972 4516 19012 4556
rect 19054 4516 19094 4556
rect 19136 4516 19176 4556
rect 33928 4516 33968 4556
rect 34010 4516 34050 4556
rect 34092 4516 34132 4556
rect 34174 4516 34214 4556
rect 34256 4516 34296 4556
rect 9484 4348 9524 4388
rect 18796 4348 18836 4388
rect 20716 4348 20756 4388
rect 24268 4348 24308 4388
rect 33388 4348 33428 4388
rect 40300 4348 40340 4388
rect 41068 4348 41108 4388
rect 4204 4264 4244 4304
rect 5068 4264 5108 4304
rect 31276 4264 31316 4304
rect 6220 4180 6260 4220
rect 23212 4180 23252 4220
rect 23500 4180 23540 4220
rect 24076 4180 24116 4220
rect 27052 4180 27092 4220
rect 29644 4180 29684 4220
rect 32812 4180 32852 4220
rect 33196 4180 33236 4220
rect 36844 4180 36884 4220
rect 40492 4180 40532 4220
rect 40876 4180 40916 4220
rect 41260 4180 41300 4220
rect 1516 4096 1556 4136
rect 2764 4096 2804 4136
rect 3532 4096 3572 4136
rect 3820 4096 3860 4136
rect 3916 4096 3956 4136
rect 4396 4096 4436 4136
rect 4588 4096 4628 4136
rect 4684 4096 4724 4136
rect 5068 4096 5108 4136
rect 5644 4096 5684 4136
rect 5740 4096 5780 4136
rect 6124 4096 6164 4136
rect 6700 4096 6740 4136
rect 7180 4101 7220 4141
rect 8044 4096 8084 4136
rect 9292 4096 9332 4136
rect 10444 4096 10484 4136
rect 11692 4096 11732 4136
rect 12076 4096 12116 4136
rect 13324 4096 13364 4136
rect 13996 4096 14036 4136
rect 14092 4096 14132 4136
rect 14476 4096 14516 4136
rect 14572 4096 14612 4136
rect 15052 4096 15092 4136
rect 15580 4105 15620 4145
rect 17356 4096 17396 4136
rect 18604 4096 18644 4136
rect 19276 4096 19316 4136
rect 20524 4096 20564 4136
rect 21100 4096 21140 4136
rect 21196 4096 21236 4136
rect 21580 4096 21620 4136
rect 21676 4096 21716 4136
rect 22156 4096 22196 4136
rect 22636 4101 22676 4141
rect 24460 4096 24500 4136
rect 25708 4096 25748 4136
rect 27532 4096 27572 4136
rect 27628 4096 27668 4136
rect 28012 4096 28052 4136
rect 28108 4096 28148 4136
rect 28588 4096 28628 4136
rect 29116 4105 29156 4145
rect 30604 4096 30644 4136
rect 30892 4096 30932 4136
rect 33580 4096 33620 4136
rect 34828 4096 34868 4136
rect 35020 4096 35060 4136
rect 36268 4096 36308 4136
rect 37228 4096 37268 4136
rect 38476 4096 38516 4136
rect 38860 4096 38900 4136
rect 40108 4096 40148 4136
rect 2956 4012 2996 4052
rect 13516 4012 13556 4052
rect 15724 4012 15764 4052
rect 29260 4012 29300 4052
rect 30988 4012 31028 4052
rect 4492 3928 4532 3968
rect 4876 3928 4916 3968
rect 7372 3928 7412 3968
rect 11884 3928 11924 3968
rect 22828 3928 22868 3968
rect 23020 3928 23060 3968
rect 23692 3928 23732 3968
rect 23884 3928 23924 3968
rect 27244 3928 27284 3968
rect 29452 3928 29492 3968
rect 32620 3928 32660 3968
rect 33004 3928 33044 3968
rect 36460 3928 36500 3968
rect 36652 3928 36692 3968
rect 38668 3928 38708 3968
rect 40684 3928 40724 3968
rect 41452 3928 41492 3968
rect 4928 3760 4968 3800
rect 5010 3760 5050 3800
rect 5092 3760 5132 3800
rect 5174 3760 5214 3800
rect 5256 3760 5296 3800
rect 20048 3760 20088 3800
rect 20130 3760 20170 3800
rect 20212 3760 20252 3800
rect 20294 3760 20334 3800
rect 20376 3760 20416 3800
rect 35168 3760 35208 3800
rect 35250 3760 35290 3800
rect 35332 3760 35372 3800
rect 35414 3760 35454 3800
rect 35496 3760 35536 3800
rect 4012 3592 4052 3632
rect 10156 3592 10196 3632
rect 12844 3592 12884 3632
rect 15628 3592 15668 3632
rect 21100 3592 21140 3632
rect 22828 3592 22868 3632
rect 29548 3592 29588 3632
rect 3340 3508 3380 3548
rect 7276 3508 7316 3548
rect 7756 3508 7796 3548
rect 18028 3508 18068 3548
rect 24652 3508 24692 3548
rect 26668 3508 26708 3548
rect 31468 3508 31508 3548
rect 33484 3508 33524 3548
rect 35884 3508 35924 3548
rect 37900 3508 37940 3548
rect 1612 3424 1652 3464
rect 2860 3424 2900 3464
rect 3244 3409 3284 3449
rect 3436 3424 3476 3464
rect 3628 3424 3668 3464
rect 3724 3424 3764 3464
rect 3916 3424 3956 3464
rect 4012 3424 4052 3464
rect 4156 3424 4196 3464
rect 4492 3424 4532 3464
rect 4588 3424 4628 3464
rect 4684 3424 4724 3464
rect 4780 3424 4820 3464
rect 4972 3424 5012 3464
rect 5068 3424 5108 3464
rect 5164 3424 5204 3464
rect 5260 3424 5300 3464
rect 5548 3424 5588 3464
rect 5644 3424 5684 3464
rect 6028 3424 6068 3464
rect 6124 3424 6164 3464
rect 6604 3424 6644 3464
rect 7084 3419 7124 3459
rect 7852 3424 7892 3464
rect 8140 3424 8180 3464
rect 8716 3424 8756 3464
rect 9964 3424 10004 3464
rect 11116 3424 11156 3464
rect 11212 3424 11252 3464
rect 12172 3424 12212 3464
rect 12652 3419 12692 3459
rect 14188 3424 14228 3464
rect 15436 3424 15476 3464
rect 16300 3424 16340 3464
rect 16396 3424 16436 3464
rect 16876 3424 16916 3464
rect 17356 3424 17396 3464
rect 17836 3419 17876 3459
rect 19660 3424 19700 3464
rect 20908 3424 20948 3464
rect 21388 3424 21428 3464
rect 22636 3424 22676 3464
rect 23212 3424 23252 3464
rect 24460 3424 24500 3464
rect 24940 3424 24980 3464
rect 25036 3424 25076 3464
rect 25420 3424 25460 3464
rect 25516 3424 25556 3464
rect 25996 3424 26036 3464
rect 26476 3410 26516 3450
rect 28108 3424 28148 3464
rect 29356 3424 29396 3464
rect 30028 3424 30068 3464
rect 31276 3424 31316 3464
rect 31756 3424 31796 3464
rect 31852 3424 31892 3464
rect 32812 3424 32852 3464
rect 33292 3410 33332 3450
rect 34444 3424 34484 3464
rect 35692 3424 35732 3464
rect 36172 3424 36212 3464
rect 36268 3424 36308 3464
rect 36748 3424 36788 3464
rect 37228 3424 37268 3464
rect 37708 3419 37748 3459
rect 38284 3424 38324 3464
rect 39532 3424 39572 3464
rect 11596 3340 11636 3380
rect 11692 3340 11732 3380
rect 16780 3340 16820 3380
rect 32236 3340 32276 3380
rect 32332 3340 32372 3380
rect 36652 3340 36692 3380
rect 39916 3340 39956 3380
rect 40108 3340 40148 3380
rect 40492 3340 40532 3380
rect 40876 3340 40916 3380
rect 41260 3340 41300 3380
rect 3052 3256 3092 3296
rect 38092 3256 38132 3296
rect 41068 3256 41108 3296
rect 7468 3172 7508 3212
rect 39724 3172 39764 3212
rect 40300 3172 40340 3212
rect 40684 3172 40724 3212
rect 41452 3172 41492 3212
rect 3688 3004 3728 3044
rect 3770 3004 3810 3044
rect 3852 3004 3892 3044
rect 3934 3004 3974 3044
rect 4016 3004 4056 3044
rect 18808 3004 18848 3044
rect 18890 3004 18930 3044
rect 18972 3004 19012 3044
rect 19054 3004 19094 3044
rect 19136 3004 19176 3044
rect 33928 3004 33968 3044
rect 34010 3004 34050 3044
rect 34092 3004 34132 3044
rect 34174 3004 34214 3044
rect 34256 3004 34296 3044
rect 2956 2836 2996 2876
rect 4876 2836 4916 2876
rect 27148 2836 27188 2876
rect 20332 2752 20372 2792
rect 24460 2752 24500 2792
rect 32908 2752 32948 2792
rect 41068 2752 41108 2792
rect 11500 2668 11540 2708
rect 14476 2668 14516 2708
rect 20716 2668 20756 2708
rect 20908 2668 20948 2708
rect 21484 2668 21524 2708
rect 22156 2668 22196 2708
rect 22924 2668 22964 2708
rect 23308 2668 23348 2708
rect 24652 2668 24692 2708
rect 25324 2668 25364 2708
rect 32716 2668 32756 2708
rect 35788 2668 35828 2708
rect 36556 2668 36596 2708
rect 38188 2668 38228 2708
rect 38572 2668 38612 2708
rect 40876 2668 40916 2708
rect 41260 2668 41300 2708
rect 1516 2584 1556 2624
rect 2764 2605 2804 2645
rect 3244 2584 3284 2624
rect 3340 2584 3380 2624
rect 3436 2584 3476 2624
rect 3532 2584 3572 2624
rect 3724 2584 3764 2624
rect 3820 2584 3860 2624
rect 4204 2584 4244 2624
rect 4300 2584 4340 2624
rect 4876 2584 4916 2624
rect 5164 2584 5204 2624
rect 5932 2584 5972 2624
rect 7180 2584 7220 2624
rect 7564 2584 7604 2624
rect 8812 2584 8852 2624
rect 9196 2584 9236 2624
rect 10444 2584 10484 2624
rect 10924 2584 10964 2624
rect 11020 2584 11060 2624
rect 11404 2584 11444 2624
rect 11980 2584 12020 2624
rect 12460 2598 12500 2638
rect 13900 2584 13940 2624
rect 13996 2584 14036 2624
rect 14380 2584 14420 2624
rect 14956 2584 14996 2624
rect 15436 2589 15476 2629
rect 15916 2584 15956 2624
rect 17164 2584 17204 2624
rect 17932 2584 17972 2624
rect 19180 2584 19220 2624
rect 19660 2584 19700 2624
rect 19948 2584 19988 2624
rect 23788 2584 23828 2624
rect 24076 2584 24116 2624
rect 24172 2584 24212 2624
rect 25708 2584 25748 2624
rect 26956 2584 26996 2624
rect 27532 2584 27572 2624
rect 28780 2584 28820 2624
rect 29164 2584 29204 2624
rect 30412 2584 30452 2624
rect 30796 2584 30836 2624
rect 32044 2584 32084 2624
rect 33100 2584 33140 2624
rect 34348 2584 34388 2624
rect 36076 2584 36116 2624
rect 36172 2584 36212 2624
rect 36652 2584 36692 2624
rect 37132 2584 37172 2624
rect 37612 2589 37652 2629
rect 39148 2584 39188 2624
rect 40396 2584 40436 2624
rect 15628 2500 15668 2540
rect 19372 2500 19412 2540
rect 20044 2500 20084 2540
rect 37804 2500 37844 2540
rect 38956 2500 38996 2540
rect 4012 2416 4052 2456
rect 4492 2416 4532 2456
rect 7372 2416 7412 2456
rect 9004 2416 9044 2456
rect 10636 2416 10676 2456
rect 12652 2416 12692 2456
rect 17356 2416 17396 2456
rect 20524 2416 20564 2456
rect 21100 2416 21140 2456
rect 21676 2416 21716 2456
rect 21964 2416 22004 2456
rect 23116 2416 23156 2456
rect 23500 2416 23540 2456
rect 24844 2416 24884 2456
rect 25516 2416 25556 2456
rect 27340 2416 27380 2456
rect 28972 2416 29012 2456
rect 30604 2416 30644 2456
rect 32524 2416 32564 2456
rect 35596 2416 35636 2456
rect 37996 2416 38036 2456
rect 38764 2416 38804 2456
rect 41452 2416 41492 2456
rect 4928 2248 4968 2288
rect 5010 2248 5050 2288
rect 5092 2248 5132 2288
rect 5174 2248 5214 2288
rect 5256 2248 5296 2288
rect 20048 2248 20088 2288
rect 20130 2248 20170 2288
rect 20212 2248 20252 2288
rect 20294 2248 20334 2288
rect 20376 2248 20416 2288
rect 35168 2248 35208 2288
rect 35250 2248 35290 2288
rect 35332 2248 35372 2288
rect 35414 2248 35454 2288
rect 35496 2248 35536 2288
rect 14860 2080 14900 2120
rect 16876 2080 16916 2120
rect 19180 2080 19220 2120
rect 22060 2080 22100 2120
rect 37036 2080 37076 2120
rect 40204 2080 40244 2120
rect 5260 1996 5300 2036
rect 7276 1996 7316 2036
rect 9580 1996 9620 2036
rect 12844 1996 12884 2036
rect 23884 1996 23924 2036
rect 26476 1996 26516 2036
rect 29452 1996 29492 2036
rect 32236 1996 32276 2036
rect 40012 1996 40052 2036
rect 2188 1912 2228 1952
rect 3436 1912 3476 1952
rect 3820 1912 3860 1952
rect 5068 1912 5108 1952
rect 5548 1912 5588 1952
rect 5644 1912 5684 1952
rect 6028 1912 6068 1952
rect 6604 1912 6644 1952
rect 7084 1907 7124 1947
rect 7852 1912 7892 1952
rect 7948 1912 7988 1952
rect 8332 1912 8372 1952
rect 8908 1912 8948 1952
rect 9388 1907 9428 1947
rect 11116 1912 11156 1952
rect 11212 1912 11252 1952
rect 12172 1912 12212 1952
rect 12652 1907 12692 1947
rect 13420 1912 13460 1952
rect 14668 1912 14708 1952
rect 15148 1912 15188 1952
rect 15244 1912 15284 1952
rect 16204 1912 16244 1952
rect 16684 1898 16724 1938
rect 17452 1912 17492 1952
rect 17548 1912 17588 1952
rect 18508 1912 18548 1952
rect 18988 1898 19028 1938
rect 20332 1912 20372 1952
rect 20428 1912 20468 1952
rect 21388 1912 21428 1952
rect 21868 1898 21908 1938
rect 22444 1912 22484 1952
rect 23692 1912 23732 1952
rect 24748 1912 24788 1952
rect 24844 1912 24884 1952
rect 25324 1912 25364 1952
rect 25804 1912 25844 1952
rect 26284 1898 26324 1938
rect 27724 1912 27764 1952
rect 27820 1912 27860 1952
rect 28780 1912 28820 1952
rect 29260 1907 29300 1947
rect 30508 1893 30548 1933
rect 30604 1893 30644 1933
rect 31084 1912 31124 1952
rect 31564 1912 31604 1952
rect 32044 1898 32084 1938
rect 33004 1912 33044 1952
rect 34252 1912 34292 1952
rect 35308 1912 35348 1952
rect 35404 1912 35444 1952
rect 35788 1912 35828 1952
rect 36364 1912 36404 1952
rect 36844 1898 36884 1938
rect 38284 1912 38324 1952
rect 38380 1912 38420 1952
rect 38764 1912 38804 1952
rect 38860 1912 38900 1952
rect 39340 1912 39380 1952
rect 39820 1902 39860 1942
rect 40396 1912 40436 1952
rect 41644 1912 41684 1952
rect 6124 1828 6164 1868
rect 8428 1828 8468 1868
rect 10636 1828 10676 1868
rect 11596 1828 11636 1868
rect 11692 1828 11732 1868
rect 13036 1828 13076 1868
rect 15628 1828 15668 1868
rect 15724 1828 15764 1868
rect 17932 1828 17972 1868
rect 18028 1828 18068 1868
rect 19852 1828 19892 1868
rect 20812 1828 20852 1868
rect 20908 1828 20948 1868
rect 24268 1828 24308 1868
rect 25228 1828 25268 1868
rect 26860 1828 26900 1868
rect 27244 1828 27284 1868
rect 28204 1828 28244 1868
rect 28300 1828 28340 1868
rect 29836 1841 29876 1881
rect 30220 1828 30260 1868
rect 30988 1828 31028 1868
rect 32620 1828 32660 1868
rect 34636 1828 34676 1868
rect 35884 1828 35924 1868
rect 37708 1828 37748 1868
rect 3628 1660 3668 1700
rect 10828 1660 10868 1700
rect 13228 1660 13268 1700
rect 20044 1660 20084 1700
rect 24076 1660 24116 1700
rect 26668 1660 26708 1700
rect 27436 1660 27476 1700
rect 29644 1660 29684 1700
rect 30028 1660 30068 1700
rect 32428 1660 32468 1700
rect 32812 1660 32852 1700
rect 34444 1660 34484 1700
rect 37516 1660 37556 1700
rect 3688 1492 3728 1532
rect 3770 1492 3810 1532
rect 3852 1492 3892 1532
rect 3934 1492 3974 1532
rect 4016 1492 4056 1532
rect 18808 1492 18848 1532
rect 18890 1492 18930 1532
rect 18972 1492 19012 1532
rect 19054 1492 19094 1532
rect 19136 1492 19176 1532
rect 33928 1492 33968 1532
rect 34010 1492 34050 1532
rect 34092 1492 34132 1532
rect 34174 1492 34214 1532
rect 34256 1492 34296 1532
rect 10540 1324 10580 1364
rect 16684 1324 16724 1364
rect 20428 1324 20468 1364
rect 22156 1324 22196 1364
rect 24940 1324 24980 1364
rect 25612 1324 25652 1364
rect 30604 1324 30644 1364
rect 38092 1324 38132 1364
rect 12172 1240 12212 1280
rect 13804 1240 13844 1280
rect 18796 1240 18836 1280
rect 33196 1240 33236 1280
rect 34828 1240 34868 1280
rect 36460 1240 36500 1280
rect 41068 1240 41108 1280
rect 5740 1156 5780 1196
rect 5836 1156 5876 1196
rect 22924 1156 22964 1196
rect 28492 1156 28532 1196
rect 30988 1156 31028 1196
rect 31756 1156 31796 1196
rect 1324 1072 1364 1112
rect 2572 1072 2612 1112
rect 3052 1072 3092 1112
rect 4300 1072 4340 1112
rect 5260 1072 5300 1112
rect 5356 1072 5396 1112
rect 6316 1072 6356 1112
rect 6796 1086 6836 1126
rect 25804 1114 25844 1154
rect 31852 1156 31892 1196
rect 39916 1156 39956 1196
rect 40108 1156 40148 1196
rect 40492 1156 40532 1196
rect 40876 1156 40916 1196
rect 41260 1156 41300 1196
rect 9100 1072 9140 1112
rect 10348 1072 10388 1112
rect 10732 1072 10772 1112
rect 11980 1072 12020 1112
rect 12364 1072 12404 1112
rect 13612 1072 13652 1112
rect 15244 1072 15284 1112
rect 16492 1072 16532 1112
rect 17356 1072 17396 1112
rect 18604 1072 18644 1112
rect 18988 1072 19028 1112
rect 20236 1072 20276 1112
rect 20716 1072 20756 1112
rect 21964 1072 22004 1112
rect 24748 1072 24788 1112
rect 27052 1072 27092 1112
rect 29164 1072 29204 1112
rect 30412 1072 30452 1112
rect 31276 1072 31316 1112
rect 23500 1030 23540 1070
rect 31372 1072 31412 1112
rect 32332 1072 32372 1112
rect 32812 1086 32852 1126
rect 33388 1072 33428 1112
rect 34636 1072 34676 1112
rect 35020 1072 35060 1112
rect 36268 1072 36308 1112
rect 36652 1072 36692 1112
rect 37900 1072 37940 1112
rect 38284 1072 38324 1112
rect 39532 1072 39572 1112
rect 4492 988 4532 1028
rect 33004 988 33044 1028
rect 2764 904 2804 944
rect 6988 904 7028 944
rect 23116 904 23156 944
rect 28684 904 28724 944
rect 30796 904 30836 944
rect 39724 904 39764 944
rect 40300 904 40340 944
rect 40684 904 40724 944
rect 41452 904 41492 944
rect 4928 736 4968 776
rect 5010 736 5050 776
rect 5092 736 5132 776
rect 5174 736 5214 776
rect 5256 736 5296 776
rect 20048 736 20088 776
rect 20130 736 20170 776
rect 20212 736 20252 776
rect 20294 736 20334 776
rect 20376 736 20416 776
rect 35168 736 35208 776
rect 35250 736 35290 776
rect 35332 736 35372 776
rect 35414 736 35454 776
rect 35496 736 35536 776
<< metal2 >>
rect 1784 10672 1864 10752
rect 2936 10672 3016 10752
rect 4088 10732 4168 10752
rect 4088 10692 4628 10732
rect 4088 10672 4196 10692
rect 1804 10604 1844 10672
rect 1804 10564 2036 10604
rect 555 10184 597 10193
rect 555 10144 556 10184
rect 596 10144 597 10184
rect 555 10135 597 10144
rect 556 7673 596 10135
rect 1516 9512 1556 9521
rect 1227 9176 1269 9185
rect 1227 9136 1228 9176
rect 1268 9136 1269 9176
rect 1227 9127 1269 9136
rect 1228 8009 1268 9127
rect 1516 8177 1556 9472
rect 1803 8840 1845 8849
rect 1803 8800 1804 8840
rect 1844 8800 1845 8840
rect 1803 8791 1845 8800
rect 1612 8672 1652 8681
rect 1515 8168 1557 8177
rect 1515 8128 1516 8168
rect 1556 8128 1557 8168
rect 1515 8119 1557 8128
rect 1227 8000 1269 8009
rect 1227 7960 1228 8000
rect 1268 7960 1269 8000
rect 1227 7951 1269 7960
rect 1420 8000 1460 8009
rect 1420 7841 1460 7960
rect 1419 7832 1461 7841
rect 1419 7792 1420 7832
rect 1460 7792 1461 7832
rect 1419 7783 1461 7792
rect 555 7664 597 7673
rect 555 7624 556 7664
rect 596 7624 597 7664
rect 555 7615 597 7624
rect 1612 7505 1652 8632
rect 1707 8504 1749 8513
rect 1707 8464 1708 8504
rect 1748 8464 1749 8504
rect 1707 8455 1749 8464
rect 1611 7496 1653 7505
rect 1611 7456 1612 7496
rect 1652 7456 1653 7496
rect 1611 7447 1653 7456
rect 1419 6824 1461 6833
rect 1419 6784 1420 6824
rect 1460 6784 1461 6824
rect 1419 6775 1461 6784
rect 1323 6152 1365 6161
rect 1323 6112 1324 6152
rect 1364 6112 1365 6152
rect 1323 6103 1365 6112
rect 1227 5984 1269 5993
rect 1227 5944 1228 5984
rect 1268 5944 1269 5984
rect 1227 5935 1269 5944
rect 1035 5816 1077 5825
rect 1035 5776 1036 5816
rect 1076 5776 1077 5816
rect 1035 5767 1077 5776
rect 1036 3221 1076 5767
rect 1131 5228 1173 5237
rect 1131 5188 1132 5228
rect 1172 5188 1173 5228
rect 1131 5179 1173 5188
rect 1035 3212 1077 3221
rect 1035 3172 1036 3212
rect 1076 3172 1077 3212
rect 1035 3163 1077 3172
rect 1132 2801 1172 5179
rect 1228 3473 1268 5935
rect 1324 5069 1364 6103
rect 1323 5060 1365 5069
rect 1323 5020 1324 5060
rect 1364 5020 1365 5060
rect 1323 5011 1365 5020
rect 1227 3464 1269 3473
rect 1227 3424 1228 3464
rect 1268 3424 1269 3464
rect 1227 3415 1269 3424
rect 1420 3044 1460 6775
rect 1708 6497 1748 8455
rect 1515 6488 1557 6497
rect 1515 6448 1516 6488
rect 1556 6448 1557 6488
rect 1515 6439 1557 6448
rect 1707 6488 1749 6497
rect 1707 6448 1708 6488
rect 1748 6448 1749 6488
rect 1707 6439 1749 6448
rect 1516 4976 1556 6439
rect 1708 6354 1748 6439
rect 1612 5648 1652 5657
rect 1804 5648 1844 8791
rect 1899 7160 1941 7169
rect 1899 7120 1900 7160
rect 1940 7120 1941 7160
rect 1899 7111 1941 7120
rect 1652 5608 1844 5648
rect 1612 5599 1652 5608
rect 1707 5060 1749 5069
rect 1707 5020 1708 5060
rect 1748 5020 1749 5060
rect 1707 5011 1749 5020
rect 1611 4976 1653 4985
rect 1516 4936 1612 4976
rect 1652 4936 1653 4976
rect 1611 4927 1653 4936
rect 1612 4842 1652 4927
rect 1516 4136 1556 4145
rect 1708 4136 1748 5011
rect 1556 4096 1748 4136
rect 1516 4087 1556 4096
rect 1900 3473 1940 7111
rect 1996 4649 2036 10564
rect 2956 9764 2996 10672
rect 4108 10648 4196 10672
rect 2956 9724 3284 9764
rect 2955 9596 2997 9605
rect 2955 9556 2956 9596
rect 2996 9556 2997 9596
rect 2955 9547 2997 9556
rect 2764 9512 2804 9521
rect 2668 9472 2764 9512
rect 2668 8681 2708 9472
rect 2764 9463 2804 9472
rect 2667 8672 2709 8681
rect 2667 8632 2668 8672
rect 2708 8632 2709 8672
rect 2667 8623 2709 8632
rect 2859 8672 2901 8681
rect 2859 8632 2860 8672
rect 2900 8632 2901 8672
rect 2859 8623 2901 8632
rect 2668 8177 2708 8623
rect 2860 8538 2900 8623
rect 2859 8252 2901 8261
rect 2859 8212 2860 8252
rect 2900 8212 2901 8252
rect 2859 8203 2901 8212
rect 2667 8168 2709 8177
rect 2667 8128 2668 8168
rect 2708 8128 2709 8168
rect 2667 8119 2709 8128
rect 2860 8168 2900 8203
rect 2668 8000 2708 8119
rect 2860 8117 2900 8128
rect 2956 8000 2996 9547
rect 3051 8588 3093 8597
rect 3051 8548 3052 8588
rect 3092 8548 3093 8588
rect 3051 8539 3093 8548
rect 3052 8454 3092 8539
rect 3052 8000 3092 8009
rect 2956 7960 3052 8000
rect 2668 6497 2708 7960
rect 2860 7748 2900 7757
rect 2860 6992 2900 7708
rect 3052 7664 3092 7960
rect 3147 7916 3189 7925
rect 3147 7876 3148 7916
rect 3188 7876 3189 7916
rect 3147 7867 3189 7876
rect 3148 7782 3188 7867
rect 3052 7624 3188 7664
rect 2955 7328 2997 7337
rect 2955 7288 2956 7328
rect 2996 7288 2997 7328
rect 2955 7279 2997 7288
rect 2956 7160 2996 7279
rect 2956 7111 2996 7120
rect 3052 7160 3092 7169
rect 3052 6992 3092 7120
rect 2860 6952 3092 6992
rect 3148 7160 3188 7624
rect 3244 7328 3284 9724
rect 4108 9680 4148 9689
rect 3915 9596 3957 9605
rect 3915 9556 3916 9596
rect 3956 9556 3957 9596
rect 3915 9547 3957 9556
rect 3340 9512 3380 9521
rect 3340 8681 3380 9472
rect 3436 9512 3476 9521
rect 3436 8933 3476 9472
rect 3532 9512 3572 9521
rect 3435 8924 3477 8933
rect 3435 8884 3436 8924
rect 3476 8884 3477 8924
rect 3532 8924 3572 9472
rect 3627 9512 3669 9521
rect 3627 9472 3628 9512
rect 3668 9472 3669 9512
rect 3627 9463 3669 9472
rect 3820 9512 3860 9521
rect 3628 9378 3668 9463
rect 3820 9353 3860 9472
rect 3916 9512 3956 9547
rect 3916 9461 3956 9472
rect 3819 9344 3861 9353
rect 3819 9304 3820 9344
rect 3860 9304 3861 9344
rect 3819 9295 3861 9304
rect 3688 9092 4056 9101
rect 3728 9052 3770 9092
rect 3810 9052 3852 9092
rect 3892 9052 3934 9092
rect 3974 9052 4016 9092
rect 3688 9043 4056 9052
rect 3628 8924 3668 8933
rect 3532 8884 3628 8924
rect 3435 8875 3477 8884
rect 3628 8875 3668 8884
rect 4011 8924 4053 8933
rect 4011 8884 4012 8924
rect 4052 8884 4053 8924
rect 4011 8875 4053 8884
rect 3339 8672 3381 8681
rect 3339 8632 3340 8672
rect 3380 8632 3381 8672
rect 3339 8623 3381 8632
rect 3532 8672 3572 8681
rect 3340 8261 3380 8623
rect 3339 8252 3381 8261
rect 3339 8212 3340 8252
rect 3380 8212 3381 8252
rect 3339 8203 3381 8212
rect 3340 8000 3380 8203
rect 3532 8168 3572 8632
rect 3627 8672 3669 8681
rect 3627 8632 3628 8672
rect 3668 8632 3669 8672
rect 3627 8623 3669 8632
rect 3820 8672 3860 8681
rect 3628 8538 3668 8623
rect 3820 8429 3860 8632
rect 4012 8672 4052 8875
rect 4012 8623 4052 8632
rect 4108 8672 4148 9640
rect 4588 9680 4628 10692
rect 5240 10672 5320 10752
rect 6392 10672 6472 10752
rect 7544 10672 7624 10752
rect 8696 10672 8776 10752
rect 8908 10692 9236 10732
rect 5260 10613 5300 10672
rect 5259 10604 5301 10613
rect 5259 10564 5260 10604
rect 5300 10564 5301 10604
rect 5259 10555 5301 10564
rect 4928 9848 5296 9857
rect 4968 9808 5010 9848
rect 5050 9808 5092 9848
rect 5132 9808 5174 9848
rect 5214 9808 5256 9848
rect 4928 9799 5296 9808
rect 5931 9764 5973 9773
rect 5931 9724 5932 9764
rect 5972 9724 5973 9764
rect 5931 9715 5973 9724
rect 4588 9631 4628 9640
rect 4203 9596 4245 9605
rect 4203 9556 4204 9596
rect 4244 9556 4245 9596
rect 4203 9547 4245 9556
rect 4108 8623 4148 8632
rect 4204 8672 4244 9547
rect 4300 9512 4340 9521
rect 4300 8840 4340 9472
rect 4395 9512 4437 9521
rect 4395 9472 4396 9512
rect 4436 9472 4437 9512
rect 4395 9463 4437 9472
rect 4492 9512 4532 9521
rect 4396 9378 4436 9463
rect 4300 8800 4436 8840
rect 4204 8623 4244 8632
rect 4300 8672 4340 8681
rect 4203 8504 4245 8513
rect 4203 8464 4204 8504
rect 4244 8464 4245 8504
rect 4203 8455 4245 8464
rect 3819 8420 3861 8429
rect 3819 8380 3820 8420
rect 3860 8380 3861 8420
rect 3819 8371 3861 8380
rect 3532 8128 3668 8168
rect 3436 8000 3476 8009
rect 3340 7960 3436 8000
rect 3436 7951 3476 7960
rect 3532 8000 3572 8009
rect 3532 7832 3572 7960
rect 3628 8000 3668 8128
rect 3628 7925 3668 7960
rect 4011 8000 4053 8009
rect 4011 7960 4012 8000
rect 4052 7960 4053 8000
rect 4011 7951 4053 7960
rect 3627 7916 3669 7925
rect 3627 7876 3628 7916
rect 3668 7876 3669 7916
rect 3627 7867 3669 7876
rect 4012 7866 4052 7951
rect 3436 7792 3572 7832
rect 3436 7505 3476 7792
rect 3820 7748 3860 7757
rect 3532 7708 3820 7748
rect 3435 7496 3477 7505
rect 3435 7456 3436 7496
rect 3476 7456 3477 7496
rect 3435 7447 3477 7456
rect 3532 7412 3572 7708
rect 3820 7699 3860 7708
rect 4107 7748 4149 7757
rect 4107 7708 4108 7748
rect 4148 7708 4149 7748
rect 4107 7699 4149 7708
rect 3688 7580 4056 7589
rect 3728 7540 3770 7580
rect 3810 7540 3852 7580
rect 3892 7540 3934 7580
rect 3974 7540 4016 7580
rect 3688 7531 4056 7540
rect 3724 7412 3764 7421
rect 4108 7412 4148 7699
rect 3532 7372 3668 7412
rect 3435 7328 3477 7337
rect 3244 7288 3380 7328
rect 3148 6665 3188 7120
rect 3243 7160 3285 7169
rect 3243 7120 3244 7160
rect 3284 7120 3285 7160
rect 3243 7111 3285 7120
rect 3244 7026 3284 7111
rect 3340 6740 3380 7288
rect 3435 7288 3436 7328
rect 3476 7288 3572 7328
rect 3435 7279 3477 7288
rect 3243 6700 3380 6740
rect 3436 7160 3476 7169
rect 3147 6656 3189 6665
rect 3147 6616 3148 6656
rect 3188 6616 3189 6656
rect 3243 6656 3283 6700
rect 3436 6656 3476 7120
rect 3532 7160 3572 7288
rect 3532 7111 3572 7120
rect 3628 7076 3668 7372
rect 3764 7372 4148 7412
rect 3724 7363 3764 7372
rect 4204 7328 4244 8455
rect 4300 7589 4340 8632
rect 4396 8597 4436 8800
rect 4395 8588 4437 8597
rect 4395 8548 4396 8588
rect 4436 8548 4437 8588
rect 4395 8539 4437 8548
rect 4395 8420 4437 8429
rect 4395 8380 4396 8420
rect 4436 8380 4437 8420
rect 4395 8371 4437 8380
rect 4299 7580 4341 7589
rect 4299 7540 4300 7580
rect 4340 7540 4341 7580
rect 4396 7580 4436 8371
rect 4492 7757 4532 9472
rect 5355 8756 5397 8765
rect 5355 8716 5356 8756
rect 5396 8716 5397 8756
rect 5355 8707 5397 8716
rect 4780 8672 4820 8681
rect 4780 8513 4820 8632
rect 4779 8504 4821 8513
rect 4779 8464 4780 8504
rect 4820 8464 4821 8504
rect 4779 8455 4821 8464
rect 4928 8336 5296 8345
rect 4968 8296 5010 8336
rect 5050 8296 5092 8336
rect 5132 8296 5174 8336
rect 5214 8296 5256 8336
rect 4928 8287 5296 8296
rect 5356 8177 5396 8707
rect 5932 8177 5972 9715
rect 6412 8840 6452 10672
rect 6316 8800 6452 8840
rect 6027 8756 6069 8765
rect 6027 8716 6028 8756
rect 6068 8716 6069 8756
rect 6027 8707 6069 8716
rect 6028 8672 6068 8707
rect 6028 8621 6068 8632
rect 6220 8504 6260 8513
rect 5355 8168 5397 8177
rect 5355 8128 5356 8168
rect 5396 8128 5397 8168
rect 5355 8119 5397 8128
rect 5931 8168 5973 8177
rect 5931 8128 5932 8168
rect 5972 8128 5973 8168
rect 5931 8119 5973 8128
rect 5260 8000 5300 8009
rect 5356 8000 5396 8119
rect 5300 7960 5396 8000
rect 5932 8000 5972 8119
rect 5260 7951 5300 7960
rect 5932 7951 5972 7960
rect 4491 7748 4533 7757
rect 4491 7708 4492 7748
rect 4532 7708 4533 7748
rect 4491 7699 4533 7708
rect 5452 7748 5492 7757
rect 4396 7540 4532 7580
rect 4299 7531 4341 7540
rect 4395 7412 4437 7421
rect 4395 7372 4396 7412
rect 4436 7372 4437 7412
rect 4395 7363 4437 7372
rect 3820 7288 4244 7328
rect 4396 7328 4436 7363
rect 3820 7244 3860 7288
rect 4396 7277 4436 7288
rect 3628 7027 3668 7036
rect 3724 7204 3860 7244
rect 3724 6992 3764 7204
rect 4203 7160 4245 7169
rect 4203 7120 4204 7160
rect 4244 7120 4245 7160
rect 4203 7111 4245 7120
rect 4396 7152 4436 7161
rect 3724 6943 3764 6952
rect 3627 6908 3669 6917
rect 3627 6868 3628 6908
rect 3668 6868 3669 6908
rect 3627 6859 3669 6868
rect 3243 6616 3284 6656
rect 3436 6616 3572 6656
rect 3147 6607 3189 6616
rect 2667 6488 2709 6497
rect 2955 6488 2997 6497
rect 2667 6448 2668 6488
rect 2708 6448 2709 6488
rect 2667 6439 2709 6448
rect 2860 6448 2956 6488
rect 2996 6448 2997 6488
rect 2475 5816 2517 5825
rect 2475 5776 2476 5816
rect 2516 5776 2517 5816
rect 2475 5767 2517 5776
rect 2283 5396 2325 5405
rect 2283 5356 2284 5396
rect 2324 5356 2325 5396
rect 2283 5347 2325 5356
rect 1995 4640 2037 4649
rect 1995 4600 1996 4640
rect 2036 4600 2037 4640
rect 1995 4591 2037 4600
rect 2187 4220 2229 4229
rect 2187 4180 2188 4220
rect 2228 4180 2229 4220
rect 2187 4171 2229 4180
rect 1611 3464 1653 3473
rect 1611 3424 1612 3464
rect 1652 3424 1653 3464
rect 1611 3415 1653 3424
rect 1899 3464 1941 3473
rect 1899 3424 1900 3464
rect 1940 3424 1941 3464
rect 1899 3415 1941 3424
rect 1612 3330 1652 3415
rect 1515 3044 1557 3053
rect 1420 3004 1516 3044
rect 1556 3004 1557 3044
rect 1515 2995 1557 3004
rect 1131 2792 1173 2801
rect 1131 2752 1132 2792
rect 1172 2752 1173 2792
rect 1131 2743 1173 2752
rect 1516 2624 1556 2995
rect 1516 2575 1556 2584
rect 2188 1952 2228 4171
rect 2284 3137 2324 5347
rect 2379 4808 2421 4817
rect 2379 4768 2380 4808
rect 2420 4768 2421 4808
rect 2379 4759 2421 4768
rect 2380 4229 2420 4759
rect 2379 4220 2421 4229
rect 2379 4180 2380 4220
rect 2420 4180 2421 4220
rect 2379 4171 2421 4180
rect 2476 3809 2516 5767
rect 2860 5648 2900 6448
rect 2955 6439 2997 6448
rect 3147 6488 3189 6497
rect 3147 6448 3148 6488
rect 3188 6448 3189 6488
rect 3147 6439 3189 6448
rect 2956 6354 2996 6439
rect 3148 6320 3188 6439
rect 3148 6271 3188 6280
rect 3244 5900 3284 6616
rect 3339 6572 3381 6581
rect 3532 6572 3572 6616
rect 3339 6532 3340 6572
rect 3380 6532 3476 6572
rect 3339 6523 3381 6532
rect 3436 6488 3476 6532
rect 3532 6523 3572 6532
rect 3436 6439 3476 6448
rect 3628 6488 3668 6859
rect 3628 6439 3668 6448
rect 3915 6488 3957 6497
rect 3915 6448 3916 6488
rect 3956 6448 3957 6488
rect 3915 6439 3957 6448
rect 4204 6488 4244 7111
rect 4396 7085 4436 7112
rect 4395 7076 4437 7085
rect 4395 7036 4396 7076
rect 4436 7036 4437 7076
rect 4395 7027 4437 7036
rect 4300 6497 4340 6582
rect 3916 6354 3956 6439
rect 4204 6245 4244 6448
rect 4299 6488 4341 6497
rect 4299 6448 4300 6488
rect 4340 6448 4341 6488
rect 4299 6439 4341 6448
rect 4299 6320 4341 6329
rect 4396 6320 4436 7027
rect 4492 6413 4532 7540
rect 5452 7505 5492 7708
rect 5163 7496 5205 7505
rect 5163 7456 5164 7496
rect 5204 7456 5205 7496
rect 5163 7447 5205 7456
rect 5451 7496 5493 7505
rect 5451 7456 5452 7496
rect 5492 7456 5493 7496
rect 5451 7447 5493 7456
rect 6027 7496 6069 7505
rect 6027 7456 6028 7496
rect 6068 7456 6069 7496
rect 6027 7447 6069 7456
rect 5164 7253 5204 7447
rect 5355 7328 5397 7337
rect 5355 7288 5356 7328
rect 5396 7288 5397 7328
rect 5355 7279 5397 7288
rect 5548 7288 5876 7328
rect 5163 7244 5205 7253
rect 5163 7204 5164 7244
rect 5204 7204 5205 7244
rect 5163 7195 5205 7204
rect 4780 7160 4820 7171
rect 5260 7169 5300 7254
rect 4780 7085 4820 7120
rect 4876 7160 4916 7169
rect 4779 7076 4821 7085
rect 4779 7036 4780 7076
rect 4820 7036 4821 7076
rect 4779 7027 4821 7036
rect 4876 7001 4916 7120
rect 5259 7160 5301 7169
rect 5259 7120 5260 7160
rect 5300 7120 5301 7160
rect 5259 7111 5301 7120
rect 5356 7160 5396 7279
rect 5452 7169 5492 7254
rect 5356 7111 5396 7120
rect 5451 7160 5493 7169
rect 5451 7120 5452 7160
rect 5492 7120 5493 7160
rect 5451 7111 5493 7120
rect 5548 7160 5588 7288
rect 5548 7111 5588 7120
rect 5740 7160 5780 7169
rect 4588 6992 4628 7001
rect 4588 6497 4628 6952
rect 4875 6992 4917 7001
rect 4875 6952 4876 6992
rect 4916 6952 4917 6992
rect 4875 6943 4917 6952
rect 5068 6992 5108 7001
rect 5451 6992 5493 7001
rect 5108 6952 5396 6992
rect 5068 6943 5108 6952
rect 4928 6824 5296 6833
rect 4968 6784 5010 6824
rect 5050 6784 5092 6824
rect 5132 6784 5174 6824
rect 5214 6784 5256 6824
rect 4928 6775 5296 6784
rect 5356 6656 5396 6952
rect 5451 6952 5452 6992
rect 5492 6952 5493 6992
rect 5451 6943 5493 6952
rect 5164 6616 5396 6656
rect 5068 6497 5108 6582
rect 4587 6488 4629 6497
rect 4587 6448 4588 6488
rect 4628 6448 4629 6488
rect 4587 6439 4629 6448
rect 4871 6488 4911 6497
rect 4491 6404 4533 6413
rect 4491 6364 4492 6404
rect 4532 6364 4533 6404
rect 4491 6355 4533 6364
rect 4299 6280 4300 6320
rect 4340 6280 4436 6320
rect 4299 6271 4341 6280
rect 4203 6236 4245 6245
rect 4203 6196 4204 6236
rect 4244 6196 4245 6236
rect 4203 6187 4245 6196
rect 3688 6068 4056 6077
rect 3728 6028 3770 6068
rect 3810 6028 3852 6068
rect 3892 6028 3934 6068
rect 3974 6028 4016 6068
rect 3688 6019 4056 6028
rect 4108 5909 4148 5994
rect 4107 5900 4149 5909
rect 3244 5860 3668 5900
rect 2667 5144 2709 5153
rect 2667 5104 2668 5144
rect 2708 5104 2709 5144
rect 2667 5095 2709 5104
rect 2475 3800 2517 3809
rect 2475 3760 2476 3800
rect 2516 3760 2517 3800
rect 2475 3751 2517 3760
rect 2283 3128 2325 3137
rect 2283 3088 2284 3128
rect 2324 3088 2325 3128
rect 2283 3079 2325 3088
rect 2668 2540 2708 5095
rect 2860 4976 2900 5608
rect 3051 5648 3093 5657
rect 3051 5608 3052 5648
rect 3092 5608 3093 5648
rect 3051 5599 3093 5608
rect 3052 5564 3092 5599
rect 3052 5513 3092 5524
rect 3628 5060 3668 5860
rect 4107 5860 4108 5900
rect 4148 5860 4149 5900
rect 4107 5851 4149 5860
rect 4300 5816 4340 6271
rect 4492 6152 4532 6355
rect 4588 6320 4628 6329
rect 4588 6236 4628 6280
rect 4871 6236 4911 6448
rect 4588 6196 4911 6236
rect 4972 6488 5012 6497
rect 4492 6112 4724 6152
rect 4300 5776 4532 5816
rect 4107 5648 4149 5657
rect 4107 5608 4108 5648
rect 4148 5608 4149 5648
rect 4107 5599 4149 5608
rect 4300 5648 4340 5776
rect 4492 5732 4532 5776
rect 4492 5692 4628 5732
rect 4300 5599 4340 5608
rect 4396 5648 4436 5657
rect 4588 5648 4628 5692
rect 4436 5608 4532 5648
rect 4396 5599 4436 5608
rect 4108 5514 4148 5599
rect 4299 5312 4341 5321
rect 4299 5272 4300 5312
rect 4340 5272 4341 5312
rect 4299 5263 4341 5272
rect 3915 5144 3957 5153
rect 3915 5104 3916 5144
rect 3956 5104 3957 5144
rect 3915 5095 3957 5104
rect 4204 5144 4244 5153
rect 4300 5144 4340 5263
rect 4244 5104 4340 5144
rect 4492 5144 4532 5608
rect 4588 5599 4628 5608
rect 4588 5144 4628 5153
rect 4492 5104 4588 5144
rect 4204 5095 4244 5104
rect 4588 5095 4628 5104
rect 3628 5011 3668 5020
rect 2764 4936 2860 4976
rect 2764 4136 2804 4936
rect 2860 4927 2900 4936
rect 3724 4976 3764 4985
rect 3051 4808 3093 4817
rect 3051 4768 3052 4808
rect 3092 4768 3093 4808
rect 3051 4759 3093 4768
rect 3339 4808 3381 4817
rect 3339 4768 3340 4808
rect 3380 4768 3381 4808
rect 3339 4759 3381 4768
rect 3052 4674 3092 4759
rect 3243 4472 3285 4481
rect 3243 4432 3244 4472
rect 3284 4432 3285 4472
rect 3243 4423 3285 4432
rect 2764 3464 2804 4096
rect 2955 4052 2997 4061
rect 2955 4012 2956 4052
rect 2996 4012 2997 4052
rect 2955 4003 2997 4012
rect 3147 4052 3189 4061
rect 3147 4012 3148 4052
rect 3188 4012 3189 4052
rect 3147 4003 3189 4012
rect 2956 3918 2996 4003
rect 2860 3464 2900 3473
rect 2764 3424 2860 3464
rect 3148 3464 3188 4003
rect 3244 3632 3284 4423
rect 3340 3809 3380 4759
rect 3724 4724 3764 4936
rect 3820 4976 3860 4985
rect 3820 4817 3860 4936
rect 3916 4976 3956 5095
rect 4108 4985 4148 5070
rect 3916 4927 3956 4936
rect 4107 4976 4149 4985
rect 4107 4936 4108 4976
rect 4148 4936 4149 4976
rect 4107 4927 4149 4936
rect 4300 4976 4340 4985
rect 3819 4808 3861 4817
rect 3819 4768 3820 4808
rect 3860 4768 3861 4808
rect 3819 4759 3861 4768
rect 3436 4684 3764 4724
rect 3339 3800 3381 3809
rect 3339 3760 3340 3800
rect 3380 3760 3381 3800
rect 3339 3751 3381 3760
rect 3436 3716 3476 4684
rect 3688 4556 4056 4565
rect 3728 4516 3770 4556
rect 3810 4516 3852 4556
rect 3892 4516 3934 4556
rect 3974 4516 4016 4556
rect 3688 4507 4056 4516
rect 4300 4481 4340 4936
rect 4396 4976 4436 4985
rect 4299 4472 4341 4481
rect 4299 4432 4300 4472
rect 4340 4432 4341 4472
rect 4299 4423 4341 4432
rect 3915 4388 3957 4397
rect 3915 4348 3916 4388
rect 3956 4348 3957 4388
rect 3915 4339 3957 4348
rect 3532 4136 3572 4147
rect 3532 4061 3572 4096
rect 3819 4136 3861 4145
rect 3819 4096 3820 4136
rect 3860 4096 3861 4136
rect 3819 4087 3861 4096
rect 3916 4136 3956 4339
rect 3916 4087 3956 4096
rect 4204 4304 4244 4313
rect 4396 4304 4436 4936
rect 4684 4976 4724 6112
rect 4875 6068 4917 6077
rect 4875 6028 4876 6068
rect 4916 6028 4917 6068
rect 4875 6019 4917 6028
rect 4876 5900 4916 6019
rect 4876 5851 4916 5860
rect 4876 5648 4916 5659
rect 4972 5657 5012 6448
rect 5067 6488 5109 6497
rect 5067 6448 5068 6488
rect 5108 6448 5109 6488
rect 5067 6439 5109 6448
rect 5164 6320 5204 6616
rect 5068 6280 5204 6320
rect 5260 6488 5300 6497
rect 4876 5573 4916 5608
rect 4971 5648 5013 5657
rect 4971 5608 4972 5648
rect 5012 5608 5013 5648
rect 4971 5599 5013 5608
rect 5068 5648 5108 6280
rect 5260 5909 5300 6448
rect 5355 6488 5397 6497
rect 5355 6448 5356 6488
rect 5396 6448 5397 6488
rect 5355 6439 5397 6448
rect 5356 6354 5396 6439
rect 5355 6236 5397 6245
rect 5355 6196 5356 6236
rect 5396 6196 5397 6236
rect 5355 6187 5397 6196
rect 5356 6102 5396 6187
rect 5452 5984 5492 6943
rect 5643 6824 5685 6833
rect 5643 6784 5644 6824
rect 5684 6784 5685 6824
rect 5643 6775 5685 6784
rect 5548 6488 5588 6497
rect 5548 6329 5588 6448
rect 5644 6488 5684 6775
rect 5740 6665 5780 7120
rect 5836 7160 5876 7288
rect 5836 7111 5876 7120
rect 5932 7160 5972 7169
rect 5932 7001 5972 7120
rect 6028 7160 6068 7447
rect 6123 7328 6165 7337
rect 6123 7288 6124 7328
rect 6164 7288 6165 7328
rect 6123 7279 6165 7288
rect 6028 7111 6068 7120
rect 5931 6992 5973 7001
rect 5931 6952 5932 6992
rect 5972 6952 5973 6992
rect 5931 6943 5973 6952
rect 6124 6824 6164 7279
rect 6220 7169 6260 8464
rect 6316 7505 6356 8800
rect 6411 8672 6453 8681
rect 6411 8632 6412 8672
rect 6452 8632 6453 8672
rect 6411 8623 6453 8632
rect 7179 8672 7221 8681
rect 7179 8632 7180 8672
rect 7220 8632 7221 8672
rect 7179 8623 7221 8632
rect 6412 8538 6452 8623
rect 7180 8261 7220 8623
rect 7179 8252 7221 8261
rect 7179 8212 7180 8252
rect 7220 8212 7221 8252
rect 7179 8203 7221 8212
rect 7180 8000 7220 8203
rect 7372 8084 7412 8095
rect 7372 8009 7412 8044
rect 7371 8000 7413 8009
rect 7180 7951 7220 7960
rect 7276 7960 7372 8000
rect 7412 7960 7413 8000
rect 6603 7580 6645 7589
rect 6603 7540 6604 7580
rect 6644 7540 6645 7580
rect 6603 7531 6645 7540
rect 6315 7496 6357 7505
rect 6315 7456 6316 7496
rect 6356 7456 6357 7496
rect 6315 7447 6357 7456
rect 6219 7160 6261 7169
rect 6219 7120 6220 7160
rect 6260 7120 6261 7160
rect 6219 7111 6261 7120
rect 6316 7160 6356 7169
rect 6356 7120 6452 7160
rect 6316 7111 6356 7120
rect 6220 7026 6260 7111
rect 6124 6784 6356 6824
rect 5739 6656 5781 6665
rect 5739 6616 5740 6656
rect 5780 6616 5781 6656
rect 5739 6607 5781 6616
rect 5836 6656 5876 6665
rect 6316 6656 6356 6784
rect 5876 6616 6164 6656
rect 5836 6607 5876 6616
rect 5547 6320 5589 6329
rect 5547 6280 5548 6320
rect 5588 6280 5589 6320
rect 5547 6271 5589 6280
rect 5644 6161 5684 6448
rect 5740 6488 5780 6497
rect 6028 6488 6068 6497
rect 5780 6448 5876 6488
rect 5740 6439 5780 6448
rect 5643 6152 5685 6161
rect 5643 6112 5644 6152
rect 5684 6112 5685 6152
rect 5643 6103 5685 6112
rect 5356 5944 5492 5984
rect 5259 5900 5301 5909
rect 5259 5860 5260 5900
rect 5300 5860 5301 5900
rect 5259 5851 5301 5860
rect 5356 5816 5396 5944
rect 5643 5900 5685 5909
rect 5643 5860 5644 5900
rect 5684 5860 5685 5900
rect 5643 5851 5685 5860
rect 5356 5767 5396 5776
rect 5068 5599 5108 5608
rect 5164 5648 5204 5657
rect 5164 5573 5204 5608
rect 5355 5648 5397 5657
rect 5644 5648 5684 5851
rect 5739 5732 5781 5741
rect 5739 5692 5740 5732
rect 5780 5692 5781 5732
rect 5739 5683 5781 5692
rect 5355 5608 5356 5648
rect 5396 5608 5397 5648
rect 5355 5599 5397 5608
rect 5548 5608 5644 5648
rect 4875 5564 4917 5573
rect 4875 5524 4876 5564
rect 4916 5524 4917 5564
rect 4875 5515 4917 5524
rect 5164 5564 5206 5573
rect 5164 5524 5165 5564
rect 5205 5524 5206 5564
rect 5164 5515 5206 5524
rect 5356 5514 5396 5599
rect 4928 5312 5296 5321
rect 4968 5272 5010 5312
rect 5050 5272 5092 5312
rect 5132 5272 5174 5312
rect 5214 5272 5256 5312
rect 4928 5263 5296 5272
rect 5355 5312 5397 5321
rect 5355 5272 5356 5312
rect 5396 5272 5397 5312
rect 5355 5263 5397 5272
rect 5259 5144 5301 5153
rect 5259 5104 5260 5144
rect 5300 5104 5301 5144
rect 5259 5095 5301 5104
rect 5068 4985 5108 5070
rect 4684 4927 4724 4936
rect 5067 4976 5109 4985
rect 5067 4936 5068 4976
rect 5108 4936 5109 4976
rect 5067 4927 5109 4936
rect 5260 4976 5300 5095
rect 5260 4927 5300 4936
rect 4491 4892 4533 4901
rect 4491 4852 4492 4892
rect 4532 4852 4533 4892
rect 4491 4843 4533 4852
rect 3531 4052 3573 4061
rect 3531 4012 3532 4052
rect 3572 4012 3573 4052
rect 3531 4003 3573 4012
rect 3820 4002 3860 4087
rect 3723 3968 3765 3977
rect 3723 3928 3724 3968
rect 3764 3928 3765 3968
rect 3723 3919 3765 3928
rect 3627 3716 3669 3725
rect 3436 3676 3572 3716
rect 3244 3592 3380 3632
rect 3340 3548 3380 3592
rect 3340 3499 3380 3508
rect 3436 3473 3476 3558
rect 3435 3464 3477 3473
rect 3148 3449 3284 3464
rect 3148 3424 3244 3449
rect 2764 2645 2804 2654
rect 2860 2624 2900 3424
rect 3435 3424 3436 3464
rect 3476 3424 3477 3464
rect 3435 3415 3477 3424
rect 3244 3400 3284 3409
rect 2955 3380 2997 3389
rect 2955 3340 2956 3380
rect 2996 3340 2997 3380
rect 2955 3331 2997 3340
rect 2956 2876 2996 3331
rect 3052 3296 3092 3305
rect 3092 3256 3380 3296
rect 3052 3247 3092 3256
rect 3243 3044 3285 3053
rect 3243 3004 3244 3044
rect 3284 3004 3285 3044
rect 3243 2995 3285 3004
rect 2956 2827 2996 2836
rect 2804 2605 2900 2624
rect 2764 2584 2900 2605
rect 2668 2500 2804 2540
rect 2188 1903 2228 1912
rect 2667 1952 2709 1961
rect 2667 1912 2668 1952
rect 2708 1912 2709 1952
rect 2667 1903 2709 1912
rect 1324 1112 1364 1121
rect 1324 953 1364 1072
rect 2571 1112 2613 1121
rect 2571 1072 2572 1112
rect 2612 1072 2613 1112
rect 2571 1063 2613 1072
rect 2572 978 2612 1063
rect 1323 944 1365 953
rect 1323 904 1324 944
rect 1364 904 1365 944
rect 2668 944 2708 1903
rect 2764 1112 2804 2500
rect 2860 1952 2900 2584
rect 3244 2624 3284 2995
rect 3340 2801 3380 3256
rect 3532 3053 3572 3676
rect 3627 3676 3628 3716
rect 3668 3676 3669 3716
rect 3627 3667 3669 3676
rect 3628 3464 3668 3667
rect 3628 3389 3668 3424
rect 3724 3464 3764 3919
rect 4011 3884 4053 3893
rect 4011 3844 4012 3884
rect 4052 3844 4053 3884
rect 4011 3835 4053 3844
rect 3915 3632 3957 3641
rect 3915 3592 3916 3632
rect 3956 3592 3957 3632
rect 3915 3583 3957 3592
rect 4012 3632 4052 3835
rect 4204 3800 4244 4264
rect 4012 3583 4052 3592
rect 4164 3760 4244 3800
rect 4300 4264 4436 4304
rect 3724 3415 3764 3424
rect 3916 3464 3956 3583
rect 4164 3473 4204 3760
rect 3916 3415 3956 3424
rect 4011 3464 4053 3473
rect 4011 3424 4012 3464
rect 4052 3424 4053 3464
rect 4011 3415 4053 3424
rect 4156 3464 4204 3473
rect 4196 3424 4204 3464
rect 4156 3415 4196 3424
rect 3627 3380 3669 3389
rect 3627 3340 3628 3380
rect 3668 3340 3669 3380
rect 3627 3331 3669 3340
rect 3628 3300 3668 3331
rect 4012 3330 4052 3415
rect 4107 3296 4149 3305
rect 4107 3256 4108 3296
rect 4148 3256 4149 3296
rect 4300 3296 4340 4264
rect 4396 4136 4436 4145
rect 4492 4136 4532 4843
rect 5164 4733 5204 4818
rect 5259 4808 5301 4817
rect 5259 4768 5260 4808
rect 5300 4768 5301 4808
rect 5259 4759 5301 4768
rect 4436 4096 4532 4136
rect 4588 4724 4628 4733
rect 4588 4136 4628 4684
rect 5163 4724 5205 4733
rect 5163 4684 5164 4724
rect 5204 4684 5205 4724
rect 5163 4675 5205 4684
rect 5163 4472 5205 4481
rect 5163 4432 5164 4472
rect 5204 4432 5205 4472
rect 5163 4423 5205 4432
rect 5068 4304 5108 4313
rect 4972 4264 5068 4304
rect 4396 3557 4436 4096
rect 4588 4087 4628 4096
rect 4684 4136 4724 4147
rect 4684 4061 4724 4096
rect 4972 4061 5012 4264
rect 5068 4255 5108 4264
rect 5068 4136 5108 4145
rect 5164 4136 5204 4423
rect 5108 4096 5204 4136
rect 5068 4087 5108 4096
rect 4683 4052 4725 4061
rect 4683 4012 4684 4052
rect 4724 4012 4725 4052
rect 4683 4003 4725 4012
rect 4971 4052 5013 4061
rect 4971 4012 4972 4052
rect 5012 4012 5013 4052
rect 4971 4003 5013 4012
rect 5260 3977 5300 4759
rect 4491 3968 4533 3977
rect 4876 3968 4916 3977
rect 4491 3928 4492 3968
rect 4532 3928 4533 3968
rect 4491 3919 4533 3928
rect 4780 3928 4876 3968
rect 4492 3834 4532 3919
rect 4587 3716 4629 3725
rect 4587 3676 4588 3716
rect 4628 3676 4629 3716
rect 4587 3667 4629 3676
rect 4395 3548 4437 3557
rect 4395 3508 4396 3548
rect 4436 3508 4437 3548
rect 4395 3499 4437 3508
rect 4492 3473 4532 3558
rect 4491 3464 4533 3473
rect 4491 3424 4492 3464
rect 4532 3424 4533 3464
rect 4491 3415 4533 3424
rect 4588 3464 4628 3667
rect 4780 3641 4820 3928
rect 4876 3919 4916 3928
rect 5259 3968 5301 3977
rect 5259 3928 5260 3968
rect 5300 3928 5301 3968
rect 5259 3919 5301 3928
rect 4928 3800 5296 3809
rect 4968 3760 5010 3800
rect 5050 3760 5092 3800
rect 5132 3760 5174 3800
rect 5214 3760 5256 3800
rect 4928 3751 5296 3760
rect 4779 3632 4821 3641
rect 4779 3592 4780 3632
rect 4820 3592 4821 3632
rect 4779 3583 4821 3592
rect 5163 3632 5205 3641
rect 5163 3592 5164 3632
rect 5204 3592 5205 3632
rect 5163 3583 5205 3592
rect 5067 3548 5109 3557
rect 5067 3508 5068 3548
rect 5108 3508 5109 3548
rect 5067 3499 5109 3508
rect 4588 3389 4628 3424
rect 4683 3464 4725 3473
rect 4683 3424 4684 3464
rect 4724 3424 4725 3464
rect 4683 3415 4725 3424
rect 4780 3464 4820 3473
rect 4587 3380 4629 3389
rect 4587 3340 4588 3380
rect 4628 3340 4629 3380
rect 4587 3331 4629 3340
rect 4684 3330 4724 3415
rect 4300 3256 4532 3296
rect 4107 3247 4149 3256
rect 3531 3044 3573 3053
rect 3531 3004 3532 3044
rect 3572 3004 3573 3044
rect 3531 2995 3573 3004
rect 3688 3044 4056 3053
rect 3728 3004 3770 3044
rect 3810 3004 3852 3044
rect 3892 3004 3934 3044
rect 3974 3004 4016 3044
rect 3688 2995 4056 3004
rect 4011 2876 4053 2885
rect 4011 2836 4012 2876
rect 4052 2836 4053 2876
rect 4011 2827 4053 2836
rect 3339 2792 3381 2801
rect 3339 2752 3340 2792
rect 3380 2752 3381 2792
rect 3339 2743 3381 2752
rect 3723 2792 3765 2801
rect 3723 2752 3724 2792
rect 3764 2752 3765 2792
rect 3723 2743 3765 2752
rect 3244 2575 3284 2584
rect 3340 2624 3380 2743
rect 3436 2633 3476 2718
rect 3531 2708 3573 2717
rect 3531 2668 3532 2708
rect 3572 2668 3573 2708
rect 3531 2659 3573 2668
rect 3340 2575 3380 2584
rect 3435 2624 3477 2633
rect 3435 2584 3436 2624
rect 3476 2584 3477 2624
rect 3435 2575 3477 2584
rect 3532 2624 3572 2659
rect 3532 2573 3572 2584
rect 3724 2624 3764 2743
rect 3819 2708 3861 2717
rect 3819 2668 3820 2708
rect 3860 2668 3861 2708
rect 3819 2659 3861 2668
rect 3724 2575 3764 2584
rect 3820 2624 3860 2659
rect 3820 2573 3860 2584
rect 4012 2456 4052 2827
rect 4108 2549 4148 3247
rect 4299 2792 4341 2801
rect 4299 2752 4300 2792
rect 4340 2752 4341 2792
rect 4299 2743 4341 2752
rect 4204 2633 4244 2718
rect 4203 2624 4245 2633
rect 4203 2584 4204 2624
rect 4244 2584 4245 2624
rect 4203 2575 4245 2584
rect 4300 2624 4340 2743
rect 4300 2575 4340 2584
rect 4107 2540 4149 2549
rect 4107 2500 4108 2540
rect 4148 2500 4149 2540
rect 4107 2491 4149 2500
rect 4012 2407 4052 2416
rect 4492 2456 4532 3256
rect 4780 2876 4820 3424
rect 4971 3464 5013 3473
rect 4971 3424 4972 3464
rect 5012 3424 5013 3464
rect 4971 3415 5013 3424
rect 5068 3464 5108 3499
rect 5164 3473 5204 3583
rect 4972 3330 5012 3415
rect 5068 3413 5108 3424
rect 5163 3464 5205 3473
rect 5163 3424 5164 3464
rect 5204 3424 5205 3464
rect 5163 3415 5205 3424
rect 5260 3464 5300 3473
rect 5356 3464 5396 5263
rect 5548 5153 5588 5608
rect 5644 5599 5684 5608
rect 5740 5648 5780 5683
rect 5836 5657 5876 6448
rect 6028 6077 6068 6448
rect 6124 6488 6164 6616
rect 6316 6607 6356 6616
rect 6124 6439 6164 6448
rect 6219 6488 6261 6497
rect 6219 6448 6220 6488
rect 6260 6448 6261 6488
rect 6219 6439 6261 6448
rect 6220 6354 6260 6439
rect 6412 6320 6452 7120
rect 6507 6992 6549 7001
rect 6507 6952 6508 6992
rect 6548 6952 6549 6992
rect 6507 6943 6549 6952
rect 6508 6858 6548 6943
rect 6508 6320 6548 6329
rect 6412 6280 6508 6320
rect 6508 6271 6548 6280
rect 6027 6068 6069 6077
rect 6027 6028 6028 6068
rect 6068 6028 6069 6068
rect 6027 6019 6069 6028
rect 5547 5144 5589 5153
rect 5547 5104 5548 5144
rect 5588 5104 5589 5144
rect 5547 5095 5589 5104
rect 5548 4976 5588 5095
rect 5548 4927 5588 4936
rect 5644 4976 5684 4985
rect 5644 4304 5684 4936
rect 5548 4264 5684 4304
rect 5548 3632 5588 4264
rect 5644 4136 5684 4147
rect 5644 4061 5684 4096
rect 5740 4136 5780 5608
rect 5835 5648 5877 5657
rect 5835 5608 5836 5648
rect 5876 5608 5877 5648
rect 5835 5599 5877 5608
rect 6124 5648 6164 5657
rect 6124 5144 6164 5608
rect 6220 5648 6260 5659
rect 6604 5648 6644 7531
rect 6891 7328 6933 7337
rect 6891 7288 6892 7328
rect 6932 7288 6933 7328
rect 6891 7279 6933 7288
rect 6795 7244 6837 7253
rect 6795 7204 6796 7244
rect 6836 7204 6837 7244
rect 6795 7195 6837 7204
rect 6796 7160 6836 7195
rect 6796 7109 6836 7120
rect 6892 7160 6932 7279
rect 6892 7111 6932 7120
rect 6988 7160 7028 7169
rect 7276 7160 7316 7960
rect 7371 7951 7413 7960
rect 7564 7757 7604 10672
rect 8716 10604 8756 10672
rect 8908 10604 8948 10692
rect 8716 10564 8948 10604
rect 9196 9680 9236 10692
rect 9196 9631 9236 9640
rect 9484 10692 9716 10732
rect 7756 9512 7796 9521
rect 7756 8840 7796 9472
rect 9004 9512 9044 9521
rect 9044 9472 9332 9512
rect 9004 9463 9044 9472
rect 7756 8800 8276 8840
rect 7660 8681 7700 8766
rect 7659 8672 7701 8681
rect 7659 8632 7660 8672
rect 7700 8632 7701 8672
rect 7659 8623 7701 8632
rect 8043 8672 8085 8681
rect 8043 8632 8044 8672
rect 8084 8632 8085 8672
rect 8043 8623 8085 8632
rect 8044 8538 8084 8623
rect 7852 8504 7892 8513
rect 7660 8464 7852 8504
rect 7563 7748 7605 7757
rect 7563 7708 7564 7748
rect 7604 7708 7605 7748
rect 7563 7699 7605 7708
rect 7563 7580 7605 7589
rect 7563 7540 7564 7580
rect 7604 7540 7605 7580
rect 7563 7531 7605 7540
rect 7028 7120 7276 7160
rect 6988 7111 7028 7120
rect 7276 7111 7316 7120
rect 7372 7160 7412 7169
rect 7412 7120 7508 7160
rect 7372 7111 7412 7120
rect 6699 6992 6741 7001
rect 6699 6952 6700 6992
rect 6740 6952 6741 6992
rect 6699 6943 6741 6952
rect 6700 6858 6740 6943
rect 6796 6616 7412 6656
rect 6796 6572 6836 6616
rect 6796 6523 6836 6532
rect 6892 6488 6932 6497
rect 7179 6488 7221 6497
rect 6932 6448 7124 6488
rect 6892 6439 6932 6448
rect 6700 5648 6740 5657
rect 6604 5608 6700 5648
rect 6220 5573 6260 5608
rect 6219 5564 6261 5573
rect 6219 5524 6220 5564
rect 6260 5524 6356 5564
rect 6219 5515 6261 5524
rect 6124 5104 6260 5144
rect 5932 5020 6164 5060
rect 5643 4052 5685 4061
rect 5643 4012 5644 4052
rect 5684 4012 5685 4052
rect 5643 4003 5685 4012
rect 5300 3424 5396 3464
rect 5452 3592 5684 3632
rect 5260 3415 5300 3424
rect 4876 2876 4916 2885
rect 4780 2836 4876 2876
rect 4876 2827 4916 2836
rect 4971 2876 5013 2885
rect 4971 2836 4972 2876
rect 5012 2836 5013 2876
rect 4971 2827 5013 2836
rect 4876 2624 4916 2633
rect 4972 2624 5012 2827
rect 4916 2584 5012 2624
rect 5164 2624 5204 3415
rect 4876 2575 4916 2584
rect 5164 2549 5204 2584
rect 5163 2540 5205 2549
rect 5163 2500 5164 2540
rect 5204 2500 5205 2540
rect 5163 2491 5205 2500
rect 4492 2407 4532 2416
rect 5355 2456 5397 2465
rect 5355 2416 5356 2456
rect 5396 2416 5397 2456
rect 5355 2407 5397 2416
rect 4928 2288 5296 2297
rect 4968 2248 5010 2288
rect 5050 2248 5092 2288
rect 5132 2248 5174 2288
rect 5214 2248 5256 2288
rect 4928 2239 5296 2248
rect 5259 2036 5301 2045
rect 5259 1996 5260 2036
rect 5300 1996 5301 2036
rect 5259 1987 5301 1996
rect 3436 1952 3476 1961
rect 2860 1912 3436 1952
rect 3436 1121 3476 1912
rect 3820 1952 3860 1961
rect 5068 1952 5108 1961
rect 3860 1912 4148 1952
rect 3820 1903 3860 1912
rect 3628 1709 3668 1794
rect 3627 1700 3669 1709
rect 3627 1660 3628 1700
rect 3668 1660 3669 1700
rect 3627 1651 3669 1660
rect 3688 1532 4056 1541
rect 3728 1492 3770 1532
rect 3810 1492 3852 1532
rect 3892 1492 3934 1532
rect 3974 1492 4016 1532
rect 3688 1483 4056 1492
rect 4108 1205 4148 1912
rect 5068 1784 5108 1912
rect 5260 1902 5300 1987
rect 5356 1784 5396 2407
rect 5068 1744 5396 1784
rect 4107 1196 4149 1205
rect 4107 1156 4108 1196
rect 4148 1156 4149 1196
rect 4107 1147 4149 1156
rect 3052 1112 3092 1121
rect 2764 1072 3052 1112
rect 3052 1063 3092 1072
rect 3435 1112 3477 1121
rect 3435 1072 3436 1112
rect 3476 1072 3477 1112
rect 3435 1063 3477 1072
rect 2764 944 2804 953
rect 2668 904 2764 944
rect 1323 895 1365 904
rect 2764 895 2804 904
rect 1324 449 1364 895
rect 1323 440 1365 449
rect 1323 400 1324 440
rect 1364 400 1365 440
rect 1323 391 1365 400
rect 4108 113 4148 1147
rect 5068 1121 5108 1744
rect 5452 1541 5492 3592
rect 5547 3464 5589 3473
rect 5547 3424 5548 3464
rect 5588 3424 5589 3464
rect 5547 3415 5589 3424
rect 5644 3464 5684 3592
rect 5644 3415 5684 3424
rect 5548 3330 5588 3415
rect 5547 1952 5589 1961
rect 5547 1912 5548 1952
rect 5588 1912 5589 1952
rect 5547 1903 5589 1912
rect 5644 1952 5684 1963
rect 5548 1818 5588 1903
rect 5644 1877 5684 1912
rect 5643 1868 5685 1877
rect 5643 1828 5644 1868
rect 5684 1828 5685 1868
rect 5643 1819 5685 1828
rect 5451 1532 5493 1541
rect 5451 1492 5452 1532
rect 5492 1492 5493 1532
rect 5451 1483 5493 1492
rect 4299 1112 4341 1121
rect 4299 1072 4300 1112
rect 4340 1072 4341 1112
rect 4299 1063 4341 1072
rect 5067 1112 5109 1121
rect 5067 1072 5068 1112
rect 5108 1072 5109 1112
rect 5067 1063 5109 1072
rect 5260 1112 5300 1123
rect 4300 978 4340 1063
rect 5260 1037 5300 1072
rect 5356 1112 5396 1121
rect 5452 1112 5492 1483
rect 5740 1196 5780 4096
rect 5835 4136 5877 4145
rect 5835 4096 5836 4136
rect 5876 4096 5877 4136
rect 5835 4087 5877 4096
rect 5836 2213 5876 4087
rect 5932 3809 5972 5020
rect 6124 4976 6164 5020
rect 6124 4927 6164 4936
rect 6028 4892 6068 4901
rect 5931 3800 5973 3809
rect 5931 3760 5932 3800
rect 5972 3760 5973 3800
rect 5931 3751 5973 3760
rect 6028 3464 6068 4852
rect 6220 4724 6260 5104
rect 6124 4684 6260 4724
rect 6124 4145 6164 4684
rect 6316 4640 6356 5524
rect 6603 5144 6645 5153
rect 6603 5104 6604 5144
rect 6644 5104 6645 5144
rect 6603 5095 6645 5104
rect 6220 4600 6356 4640
rect 6604 4976 6644 5095
rect 6220 4220 6260 4600
rect 6220 4171 6260 4180
rect 6123 4136 6165 4145
rect 6123 4096 6124 4136
rect 6164 4096 6165 4136
rect 6123 4087 6165 4096
rect 6124 4002 6164 4087
rect 6219 3800 6261 3809
rect 6219 3760 6220 3800
rect 6260 3760 6261 3800
rect 6219 3751 6261 3760
rect 5931 3212 5973 3221
rect 5931 3172 5932 3212
rect 5972 3172 5973 3212
rect 5931 3163 5973 3172
rect 5932 2633 5972 3163
rect 5931 2624 5973 2633
rect 5931 2584 5932 2624
rect 5972 2584 5973 2624
rect 5931 2575 5973 2584
rect 6028 2372 6068 3424
rect 6124 3464 6164 3492
rect 6220 3464 6260 3751
rect 6604 3464 6644 4936
rect 6164 3424 6260 3464
rect 6124 3415 6164 3424
rect 5932 2332 6068 2372
rect 5835 2204 5877 2213
rect 5835 2164 5836 2204
rect 5876 2164 5877 2204
rect 5835 2155 5877 2164
rect 5932 1877 5972 2332
rect 6027 2204 6069 2213
rect 6027 2164 6028 2204
rect 6068 2164 6069 2204
rect 6027 2155 6069 2164
rect 6028 1952 6068 2155
rect 6028 1903 6068 1912
rect 6124 1877 6164 1962
rect 5931 1868 5973 1877
rect 5931 1828 5932 1868
rect 5972 1828 5973 1868
rect 5931 1819 5973 1828
rect 6123 1868 6165 1877
rect 6123 1828 6124 1868
rect 6164 1828 6165 1868
rect 6123 1819 6165 1828
rect 6220 1700 6260 3424
rect 6508 3424 6604 3464
rect 6508 1877 6548 3424
rect 6604 3415 6644 3424
rect 6700 4136 6740 5608
rect 6987 5648 7029 5657
rect 6987 5608 6988 5648
rect 7028 5608 7029 5648
rect 6987 5599 7029 5608
rect 6988 4976 7028 5599
rect 7084 5060 7124 6448
rect 7179 6448 7180 6488
rect 7220 6448 7221 6488
rect 7179 6439 7221 6448
rect 7180 6354 7220 6439
rect 7180 5657 7220 5743
rect 7179 5653 7221 5657
rect 7179 5608 7180 5653
rect 7220 5608 7221 5653
rect 7179 5599 7221 5608
rect 7372 5564 7412 6616
rect 7468 5573 7508 7120
rect 7564 6581 7604 7531
rect 7660 7253 7700 8464
rect 7852 8455 7892 8464
rect 7852 8000 7892 8009
rect 7852 7673 7892 7960
rect 7947 8000 7989 8009
rect 7947 7960 7948 8000
rect 7988 7960 7989 8000
rect 7947 7951 7989 7960
rect 8044 8000 8084 8009
rect 7948 7866 7988 7951
rect 7851 7664 7893 7673
rect 7851 7624 7852 7664
rect 7892 7624 7893 7664
rect 7851 7615 7893 7624
rect 8044 7589 8084 7960
rect 8140 8000 8180 8009
rect 8043 7580 8085 7589
rect 8043 7540 8044 7580
rect 8084 7540 8085 7580
rect 8043 7531 8085 7540
rect 7755 7496 7797 7505
rect 7755 7456 7756 7496
rect 7796 7456 7797 7496
rect 7755 7447 7797 7456
rect 7659 7244 7701 7253
rect 7659 7204 7660 7244
rect 7700 7204 7701 7244
rect 7659 7195 7701 7204
rect 7756 7244 7796 7447
rect 7756 7195 7796 7204
rect 7851 7160 7893 7169
rect 7851 7120 7852 7160
rect 7892 7120 7893 7160
rect 7851 7111 7893 7120
rect 7659 7076 7701 7085
rect 7659 7036 7660 7076
rect 7700 7036 7701 7076
rect 7659 7027 7701 7036
rect 7563 6572 7605 6581
rect 7563 6532 7564 6572
rect 7604 6532 7605 6572
rect 7563 6523 7605 6532
rect 7564 6488 7604 6523
rect 7564 6438 7604 6448
rect 7660 6413 7700 7027
rect 7852 7026 7892 7111
rect 8140 6833 8180 7960
rect 8236 7085 8276 8800
rect 9292 8672 9332 9472
rect 9484 8840 9524 10692
rect 9676 10604 9716 10692
rect 9848 10672 9928 10752
rect 10348 10692 10868 10732
rect 9868 10604 9908 10672
rect 9676 10564 9908 10604
rect 10251 9512 10293 9521
rect 10251 9472 10252 9512
rect 10292 9472 10293 9512
rect 10251 9463 10293 9472
rect 10252 9378 10292 9463
rect 9484 8791 9524 8800
rect 9675 8840 9717 8849
rect 9675 8800 9676 8840
rect 9716 8800 9717 8840
rect 9675 8791 9717 8800
rect 9676 8681 9716 8791
rect 8427 8588 8469 8597
rect 8427 8548 8428 8588
rect 8468 8548 8469 8588
rect 8427 8539 8469 8548
rect 8332 8168 8372 8177
rect 8332 7337 8372 8128
rect 8331 7328 8373 7337
rect 8331 7288 8332 7328
rect 8372 7288 8373 7328
rect 8331 7279 8373 7288
rect 8332 7160 8372 7169
rect 8235 7076 8277 7085
rect 8235 7036 8236 7076
rect 8276 7036 8277 7076
rect 8235 7027 8277 7036
rect 8332 6917 8372 7120
rect 8331 6908 8373 6917
rect 8331 6868 8332 6908
rect 8372 6868 8373 6908
rect 8331 6859 8373 6868
rect 8139 6824 8181 6833
rect 8139 6784 8140 6824
rect 8180 6784 8181 6824
rect 8139 6775 8181 6784
rect 7659 6404 7701 6413
rect 7659 6364 7660 6404
rect 7700 6364 7701 6404
rect 7659 6355 7701 6364
rect 7372 5515 7412 5524
rect 7467 5564 7509 5573
rect 7467 5524 7468 5564
rect 7508 5524 7509 5564
rect 7467 5515 7509 5524
rect 7563 5480 7605 5489
rect 7563 5440 7564 5480
rect 7604 5440 7605 5480
rect 7563 5431 7605 5440
rect 7276 5060 7316 5069
rect 7084 5020 7276 5060
rect 7276 5011 7316 5020
rect 6988 4966 7124 4976
rect 6988 4936 7084 4966
rect 7084 4917 7124 4926
rect 6603 2288 6645 2297
rect 6700 2288 6740 4096
rect 7180 4141 7220 4150
rect 7083 3548 7125 3557
rect 7180 3548 7220 4101
rect 7371 3968 7413 3977
rect 7371 3928 7372 3968
rect 7412 3928 7413 3968
rect 7371 3919 7413 3928
rect 7372 3834 7412 3919
rect 7083 3508 7084 3548
rect 7124 3508 7220 3548
rect 7275 3548 7317 3557
rect 7275 3508 7276 3548
rect 7316 3508 7317 3548
rect 7083 3499 7125 3508
rect 7275 3499 7317 3508
rect 7084 3459 7124 3499
rect 7084 3410 7124 3419
rect 7276 3414 7316 3499
rect 7468 3212 7508 3221
rect 7180 2633 7220 2718
rect 7468 2717 7508 3172
rect 7564 2801 7604 5431
rect 7563 2792 7605 2801
rect 7563 2752 7564 2792
rect 7604 2752 7605 2792
rect 7563 2743 7605 2752
rect 7467 2708 7509 2717
rect 7467 2668 7468 2708
rect 7508 2668 7509 2708
rect 7467 2659 7509 2668
rect 7179 2624 7221 2633
rect 7179 2584 7180 2624
rect 7220 2584 7221 2624
rect 7179 2575 7221 2584
rect 7564 2624 7604 2743
rect 7564 2575 7604 2584
rect 6603 2248 6604 2288
rect 6644 2248 6740 2288
rect 7372 2456 7412 2465
rect 6603 2239 6645 2248
rect 6604 1952 6644 2239
rect 7083 2036 7125 2045
rect 7083 1996 7084 2036
rect 7124 1996 7125 2036
rect 7083 1987 7125 1996
rect 7275 2036 7317 2045
rect 7275 1996 7276 2036
rect 7316 1996 7317 2036
rect 7275 1987 7317 1996
rect 6604 1903 6644 1912
rect 7084 1947 7124 1987
rect 7084 1898 7124 1907
rect 7276 1902 7316 1987
rect 7372 1961 7412 2416
rect 7660 2129 7700 6355
rect 8428 5657 8468 8539
rect 8811 8168 8853 8177
rect 8811 8128 8812 8168
rect 8852 8128 8853 8168
rect 8811 8119 8853 8128
rect 8524 8000 8564 8009
rect 8332 5648 8372 5657
rect 8427 5648 8469 5657
rect 8372 5608 8428 5648
rect 8468 5608 8469 5648
rect 8332 5599 8372 5608
rect 8427 5599 8469 5608
rect 8428 5514 8468 5599
rect 8428 4976 8468 4985
rect 8428 4397 8468 4936
rect 8524 4817 8564 7960
rect 8620 8000 8660 8009
rect 8620 7589 8660 7960
rect 8812 7589 8852 8119
rect 9292 8009 9332 8632
rect 9675 8672 9717 8681
rect 9675 8632 9676 8672
rect 9716 8632 9717 8672
rect 9675 8623 9717 8632
rect 9676 8538 9716 8623
rect 10059 8252 10101 8261
rect 10059 8212 10060 8252
rect 10100 8212 10101 8252
rect 10059 8203 10101 8212
rect 8908 8000 8948 8009
rect 9099 8000 9141 8009
rect 8948 7960 9100 8000
rect 9140 7960 9141 8000
rect 8908 7951 8948 7960
rect 9099 7951 9141 7960
rect 9291 8000 9333 8009
rect 9291 7960 9292 8000
rect 9332 7960 9428 8000
rect 9291 7951 9333 7960
rect 8619 7580 8661 7589
rect 8619 7540 8620 7580
rect 8660 7540 8661 7580
rect 8619 7531 8661 7540
rect 8811 7580 8853 7589
rect 8811 7540 8812 7580
rect 8852 7540 8853 7580
rect 8811 7531 8853 7540
rect 8620 7160 8660 7531
rect 8860 7169 8900 7178
rect 8620 7129 8860 7160
rect 9003 7160 9045 7169
rect 8900 7129 8948 7160
rect 8620 7120 8948 7129
rect 8811 6656 8853 6665
rect 8811 6616 8812 6656
rect 8852 6616 8853 6656
rect 8908 6656 8948 7120
rect 9003 7120 9004 7160
rect 9044 7120 9045 7160
rect 9003 7111 9045 7120
rect 9004 7076 9044 7111
rect 9004 7025 9044 7036
rect 9004 6656 9044 6665
rect 8908 6616 9004 6656
rect 8811 6607 8853 6616
rect 9004 6607 9044 6616
rect 8812 6488 8852 6607
rect 8812 6439 8852 6448
rect 9100 5237 9140 7951
rect 9291 7664 9333 7673
rect 9291 7624 9292 7664
rect 9332 7624 9333 7664
rect 9291 7615 9333 7624
rect 9196 7160 9236 7169
rect 9196 7001 9236 7120
rect 9292 7160 9332 7615
rect 9292 7111 9332 7120
rect 9195 6992 9237 7001
rect 9195 6952 9196 6992
rect 9236 6952 9237 6992
rect 9195 6943 9237 6952
rect 9291 6740 9333 6749
rect 9291 6700 9292 6740
rect 9332 6700 9333 6740
rect 9291 6691 9333 6700
rect 9099 5228 9141 5237
rect 9099 5188 9100 5228
rect 9140 5188 9141 5228
rect 9099 5179 9141 5188
rect 8716 4976 8756 4985
rect 8620 4936 8716 4976
rect 8523 4808 8565 4817
rect 8523 4768 8524 4808
rect 8564 4768 8565 4808
rect 8523 4759 8565 4768
rect 8235 4388 8277 4397
rect 8235 4348 8236 4388
rect 8276 4348 8277 4388
rect 8235 4339 8277 4348
rect 8427 4388 8469 4397
rect 8427 4348 8428 4388
rect 8468 4348 8469 4388
rect 8427 4339 8469 4348
rect 8236 4229 8276 4339
rect 8043 4220 8085 4229
rect 8043 4180 8044 4220
rect 8084 4180 8085 4220
rect 8043 4171 8085 4180
rect 8235 4220 8277 4229
rect 8235 4180 8236 4220
rect 8276 4180 8277 4220
rect 8235 4171 8277 4180
rect 8044 4136 8084 4171
rect 7755 3968 7797 3977
rect 7755 3928 7756 3968
rect 7796 3928 7797 3968
rect 7755 3919 7797 3928
rect 7756 3548 7796 3919
rect 8044 3893 8084 4096
rect 8043 3884 8085 3893
rect 8043 3844 8044 3884
rect 8084 3844 8085 3884
rect 8043 3835 8085 3844
rect 7756 3499 7796 3508
rect 7851 3548 7893 3557
rect 7851 3508 7852 3548
rect 7892 3508 7893 3548
rect 7851 3499 7893 3508
rect 7852 3464 7892 3499
rect 8620 3473 8660 4936
rect 8716 4927 8756 4936
rect 8812 4976 8852 4985
rect 8812 4808 8852 4936
rect 9292 4976 9332 6691
rect 9292 4927 9332 4936
rect 8716 4768 8852 4808
rect 8716 4649 8756 4768
rect 9100 4724 9140 4733
rect 8715 4640 8757 4649
rect 8715 4600 8716 4640
rect 8756 4600 8757 4640
rect 8715 4591 8757 4600
rect 7852 3413 7892 3424
rect 8139 3464 8181 3473
rect 8139 3424 8140 3464
rect 8180 3424 8181 3464
rect 8139 3415 8181 3424
rect 8619 3464 8661 3473
rect 8619 3424 8620 3464
rect 8660 3424 8661 3464
rect 8619 3415 8661 3424
rect 8716 3464 8756 3473
rect 8140 3330 8180 3415
rect 8716 3389 8756 3424
rect 8715 3380 8757 3389
rect 8715 3340 8716 3380
rect 8756 3340 8757 3380
rect 8715 3331 8757 3340
rect 8716 3137 8756 3331
rect 8715 3128 8757 3137
rect 8715 3088 8716 3128
rect 8756 3088 8757 3128
rect 8715 3079 8757 3088
rect 8812 2633 8852 2718
rect 9100 2633 9140 4684
rect 9388 4145 9428 7960
rect 9963 7748 10005 7757
rect 9963 7708 9964 7748
rect 10004 7708 10005 7748
rect 9963 7699 10005 7708
rect 9675 7328 9717 7337
rect 9675 7288 9676 7328
rect 9716 7288 9717 7328
rect 9675 7279 9717 7288
rect 9676 7160 9716 7279
rect 9772 7169 9812 7254
rect 9676 7111 9716 7120
rect 9771 7160 9813 7169
rect 9771 7120 9772 7160
rect 9812 7120 9813 7160
rect 9771 7111 9813 7120
rect 9868 7160 9908 7169
rect 9484 6992 9524 7001
rect 9868 6992 9908 7120
rect 9964 7160 10004 7699
rect 10060 7673 10100 8203
rect 10348 8168 10388 10692
rect 10828 10604 10868 10692
rect 11000 10672 11080 10752
rect 12152 10672 12232 10752
rect 13304 10672 13384 10752
rect 14456 10672 14536 10752
rect 15608 10672 15688 10752
rect 16760 10672 16840 10752
rect 17912 10688 17992 10752
rect 17912 10672 17932 10688
rect 11020 10604 11060 10672
rect 10828 10564 11060 10604
rect 11595 10604 11637 10613
rect 11595 10564 11596 10604
rect 11636 10564 11637 10604
rect 11595 10555 11637 10564
rect 11500 9512 11540 9521
rect 11500 8849 11540 9472
rect 11499 8840 11541 8849
rect 11499 8800 11500 8840
rect 11540 8800 11541 8840
rect 11499 8791 11541 8800
rect 10924 8672 10964 8681
rect 10348 8119 10388 8128
rect 10539 8168 10581 8177
rect 10539 8128 10540 8168
rect 10580 8128 10581 8168
rect 10539 8119 10581 8128
rect 10155 8000 10197 8009
rect 10155 7960 10156 8000
rect 10196 7960 10197 8000
rect 10155 7951 10197 7960
rect 10540 8000 10580 8119
rect 10924 8009 10964 8632
rect 11116 8504 11156 8513
rect 11156 8464 11348 8504
rect 11116 8455 11156 8464
rect 10156 7866 10196 7951
rect 10540 7925 10580 7960
rect 10923 8000 10965 8009
rect 10923 7960 10924 8000
rect 10964 7960 10965 8000
rect 10923 7951 10965 7960
rect 11115 8000 11157 8009
rect 11115 7960 11116 8000
rect 11156 7960 11157 8000
rect 11115 7951 11157 7960
rect 10539 7916 10581 7925
rect 10539 7876 10540 7916
rect 10580 7876 10581 7916
rect 10539 7867 10581 7876
rect 10059 7664 10101 7673
rect 10059 7624 10060 7664
rect 10100 7624 10101 7664
rect 10059 7615 10101 7624
rect 9964 7111 10004 7120
rect 9524 6952 9908 6992
rect 9484 6943 9524 6952
rect 9771 6740 9813 6749
rect 10060 6740 10100 7615
rect 9771 6700 9772 6740
rect 9812 6700 10100 6740
rect 9771 6691 9813 6700
rect 9867 6572 9909 6581
rect 9867 6532 9868 6572
rect 9908 6532 9909 6572
rect 9867 6523 9909 6532
rect 9579 6488 9621 6497
rect 9579 6448 9580 6488
rect 9620 6448 9621 6488
rect 9579 6439 9621 6448
rect 9868 6488 9908 6523
rect 11116 6497 11156 7951
rect 11308 7160 11348 8464
rect 11500 7925 11540 8791
rect 11499 7916 11541 7925
rect 11499 7876 11500 7916
rect 11540 7876 11541 7916
rect 11499 7867 11541 7876
rect 11404 7169 11444 7254
rect 11308 7111 11348 7120
rect 11403 7160 11445 7169
rect 11403 7120 11404 7160
rect 11444 7120 11445 7160
rect 11403 7111 11445 7120
rect 11596 7001 11636 10555
rect 12172 9689 12212 10672
rect 11691 9680 11733 9689
rect 11691 9640 11692 9680
rect 11732 9640 11733 9680
rect 11691 9631 11733 9640
rect 12171 9680 12213 9689
rect 12171 9640 12172 9680
rect 12212 9640 12213 9680
rect 12171 9631 12213 9640
rect 13324 9680 13364 10672
rect 14476 9680 14516 10672
rect 13324 9631 13364 9640
rect 13900 9640 14516 9680
rect 11692 9546 11732 9631
rect 11884 9512 11924 9521
rect 11884 8429 11924 9472
rect 13132 9512 13172 9521
rect 12555 9344 12597 9353
rect 12555 9304 12556 9344
rect 12596 9304 12597 9344
rect 12555 9295 12597 9304
rect 12459 8756 12501 8765
rect 12459 8716 12460 8756
rect 12500 8716 12501 8756
rect 12459 8707 12501 8716
rect 12460 8672 12500 8707
rect 12171 8504 12213 8513
rect 12171 8464 12172 8504
rect 12212 8464 12213 8504
rect 12171 8455 12213 8464
rect 11883 8420 11925 8429
rect 11883 8380 11884 8420
rect 11924 8380 11925 8420
rect 11883 8371 11925 8380
rect 11788 8000 11828 8011
rect 11788 7925 11828 7960
rect 11787 7916 11829 7925
rect 11787 7876 11788 7916
rect 11828 7876 11829 7916
rect 11787 7867 11829 7876
rect 11884 7328 11924 8371
rect 12172 8000 12212 8455
rect 11979 7748 12021 7757
rect 11979 7708 11980 7748
rect 12020 7708 12021 7748
rect 11979 7699 12021 7708
rect 11980 7614 12020 7699
rect 11884 7288 12020 7328
rect 11691 7160 11733 7169
rect 11691 7120 11692 7160
rect 11732 7120 11733 7160
rect 11691 7111 11733 7120
rect 11788 7160 11828 7169
rect 11595 6992 11637 7001
rect 11595 6952 11596 6992
rect 11636 6952 11637 6992
rect 11595 6943 11637 6952
rect 11595 6824 11637 6833
rect 11500 6784 11596 6824
rect 11636 6784 11637 6824
rect 9580 5648 9620 6439
rect 9868 6437 9908 6448
rect 11115 6488 11157 6497
rect 11115 6448 11116 6488
rect 11156 6448 11157 6488
rect 11115 6439 11157 6448
rect 11116 6354 11156 6439
rect 11307 6236 11349 6245
rect 11307 6196 11308 6236
rect 11348 6196 11349 6236
rect 11307 6187 11349 6196
rect 11211 6152 11253 6161
rect 11211 6112 11212 6152
rect 11252 6112 11253 6152
rect 11211 6103 11253 6112
rect 10251 5900 10293 5909
rect 10251 5860 10252 5900
rect 10292 5860 10293 5900
rect 10251 5851 10293 5860
rect 9580 5599 9620 5608
rect 10060 5648 10100 5657
rect 9772 5564 9812 5573
rect 10060 5564 10100 5608
rect 9812 5524 10100 5564
rect 10156 5648 10196 5657
rect 9772 5515 9812 5524
rect 10156 4892 10196 5608
rect 10252 5153 10292 5851
rect 10539 5732 10581 5741
rect 10539 5692 10540 5732
rect 10580 5692 10581 5732
rect 10539 5683 10581 5692
rect 10827 5732 10869 5741
rect 10827 5692 10828 5732
rect 10868 5692 10869 5732
rect 10827 5683 10869 5692
rect 10540 5598 10580 5683
rect 10636 5648 10676 5657
rect 10251 5144 10293 5153
rect 10251 5104 10252 5144
rect 10292 5104 10293 5144
rect 10251 5095 10293 5104
rect 10540 4976 10580 4985
rect 10156 4852 10388 4892
rect 10251 4724 10293 4733
rect 10251 4684 10252 4724
rect 10292 4684 10293 4724
rect 10251 4675 10293 4684
rect 9483 4388 9525 4397
rect 9483 4348 9484 4388
rect 9524 4348 9525 4388
rect 9483 4339 9525 4348
rect 9484 4254 9524 4339
rect 9292 4136 9332 4145
rect 9387 4136 9429 4145
rect 9332 4096 9388 4136
rect 9428 4096 9429 4136
rect 9292 4087 9332 4096
rect 9387 4087 9429 4096
rect 9963 4136 10005 4145
rect 9963 4096 9964 4136
rect 10004 4096 10005 4136
rect 9963 4087 10005 4096
rect 9388 4002 9428 4087
rect 9867 3464 9909 3473
rect 9867 3424 9868 3464
rect 9908 3424 9909 3464
rect 9867 3415 9909 3424
rect 9964 3464 10004 4087
rect 10252 3809 10292 4675
rect 10251 3800 10293 3809
rect 10251 3760 10252 3800
rect 10292 3760 10293 3800
rect 10251 3751 10293 3760
rect 10155 3632 10197 3641
rect 10155 3592 10156 3632
rect 10196 3592 10197 3632
rect 10155 3583 10197 3592
rect 10156 3498 10196 3583
rect 9964 3415 10004 3424
rect 9868 3296 9908 3415
rect 9868 3256 10004 3296
rect 9964 2960 10004 3256
rect 9964 2920 10100 2960
rect 8811 2624 8853 2633
rect 8811 2584 8812 2624
rect 8852 2584 8853 2624
rect 8811 2575 8853 2584
rect 9099 2624 9141 2633
rect 9099 2584 9100 2624
rect 9140 2584 9141 2624
rect 9099 2575 9141 2584
rect 9196 2624 9236 2633
rect 9196 2540 9236 2584
rect 9675 2624 9717 2633
rect 9675 2584 9676 2624
rect 9716 2584 9717 2624
rect 9675 2575 9717 2584
rect 9196 2500 9524 2540
rect 9004 2456 9044 2465
rect 9044 2416 9428 2456
rect 9004 2407 9044 2416
rect 8907 2288 8949 2297
rect 8907 2248 8908 2288
rect 8948 2248 8949 2288
rect 8907 2239 8949 2248
rect 8331 2204 8373 2213
rect 8331 2164 8332 2204
rect 8372 2164 8373 2204
rect 8331 2155 8373 2164
rect 7659 2120 7701 2129
rect 7659 2080 7660 2120
rect 7700 2080 7701 2120
rect 7659 2071 7701 2080
rect 8139 2120 8181 2129
rect 8139 2080 8140 2120
rect 8180 2080 8181 2120
rect 8139 2071 8181 2080
rect 7371 1952 7413 1961
rect 7371 1912 7372 1952
rect 7412 1912 7413 1952
rect 7371 1903 7413 1912
rect 7851 1952 7893 1961
rect 7851 1912 7852 1952
rect 7892 1912 7893 1952
rect 7851 1903 7893 1912
rect 7948 1952 7988 1961
rect 6507 1868 6549 1877
rect 6507 1828 6508 1868
rect 6548 1828 6549 1868
rect 6507 1819 6549 1828
rect 7852 1818 7892 1903
rect 7948 1793 7988 1912
rect 7947 1784 7989 1793
rect 7947 1744 7948 1784
rect 7988 1744 7989 1784
rect 7947 1735 7989 1744
rect 5740 1147 5780 1156
rect 5836 1660 6260 1700
rect 6795 1700 6837 1709
rect 6795 1660 6796 1700
rect 6836 1660 6837 1700
rect 5836 1196 5876 1660
rect 6795 1651 6837 1660
rect 5836 1147 5876 1156
rect 6796 1126 6836 1651
rect 8140 1625 8180 2071
rect 8332 1961 8372 2155
rect 8331 1952 8373 1961
rect 8331 1912 8332 1952
rect 8372 1912 8373 1952
rect 8331 1903 8373 1912
rect 8908 1952 8948 2239
rect 8908 1903 8948 1912
rect 9388 1947 9428 2416
rect 9484 2129 9524 2500
rect 9483 2120 9525 2129
rect 9483 2080 9484 2120
rect 9524 2080 9525 2120
rect 9483 2071 9525 2080
rect 9579 2036 9621 2045
rect 9579 1996 9580 2036
rect 9620 1996 9621 2036
rect 9579 1987 9621 1996
rect 8332 1818 8372 1903
rect 9388 1898 9428 1907
rect 9580 1902 9620 1987
rect 8427 1868 8469 1877
rect 8427 1828 8428 1868
rect 8468 1828 8469 1868
rect 8427 1819 8469 1828
rect 8139 1616 8181 1625
rect 8139 1576 8140 1616
rect 8180 1576 8181 1616
rect 8139 1567 8181 1576
rect 8428 1541 8468 1819
rect 8427 1532 8469 1541
rect 8427 1492 8428 1532
rect 8468 1492 8469 1532
rect 8427 1483 8469 1492
rect 9099 1280 9141 1289
rect 9099 1240 9100 1280
rect 9140 1240 9141 1280
rect 9099 1231 9141 1240
rect 5396 1072 5492 1112
rect 6315 1112 6357 1121
rect 6315 1072 6316 1112
rect 6356 1072 6357 1112
rect 6796 1077 6836 1086
rect 9100 1112 9140 1231
rect 5356 1063 5396 1072
rect 6315 1063 6357 1072
rect 9100 1063 9140 1072
rect 4491 1028 4533 1037
rect 4491 988 4492 1028
rect 4532 988 4533 1028
rect 4491 979 4533 988
rect 5259 1028 5301 1037
rect 5259 988 5260 1028
rect 5300 988 5301 1028
rect 5259 979 5301 988
rect 4492 894 4532 979
rect 6316 978 6356 1063
rect 6987 944 7029 953
rect 6987 904 6988 944
rect 7028 904 7029 944
rect 6987 895 7029 904
rect 6988 810 7028 895
rect 4928 776 5296 785
rect 4968 736 5010 776
rect 5050 736 5092 776
rect 5132 736 5174 776
rect 5214 736 5256 776
rect 4928 727 5296 736
rect 4107 104 4149 113
rect 4107 64 4108 104
rect 4148 64 4149 104
rect 9483 104 9525 113
rect 9483 80 9484 104
rect 4107 55 4149 64
rect 9464 64 9484 80
rect 9524 80 9525 104
rect 9676 80 9716 2575
rect 9867 2204 9909 2213
rect 9867 2164 9868 2204
rect 9908 2164 9909 2204
rect 9867 2155 9909 2164
rect 9868 80 9908 2155
rect 10060 80 10100 2920
rect 10155 1700 10197 1709
rect 10155 1660 10156 1700
rect 10196 1660 10197 1700
rect 10155 1651 10197 1660
rect 10156 1448 10196 1651
rect 10252 1625 10292 3751
rect 10348 3128 10388 4852
rect 10540 4817 10580 4936
rect 10539 4808 10581 4817
rect 10539 4768 10540 4808
rect 10580 4768 10581 4808
rect 10539 4759 10581 4768
rect 10444 4136 10484 4147
rect 10444 4061 10484 4096
rect 10443 4052 10485 4061
rect 10443 4012 10444 4052
rect 10484 4012 10485 4052
rect 10443 4003 10485 4012
rect 10348 3088 10484 3128
rect 10444 2960 10484 3088
rect 10348 2920 10484 2960
rect 10348 1877 10388 2920
rect 10444 2624 10484 2633
rect 10540 2624 10580 4759
rect 10636 4733 10676 5608
rect 10635 4724 10677 4733
rect 10635 4684 10636 4724
rect 10676 4684 10677 4724
rect 10635 4675 10677 4684
rect 10732 4724 10772 4733
rect 10732 3557 10772 4684
rect 10731 3548 10773 3557
rect 10731 3508 10732 3548
rect 10772 3508 10773 3548
rect 10731 3499 10773 3508
rect 10484 2584 10580 2624
rect 10444 2575 10484 2584
rect 10828 2540 10868 5683
rect 11116 5648 11156 5657
rect 11116 5573 11156 5608
rect 11115 5564 11157 5573
rect 11115 5524 11116 5564
rect 11156 5524 11157 5564
rect 11115 5515 11157 5524
rect 11116 5144 11156 5515
rect 11020 5104 11156 5144
rect 10923 3632 10965 3641
rect 10923 3592 10924 3632
rect 10964 3592 10965 3632
rect 10923 3583 10965 3592
rect 10924 2624 10964 3583
rect 10924 2575 10964 2584
rect 11020 2624 11060 5104
rect 11115 4976 11157 4985
rect 11115 4936 11116 4976
rect 11156 4936 11157 4976
rect 11115 4927 11157 4936
rect 11116 4842 11156 4927
rect 11212 3641 11252 6103
rect 11308 6102 11348 6187
rect 11307 3716 11349 3725
rect 11307 3676 11308 3716
rect 11348 3676 11349 3716
rect 11307 3667 11349 3676
rect 11211 3632 11253 3641
rect 11211 3592 11212 3632
rect 11252 3592 11253 3632
rect 11211 3583 11253 3592
rect 11115 3548 11157 3557
rect 11115 3508 11116 3548
rect 11156 3508 11157 3548
rect 11115 3499 11157 3508
rect 11116 3464 11156 3499
rect 11116 3413 11156 3424
rect 11211 3464 11253 3473
rect 11211 3424 11212 3464
rect 11252 3424 11253 3464
rect 11211 3415 11253 3424
rect 11212 3330 11252 3415
rect 11308 3128 11348 3667
rect 11500 3632 11540 6784
rect 11595 6775 11637 6784
rect 11595 6236 11637 6245
rect 11595 6196 11596 6236
rect 11636 6196 11637 6236
rect 11595 6187 11637 6196
rect 11596 5662 11636 6187
rect 11596 5613 11636 5622
rect 11692 5228 11732 7111
rect 11788 5648 11828 7120
rect 11883 7160 11925 7169
rect 11883 7120 11884 7160
rect 11924 7120 11925 7160
rect 11883 7111 11925 7120
rect 11884 6917 11924 7111
rect 11883 6908 11925 6917
rect 11883 6868 11884 6908
rect 11924 6868 11925 6908
rect 11883 6859 11925 6868
rect 11980 6077 12020 7288
rect 12172 6488 12212 7960
rect 12364 7160 12404 7169
rect 12364 6833 12404 7120
rect 12363 6824 12405 6833
rect 12363 6784 12364 6824
rect 12404 6784 12405 6824
rect 12363 6775 12405 6784
rect 12268 6488 12308 6497
rect 12172 6448 12268 6488
rect 12075 6404 12117 6413
rect 12075 6364 12076 6404
rect 12116 6364 12117 6404
rect 12075 6355 12117 6364
rect 11979 6068 12021 6077
rect 11979 6028 11980 6068
rect 12020 6028 12021 6068
rect 11979 6019 12021 6028
rect 11788 5608 11924 5648
rect 11787 5480 11829 5489
rect 11787 5440 11788 5480
rect 11828 5440 11829 5480
rect 11787 5431 11829 5440
rect 11788 5346 11828 5431
rect 11692 5188 11828 5228
rect 11691 4136 11733 4145
rect 11691 4096 11692 4136
rect 11732 4096 11733 4136
rect 11691 4087 11733 4096
rect 11692 4002 11732 4087
rect 10732 2500 10868 2540
rect 10539 2456 10581 2465
rect 10539 2416 10540 2456
rect 10580 2416 10581 2456
rect 10539 2407 10581 2416
rect 10636 2456 10676 2465
rect 10443 2372 10485 2381
rect 10443 2332 10444 2372
rect 10484 2332 10485 2372
rect 10443 2323 10485 2332
rect 10347 1868 10389 1877
rect 10347 1828 10348 1868
rect 10388 1828 10389 1868
rect 10347 1819 10389 1828
rect 10348 1709 10388 1819
rect 10444 1793 10484 2323
rect 10540 1868 10580 2407
rect 10636 2129 10676 2416
rect 10635 2120 10677 2129
rect 10635 2080 10636 2120
rect 10676 2080 10677 2120
rect 10635 2071 10677 2080
rect 10636 1868 10676 1877
rect 10540 1828 10636 1868
rect 10636 1819 10676 1828
rect 10443 1784 10485 1793
rect 10443 1744 10444 1784
rect 10484 1744 10485 1784
rect 10443 1735 10485 1744
rect 10347 1700 10389 1709
rect 10347 1660 10348 1700
rect 10388 1660 10389 1700
rect 10347 1651 10389 1660
rect 10251 1616 10293 1625
rect 10251 1576 10252 1616
rect 10292 1576 10293 1616
rect 10251 1567 10293 1576
rect 10156 1408 10292 1448
rect 10155 1280 10197 1289
rect 10155 1240 10156 1280
rect 10196 1240 10197 1280
rect 10155 1231 10197 1240
rect 10156 1121 10196 1231
rect 10155 1112 10197 1121
rect 10155 1072 10156 1112
rect 10196 1072 10197 1112
rect 10155 1063 10197 1072
rect 10252 80 10292 1408
rect 10348 1112 10388 1121
rect 10348 953 10388 1072
rect 10347 944 10389 953
rect 10347 904 10348 944
rect 10388 904 10389 944
rect 10347 895 10389 904
rect 10444 80 10484 1735
rect 10732 1625 10772 2500
rect 11020 1784 11060 2584
rect 11212 3088 11348 3128
rect 11404 3592 11540 3632
rect 11212 2381 11252 3088
rect 11404 2792 11444 3592
rect 11308 2752 11444 2792
rect 11596 3380 11636 3389
rect 11211 2372 11253 2381
rect 11211 2332 11212 2372
rect 11252 2332 11253 2372
rect 11211 2323 11253 2332
rect 10924 1744 11060 1784
rect 11116 1952 11156 1961
rect 10827 1700 10869 1709
rect 10827 1660 10828 1700
rect 10868 1660 10869 1700
rect 10827 1651 10869 1660
rect 10539 1616 10581 1625
rect 10731 1616 10773 1625
rect 10539 1576 10540 1616
rect 10580 1576 10676 1616
rect 10539 1567 10581 1576
rect 10539 1364 10581 1373
rect 10539 1324 10540 1364
rect 10580 1324 10581 1364
rect 10539 1315 10581 1324
rect 10540 1230 10580 1315
rect 10636 80 10676 1576
rect 10731 1576 10732 1616
rect 10772 1576 10773 1616
rect 10731 1567 10773 1576
rect 10828 1566 10868 1651
rect 10827 1448 10869 1457
rect 10827 1408 10828 1448
rect 10868 1408 10869 1448
rect 10827 1399 10869 1408
rect 10731 1196 10773 1205
rect 10731 1156 10732 1196
rect 10772 1156 10773 1196
rect 10731 1147 10773 1156
rect 10732 1112 10772 1147
rect 10732 1061 10772 1072
rect 10828 80 10868 1399
rect 10924 1289 10964 1744
rect 11019 1616 11061 1625
rect 11019 1576 11020 1616
rect 11060 1576 11061 1616
rect 11019 1567 11061 1576
rect 10923 1280 10965 1289
rect 10923 1240 10924 1280
rect 10964 1240 10965 1280
rect 10923 1231 10965 1240
rect 11020 80 11060 1567
rect 11116 1373 11156 1912
rect 11212 1952 11252 1961
rect 11308 1952 11348 2752
rect 11500 2708 11540 2717
rect 11596 2708 11636 3340
rect 11540 2668 11636 2708
rect 11500 2659 11540 2668
rect 11252 1912 11348 1952
rect 11404 2624 11444 2633
rect 11404 2540 11444 2584
rect 11499 2540 11541 2549
rect 11404 2500 11500 2540
rect 11540 2500 11541 2540
rect 11212 1625 11252 1912
rect 11404 1868 11444 2500
rect 11499 2491 11541 2500
rect 11596 2036 11636 2668
rect 11692 3380 11732 3389
rect 11692 2549 11732 3340
rect 11691 2540 11733 2549
rect 11691 2500 11692 2540
rect 11732 2500 11733 2540
rect 11691 2491 11733 2500
rect 11788 2297 11828 5188
rect 11884 4145 11924 5608
rect 11979 4472 12021 4481
rect 11979 4432 11980 4472
rect 12020 4432 12021 4472
rect 11979 4423 12021 4432
rect 11980 4229 12020 4423
rect 12076 4388 12116 6355
rect 12172 4985 12212 6448
rect 12268 6439 12308 6448
rect 12460 5993 12500 8632
rect 12556 8513 12596 9295
rect 13132 8849 13172 9472
rect 13131 8840 13173 8849
rect 13131 8800 13132 8840
rect 13172 8800 13173 8840
rect 13131 8791 13173 8800
rect 13515 8840 13557 8849
rect 13515 8800 13516 8840
rect 13556 8800 13557 8840
rect 13515 8791 13557 8800
rect 13707 8840 13749 8849
rect 13707 8800 13708 8840
rect 13748 8800 13749 8840
rect 13707 8791 13749 8800
rect 13900 8840 13940 9640
rect 14667 9512 14709 9521
rect 14667 9472 14668 9512
rect 14708 9472 14709 9512
rect 14667 9463 14709 9472
rect 15244 9512 15284 9523
rect 14283 8924 14325 8933
rect 14283 8884 14284 8924
rect 14324 8884 14325 8924
rect 14283 8875 14325 8884
rect 13900 8791 13940 8800
rect 12555 8504 12597 8513
rect 12555 8464 12556 8504
rect 12596 8464 12597 8504
rect 12555 8455 12597 8464
rect 13420 8000 13460 8011
rect 13420 7925 13460 7960
rect 13419 7916 13461 7925
rect 13419 7876 13420 7916
rect 13460 7876 13461 7916
rect 13419 7867 13461 7876
rect 12843 7748 12885 7757
rect 12843 7708 12844 7748
rect 12884 7708 12885 7748
rect 12843 7699 12885 7708
rect 12555 7328 12597 7337
rect 12555 7288 12556 7328
rect 12596 7288 12597 7328
rect 12555 7279 12597 7288
rect 12459 5984 12501 5993
rect 12459 5944 12460 5984
rect 12500 5944 12501 5984
rect 12459 5935 12501 5944
rect 12171 4976 12213 4985
rect 12171 4936 12172 4976
rect 12212 4936 12213 4976
rect 12171 4927 12213 4936
rect 12364 4976 12404 4985
rect 12364 4817 12404 4936
rect 12556 4892 12596 7279
rect 12844 7174 12884 7699
rect 13131 7580 13173 7589
rect 13131 7540 13132 7580
rect 13172 7540 13173 7580
rect 13131 7531 13173 7540
rect 12844 7125 12884 7134
rect 13035 6992 13077 7001
rect 13035 6952 13036 6992
rect 13076 6952 13077 6992
rect 13035 6943 13077 6952
rect 13036 6858 13076 6943
rect 13132 5648 13172 7531
rect 13419 7244 13461 7253
rect 13419 7204 13420 7244
rect 13460 7204 13461 7244
rect 13419 7195 13461 7204
rect 13132 5599 13172 5608
rect 12460 4852 12596 4892
rect 12363 4808 12405 4817
rect 12363 4768 12364 4808
rect 12404 4768 12405 4808
rect 12363 4759 12405 4768
rect 12267 4472 12309 4481
rect 12267 4432 12268 4472
rect 12308 4432 12309 4472
rect 12267 4423 12309 4432
rect 12076 4348 12212 4388
rect 11979 4220 12021 4229
rect 11979 4180 11980 4220
rect 12020 4180 12021 4220
rect 11979 4171 12021 4180
rect 12076 4145 12116 4230
rect 11883 4136 11925 4145
rect 11883 4096 11884 4136
rect 11924 4096 11925 4136
rect 11883 4087 11925 4096
rect 12075 4136 12117 4145
rect 12075 4096 12076 4136
rect 12116 4096 12117 4136
rect 12075 4087 12117 4096
rect 11979 4052 12021 4061
rect 11979 4012 11980 4052
rect 12020 4012 12021 4052
rect 11979 4003 12021 4012
rect 11883 3968 11925 3977
rect 11883 3928 11884 3968
rect 11924 3928 11925 3968
rect 11883 3919 11925 3928
rect 11884 3834 11924 3919
rect 11883 3632 11925 3641
rect 11883 3592 11884 3632
rect 11924 3592 11925 3632
rect 11883 3583 11925 3592
rect 11884 2960 11924 3583
rect 11980 3128 12020 4003
rect 12172 3884 12212 4348
rect 12076 3844 12212 3884
rect 12268 3884 12308 4423
rect 12364 4145 12404 4759
rect 12460 4556 12500 4852
rect 12556 4724 12596 4733
rect 12596 4684 12692 4724
rect 12556 4675 12596 4684
rect 12460 4516 12596 4556
rect 12363 4136 12405 4145
rect 12363 4096 12364 4136
rect 12404 4096 12405 4136
rect 12363 4087 12405 4096
rect 12459 3968 12501 3977
rect 12459 3928 12460 3968
rect 12500 3928 12501 3968
rect 12459 3919 12501 3928
rect 12268 3844 12404 3884
rect 12076 3641 12116 3844
rect 12075 3632 12117 3641
rect 12075 3592 12076 3632
rect 12116 3592 12117 3632
rect 12075 3583 12117 3592
rect 12171 3548 12213 3557
rect 12171 3508 12172 3548
rect 12212 3508 12213 3548
rect 12171 3499 12213 3508
rect 12172 3464 12212 3499
rect 12172 3413 12212 3424
rect 11980 3088 12308 3128
rect 11884 2920 12116 2960
rect 11980 2717 12020 2719
rect 11979 2708 12021 2717
rect 11979 2668 11980 2708
rect 12020 2668 12021 2708
rect 11979 2659 12021 2668
rect 11980 2624 12020 2659
rect 11980 2575 12020 2584
rect 11787 2288 11829 2297
rect 11787 2248 11788 2288
rect 11828 2248 11829 2288
rect 11787 2239 11829 2248
rect 11596 1996 11732 2036
rect 11596 1868 11636 1877
rect 11404 1828 11596 1868
rect 11211 1616 11253 1625
rect 11211 1576 11212 1616
rect 11252 1576 11253 1616
rect 11211 1567 11253 1576
rect 11404 1457 11444 1828
rect 11596 1819 11636 1828
rect 11692 1868 11732 1996
rect 11692 1541 11732 1828
rect 11691 1532 11733 1541
rect 11691 1492 11692 1532
rect 11732 1492 11733 1532
rect 11691 1483 11733 1492
rect 11211 1448 11253 1457
rect 11211 1408 11212 1448
rect 11252 1408 11253 1448
rect 11211 1399 11253 1408
rect 11403 1448 11445 1457
rect 11403 1408 11404 1448
rect 11444 1408 11445 1448
rect 11403 1399 11445 1408
rect 11115 1364 11157 1373
rect 11115 1324 11116 1364
rect 11156 1324 11157 1364
rect 11115 1315 11157 1324
rect 11212 80 11252 1399
rect 11595 1364 11637 1373
rect 11595 1324 11596 1364
rect 11636 1324 11637 1364
rect 11595 1315 11637 1324
rect 11403 1280 11445 1289
rect 11403 1240 11404 1280
rect 11444 1240 11445 1280
rect 11403 1231 11445 1240
rect 11404 80 11444 1231
rect 11596 80 11636 1315
rect 11788 80 11828 2239
rect 11980 1112 12020 1121
rect 11884 1072 11980 1112
rect 11884 785 11924 1072
rect 11980 1063 12020 1072
rect 12076 944 12116 2920
rect 12171 2708 12213 2717
rect 12171 2668 12172 2708
rect 12212 2668 12213 2708
rect 12171 2659 12213 2668
rect 12172 1952 12212 2659
rect 12172 1903 12212 1912
rect 12172 1280 12212 1291
rect 12172 1205 12212 1240
rect 12171 1196 12213 1205
rect 12171 1156 12172 1196
rect 12212 1156 12213 1196
rect 12171 1147 12213 1156
rect 11980 904 12116 944
rect 11883 776 11925 785
rect 11883 736 11884 776
rect 11924 736 11925 776
rect 11883 727 11925 736
rect 11980 80 12020 904
rect 12268 776 12308 3088
rect 12364 2540 12404 3844
rect 12460 2638 12500 3919
rect 12460 2589 12500 2598
rect 12364 2500 12500 2540
rect 12363 1112 12405 1121
rect 12363 1072 12364 1112
rect 12404 1072 12405 1112
rect 12363 1063 12405 1072
rect 12364 978 12404 1063
rect 12460 860 12500 2500
rect 12172 736 12308 776
rect 12364 820 12500 860
rect 12172 80 12212 736
rect 12364 80 12404 820
rect 12556 80 12596 4516
rect 12652 3459 12692 4684
rect 13420 4565 13460 7195
rect 13516 6488 13556 8791
rect 13708 8672 13748 8791
rect 13708 8623 13748 8632
rect 14092 8672 14132 8683
rect 14092 8597 14132 8632
rect 14091 8588 14133 8597
rect 14091 8548 14092 8588
rect 14132 8548 14133 8588
rect 14091 8539 14133 8548
rect 13803 8000 13845 8009
rect 13803 7960 13804 8000
rect 13844 7960 13845 8000
rect 13803 7951 13845 7960
rect 13804 7866 13844 7951
rect 13612 7748 13652 7757
rect 13652 7708 13844 7748
rect 13612 7699 13652 7708
rect 13804 7160 13844 7708
rect 14284 7244 14324 8875
rect 14475 8588 14517 8597
rect 14475 8548 14476 8588
rect 14516 8548 14517 8588
rect 14475 8539 14517 8548
rect 14092 7204 14284 7244
rect 13804 7111 13844 7120
rect 13900 7160 13940 7169
rect 13900 6917 13940 7120
rect 13899 6908 13941 6917
rect 13899 6868 13900 6908
rect 13940 6868 13941 6908
rect 13899 6859 13941 6868
rect 13516 5657 13556 6448
rect 13900 6413 13940 6859
rect 13899 6404 13941 6413
rect 13899 6364 13900 6404
rect 13940 6364 13941 6404
rect 13899 6355 13941 6364
rect 13708 6236 13748 6245
rect 13748 6196 13940 6236
rect 13708 6187 13748 6196
rect 13515 5648 13557 5657
rect 13515 5608 13516 5648
rect 13556 5608 13557 5648
rect 13515 5599 13557 5608
rect 13900 4976 13940 6196
rect 13900 4927 13940 4936
rect 13996 4976 14036 4985
rect 13611 4892 13653 4901
rect 13611 4852 13612 4892
rect 13652 4852 13653 4892
rect 13611 4843 13653 4852
rect 12747 4556 12789 4565
rect 12747 4516 12748 4556
rect 12788 4516 12789 4556
rect 12747 4507 12789 4516
rect 13419 4556 13461 4565
rect 13419 4516 13420 4556
rect 13460 4516 13461 4556
rect 13419 4507 13461 4516
rect 12652 3410 12692 3419
rect 12651 2456 12693 2465
rect 12651 2416 12652 2456
rect 12692 2416 12693 2456
rect 12651 2407 12693 2416
rect 12652 2322 12692 2407
rect 12651 2120 12693 2129
rect 12651 2080 12652 2120
rect 12692 2080 12693 2120
rect 12651 2071 12693 2080
rect 12652 1947 12692 2071
rect 12652 1898 12692 1907
rect 12748 80 12788 4507
rect 13323 4136 13365 4145
rect 13323 4096 13324 4136
rect 13364 4096 13365 4136
rect 13323 4087 13365 4096
rect 13324 4002 13364 4087
rect 13515 4052 13557 4061
rect 13515 4012 13516 4052
rect 13556 4012 13557 4052
rect 13515 4003 13557 4012
rect 13516 3918 13556 4003
rect 12843 3632 12885 3641
rect 12843 3592 12844 3632
rect 12884 3592 12885 3632
rect 12843 3583 12885 3592
rect 12844 3498 12884 3583
rect 13419 3212 13461 3221
rect 13419 3172 13420 3212
rect 13460 3172 13461 3212
rect 13419 3163 13461 3172
rect 13131 2876 13173 2885
rect 13131 2836 13132 2876
rect 13172 2836 13173 2876
rect 13131 2827 13173 2836
rect 13035 2456 13077 2465
rect 13035 2416 13036 2456
rect 13076 2416 13077 2456
rect 13035 2407 13077 2416
rect 12843 2036 12885 2045
rect 12843 1996 12844 2036
rect 12884 1996 12885 2036
rect 12843 1987 12885 1996
rect 12844 1902 12884 1987
rect 13036 1868 13076 2407
rect 13036 1819 13076 1828
rect 13035 1700 13077 1709
rect 13035 1660 13036 1700
rect 13076 1660 13077 1700
rect 13035 1651 13077 1660
rect 12939 1616 12981 1625
rect 12939 1576 12940 1616
rect 12980 1576 12981 1616
rect 12939 1567 12981 1576
rect 12940 80 12980 1567
rect 13036 869 13076 1651
rect 13035 860 13077 869
rect 13035 820 13036 860
rect 13076 820 13077 860
rect 13035 811 13077 820
rect 13132 80 13172 2827
rect 13420 2633 13460 3163
rect 13419 2624 13461 2633
rect 13419 2584 13420 2624
rect 13460 2584 13461 2624
rect 13419 2575 13461 2584
rect 13420 1952 13460 2575
rect 13612 2540 13652 4843
rect 13996 4733 14036 4936
rect 13995 4724 14037 4733
rect 13995 4684 13996 4724
rect 14036 4684 14037 4724
rect 13995 4675 14037 4684
rect 14092 4481 14132 7204
rect 14284 7195 14324 7204
rect 14379 7244 14421 7253
rect 14379 7204 14380 7244
rect 14420 7204 14421 7244
rect 14379 7195 14421 7204
rect 14380 7110 14420 7195
rect 14187 7076 14229 7085
rect 14187 7036 14188 7076
rect 14228 7036 14229 7076
rect 14187 7027 14229 7036
rect 14091 4472 14133 4481
rect 14091 4432 14092 4472
rect 14132 4432 14133 4472
rect 14091 4423 14133 4432
rect 13996 4136 14036 4147
rect 13996 4061 14036 4096
rect 14092 4136 14132 4145
rect 13995 4052 14037 4061
rect 13995 4012 13996 4052
rect 14036 4012 14037 4052
rect 13995 4003 14037 4012
rect 14092 3977 14132 4096
rect 14091 3968 14133 3977
rect 14091 3928 14092 3968
rect 14132 3928 14133 3968
rect 14091 3919 14133 3928
rect 14188 3632 14228 7027
rect 14283 6656 14325 6665
rect 14283 6616 14284 6656
rect 14324 6616 14325 6656
rect 14283 6607 14325 6616
rect 14092 3592 14228 3632
rect 14284 3632 14324 6607
rect 14379 5648 14421 5657
rect 14379 5608 14380 5648
rect 14420 5608 14421 5648
rect 14379 5599 14421 5608
rect 14380 5514 14420 5599
rect 14476 5228 14516 8539
rect 14668 6749 14708 9463
rect 15244 9437 15284 9472
rect 15243 9428 15285 9437
rect 15243 9388 15244 9428
rect 15284 9388 15285 9428
rect 15243 9379 15285 9388
rect 15339 8840 15381 8849
rect 15339 8800 15340 8840
rect 15380 8800 15381 8840
rect 15339 8791 15381 8800
rect 15532 8840 15572 8849
rect 15628 8840 15668 10672
rect 16684 9680 16724 9689
rect 16780 9680 16820 10672
rect 17931 10648 17932 10672
rect 17972 10672 17992 10688
rect 19064 10672 19144 10752
rect 19276 10692 19508 10732
rect 17972 10648 17973 10672
rect 17931 10639 17973 10648
rect 19084 10604 19124 10672
rect 19276 10604 19316 10692
rect 19084 10564 19316 10604
rect 16724 9640 16820 9680
rect 19468 9680 19508 10692
rect 20216 10672 20296 10752
rect 21368 10672 21448 10752
rect 22520 10672 22600 10752
rect 23672 10672 23752 10752
rect 24824 10672 24904 10752
rect 25976 10672 26056 10752
rect 27128 10672 27208 10752
rect 28280 10672 28360 10752
rect 29259 10688 29301 10697
rect 20236 10016 20276 10672
rect 16684 9631 16724 9640
rect 19468 9631 19508 9640
rect 19948 9976 20276 10016
rect 16492 9512 16532 9521
rect 16492 8849 16532 9472
rect 17836 9512 17876 9521
rect 15572 8800 15668 8840
rect 16491 8840 16533 8849
rect 16491 8800 16492 8840
rect 16532 8800 16533 8840
rect 15532 8791 15572 8800
rect 16491 8791 16533 8800
rect 17163 8840 17205 8849
rect 17163 8800 17164 8840
rect 17204 8800 17205 8840
rect 17163 8791 17205 8800
rect 15340 8672 15380 8791
rect 15340 8623 15380 8632
rect 15915 8672 15957 8681
rect 15915 8632 15916 8672
rect 15956 8632 15957 8672
rect 15915 8623 15957 8632
rect 16683 8672 16725 8681
rect 16683 8632 16684 8672
rect 16724 8632 16725 8672
rect 16683 8623 16725 8632
rect 17164 8672 17204 8791
rect 17644 8672 17684 8681
rect 17204 8632 17300 8672
rect 17164 8623 17204 8632
rect 15916 8538 15956 8623
rect 16107 8084 16149 8093
rect 16107 8044 16108 8084
rect 16148 8044 16149 8084
rect 16107 8035 16149 8044
rect 15051 8000 15093 8009
rect 15051 7960 15052 8000
rect 15092 7960 15093 8000
rect 15051 7951 15093 7960
rect 16108 8000 16148 8035
rect 15052 7866 15092 7951
rect 16108 7949 16148 7960
rect 16011 7916 16053 7925
rect 16011 7876 16012 7916
rect 16052 7876 16053 7916
rect 16011 7867 16053 7876
rect 15244 7748 15284 7757
rect 15284 7708 15380 7748
rect 15244 7699 15284 7708
rect 14763 7580 14805 7589
rect 14763 7540 14764 7580
rect 14804 7540 14805 7580
rect 14763 7531 14805 7540
rect 14667 6740 14709 6749
rect 14667 6700 14668 6740
rect 14708 6700 14709 6740
rect 14667 6691 14709 6700
rect 14668 5648 14708 6691
rect 14764 6497 14804 7531
rect 15340 7174 15380 7708
rect 14860 7160 14900 7169
rect 15340 7125 15380 7134
rect 14763 6488 14805 6497
rect 14763 6448 14764 6488
rect 14804 6448 14805 6488
rect 14763 6439 14805 6448
rect 14764 6354 14804 6439
rect 14764 5648 14804 5657
rect 14668 5608 14764 5648
rect 14764 5599 14804 5608
rect 14571 5480 14613 5489
rect 14860 5480 14900 7120
rect 15532 6992 15572 7001
rect 15532 5573 15572 6952
rect 16012 6488 16052 7867
rect 16299 7412 16341 7421
rect 16299 7372 16300 7412
rect 16340 7372 16341 7412
rect 16299 7363 16341 7372
rect 16300 7169 16340 7363
rect 16299 7160 16341 7169
rect 16299 7120 16300 7160
rect 16340 7120 16341 7160
rect 16299 7111 16341 7120
rect 16300 7026 16340 7111
rect 15916 6448 16012 6488
rect 15819 5816 15861 5825
rect 15819 5776 15820 5816
rect 15860 5776 15861 5816
rect 15819 5767 15861 5776
rect 15531 5564 15573 5573
rect 15531 5524 15532 5564
rect 15572 5524 15573 5564
rect 15531 5515 15573 5524
rect 14571 5440 14572 5480
rect 14612 5440 14613 5480
rect 14571 5431 14613 5440
rect 14764 5440 14900 5480
rect 15435 5480 15477 5489
rect 15435 5440 15436 5480
rect 15476 5440 15477 5480
rect 14572 5346 14612 5431
rect 14476 5188 14708 5228
rect 14380 4892 14420 4901
rect 14380 4136 14420 4852
rect 14476 4892 14516 4901
rect 14516 4852 14612 4892
rect 14476 4843 14516 4852
rect 14476 4136 14516 4145
rect 14380 4096 14476 4136
rect 14284 3592 14420 3632
rect 13995 3464 14037 3473
rect 13995 3424 13996 3464
rect 14036 3424 14037 3464
rect 13995 3415 14037 3424
rect 13707 2624 13749 2633
rect 13707 2584 13708 2624
rect 13748 2584 13749 2624
rect 13707 2575 13749 2584
rect 13900 2624 13940 2633
rect 13420 1903 13460 1912
rect 13516 2500 13652 2540
rect 13227 1700 13269 1709
rect 13227 1660 13228 1700
rect 13268 1660 13269 1700
rect 13227 1651 13269 1660
rect 13228 1566 13268 1651
rect 13323 1616 13365 1625
rect 13323 1576 13324 1616
rect 13364 1576 13365 1616
rect 13323 1567 13365 1576
rect 13324 80 13364 1567
rect 13516 80 13556 2500
rect 13612 1112 13652 1121
rect 13612 953 13652 1072
rect 13611 944 13653 953
rect 13611 904 13612 944
rect 13652 904 13653 944
rect 13611 895 13653 904
rect 13708 80 13748 2575
rect 13804 1280 13844 1289
rect 13900 1280 13940 2584
rect 13996 2624 14036 3415
rect 13996 2575 14036 2584
rect 13995 2120 14037 2129
rect 13995 2080 13996 2120
rect 14036 2080 14037 2120
rect 13995 2071 14037 2080
rect 13844 1240 13940 1280
rect 13804 1231 13844 1240
rect 13996 1196 14036 2071
rect 13900 1156 14036 1196
rect 13900 80 13940 1156
rect 14092 80 14132 3592
rect 14187 3464 14229 3473
rect 14187 3424 14188 3464
rect 14228 3424 14229 3464
rect 14187 3415 14229 3424
rect 14188 3330 14228 3415
rect 14380 3380 14420 3592
rect 14284 3340 14420 3380
rect 14284 80 14324 3340
rect 14476 3137 14516 4096
rect 14572 4136 14612 4852
rect 14475 3128 14517 3137
rect 14475 3088 14476 3128
rect 14516 3088 14517 3128
rect 14475 3079 14517 3088
rect 14475 2708 14517 2717
rect 14475 2668 14476 2708
rect 14516 2668 14517 2708
rect 14475 2659 14517 2668
rect 14380 2624 14420 2633
rect 14380 281 14420 2584
rect 14476 2574 14516 2659
rect 14572 1793 14612 4096
rect 14668 2129 14708 5188
rect 14764 2885 14804 5440
rect 15435 5431 15477 5440
rect 14859 5312 14901 5321
rect 14859 5272 14860 5312
rect 14900 5272 14901 5312
rect 14859 5263 14901 5272
rect 14860 3632 14900 5263
rect 14956 4976 14996 4985
rect 14996 4936 15092 4976
rect 14956 4927 14996 4936
rect 15052 4136 15092 4936
rect 15436 4971 15476 5431
rect 15723 5144 15765 5153
rect 15723 5104 15724 5144
rect 15764 5104 15765 5144
rect 15723 5095 15765 5104
rect 15436 4922 15476 4931
rect 15628 5060 15668 5069
rect 15628 4817 15668 5020
rect 15627 4808 15669 4817
rect 15627 4768 15628 4808
rect 15668 4768 15669 4808
rect 15627 4759 15669 4768
rect 15580 4145 15620 4154
rect 15052 3809 15092 4096
rect 15147 4136 15189 4145
rect 15147 4096 15148 4136
rect 15188 4096 15189 4136
rect 15620 4105 15668 4136
rect 15580 4096 15668 4105
rect 15147 4087 15189 4096
rect 15051 3800 15093 3809
rect 15051 3760 15052 3800
rect 15092 3760 15093 3800
rect 15051 3751 15093 3760
rect 14860 3592 15092 3632
rect 14955 3464 14997 3473
rect 14955 3424 14956 3464
rect 14996 3424 14997 3464
rect 14955 3415 14997 3424
rect 14763 2876 14805 2885
rect 14763 2836 14764 2876
rect 14804 2836 14805 2876
rect 14763 2827 14805 2836
rect 14956 2624 14996 3415
rect 14763 2456 14805 2465
rect 14763 2416 14764 2456
rect 14804 2416 14805 2456
rect 14763 2407 14805 2416
rect 14667 2120 14709 2129
rect 14667 2080 14668 2120
rect 14708 2080 14709 2120
rect 14667 2071 14709 2080
rect 14668 1952 14708 1961
rect 14764 1952 14804 2407
rect 14859 2120 14901 2129
rect 14859 2080 14860 2120
rect 14900 2080 14901 2120
rect 14859 2071 14901 2080
rect 14860 1986 14900 2071
rect 14956 1961 14996 2584
rect 14708 1912 14804 1952
rect 14955 1952 14997 1961
rect 14955 1912 14956 1952
rect 14996 1912 14997 1952
rect 14571 1784 14613 1793
rect 14571 1744 14572 1784
rect 14612 1744 14613 1784
rect 14571 1735 14613 1744
rect 14475 1448 14517 1457
rect 14475 1408 14476 1448
rect 14516 1408 14517 1448
rect 14475 1399 14517 1408
rect 14379 272 14421 281
rect 14379 232 14380 272
rect 14420 232 14421 272
rect 14379 223 14421 232
rect 14476 80 14516 1399
rect 14668 953 14708 1912
rect 14955 1903 14997 1912
rect 14859 1280 14901 1289
rect 14859 1240 14860 1280
rect 14900 1240 14901 1280
rect 14859 1231 14901 1240
rect 14667 944 14709 953
rect 14667 904 14668 944
rect 14708 904 14709 944
rect 14667 895 14709 904
rect 14667 356 14709 365
rect 14667 316 14668 356
rect 14708 316 14709 356
rect 14667 307 14709 316
rect 14668 80 14708 307
rect 14860 80 14900 1231
rect 15052 80 15092 3592
rect 15148 3305 15188 4087
rect 15628 3632 15668 4096
rect 15724 4052 15764 5095
rect 15724 4003 15764 4012
rect 15628 3583 15668 3592
rect 15820 3548 15860 5767
rect 15916 4145 15956 6448
rect 16012 6439 16052 6448
rect 16204 6236 16244 6245
rect 16244 6196 16340 6236
rect 16204 6187 16244 6196
rect 16011 5648 16053 5657
rect 16011 5608 16012 5648
rect 16052 5608 16053 5648
rect 16011 5599 16053 5608
rect 16012 5321 16052 5599
rect 16204 5480 16244 5489
rect 16011 5312 16053 5321
rect 16011 5272 16012 5312
rect 16052 5272 16053 5312
rect 16011 5263 16053 5272
rect 16204 4985 16244 5440
rect 16203 4976 16245 4985
rect 16203 4936 16204 4976
rect 16244 4936 16245 4976
rect 16203 4927 16245 4936
rect 15915 4136 15957 4145
rect 15915 4096 15916 4136
rect 15956 4096 15957 4136
rect 15915 4087 15957 4096
rect 15724 3508 15860 3548
rect 15436 3464 15476 3473
rect 15724 3464 15764 3508
rect 15436 3305 15476 3424
rect 15532 3424 15764 3464
rect 16300 3464 16340 6196
rect 16395 5648 16437 5657
rect 16395 5608 16396 5648
rect 16436 5608 16437 5648
rect 16395 5599 16437 5608
rect 16396 5514 16436 5599
rect 16587 4220 16629 4229
rect 16587 4180 16588 4220
rect 16628 4180 16629 4220
rect 16587 4171 16629 4180
rect 15147 3296 15189 3305
rect 15147 3256 15148 3296
rect 15188 3256 15189 3296
rect 15147 3247 15189 3256
rect 15435 3296 15477 3305
rect 15435 3256 15436 3296
rect 15476 3256 15477 3296
rect 15435 3247 15477 3256
rect 15148 2549 15188 3247
rect 15243 3128 15285 3137
rect 15243 3088 15244 3128
rect 15284 3088 15285 3128
rect 15243 3079 15285 3088
rect 15244 2633 15284 3079
rect 15243 2624 15285 2633
rect 15243 2584 15244 2624
rect 15284 2584 15285 2624
rect 15243 2575 15285 2584
rect 15436 2629 15476 2638
rect 15147 2540 15189 2549
rect 15147 2500 15148 2540
rect 15188 2500 15189 2540
rect 15147 2491 15189 2500
rect 15148 1952 15188 1961
rect 15148 1205 15188 1912
rect 15244 1952 15284 2575
rect 15436 2129 15476 2589
rect 15435 2120 15477 2129
rect 15435 2080 15436 2120
rect 15476 2080 15477 2120
rect 15435 2071 15477 2080
rect 15244 1903 15284 1912
rect 15339 1280 15381 1289
rect 15532 1280 15572 3424
rect 16300 3415 16340 3424
rect 16395 3464 16437 3473
rect 16395 3424 16396 3464
rect 16436 3424 16437 3464
rect 16395 3415 16437 3424
rect 15627 2876 15669 2885
rect 15627 2836 15628 2876
rect 15668 2836 15669 2876
rect 15627 2827 15669 2836
rect 15628 2540 15668 2827
rect 15723 2708 15765 2717
rect 15723 2668 15724 2708
rect 15764 2668 15765 2708
rect 15723 2659 15765 2668
rect 15628 2491 15668 2500
rect 15628 1868 15668 1879
rect 15628 1793 15668 1828
rect 15724 1868 15764 2659
rect 15916 2633 15956 2718
rect 15915 2624 15957 2633
rect 15915 2584 15916 2624
rect 15956 2584 15957 2624
rect 15915 2575 15957 2584
rect 16203 1952 16245 1961
rect 16203 1912 16204 1952
rect 16244 1912 16245 1952
rect 16203 1903 16245 1912
rect 15627 1784 15669 1793
rect 15627 1744 15628 1784
rect 15668 1744 15669 1784
rect 15627 1735 15669 1744
rect 15724 1457 15764 1828
rect 16204 1818 16244 1903
rect 15723 1448 15765 1457
rect 15723 1408 15724 1448
rect 15764 1408 15765 1448
rect 15723 1399 15765 1408
rect 16299 1364 16341 1373
rect 16299 1324 16300 1364
rect 16340 1324 16341 1364
rect 16299 1315 16341 1324
rect 15339 1240 15340 1280
rect 15380 1240 15381 1280
rect 15339 1231 15381 1240
rect 15436 1240 15572 1280
rect 15147 1196 15189 1205
rect 15147 1156 15148 1196
rect 15188 1156 15189 1196
rect 15147 1147 15189 1156
rect 15243 1112 15285 1121
rect 15243 1072 15244 1112
rect 15284 1072 15285 1112
rect 15243 1063 15285 1072
rect 15244 978 15284 1063
rect 15340 860 15380 1231
rect 15244 820 15380 860
rect 15244 80 15284 820
rect 15436 80 15476 1240
rect 16300 1112 16340 1315
rect 16396 1289 16436 3415
rect 16395 1280 16437 1289
rect 16395 1240 16396 1280
rect 16436 1240 16437 1280
rect 16395 1231 16437 1240
rect 16492 1112 16532 1121
rect 16300 1072 16436 1112
rect 15627 944 15669 953
rect 15627 904 15628 944
rect 15668 904 15669 944
rect 15627 895 15669 904
rect 15628 80 15668 895
rect 15819 692 15861 701
rect 15819 652 15820 692
rect 15860 652 15861 692
rect 15819 643 15861 652
rect 15820 80 15860 643
rect 16203 440 16245 449
rect 16203 400 16204 440
rect 16244 400 16245 440
rect 16203 391 16245 400
rect 16011 272 16053 281
rect 16011 232 16012 272
rect 16052 232 16053 272
rect 16011 223 16053 232
rect 16012 80 16052 223
rect 16204 80 16244 391
rect 16396 80 16436 1072
rect 16492 785 16532 1072
rect 16491 776 16533 785
rect 16491 736 16492 776
rect 16532 736 16533 776
rect 16491 727 16533 736
rect 16588 80 16628 4171
rect 16684 3053 16724 8623
rect 17260 8168 17300 8632
rect 17356 8588 17396 8597
rect 17644 8588 17684 8632
rect 17396 8548 17684 8588
rect 17740 8672 17780 8681
rect 17356 8539 17396 8548
rect 17260 8128 17492 8168
rect 17260 8044 17396 8084
rect 17260 7925 17300 8044
rect 17356 8000 17396 8044
rect 17356 7951 17396 7960
rect 17452 7925 17492 8128
rect 17259 7916 17301 7925
rect 17259 7876 17260 7916
rect 17300 7876 17301 7916
rect 17259 7867 17301 7876
rect 17451 7916 17493 7925
rect 17451 7876 17452 7916
rect 17492 7876 17493 7916
rect 17451 7867 17493 7876
rect 17355 7832 17397 7841
rect 17355 7792 17356 7832
rect 17396 7792 17397 7832
rect 17355 7783 17397 7792
rect 17356 6329 17396 7783
rect 17452 7160 17492 7867
rect 17548 7748 17588 7757
rect 17588 7708 17684 7748
rect 17548 7699 17588 7708
rect 17548 7160 17588 7169
rect 17452 7120 17548 7160
rect 17548 7111 17588 7120
rect 17547 6488 17589 6497
rect 17547 6448 17548 6488
rect 17588 6448 17589 6488
rect 17547 6439 17589 6448
rect 17451 6404 17493 6413
rect 17451 6364 17452 6404
rect 17492 6364 17493 6404
rect 17451 6355 17493 6364
rect 17355 6320 17397 6329
rect 17355 6280 17356 6320
rect 17396 6280 17397 6320
rect 17355 6271 17397 6280
rect 17163 5648 17205 5657
rect 17163 5608 17164 5648
rect 17204 5608 17205 5648
rect 17163 5599 17205 5608
rect 17164 5069 17204 5599
rect 17163 5060 17205 5069
rect 17163 5020 17164 5060
rect 17204 5020 17205 5060
rect 17163 5011 17205 5020
rect 16779 4976 16821 4985
rect 16779 4936 16780 4976
rect 16820 4936 16821 4976
rect 16779 4927 16821 4936
rect 16876 4976 16916 4985
rect 16780 4842 16820 4927
rect 16876 3725 16916 4936
rect 16971 4892 17013 4901
rect 16971 4852 16972 4892
rect 17012 4852 17013 4892
rect 16971 4843 17013 4852
rect 16972 4061 17012 4843
rect 17067 4640 17109 4649
rect 17067 4600 17068 4640
rect 17108 4600 17109 4640
rect 17067 4591 17109 4600
rect 16971 4052 17013 4061
rect 16971 4012 16972 4052
rect 17012 4012 17013 4052
rect 16971 4003 17013 4012
rect 16971 3800 17013 3809
rect 16971 3760 16972 3800
rect 17012 3760 17013 3800
rect 16971 3751 17013 3760
rect 16875 3716 16917 3725
rect 16875 3676 16876 3716
rect 16916 3676 16917 3716
rect 16875 3667 16917 3676
rect 16876 3464 16916 3473
rect 16972 3464 17012 3751
rect 16916 3424 17012 3464
rect 16876 3415 16916 3424
rect 16780 3380 16820 3389
rect 16683 3044 16725 3053
rect 16683 3004 16684 3044
rect 16724 3004 16725 3044
rect 16683 2995 16725 3004
rect 16780 2717 16820 3340
rect 17068 3296 17108 4591
rect 17164 4136 17204 5011
rect 17259 4892 17301 4901
rect 17259 4852 17260 4892
rect 17300 4852 17301 4892
rect 17259 4843 17301 4852
rect 17356 4892 17396 4901
rect 17260 4758 17300 4843
rect 17356 4313 17396 4852
rect 17355 4304 17397 4313
rect 17355 4264 17356 4304
rect 17396 4264 17397 4304
rect 17355 4255 17397 4264
rect 17356 4136 17396 4145
rect 17164 4096 17356 4136
rect 17356 4087 17396 4096
rect 17452 3968 17492 6355
rect 16876 3256 17108 3296
rect 17260 3928 17492 3968
rect 16779 2708 16821 2717
rect 16779 2668 16780 2708
rect 16820 2668 16821 2708
rect 16779 2659 16821 2668
rect 16876 2120 16916 3256
rect 16971 3044 17013 3053
rect 16971 3004 16972 3044
rect 17012 3004 17013 3044
rect 16971 2995 17013 3004
rect 16876 2071 16916 2080
rect 16684 1938 16724 1947
rect 16684 1364 16724 1898
rect 16779 1784 16821 1793
rect 16779 1744 16780 1784
rect 16820 1744 16821 1784
rect 16779 1735 16821 1744
rect 16684 1315 16724 1324
rect 16780 80 16820 1735
rect 16972 80 17012 2995
rect 17164 2633 17204 2718
rect 17163 2624 17205 2633
rect 17163 2584 17164 2624
rect 17204 2584 17205 2624
rect 17163 2575 17205 2584
rect 17163 2120 17205 2129
rect 17163 2080 17164 2120
rect 17204 2080 17205 2120
rect 17163 2071 17205 2080
rect 17164 80 17204 2071
rect 17260 944 17300 3928
rect 17355 3548 17397 3557
rect 17355 3508 17356 3548
rect 17396 3508 17397 3548
rect 17355 3499 17397 3508
rect 17356 3464 17396 3499
rect 17356 2969 17396 3424
rect 17355 2960 17397 2969
rect 17355 2920 17356 2960
rect 17396 2920 17397 2960
rect 17355 2911 17397 2920
rect 17548 2540 17588 6439
rect 17644 5816 17684 7708
rect 17740 7160 17780 8632
rect 17836 8261 17876 9472
rect 19084 9512 19124 9521
rect 19084 9428 19124 9472
rect 19660 9428 19700 9437
rect 19084 9388 19412 9428
rect 19276 9260 19316 9269
rect 18808 9092 19176 9101
rect 18848 9052 18890 9092
rect 18930 9052 18972 9092
rect 19012 9052 19054 9092
rect 19094 9052 19136 9092
rect 18808 9043 19176 9052
rect 19083 8840 19125 8849
rect 19083 8800 19084 8840
rect 19124 8800 19125 8840
rect 19083 8791 19125 8800
rect 18124 8672 18164 8683
rect 18124 8597 18164 8632
rect 18219 8672 18261 8681
rect 18699 8672 18741 8681
rect 18219 8632 18220 8672
rect 18260 8632 18261 8672
rect 18219 8623 18261 8632
rect 18604 8632 18700 8672
rect 18740 8632 18741 8672
rect 18123 8588 18165 8597
rect 18123 8548 18124 8588
rect 18164 8548 18165 8588
rect 18123 8539 18165 8548
rect 18220 8261 18260 8623
rect 17835 8252 17877 8261
rect 17835 8212 17836 8252
rect 17876 8212 17877 8252
rect 17835 8203 17877 8212
rect 18219 8252 18261 8261
rect 18219 8212 18220 8252
rect 18260 8212 18261 8252
rect 18219 8203 18261 8212
rect 17835 8084 17877 8093
rect 17835 8044 17836 8084
rect 17876 8044 17877 8084
rect 17835 8035 17877 8044
rect 17836 8000 17876 8035
rect 17836 7841 17876 7960
rect 17835 7832 17877 7841
rect 17835 7792 17836 7832
rect 17876 7792 17877 7832
rect 17835 7783 17877 7792
rect 17740 7120 17876 7160
rect 17740 6992 17780 7001
rect 17740 6749 17780 6952
rect 17739 6740 17781 6749
rect 17739 6700 17740 6740
rect 17780 6700 17781 6740
rect 17739 6691 17781 6700
rect 17836 5909 17876 7120
rect 17931 6740 17973 6749
rect 17931 6700 17932 6740
rect 17972 6700 17973 6740
rect 17931 6691 17973 6700
rect 17932 6488 17972 6691
rect 18411 6656 18453 6665
rect 18411 6616 18412 6656
rect 18452 6616 18453 6656
rect 18411 6607 18453 6616
rect 17932 6439 17972 6448
rect 18028 6488 18068 6497
rect 17931 6320 17973 6329
rect 17931 6280 17932 6320
rect 17972 6280 17973 6320
rect 17931 6271 17973 6280
rect 17835 5900 17877 5909
rect 17835 5860 17836 5900
rect 17876 5860 17877 5900
rect 17835 5851 17877 5860
rect 17644 5776 17780 5816
rect 17644 5648 17684 5657
rect 17644 5321 17684 5608
rect 17643 5312 17685 5321
rect 17643 5272 17644 5312
rect 17684 5272 17685 5312
rect 17643 5263 17685 5272
rect 17644 4901 17684 5263
rect 17643 4892 17685 4901
rect 17643 4852 17644 4892
rect 17684 4852 17685 4892
rect 17643 4843 17685 4852
rect 17740 4808 17780 5776
rect 17932 5648 17972 6271
rect 18028 6161 18068 6448
rect 18412 6488 18452 6607
rect 18412 6439 18452 6448
rect 18507 6404 18549 6413
rect 18507 6364 18508 6404
rect 18548 6364 18549 6404
rect 18507 6355 18549 6364
rect 18508 6270 18548 6355
rect 18027 6152 18069 6161
rect 18027 6112 18028 6152
rect 18068 6112 18069 6152
rect 18027 6103 18069 6112
rect 18028 5648 18068 5657
rect 17932 5608 18028 5648
rect 18028 5599 18068 5608
rect 17836 5480 17876 5489
rect 17876 5440 18356 5480
rect 17836 5431 17876 5440
rect 17835 5312 17877 5321
rect 17835 5272 17836 5312
rect 17876 5272 17877 5312
rect 17835 5263 17877 5272
rect 18123 5312 18165 5321
rect 18123 5272 18124 5312
rect 18164 5272 18165 5312
rect 18123 5263 18165 5272
rect 17836 4976 17876 5263
rect 17836 4927 17876 4936
rect 17740 4768 17876 4808
rect 17836 3459 17876 4768
rect 18027 3548 18069 3557
rect 18027 3508 18028 3548
rect 18068 3508 18069 3548
rect 18027 3499 18069 3508
rect 17836 3410 17876 3419
rect 18028 3414 18068 3499
rect 17643 3296 17685 3305
rect 17643 3256 17644 3296
rect 17684 3256 17685 3296
rect 17643 3247 17685 3256
rect 17644 2633 17684 3247
rect 17931 2792 17973 2801
rect 17931 2752 17932 2792
rect 17972 2752 17973 2792
rect 17931 2743 17973 2752
rect 17643 2624 17685 2633
rect 17643 2584 17644 2624
rect 17684 2584 17685 2624
rect 17643 2575 17685 2584
rect 17932 2624 17972 2743
rect 17932 2575 17972 2584
rect 17452 2500 17588 2540
rect 17356 2456 17396 2465
rect 17356 1952 17396 2416
rect 17452 2129 17492 2500
rect 17451 2120 17493 2129
rect 17451 2080 17452 2120
rect 17492 2080 17493 2120
rect 17451 2071 17493 2080
rect 17452 1952 17492 1961
rect 17356 1912 17452 1952
rect 17452 1903 17492 1912
rect 17547 1952 17589 1961
rect 17547 1912 17548 1952
rect 17588 1912 17589 1952
rect 17547 1903 17589 1912
rect 17548 1818 17588 1903
rect 17932 1877 17972 1962
rect 17739 1868 17781 1877
rect 17739 1828 17740 1868
rect 17780 1828 17781 1868
rect 17739 1819 17781 1828
rect 17931 1868 17973 1877
rect 17931 1828 17932 1868
rect 17972 1828 17973 1868
rect 17931 1819 17973 1828
rect 18028 1868 18068 1879
rect 17740 1625 17780 1819
rect 18028 1793 18068 1828
rect 18027 1784 18069 1793
rect 18027 1744 18028 1784
rect 18068 1744 18069 1784
rect 18027 1735 18069 1744
rect 17739 1616 17781 1625
rect 17739 1576 17740 1616
rect 17780 1576 17781 1616
rect 17739 1567 17781 1576
rect 17931 1616 17973 1625
rect 17931 1576 17932 1616
rect 17972 1576 17973 1616
rect 17931 1567 17973 1576
rect 17547 1532 17589 1541
rect 17547 1492 17548 1532
rect 17588 1492 17589 1532
rect 17547 1483 17589 1492
rect 17356 1121 17396 1206
rect 17355 1112 17397 1121
rect 17355 1072 17356 1112
rect 17396 1072 17397 1112
rect 17355 1063 17397 1072
rect 17260 904 17396 944
rect 17356 80 17396 904
rect 17548 80 17588 1483
rect 17739 1196 17781 1205
rect 17739 1156 17740 1196
rect 17780 1156 17781 1196
rect 17739 1147 17781 1156
rect 17740 80 17780 1147
rect 17932 80 17972 1567
rect 18124 80 18164 5263
rect 18316 4971 18356 5440
rect 18411 5228 18453 5237
rect 18411 5188 18412 5228
rect 18452 5188 18453 5228
rect 18411 5179 18453 5188
rect 18316 4922 18356 4931
rect 18219 4892 18261 4901
rect 18219 4852 18220 4892
rect 18260 4852 18261 4892
rect 18219 4843 18261 4852
rect 18220 4145 18260 4843
rect 18219 4136 18261 4145
rect 18219 4096 18220 4136
rect 18260 4096 18261 4136
rect 18219 4087 18261 4096
rect 18412 3884 18452 5179
rect 18507 5060 18549 5069
rect 18507 5020 18508 5060
rect 18548 5020 18549 5060
rect 18507 5011 18549 5020
rect 18508 4926 18548 5011
rect 18604 4808 18644 8632
rect 18699 8623 18741 8632
rect 18700 8538 18740 8623
rect 19084 8093 19124 8791
rect 19276 8756 19316 9220
rect 19372 8849 19412 9388
rect 19371 8840 19413 8849
rect 19371 8800 19372 8840
rect 19412 8800 19413 8840
rect 19371 8791 19413 8800
rect 19228 8716 19316 8756
rect 19228 8714 19268 8716
rect 19228 8665 19268 8674
rect 19372 8504 19412 8513
rect 19083 8084 19125 8093
rect 19083 8044 19084 8084
rect 19124 8044 19125 8084
rect 19083 8035 19125 8044
rect 19084 8000 19124 8035
rect 19084 7925 19124 7960
rect 19372 7925 19412 8464
rect 19083 7916 19125 7925
rect 19083 7876 19084 7916
rect 19124 7876 19125 7916
rect 19083 7867 19125 7876
rect 19371 7916 19413 7925
rect 19371 7876 19372 7916
rect 19412 7876 19413 7916
rect 19371 7867 19413 7876
rect 19276 7748 19316 7757
rect 18808 7580 19176 7589
rect 18848 7540 18890 7580
rect 18930 7540 18972 7580
rect 19012 7540 19054 7580
rect 19094 7540 19136 7580
rect 18808 7531 19176 7540
rect 19276 7160 19316 7708
rect 19563 7748 19605 7757
rect 19660 7748 19700 9388
rect 19948 8840 19988 9976
rect 20048 9848 20416 9857
rect 20088 9808 20130 9848
rect 20170 9808 20212 9848
rect 20252 9808 20294 9848
rect 20334 9808 20376 9848
rect 20048 9799 20416 9808
rect 21388 9680 21428 10672
rect 21388 9631 21428 9640
rect 22444 9512 22484 9521
rect 22348 9472 22444 9512
rect 21196 9428 21236 9437
rect 20044 8840 20084 8849
rect 19948 8800 20044 8840
rect 21196 8840 21236 9388
rect 22059 8924 22101 8933
rect 22059 8884 22060 8924
rect 22100 8884 22101 8924
rect 22059 8875 22101 8884
rect 21196 8800 21524 8840
rect 20044 8791 20084 8800
rect 19852 8756 19892 8765
rect 19852 8009 19892 8716
rect 20236 8672 20276 8681
rect 20236 8513 20276 8632
rect 21484 8672 21524 8800
rect 20235 8504 20277 8513
rect 20235 8464 20236 8504
rect 20276 8464 20277 8504
rect 20235 8455 20277 8464
rect 21484 8429 21524 8632
rect 21964 8672 22004 8681
rect 21676 8588 21716 8597
rect 21964 8588 22004 8632
rect 22060 8672 22100 8875
rect 22060 8623 22100 8632
rect 21716 8548 22004 8588
rect 21676 8539 21716 8548
rect 22348 8513 22388 9472
rect 22444 9463 22484 9472
rect 22540 8840 22580 10672
rect 23692 10529 23732 10672
rect 23691 10520 23733 10529
rect 23691 10480 23692 10520
rect 23732 10480 23733 10520
rect 23691 10471 23733 10480
rect 24844 10025 24884 10672
rect 24843 10016 24885 10025
rect 24843 9976 24844 10016
rect 24884 9976 24885 10016
rect 24843 9967 24885 9976
rect 24267 9680 24309 9689
rect 24267 9640 24268 9680
rect 24308 9640 24309 9680
rect 24267 9631 24309 9640
rect 24268 9521 24308 9631
rect 23692 9512 23732 9521
rect 23019 8840 23061 8849
rect 23692 8840 23732 9472
rect 24267 9512 24309 9521
rect 24267 9472 24268 9512
rect 24308 9472 24309 9512
rect 24267 9463 24309 9472
rect 25516 9512 25556 9521
rect 24268 9378 24308 9463
rect 25516 9344 25556 9472
rect 25324 9304 25556 9344
rect 23884 9260 23924 9269
rect 22540 8800 22676 8840
rect 22443 8756 22485 8765
rect 22443 8716 22444 8756
rect 22484 8716 22485 8756
rect 22443 8707 22485 8716
rect 22444 8622 22484 8707
rect 22539 8672 22581 8681
rect 22539 8632 22540 8672
rect 22580 8632 22581 8672
rect 22539 8623 22581 8632
rect 22347 8504 22389 8513
rect 22347 8464 22348 8504
rect 22388 8464 22389 8504
rect 22347 8455 22389 8464
rect 20715 8420 20757 8429
rect 20715 8380 20716 8420
rect 20756 8380 20757 8420
rect 20715 8371 20757 8380
rect 21483 8420 21525 8429
rect 21483 8380 21484 8420
rect 21524 8380 21525 8420
rect 21483 8371 21525 8380
rect 20048 8336 20416 8345
rect 20088 8296 20130 8336
rect 20170 8296 20212 8336
rect 20252 8296 20294 8336
rect 20334 8296 20376 8336
rect 20048 8287 20416 8296
rect 19563 7708 19564 7748
rect 19604 7708 19700 7748
rect 19756 8000 19796 8009
rect 19563 7699 19605 7708
rect 19276 7111 19316 7120
rect 19371 7160 19413 7169
rect 19371 7120 19372 7160
rect 19412 7120 19413 7160
rect 19371 7111 19413 7120
rect 19372 7026 19412 7111
rect 18988 6488 19028 6499
rect 18988 6413 19028 6448
rect 19468 6474 19508 6483
rect 18987 6404 19029 6413
rect 18987 6364 18988 6404
rect 19028 6364 19029 6404
rect 18987 6355 19029 6364
rect 18808 6068 19176 6077
rect 18848 6028 18890 6068
rect 18930 6028 18972 6068
rect 19012 6028 19054 6068
rect 19094 6028 19136 6068
rect 18808 6019 19176 6028
rect 19468 5900 19508 6434
rect 19564 5993 19604 7699
rect 19756 7673 19796 7960
rect 19851 8000 19893 8009
rect 19851 7960 19852 8000
rect 19892 7960 19893 8000
rect 19851 7951 19893 7960
rect 19755 7664 19797 7673
rect 19755 7624 19756 7664
rect 19796 7624 19797 7664
rect 19755 7615 19797 7624
rect 19851 7328 19893 7337
rect 19851 7288 19852 7328
rect 19892 7288 19893 7328
rect 19756 7253 19796 7284
rect 19851 7279 19893 7288
rect 19755 7244 19797 7253
rect 19755 7204 19756 7244
rect 19796 7204 19797 7244
rect 19755 7195 19797 7204
rect 19756 7160 19796 7195
rect 19756 7085 19796 7120
rect 19852 7160 19892 7279
rect 19755 7076 19797 7085
rect 19755 7036 19756 7076
rect 19796 7036 19797 7076
rect 19755 7027 19797 7036
rect 19852 6740 19892 7120
rect 20332 7160 20372 7169
rect 20372 7120 20564 7160
rect 20332 7111 20372 7120
rect 20048 6824 20416 6833
rect 20088 6784 20130 6824
rect 20170 6784 20212 6824
rect 20252 6784 20294 6824
rect 20334 6784 20376 6824
rect 20048 6775 20416 6784
rect 19756 6700 19892 6740
rect 19660 6572 19700 6581
rect 19563 5984 19605 5993
rect 19563 5944 19564 5984
rect 19604 5944 19605 5984
rect 19563 5935 19605 5944
rect 19468 5851 19508 5860
rect 19660 5741 19700 6532
rect 19756 6497 19796 6700
rect 20524 6581 20564 7120
rect 19851 6572 19893 6581
rect 19851 6532 19852 6572
rect 19892 6532 19893 6572
rect 19851 6523 19893 6532
rect 20523 6572 20565 6581
rect 20523 6532 20524 6572
rect 20564 6532 20660 6572
rect 20523 6523 20565 6532
rect 19755 6488 19797 6497
rect 19755 6448 19756 6488
rect 19796 6448 19797 6488
rect 19755 6439 19797 6448
rect 19852 6488 19892 6523
rect 19852 6437 19892 6448
rect 19659 5732 19701 5741
rect 19659 5692 19660 5732
rect 19700 5692 19701 5732
rect 19659 5683 19701 5692
rect 20235 5732 20277 5741
rect 20235 5692 20236 5732
rect 20276 5692 20277 5732
rect 20235 5683 20277 5692
rect 19276 5648 19316 5657
rect 19180 5608 19276 5648
rect 18699 5312 18741 5321
rect 18699 5272 18700 5312
rect 18740 5272 18741 5312
rect 18699 5263 18741 5272
rect 18700 5153 18740 5263
rect 18699 5144 18741 5153
rect 18699 5104 18700 5144
rect 18740 5104 18741 5144
rect 18699 5095 18741 5104
rect 18796 4976 18836 4985
rect 18316 3844 18452 3884
rect 18508 4768 18644 4808
rect 18700 4936 18796 4976
rect 18219 3800 18261 3809
rect 18219 3760 18220 3800
rect 18260 3760 18261 3800
rect 18219 3751 18261 3760
rect 18220 1112 18260 3751
rect 18316 1196 18356 3844
rect 18508 2540 18548 4768
rect 18700 4388 18740 4936
rect 18796 4927 18836 4936
rect 18892 4976 18932 4985
rect 18892 4733 18932 4936
rect 19083 4892 19125 4901
rect 19180 4892 19220 5608
rect 19276 5599 19316 5608
rect 20236 5598 20276 5683
rect 20428 5480 20468 5489
rect 20468 5440 20564 5480
rect 20428 5431 20468 5440
rect 20524 5321 20564 5440
rect 20048 5312 20416 5321
rect 20088 5272 20130 5312
rect 20170 5272 20212 5312
rect 20252 5272 20294 5312
rect 20334 5272 20376 5312
rect 20048 5263 20416 5272
rect 20523 5312 20565 5321
rect 20523 5272 20524 5312
rect 20564 5272 20565 5312
rect 20523 5263 20565 5272
rect 20620 5237 20660 6532
rect 20716 5405 20756 8371
rect 21003 8084 21045 8093
rect 21003 8044 21004 8084
rect 21044 8044 21045 8084
rect 21003 8035 21045 8044
rect 21004 8000 21044 8035
rect 21004 7949 21044 7960
rect 21196 7748 21236 7757
rect 20908 7708 21196 7748
rect 20908 7244 20948 7708
rect 21196 7699 21236 7708
rect 21388 7748 21428 7757
rect 21388 7412 21428 7708
rect 21484 7664 21524 8371
rect 22540 8345 22580 8623
rect 22539 8336 22581 8345
rect 22539 8296 22540 8336
rect 22580 8296 22581 8336
rect 22539 8287 22581 8296
rect 22540 8168 22580 8177
rect 22636 8168 22676 8800
rect 23019 8800 23020 8840
rect 23060 8800 23061 8840
rect 23019 8791 23061 8800
rect 23308 8800 23732 8840
rect 23788 9220 23884 9260
rect 23020 8672 23060 8791
rect 22827 8252 22869 8261
rect 22827 8212 22828 8252
rect 22868 8212 22869 8252
rect 22827 8203 22869 8212
rect 22580 8128 22676 8168
rect 22540 8119 22580 8128
rect 22347 8084 22389 8093
rect 22347 8044 22348 8084
rect 22388 8044 22389 8084
rect 22347 8035 22389 8044
rect 21579 7916 21621 7925
rect 21579 7876 21580 7916
rect 21620 7876 21621 7916
rect 21579 7867 21621 7876
rect 22348 7916 22388 8035
rect 22828 8000 22868 8203
rect 23020 8009 23060 8632
rect 23308 8429 23348 8800
rect 23548 8681 23588 8690
rect 23788 8672 23828 9220
rect 23884 9211 23924 9220
rect 23588 8641 23828 8672
rect 23548 8632 23828 8641
rect 24363 8588 24405 8597
rect 24363 8548 24364 8588
rect 24404 8548 24405 8588
rect 24363 8539 24405 8548
rect 23692 8504 23732 8513
rect 23404 8464 23692 8504
rect 23307 8420 23349 8429
rect 23307 8380 23308 8420
rect 23348 8380 23349 8420
rect 23307 8371 23349 8380
rect 22828 7951 22868 7960
rect 23019 8000 23061 8009
rect 23019 7960 23020 8000
rect 23060 7960 23061 8000
rect 23019 7951 23061 7960
rect 22348 7867 22388 7876
rect 21580 7782 21620 7867
rect 21484 7624 21620 7664
rect 21388 7372 21524 7412
rect 20860 7204 20948 7244
rect 21004 7288 21428 7328
rect 20860 7202 20900 7204
rect 20860 7153 20900 7162
rect 21004 7076 21044 7288
rect 21388 7244 21428 7288
rect 21388 7195 21428 7204
rect 21004 7027 21044 7036
rect 21099 7076 21141 7085
rect 21484 7076 21524 7372
rect 21580 7085 21620 7624
rect 23404 7244 23444 8464
rect 23692 8455 23732 8464
rect 24364 8429 24404 8539
rect 25324 8513 25364 9304
rect 25708 9260 25748 9269
rect 25420 9220 25708 9260
rect 25420 8672 25460 9220
rect 25708 9211 25748 9220
rect 25996 9101 26036 10672
rect 27148 10109 27188 10672
rect 27147 10100 27189 10109
rect 27147 10060 27148 10100
rect 27188 10060 27189 10100
rect 27147 10051 27189 10060
rect 27724 9512 27764 9521
rect 25995 9092 26037 9101
rect 25995 9052 25996 9092
rect 26036 9052 26037 9092
rect 25995 9043 26037 9052
rect 25515 8756 25557 8765
rect 25515 8716 25516 8756
rect 25556 8716 25557 8756
rect 25515 8707 25557 8716
rect 25420 8623 25460 8632
rect 25516 8672 25556 8707
rect 27004 8681 27044 8690
rect 25516 8621 25556 8632
rect 25899 8672 25941 8681
rect 25899 8632 25900 8672
rect 25940 8632 25941 8672
rect 25899 8623 25941 8632
rect 25996 8672 26036 8681
rect 26476 8672 26516 8681
rect 25900 8538 25940 8623
rect 25323 8504 25365 8513
rect 25323 8464 25324 8504
rect 25364 8464 25365 8504
rect 25323 8455 25365 8464
rect 24075 8420 24117 8429
rect 24075 8380 24076 8420
rect 24116 8380 24117 8420
rect 24075 8371 24117 8380
rect 24363 8420 24405 8429
rect 24363 8380 24364 8420
rect 24404 8380 24405 8420
rect 24363 8371 24405 8380
rect 24076 8000 24116 8371
rect 24076 7951 24116 7960
rect 23883 7748 23925 7757
rect 23883 7708 23884 7748
rect 23924 7708 23925 7748
rect 23883 7699 23925 7708
rect 24267 7748 24309 7757
rect 24267 7708 24268 7748
rect 24308 7708 24309 7748
rect 24267 7699 24309 7708
rect 23404 7195 23444 7204
rect 21675 7160 21717 7169
rect 21675 7120 21676 7160
rect 21716 7120 21717 7160
rect 21675 7111 21717 7120
rect 21099 7036 21100 7076
rect 21140 7036 21141 7076
rect 21099 7027 21141 7036
rect 21388 7036 21524 7076
rect 21579 7076 21621 7085
rect 21579 7036 21580 7076
rect 21620 7036 21621 7076
rect 21003 6908 21045 6917
rect 21003 6868 21004 6908
rect 21044 6868 21045 6908
rect 21003 6859 21045 6868
rect 20715 5396 20757 5405
rect 20715 5356 20716 5396
rect 20756 5356 20757 5396
rect 20715 5347 20757 5356
rect 20619 5228 20661 5237
rect 20619 5188 20620 5228
rect 20660 5188 20661 5228
rect 20619 5179 20661 5188
rect 20524 5144 20564 5153
rect 20524 5060 20564 5104
rect 20524 5020 20852 5060
rect 19852 4976 19892 4985
rect 19892 4936 19988 4976
rect 19852 4927 19892 4936
rect 19083 4852 19084 4892
rect 19124 4852 19220 4892
rect 19275 4892 19317 4901
rect 19275 4852 19276 4892
rect 19316 4852 19317 4892
rect 19083 4843 19125 4852
rect 19275 4843 19317 4852
rect 19372 4892 19412 4901
rect 19276 4758 19316 4843
rect 19372 4733 19412 4852
rect 18891 4724 18933 4733
rect 18891 4684 18892 4724
rect 18932 4684 18933 4724
rect 18891 4675 18933 4684
rect 19371 4724 19413 4733
rect 19371 4684 19372 4724
rect 19412 4684 19413 4724
rect 19371 4675 19413 4684
rect 18808 4556 19176 4565
rect 18848 4516 18890 4556
rect 18930 4516 18972 4556
rect 19012 4516 19054 4556
rect 19094 4516 19136 4556
rect 18808 4507 19176 4516
rect 18796 4388 18836 4397
rect 18700 4348 18796 4388
rect 18796 4339 18836 4348
rect 19948 4313 19988 4936
rect 20380 4934 20420 4943
rect 20380 4892 20420 4894
rect 20715 4892 20757 4901
rect 20380 4852 20660 4892
rect 20043 4724 20085 4733
rect 20043 4684 20044 4724
rect 20084 4684 20085 4724
rect 20043 4675 20085 4684
rect 18603 4304 18645 4313
rect 18603 4264 18604 4304
rect 18644 4264 18645 4304
rect 18603 4255 18645 4264
rect 19371 4304 19413 4313
rect 19371 4264 19372 4304
rect 19412 4264 19413 4304
rect 19371 4255 19413 4264
rect 19563 4304 19605 4313
rect 19563 4264 19564 4304
rect 19604 4264 19605 4304
rect 19563 4255 19605 4264
rect 19947 4304 19989 4313
rect 19947 4264 19948 4304
rect 19988 4264 19989 4304
rect 19947 4255 19989 4264
rect 18604 4145 18644 4255
rect 18603 4136 18645 4145
rect 18603 4096 18604 4136
rect 18644 4096 18645 4136
rect 18603 4087 18645 4096
rect 19275 4136 19317 4145
rect 19275 4096 19276 4136
rect 19316 4096 19317 4136
rect 19275 4087 19317 4096
rect 18604 4002 18644 4087
rect 19276 4002 19316 4087
rect 18808 3044 19176 3053
rect 18848 3004 18890 3044
rect 18930 3004 18972 3044
rect 19012 3004 19054 3044
rect 19094 3004 19136 3044
rect 18808 2995 19176 3004
rect 19372 2876 19412 4255
rect 19564 4145 19604 4255
rect 19563 4136 19605 4145
rect 19563 4096 19564 4136
rect 19604 4096 19605 4136
rect 19563 4087 19605 4096
rect 19659 3800 19701 3809
rect 19659 3760 19660 3800
rect 19700 3760 19701 3800
rect 19659 3751 19701 3760
rect 19660 3464 19700 3751
rect 19660 3415 19700 3424
rect 19948 3053 19988 4255
rect 20044 3977 20084 4675
rect 20620 4388 20660 4852
rect 20715 4852 20716 4892
rect 20756 4852 20757 4892
rect 20715 4843 20757 4852
rect 20716 4758 20756 4843
rect 20716 4388 20756 4397
rect 20620 4348 20716 4388
rect 20716 4339 20756 4348
rect 20524 4145 20564 4230
rect 20523 4136 20565 4145
rect 20523 4096 20524 4136
rect 20564 4096 20565 4136
rect 20523 4087 20565 4096
rect 20043 3968 20085 3977
rect 20043 3928 20044 3968
rect 20084 3928 20085 3968
rect 20043 3919 20085 3928
rect 20048 3800 20416 3809
rect 20088 3760 20130 3800
rect 20170 3760 20212 3800
rect 20252 3760 20294 3800
rect 20334 3760 20376 3800
rect 20048 3751 20416 3760
rect 19947 3044 19989 3053
rect 19947 3004 19948 3044
rect 19988 3004 19989 3044
rect 19947 2995 19989 3004
rect 20235 3044 20277 3053
rect 20235 3004 20236 3044
rect 20276 3004 20277 3044
rect 20235 2995 20277 3004
rect 20139 2960 20181 2969
rect 20139 2920 20140 2960
rect 20180 2920 20181 2960
rect 20139 2911 20181 2920
rect 19180 2836 19412 2876
rect 18603 2624 18645 2633
rect 18603 2584 18604 2624
rect 18644 2584 18645 2624
rect 18603 2575 18645 2584
rect 19180 2624 19220 2836
rect 19755 2792 19797 2801
rect 19755 2752 19756 2792
rect 19796 2752 19892 2792
rect 19755 2743 19797 2752
rect 19275 2708 19317 2717
rect 19275 2668 19276 2708
rect 19316 2668 19317 2708
rect 19275 2659 19317 2668
rect 19180 2575 19220 2584
rect 18412 2500 18548 2540
rect 18412 1280 18452 2500
rect 18508 1952 18548 1961
rect 18508 1625 18548 1912
rect 18507 1616 18549 1625
rect 18507 1576 18508 1616
rect 18548 1576 18549 1616
rect 18507 1567 18549 1576
rect 18604 1457 18644 2575
rect 18891 2288 18933 2297
rect 18891 2248 18892 2288
rect 18932 2248 18933 2288
rect 18891 2239 18933 2248
rect 18892 2129 18932 2239
rect 18891 2120 18933 2129
rect 18891 2080 18892 2120
rect 18932 2080 18933 2120
rect 18891 2071 18933 2080
rect 19180 2120 19220 2129
rect 19276 2120 19316 2659
rect 19372 2549 19412 2634
rect 19563 2624 19605 2633
rect 19660 2624 19700 2633
rect 19563 2584 19564 2624
rect 19604 2584 19660 2624
rect 19563 2575 19605 2584
rect 19660 2575 19700 2584
rect 19755 2624 19797 2633
rect 19755 2584 19756 2624
rect 19796 2584 19797 2624
rect 19755 2575 19797 2584
rect 19371 2540 19413 2549
rect 19371 2500 19372 2540
rect 19412 2500 19413 2540
rect 19371 2491 19413 2500
rect 19756 2129 19796 2575
rect 19852 2540 19892 2752
rect 19948 2624 19988 2633
rect 20140 2624 20180 2911
rect 19948 2540 19988 2584
rect 19852 2500 19988 2540
rect 19948 2381 19988 2500
rect 20044 2584 20180 2624
rect 20044 2540 20084 2584
rect 20236 2549 20276 2995
rect 20332 2792 20372 2801
rect 20044 2491 20084 2500
rect 20235 2540 20277 2549
rect 20235 2500 20236 2540
rect 20276 2500 20277 2540
rect 20235 2491 20277 2500
rect 20332 2465 20372 2752
rect 20716 2708 20756 2717
rect 20812 2708 20852 5020
rect 20908 4724 20948 4733
rect 20908 3641 20948 4684
rect 21004 4388 21044 6859
rect 21100 6488 21140 7027
rect 21100 6439 21140 6448
rect 21196 6992 21236 7001
rect 21196 5237 21236 6952
rect 21291 6656 21333 6665
rect 21291 6616 21292 6656
rect 21332 6616 21333 6656
rect 21291 6607 21333 6616
rect 21292 6522 21332 6607
rect 21195 5228 21237 5237
rect 21195 5188 21196 5228
rect 21236 5188 21237 5228
rect 21195 5179 21237 5188
rect 21099 4892 21141 4901
rect 21099 4852 21100 4892
rect 21140 4852 21141 4892
rect 21099 4843 21141 4852
rect 21100 4758 21140 4843
rect 21292 4817 21332 4902
rect 21291 4808 21333 4817
rect 21291 4768 21292 4808
rect 21332 4768 21333 4808
rect 21291 4759 21333 4768
rect 21291 4556 21333 4565
rect 21291 4516 21292 4556
rect 21332 4516 21333 4556
rect 21291 4507 21333 4516
rect 21004 4348 21236 4388
rect 21100 4136 21140 4145
rect 20907 3632 20949 3641
rect 20907 3592 20908 3632
rect 20948 3592 20949 3632
rect 20907 3583 20949 3592
rect 21100 3632 21140 4096
rect 21196 4136 21236 4348
rect 21292 4145 21332 4507
rect 21196 4087 21236 4096
rect 21291 4136 21333 4145
rect 21291 4096 21292 4136
rect 21332 4096 21333 4136
rect 21291 4087 21333 4096
rect 21195 3968 21237 3977
rect 21195 3928 21196 3968
rect 21236 3928 21237 3968
rect 21195 3919 21237 3928
rect 21100 3583 21140 3592
rect 20908 3464 20948 3475
rect 20908 3389 20948 3424
rect 21003 3464 21045 3473
rect 21003 3424 21004 3464
rect 21044 3424 21045 3464
rect 21003 3415 21045 3424
rect 20907 3380 20949 3389
rect 20907 3340 20908 3380
rect 20948 3340 20949 3380
rect 20907 3331 20949 3340
rect 20756 2668 20852 2708
rect 20907 2708 20949 2717
rect 20907 2668 20908 2708
rect 20948 2668 20949 2708
rect 20716 2659 20756 2668
rect 20907 2659 20949 2668
rect 20908 2574 20948 2659
rect 20331 2456 20373 2465
rect 20331 2416 20332 2456
rect 20372 2416 20373 2456
rect 20331 2407 20373 2416
rect 20524 2456 20564 2465
rect 19947 2372 19989 2381
rect 19947 2332 19948 2372
rect 19988 2332 19989 2372
rect 19947 2323 19989 2332
rect 19851 2288 19893 2297
rect 19851 2248 19852 2288
rect 19892 2248 19893 2288
rect 19851 2239 19893 2248
rect 20048 2288 20416 2297
rect 20088 2248 20130 2288
rect 20170 2248 20212 2288
rect 20252 2248 20294 2288
rect 20334 2248 20376 2288
rect 20048 2239 20416 2248
rect 19220 2080 19316 2120
rect 19755 2120 19797 2129
rect 19755 2080 19756 2120
rect 19796 2080 19797 2120
rect 19180 2071 19220 2080
rect 19755 2071 19797 2080
rect 19371 1952 19413 1961
rect 18988 1938 19028 1947
rect 19371 1912 19372 1952
rect 19412 1912 19413 1952
rect 19371 1903 19413 1912
rect 18988 1700 19028 1898
rect 18700 1660 19028 1700
rect 19275 1700 19317 1709
rect 19275 1660 19276 1700
rect 19316 1660 19317 1700
rect 18603 1448 18645 1457
rect 18603 1408 18604 1448
rect 18644 1408 18645 1448
rect 18603 1399 18645 1408
rect 18412 1240 18548 1280
rect 18316 1156 18452 1196
rect 18220 1072 18356 1112
rect 18316 80 18356 1072
rect 18412 953 18452 1156
rect 18411 944 18453 953
rect 18411 904 18412 944
rect 18452 904 18453 944
rect 18411 895 18453 904
rect 18508 80 18548 1240
rect 18604 1112 18644 1399
rect 18700 1280 18740 1660
rect 19275 1651 19317 1660
rect 18808 1532 19176 1541
rect 18848 1492 18890 1532
rect 18930 1492 18972 1532
rect 19012 1492 19054 1532
rect 19094 1492 19136 1532
rect 18808 1483 19176 1492
rect 18891 1364 18933 1373
rect 18891 1324 18892 1364
rect 18932 1324 18933 1364
rect 18891 1315 18933 1324
rect 18796 1280 18836 1289
rect 18700 1240 18796 1280
rect 18796 1231 18836 1240
rect 18604 1063 18644 1072
rect 18699 944 18741 953
rect 18699 904 18700 944
rect 18740 904 18741 944
rect 18699 895 18741 904
rect 18700 80 18740 895
rect 18892 80 18932 1315
rect 19083 1280 19125 1289
rect 19083 1240 19084 1280
rect 19124 1240 19125 1280
rect 19083 1231 19125 1240
rect 18987 1112 19029 1121
rect 18987 1072 18988 1112
rect 19028 1072 19029 1112
rect 18987 1063 19029 1072
rect 18988 617 19028 1063
rect 18987 608 19029 617
rect 18987 568 18988 608
rect 19028 568 19029 608
rect 18987 559 19029 568
rect 19084 80 19124 1231
rect 19276 953 19316 1651
rect 19275 944 19317 953
rect 19275 904 19276 944
rect 19316 904 19317 944
rect 19275 895 19317 904
rect 19372 776 19412 1903
rect 19852 1868 19892 2239
rect 20427 2120 20469 2129
rect 20427 2080 20428 2120
rect 20468 2080 20469 2120
rect 20427 2071 20469 2080
rect 20332 1952 20372 1961
rect 19852 1819 19892 1828
rect 20235 1868 20277 1877
rect 20235 1828 20236 1868
rect 20276 1828 20277 1868
rect 20235 1819 20277 1828
rect 19659 1700 19701 1709
rect 20044 1700 20084 1709
rect 19659 1660 19660 1700
rect 19700 1660 19701 1700
rect 19659 1651 19701 1660
rect 19948 1660 20044 1700
rect 19660 1373 19700 1651
rect 19659 1364 19701 1373
rect 19659 1324 19660 1364
rect 19700 1324 19701 1364
rect 19659 1315 19701 1324
rect 19659 860 19701 869
rect 19659 820 19660 860
rect 19700 820 19701 860
rect 19659 811 19701 820
rect 19276 736 19412 776
rect 19276 80 19316 736
rect 19660 80 19700 811
rect 19851 608 19893 617
rect 19851 568 19852 608
rect 19892 568 19893 608
rect 19948 608 19988 1660
rect 20044 1651 20084 1660
rect 20043 1448 20085 1457
rect 20043 1408 20044 1448
rect 20084 1408 20085 1448
rect 20043 1399 20085 1408
rect 20044 1070 20084 1399
rect 20236 1364 20276 1819
rect 20140 1324 20276 1364
rect 20332 1364 20372 1912
rect 20428 1952 20468 2071
rect 20428 1903 20468 1912
rect 20428 1364 20468 1373
rect 20332 1324 20428 1364
rect 20140 1205 20180 1324
rect 20428 1315 20468 1324
rect 20139 1196 20181 1205
rect 20139 1156 20140 1196
rect 20180 1156 20181 1196
rect 20139 1147 20181 1156
rect 20236 1112 20276 1121
rect 20331 1112 20373 1121
rect 20276 1072 20332 1112
rect 20372 1072 20373 1112
rect 20236 1070 20276 1072
rect 20044 1030 20276 1070
rect 20331 1063 20373 1072
rect 20048 776 20416 785
rect 20088 736 20130 776
rect 20170 736 20212 776
rect 20252 736 20294 776
rect 20334 736 20376 776
rect 20048 727 20416 736
rect 20524 608 20564 2416
rect 20715 2456 20757 2465
rect 20715 2416 20716 2456
rect 20756 2416 20757 2456
rect 20715 2407 20757 2416
rect 20716 1961 20756 2407
rect 20715 1952 20757 1961
rect 20715 1912 20716 1952
rect 20756 1912 20757 1952
rect 20715 1903 20757 1912
rect 20812 1868 20852 1877
rect 20812 1709 20852 1828
rect 20907 1868 20949 1877
rect 20907 1828 20908 1868
rect 20948 1828 20949 1868
rect 20907 1819 20949 1828
rect 20908 1734 20948 1819
rect 20811 1700 20853 1709
rect 20811 1660 20812 1700
rect 20852 1660 20853 1700
rect 20811 1651 20853 1660
rect 20811 1364 20853 1373
rect 20811 1324 20812 1364
rect 20852 1324 20853 1364
rect 20811 1315 20853 1324
rect 20715 1280 20757 1289
rect 20715 1240 20716 1280
rect 20756 1240 20757 1280
rect 20715 1231 20757 1240
rect 20716 1112 20756 1231
rect 20716 1063 20756 1072
rect 20619 776 20661 785
rect 20619 736 20620 776
rect 20660 736 20661 776
rect 20619 727 20661 736
rect 19948 568 20084 608
rect 19851 559 19893 568
rect 19852 80 19892 559
rect 20044 80 20084 568
rect 20428 568 20564 608
rect 20235 188 20277 197
rect 20235 148 20236 188
rect 20276 148 20277 188
rect 20235 139 20277 148
rect 20236 80 20276 139
rect 20428 80 20468 568
rect 20620 80 20660 727
rect 20812 80 20852 1315
rect 21004 80 21044 3415
rect 21100 2456 21140 2465
rect 21100 1205 21140 2416
rect 21196 1877 21236 3919
rect 21388 3809 21428 7036
rect 21579 7027 21621 7036
rect 21579 6656 21621 6665
rect 21579 6616 21580 6656
rect 21620 6616 21621 6656
rect 21579 6607 21621 6616
rect 21580 6488 21620 6607
rect 21580 6439 21620 6448
rect 21676 6488 21716 7111
rect 23212 6992 23252 7001
rect 22732 6952 23212 6992
rect 22059 6740 22101 6749
rect 22059 6700 22060 6740
rect 22100 6700 22101 6740
rect 22059 6691 22101 6700
rect 21676 6439 21716 6448
rect 22060 6488 22100 6691
rect 22060 6439 22100 6448
rect 22635 6488 22677 6497
rect 22635 6448 22636 6488
rect 22676 6448 22677 6488
rect 22635 6439 22677 6448
rect 22155 6404 22197 6413
rect 22155 6364 22156 6404
rect 22196 6364 22197 6404
rect 22155 6355 22197 6364
rect 22156 6270 22196 6355
rect 22636 6354 22676 6439
rect 22059 5732 22101 5741
rect 22059 5692 22060 5732
rect 22100 5692 22101 5732
rect 22059 5683 22101 5692
rect 21675 5648 21717 5657
rect 21675 5608 21676 5648
rect 21716 5608 21717 5648
rect 21675 5599 21717 5608
rect 22060 5648 22100 5683
rect 21676 4976 21716 5599
rect 22060 5597 22100 5608
rect 22155 5228 22197 5237
rect 22155 5188 22156 5228
rect 22196 5188 22197 5228
rect 22155 5179 22197 5188
rect 21676 4927 21716 4936
rect 21483 4808 21525 4817
rect 21483 4768 21484 4808
rect 21524 4768 21525 4808
rect 21483 4759 21525 4768
rect 21387 3800 21429 3809
rect 21387 3760 21388 3800
rect 21428 3760 21429 3800
rect 21387 3751 21429 3760
rect 21291 3632 21333 3641
rect 21291 3592 21292 3632
rect 21332 3592 21333 3632
rect 21484 3632 21524 4759
rect 21580 4136 21620 4147
rect 21580 4061 21620 4096
rect 21675 4136 21717 4145
rect 21675 4096 21676 4136
rect 21716 4096 21717 4136
rect 21675 4087 21717 4096
rect 22156 4136 22196 5179
rect 22347 4388 22389 4397
rect 22347 4348 22348 4388
rect 22388 4348 22389 4388
rect 22347 4339 22389 4348
rect 22156 4087 22196 4096
rect 21579 4052 21621 4061
rect 21579 4012 21580 4052
rect 21620 4012 21621 4052
rect 21579 4003 21621 4012
rect 21676 4002 21716 4087
rect 21484 3592 21620 3632
rect 21291 3583 21333 3592
rect 21195 1868 21237 1877
rect 21195 1828 21196 1868
rect 21236 1828 21237 1868
rect 21195 1819 21237 1828
rect 21195 1280 21237 1289
rect 21195 1240 21196 1280
rect 21236 1240 21237 1280
rect 21292 1280 21332 3583
rect 21388 3464 21428 3473
rect 21483 3464 21525 3473
rect 21428 3424 21484 3464
rect 21524 3424 21525 3464
rect 21388 3415 21428 3424
rect 21483 3415 21525 3424
rect 21484 2708 21524 2717
rect 21484 2045 21524 2668
rect 21483 2036 21525 2045
rect 21483 1996 21484 2036
rect 21524 1996 21525 2036
rect 21483 1987 21525 1996
rect 21387 1952 21429 1961
rect 21387 1912 21388 1952
rect 21428 1912 21429 1952
rect 21387 1903 21429 1912
rect 21388 1818 21428 1903
rect 21292 1240 21428 1280
rect 21195 1231 21237 1240
rect 21099 1196 21141 1205
rect 21099 1156 21100 1196
rect 21140 1156 21141 1196
rect 21099 1147 21141 1156
rect 21196 80 21236 1231
rect 21388 80 21428 1240
rect 21580 80 21620 3592
rect 22156 2708 22196 2717
rect 21676 2456 21716 2465
rect 21676 1037 21716 2416
rect 21964 2456 22004 2465
rect 21868 1938 21908 1947
rect 21868 1373 21908 1898
rect 21867 1364 21909 1373
rect 21867 1324 21868 1364
rect 21908 1324 21909 1364
rect 21964 1364 22004 2416
rect 22060 2120 22100 2129
rect 22156 2120 22196 2668
rect 22100 2080 22196 2120
rect 22060 2071 22100 2080
rect 22155 1364 22197 1373
rect 21964 1324 22100 1364
rect 21867 1315 21909 1324
rect 21771 1196 21813 1205
rect 21771 1156 21772 1196
rect 21812 1156 21813 1196
rect 21771 1147 21813 1156
rect 21675 1028 21717 1037
rect 21675 988 21676 1028
rect 21716 988 21717 1028
rect 21675 979 21717 988
rect 21772 80 21812 1147
rect 21964 1121 22004 1206
rect 21963 1112 22005 1121
rect 21963 1072 21964 1112
rect 22004 1072 22005 1112
rect 21963 1063 22005 1072
rect 22060 944 22100 1324
rect 22155 1324 22156 1364
rect 22196 1324 22197 1364
rect 22155 1315 22197 1324
rect 22156 1230 22196 1315
rect 22155 1028 22197 1037
rect 22155 988 22156 1028
rect 22196 988 22197 1028
rect 22155 979 22197 988
rect 21964 904 22100 944
rect 21964 80 22004 904
rect 22156 80 22196 979
rect 22348 80 22388 4339
rect 22636 4141 22676 4150
rect 22636 3641 22676 4101
rect 22635 3632 22677 3641
rect 22635 3592 22636 3632
rect 22676 3592 22677 3632
rect 22635 3583 22677 3592
rect 22443 3464 22485 3473
rect 22443 3424 22444 3464
rect 22484 3424 22485 3464
rect 22443 3415 22485 3424
rect 22635 3464 22677 3473
rect 22635 3424 22636 3464
rect 22676 3424 22677 3464
rect 22635 3415 22677 3424
rect 22444 3305 22484 3415
rect 22636 3330 22676 3415
rect 22443 3296 22485 3305
rect 22443 3256 22444 3296
rect 22484 3256 22485 3296
rect 22443 3247 22485 3256
rect 22444 1952 22484 3247
rect 22444 1903 22484 1912
rect 22539 356 22581 365
rect 22539 316 22540 356
rect 22580 316 22581 356
rect 22539 307 22581 316
rect 22540 80 22580 307
rect 22732 80 22772 6952
rect 23212 6943 23252 6952
rect 23308 6572 23348 6581
rect 23348 6532 23732 6572
rect 23308 6523 23348 6532
rect 23164 6446 23204 6455
rect 23164 6404 23204 6406
rect 23692 6404 23732 6532
rect 23164 6364 23444 6404
rect 23404 5900 23444 6364
rect 23692 6355 23732 6364
rect 23500 6236 23540 6245
rect 23540 6196 23636 6236
rect 23500 6187 23540 6196
rect 23500 5900 23540 5909
rect 23404 5860 23500 5900
rect 23500 5851 23540 5860
rect 23308 5648 23348 5657
rect 23308 5321 23348 5608
rect 22923 5312 22965 5321
rect 22923 5272 22924 5312
rect 22964 5272 22965 5312
rect 22923 5263 22965 5272
rect 23307 5312 23349 5321
rect 23307 5272 23308 5312
rect 23348 5272 23349 5312
rect 23307 5263 23349 5272
rect 22924 4985 22964 5263
rect 23499 5144 23541 5153
rect 23499 5104 23500 5144
rect 23540 5104 23541 5144
rect 23499 5095 23541 5104
rect 23019 5060 23061 5069
rect 23019 5020 23020 5060
rect 23060 5020 23061 5060
rect 23019 5011 23061 5020
rect 23116 5060 23156 5069
rect 23156 5020 23444 5060
rect 23116 5011 23156 5020
rect 22923 4976 22965 4985
rect 22923 4936 22924 4976
rect 22964 4936 22965 4976
rect 22923 4927 22965 4936
rect 22924 4842 22964 4927
rect 23020 4220 23060 5011
rect 23404 4976 23444 5020
rect 23404 4927 23444 4936
rect 23500 4976 23540 5095
rect 23500 4388 23540 4936
rect 23596 4397 23636 6196
rect 23884 5648 23924 7699
rect 24268 7614 24308 7699
rect 24171 7160 24213 7169
rect 24171 7120 24172 7160
rect 24212 7120 24213 7160
rect 24171 7111 24213 7120
rect 24172 6665 24212 7111
rect 24171 6656 24213 6665
rect 24171 6616 24172 6656
rect 24212 6616 24213 6656
rect 24171 6607 24213 6616
rect 24364 6488 24404 8371
rect 25996 8168 26036 8632
rect 25228 8128 25460 8168
rect 24939 8084 24981 8093
rect 24939 8044 24940 8084
rect 24980 8044 24981 8084
rect 24939 8035 24981 8044
rect 24555 7916 24597 7925
rect 24555 7876 24556 7916
rect 24596 7876 24597 7916
rect 24555 7867 24597 7876
rect 24364 6439 24404 6448
rect 24459 6068 24501 6077
rect 24459 6028 24460 6068
rect 24500 6028 24501 6068
rect 24459 6019 24501 6028
rect 24460 5732 24500 6019
rect 24460 5683 24500 5692
rect 23884 5599 23924 5608
rect 23980 5648 24020 5657
rect 23980 5153 24020 5608
rect 24364 5648 24404 5657
rect 23979 5144 24021 5153
rect 23979 5104 23980 5144
rect 24020 5104 24021 5144
rect 23979 5095 24021 5104
rect 23980 4985 24020 5016
rect 23979 4976 24021 4985
rect 23979 4936 23980 4976
rect 24020 4936 24021 4976
rect 23979 4927 24021 4936
rect 23883 4892 23925 4901
rect 23883 4852 23884 4892
rect 23924 4852 23925 4892
rect 23883 4843 23925 4852
rect 23980 4892 24020 4927
rect 23884 4758 23924 4843
rect 23691 4556 23733 4565
rect 23691 4516 23692 4556
rect 23732 4516 23733 4556
rect 23691 4507 23733 4516
rect 23308 4348 23540 4388
rect 23595 4388 23637 4397
rect 23595 4348 23596 4388
rect 23636 4348 23637 4388
rect 23212 4220 23252 4229
rect 23020 4180 23212 4220
rect 23212 4171 23252 4180
rect 23308 4052 23348 4348
rect 23595 4339 23637 4348
rect 23500 4220 23540 4229
rect 23116 4012 23348 4052
rect 23404 4180 23500 4220
rect 22828 3968 22868 3977
rect 23020 3968 23060 3977
rect 22868 3928 22964 3968
rect 22828 3919 22868 3928
rect 22827 3632 22869 3641
rect 22827 3592 22828 3632
rect 22868 3592 22869 3632
rect 22827 3583 22869 3592
rect 22828 3498 22868 3583
rect 22924 2708 22964 3928
rect 22924 2659 22964 2668
rect 22924 1205 22964 1290
rect 22923 1196 22965 1205
rect 22923 1156 22924 1196
rect 22964 1156 22965 1196
rect 22923 1147 22965 1156
rect 23020 1028 23060 3928
rect 23116 3053 23156 4012
rect 23404 3809 23444 4180
rect 23500 4171 23540 4180
rect 23692 4136 23732 4507
rect 23980 4313 24020 4852
rect 24075 4892 24117 4901
rect 24075 4852 24076 4892
rect 24116 4852 24117 4892
rect 24075 4843 24117 4852
rect 24076 4481 24116 4843
rect 24267 4808 24309 4817
rect 24267 4768 24268 4808
rect 24308 4768 24309 4808
rect 24267 4759 24309 4768
rect 24171 4640 24213 4649
rect 24171 4600 24172 4640
rect 24212 4600 24213 4640
rect 24171 4591 24213 4600
rect 24075 4472 24117 4481
rect 24075 4432 24076 4472
rect 24116 4432 24117 4472
rect 24075 4423 24117 4432
rect 23979 4304 24021 4313
rect 23979 4264 23980 4304
rect 24020 4264 24021 4304
rect 23979 4255 24021 4264
rect 24075 4220 24117 4229
rect 24075 4180 24076 4220
rect 24116 4180 24117 4220
rect 24075 4171 24117 4180
rect 23596 4096 23732 4136
rect 23403 3800 23445 3809
rect 23403 3760 23404 3800
rect 23444 3760 23445 3800
rect 23403 3751 23445 3760
rect 23307 3548 23349 3557
rect 23307 3508 23308 3548
rect 23348 3508 23349 3548
rect 23307 3499 23349 3508
rect 23499 3548 23541 3557
rect 23499 3508 23500 3548
rect 23540 3508 23541 3548
rect 23499 3499 23541 3508
rect 23211 3464 23253 3473
rect 23211 3424 23212 3464
rect 23252 3424 23253 3464
rect 23211 3415 23253 3424
rect 23212 3330 23252 3415
rect 23115 3044 23157 3053
rect 23115 3004 23116 3044
rect 23156 3004 23157 3044
rect 23115 2995 23157 3004
rect 23211 2792 23253 2801
rect 23211 2752 23212 2792
rect 23252 2752 23253 2792
rect 23211 2743 23253 2752
rect 23212 2540 23252 2743
rect 23308 2708 23348 3499
rect 23308 2659 23348 2668
rect 23500 2633 23540 3499
rect 23596 3296 23636 4096
rect 24076 4086 24116 4171
rect 23692 3968 23732 3977
rect 23884 3968 23924 3977
rect 23692 3557 23732 3928
rect 23788 3928 23884 3968
rect 23691 3548 23733 3557
rect 23691 3508 23692 3548
rect 23732 3508 23733 3548
rect 23691 3499 23733 3508
rect 23596 3256 23732 3296
rect 23595 2960 23637 2969
rect 23595 2920 23596 2960
rect 23636 2920 23637 2960
rect 23595 2911 23637 2920
rect 23499 2624 23541 2633
rect 23499 2584 23500 2624
rect 23540 2584 23541 2624
rect 23499 2575 23541 2584
rect 23212 2500 23348 2540
rect 23116 2456 23156 2465
rect 23156 2416 23252 2456
rect 23116 2407 23156 2416
rect 22924 988 23060 1028
rect 22924 80 22964 988
rect 23116 953 23156 1038
rect 23115 944 23157 953
rect 23115 904 23116 944
rect 23156 904 23157 944
rect 23115 895 23157 904
rect 23212 776 23252 2416
rect 23308 1205 23348 2500
rect 23500 2456 23540 2465
rect 23403 2120 23445 2129
rect 23403 2080 23404 2120
rect 23444 2080 23445 2120
rect 23403 2071 23445 2080
rect 23307 1196 23349 1205
rect 23307 1156 23308 1196
rect 23348 1156 23349 1196
rect 23307 1147 23349 1156
rect 23404 776 23444 2071
rect 23500 1709 23540 2416
rect 23499 1700 23541 1709
rect 23499 1660 23500 1700
rect 23540 1660 23541 1700
rect 23499 1651 23541 1660
rect 23499 1280 23541 1289
rect 23499 1240 23500 1280
rect 23540 1240 23541 1280
rect 23499 1231 23541 1240
rect 23500 1070 23540 1231
rect 23500 1021 23540 1030
rect 23596 944 23636 2911
rect 23692 1952 23732 3256
rect 23788 2969 23828 3928
rect 23884 3919 23924 3928
rect 23979 3884 24021 3893
rect 23979 3844 23980 3884
rect 24020 3844 24021 3884
rect 23979 3835 24021 3844
rect 23883 3800 23925 3809
rect 23883 3760 23884 3800
rect 23924 3760 23925 3800
rect 23883 3751 23925 3760
rect 23787 2960 23829 2969
rect 23787 2920 23788 2960
rect 23828 2920 23829 2960
rect 23787 2911 23829 2920
rect 23788 2624 23828 2633
rect 23788 2036 23828 2584
rect 23884 2297 23924 3751
rect 23883 2288 23925 2297
rect 23883 2248 23884 2288
rect 23924 2248 23925 2288
rect 23883 2239 23925 2248
rect 23884 2036 23924 2045
rect 23788 1996 23884 2036
rect 23884 1987 23924 1996
rect 23692 1903 23732 1912
rect 23691 1700 23733 1709
rect 23691 1660 23692 1700
rect 23732 1660 23733 1700
rect 23691 1651 23733 1660
rect 23883 1700 23925 1709
rect 23883 1660 23884 1700
rect 23924 1660 23925 1700
rect 23883 1651 23925 1660
rect 23692 1289 23732 1651
rect 23691 1280 23733 1289
rect 23691 1240 23692 1280
rect 23732 1240 23733 1280
rect 23691 1231 23733 1240
rect 23116 736 23252 776
rect 23308 736 23444 776
rect 23500 904 23636 944
rect 23691 944 23733 953
rect 23691 904 23692 944
rect 23732 904 23733 944
rect 23116 80 23156 736
rect 23308 80 23348 736
rect 23500 80 23540 904
rect 23691 895 23733 904
rect 23692 80 23732 895
rect 23884 80 23924 1651
rect 23980 365 24020 3835
rect 24172 3389 24212 4591
rect 24268 4388 24308 4759
rect 24364 4733 24404 5608
rect 24460 4976 24500 4987
rect 24460 4901 24500 4936
rect 24459 4892 24501 4901
rect 24459 4852 24460 4892
rect 24500 4852 24501 4892
rect 24459 4843 24501 4852
rect 24363 4724 24405 4733
rect 24363 4684 24364 4724
rect 24404 4684 24405 4724
rect 24363 4675 24405 4684
rect 24268 4339 24308 4348
rect 24460 4136 24500 4145
rect 24460 3809 24500 4096
rect 24459 3800 24501 3809
rect 24459 3760 24460 3800
rect 24500 3760 24501 3800
rect 24459 3751 24501 3760
rect 24459 3464 24501 3473
rect 24459 3424 24460 3464
rect 24500 3424 24501 3464
rect 24459 3415 24501 3424
rect 24171 3380 24213 3389
rect 24171 3340 24172 3380
rect 24212 3340 24213 3380
rect 24171 3331 24213 3340
rect 24460 3330 24500 3415
rect 24075 3044 24117 3053
rect 24075 3004 24076 3044
rect 24116 3004 24117 3044
rect 24075 2995 24117 3004
rect 24076 2624 24116 2995
rect 24171 2960 24213 2969
rect 24171 2920 24172 2960
rect 24212 2920 24213 2960
rect 24171 2911 24213 2920
rect 24076 2575 24116 2584
rect 24172 2624 24212 2911
rect 24460 2792 24500 2801
rect 24172 2575 24212 2584
rect 24268 2752 24460 2792
rect 24268 1868 24308 2752
rect 24460 2743 24500 2752
rect 24459 2624 24501 2633
rect 24459 2584 24460 2624
rect 24500 2584 24501 2624
rect 24459 2575 24501 2584
rect 24268 1819 24308 1828
rect 24076 1700 24116 1709
rect 24116 1660 24212 1700
rect 24076 1651 24116 1660
rect 24075 1280 24117 1289
rect 24075 1240 24076 1280
rect 24116 1240 24117 1280
rect 24075 1231 24117 1240
rect 23979 356 24021 365
rect 23979 316 23980 356
rect 24020 316 24021 356
rect 23979 307 24021 316
rect 24076 80 24116 1231
rect 24172 617 24212 1660
rect 24267 1280 24309 1289
rect 24267 1240 24268 1280
rect 24308 1240 24309 1280
rect 24267 1231 24309 1240
rect 24171 608 24213 617
rect 24171 568 24172 608
rect 24212 568 24213 608
rect 24171 559 24213 568
rect 24268 80 24308 1231
rect 24460 80 24500 2575
rect 24556 2540 24596 7867
rect 24940 5648 24980 8035
rect 25228 6917 25268 8128
rect 25324 8000 25364 8009
rect 25324 7496 25364 7960
rect 25420 8000 25460 8128
rect 25420 7951 25460 7960
rect 25804 8128 26036 8168
rect 26380 8632 26476 8672
rect 25804 7916 25844 8128
rect 26380 8093 26420 8632
rect 26476 8623 26516 8632
rect 26571 8672 26613 8681
rect 26571 8632 26572 8672
rect 26612 8632 26613 8672
rect 27531 8672 27573 8681
rect 27044 8641 27284 8672
rect 27004 8632 27284 8641
rect 26571 8623 26613 8632
rect 26379 8084 26421 8093
rect 26379 8044 26380 8084
rect 26420 8044 26421 8084
rect 26379 8035 26421 8044
rect 25899 8000 25941 8009
rect 25899 7960 25900 8000
rect 25940 7960 25941 8000
rect 25899 7951 25941 7960
rect 26380 8000 26420 8035
rect 25324 7456 25652 7496
rect 25612 7412 25652 7456
rect 25612 7363 25652 7372
rect 25419 7160 25461 7169
rect 25419 7120 25420 7160
rect 25460 7120 25461 7160
rect 25419 7111 25461 7120
rect 25611 7160 25653 7169
rect 25611 7120 25612 7160
rect 25652 7120 25653 7160
rect 25611 7111 25653 7120
rect 25420 7026 25460 7111
rect 25227 6908 25269 6917
rect 25227 6868 25228 6908
rect 25268 6868 25269 6908
rect 25227 6859 25269 6868
rect 25228 5825 25268 6859
rect 25612 6488 25652 7111
rect 25804 6488 25844 7876
rect 25900 7866 25940 7951
rect 26380 7949 26420 7960
rect 26379 7748 26421 7757
rect 26379 7708 26380 7748
rect 26420 7708 26421 7748
rect 26379 7699 26421 7708
rect 26283 7580 26325 7589
rect 26283 7540 26284 7580
rect 26324 7540 26325 7580
rect 26283 7531 26325 7540
rect 26284 7412 26324 7531
rect 26284 7363 26324 7372
rect 25900 7244 25940 7253
rect 25900 7001 25940 7204
rect 25899 6992 25941 7001
rect 25899 6952 25900 6992
rect 25940 6952 25941 6992
rect 25899 6943 25941 6952
rect 26092 6992 26132 7001
rect 26283 6992 26325 7001
rect 26132 6952 26228 6992
rect 26092 6943 26132 6952
rect 25995 6740 26037 6749
rect 25995 6700 25996 6740
rect 26036 6700 26037 6740
rect 25995 6691 26037 6700
rect 25804 6448 25940 6488
rect 25612 6439 25652 6448
rect 25323 6404 25365 6413
rect 25323 6364 25324 6404
rect 25364 6364 25365 6404
rect 25323 6355 25365 6364
rect 25227 5816 25269 5825
rect 25227 5776 25228 5816
rect 25268 5776 25269 5816
rect 25227 5767 25269 5776
rect 24844 5608 24940 5648
rect 24747 5396 24789 5405
rect 24747 5356 24748 5396
rect 24788 5356 24789 5396
rect 24747 5347 24789 5356
rect 24748 3725 24788 5347
rect 24844 4901 24884 5608
rect 24940 5599 24980 5608
rect 25324 5564 25364 6355
rect 25804 6236 25844 6245
rect 25612 6196 25804 6236
rect 25468 5690 25508 5699
rect 25612 5690 25652 6196
rect 25804 6187 25844 6196
rect 25508 5650 25652 5690
rect 25468 5641 25508 5650
rect 25324 5524 25460 5564
rect 25132 5060 25172 5069
rect 24940 4962 24980 4971
rect 24843 4892 24885 4901
rect 24843 4852 24844 4892
rect 24884 4852 24885 4892
rect 24843 4843 24885 4852
rect 24940 4817 24980 4922
rect 24939 4808 24981 4817
rect 24939 4768 24940 4808
rect 24980 4768 24981 4808
rect 24939 4759 24981 4768
rect 25132 4229 25172 5020
rect 25324 4724 25364 4733
rect 25228 4684 25324 4724
rect 25131 4220 25173 4229
rect 25131 4180 25132 4220
rect 25172 4180 25173 4220
rect 25131 4171 25173 4180
rect 24747 3716 24789 3725
rect 24747 3676 24748 3716
rect 24788 3676 24789 3716
rect 24747 3667 24789 3676
rect 24652 3548 24692 3557
rect 24692 3508 24980 3548
rect 24652 3499 24692 3508
rect 24940 3464 24980 3508
rect 24940 3415 24980 3424
rect 25036 3464 25076 3473
rect 25076 3424 25172 3464
rect 25036 3415 25076 3424
rect 24651 3380 24693 3389
rect 24651 3340 24652 3380
rect 24692 3340 24693 3380
rect 24651 3331 24693 3340
rect 24652 2708 24692 3331
rect 25132 2801 25172 3424
rect 24747 2792 24789 2801
rect 24747 2752 24748 2792
rect 24788 2752 24789 2792
rect 24747 2743 24789 2752
rect 25131 2792 25173 2801
rect 25131 2752 25132 2792
rect 25172 2752 25173 2792
rect 25131 2743 25173 2752
rect 24652 2659 24692 2668
rect 24556 2500 24692 2540
rect 24555 2288 24597 2297
rect 24555 2248 24556 2288
rect 24596 2248 24597 2288
rect 24555 2239 24597 2248
rect 24556 953 24596 2239
rect 24555 944 24597 953
rect 24555 904 24556 944
rect 24596 904 24597 944
rect 24555 895 24597 904
rect 24652 80 24692 2500
rect 24748 2288 24788 2743
rect 24844 2456 24884 2465
rect 24884 2416 24980 2456
rect 24844 2407 24884 2416
rect 24940 2297 24980 2416
rect 24939 2288 24981 2297
rect 24748 2248 24884 2288
rect 24748 1952 24788 1961
rect 24748 1700 24788 1912
rect 24844 1952 24884 2248
rect 24939 2248 24940 2288
rect 24980 2248 24981 2288
rect 24939 2239 24981 2248
rect 25228 2036 25268 4684
rect 25324 4675 25364 4684
rect 25323 3548 25365 3557
rect 25323 3508 25324 3548
rect 25364 3508 25365 3548
rect 25323 3499 25365 3508
rect 25324 2708 25364 3499
rect 25420 3464 25460 5524
rect 25612 5480 25652 5489
rect 25516 5440 25612 5480
rect 25516 4892 25556 5440
rect 25612 5431 25652 5440
rect 25611 5144 25653 5153
rect 25611 5104 25612 5144
rect 25652 5104 25653 5144
rect 25611 5095 25653 5104
rect 25516 4843 25556 4852
rect 25515 3632 25557 3641
rect 25515 3592 25516 3632
rect 25556 3592 25557 3632
rect 25515 3583 25557 3592
rect 25420 3415 25460 3424
rect 25516 3464 25556 3583
rect 25516 3415 25556 3424
rect 25612 3212 25652 5095
rect 25900 4985 25940 6448
rect 25899 4976 25941 4985
rect 25899 4936 25900 4976
rect 25940 4936 25941 4976
rect 25899 4927 25941 4936
rect 25707 4892 25749 4901
rect 25707 4852 25708 4892
rect 25748 4852 25749 4892
rect 25707 4843 25749 4852
rect 25708 4229 25748 4843
rect 25707 4220 25749 4229
rect 25707 4180 25708 4220
rect 25748 4180 25749 4220
rect 25707 4171 25749 4180
rect 25708 4136 25748 4171
rect 25708 4085 25748 4096
rect 25707 3716 25749 3725
rect 25707 3676 25708 3716
rect 25748 3676 25749 3716
rect 25707 3667 25749 3676
rect 25324 2659 25364 2668
rect 25420 3172 25652 3212
rect 24844 1903 24884 1912
rect 25132 1996 25268 2036
rect 24748 1660 24980 1700
rect 24940 1364 24980 1660
rect 24940 1315 24980 1324
rect 25132 1289 25172 1996
rect 25324 1961 25364 2046
rect 25323 1952 25365 1961
rect 25323 1912 25324 1952
rect 25364 1912 25365 1952
rect 25323 1903 25365 1912
rect 25228 1868 25268 1877
rect 25131 1280 25173 1289
rect 25131 1240 25132 1280
rect 25172 1240 25173 1280
rect 25131 1231 25173 1240
rect 24747 1196 24789 1205
rect 24747 1156 24748 1196
rect 24788 1156 24789 1196
rect 24747 1147 24789 1156
rect 24748 1112 24788 1147
rect 24748 1061 24788 1072
rect 24843 944 24885 953
rect 24843 904 24844 944
rect 24884 904 24885 944
rect 24843 895 24885 904
rect 24844 80 24884 895
rect 25035 860 25077 869
rect 25035 820 25036 860
rect 25076 820 25077 860
rect 25035 811 25077 820
rect 25036 80 25076 811
rect 25228 785 25268 1828
rect 25323 1700 25365 1709
rect 25323 1660 25324 1700
rect 25364 1660 25365 1700
rect 25323 1651 25365 1660
rect 25227 776 25269 785
rect 25227 736 25228 776
rect 25268 736 25269 776
rect 25227 727 25269 736
rect 25324 608 25364 1651
rect 25228 568 25364 608
rect 25228 80 25268 568
rect 25420 80 25460 3172
rect 25708 2969 25748 3667
rect 25996 3641 26036 6691
rect 26092 6236 26132 6245
rect 26092 3977 26132 6196
rect 26188 4808 26228 6952
rect 26283 6952 26284 6992
rect 26324 6952 26325 6992
rect 26283 6943 26325 6952
rect 26284 6749 26324 6943
rect 26283 6740 26325 6749
rect 26283 6700 26284 6740
rect 26324 6700 26325 6740
rect 26283 6691 26325 6700
rect 26284 6404 26324 6413
rect 26380 6404 26420 7699
rect 26475 7160 26517 7169
rect 26572 7160 26612 8623
rect 27244 8588 27284 8632
rect 27531 8632 27532 8672
rect 27572 8632 27573 8672
rect 27531 8623 27573 8632
rect 27340 8588 27380 8597
rect 27244 8548 27340 8588
rect 27340 8539 27380 8548
rect 27532 8538 27572 8623
rect 27148 8504 27188 8513
rect 27188 8464 27284 8504
rect 27148 8455 27188 8464
rect 27052 8084 27092 8093
rect 26860 7986 26900 7995
rect 26860 7589 26900 7946
rect 27052 7757 27092 8044
rect 27147 7916 27189 7925
rect 27147 7876 27148 7916
rect 27188 7876 27189 7916
rect 27244 7916 27284 8464
rect 27724 7925 27764 9472
rect 28300 8933 28340 10672
rect 29259 10648 29260 10688
rect 29300 10648 29301 10688
rect 29432 10672 29512 10752
rect 30584 10672 30664 10752
rect 31736 10732 31816 10752
rect 31736 10692 32564 10732
rect 31736 10672 31844 10692
rect 29259 10639 29301 10648
rect 28972 9512 29012 9521
rect 28299 8924 28341 8933
rect 28299 8884 28300 8924
rect 28340 8884 28341 8924
rect 28299 8875 28341 8884
rect 28780 8672 28820 8683
rect 28780 8597 28820 8632
rect 28779 8588 28821 8597
rect 28779 8548 28780 8588
rect 28820 8548 28821 8588
rect 28779 8539 28821 8548
rect 28683 8000 28725 8009
rect 28683 7960 28684 8000
rect 28724 7960 28725 8000
rect 28683 7951 28725 7960
rect 28780 8000 28820 8009
rect 27436 7916 27476 7925
rect 27244 7876 27436 7916
rect 27147 7867 27189 7876
rect 27436 7867 27476 7876
rect 27723 7916 27765 7925
rect 27723 7876 27724 7916
rect 27764 7876 27765 7916
rect 27723 7867 27765 7876
rect 28395 7916 28437 7925
rect 28395 7876 28396 7916
rect 28436 7876 28437 7916
rect 28395 7867 28437 7876
rect 27051 7748 27093 7757
rect 27051 7708 27052 7748
rect 27092 7708 27093 7748
rect 27148 7748 27188 7867
rect 27244 7748 27284 7757
rect 27148 7708 27244 7748
rect 27051 7699 27093 7708
rect 27244 7699 27284 7708
rect 26859 7580 26901 7589
rect 26859 7540 26860 7580
rect 26900 7540 26901 7580
rect 26859 7531 26901 7540
rect 27723 7412 27765 7421
rect 27723 7372 27724 7412
rect 27764 7372 27765 7412
rect 27723 7363 27765 7372
rect 27724 7169 27764 7363
rect 26475 7120 26476 7160
rect 26516 7120 26612 7160
rect 26475 7111 26517 7120
rect 26476 7026 26516 7111
rect 26324 6364 26420 6404
rect 26476 6488 26516 6497
rect 26284 6355 26324 6364
rect 26476 5909 26516 6448
rect 26475 5900 26517 5909
rect 26475 5860 26476 5900
rect 26516 5860 26517 5900
rect 26475 5851 26517 5860
rect 26476 5741 26516 5851
rect 26475 5732 26517 5741
rect 26475 5692 26476 5732
rect 26516 5692 26517 5732
rect 26475 5683 26517 5692
rect 26380 4985 26420 5070
rect 26379 4976 26421 4985
rect 26379 4936 26380 4976
rect 26420 4936 26421 4976
rect 26379 4927 26421 4936
rect 26188 4768 26420 4808
rect 26091 3968 26133 3977
rect 26091 3928 26092 3968
rect 26132 3928 26133 3968
rect 26091 3919 26133 3928
rect 26091 3800 26133 3809
rect 26091 3760 26092 3800
rect 26132 3760 26133 3800
rect 26091 3751 26133 3760
rect 25995 3632 26037 3641
rect 25995 3592 25996 3632
rect 26036 3592 26037 3632
rect 25995 3583 26037 3592
rect 25995 3464 26037 3473
rect 25995 3424 25996 3464
rect 26036 3424 26037 3464
rect 25995 3415 26037 3424
rect 25996 3053 26036 3415
rect 25803 3044 25845 3053
rect 25803 3004 25804 3044
rect 25844 3004 25845 3044
rect 25803 2995 25845 3004
rect 25995 3044 26037 3053
rect 25995 3004 25996 3044
rect 26036 3004 26037 3044
rect 25995 2995 26037 3004
rect 25707 2960 25749 2969
rect 25707 2920 25708 2960
rect 25748 2920 25749 2960
rect 25707 2911 25749 2920
rect 25708 2624 25748 2911
rect 25708 2575 25748 2584
rect 25516 2456 25556 2465
rect 25516 944 25556 2416
rect 25804 1952 25844 2995
rect 26092 2540 26132 3751
rect 26283 3212 26325 3221
rect 26283 3172 26284 3212
rect 26324 3172 26325 3212
rect 26283 3163 26325 3172
rect 26187 2708 26229 2717
rect 26187 2668 26188 2708
rect 26228 2668 26229 2708
rect 26187 2659 26229 2668
rect 25804 1903 25844 1912
rect 25996 2500 26132 2540
rect 25611 1364 25653 1373
rect 25611 1324 25612 1364
rect 25652 1324 25653 1364
rect 25611 1315 25653 1324
rect 25612 1230 25652 1315
rect 25707 1196 25749 1205
rect 25707 1156 25708 1196
rect 25748 1156 25844 1196
rect 25707 1147 25749 1156
rect 25804 1154 25844 1156
rect 25804 1105 25844 1114
rect 25516 904 25844 944
rect 25611 272 25653 281
rect 25611 232 25612 272
rect 25652 232 25653 272
rect 25611 223 25653 232
rect 25612 80 25652 223
rect 25804 80 25844 904
rect 25996 80 26036 2500
rect 26091 2204 26133 2213
rect 26091 2164 26092 2204
rect 26132 2164 26133 2204
rect 26091 2155 26133 2164
rect 26092 1205 26132 2155
rect 26091 1196 26133 1205
rect 26091 1156 26092 1196
rect 26132 1156 26133 1196
rect 26091 1147 26133 1156
rect 26188 80 26228 2659
rect 26284 2036 26324 3163
rect 26380 2213 26420 4768
rect 26572 3725 26612 7120
rect 27723 7160 27765 7169
rect 27723 7120 27724 7160
rect 27764 7120 27765 7160
rect 27723 7111 27765 7120
rect 27724 7026 27764 7111
rect 27724 6532 28052 6572
rect 27724 6488 27764 6532
rect 27724 6404 27764 6448
rect 28012 6413 28052 6532
rect 28299 6488 28341 6497
rect 28299 6448 28300 6488
rect 28340 6448 28341 6488
rect 28299 6439 28341 6448
rect 27532 6364 27764 6404
rect 28011 6404 28053 6413
rect 28011 6364 28012 6404
rect 28052 6364 28053 6404
rect 26955 6320 26997 6329
rect 26955 6280 26956 6320
rect 26996 6280 26997 6320
rect 26955 6271 26997 6280
rect 26860 5732 26900 5741
rect 26860 5573 26900 5692
rect 26859 5564 26901 5573
rect 26859 5524 26860 5564
rect 26900 5524 26901 5564
rect 26859 5515 26901 5524
rect 26571 3716 26613 3725
rect 26571 3676 26572 3716
rect 26612 3676 26613 3716
rect 26571 3667 26613 3676
rect 26667 3548 26709 3557
rect 26667 3508 26668 3548
rect 26708 3508 26709 3548
rect 26667 3499 26709 3508
rect 26476 3450 26516 3459
rect 26668 3414 26708 3499
rect 26476 3053 26516 3410
rect 26859 3380 26901 3389
rect 26859 3340 26860 3380
rect 26900 3340 26901 3380
rect 26859 3331 26901 3340
rect 26475 3044 26517 3053
rect 26475 3004 26476 3044
rect 26516 3004 26517 3044
rect 26475 2995 26517 3004
rect 26860 2540 26900 3331
rect 26956 2876 26996 6271
rect 27052 5480 27092 5489
rect 27092 5440 27476 5480
rect 27052 5431 27092 5440
rect 27051 5060 27093 5069
rect 27051 5020 27052 5060
rect 27092 5020 27093 5060
rect 27051 5011 27093 5020
rect 27052 4220 27092 5011
rect 27052 4171 27092 4180
rect 27244 3968 27284 3977
rect 27147 3044 27189 3053
rect 27147 3004 27148 3044
rect 27188 3004 27189 3044
rect 27147 2995 27189 3004
rect 27148 2876 27188 2995
rect 26956 2836 27092 2876
rect 26956 2624 26996 2633
rect 26956 2540 26996 2584
rect 26860 2500 26996 2540
rect 27052 2540 27092 2836
rect 27148 2827 27188 2836
rect 27244 2549 27284 3928
rect 27243 2540 27285 2549
rect 27052 2500 27188 2540
rect 26379 2204 26421 2213
rect 26379 2164 26380 2204
rect 26420 2164 26421 2204
rect 26379 2155 26421 2164
rect 26476 2036 26516 2045
rect 26284 1996 26420 2036
rect 26284 1938 26324 1947
rect 26284 1373 26324 1898
rect 26283 1364 26325 1373
rect 26283 1324 26284 1364
rect 26324 1324 26325 1364
rect 26283 1315 26325 1324
rect 26380 80 26420 1996
rect 26516 1996 26900 2036
rect 26476 1987 26516 1996
rect 26860 1868 26900 1996
rect 26860 1819 26900 1828
rect 26668 1700 26708 1709
rect 26668 869 26708 1660
rect 26763 1616 26805 1625
rect 26956 1616 26996 2500
rect 26763 1576 26764 1616
rect 26804 1576 26805 1616
rect 26763 1567 26805 1576
rect 26860 1576 26996 1616
rect 26667 860 26709 869
rect 26667 820 26668 860
rect 26708 820 26709 860
rect 26667 811 26709 820
rect 26571 776 26613 785
rect 26571 736 26572 776
rect 26612 736 26613 776
rect 26571 727 26613 736
rect 26572 80 26612 727
rect 26764 80 26804 1567
rect 26860 1373 26900 1576
rect 26859 1364 26901 1373
rect 26859 1324 26860 1364
rect 26900 1324 26901 1364
rect 26859 1315 26901 1324
rect 26955 1280 26997 1289
rect 26955 1240 26956 1280
rect 26996 1240 26997 1280
rect 26955 1231 26997 1240
rect 26956 80 26996 1231
rect 27052 1112 27092 1121
rect 27052 701 27092 1072
rect 27051 692 27093 701
rect 27051 652 27052 692
rect 27092 652 27093 692
rect 27051 643 27093 652
rect 27052 533 27092 643
rect 27051 524 27093 533
rect 27051 484 27052 524
rect 27092 484 27093 524
rect 27051 475 27093 484
rect 27148 80 27188 2500
rect 27243 2500 27244 2540
rect 27284 2500 27285 2540
rect 27243 2491 27285 2500
rect 27340 2456 27380 2465
rect 27340 1961 27380 2416
rect 27339 1952 27381 1961
rect 27339 1912 27340 1952
rect 27380 1912 27381 1952
rect 27339 1903 27381 1912
rect 27243 1868 27285 1877
rect 27243 1828 27244 1868
rect 27284 1828 27285 1868
rect 27436 1868 27476 5440
rect 27532 4976 27572 6364
rect 28011 6355 28053 6364
rect 28300 6354 28340 6439
rect 27916 6320 27956 6329
rect 27628 6280 27916 6320
rect 27628 5648 27668 6280
rect 27916 6271 27956 6280
rect 27628 5599 27668 5608
rect 27724 5648 27764 5657
rect 27724 5489 27764 5608
rect 28108 5648 28148 5657
rect 27723 5480 27765 5489
rect 27723 5440 27724 5480
rect 27764 5440 27765 5480
rect 27723 5431 27765 5440
rect 27628 4976 27668 4985
rect 27532 4936 27628 4976
rect 27532 4388 27572 4936
rect 27628 4927 27668 4936
rect 27820 4724 27860 4733
rect 27532 4348 27668 4388
rect 27628 4304 27668 4348
rect 27628 4264 27764 4304
rect 27531 4220 27573 4229
rect 27531 4180 27532 4220
rect 27572 4180 27573 4220
rect 27531 4171 27573 4180
rect 27532 4136 27572 4171
rect 27532 4085 27572 4096
rect 27628 4136 27668 4147
rect 27628 4061 27668 4096
rect 27627 4052 27669 4061
rect 27627 4012 27628 4052
rect 27668 4012 27669 4052
rect 27627 4003 27669 4012
rect 27724 3884 27764 4264
rect 27820 4229 27860 4684
rect 27819 4220 27861 4229
rect 27819 4180 27820 4220
rect 27860 4180 27861 4220
rect 27819 4171 27861 4180
rect 28011 4136 28053 4145
rect 28011 4096 28012 4136
rect 28052 4096 28053 4136
rect 28011 4087 28053 4096
rect 28108 4136 28148 5608
rect 28204 5648 28244 5657
rect 28204 5237 28244 5608
rect 28203 5228 28245 5237
rect 28203 5188 28204 5228
rect 28244 5188 28245 5228
rect 28203 5179 28245 5188
rect 28299 4640 28341 4649
rect 28299 4600 28300 4640
rect 28340 4600 28341 4640
rect 28299 4591 28341 4600
rect 28148 4096 28244 4136
rect 28108 4087 28148 4096
rect 28012 4002 28052 4087
rect 27628 3844 27764 3884
rect 27531 3716 27573 3725
rect 27531 3676 27532 3716
rect 27572 3676 27573 3716
rect 27531 3667 27573 3676
rect 27532 2801 27572 3667
rect 27628 3389 27668 3844
rect 28108 3464 28148 3473
rect 27627 3380 27669 3389
rect 27627 3340 27628 3380
rect 27668 3340 27669 3380
rect 27627 3331 27669 3340
rect 28108 3305 28148 3424
rect 28107 3296 28149 3305
rect 28107 3256 28108 3296
rect 28148 3256 28149 3296
rect 28107 3247 28149 3256
rect 27531 2792 27573 2801
rect 27531 2752 27532 2792
rect 27572 2752 27573 2792
rect 27531 2743 27573 2752
rect 27532 2624 27572 2743
rect 27532 2575 27572 2584
rect 28204 2540 28244 4096
rect 28300 3305 28340 4591
rect 28396 4481 28436 7867
rect 28684 7866 28724 7951
rect 28780 7505 28820 7960
rect 28779 7496 28821 7505
rect 28779 7456 28780 7496
rect 28820 7456 28821 7496
rect 28779 7447 28821 7456
rect 28875 7244 28917 7253
rect 28875 7204 28876 7244
rect 28916 7204 28917 7244
rect 28875 7195 28917 7204
rect 28876 7160 28916 7195
rect 28972 7169 29012 9472
rect 29164 9260 29204 9269
rect 29164 8093 29204 9220
rect 29260 8840 29300 10639
rect 29452 9941 29492 10672
rect 29739 10520 29781 10529
rect 29739 10480 29740 10520
rect 29780 10480 29781 10520
rect 29739 10471 29781 10480
rect 29451 9932 29493 9941
rect 29451 9892 29452 9932
rect 29492 9892 29493 9932
rect 29451 9883 29493 9892
rect 29548 9512 29588 9521
rect 29260 8791 29300 8800
rect 29452 9472 29548 9512
rect 29452 8756 29492 9472
rect 29548 9463 29588 9472
rect 29740 8840 29780 10471
rect 30604 9680 30644 10672
rect 31756 10648 31844 10672
rect 32427 10100 32469 10109
rect 32427 10060 32428 10100
rect 32468 10060 32469 10100
rect 32427 10051 32469 10060
rect 32043 10016 32085 10025
rect 32043 9976 32044 10016
rect 32084 9976 32085 10016
rect 32043 9967 32085 9976
rect 32044 9680 32084 9967
rect 30604 9640 30932 9680
rect 29835 9512 29877 9521
rect 29835 9472 29836 9512
rect 29876 9472 29877 9512
rect 29835 9463 29877 9472
rect 30508 9512 30548 9521
rect 30796 9512 30836 9521
rect 30548 9472 30796 9512
rect 30508 9463 30548 9472
rect 30796 9463 30836 9472
rect 29740 8791 29780 8800
rect 29452 8707 29492 8716
rect 29163 8084 29205 8093
rect 29163 8044 29164 8084
rect 29204 8044 29205 8084
rect 29163 8035 29205 8044
rect 29740 8000 29780 8009
rect 29164 7916 29204 7925
rect 29164 7589 29204 7876
rect 29259 7916 29301 7925
rect 29259 7876 29260 7916
rect 29300 7876 29301 7916
rect 29259 7867 29301 7876
rect 29163 7580 29205 7589
rect 29163 7540 29164 7580
rect 29204 7540 29205 7580
rect 29163 7531 29205 7540
rect 28876 6320 28916 7120
rect 28971 7160 29013 7169
rect 28971 7120 28972 7160
rect 29012 7120 29108 7160
rect 28971 7111 29013 7120
rect 28971 6740 29013 6749
rect 28971 6700 28972 6740
rect 29012 6700 29013 6740
rect 28971 6691 29013 6700
rect 28972 6320 29012 6691
rect 28876 6280 29012 6320
rect 28779 5816 28821 5825
rect 28779 5776 28780 5816
rect 28820 5776 28821 5816
rect 28779 5767 28821 5776
rect 28695 5662 28735 5670
rect 28780 5662 28820 5767
rect 28588 5661 28820 5662
rect 28588 5622 28695 5661
rect 28395 4472 28437 4481
rect 28395 4432 28396 4472
rect 28436 4432 28437 4472
rect 28395 4423 28437 4432
rect 28588 4136 28628 5622
rect 28735 5622 28820 5661
rect 28695 5612 28735 5621
rect 29068 5144 29108 7120
rect 29164 7085 29204 7531
rect 29260 7337 29300 7867
rect 29259 7328 29301 7337
rect 29259 7288 29260 7328
rect 29300 7288 29301 7328
rect 29259 7279 29301 7288
rect 29163 7076 29205 7085
rect 29163 7036 29164 7076
rect 29204 7036 29205 7076
rect 29163 7027 29205 7036
rect 29740 6581 29780 7960
rect 29739 6572 29781 6581
rect 29739 6532 29740 6572
rect 29780 6532 29781 6572
rect 29739 6523 29781 6532
rect 29548 6488 29588 6499
rect 29548 6413 29588 6448
rect 29547 6404 29589 6413
rect 29547 6364 29548 6404
rect 29588 6364 29589 6404
rect 29547 6355 29589 6364
rect 29740 6236 29780 6245
rect 29260 6196 29740 6236
rect 29260 5732 29300 6196
rect 29740 6187 29780 6196
rect 29212 5692 29300 5732
rect 29740 5732 29780 5741
rect 29212 5690 29252 5692
rect 29212 5641 29252 5650
rect 29740 5648 29780 5692
rect 29452 5608 29780 5648
rect 29356 5564 29396 5573
rect 29452 5564 29492 5608
rect 29396 5524 29492 5564
rect 29356 5515 29396 5524
rect 29548 5480 29588 5489
rect 29548 5153 29588 5440
rect 28588 3473 28628 4096
rect 28972 5104 29108 5144
rect 29547 5144 29589 5153
rect 29547 5104 29548 5144
rect 29588 5104 29589 5144
rect 28779 3632 28821 3641
rect 28779 3592 28780 3632
rect 28820 3592 28821 3632
rect 28779 3583 28821 3592
rect 28587 3464 28629 3473
rect 28587 3424 28588 3464
rect 28628 3424 28629 3464
rect 28587 3415 28629 3424
rect 28299 3296 28341 3305
rect 28299 3256 28300 3296
rect 28340 3256 28341 3296
rect 28299 3247 28341 3256
rect 28780 2633 28820 3583
rect 28972 2801 29012 5104
rect 29547 5095 29589 5104
rect 29067 4976 29109 4985
rect 29067 4936 29068 4976
rect 29108 4936 29109 4976
rect 29067 4927 29109 4936
rect 29068 4842 29108 4927
rect 29644 4220 29684 4229
rect 29116 4145 29156 4154
rect 29644 4136 29684 4180
rect 29156 4105 29204 4136
rect 29116 4096 29204 4105
rect 29067 3968 29109 3977
rect 29067 3928 29068 3968
rect 29108 3928 29109 3968
rect 29067 3919 29109 3928
rect 28971 2792 29013 2801
rect 28971 2752 28972 2792
rect 29012 2752 29013 2792
rect 28971 2743 29013 2752
rect 28779 2624 28821 2633
rect 28779 2584 28780 2624
rect 28820 2584 28821 2624
rect 28779 2575 28821 2584
rect 28108 2500 28244 2540
rect 27915 2456 27957 2465
rect 27915 2416 27916 2456
rect 27956 2416 27957 2456
rect 27915 2407 27957 2416
rect 27819 2372 27861 2381
rect 27819 2332 27820 2372
rect 27860 2332 27861 2372
rect 27819 2323 27861 2332
rect 27723 1952 27765 1961
rect 27723 1912 27724 1952
rect 27764 1912 27765 1952
rect 27723 1903 27765 1912
rect 27820 1952 27860 2323
rect 27820 1903 27860 1912
rect 27436 1828 27572 1868
rect 27243 1819 27285 1828
rect 27244 1734 27284 1819
rect 27436 1700 27476 1709
rect 27339 1196 27381 1205
rect 27339 1156 27340 1196
rect 27380 1156 27381 1196
rect 27339 1147 27381 1156
rect 27340 80 27380 1147
rect 27436 953 27476 1660
rect 27435 944 27477 953
rect 27435 904 27436 944
rect 27476 904 27477 944
rect 27435 895 27477 904
rect 27532 80 27572 1828
rect 27724 1818 27764 1903
rect 27916 1280 27956 2407
rect 28011 2372 28053 2381
rect 28011 2332 28012 2372
rect 28052 2332 28053 2372
rect 28011 2323 28053 2332
rect 28012 1541 28052 2323
rect 28108 2045 28148 2500
rect 28587 2456 28629 2465
rect 28587 2416 28588 2456
rect 28628 2416 28629 2456
rect 28587 2407 28629 2416
rect 28972 2456 29012 2465
rect 28395 2120 28437 2129
rect 28395 2080 28396 2120
rect 28436 2080 28437 2120
rect 28395 2071 28437 2080
rect 28107 2036 28149 2045
rect 28107 1996 28108 2036
rect 28148 1996 28149 2036
rect 28107 1987 28149 1996
rect 28204 1868 28244 1877
rect 28011 1532 28053 1541
rect 28011 1492 28012 1532
rect 28052 1492 28053 1532
rect 28011 1483 28053 1492
rect 28204 1373 28244 1828
rect 28300 1868 28340 1879
rect 28300 1793 28340 1828
rect 28299 1784 28341 1793
rect 28299 1744 28300 1784
rect 28340 1744 28341 1784
rect 28299 1735 28341 1744
rect 28396 1541 28436 2071
rect 28395 1532 28437 1541
rect 28395 1492 28396 1532
rect 28436 1492 28437 1532
rect 28395 1483 28437 1492
rect 28203 1364 28245 1373
rect 28203 1324 28204 1364
rect 28244 1324 28245 1364
rect 28203 1315 28245 1324
rect 27724 1240 27956 1280
rect 27724 80 27764 1240
rect 28492 1196 28532 1205
rect 28492 1037 28532 1156
rect 28491 1028 28533 1037
rect 28491 988 28492 1028
rect 28532 988 28533 1028
rect 28491 979 28533 988
rect 27915 944 27957 953
rect 27915 904 27916 944
rect 27956 904 27957 944
rect 27915 895 27957 904
rect 27916 80 27956 895
rect 28588 860 28628 2407
rect 28779 2372 28821 2381
rect 28779 2332 28780 2372
rect 28820 2332 28821 2372
rect 28779 2323 28821 2332
rect 28780 1952 28820 2323
rect 28875 2204 28917 2213
rect 28875 2164 28876 2204
rect 28916 2164 28917 2204
rect 28875 2155 28917 2164
rect 28780 1903 28820 1912
rect 28683 944 28725 953
rect 28683 904 28684 944
rect 28724 904 28725 944
rect 28683 895 28725 904
rect 28492 820 28628 860
rect 28107 440 28149 449
rect 28107 400 28108 440
rect 28148 400 28149 440
rect 28107 391 28149 400
rect 28108 80 28148 391
rect 28299 104 28341 113
rect 28299 80 28300 104
rect 9524 64 9544 80
rect 9464 0 9544 64
rect 9656 0 9736 80
rect 9848 0 9928 80
rect 10040 0 10120 80
rect 10232 0 10312 80
rect 10424 0 10504 80
rect 10616 0 10696 80
rect 10808 0 10888 80
rect 11000 0 11080 80
rect 11192 0 11272 80
rect 11384 0 11464 80
rect 11576 0 11656 80
rect 11768 0 11848 80
rect 11960 0 12040 80
rect 12152 0 12232 80
rect 12344 0 12424 80
rect 12536 0 12616 80
rect 12728 0 12808 80
rect 12920 0 13000 80
rect 13112 0 13192 80
rect 13304 0 13384 80
rect 13496 0 13576 80
rect 13688 0 13768 80
rect 13880 0 13960 80
rect 14072 0 14152 80
rect 14264 0 14344 80
rect 14456 0 14536 80
rect 14648 0 14728 80
rect 14840 0 14920 80
rect 15032 0 15112 80
rect 15224 0 15304 80
rect 15416 0 15496 80
rect 15608 0 15688 80
rect 15800 0 15880 80
rect 15992 0 16072 80
rect 16184 0 16264 80
rect 16376 0 16456 80
rect 16568 0 16648 80
rect 16760 0 16840 80
rect 16952 0 17032 80
rect 17144 0 17224 80
rect 17336 0 17416 80
rect 17528 0 17608 80
rect 17720 0 17800 80
rect 17912 0 17992 80
rect 18104 0 18184 80
rect 18296 0 18376 80
rect 18488 0 18568 80
rect 18680 0 18760 80
rect 18872 0 18952 80
rect 19064 0 19144 80
rect 19256 0 19336 80
rect 19448 0 19528 80
rect 19640 0 19720 80
rect 19832 0 19912 80
rect 20024 0 20104 80
rect 20216 0 20296 80
rect 20408 0 20488 80
rect 20600 0 20680 80
rect 20792 0 20872 80
rect 20984 0 21064 80
rect 21176 0 21256 80
rect 21368 0 21448 80
rect 21560 0 21640 80
rect 21752 0 21832 80
rect 21944 0 22024 80
rect 22136 0 22216 80
rect 22328 0 22408 80
rect 22520 0 22600 80
rect 22712 0 22792 80
rect 22904 0 22984 80
rect 23096 0 23176 80
rect 23288 0 23368 80
rect 23480 0 23560 80
rect 23672 0 23752 80
rect 23864 0 23944 80
rect 24056 0 24136 80
rect 24248 0 24328 80
rect 24440 0 24520 80
rect 24632 0 24712 80
rect 24824 0 24904 80
rect 25016 0 25096 80
rect 25208 0 25288 80
rect 25400 0 25480 80
rect 25592 0 25672 80
rect 25784 0 25864 80
rect 25976 0 26056 80
rect 26168 0 26248 80
rect 26360 0 26440 80
rect 26552 0 26632 80
rect 26744 0 26824 80
rect 26936 0 27016 80
rect 27128 0 27208 80
rect 27320 0 27400 80
rect 27512 0 27592 80
rect 27704 0 27784 80
rect 27896 0 27976 80
rect 28088 0 28168 80
rect 28280 64 28300 80
rect 28340 80 28341 104
rect 28492 80 28532 820
rect 28684 810 28724 895
rect 28683 356 28725 365
rect 28683 316 28684 356
rect 28724 316 28725 356
rect 28683 307 28725 316
rect 28684 80 28724 307
rect 28876 80 28916 2155
rect 28972 1961 29012 2416
rect 28971 1952 29013 1961
rect 28971 1912 28972 1952
rect 29012 1912 29013 1952
rect 28971 1903 29013 1912
rect 29068 80 29108 3919
rect 29164 3632 29204 4096
rect 29356 4096 29684 4136
rect 29260 4052 29300 4061
rect 29356 4052 29396 4096
rect 29300 4012 29396 4052
rect 29260 4003 29300 4012
rect 29452 3968 29492 3977
rect 29492 3928 29684 3968
rect 29452 3919 29492 3928
rect 29548 3632 29588 3641
rect 29164 3592 29548 3632
rect 29548 3583 29588 3592
rect 29356 3464 29396 3473
rect 29356 3389 29396 3424
rect 29355 3380 29397 3389
rect 29355 3340 29356 3380
rect 29396 3340 29397 3380
rect 29355 3331 29397 3340
rect 29356 3053 29396 3331
rect 29355 3044 29397 3053
rect 29355 3004 29356 3044
rect 29396 3004 29397 3044
rect 29355 2995 29397 3004
rect 29163 2792 29205 2801
rect 29163 2752 29164 2792
rect 29204 2752 29205 2792
rect 29163 2743 29205 2752
rect 29164 2624 29204 2743
rect 29164 2575 29204 2584
rect 29259 1952 29301 1961
rect 29259 1907 29260 1952
rect 29300 1907 29301 1952
rect 29259 1903 29301 1907
rect 29260 1817 29300 1903
rect 29163 1112 29205 1121
rect 29163 1072 29164 1112
rect 29204 1072 29205 1112
rect 29163 1063 29205 1072
rect 29164 978 29204 1063
rect 29356 1037 29396 2995
rect 29644 2633 29684 3928
rect 29643 2624 29685 2633
rect 29643 2584 29644 2624
rect 29684 2584 29685 2624
rect 29643 2575 29685 2584
rect 29836 2540 29876 9463
rect 30603 9092 30645 9101
rect 30603 9052 30604 9092
rect 30644 9052 30645 9092
rect 30603 9043 30645 9052
rect 29740 2500 29876 2540
rect 29932 8756 29972 8765
rect 29452 2036 29492 2045
rect 29452 1877 29492 1996
rect 29451 1868 29493 1877
rect 29451 1828 29452 1868
rect 29492 1828 29493 1868
rect 29451 1819 29493 1828
rect 29644 1700 29684 1709
rect 29452 1660 29644 1700
rect 29355 1028 29397 1037
rect 29355 988 29356 1028
rect 29396 988 29397 1028
rect 29355 979 29397 988
rect 29259 944 29301 953
rect 29259 904 29260 944
rect 29300 904 29301 944
rect 29259 895 29301 904
rect 29260 80 29300 895
rect 29452 80 29492 1660
rect 29644 1651 29684 1660
rect 29740 1532 29780 2500
rect 29932 2297 29972 8716
rect 30027 8672 30069 8681
rect 30124 8672 30164 8681
rect 30027 8632 30028 8672
rect 30068 8632 30124 8672
rect 30027 8623 30069 8632
rect 30124 8623 30164 8632
rect 30028 6908 30068 8623
rect 30412 8084 30452 8093
rect 30452 8044 30548 8084
rect 30412 8035 30452 8044
rect 30268 7958 30308 7967
rect 30268 7916 30308 7918
rect 30268 7876 30356 7916
rect 30316 7412 30356 7876
rect 30316 7363 30356 7372
rect 30508 7244 30548 8044
rect 30604 7832 30644 9043
rect 30892 8849 30932 9640
rect 32044 9631 32084 9640
rect 32428 9680 32468 10051
rect 32428 9631 32468 9640
rect 31659 9512 31701 9521
rect 31659 9472 31660 9512
rect 31700 9472 31701 9512
rect 31659 9463 31701 9472
rect 31660 9378 31700 9463
rect 32235 9428 32277 9437
rect 32235 9388 32236 9428
rect 32276 9388 32277 9428
rect 32235 9379 32277 9388
rect 32236 9294 32276 9379
rect 31755 8924 31797 8933
rect 31755 8884 31756 8924
rect 31796 8884 31797 8924
rect 31755 8875 31797 8884
rect 30891 8840 30933 8849
rect 30891 8800 30892 8840
rect 30932 8800 30933 8840
rect 30891 8791 30933 8800
rect 31756 8840 31796 8875
rect 31756 8789 31796 8800
rect 32139 8840 32181 8849
rect 32139 8800 32140 8840
rect 32180 8800 32181 8840
rect 32139 8791 32181 8800
rect 32524 8840 32564 10692
rect 32888 10672 32968 10752
rect 34040 10672 34120 10752
rect 35192 10672 35272 10752
rect 36344 10672 36424 10752
rect 37496 10672 37576 10752
rect 38648 10672 38728 10752
rect 39800 10672 39880 10752
rect 40396 10692 40906 10732
rect 32811 9932 32853 9941
rect 32811 9892 32812 9932
rect 32852 9892 32853 9932
rect 32811 9883 32853 9892
rect 32812 9680 32852 9883
rect 32812 9631 32852 9640
rect 32620 9428 32660 9437
rect 32620 9017 32660 9388
rect 32619 9008 32661 9017
rect 32619 8968 32620 9008
rect 32660 8968 32661 9008
rect 32619 8959 32661 8968
rect 32524 8791 32564 8800
rect 32908 8840 32948 10672
rect 34060 9512 34100 10672
rect 35212 10016 35252 10672
rect 35020 9976 35252 10016
rect 34539 9512 34581 9521
rect 34060 9472 34388 9512
rect 32908 8791 32948 8800
rect 33004 9428 33044 9437
rect 31948 8756 31988 8765
rect 31372 8672 31412 8681
rect 31083 8504 31125 8513
rect 31083 8464 31084 8504
rect 31124 8464 31125 8504
rect 31083 8455 31125 8464
rect 31084 8000 31124 8455
rect 31084 7951 31124 7960
rect 31180 8000 31220 8009
rect 30604 7783 30644 7792
rect 30796 7916 30836 7925
rect 30700 7244 30740 7253
rect 30508 7204 30700 7244
rect 30700 7195 30740 7204
rect 30123 7160 30165 7169
rect 30123 7120 30124 7160
rect 30164 7120 30165 7160
rect 30123 7111 30165 7120
rect 30124 7026 30164 7111
rect 30508 6992 30548 7001
rect 30412 6952 30508 6992
rect 30028 6868 30164 6908
rect 30027 6740 30069 6749
rect 30027 6700 30028 6740
rect 30068 6700 30069 6740
rect 30027 6691 30069 6700
rect 30028 3464 30068 6691
rect 30124 6161 30164 6868
rect 30219 6572 30261 6581
rect 30219 6532 30220 6572
rect 30260 6532 30261 6572
rect 30219 6523 30261 6532
rect 30123 6152 30165 6161
rect 30123 6112 30124 6152
rect 30164 6112 30165 6152
rect 30123 6103 30165 6112
rect 30124 5648 30164 5657
rect 30124 5489 30164 5608
rect 30123 5480 30165 5489
rect 30123 5440 30124 5480
rect 30164 5440 30165 5480
rect 30123 5431 30165 5440
rect 30123 5312 30165 5321
rect 30123 5272 30124 5312
rect 30164 5272 30165 5312
rect 30123 5263 30165 5272
rect 30028 3305 30068 3424
rect 30027 3296 30069 3305
rect 30027 3256 30028 3296
rect 30068 3256 30069 3296
rect 30027 3247 30069 3256
rect 30124 3128 30164 5263
rect 30028 3088 30164 3128
rect 29931 2288 29973 2297
rect 29931 2248 29932 2288
rect 29972 2248 29973 2288
rect 29931 2239 29973 2248
rect 29835 2036 29877 2045
rect 29835 1996 29836 2036
rect 29876 1996 29877 2036
rect 29835 1987 29877 1996
rect 29836 1881 29876 1987
rect 30028 1868 30068 3088
rect 30220 2960 30260 6523
rect 30316 4976 30356 4985
rect 30316 4565 30356 4936
rect 30315 4556 30357 4565
rect 30315 4516 30316 4556
rect 30356 4516 30357 4556
rect 30315 4507 30357 4516
rect 30124 2920 30260 2960
rect 30124 2633 30164 2920
rect 30219 2792 30261 2801
rect 30219 2752 30220 2792
rect 30260 2752 30261 2792
rect 30219 2743 30261 2752
rect 30123 2624 30165 2633
rect 30123 2584 30124 2624
rect 30164 2584 30165 2624
rect 30123 2575 30165 2584
rect 30220 2036 30260 2743
rect 29836 1832 29876 1841
rect 29932 1828 30068 1868
rect 30124 1996 30260 2036
rect 29932 1784 29972 1828
rect 29644 1492 29780 1532
rect 29836 1744 29972 1784
rect 29644 80 29684 1492
rect 29836 80 29876 1744
rect 30028 1700 30068 1709
rect 30028 1541 30068 1660
rect 30124 1616 30164 1996
rect 30219 1868 30261 1877
rect 30219 1828 30220 1868
rect 30260 1828 30261 1868
rect 30219 1819 30261 1828
rect 30220 1734 30260 1819
rect 30124 1576 30260 1616
rect 30027 1532 30069 1541
rect 30027 1492 30028 1532
rect 30068 1492 30069 1532
rect 30027 1483 30069 1492
rect 30027 1028 30069 1037
rect 30027 988 30028 1028
rect 30068 988 30069 1028
rect 30027 979 30069 988
rect 30028 80 30068 979
rect 30220 80 30260 1576
rect 30316 944 30356 4507
rect 30412 3893 30452 6952
rect 30508 6943 30548 6952
rect 30507 6572 30549 6581
rect 30507 6532 30508 6572
rect 30548 6532 30549 6572
rect 30507 6523 30549 6532
rect 30508 6488 30548 6523
rect 30508 6437 30548 6448
rect 30508 4724 30548 4733
rect 30548 4684 30644 4724
rect 30508 4675 30548 4684
rect 30604 4136 30644 4684
rect 30604 4087 30644 4096
rect 30796 3968 30836 7876
rect 31180 4892 31220 7960
rect 31372 7169 31412 8632
rect 31563 8504 31605 8513
rect 31563 8464 31564 8504
rect 31604 8464 31605 8504
rect 31563 8455 31605 8464
rect 31564 8370 31604 8455
rect 31755 8084 31797 8093
rect 31755 8044 31756 8084
rect 31796 8044 31797 8084
rect 31755 8035 31797 8044
rect 31563 7916 31605 7925
rect 31563 7876 31564 7916
rect 31604 7876 31605 7916
rect 31563 7867 31605 7876
rect 31660 7916 31700 7925
rect 31564 7782 31604 7867
rect 31660 7589 31700 7876
rect 31659 7580 31701 7589
rect 31659 7540 31660 7580
rect 31700 7540 31701 7580
rect 31659 7531 31701 7540
rect 31371 7160 31413 7169
rect 31371 7120 31372 7160
rect 31412 7120 31413 7160
rect 31371 7111 31413 7120
rect 31660 7160 31700 7171
rect 31275 6404 31317 6413
rect 31372 6404 31412 7111
rect 31660 7085 31700 7120
rect 31659 7076 31701 7085
rect 31659 7036 31660 7076
rect 31700 7036 31701 7076
rect 31659 7027 31701 7036
rect 31756 6824 31796 8035
rect 31660 6784 31796 6824
rect 31467 6488 31509 6497
rect 31467 6448 31468 6488
rect 31508 6448 31509 6488
rect 31467 6439 31509 6448
rect 31275 6364 31276 6404
rect 31316 6364 31412 6404
rect 31275 6355 31317 6364
rect 31372 5648 31412 6364
rect 31372 5599 31412 5608
rect 31468 5480 31508 6439
rect 31563 5564 31605 5573
rect 31563 5524 31564 5564
rect 31604 5524 31605 5564
rect 31563 5515 31605 5524
rect 30508 3928 30836 3968
rect 30892 4852 31220 4892
rect 31372 5440 31508 5480
rect 30892 4136 30932 4852
rect 31276 4304 31316 4313
rect 30411 3884 30453 3893
rect 30411 3844 30412 3884
rect 30452 3844 30453 3884
rect 30411 3835 30453 3844
rect 30411 3128 30453 3137
rect 30411 3088 30412 3128
rect 30452 3088 30453 3128
rect 30411 3079 30453 3088
rect 30412 2624 30452 3079
rect 30412 2575 30452 2584
rect 30411 2288 30453 2297
rect 30411 2248 30412 2288
rect 30452 2248 30453 2288
rect 30411 2239 30453 2248
rect 30412 1280 30452 2239
rect 30508 2036 30548 3928
rect 30795 3716 30837 3725
rect 30795 3676 30796 3716
rect 30836 3676 30837 3716
rect 30795 3667 30837 3676
rect 30796 3053 30836 3667
rect 30795 3044 30837 3053
rect 30795 3004 30796 3044
rect 30836 3004 30837 3044
rect 30795 2995 30837 3004
rect 30796 2624 30836 2995
rect 30796 2575 30836 2584
rect 30892 2549 30932 4096
rect 31180 4264 31276 4304
rect 30988 4052 31028 4061
rect 30988 3893 31028 4012
rect 30987 3884 31029 3893
rect 30987 3844 30988 3884
rect 31028 3844 31029 3884
rect 30987 3835 31029 3844
rect 30891 2540 30933 2549
rect 30891 2500 30892 2540
rect 30932 2500 30933 2540
rect 30891 2491 30933 2500
rect 31083 2540 31125 2549
rect 31083 2500 31084 2540
rect 31124 2500 31125 2540
rect 31083 2491 31125 2500
rect 30604 2456 30644 2465
rect 30604 2120 30644 2416
rect 30604 2080 30932 2120
rect 30508 1996 30740 2036
rect 30508 1933 30548 1942
rect 30508 1364 30548 1893
rect 30604 1933 30644 1942
rect 30604 1877 30644 1893
rect 30603 1868 30645 1877
rect 30603 1828 30604 1868
rect 30644 1828 30645 1868
rect 30603 1819 30645 1828
rect 30604 1798 30644 1819
rect 30604 1364 30644 1373
rect 30508 1324 30604 1364
rect 30604 1315 30644 1324
rect 30412 1240 30548 1280
rect 30508 1196 30548 1240
rect 30508 1156 30644 1196
rect 30412 1112 30452 1121
rect 30412 1028 30452 1072
rect 30507 1028 30549 1037
rect 30412 988 30508 1028
rect 30548 988 30549 1028
rect 30507 979 30549 988
rect 30316 904 30452 944
rect 30412 80 30452 904
rect 30604 80 30644 1156
rect 30700 869 30740 1996
rect 30892 1028 30932 2080
rect 31084 1952 31124 2491
rect 31084 1903 31124 1912
rect 30987 1868 31029 1877
rect 30987 1828 30988 1868
rect 31028 1828 31029 1868
rect 30987 1819 31029 1828
rect 30988 1734 31028 1819
rect 30988 1196 31028 1205
rect 31180 1196 31220 4264
rect 31276 4255 31316 4264
rect 31275 3716 31317 3725
rect 31275 3676 31276 3716
rect 31316 3676 31317 3716
rect 31275 3667 31317 3676
rect 31276 3464 31316 3667
rect 31276 3415 31316 3424
rect 31275 2120 31317 2129
rect 31275 2080 31276 2120
rect 31316 2080 31317 2120
rect 31275 2071 31317 2080
rect 31276 1364 31316 2071
rect 31372 1868 31412 5440
rect 31564 5430 31604 5515
rect 31563 3884 31605 3893
rect 31563 3844 31564 3884
rect 31604 3844 31605 3884
rect 31563 3835 31605 3844
rect 31467 3548 31509 3557
rect 31467 3508 31468 3548
rect 31508 3508 31509 3548
rect 31467 3499 31509 3508
rect 31468 3414 31508 3499
rect 31564 1961 31604 3835
rect 31563 1952 31605 1961
rect 31563 1912 31564 1952
rect 31604 1912 31605 1952
rect 31563 1903 31605 1912
rect 31372 1828 31508 1868
rect 31371 1364 31413 1373
rect 31276 1324 31372 1364
rect 31412 1324 31413 1364
rect 31371 1315 31413 1324
rect 31028 1156 31220 1196
rect 30988 1147 31028 1156
rect 31276 1112 31316 1121
rect 31276 1028 31316 1072
rect 31372 1112 31412 1315
rect 31372 1063 31412 1072
rect 30892 988 31316 1028
rect 30796 944 30836 953
rect 31468 944 31508 1828
rect 31660 1784 31700 6784
rect 31756 6446 31796 6499
rect 31948 6497 31988 8716
rect 32140 8706 32180 8791
rect 32332 8756 32372 8765
rect 32236 8716 32332 8756
rect 32140 8000 32180 8011
rect 32140 7925 32180 7960
rect 32139 7916 32181 7925
rect 32139 7876 32140 7916
rect 32180 7876 32181 7916
rect 32139 7867 32181 7876
rect 31755 6406 31756 6413
rect 31947 6488 31989 6497
rect 31947 6448 31948 6488
rect 31988 6448 31989 6488
rect 31947 6439 31989 6448
rect 31796 6406 31797 6413
rect 31755 6404 31797 6406
rect 31755 6364 31756 6404
rect 31796 6364 31797 6404
rect 31755 6355 31797 6364
rect 31755 6236 31797 6245
rect 31755 6196 31756 6236
rect 31796 6196 31797 6236
rect 31755 6187 31797 6196
rect 31948 6236 31988 6245
rect 32139 6236 32181 6245
rect 31988 6196 32084 6236
rect 31948 6187 31988 6196
rect 31756 3809 31796 6187
rect 31852 5648 31892 5659
rect 31948 5657 31988 5742
rect 31852 5573 31892 5608
rect 31947 5648 31989 5657
rect 31947 5608 31948 5648
rect 31988 5608 31989 5648
rect 31947 5599 31989 5608
rect 31851 5564 31893 5573
rect 31851 5524 31852 5564
rect 31892 5524 31893 5564
rect 31851 5515 31893 5524
rect 32044 5480 32084 6196
rect 32139 6196 32140 6236
rect 32180 6196 32181 6236
rect 32139 6187 32181 6196
rect 32140 6102 32180 6187
rect 32139 5648 32181 5657
rect 32139 5608 32140 5648
rect 32180 5608 32181 5648
rect 32139 5599 32181 5608
rect 31948 5440 32084 5480
rect 31948 4976 31988 5440
rect 31948 4927 31988 4936
rect 32044 4976 32084 4985
rect 32140 4976 32180 5599
rect 32084 4936 32180 4976
rect 32044 4927 32084 4936
rect 31947 4808 31989 4817
rect 31947 4768 31948 4808
rect 31988 4768 31989 4808
rect 31947 4759 31989 4768
rect 31755 3800 31797 3809
rect 31755 3760 31756 3800
rect 31796 3760 31797 3800
rect 31755 3751 31797 3760
rect 31755 3548 31797 3557
rect 31755 3508 31756 3548
rect 31796 3508 31797 3548
rect 31755 3499 31797 3508
rect 31756 3464 31796 3499
rect 31756 3413 31796 3424
rect 31851 3464 31893 3473
rect 31851 3424 31852 3464
rect 31892 3424 31893 3464
rect 31851 3415 31893 3424
rect 31852 3330 31892 3415
rect 31851 2624 31893 2633
rect 31851 2584 31852 2624
rect 31892 2584 31893 2624
rect 31851 2575 31893 2584
rect 30836 904 30932 944
rect 30796 895 30836 904
rect 30699 860 30741 869
rect 30699 820 30700 860
rect 30740 820 30741 860
rect 30699 811 30741 820
rect 30795 776 30837 785
rect 30795 736 30796 776
rect 30836 736 30837 776
rect 30795 727 30837 736
rect 30796 80 30836 727
rect 30892 197 30932 904
rect 31372 904 31508 944
rect 31564 1744 31700 1784
rect 31755 1784 31797 1793
rect 31755 1744 31756 1784
rect 31796 1744 31797 1784
rect 30987 860 31029 869
rect 30987 820 30988 860
rect 31028 820 31029 860
rect 30987 811 31029 820
rect 30891 188 30933 197
rect 30891 148 30892 188
rect 30932 148 30933 188
rect 30891 139 30933 148
rect 30988 80 31028 811
rect 31179 776 31221 785
rect 31179 736 31180 776
rect 31220 736 31221 776
rect 31179 727 31221 736
rect 31180 80 31220 727
rect 31372 80 31412 904
rect 31564 80 31604 1744
rect 31755 1735 31797 1744
rect 31659 1280 31701 1289
rect 31659 1240 31660 1280
rect 31700 1240 31701 1280
rect 31659 1231 31701 1240
rect 31660 869 31700 1231
rect 31756 1196 31796 1735
rect 31756 1147 31796 1156
rect 31852 1196 31892 2575
rect 31852 1147 31892 1156
rect 31948 1028 31988 4759
rect 32043 3800 32085 3809
rect 32043 3760 32044 3800
rect 32084 3760 32085 3800
rect 32043 3751 32085 3760
rect 32044 3641 32084 3751
rect 32043 3632 32085 3641
rect 32043 3592 32044 3632
rect 32084 3592 32085 3632
rect 32043 3583 32085 3592
rect 32044 2624 32084 3583
rect 32044 2575 32084 2584
rect 32140 2456 32180 4936
rect 32236 4817 32276 8716
rect 32332 8707 32372 8716
rect 32716 8756 32756 8765
rect 32620 7986 32660 7995
rect 32523 7916 32565 7925
rect 32523 7876 32524 7916
rect 32564 7876 32565 7916
rect 32523 7867 32565 7876
rect 32524 7757 32564 7867
rect 32523 7748 32565 7757
rect 32523 7708 32524 7748
rect 32564 7708 32565 7748
rect 32523 7699 32565 7708
rect 32427 7580 32469 7589
rect 32427 7540 32428 7580
rect 32468 7540 32469 7580
rect 32427 7531 32469 7540
rect 32331 6404 32373 6413
rect 32331 6364 32332 6404
rect 32372 6364 32373 6404
rect 32331 6355 32373 6364
rect 32332 6270 32372 6355
rect 32332 5648 32372 5657
rect 32332 4892 32372 5608
rect 32428 5648 32468 7531
rect 32524 7412 32564 7699
rect 32620 7589 32660 7946
rect 32619 7580 32661 7589
rect 32619 7540 32620 7580
rect 32660 7540 32661 7580
rect 32619 7531 32661 7540
rect 32524 7372 32660 7412
rect 32523 6740 32565 6749
rect 32523 6700 32524 6740
rect 32564 6700 32565 6740
rect 32523 6691 32565 6700
rect 32428 5060 32468 5608
rect 32524 6488 32564 6691
rect 32524 5237 32564 6448
rect 32523 5228 32565 5237
rect 32523 5188 32524 5228
rect 32564 5188 32565 5228
rect 32523 5179 32565 5188
rect 32428 5020 32564 5060
rect 32427 4892 32469 4901
rect 32332 4852 32428 4892
rect 32468 4852 32469 4892
rect 32427 4843 32469 4852
rect 32524 4892 32564 5020
rect 32235 4808 32277 4817
rect 32235 4768 32236 4808
rect 32276 4768 32277 4808
rect 32235 4759 32277 4768
rect 32428 4758 32468 4843
rect 32524 4817 32564 4852
rect 32523 4808 32565 4817
rect 32523 4768 32524 4808
rect 32564 4768 32565 4808
rect 32523 4759 32565 4768
rect 32620 4640 32660 7372
rect 32428 4600 32660 4640
rect 32428 3893 32468 4600
rect 32620 3968 32660 3977
rect 32524 3928 32620 3968
rect 32427 3884 32469 3893
rect 32427 3844 32428 3884
rect 32468 3844 32469 3884
rect 32427 3835 32469 3844
rect 32236 3380 32276 3389
rect 32236 2633 32276 3340
rect 32332 3380 32372 3389
rect 32235 2624 32277 2633
rect 32235 2584 32236 2624
rect 32276 2584 32277 2624
rect 32235 2575 32277 2584
rect 32044 2416 32180 2456
rect 32044 2129 32084 2416
rect 32332 2381 32372 3340
rect 32427 3212 32469 3221
rect 32427 3172 32428 3212
rect 32468 3172 32469 3212
rect 32427 3163 32469 3172
rect 32428 2456 32468 3163
rect 32524 2633 32564 3928
rect 32620 3919 32660 3928
rect 32716 3800 32756 8716
rect 33004 8093 33044 9388
rect 33388 9344 33428 9353
rect 33428 9304 33716 9344
rect 33388 9295 33428 9304
rect 33100 8756 33140 8765
rect 33140 8716 33236 8756
rect 33100 8707 33140 8716
rect 32812 8084 32852 8093
rect 32812 6413 32852 8044
rect 33003 8084 33045 8093
rect 33003 8044 33004 8084
rect 33044 8044 33045 8084
rect 33003 8035 33045 8044
rect 33099 7916 33141 7925
rect 33099 7876 33100 7916
rect 33140 7876 33141 7916
rect 33099 7867 33141 7876
rect 33100 7782 33140 7867
rect 33099 7580 33141 7589
rect 33099 7540 33100 7580
rect 33140 7540 33141 7580
rect 33099 7531 33141 7540
rect 33100 7412 33140 7531
rect 33100 7363 33140 7372
rect 32907 7160 32949 7169
rect 32907 7120 32908 7160
rect 32948 7120 32949 7160
rect 32907 7111 32949 7120
rect 32908 7026 32948 7111
rect 32811 6404 32853 6413
rect 32811 6364 32812 6404
rect 32852 6364 32853 6404
rect 32811 6355 32853 6364
rect 32907 5732 32949 5741
rect 32907 5692 32908 5732
rect 32948 5692 32949 5732
rect 32907 5683 32949 5692
rect 33099 5732 33141 5741
rect 33099 5692 33100 5732
rect 33140 5692 33141 5732
rect 33099 5683 33141 5692
rect 32908 5648 32948 5683
rect 32908 5597 32948 5608
rect 33004 4976 33044 4985
rect 33100 4976 33140 5683
rect 33196 5657 33236 8716
rect 33676 8672 33716 9304
rect 34252 9269 34292 9354
rect 34251 9260 34293 9269
rect 34251 9220 34252 9260
rect 34292 9220 34293 9260
rect 34251 9211 34293 9220
rect 33928 9092 34296 9101
rect 33968 9052 34010 9092
rect 34050 9052 34092 9092
rect 34132 9052 34174 9092
rect 34214 9052 34256 9092
rect 33928 9043 34296 9052
rect 33964 8672 34004 8681
rect 33676 8632 33964 8672
rect 33964 8623 34004 8632
rect 33580 8588 33620 8597
rect 33291 8168 33333 8177
rect 33291 8128 33292 8168
rect 33332 8128 33333 8168
rect 33291 8119 33333 8128
rect 33292 8034 33332 8119
rect 33580 8009 33620 8548
rect 34348 8177 34388 9472
rect 34539 9472 34540 9512
rect 34580 9472 34581 9512
rect 34539 9463 34581 9472
rect 34540 9378 34580 9463
rect 34828 9344 34868 9353
rect 34732 9304 34828 9344
rect 34347 8168 34389 8177
rect 34347 8128 34348 8168
rect 34388 8128 34389 8168
rect 34347 8119 34389 8128
rect 33675 8084 33717 8093
rect 33675 8044 33676 8084
rect 33716 8044 33717 8084
rect 33675 8035 33717 8044
rect 33579 8000 33621 8009
rect 33579 7960 33580 8000
rect 33620 7960 33621 8000
rect 33579 7951 33621 7960
rect 33291 7916 33333 7925
rect 33291 7876 33292 7916
rect 33332 7876 33333 7916
rect 33291 7867 33333 7876
rect 33292 5741 33332 7867
rect 33387 7832 33429 7841
rect 33387 7792 33388 7832
rect 33428 7792 33429 7832
rect 33387 7783 33429 7792
rect 33388 7160 33428 7783
rect 33388 7111 33428 7120
rect 33387 6236 33429 6245
rect 33387 6196 33388 6236
rect 33428 6196 33429 6236
rect 33387 6187 33429 6196
rect 33291 5732 33333 5741
rect 33291 5692 33292 5732
rect 33332 5692 33333 5732
rect 33291 5683 33333 5692
rect 33388 5662 33428 6187
rect 33195 5648 33237 5657
rect 33195 5608 33196 5648
rect 33236 5608 33237 5648
rect 33388 5613 33428 5622
rect 33195 5599 33237 5608
rect 33580 5480 33620 5489
rect 33044 4936 33140 4976
rect 33196 5440 33580 5480
rect 33004 4927 33044 4936
rect 32811 4220 32853 4229
rect 32811 4180 32812 4220
rect 32852 4180 32853 4220
rect 32811 4171 32853 4180
rect 33196 4220 33236 5440
rect 33580 5431 33620 5440
rect 33676 5321 33716 8035
rect 34060 8000 34100 8009
rect 34060 7748 34100 7960
rect 34444 8000 34484 8009
rect 34732 8000 34772 9304
rect 34828 9295 34868 9304
rect 34827 9176 34869 9185
rect 34827 9136 34828 9176
rect 34868 9136 34869 9176
rect 34827 9127 34869 9136
rect 34828 8672 34868 9127
rect 35020 8849 35060 9976
rect 35168 9848 35536 9857
rect 35208 9808 35250 9848
rect 35290 9808 35332 9848
rect 35372 9808 35414 9848
rect 35454 9808 35496 9848
rect 35168 9799 35536 9808
rect 35211 9512 35253 9521
rect 35211 9472 35212 9512
rect 35252 9472 35253 9512
rect 35211 9463 35253 9472
rect 36171 9512 36213 9521
rect 36171 9472 36172 9512
rect 36212 9472 36213 9512
rect 36171 9463 36213 9472
rect 35212 9378 35252 9463
rect 36172 9378 36212 9463
rect 35884 9260 35924 9269
rect 35884 9101 35924 9220
rect 35883 9092 35925 9101
rect 35883 9052 35884 9092
rect 35924 9052 35925 9092
rect 35883 9043 35925 9052
rect 36364 8924 36404 10672
rect 37516 10016 37556 10672
rect 37516 9976 37748 10016
rect 37708 9680 37748 9976
rect 37708 9631 37748 9640
rect 36555 9596 36597 9605
rect 36555 9556 36556 9596
rect 36596 9556 36597 9596
rect 36555 9547 36597 9556
rect 36556 9512 36596 9547
rect 36556 9461 36596 9472
rect 36843 9512 36885 9521
rect 36843 9472 36844 9512
rect 36884 9472 36885 9512
rect 36843 9463 36885 9472
rect 36844 9344 36884 9463
rect 37900 9428 37940 9437
rect 36844 9295 36884 9304
rect 37804 9388 37900 9428
rect 36843 9092 36885 9101
rect 36843 9052 36844 9092
rect 36884 9052 36885 9092
rect 36843 9043 36885 9052
rect 36364 8884 36500 8924
rect 35019 8840 35061 8849
rect 35019 8800 35020 8840
rect 35060 8800 35061 8840
rect 35019 8791 35061 8800
rect 36171 8840 36213 8849
rect 36171 8800 36172 8840
rect 36212 8800 36213 8840
rect 36460 8840 36500 8884
rect 36556 8840 36596 8849
rect 36460 8800 36556 8840
rect 36171 8791 36213 8800
rect 36556 8791 36596 8800
rect 36172 8706 36212 8791
rect 36364 8756 36404 8765
rect 36268 8716 36364 8756
rect 34828 8623 34868 8632
rect 35980 8504 36020 8513
rect 35168 8336 35536 8345
rect 35208 8296 35250 8336
rect 35290 8296 35332 8336
rect 35372 8296 35414 8336
rect 35454 8296 35496 8336
rect 35168 8287 35536 8296
rect 34484 7960 34772 8000
rect 35307 8000 35349 8009
rect 35307 7960 35308 8000
rect 35348 7960 35349 8000
rect 34444 7951 34484 7960
rect 35307 7951 35349 7960
rect 35308 7866 35348 7951
rect 34060 7708 34772 7748
rect 33928 7580 34296 7589
rect 33968 7540 34010 7580
rect 34050 7540 34092 7580
rect 34132 7540 34174 7580
rect 34214 7540 34256 7580
rect 33928 7531 34296 7540
rect 33771 7160 33813 7169
rect 33771 7120 33772 7160
rect 33812 7120 33813 7160
rect 33771 7111 33813 7120
rect 34635 7160 34677 7169
rect 34635 7120 34636 7160
rect 34676 7120 34677 7160
rect 34635 7111 34677 7120
rect 33772 6488 33812 7111
rect 34347 7076 34389 7085
rect 34347 7036 34348 7076
rect 34388 7036 34389 7076
rect 34347 7027 34389 7036
rect 33772 6439 33812 6448
rect 33964 6245 34004 6330
rect 33963 6236 34005 6245
rect 33963 6196 33964 6236
rect 34004 6196 34005 6236
rect 33963 6187 34005 6196
rect 33928 6068 34296 6077
rect 33968 6028 34010 6068
rect 34050 6028 34092 6068
rect 34132 6028 34174 6068
rect 34214 6028 34256 6068
rect 33928 6019 34296 6028
rect 34348 5900 34388 7027
rect 34636 7026 34676 7111
rect 34156 5860 34388 5900
rect 33771 5648 33813 5657
rect 33771 5608 33772 5648
rect 33812 5608 33813 5648
rect 33771 5599 33813 5608
rect 33291 5312 33333 5321
rect 33291 5272 33292 5312
rect 33332 5272 33333 5312
rect 33291 5263 33333 5272
rect 33675 5312 33717 5321
rect 33675 5272 33676 5312
rect 33716 5272 33717 5312
rect 33675 5263 33717 5272
rect 33196 4171 33236 4180
rect 32812 4086 32852 4171
rect 33004 3968 33044 3977
rect 32811 3884 32853 3893
rect 32811 3844 32812 3884
rect 32852 3844 32853 3884
rect 32811 3835 32853 3844
rect 32620 3760 32756 3800
rect 32523 2624 32565 2633
rect 32523 2584 32524 2624
rect 32564 2584 32565 2624
rect 32523 2575 32565 2584
rect 32524 2456 32564 2465
rect 32428 2416 32524 2456
rect 32524 2407 32564 2416
rect 32331 2372 32373 2381
rect 32331 2332 32332 2372
rect 32372 2332 32373 2372
rect 32331 2323 32373 2332
rect 32043 2120 32085 2129
rect 32043 2080 32044 2120
rect 32084 2080 32085 2120
rect 32620 2120 32660 3760
rect 32812 3464 32852 3835
rect 32812 3415 32852 3424
rect 33004 2885 33044 3928
rect 33099 3716 33141 3725
rect 33099 3676 33100 3716
rect 33140 3676 33141 3716
rect 33099 3667 33141 3676
rect 33003 2876 33045 2885
rect 33003 2836 33004 2876
rect 33044 2836 33045 2876
rect 33003 2827 33045 2836
rect 32907 2792 32949 2801
rect 32907 2752 32908 2792
rect 32948 2752 32949 2792
rect 32907 2743 32949 2752
rect 32716 2708 32756 2717
rect 32756 2668 32852 2708
rect 32716 2659 32756 2668
rect 32812 2540 32852 2668
rect 32908 2658 32948 2743
rect 33100 2624 33140 3667
rect 33292 3548 33332 5263
rect 33579 5228 33621 5237
rect 33579 5188 33580 5228
rect 33620 5188 33621 5228
rect 33579 5179 33621 5188
rect 33484 4962 33524 4971
rect 33388 4388 33428 4397
rect 33484 4388 33524 4922
rect 33428 4348 33524 4388
rect 33388 4339 33428 4348
rect 33580 4304 33620 5179
rect 33484 4264 33620 4304
rect 33676 5060 33716 5069
rect 33484 3884 33524 4264
rect 33676 4229 33716 5020
rect 33675 4220 33717 4229
rect 33675 4180 33676 4220
rect 33716 4180 33717 4220
rect 33675 4171 33717 4180
rect 33579 4136 33621 4145
rect 33579 4096 33580 4136
rect 33620 4096 33621 4136
rect 33579 4087 33621 4096
rect 33580 4002 33620 4087
rect 33484 3844 33716 3884
rect 33100 2540 33140 2584
rect 32812 2500 32948 2540
rect 32620 2080 32756 2120
rect 32043 2071 32085 2080
rect 32236 2036 32276 2045
rect 32276 1996 32660 2036
rect 32236 1987 32276 1996
rect 32044 1938 32084 1947
rect 32044 1289 32084 1898
rect 32523 1868 32565 1877
rect 32523 1828 32524 1868
rect 32564 1828 32565 1868
rect 32523 1819 32565 1828
rect 32620 1868 32660 1996
rect 32620 1819 32660 1828
rect 32331 1784 32373 1793
rect 32331 1744 32332 1784
rect 32372 1744 32373 1784
rect 32331 1735 32373 1744
rect 32139 1364 32181 1373
rect 32139 1324 32140 1364
rect 32180 1324 32181 1364
rect 32139 1315 32181 1324
rect 32043 1280 32085 1289
rect 32043 1240 32044 1280
rect 32084 1240 32085 1280
rect 32043 1231 32085 1240
rect 31756 988 31988 1028
rect 31659 860 31701 869
rect 31659 820 31660 860
rect 31700 820 31701 860
rect 31659 811 31701 820
rect 31756 80 31796 988
rect 31947 608 31989 617
rect 31947 568 31948 608
rect 31988 568 31989 608
rect 31947 559 31989 568
rect 31948 80 31988 559
rect 32140 80 32180 1315
rect 32332 1112 32372 1735
rect 32427 1700 32469 1709
rect 32427 1660 32428 1700
rect 32468 1660 32469 1700
rect 32427 1651 32469 1660
rect 32428 1566 32468 1651
rect 32332 1063 32372 1072
rect 32331 692 32373 701
rect 32331 652 32332 692
rect 32372 652 32373 692
rect 32331 643 32373 652
rect 32332 80 32372 643
rect 32524 80 32564 1819
rect 32619 1700 32661 1709
rect 32619 1660 32620 1700
rect 32660 1660 32661 1700
rect 32619 1651 32661 1660
rect 32620 1373 32660 1651
rect 32619 1364 32661 1373
rect 32619 1324 32620 1364
rect 32660 1324 32661 1364
rect 32619 1315 32661 1324
rect 32716 617 32756 2080
rect 32812 1700 32852 1709
rect 32812 1126 32852 1660
rect 32812 1077 32852 1086
rect 32908 1028 32948 2500
rect 33004 2500 33140 2540
rect 33196 3508 33332 3548
rect 33483 3548 33525 3557
rect 33483 3508 33484 3548
rect 33524 3508 33525 3548
rect 33196 2540 33236 3508
rect 33483 3499 33525 3508
rect 33292 3450 33332 3459
rect 33484 3414 33524 3499
rect 33292 2801 33332 3410
rect 33483 2876 33525 2885
rect 33483 2836 33484 2876
rect 33524 2836 33525 2876
rect 33483 2827 33525 2836
rect 33291 2792 33333 2801
rect 33291 2752 33292 2792
rect 33332 2752 33333 2792
rect 33291 2743 33333 2752
rect 33196 2500 33428 2540
rect 33004 1961 33044 2500
rect 33388 2456 33428 2500
rect 33100 2416 33428 2456
rect 33003 1952 33045 1961
rect 33003 1912 33004 1952
rect 33044 1912 33045 1952
rect 33003 1903 33045 1912
rect 33004 1818 33044 1903
rect 33004 1028 33044 1037
rect 32908 988 33004 1028
rect 33004 979 33044 988
rect 32907 776 32949 785
rect 32907 736 32908 776
rect 32948 736 32949 776
rect 32907 727 32949 736
rect 32715 608 32757 617
rect 32715 568 32716 608
rect 32756 568 32757 608
rect 32715 559 32757 568
rect 32715 188 32757 197
rect 32715 148 32716 188
rect 32756 148 32757 188
rect 32715 139 32757 148
rect 32716 80 32756 139
rect 32908 80 32948 727
rect 33100 80 33140 2416
rect 33291 2036 33333 2045
rect 33291 1996 33292 2036
rect 33332 1996 33333 2036
rect 33291 1987 33333 1996
rect 33195 1280 33237 1289
rect 33195 1240 33196 1280
rect 33236 1240 33237 1280
rect 33195 1231 33237 1240
rect 33196 1146 33236 1231
rect 33292 785 33332 1987
rect 33387 1952 33429 1961
rect 33387 1912 33388 1952
rect 33428 1912 33429 1952
rect 33387 1903 33429 1912
rect 33388 1112 33428 1903
rect 33484 1121 33524 2827
rect 33579 2372 33621 2381
rect 33579 2332 33580 2372
rect 33620 2332 33621 2372
rect 33579 2323 33621 2332
rect 33388 1063 33428 1072
rect 33483 1112 33525 1121
rect 33483 1072 33484 1112
rect 33524 1072 33525 1112
rect 33483 1063 33525 1072
rect 33291 776 33333 785
rect 33291 736 33292 776
rect 33332 736 33333 776
rect 33291 727 33333 736
rect 33580 608 33620 2323
rect 33292 568 33620 608
rect 33292 80 33332 568
rect 33484 80 33572 104
rect 28340 64 28360 80
rect 28280 0 28360 64
rect 28472 0 28552 80
rect 28664 0 28744 80
rect 28856 0 28936 80
rect 29048 0 29128 80
rect 29240 0 29320 80
rect 29432 0 29512 80
rect 29624 0 29704 80
rect 29816 0 29896 80
rect 30008 0 30088 80
rect 30200 0 30280 80
rect 30392 0 30472 80
rect 30584 0 30664 80
rect 30776 0 30856 80
rect 30968 0 31048 80
rect 31160 0 31240 80
rect 31352 0 31432 80
rect 31544 0 31624 80
rect 31736 0 31816 80
rect 31928 0 32008 80
rect 32120 0 32200 80
rect 32312 0 32392 80
rect 32504 0 32584 80
rect 32696 0 32776 80
rect 32888 0 32968 80
rect 33080 0 33160 80
rect 33272 0 33352 80
rect 33464 60 33572 80
rect 33676 60 33716 3844
rect 33772 1877 33812 5599
rect 34156 4985 34196 5860
rect 34539 5732 34581 5741
rect 34539 5692 34540 5732
rect 34580 5692 34581 5732
rect 34539 5683 34581 5692
rect 34155 4976 34197 4985
rect 34155 4936 34156 4976
rect 34196 4936 34197 4976
rect 34155 4927 34197 4936
rect 34156 4842 34196 4927
rect 34443 4808 34485 4817
rect 34443 4768 34444 4808
rect 34484 4768 34485 4808
rect 34443 4759 34485 4768
rect 33928 4556 34296 4565
rect 33968 4516 34010 4556
rect 34050 4516 34092 4556
rect 34132 4516 34174 4556
rect 34214 4516 34256 4556
rect 33928 4507 34296 4516
rect 34347 4388 34389 4397
rect 34347 4348 34348 4388
rect 34388 4348 34389 4388
rect 34347 4339 34389 4348
rect 33928 3044 34296 3053
rect 33968 3004 34010 3044
rect 34050 3004 34092 3044
rect 34132 3004 34174 3044
rect 34214 3004 34256 3044
rect 33928 2995 34296 3004
rect 34348 2885 34388 4339
rect 34444 3809 34484 4759
rect 34443 3800 34485 3809
rect 34443 3760 34444 3800
rect 34484 3760 34485 3800
rect 34443 3751 34485 3760
rect 34443 3464 34485 3473
rect 34443 3424 34444 3464
rect 34484 3424 34485 3464
rect 34443 3415 34485 3424
rect 34444 3330 34484 3415
rect 34540 3221 34580 5683
rect 34635 3548 34677 3557
rect 34635 3508 34636 3548
rect 34676 3508 34677 3548
rect 34635 3499 34677 3508
rect 34539 3212 34581 3221
rect 34539 3172 34540 3212
rect 34580 3172 34581 3212
rect 34539 3163 34581 3172
rect 34347 2876 34389 2885
rect 34347 2836 34348 2876
rect 34388 2836 34389 2876
rect 34347 2827 34389 2836
rect 34251 2792 34293 2801
rect 34251 2752 34252 2792
rect 34292 2752 34293 2792
rect 34251 2743 34293 2752
rect 34252 1952 34292 2743
rect 34348 2624 34388 2827
rect 34540 2801 34580 3163
rect 34539 2792 34581 2801
rect 34539 2752 34540 2792
rect 34580 2752 34581 2792
rect 34539 2743 34581 2752
rect 34348 2575 34388 2584
rect 34252 1903 34292 1912
rect 33771 1868 33813 1877
rect 33771 1828 33772 1868
rect 33812 1828 33813 1868
rect 33771 1819 33813 1828
rect 34636 1868 34676 3499
rect 34732 2633 34772 7708
rect 35116 7160 35156 7169
rect 34828 7076 34868 7085
rect 35116 7076 35156 7120
rect 34868 7036 35156 7076
rect 35212 7160 35252 7169
rect 34828 7027 34868 7036
rect 35212 6992 35252 7120
rect 35020 6952 35252 6992
rect 35596 7160 35636 7169
rect 35020 5993 35060 6952
rect 35168 6824 35536 6833
rect 35208 6784 35250 6824
rect 35290 6784 35332 6824
rect 35372 6784 35414 6824
rect 35454 6784 35496 6824
rect 35168 6775 35536 6784
rect 35019 5984 35061 5993
rect 35019 5944 35020 5984
rect 35060 5944 35061 5984
rect 35019 5935 35061 5944
rect 35403 5984 35445 5993
rect 35403 5944 35404 5984
rect 35444 5944 35445 5984
rect 35403 5935 35445 5944
rect 34827 5900 34869 5909
rect 34827 5860 34828 5900
rect 34868 5860 34869 5900
rect 34827 5851 34869 5860
rect 34828 4145 34868 5851
rect 35404 5657 35444 5935
rect 35308 5648 35348 5657
rect 35308 5480 35348 5608
rect 35403 5648 35445 5657
rect 35403 5608 35404 5648
rect 35444 5608 35445 5648
rect 35596 5648 35636 7120
rect 35692 7160 35732 7169
rect 35692 6917 35732 7120
rect 35691 6908 35733 6917
rect 35691 6868 35692 6908
rect 35732 6868 35733 6908
rect 35691 6859 35733 6868
rect 35883 6908 35925 6917
rect 35883 6868 35884 6908
rect 35924 6868 35925 6908
rect 35883 6859 35925 6868
rect 35884 5732 35924 6859
rect 35980 5825 36020 8464
rect 36171 7748 36213 7757
rect 36171 7708 36172 7748
rect 36212 7708 36213 7748
rect 36171 7699 36213 7708
rect 36172 7160 36212 7699
rect 36172 7111 36212 7120
rect 36075 6152 36117 6161
rect 36075 6112 36076 6152
rect 36116 6112 36117 6152
rect 36075 6103 36117 6112
rect 35979 5816 36021 5825
rect 35979 5776 35980 5816
rect 36020 5776 36021 5816
rect 35979 5767 36021 5776
rect 35884 5683 35924 5692
rect 35788 5648 35828 5657
rect 35596 5608 35788 5648
rect 35403 5599 35445 5608
rect 35308 5440 35636 5480
rect 35168 5312 35536 5321
rect 35208 5272 35250 5312
rect 35290 5272 35332 5312
rect 35372 5272 35414 5312
rect 35454 5272 35496 5312
rect 35168 5263 35536 5272
rect 35596 5144 35636 5440
rect 35788 5405 35828 5608
rect 35787 5396 35829 5405
rect 35787 5356 35788 5396
rect 35828 5356 35829 5396
rect 35787 5347 35829 5356
rect 35596 5095 35636 5104
rect 35787 5144 35829 5153
rect 35787 5104 35788 5144
rect 35828 5104 35829 5144
rect 35787 5095 35829 5104
rect 35404 4976 35444 4985
rect 35019 4472 35061 4481
rect 35019 4432 35020 4472
rect 35060 4432 35061 4472
rect 35019 4423 35061 4432
rect 34827 4136 34869 4145
rect 34827 4096 34828 4136
rect 34868 4096 34869 4136
rect 34827 4087 34869 4096
rect 35020 4136 35060 4423
rect 35404 4229 35444 4936
rect 35595 4892 35637 4901
rect 35595 4852 35596 4892
rect 35636 4852 35637 4892
rect 35595 4843 35637 4852
rect 35403 4220 35445 4229
rect 35403 4180 35404 4220
rect 35444 4180 35445 4220
rect 35403 4171 35445 4180
rect 35020 4087 35060 4096
rect 34828 4002 34868 4087
rect 35168 3800 35536 3809
rect 35208 3760 35250 3800
rect 35290 3760 35332 3800
rect 35372 3760 35414 3800
rect 35454 3760 35496 3800
rect 35168 3751 35536 3760
rect 35211 3044 35253 3053
rect 35211 3004 35212 3044
rect 35252 3004 35253 3044
rect 35211 2995 35253 3004
rect 35212 2633 35252 2995
rect 34731 2624 34773 2633
rect 34731 2584 34732 2624
rect 34772 2584 34773 2624
rect 34731 2575 34773 2584
rect 35211 2624 35253 2633
rect 35211 2584 35212 2624
rect 35252 2584 35253 2624
rect 35596 2624 35636 4843
rect 35691 3716 35733 3725
rect 35691 3676 35692 3716
rect 35732 3676 35733 3716
rect 35691 3667 35733 3676
rect 35692 3464 35732 3667
rect 35788 3473 35828 5095
rect 35884 4976 35924 4985
rect 36076 4976 36116 6103
rect 36268 5480 36308 8716
rect 36364 8707 36404 8716
rect 36748 8756 36788 8765
rect 36459 7748 36501 7757
rect 36459 7708 36460 7748
rect 36500 7708 36501 7748
rect 36459 7699 36501 7708
rect 36652 7748 36692 7757
rect 36363 6320 36405 6329
rect 36363 6280 36364 6320
rect 36404 6280 36405 6320
rect 36363 6271 36405 6280
rect 36364 6186 36404 6271
rect 36364 5648 36404 5657
rect 36460 5648 36500 7699
rect 36652 7174 36692 7708
rect 36652 7125 36692 7134
rect 36555 6404 36597 6413
rect 36555 6364 36556 6404
rect 36596 6364 36597 6404
rect 36555 6355 36597 6364
rect 36556 6270 36596 6355
rect 36404 5608 36500 5648
rect 36364 5599 36404 5608
rect 36748 5573 36788 8716
rect 36844 8504 36884 9043
rect 36940 8672 36980 8681
rect 36980 8632 37076 8672
rect 36940 8623 36980 8632
rect 36844 8464 36980 8504
rect 36844 8000 36884 8011
rect 36844 7925 36884 7960
rect 36843 7916 36885 7925
rect 36843 7876 36844 7916
rect 36884 7876 36885 7916
rect 36843 7867 36885 7876
rect 36844 6992 36884 7001
rect 36844 6413 36884 6952
rect 36940 6488 36980 8464
rect 37036 7421 37076 8632
rect 37323 8000 37365 8009
rect 37323 7960 37324 8000
rect 37364 7960 37365 8000
rect 37323 7951 37365 7960
rect 37035 7412 37077 7421
rect 37035 7372 37036 7412
rect 37076 7372 37077 7412
rect 37035 7363 37077 7372
rect 37324 6656 37364 7951
rect 37324 6607 37364 6616
rect 36940 6439 36980 6448
rect 36843 6404 36885 6413
rect 36843 6364 36844 6404
rect 36884 6364 36885 6404
rect 36843 6355 36885 6364
rect 36892 5657 36932 5666
rect 36932 5617 37364 5648
rect 36892 5608 37364 5617
rect 36747 5564 36789 5573
rect 36747 5524 36748 5564
rect 36788 5524 36789 5564
rect 36747 5515 36789 5524
rect 37036 5480 37076 5489
rect 36268 5440 36404 5480
rect 35924 4936 36116 4976
rect 35884 4229 35924 4936
rect 35883 4220 35925 4229
rect 35883 4180 35884 4220
rect 35924 4180 35925 4220
rect 35883 4171 35925 4180
rect 36267 4136 36309 4145
rect 36267 4096 36268 4136
rect 36308 4096 36309 4136
rect 36267 4087 36309 4096
rect 36268 4002 36308 4087
rect 35884 3548 35924 3557
rect 35924 3508 36212 3548
rect 35884 3499 35924 3508
rect 35692 3415 35732 3424
rect 35787 3464 35829 3473
rect 35787 3424 35788 3464
rect 35828 3424 35829 3464
rect 35787 3415 35829 3424
rect 36172 3464 36212 3508
rect 36172 3415 36212 3424
rect 36268 3464 36308 3473
rect 35883 3380 35925 3389
rect 35883 3340 35884 3380
rect 35924 3340 35925 3380
rect 35883 3331 35925 3340
rect 35884 2717 35924 3331
rect 35788 2708 35828 2717
rect 35596 2584 35732 2624
rect 35211 2575 35253 2584
rect 35596 2456 35636 2465
rect 35168 2288 35536 2297
rect 35208 2248 35250 2288
rect 35290 2248 35332 2288
rect 35372 2248 35414 2288
rect 35454 2248 35496 2288
rect 35168 2239 35536 2248
rect 34636 1819 34676 1828
rect 35308 1952 35348 1961
rect 34444 1700 34484 1709
rect 33928 1532 34296 1541
rect 33968 1492 34010 1532
rect 34050 1492 34092 1532
rect 34132 1492 34174 1532
rect 34214 1492 34256 1532
rect 33928 1483 34296 1492
rect 34444 281 34484 1660
rect 35308 1289 35348 1912
rect 35403 1952 35445 1961
rect 35403 1912 35404 1952
rect 35444 1912 35445 1952
rect 35403 1903 35445 1912
rect 35404 1818 35444 1903
rect 34827 1280 34869 1289
rect 34827 1240 34828 1280
rect 34868 1240 34869 1280
rect 34827 1231 34869 1240
rect 35307 1280 35349 1289
rect 35307 1240 35308 1280
rect 35348 1240 35349 1280
rect 35307 1231 35349 1240
rect 34828 1146 34868 1231
rect 34635 1112 34677 1121
rect 34635 1072 34636 1112
rect 34676 1072 34677 1112
rect 34635 1063 34677 1072
rect 35020 1112 35060 1121
rect 34636 978 34676 1063
rect 35020 701 35060 1072
rect 35168 776 35536 785
rect 35208 736 35250 776
rect 35290 736 35332 776
rect 35372 736 35414 776
rect 35454 736 35496 776
rect 35168 727 35536 736
rect 35019 692 35061 701
rect 35019 652 35020 692
rect 35060 652 35061 692
rect 35019 643 35061 652
rect 35596 449 35636 2416
rect 35692 1961 35732 2584
rect 35788 2297 35828 2668
rect 35883 2708 35925 2717
rect 35883 2668 35884 2708
rect 35924 2668 35925 2708
rect 35883 2659 35925 2668
rect 35787 2288 35829 2297
rect 35787 2248 35788 2288
rect 35828 2248 35829 2288
rect 35787 2239 35829 2248
rect 35884 2036 35924 2659
rect 36076 2633 36116 2718
rect 36075 2624 36117 2633
rect 36075 2584 36076 2624
rect 36116 2584 36117 2624
rect 36075 2575 36117 2584
rect 36172 2624 36212 2633
rect 36268 2624 36308 3424
rect 36364 3137 36404 5440
rect 36844 5440 37036 5480
rect 36844 4220 36884 5440
rect 37036 5431 37076 5440
rect 37324 5144 37364 5608
rect 37324 5095 37364 5104
rect 36844 4171 36884 4180
rect 37132 4976 37172 4985
rect 37132 4145 37172 4936
rect 36939 4136 36981 4145
rect 36939 4096 36940 4136
rect 36980 4096 36981 4136
rect 36939 4087 36981 4096
rect 37131 4136 37173 4145
rect 37131 4096 37132 4136
rect 37172 4096 37173 4136
rect 37131 4087 37173 4096
rect 37228 4136 37268 4145
rect 37268 4096 37364 4136
rect 37228 4087 37268 4096
rect 36460 3968 36500 3977
rect 36363 3128 36405 3137
rect 36363 3088 36364 3128
rect 36404 3088 36405 3128
rect 36363 3079 36405 3088
rect 36363 2792 36405 2801
rect 36363 2752 36364 2792
rect 36404 2752 36405 2792
rect 36363 2743 36405 2752
rect 36212 2584 36308 2624
rect 35788 1996 35924 2036
rect 35691 1952 35733 1961
rect 35691 1912 35692 1952
rect 35732 1912 35733 1952
rect 35691 1903 35733 1912
rect 35788 1952 35828 1996
rect 35788 1903 35828 1912
rect 36172 1877 36212 2584
rect 36364 1952 36404 2743
rect 36460 2633 36500 3928
rect 36651 3968 36693 3977
rect 36651 3928 36652 3968
rect 36692 3928 36693 3968
rect 36651 3919 36693 3928
rect 36652 3834 36692 3919
rect 36747 3632 36789 3641
rect 36747 3592 36748 3632
rect 36788 3592 36789 3632
rect 36747 3583 36789 3592
rect 36748 3464 36788 3583
rect 36555 3380 36597 3389
rect 36555 3340 36556 3380
rect 36596 3340 36597 3380
rect 36555 3331 36597 3340
rect 36652 3380 36692 3389
rect 36556 2969 36596 3331
rect 36555 2960 36597 2969
rect 36555 2920 36556 2960
rect 36596 2920 36597 2960
rect 36555 2911 36597 2920
rect 36652 2792 36692 3340
rect 36748 2801 36788 3424
rect 36574 2752 36692 2792
rect 36747 2792 36789 2801
rect 36747 2752 36748 2792
rect 36788 2752 36789 2792
rect 36574 2717 36614 2752
rect 36747 2743 36789 2752
rect 36555 2708 36614 2717
rect 36555 2668 36556 2708
rect 36596 2668 36614 2708
rect 36555 2659 36597 2668
rect 36459 2624 36501 2633
rect 36459 2584 36460 2624
rect 36500 2584 36501 2624
rect 36459 2575 36501 2584
rect 36556 2574 36596 2659
rect 36652 2624 36692 2633
rect 36748 2624 36788 2743
rect 36692 2584 36788 2624
rect 36652 2575 36692 2584
rect 36364 1903 36404 1912
rect 36844 1938 36884 1947
rect 35883 1868 35925 1877
rect 35883 1828 35884 1868
rect 35924 1828 35925 1868
rect 35883 1819 35925 1828
rect 36171 1868 36213 1877
rect 36171 1828 36172 1868
rect 36212 1828 36213 1868
rect 36171 1819 36213 1828
rect 35884 1734 35924 1819
rect 36844 1289 36884 1898
rect 36459 1280 36501 1289
rect 36459 1240 36460 1280
rect 36500 1240 36501 1280
rect 36459 1231 36501 1240
rect 36843 1280 36885 1289
rect 36843 1240 36844 1280
rect 36884 1240 36885 1280
rect 36843 1231 36885 1240
rect 36460 1146 36500 1231
rect 36267 1112 36309 1121
rect 36267 1072 36268 1112
rect 36308 1072 36309 1112
rect 36267 1063 36309 1072
rect 36652 1112 36692 1121
rect 36940 1112 36980 4087
rect 37228 3464 37268 3473
rect 37131 3044 37173 3053
rect 37228 3044 37268 3424
rect 37324 3389 37364 4096
rect 37708 3473 37748 3554
rect 37707 3464 37749 3473
rect 37707 3419 37708 3464
rect 37748 3419 37749 3464
rect 37707 3415 37749 3419
rect 37708 3410 37748 3415
rect 37323 3380 37365 3389
rect 37323 3340 37324 3380
rect 37364 3340 37365 3380
rect 37804 3380 37844 9388
rect 37900 9379 37940 9388
rect 38668 8840 38708 10672
rect 39820 9596 39860 10672
rect 40011 9848 40053 9857
rect 40011 9808 40012 9848
rect 40052 9808 40053 9848
rect 40011 9799 40053 9808
rect 39148 9556 39860 9596
rect 38764 8840 38804 8849
rect 38668 8800 38764 8840
rect 38764 8791 38804 8800
rect 39148 8840 39188 9556
rect 39148 8791 39188 8800
rect 40012 8840 40052 9799
rect 40012 8791 40052 8800
rect 40396 8840 40436 10692
rect 40866 10688 40906 10692
rect 40952 10688 41032 10752
rect 40866 10672 41032 10688
rect 40866 10648 41012 10672
rect 40683 10520 40725 10529
rect 40683 10480 40684 10520
rect 40724 10480 40725 10520
rect 40683 10471 40725 10480
rect 40684 9680 40724 10471
rect 41451 10184 41493 10193
rect 41451 10144 41452 10184
rect 41492 10144 41493 10184
rect 41451 10135 41493 10144
rect 40684 9631 40724 9640
rect 41259 9680 41301 9689
rect 41259 9640 41260 9680
rect 41300 9640 41301 9680
rect 41259 9631 41301 9640
rect 41452 9680 41492 10135
rect 41452 9631 41492 9640
rect 41067 9512 41109 9521
rect 41067 9472 41068 9512
rect 41108 9472 41109 9512
rect 41067 9463 41109 9472
rect 40396 8791 40436 8800
rect 40492 9428 40532 9437
rect 38475 8756 38517 8765
rect 38475 8716 38476 8756
rect 38516 8716 38517 8756
rect 38475 8707 38517 8716
rect 38572 8756 38612 8765
rect 38188 8672 38228 8681
rect 38188 8588 38228 8632
rect 37900 8548 38228 8588
rect 37900 7925 37940 8548
rect 38380 8504 38420 8513
rect 37996 8464 38380 8504
rect 37899 7916 37941 7925
rect 37899 7876 37900 7916
rect 37940 7876 37941 7916
rect 37899 7867 37941 7876
rect 37900 6413 37940 7867
rect 37996 7160 38036 8464
rect 38380 8455 38420 8464
rect 38091 8000 38133 8009
rect 38091 7960 38092 8000
rect 38132 7960 38133 8000
rect 38091 7951 38133 7960
rect 38092 7673 38132 7951
rect 38091 7664 38133 7673
rect 38091 7624 38092 7664
rect 38132 7624 38133 7664
rect 38091 7615 38133 7624
rect 38476 7244 38516 8707
rect 38572 8093 38612 8716
rect 38956 8756 38996 8765
rect 38571 8084 38613 8093
rect 38571 8044 38572 8084
rect 38612 8044 38613 8084
rect 38571 8035 38613 8044
rect 37996 7111 38036 7120
rect 38092 7160 38132 7169
rect 38132 7120 38420 7160
rect 38092 7111 38132 7120
rect 37995 6488 38037 6497
rect 37995 6448 37996 6488
rect 38036 6448 38037 6488
rect 37995 6439 38037 6448
rect 37899 6404 37941 6413
rect 37899 6364 37900 6404
rect 37940 6364 37941 6404
rect 37899 6355 37941 6364
rect 37996 6354 38036 6439
rect 38091 6404 38133 6413
rect 38091 6364 38092 6404
rect 38132 6364 38133 6404
rect 38091 6355 38133 6364
rect 38092 3725 38132 6355
rect 38380 5144 38420 7120
rect 38188 5104 38420 5144
rect 38188 4061 38228 5104
rect 38284 4976 38324 4985
rect 38187 4052 38229 4061
rect 38187 4012 38188 4052
rect 38228 4012 38229 4052
rect 38187 4003 38229 4012
rect 38284 3977 38324 4936
rect 38380 4976 38420 5104
rect 38380 4927 38420 4936
rect 38476 4976 38516 7204
rect 38571 7160 38613 7169
rect 38571 7120 38572 7160
rect 38612 7120 38613 7160
rect 38571 7111 38613 7120
rect 38859 7160 38901 7169
rect 38859 7120 38860 7160
rect 38900 7120 38901 7160
rect 38859 7111 38901 7120
rect 38572 7026 38612 7111
rect 38764 4976 38804 4985
rect 38476 4936 38764 4976
rect 38476 4304 38516 4936
rect 38764 4927 38804 4936
rect 38860 4892 38900 7111
rect 38860 4472 38900 4852
rect 38764 4432 38900 4472
rect 38476 4264 38612 4304
rect 38475 4136 38517 4145
rect 38475 4096 38476 4136
rect 38516 4096 38517 4136
rect 38475 4087 38517 4096
rect 38379 4052 38421 4061
rect 38379 4012 38380 4052
rect 38420 4012 38421 4052
rect 38379 4003 38421 4012
rect 38283 3968 38325 3977
rect 38283 3928 38284 3968
rect 38324 3928 38325 3968
rect 38283 3919 38325 3928
rect 38091 3716 38133 3725
rect 38091 3676 38092 3716
rect 38132 3676 38133 3716
rect 38091 3667 38133 3676
rect 38283 3716 38325 3725
rect 38283 3676 38284 3716
rect 38324 3676 38325 3716
rect 38283 3667 38325 3676
rect 37900 3548 37940 3557
rect 37940 3508 38228 3548
rect 37900 3499 37940 3508
rect 37804 3340 37940 3380
rect 37323 3331 37365 3340
rect 37131 3004 37132 3044
rect 37172 3004 37268 3044
rect 37131 2995 37173 3004
rect 37132 2624 37172 2995
rect 37612 2633 37652 2719
rect 37132 2575 37172 2584
rect 37611 2629 37653 2633
rect 37611 2584 37612 2629
rect 37652 2584 37653 2629
rect 37611 2575 37653 2584
rect 37804 2540 37844 2568
rect 37708 2500 37804 2540
rect 37035 2288 37077 2297
rect 37035 2248 37036 2288
rect 37076 2248 37077 2288
rect 37035 2239 37077 2248
rect 37036 2120 37076 2239
rect 37036 2071 37076 2080
rect 37708 1868 37748 2500
rect 37804 2491 37844 2500
rect 37900 2045 37940 3340
rect 38091 3296 38133 3305
rect 38091 3256 38092 3296
rect 38132 3256 38133 3296
rect 38091 3247 38133 3256
rect 38092 3162 38132 3247
rect 38188 2708 38228 3508
rect 38284 3464 38324 3667
rect 38284 3415 38324 3424
rect 38188 2659 38228 2668
rect 37996 2456 38036 2465
rect 37899 2036 37941 2045
rect 37899 1996 37900 2036
rect 37940 1996 37941 2036
rect 37899 1987 37941 1996
rect 37708 1819 37748 1828
rect 36692 1072 36980 1112
rect 36268 953 36308 1063
rect 36267 944 36309 953
rect 36267 904 36268 944
rect 36308 904 36309 944
rect 36267 895 36309 904
rect 36652 701 36692 1072
rect 36940 953 36980 1072
rect 37516 1700 37556 1709
rect 36939 944 36981 953
rect 36939 904 36940 944
rect 36980 904 36981 944
rect 36939 895 36981 904
rect 36651 692 36693 701
rect 36651 652 36652 692
rect 36692 652 36693 692
rect 36651 643 36693 652
rect 35595 440 35637 449
rect 35595 400 35596 440
rect 35636 400 35637 440
rect 35595 391 35637 400
rect 37516 365 37556 1660
rect 37996 1625 38036 2416
rect 38284 1952 38324 1961
rect 37995 1616 38037 1625
rect 37995 1576 37996 1616
rect 38036 1576 38037 1616
rect 37995 1567 38037 1576
rect 38092 1364 38132 1373
rect 38284 1364 38324 1912
rect 38380 1952 38420 4003
rect 38476 4002 38516 4087
rect 38572 3212 38612 4264
rect 38667 3968 38709 3977
rect 38667 3928 38668 3968
rect 38708 3928 38709 3968
rect 38667 3919 38709 3928
rect 38668 3834 38708 3919
rect 38572 3172 38708 3212
rect 38380 1903 38420 1912
rect 38572 2708 38612 2717
rect 38132 1324 38324 1364
rect 38092 1315 38132 1324
rect 38572 1205 38612 2668
rect 38668 1952 38708 3172
rect 38764 3128 38804 4432
rect 38859 4304 38901 4313
rect 38859 4264 38860 4304
rect 38900 4264 38901 4304
rect 38859 4255 38901 4264
rect 38860 4136 38900 4255
rect 38860 4061 38900 4096
rect 38859 4052 38901 4061
rect 38859 4012 38860 4052
rect 38900 4012 38901 4052
rect 38859 4003 38901 4012
rect 38956 3548 38996 8716
rect 39819 8756 39861 8765
rect 39819 8716 39820 8756
rect 39860 8716 39861 8756
rect 39819 8707 39861 8716
rect 40204 8756 40244 8765
rect 39820 8622 39860 8707
rect 39052 7160 39092 7169
rect 39052 5825 39092 7120
rect 39532 7165 39572 7174
rect 39436 6656 39476 6665
rect 39532 6656 39572 7125
rect 39476 6616 39572 6656
rect 39724 6992 39764 7001
rect 39436 6607 39476 6616
rect 39244 6488 39284 6499
rect 39244 6413 39284 6448
rect 39243 6404 39285 6413
rect 39243 6364 39244 6404
rect 39284 6364 39285 6404
rect 39724 6404 39764 6952
rect 39820 6404 39860 6413
rect 39724 6364 39820 6404
rect 39243 6355 39285 6364
rect 39820 6355 39860 6364
rect 39627 6320 39669 6329
rect 39627 6280 39628 6320
rect 39668 6280 39669 6320
rect 39627 6271 39669 6280
rect 39628 6186 39668 6271
rect 39051 5816 39093 5825
rect 39051 5776 39052 5816
rect 39092 5776 39093 5816
rect 39051 5767 39093 5776
rect 39052 4976 39092 5767
rect 39435 5648 39477 5657
rect 39435 5608 39436 5648
rect 39476 5608 39477 5648
rect 39435 5599 39477 5608
rect 39340 4976 39380 4985
rect 39052 4936 39340 4976
rect 39340 4927 39380 4936
rect 39147 4136 39189 4145
rect 39147 4096 39148 4136
rect 39188 4096 39189 4136
rect 39147 4087 39189 4096
rect 38956 3508 39092 3548
rect 38764 3088 38900 3128
rect 38764 2456 38804 2465
rect 38764 2129 38804 2416
rect 38763 2120 38805 2129
rect 38763 2080 38764 2120
rect 38804 2080 38805 2120
rect 38763 2071 38805 2080
rect 38764 1952 38804 1961
rect 38668 1912 38764 1952
rect 38764 1903 38804 1912
rect 38860 1952 38900 3088
rect 38956 2549 38996 2634
rect 38955 2540 38997 2549
rect 38955 2500 38956 2540
rect 38996 2500 38997 2540
rect 38955 2491 38997 2500
rect 39052 2381 39092 3508
rect 39148 2624 39188 4087
rect 39148 2575 39188 2584
rect 39436 2540 39476 5599
rect 40204 5237 40244 8716
rect 40492 8597 40532 9388
rect 40875 9428 40917 9437
rect 40875 9388 40876 9428
rect 40916 9388 40917 9428
rect 40875 9379 40917 9388
rect 40876 9294 40916 9379
rect 41068 9344 41108 9463
rect 41260 9428 41300 9631
rect 41260 9379 41300 9388
rect 41068 9295 41108 9304
rect 41451 9092 41493 9101
rect 41451 9052 41452 9092
rect 41492 9052 41493 9092
rect 41451 9043 41493 9052
rect 41067 8840 41109 8849
rect 41067 8800 41068 8840
rect 41108 8800 41109 8840
rect 41067 8791 41109 8800
rect 41452 8840 41492 9043
rect 41452 8791 41492 8800
rect 40876 8756 40916 8765
rect 40491 8588 40533 8597
rect 40491 8548 40492 8588
rect 40532 8548 40533 8588
rect 40491 8539 40533 8548
rect 40876 8429 40916 8716
rect 41068 8706 41108 8791
rect 41260 8756 41300 8765
rect 40875 8420 40917 8429
rect 40875 8380 40876 8420
rect 40916 8380 40917 8420
rect 40875 8371 40917 8380
rect 41260 8261 41300 8716
rect 41451 8504 41493 8513
rect 41451 8464 41452 8504
rect 41492 8464 41493 8504
rect 41451 8455 41493 8464
rect 41259 8252 41301 8261
rect 41259 8212 41260 8252
rect 41300 8212 41301 8252
rect 41259 8203 41301 8212
rect 40683 8168 40725 8177
rect 40683 8128 40684 8168
rect 40724 8128 40725 8168
rect 40683 8119 40725 8128
rect 41452 8168 41492 8455
rect 41452 8119 41492 8128
rect 40684 8034 40724 8119
rect 40491 7916 40533 7925
rect 40876 7916 40916 7925
rect 40491 7876 40492 7916
rect 40532 7876 40533 7916
rect 40491 7867 40533 7876
rect 40780 7876 40876 7916
rect 40492 7782 40532 7867
rect 40683 7496 40725 7505
rect 40683 7456 40684 7496
rect 40724 7456 40725 7496
rect 40683 7447 40725 7456
rect 40491 7412 40533 7421
rect 40491 7372 40492 7412
rect 40532 7372 40533 7412
rect 40491 7363 40533 7372
rect 40684 7412 40724 7447
rect 40492 7244 40532 7363
rect 40684 7361 40724 7372
rect 40492 7195 40532 7204
rect 40683 6824 40725 6833
rect 40683 6784 40684 6824
rect 40724 6784 40725 6824
rect 40683 6775 40725 6784
rect 40684 6656 40724 6775
rect 40684 6607 40724 6616
rect 40780 6497 40820 7876
rect 40876 7867 40916 7876
rect 41259 7916 41301 7925
rect 41259 7876 41260 7916
rect 41300 7876 41301 7916
rect 41259 7867 41301 7876
rect 41067 7832 41109 7841
rect 41067 7792 41068 7832
rect 41108 7792 41109 7832
rect 41067 7783 41109 7792
rect 41068 7698 41108 7783
rect 41260 7782 41300 7867
rect 40876 7244 40916 7253
rect 40916 7204 41012 7244
rect 40876 7195 40916 7204
rect 40875 6740 40917 6749
rect 40875 6700 40876 6740
rect 40916 6700 40917 6740
rect 40875 6691 40917 6700
rect 40779 6488 40821 6497
rect 40779 6448 40780 6488
rect 40820 6448 40821 6488
rect 40779 6439 40821 6448
rect 40492 6404 40532 6413
rect 40396 6364 40492 6404
rect 40203 5228 40245 5237
rect 40203 5188 40204 5228
rect 40244 5188 40245 5228
rect 40203 5179 40245 5188
rect 40396 5153 40436 6364
rect 40492 6355 40532 6364
rect 40876 6404 40916 6691
rect 40876 6355 40916 6364
rect 40683 5816 40725 5825
rect 40683 5776 40684 5816
rect 40724 5776 40725 5816
rect 40683 5767 40725 5776
rect 40491 5732 40533 5741
rect 40491 5692 40492 5732
rect 40532 5692 40533 5732
rect 40491 5683 40533 5692
rect 40492 5598 40532 5683
rect 40684 5682 40724 5767
rect 40876 5732 40916 5741
rect 40876 5489 40916 5692
rect 40875 5480 40917 5489
rect 40875 5440 40876 5480
rect 40916 5440 40917 5480
rect 40875 5431 40917 5440
rect 40395 5144 40437 5153
rect 40395 5104 40396 5144
rect 40436 5104 40437 5144
rect 40395 5095 40437 5104
rect 40683 5144 40725 5153
rect 40683 5104 40684 5144
rect 40724 5104 40725 5144
rect 40683 5095 40725 5104
rect 40012 5060 40052 5069
rect 39820 4962 39860 4971
rect 39820 4397 39860 4922
rect 39819 4388 39861 4397
rect 39819 4348 39820 4388
rect 39860 4348 39861 4388
rect 39819 4339 39861 4348
rect 39531 3548 39573 3557
rect 39531 3508 39532 3548
rect 39572 3508 39573 3548
rect 39531 3499 39573 3508
rect 39532 3464 39572 3499
rect 39532 3413 39572 3424
rect 39916 3380 39956 3389
rect 40012 3380 40052 5020
rect 40395 4976 40437 4985
rect 40395 4936 40396 4976
rect 40436 4936 40437 4976
rect 40395 4927 40437 4936
rect 40299 4388 40341 4397
rect 40299 4348 40300 4388
rect 40340 4348 40341 4388
rect 40299 4339 40341 4348
rect 40300 4254 40340 4339
rect 40396 4220 40436 4927
rect 40492 4892 40532 4901
rect 40492 4649 40532 4852
rect 40684 4808 40724 5095
rect 40875 4892 40917 4901
rect 40875 4852 40876 4892
rect 40916 4852 40917 4892
rect 40875 4843 40917 4852
rect 40684 4759 40724 4768
rect 40876 4758 40916 4843
rect 40491 4640 40533 4649
rect 40491 4600 40492 4640
rect 40532 4600 40533 4640
rect 40491 4591 40533 4600
rect 40492 4220 40532 4229
rect 40396 4180 40492 4220
rect 40492 4171 40532 4180
rect 40875 4220 40917 4229
rect 40875 4180 40876 4220
rect 40916 4180 40917 4220
rect 40875 4171 40917 4180
rect 40107 4136 40149 4145
rect 40107 4096 40108 4136
rect 40148 4096 40149 4136
rect 40107 4087 40149 4096
rect 40683 4136 40725 4145
rect 40683 4096 40684 4136
rect 40724 4096 40725 4136
rect 40683 4087 40725 4096
rect 40108 3809 40148 4087
rect 40684 3968 40724 4087
rect 40876 4086 40916 4171
rect 40684 3919 40724 3928
rect 40107 3800 40149 3809
rect 40107 3760 40108 3800
rect 40148 3760 40149 3800
rect 40107 3751 40149 3760
rect 40587 3800 40629 3809
rect 40587 3760 40588 3800
rect 40628 3760 40629 3800
rect 40587 3751 40629 3760
rect 40491 3632 40533 3641
rect 40491 3592 40492 3632
rect 40532 3592 40533 3632
rect 40491 3583 40533 3592
rect 39956 3340 40052 3380
rect 40108 3380 40148 3389
rect 40492 3380 40532 3583
rect 39916 3331 39956 3340
rect 39244 2500 39476 2540
rect 39724 3212 39764 3221
rect 39051 2372 39093 2381
rect 39051 2332 39052 2372
rect 39092 2332 39093 2372
rect 39051 2323 39093 2332
rect 38955 2120 38997 2129
rect 38955 2080 38956 2120
rect 38996 2080 38997 2120
rect 38955 2071 38997 2080
rect 38860 1903 38900 1912
rect 38956 1457 38996 2071
rect 39244 1952 39284 2500
rect 39724 2213 39764 3172
rect 40108 2288 40148 3340
rect 40396 3340 40492 3380
rect 39820 2248 40148 2288
rect 40300 3212 40340 3221
rect 39723 2204 39765 2213
rect 39723 2164 39724 2204
rect 39764 2164 39765 2204
rect 39723 2155 39765 2164
rect 39820 2036 39860 2248
rect 39916 2164 40244 2204
rect 39916 2036 39956 2164
rect 40204 2120 40244 2164
rect 40204 2071 40244 2080
rect 39724 1996 39860 2036
rect 39905 1996 39956 2036
rect 40012 2036 40052 2045
rect 39340 1952 39380 1961
rect 39244 1912 39340 1952
rect 39340 1903 39380 1912
rect 38955 1448 38997 1457
rect 38955 1408 38956 1448
rect 38996 1408 38997 1448
rect 38955 1399 38997 1408
rect 38571 1196 38613 1205
rect 38571 1156 38572 1196
rect 38612 1156 38613 1196
rect 38571 1147 38613 1156
rect 39531 1196 39573 1205
rect 39531 1156 39532 1196
rect 39572 1156 39573 1196
rect 39531 1147 39573 1156
rect 37900 1112 37940 1121
rect 37900 869 37940 1072
rect 38284 1112 38324 1121
rect 38284 953 38324 1072
rect 39532 1112 39572 1147
rect 39724 1121 39764 1996
rect 39905 1952 39945 1996
rect 39820 1942 39945 1952
rect 39860 1912 39945 1942
rect 39820 1893 39860 1902
rect 39916 1196 39956 1205
rect 40012 1196 40052 1996
rect 39956 1156 40052 1196
rect 40108 1196 40148 1205
rect 39916 1147 39956 1156
rect 39532 1061 39572 1072
rect 39723 1112 39765 1121
rect 39723 1072 39724 1112
rect 39764 1072 39765 1112
rect 39723 1063 39765 1072
rect 38283 944 38325 953
rect 38283 904 38284 944
rect 38324 904 38325 944
rect 38283 895 38325 904
rect 39724 944 39764 953
rect 37899 860 37941 869
rect 37899 820 37900 860
rect 37940 820 37941 860
rect 37899 811 37941 820
rect 37515 356 37557 365
rect 37515 316 37516 356
rect 37556 316 37557 356
rect 37515 307 37557 316
rect 34443 272 34485 281
rect 34443 232 34444 272
rect 34484 232 34485 272
rect 34443 223 34485 232
rect 39724 113 39764 904
rect 40108 869 40148 1156
rect 40300 1121 40340 3172
rect 40396 2624 40436 3340
rect 40492 3331 40532 3340
rect 40396 2575 40436 2584
rect 40588 2456 40628 3751
rect 40972 3557 41012 7204
rect 41067 7160 41109 7169
rect 41067 7120 41068 7160
rect 41108 7120 41109 7160
rect 41067 7111 41109 7120
rect 41068 6992 41108 7111
rect 41068 6943 41108 6952
rect 41067 6488 41109 6497
rect 41067 6448 41068 6488
rect 41108 6448 41109 6488
rect 41067 6439 41109 6448
rect 41068 6320 41108 6439
rect 41163 6404 41205 6413
rect 41163 6364 41164 6404
rect 41204 6364 41205 6404
rect 41163 6355 41205 6364
rect 41068 6271 41108 6280
rect 41067 6152 41109 6161
rect 41067 6112 41068 6152
rect 41108 6112 41109 6152
rect 41067 6103 41109 6112
rect 41068 5900 41108 6103
rect 41068 5851 41108 5860
rect 41067 5480 41109 5489
rect 41067 5440 41068 5480
rect 41108 5440 41109 5480
rect 41067 5431 41109 5440
rect 41068 4808 41108 5431
rect 41068 4759 41108 4768
rect 41067 4472 41109 4481
rect 41067 4432 41068 4472
rect 41108 4432 41109 4472
rect 41067 4423 41109 4432
rect 41068 4388 41108 4423
rect 41068 4337 41108 4348
rect 40971 3548 41013 3557
rect 40971 3508 40972 3548
rect 41012 3508 41013 3548
rect 40971 3499 41013 3508
rect 41067 3464 41109 3473
rect 41067 3424 41068 3464
rect 41108 3424 41109 3464
rect 41067 3415 41109 3424
rect 40875 3380 40917 3389
rect 40875 3340 40876 3380
rect 40916 3340 40917 3380
rect 40875 3331 40917 3340
rect 40876 3246 40916 3331
rect 41068 3296 41108 3415
rect 41164 3380 41204 6355
rect 41260 4892 41300 4901
rect 41260 4733 41300 4852
rect 41451 4808 41493 4817
rect 41451 4768 41452 4808
rect 41492 4768 41493 4808
rect 41451 4759 41493 4768
rect 41259 4724 41301 4733
rect 41259 4684 41260 4724
rect 41300 4684 41301 4724
rect 41259 4675 41301 4684
rect 41452 4674 41492 4759
rect 41260 4220 41300 4229
rect 41260 4061 41300 4180
rect 41259 4052 41301 4061
rect 41259 4012 41260 4052
rect 41300 4012 41301 4052
rect 41259 4003 41301 4012
rect 41452 3968 41492 3977
rect 41452 3809 41492 3928
rect 41451 3800 41493 3809
rect 41451 3760 41452 3800
rect 41492 3760 41493 3800
rect 41451 3751 41493 3760
rect 41260 3380 41300 3389
rect 41164 3340 41260 3380
rect 41260 3331 41300 3340
rect 41068 3247 41108 3256
rect 40683 3212 40725 3221
rect 40683 3172 40684 3212
rect 40724 3172 40725 3212
rect 40683 3163 40725 3172
rect 41452 3212 41492 3221
rect 41492 3172 41588 3212
rect 41452 3163 41492 3172
rect 40684 3078 40724 3163
rect 41259 3044 41301 3053
rect 41259 3004 41260 3044
rect 41300 3004 41301 3044
rect 41259 2995 41301 3004
rect 40875 2876 40917 2885
rect 40875 2836 40876 2876
rect 40916 2836 40917 2876
rect 40875 2827 40917 2836
rect 40876 2708 40916 2827
rect 41067 2792 41109 2801
rect 41067 2752 41068 2792
rect 41108 2752 41109 2792
rect 41067 2743 41109 2752
rect 40876 2659 40916 2668
rect 41068 2658 41108 2743
rect 41260 2708 41300 2995
rect 41260 2659 41300 2668
rect 40396 2416 40628 2456
rect 41451 2456 41493 2465
rect 41451 2416 41452 2456
rect 41492 2416 41493 2456
rect 40396 1952 40436 2416
rect 41451 2407 41493 2416
rect 41452 2322 41492 2407
rect 41548 2129 41588 3172
rect 41547 2120 41589 2129
rect 41547 2080 41548 2120
rect 41588 2080 41589 2120
rect 41547 2071 41589 2080
rect 40396 1903 40436 1912
rect 41644 1952 41684 1961
rect 41067 1784 41109 1793
rect 41067 1744 41068 1784
rect 41108 1744 41109 1784
rect 41067 1735 41109 1744
rect 40876 1289 40916 1320
rect 40875 1280 40917 1289
rect 40875 1240 40876 1280
rect 40916 1240 40917 1280
rect 40875 1231 40917 1240
rect 41068 1280 41108 1735
rect 41644 1289 41684 1912
rect 41068 1231 41108 1240
rect 41643 1280 41685 1289
rect 41643 1240 41644 1280
rect 41684 1240 41685 1280
rect 41643 1231 41685 1240
rect 40491 1196 40533 1205
rect 40491 1156 40492 1196
rect 40532 1156 40533 1196
rect 40491 1147 40533 1156
rect 40876 1196 40916 1231
rect 40299 1112 40341 1121
rect 40299 1072 40300 1112
rect 40340 1072 40341 1112
rect 40299 1063 40341 1072
rect 40492 1062 40532 1147
rect 40876 1037 40916 1156
rect 41259 1196 41301 1205
rect 41259 1156 41260 1196
rect 41300 1156 41301 1196
rect 41259 1147 41301 1156
rect 41260 1062 41300 1147
rect 40875 1028 40917 1037
rect 40875 988 40876 1028
rect 40916 988 40917 1028
rect 40875 979 40917 988
rect 40300 944 40340 953
rect 40107 860 40149 869
rect 40107 820 40108 860
rect 40148 820 40149 860
rect 40107 811 40149 820
rect 40300 785 40340 904
rect 40684 944 40724 953
rect 40299 776 40341 785
rect 40299 736 40300 776
rect 40340 736 40341 776
rect 40299 727 40341 736
rect 40684 449 40724 904
rect 41452 944 41492 953
rect 40683 440 40725 449
rect 40683 400 40684 440
rect 40724 400 40725 440
rect 40683 391 40725 400
rect 41452 113 41492 904
rect 33464 20 33716 60
rect 39723 104 39765 113
rect 39723 64 39724 104
rect 39764 64 39765 104
rect 39723 55 39765 64
rect 41451 104 41493 113
rect 41451 64 41452 104
rect 41492 64 41493 104
rect 41451 55 41493 64
rect 33464 0 33544 20
<< via2 >>
rect 556 10144 596 10184
rect 1228 9136 1268 9176
rect 1804 8800 1844 8840
rect 1516 8128 1556 8168
rect 1228 7960 1268 8000
rect 1420 7792 1460 7832
rect 556 7624 596 7664
rect 1708 8464 1748 8504
rect 1612 7456 1652 7496
rect 1420 6784 1460 6824
rect 1324 6112 1364 6152
rect 1228 5944 1268 5984
rect 1036 5776 1076 5816
rect 1132 5188 1172 5228
rect 1036 3172 1076 3212
rect 1324 5020 1364 5060
rect 1228 3424 1268 3464
rect 1516 6448 1556 6488
rect 1708 6448 1748 6488
rect 1900 7120 1940 7160
rect 1708 5020 1748 5060
rect 1612 4936 1652 4976
rect 2956 9556 2996 9596
rect 2668 8632 2708 8672
rect 2860 8632 2900 8672
rect 2860 8212 2900 8252
rect 2668 8128 2708 8168
rect 3052 8548 3092 8588
rect 3148 7876 3188 7916
rect 2956 7288 2996 7328
rect 3916 9556 3956 9596
rect 3436 8884 3476 8924
rect 3628 9472 3668 9512
rect 3820 9304 3860 9344
rect 3688 9052 3728 9092
rect 3770 9052 3810 9092
rect 3852 9052 3892 9092
rect 3934 9052 3974 9092
rect 4016 9052 4056 9092
rect 4012 8884 4052 8924
rect 3340 8632 3380 8672
rect 3340 8212 3380 8252
rect 3628 8632 3668 8672
rect 5260 10564 5300 10604
rect 4928 9808 4968 9848
rect 5010 9808 5050 9848
rect 5092 9808 5132 9848
rect 5174 9808 5214 9848
rect 5256 9808 5296 9848
rect 5932 9724 5972 9764
rect 4204 9556 4244 9596
rect 4396 9472 4436 9512
rect 4204 8464 4244 8504
rect 3820 8380 3860 8420
rect 4012 7960 4052 8000
rect 3628 7876 3668 7916
rect 3436 7456 3476 7496
rect 4108 7708 4148 7748
rect 3688 7540 3728 7580
rect 3770 7540 3810 7580
rect 3852 7540 3892 7580
rect 3934 7540 3974 7580
rect 4016 7540 4056 7580
rect 3244 7120 3284 7160
rect 3436 7288 3476 7328
rect 3148 6616 3188 6656
rect 4396 8548 4436 8588
rect 4396 8380 4436 8420
rect 4300 7540 4340 7580
rect 5356 8716 5396 8756
rect 4780 8464 4820 8504
rect 4928 8296 4968 8336
rect 5010 8296 5050 8336
rect 5092 8296 5132 8336
rect 5174 8296 5214 8336
rect 5256 8296 5296 8336
rect 6028 8716 6068 8756
rect 5356 8128 5396 8168
rect 5932 8128 5972 8168
rect 4492 7708 4532 7748
rect 4396 7372 4436 7412
rect 4204 7120 4244 7160
rect 3628 6868 3668 6908
rect 2668 6448 2708 6488
rect 2956 6448 2996 6488
rect 2476 5776 2516 5816
rect 2284 5356 2324 5396
rect 1996 4600 2036 4640
rect 2188 4180 2228 4220
rect 1612 3424 1652 3464
rect 1900 3424 1940 3464
rect 1516 3004 1556 3044
rect 1132 2752 1172 2792
rect 2380 4768 2420 4808
rect 2380 4180 2420 4220
rect 3148 6448 3188 6488
rect 3340 6532 3380 6572
rect 3916 6448 3956 6488
rect 4396 7036 4436 7076
rect 4300 6448 4340 6488
rect 5164 7456 5204 7496
rect 5452 7456 5492 7496
rect 6028 7456 6068 7496
rect 5356 7288 5396 7328
rect 5164 7204 5204 7244
rect 4780 7036 4820 7076
rect 5260 7120 5300 7160
rect 5452 7120 5492 7160
rect 4876 6952 4916 6992
rect 4928 6784 4968 6824
rect 5010 6784 5050 6824
rect 5092 6784 5132 6824
rect 5174 6784 5214 6824
rect 5256 6784 5296 6824
rect 5452 6952 5492 6992
rect 4588 6448 4628 6488
rect 4492 6364 4532 6404
rect 4300 6280 4340 6320
rect 4204 6196 4244 6236
rect 3688 6028 3728 6068
rect 3770 6028 3810 6068
rect 3852 6028 3892 6068
rect 3934 6028 3974 6068
rect 4016 6028 4056 6068
rect 2668 5104 2708 5144
rect 2476 3760 2516 3800
rect 2284 3088 2324 3128
rect 3052 5608 3092 5648
rect 4108 5860 4148 5900
rect 4108 5608 4148 5648
rect 4300 5272 4340 5312
rect 3916 5104 3956 5144
rect 3052 4768 3092 4808
rect 3340 4768 3380 4808
rect 3244 4432 3284 4472
rect 2956 4012 2996 4052
rect 3148 4012 3188 4052
rect 4108 4936 4148 4976
rect 3820 4768 3860 4808
rect 3340 3760 3380 3800
rect 3688 4516 3728 4556
rect 3770 4516 3810 4556
rect 3852 4516 3892 4556
rect 3934 4516 3974 4556
rect 4016 4516 4056 4556
rect 4300 4432 4340 4472
rect 3916 4348 3956 4388
rect 3820 4096 3860 4136
rect 4876 6028 4916 6068
rect 5068 6448 5108 6488
rect 4972 5608 5012 5648
rect 5356 6448 5396 6488
rect 5356 6196 5396 6236
rect 5644 6784 5684 6824
rect 6124 7288 6164 7328
rect 5932 6952 5972 6992
rect 6412 8632 6452 8672
rect 7180 8632 7220 8672
rect 7180 8212 7220 8252
rect 7372 7960 7412 8000
rect 6604 7540 6644 7580
rect 6316 7456 6356 7496
rect 6220 7120 6260 7160
rect 5740 6616 5780 6656
rect 5548 6280 5588 6320
rect 5644 6112 5684 6152
rect 5260 5860 5300 5900
rect 5644 5860 5684 5900
rect 5740 5692 5780 5732
rect 5356 5608 5396 5648
rect 4876 5524 4916 5564
rect 5165 5524 5205 5564
rect 4928 5272 4968 5312
rect 5010 5272 5050 5312
rect 5092 5272 5132 5312
rect 5174 5272 5214 5312
rect 5256 5272 5296 5312
rect 5356 5272 5396 5312
rect 5260 5104 5300 5144
rect 5068 4936 5108 4976
rect 4492 4852 4532 4892
rect 3532 4012 3572 4052
rect 3724 3928 3764 3968
rect 3436 3424 3476 3464
rect 2956 3340 2996 3380
rect 3244 3004 3284 3044
rect 2668 1912 2708 1952
rect 2572 1072 2612 1112
rect 1324 904 1364 944
rect 3628 3676 3668 3716
rect 4012 3844 4052 3884
rect 3916 3592 3956 3632
rect 4012 3424 4052 3464
rect 3628 3340 3668 3380
rect 4108 3256 4148 3296
rect 5260 4768 5300 4808
rect 5164 4684 5204 4724
rect 5164 4432 5204 4472
rect 4684 4012 4724 4052
rect 4972 4012 5012 4052
rect 4492 3928 4532 3968
rect 4588 3676 4628 3716
rect 4396 3508 4436 3548
rect 4492 3424 4532 3464
rect 5260 3928 5300 3968
rect 4928 3760 4968 3800
rect 5010 3760 5050 3800
rect 5092 3760 5132 3800
rect 5174 3760 5214 3800
rect 5256 3760 5296 3800
rect 4780 3592 4820 3632
rect 5164 3592 5204 3632
rect 5068 3508 5108 3548
rect 4684 3424 4724 3464
rect 4588 3340 4628 3380
rect 3532 3004 3572 3044
rect 3688 3004 3728 3044
rect 3770 3004 3810 3044
rect 3852 3004 3892 3044
rect 3934 3004 3974 3044
rect 4016 3004 4056 3044
rect 4012 2836 4052 2876
rect 3340 2752 3380 2792
rect 3724 2752 3764 2792
rect 3532 2668 3572 2708
rect 3436 2584 3476 2624
rect 3820 2668 3860 2708
rect 4300 2752 4340 2792
rect 4204 2584 4244 2624
rect 4108 2500 4148 2540
rect 4972 3424 5012 3464
rect 5164 3424 5204 3464
rect 6220 6448 6260 6488
rect 6508 6952 6548 6992
rect 6028 6028 6068 6068
rect 5548 5104 5588 5144
rect 5836 5608 5876 5648
rect 6892 7288 6932 7328
rect 6796 7204 6836 7244
rect 7660 8632 7700 8672
rect 8044 8632 8084 8672
rect 7564 7708 7604 7748
rect 7564 7540 7604 7580
rect 6700 6952 6740 6992
rect 6220 5524 6260 5564
rect 5644 4012 5684 4052
rect 4972 2836 5012 2876
rect 5164 2500 5204 2540
rect 5356 2416 5396 2456
rect 4928 2248 4968 2288
rect 5010 2248 5050 2288
rect 5092 2248 5132 2288
rect 5174 2248 5214 2288
rect 5256 2248 5296 2288
rect 5260 1996 5300 2036
rect 3628 1660 3668 1700
rect 3688 1492 3728 1532
rect 3770 1492 3810 1532
rect 3852 1492 3892 1532
rect 3934 1492 3974 1532
rect 4016 1492 4056 1532
rect 4108 1156 4148 1196
rect 3436 1072 3476 1112
rect 1324 400 1364 440
rect 5548 3424 5588 3464
rect 5548 1912 5588 1952
rect 5644 1828 5684 1868
rect 5452 1492 5492 1532
rect 4300 1072 4340 1112
rect 5068 1072 5108 1112
rect 5836 4096 5876 4136
rect 5932 3760 5972 3800
rect 6604 5104 6644 5144
rect 6124 4096 6164 4136
rect 6220 3760 6260 3800
rect 5932 3172 5972 3212
rect 5932 2584 5972 2624
rect 5836 2164 5876 2204
rect 6028 2164 6068 2204
rect 5932 1828 5972 1868
rect 6124 1828 6164 1868
rect 6988 5608 7028 5648
rect 7180 6448 7220 6488
rect 7180 5613 7220 5648
rect 7180 5608 7220 5613
rect 7948 7960 7988 8000
rect 7852 7624 7892 7664
rect 8044 7540 8084 7580
rect 7756 7456 7796 7496
rect 7660 7204 7700 7244
rect 7852 7120 7892 7160
rect 7660 7036 7700 7076
rect 7564 6532 7604 6572
rect 10252 9472 10292 9512
rect 9676 8800 9716 8840
rect 8428 8548 8468 8588
rect 8332 7288 8372 7328
rect 8236 7036 8276 7076
rect 8332 6868 8372 6908
rect 8140 6784 8180 6824
rect 7660 6364 7700 6404
rect 7468 5524 7508 5564
rect 7564 5440 7604 5480
rect 7372 3928 7412 3968
rect 7084 3508 7124 3548
rect 7276 3508 7316 3548
rect 7564 2752 7604 2792
rect 7468 2668 7508 2708
rect 7180 2584 7220 2624
rect 6604 2248 6644 2288
rect 7084 1996 7124 2036
rect 7276 1996 7316 2036
rect 8812 8128 8852 8168
rect 8428 5608 8468 5648
rect 9676 8632 9716 8672
rect 10060 8212 10100 8252
rect 9100 7960 9140 8000
rect 9292 7960 9332 8000
rect 8620 7540 8660 7580
rect 8812 7540 8852 7580
rect 8812 6616 8852 6656
rect 9004 7120 9044 7160
rect 9292 7624 9332 7664
rect 9196 6952 9236 6992
rect 9292 6700 9332 6740
rect 9100 5188 9140 5228
rect 8524 4768 8564 4808
rect 8236 4348 8276 4388
rect 8428 4348 8468 4388
rect 8044 4180 8084 4220
rect 8236 4180 8276 4220
rect 7756 3928 7796 3968
rect 8044 3844 8084 3884
rect 7852 3508 7892 3548
rect 8716 4600 8756 4640
rect 8140 3424 8180 3464
rect 8620 3424 8660 3464
rect 8716 3340 8756 3380
rect 8716 3088 8756 3128
rect 9964 7708 10004 7748
rect 9676 7288 9716 7328
rect 9772 7120 9812 7160
rect 11596 10564 11636 10604
rect 11500 8800 11540 8840
rect 10540 8128 10580 8168
rect 10156 7960 10196 8000
rect 10924 7960 10964 8000
rect 11116 7960 11156 8000
rect 10540 7876 10580 7916
rect 10060 7624 10100 7664
rect 9772 6700 9812 6740
rect 9868 6532 9908 6572
rect 9580 6448 9620 6488
rect 11500 7876 11540 7916
rect 11404 7120 11444 7160
rect 11692 9640 11732 9680
rect 12172 9640 12212 9680
rect 12556 9304 12596 9344
rect 12460 8716 12500 8756
rect 12172 8464 12212 8504
rect 11884 8380 11924 8420
rect 11788 7876 11828 7916
rect 11980 7708 12020 7748
rect 11692 7120 11732 7160
rect 11596 6952 11636 6992
rect 11596 6784 11636 6824
rect 11116 6448 11156 6488
rect 11308 6196 11348 6236
rect 11212 6112 11252 6152
rect 10252 5860 10292 5900
rect 10540 5692 10580 5732
rect 10828 5692 10868 5732
rect 10252 5104 10292 5144
rect 10252 4684 10292 4724
rect 9484 4348 9524 4388
rect 9388 4096 9428 4136
rect 9964 4096 10004 4136
rect 9868 3424 9908 3464
rect 10252 3760 10292 3800
rect 10156 3592 10196 3632
rect 8812 2584 8852 2624
rect 9100 2584 9140 2624
rect 9676 2584 9716 2624
rect 8908 2248 8948 2288
rect 8332 2164 8372 2204
rect 7660 2080 7700 2120
rect 8140 2080 8180 2120
rect 7372 1912 7412 1952
rect 7852 1912 7892 1952
rect 6508 1828 6548 1868
rect 7948 1744 7988 1784
rect 6796 1660 6836 1700
rect 8332 1912 8372 1952
rect 9484 2080 9524 2120
rect 9580 1996 9620 2036
rect 8428 1828 8468 1868
rect 8140 1576 8180 1616
rect 8428 1492 8468 1532
rect 9100 1240 9140 1280
rect 6316 1072 6356 1112
rect 4492 988 4532 1028
rect 5260 988 5300 1028
rect 6988 904 7028 944
rect 4928 736 4968 776
rect 5010 736 5050 776
rect 5092 736 5132 776
rect 5174 736 5214 776
rect 5256 736 5296 776
rect 4108 64 4148 104
rect 9484 64 9524 104
rect 9868 2164 9908 2204
rect 10156 1660 10196 1700
rect 10540 4768 10580 4808
rect 10444 4012 10484 4052
rect 10636 4684 10676 4724
rect 10732 3508 10772 3548
rect 11116 5524 11156 5564
rect 10924 3592 10964 3632
rect 11116 4936 11156 4976
rect 11308 3676 11348 3716
rect 11212 3592 11252 3632
rect 11116 3508 11156 3548
rect 11212 3424 11252 3464
rect 11596 6196 11636 6236
rect 11884 7120 11924 7160
rect 11884 6868 11924 6908
rect 12364 6784 12404 6824
rect 12076 6364 12116 6404
rect 11980 6028 12020 6068
rect 11788 5440 11828 5480
rect 11692 4096 11732 4136
rect 10540 2416 10580 2456
rect 10444 2332 10484 2372
rect 10348 1828 10388 1868
rect 10636 2080 10676 2120
rect 10444 1744 10484 1784
rect 10348 1660 10388 1700
rect 10252 1576 10292 1616
rect 10156 1240 10196 1280
rect 10156 1072 10196 1112
rect 10348 904 10388 944
rect 11212 2332 11252 2372
rect 10828 1660 10868 1700
rect 10540 1576 10580 1616
rect 10540 1324 10580 1364
rect 10732 1576 10772 1616
rect 10828 1408 10868 1448
rect 10732 1156 10772 1196
rect 11020 1576 11060 1616
rect 10924 1240 10964 1280
rect 11500 2500 11540 2540
rect 11692 2500 11732 2540
rect 11980 4432 12020 4472
rect 13132 8800 13172 8840
rect 13516 8800 13556 8840
rect 13708 8800 13748 8840
rect 14668 9472 14708 9512
rect 14284 8884 14324 8924
rect 12556 8464 12596 8504
rect 13420 7876 13460 7916
rect 12844 7708 12884 7748
rect 12556 7288 12596 7328
rect 12460 5944 12500 5984
rect 12172 4936 12212 4976
rect 13132 7540 13172 7580
rect 13036 6952 13076 6992
rect 13420 7204 13460 7244
rect 12364 4768 12404 4808
rect 12268 4432 12308 4472
rect 11980 4180 12020 4220
rect 11884 4096 11924 4136
rect 12076 4096 12116 4136
rect 11980 4012 12020 4052
rect 11884 3928 11924 3968
rect 11884 3592 11924 3632
rect 12364 4096 12404 4136
rect 12460 3928 12500 3968
rect 12076 3592 12116 3632
rect 12172 3508 12212 3548
rect 11980 2668 12020 2708
rect 11788 2248 11828 2288
rect 11212 1576 11252 1616
rect 11692 1492 11732 1532
rect 11212 1408 11252 1448
rect 11404 1408 11444 1448
rect 11116 1324 11156 1364
rect 11596 1324 11636 1364
rect 11404 1240 11444 1280
rect 12172 2668 12212 2708
rect 12172 1156 12212 1196
rect 11884 736 11924 776
rect 12364 1072 12404 1112
rect 14092 8548 14132 8588
rect 13804 7960 13844 8000
rect 14476 8548 14516 8588
rect 13900 6868 13940 6908
rect 13900 6364 13940 6404
rect 13516 5608 13556 5648
rect 13612 4852 13652 4892
rect 12748 4516 12788 4556
rect 13420 4516 13460 4556
rect 12652 2416 12692 2456
rect 12652 2080 12692 2120
rect 13324 4096 13364 4136
rect 13516 4012 13556 4052
rect 12844 3592 12884 3632
rect 13420 3172 13460 3212
rect 13132 2836 13172 2876
rect 13036 2416 13076 2456
rect 12844 1996 12884 2036
rect 13036 1660 13076 1700
rect 12940 1576 12980 1616
rect 13036 820 13076 860
rect 13420 2584 13460 2624
rect 13996 4684 14036 4724
rect 14380 7204 14420 7244
rect 14188 7036 14228 7076
rect 14092 4432 14132 4472
rect 13996 4012 14036 4052
rect 14092 3928 14132 3968
rect 14284 6616 14324 6656
rect 14380 5608 14420 5648
rect 15244 9388 15284 9428
rect 15340 8800 15380 8840
rect 17932 10648 17972 10688
rect 16492 8800 16532 8840
rect 17164 8800 17204 8840
rect 15916 8632 15956 8672
rect 16684 8632 16724 8672
rect 16108 8044 16148 8084
rect 15052 7960 15092 8000
rect 16012 7876 16052 7916
rect 14764 7540 14804 7580
rect 14668 6700 14708 6740
rect 14764 6448 14804 6488
rect 16300 7372 16340 7412
rect 16300 7120 16340 7160
rect 15820 5776 15860 5816
rect 15532 5524 15572 5564
rect 14572 5440 14612 5480
rect 15436 5440 15476 5480
rect 13996 3424 14036 3464
rect 13708 2584 13748 2624
rect 13228 1660 13268 1700
rect 13324 1576 13364 1616
rect 13612 904 13652 944
rect 13996 2080 14036 2120
rect 14188 3424 14228 3464
rect 14476 3088 14516 3128
rect 14476 2668 14516 2708
rect 14860 5272 14900 5312
rect 15724 5104 15764 5144
rect 15628 4768 15668 4808
rect 15148 4096 15188 4136
rect 15052 3760 15092 3800
rect 14956 3424 14996 3464
rect 14764 2836 14804 2876
rect 14764 2416 14804 2456
rect 14668 2080 14708 2120
rect 14860 2080 14900 2120
rect 14956 1912 14996 1952
rect 14572 1744 14612 1784
rect 14476 1408 14516 1448
rect 14380 232 14420 272
rect 14860 1240 14900 1280
rect 14668 904 14708 944
rect 14668 316 14708 356
rect 16012 5608 16052 5648
rect 16012 5272 16052 5312
rect 16204 4936 16244 4976
rect 15916 4096 15956 4136
rect 16396 5608 16436 5648
rect 16588 4180 16628 4220
rect 15148 3256 15188 3296
rect 15436 3256 15476 3296
rect 15244 3088 15284 3128
rect 15244 2584 15284 2624
rect 15148 2500 15188 2540
rect 15436 2080 15476 2120
rect 16396 3424 16436 3464
rect 15628 2836 15668 2876
rect 15724 2668 15764 2708
rect 15916 2584 15956 2624
rect 16204 1912 16244 1952
rect 15628 1744 15668 1784
rect 15724 1408 15764 1448
rect 16300 1324 16340 1364
rect 15340 1240 15380 1280
rect 15148 1156 15188 1196
rect 15244 1072 15284 1112
rect 16396 1240 16436 1280
rect 15628 904 15668 944
rect 15820 652 15860 692
rect 16204 400 16244 440
rect 16012 232 16052 272
rect 16492 736 16532 776
rect 17260 7876 17300 7916
rect 17452 7876 17492 7916
rect 17356 7792 17396 7832
rect 17548 6448 17588 6488
rect 17452 6364 17492 6404
rect 17356 6280 17396 6320
rect 17164 5608 17204 5648
rect 17164 5020 17204 5060
rect 16780 4936 16820 4976
rect 16972 4852 17012 4892
rect 17068 4600 17108 4640
rect 16972 4012 17012 4052
rect 16972 3760 17012 3800
rect 16876 3676 16916 3716
rect 16684 3004 16724 3044
rect 17260 4852 17300 4892
rect 17356 4264 17396 4304
rect 16780 2668 16820 2708
rect 16972 3004 17012 3044
rect 16780 1744 16820 1784
rect 17164 2584 17204 2624
rect 17164 2080 17204 2120
rect 17356 3508 17396 3548
rect 17356 2920 17396 2960
rect 18808 9052 18848 9092
rect 18890 9052 18930 9092
rect 18972 9052 19012 9092
rect 19054 9052 19094 9092
rect 19136 9052 19176 9092
rect 19084 8800 19124 8840
rect 18220 8632 18260 8672
rect 18700 8632 18740 8672
rect 18124 8548 18164 8588
rect 17836 8212 17876 8252
rect 18220 8212 18260 8252
rect 17836 8044 17876 8084
rect 17836 7792 17876 7832
rect 17740 6700 17780 6740
rect 17932 6700 17972 6740
rect 18412 6616 18452 6656
rect 17932 6280 17972 6320
rect 17836 5860 17876 5900
rect 17644 5272 17684 5312
rect 17644 4852 17684 4892
rect 18508 6364 18548 6404
rect 18028 6112 18068 6152
rect 17836 5272 17876 5312
rect 18124 5272 18164 5312
rect 18028 3508 18068 3548
rect 17644 3256 17684 3296
rect 17932 2752 17972 2792
rect 17644 2584 17684 2624
rect 17452 2080 17492 2120
rect 17548 1912 17588 1952
rect 17740 1828 17780 1868
rect 17932 1828 17972 1868
rect 18028 1744 18068 1784
rect 17740 1576 17780 1616
rect 17932 1576 17972 1616
rect 17548 1492 17588 1532
rect 17356 1072 17396 1112
rect 17740 1156 17780 1196
rect 18412 5188 18452 5228
rect 18220 4852 18260 4892
rect 18220 4096 18260 4136
rect 18508 5020 18548 5060
rect 19372 8800 19412 8840
rect 19084 8044 19124 8084
rect 19084 7876 19124 7916
rect 19372 7876 19412 7916
rect 18808 7540 18848 7580
rect 18890 7540 18930 7580
rect 18972 7540 19012 7580
rect 19054 7540 19094 7580
rect 19136 7540 19176 7580
rect 20048 9808 20088 9848
rect 20130 9808 20170 9848
rect 20212 9808 20252 9848
rect 20294 9808 20334 9848
rect 20376 9808 20416 9848
rect 22060 8884 22100 8924
rect 20236 8464 20276 8504
rect 23692 10480 23732 10520
rect 24844 9976 24884 10016
rect 24268 9640 24308 9680
rect 24268 9472 24308 9512
rect 22444 8716 22484 8756
rect 22540 8632 22580 8672
rect 22348 8464 22388 8504
rect 20716 8380 20756 8420
rect 21484 8380 21524 8420
rect 20048 8296 20088 8336
rect 20130 8296 20170 8336
rect 20212 8296 20252 8336
rect 20294 8296 20334 8336
rect 20376 8296 20416 8336
rect 19564 7708 19604 7748
rect 19372 7120 19412 7160
rect 18988 6364 19028 6404
rect 18808 6028 18848 6068
rect 18890 6028 18930 6068
rect 18972 6028 19012 6068
rect 19054 6028 19094 6068
rect 19136 6028 19176 6068
rect 19852 7960 19892 8000
rect 19756 7624 19796 7664
rect 19852 7288 19892 7328
rect 19756 7204 19796 7244
rect 19756 7036 19796 7076
rect 20048 6784 20088 6824
rect 20130 6784 20170 6824
rect 20212 6784 20252 6824
rect 20294 6784 20334 6824
rect 20376 6784 20416 6824
rect 19564 5944 19604 5984
rect 19852 6532 19892 6572
rect 20524 6532 20564 6572
rect 19756 6448 19796 6488
rect 19660 5692 19700 5732
rect 20236 5692 20276 5732
rect 18700 5272 18740 5312
rect 18700 5104 18740 5144
rect 18220 3760 18260 3800
rect 20048 5272 20088 5312
rect 20130 5272 20170 5312
rect 20212 5272 20252 5312
rect 20294 5272 20334 5312
rect 20376 5272 20416 5312
rect 20524 5272 20564 5312
rect 21004 8044 21044 8084
rect 22540 8296 22580 8336
rect 23020 8800 23060 8840
rect 22828 8212 22868 8252
rect 22348 8044 22388 8084
rect 21580 7876 21620 7916
rect 24364 8548 24404 8588
rect 23308 8380 23348 8420
rect 23020 7960 23060 8000
rect 27148 10060 27188 10100
rect 25996 9052 26036 9092
rect 25516 8716 25556 8756
rect 25900 8632 25940 8672
rect 25324 8464 25364 8504
rect 24076 8380 24116 8420
rect 24364 8380 24404 8420
rect 23884 7708 23924 7748
rect 24268 7708 24308 7748
rect 21676 7120 21716 7160
rect 21100 7036 21140 7076
rect 21580 7036 21620 7076
rect 21004 6868 21044 6908
rect 20716 5356 20756 5396
rect 20620 5188 20660 5228
rect 19084 4852 19124 4892
rect 19276 4852 19316 4892
rect 18892 4684 18932 4724
rect 19372 4684 19412 4724
rect 18808 4516 18848 4556
rect 18890 4516 18930 4556
rect 18972 4516 19012 4556
rect 19054 4516 19094 4556
rect 19136 4516 19176 4556
rect 20044 4684 20084 4724
rect 18604 4264 18644 4304
rect 19372 4264 19412 4304
rect 19564 4264 19604 4304
rect 19948 4264 19988 4304
rect 18604 4096 18644 4136
rect 19276 4096 19316 4136
rect 18808 3004 18848 3044
rect 18890 3004 18930 3044
rect 18972 3004 19012 3044
rect 19054 3004 19094 3044
rect 19136 3004 19176 3044
rect 19564 4096 19604 4136
rect 19660 3760 19700 3800
rect 20716 4852 20756 4892
rect 20524 4096 20564 4136
rect 20044 3928 20084 3968
rect 20048 3760 20088 3800
rect 20130 3760 20170 3800
rect 20212 3760 20252 3800
rect 20294 3760 20334 3800
rect 20376 3760 20416 3800
rect 19948 3004 19988 3044
rect 20236 3004 20276 3044
rect 20140 2920 20180 2960
rect 18604 2584 18644 2624
rect 19756 2752 19796 2792
rect 19276 2668 19316 2708
rect 18508 1576 18548 1616
rect 18892 2248 18932 2288
rect 18892 2080 18932 2120
rect 19564 2584 19604 2624
rect 19756 2584 19796 2624
rect 19372 2500 19412 2540
rect 20236 2500 20276 2540
rect 21292 6616 21332 6656
rect 21196 5188 21236 5228
rect 21100 4852 21140 4892
rect 21292 4768 21332 4808
rect 21292 4516 21332 4556
rect 20908 3592 20948 3632
rect 21292 4096 21332 4136
rect 21196 3928 21236 3968
rect 21004 3424 21044 3464
rect 20908 3340 20948 3380
rect 20908 2668 20948 2708
rect 20332 2416 20372 2456
rect 19948 2332 19988 2372
rect 19852 2248 19892 2288
rect 20048 2248 20088 2288
rect 20130 2248 20170 2288
rect 20212 2248 20252 2288
rect 20294 2248 20334 2288
rect 20376 2248 20416 2288
rect 19756 2080 19796 2120
rect 19372 1912 19412 1952
rect 19276 1660 19316 1700
rect 18604 1408 18644 1448
rect 18412 904 18452 944
rect 18808 1492 18848 1532
rect 18890 1492 18930 1532
rect 18972 1492 19012 1532
rect 19054 1492 19094 1532
rect 19136 1492 19176 1532
rect 18892 1324 18932 1364
rect 18700 904 18740 944
rect 19084 1240 19124 1280
rect 18988 1072 19028 1112
rect 18988 568 19028 608
rect 19276 904 19316 944
rect 20428 2080 20468 2120
rect 20236 1828 20276 1868
rect 19660 1660 19700 1700
rect 19660 1324 19700 1364
rect 19660 820 19700 860
rect 19852 568 19892 608
rect 20044 1408 20084 1448
rect 20140 1156 20180 1196
rect 20332 1072 20372 1112
rect 20048 736 20088 776
rect 20130 736 20170 776
rect 20212 736 20252 776
rect 20294 736 20334 776
rect 20376 736 20416 776
rect 20716 2416 20756 2456
rect 20716 1912 20756 1952
rect 20908 1828 20948 1868
rect 20812 1660 20852 1700
rect 20812 1324 20852 1364
rect 20716 1240 20756 1280
rect 20620 736 20660 776
rect 20236 148 20276 188
rect 21580 6616 21620 6656
rect 22060 6700 22100 6740
rect 22636 6448 22676 6488
rect 22156 6364 22196 6404
rect 22060 5692 22100 5732
rect 21676 5608 21716 5648
rect 22156 5188 22196 5228
rect 21484 4768 21524 4808
rect 21388 3760 21428 3800
rect 21292 3592 21332 3632
rect 21676 4096 21716 4136
rect 22348 4348 22388 4388
rect 21580 4012 21620 4052
rect 21196 1828 21236 1868
rect 21196 1240 21236 1280
rect 21484 3424 21524 3464
rect 21484 1996 21524 2036
rect 21388 1912 21428 1952
rect 21100 1156 21140 1196
rect 21868 1324 21908 1364
rect 21772 1156 21812 1196
rect 21676 988 21716 1028
rect 21964 1072 22004 1112
rect 22156 1324 22196 1364
rect 22156 988 22196 1028
rect 22636 3592 22676 3632
rect 22444 3424 22484 3464
rect 22636 3424 22676 3464
rect 22444 3256 22484 3296
rect 22540 316 22580 356
rect 22924 5272 22964 5312
rect 23308 5272 23348 5312
rect 23500 5104 23540 5144
rect 23020 5020 23060 5060
rect 22924 4936 22964 4976
rect 24172 7120 24212 7160
rect 24172 6616 24212 6656
rect 24940 8044 24980 8084
rect 24556 7876 24596 7916
rect 24460 6028 24500 6068
rect 23980 5104 24020 5144
rect 23980 4936 24020 4976
rect 23884 4852 23924 4892
rect 23692 4516 23732 4556
rect 23596 4348 23636 4388
rect 22828 3592 22868 3632
rect 22924 1156 22964 1196
rect 24076 4852 24116 4892
rect 24268 4768 24308 4808
rect 24172 4600 24212 4640
rect 24076 4432 24116 4472
rect 23980 4264 24020 4304
rect 24076 4180 24116 4220
rect 23404 3760 23444 3800
rect 23308 3508 23348 3548
rect 23500 3508 23540 3548
rect 23212 3424 23252 3464
rect 23116 3004 23156 3044
rect 23212 2752 23252 2792
rect 23692 3508 23732 3548
rect 23596 2920 23636 2960
rect 23500 2584 23540 2624
rect 23116 904 23156 944
rect 23404 2080 23444 2120
rect 23308 1156 23348 1196
rect 23500 1660 23540 1700
rect 23500 1240 23540 1280
rect 23980 3844 24020 3884
rect 23884 3760 23924 3800
rect 23788 2920 23828 2960
rect 23884 2248 23924 2288
rect 23692 1660 23732 1700
rect 23884 1660 23924 1700
rect 23692 1240 23732 1280
rect 23692 904 23732 944
rect 24460 4852 24500 4892
rect 24364 4684 24404 4724
rect 24460 3760 24500 3800
rect 24460 3424 24500 3464
rect 24172 3340 24212 3380
rect 24076 3004 24116 3044
rect 24172 2920 24212 2960
rect 24460 2584 24500 2624
rect 24076 1240 24116 1280
rect 23980 316 24020 356
rect 24268 1240 24308 1280
rect 24172 568 24212 608
rect 26572 8632 26612 8672
rect 26380 8044 26420 8084
rect 25900 7960 25940 8000
rect 25420 7120 25460 7160
rect 25612 7120 25652 7160
rect 25228 6868 25268 6908
rect 26380 7708 26420 7748
rect 26284 7540 26324 7580
rect 25900 6952 25940 6992
rect 25996 6700 26036 6740
rect 25324 6364 25364 6404
rect 25228 5776 25268 5816
rect 24748 5356 24788 5396
rect 24844 4852 24884 4892
rect 24940 4768 24980 4808
rect 25132 4180 25172 4220
rect 24748 3676 24788 3716
rect 24652 3340 24692 3380
rect 24748 2752 24788 2792
rect 25132 2752 25172 2792
rect 24556 2248 24596 2288
rect 24556 904 24596 944
rect 24940 2248 24980 2288
rect 25324 3508 25364 3548
rect 25612 5104 25652 5144
rect 25516 3592 25556 3632
rect 25900 4936 25940 4976
rect 25708 4852 25748 4892
rect 25708 4180 25748 4220
rect 25708 3676 25748 3716
rect 25324 1912 25364 1952
rect 25132 1240 25172 1280
rect 24748 1156 24788 1196
rect 24844 904 24884 944
rect 25036 820 25076 860
rect 25324 1660 25364 1700
rect 25228 736 25268 776
rect 26284 6952 26324 6992
rect 26284 6700 26324 6740
rect 27532 8632 27572 8672
rect 27148 7876 27188 7916
rect 29260 10648 29300 10688
rect 28300 8884 28340 8924
rect 28780 8548 28820 8588
rect 28684 7960 28724 8000
rect 27724 7876 27764 7916
rect 28396 7876 28436 7916
rect 27052 7708 27092 7748
rect 26860 7540 26900 7580
rect 27724 7372 27764 7412
rect 26476 7120 26516 7160
rect 26476 5860 26516 5900
rect 26476 5692 26516 5732
rect 26380 4936 26420 4976
rect 26092 3928 26132 3968
rect 26092 3760 26132 3800
rect 25996 3592 26036 3632
rect 25996 3424 26036 3464
rect 25804 3004 25844 3044
rect 25996 3004 26036 3044
rect 25708 2920 25748 2960
rect 26284 3172 26324 3212
rect 26188 2668 26228 2708
rect 25612 1324 25652 1364
rect 25708 1156 25748 1196
rect 25612 232 25652 272
rect 26092 2164 26132 2204
rect 26092 1156 26132 1196
rect 27724 7120 27764 7160
rect 28300 6448 28340 6488
rect 28012 6364 28052 6404
rect 26956 6280 26996 6320
rect 26860 5524 26900 5564
rect 26572 3676 26612 3716
rect 26668 3508 26708 3548
rect 26860 3340 26900 3380
rect 26476 3004 26516 3044
rect 27052 5020 27092 5060
rect 27148 3004 27188 3044
rect 26380 2164 26420 2204
rect 26284 1324 26324 1364
rect 26764 1576 26804 1616
rect 26668 820 26708 860
rect 26572 736 26612 776
rect 26860 1324 26900 1364
rect 26956 1240 26996 1280
rect 27052 652 27092 692
rect 27052 484 27092 524
rect 27244 2500 27284 2540
rect 27340 1912 27380 1952
rect 27244 1828 27284 1868
rect 27724 5440 27764 5480
rect 27532 4180 27572 4220
rect 27628 4012 27668 4052
rect 27820 4180 27860 4220
rect 28012 4096 28052 4136
rect 28204 5188 28244 5228
rect 28300 4600 28340 4640
rect 27532 3676 27572 3716
rect 27628 3340 27668 3380
rect 28108 3256 28148 3296
rect 27532 2752 27572 2792
rect 28780 7456 28820 7496
rect 28876 7204 28916 7244
rect 29740 10480 29780 10520
rect 29452 9892 29492 9932
rect 32428 10060 32468 10100
rect 32044 9976 32084 10016
rect 29836 9472 29876 9512
rect 29164 8044 29204 8084
rect 29260 7876 29300 7916
rect 29164 7540 29204 7580
rect 28972 7120 29012 7160
rect 28972 6700 29012 6740
rect 28780 5776 28820 5816
rect 28396 4432 28436 4472
rect 29260 7288 29300 7328
rect 29164 7036 29204 7076
rect 29740 6532 29780 6572
rect 29548 6364 29588 6404
rect 29548 5104 29588 5144
rect 28780 3592 28820 3632
rect 28588 3424 28628 3464
rect 28300 3256 28340 3296
rect 29068 4936 29108 4976
rect 29068 3928 29108 3968
rect 28972 2752 29012 2792
rect 28780 2584 28820 2624
rect 27916 2416 27956 2456
rect 27820 2332 27860 2372
rect 27724 1912 27764 1952
rect 27340 1156 27380 1196
rect 27436 904 27476 944
rect 28012 2332 28052 2372
rect 28588 2416 28628 2456
rect 28396 2080 28436 2120
rect 28108 1996 28148 2036
rect 28012 1492 28052 1532
rect 28300 1744 28340 1784
rect 28396 1492 28436 1532
rect 28204 1324 28244 1364
rect 28492 988 28532 1028
rect 27916 904 27956 944
rect 28780 2332 28820 2372
rect 28876 2164 28916 2204
rect 28684 904 28724 944
rect 28108 400 28148 440
rect 28300 64 28340 104
rect 28684 316 28724 356
rect 28972 1912 29012 1952
rect 29356 3340 29396 3380
rect 29356 3004 29396 3044
rect 29164 2752 29204 2792
rect 29260 1947 29300 1952
rect 29260 1912 29300 1947
rect 29164 1072 29204 1112
rect 29644 2584 29684 2624
rect 30604 9052 30644 9092
rect 29452 1828 29492 1868
rect 29356 988 29396 1028
rect 29260 904 29300 944
rect 30028 8632 30068 8672
rect 31660 9472 31700 9512
rect 32236 9388 32276 9428
rect 31756 8884 31796 8924
rect 30892 8800 30932 8840
rect 32140 8800 32180 8840
rect 32812 9892 32852 9932
rect 32620 8968 32660 9008
rect 31084 8464 31124 8504
rect 30124 7120 30164 7160
rect 30028 6700 30068 6740
rect 30220 6532 30260 6572
rect 30124 6112 30164 6152
rect 30124 5440 30164 5480
rect 30124 5272 30164 5312
rect 30028 3256 30068 3296
rect 29932 2248 29972 2288
rect 29836 1996 29876 2036
rect 30316 4516 30356 4556
rect 30220 2752 30260 2792
rect 30124 2584 30164 2624
rect 30220 1828 30260 1868
rect 30028 1492 30068 1532
rect 30028 988 30068 1028
rect 30508 6532 30548 6572
rect 31564 8464 31604 8504
rect 31756 8044 31796 8084
rect 31564 7876 31604 7916
rect 31660 7540 31700 7580
rect 31372 7120 31412 7160
rect 31660 7036 31700 7076
rect 31468 6448 31508 6488
rect 31276 6364 31316 6404
rect 31564 5524 31604 5564
rect 30412 3844 30452 3884
rect 30412 3088 30452 3128
rect 30412 2248 30452 2288
rect 30796 3676 30836 3716
rect 30796 3004 30836 3044
rect 30988 3844 31028 3884
rect 30892 2500 30932 2540
rect 31084 2500 31124 2540
rect 30604 1828 30644 1868
rect 30508 988 30548 1028
rect 30988 1828 31028 1868
rect 31276 3676 31316 3716
rect 31276 2080 31316 2120
rect 31564 3844 31604 3884
rect 31468 3508 31508 3548
rect 31564 1912 31604 1952
rect 31372 1324 31412 1364
rect 32140 7876 32180 7916
rect 31948 6448 31988 6488
rect 31756 6364 31796 6404
rect 31756 6196 31796 6236
rect 31948 5608 31988 5648
rect 31852 5524 31892 5564
rect 32140 6196 32180 6236
rect 32140 5608 32180 5648
rect 31948 4768 31988 4808
rect 31756 3760 31796 3800
rect 31756 3508 31796 3548
rect 31852 3424 31892 3464
rect 31852 2584 31892 2624
rect 30700 820 30740 860
rect 30796 736 30836 776
rect 31756 1744 31796 1784
rect 30988 820 31028 860
rect 30892 148 30932 188
rect 31180 736 31220 776
rect 31660 1240 31700 1280
rect 32044 3760 32084 3800
rect 32044 3592 32084 3632
rect 32524 7876 32564 7916
rect 32524 7708 32564 7748
rect 32428 7540 32468 7580
rect 32332 6364 32372 6404
rect 32620 7540 32660 7580
rect 32524 6700 32564 6740
rect 32524 5188 32564 5228
rect 32428 4852 32468 4892
rect 32236 4768 32276 4808
rect 32524 4768 32564 4808
rect 32428 3844 32468 3884
rect 32236 2584 32276 2624
rect 32428 3172 32468 3212
rect 33004 8044 33044 8084
rect 33100 7876 33140 7916
rect 33100 7540 33140 7580
rect 32908 7120 32948 7160
rect 32812 6364 32852 6404
rect 32908 5692 32948 5732
rect 33100 5692 33140 5732
rect 34252 9220 34292 9260
rect 33928 9052 33968 9092
rect 34010 9052 34050 9092
rect 34092 9052 34132 9092
rect 34174 9052 34214 9092
rect 34256 9052 34296 9092
rect 33292 8128 33332 8168
rect 34540 9472 34580 9512
rect 34348 8128 34388 8168
rect 33676 8044 33716 8084
rect 33580 7960 33620 8000
rect 33292 7876 33332 7916
rect 33388 7792 33428 7832
rect 33388 6196 33428 6236
rect 33292 5692 33332 5732
rect 33196 5608 33236 5648
rect 32812 4180 32852 4220
rect 34828 9136 34868 9176
rect 35168 9808 35208 9848
rect 35250 9808 35290 9848
rect 35332 9808 35372 9848
rect 35414 9808 35454 9848
rect 35496 9808 35536 9848
rect 35212 9472 35252 9512
rect 36172 9472 36212 9512
rect 35884 9052 35924 9092
rect 36556 9556 36596 9596
rect 36844 9472 36884 9512
rect 36844 9052 36884 9092
rect 35020 8800 35060 8840
rect 36172 8800 36212 8840
rect 35168 8296 35208 8336
rect 35250 8296 35290 8336
rect 35332 8296 35372 8336
rect 35414 8296 35454 8336
rect 35496 8296 35536 8336
rect 35308 7960 35348 8000
rect 33928 7540 33968 7580
rect 34010 7540 34050 7580
rect 34092 7540 34132 7580
rect 34174 7540 34214 7580
rect 34256 7540 34296 7580
rect 33772 7120 33812 7160
rect 34636 7120 34676 7160
rect 34348 7036 34388 7076
rect 33964 6196 34004 6236
rect 33928 6028 33968 6068
rect 34010 6028 34050 6068
rect 34092 6028 34132 6068
rect 34174 6028 34214 6068
rect 34256 6028 34296 6068
rect 33772 5608 33812 5648
rect 33292 5272 33332 5312
rect 33676 5272 33716 5312
rect 32812 3844 32852 3884
rect 32524 2584 32564 2624
rect 32332 2332 32372 2372
rect 32044 2080 32084 2120
rect 33100 3676 33140 3716
rect 33004 2836 33044 2876
rect 32908 2752 32948 2792
rect 33580 5188 33620 5228
rect 33676 4180 33716 4220
rect 33580 4096 33620 4136
rect 32524 1828 32564 1868
rect 32332 1744 32372 1784
rect 32140 1324 32180 1364
rect 32044 1240 32084 1280
rect 31660 820 31700 860
rect 31948 568 31988 608
rect 32428 1660 32468 1700
rect 32332 652 32372 692
rect 32620 1660 32660 1700
rect 32620 1324 32660 1364
rect 33484 3508 33524 3548
rect 33484 2836 33524 2876
rect 33292 2752 33332 2792
rect 33004 1912 33044 1952
rect 32908 736 32948 776
rect 32716 568 32756 608
rect 32716 148 32756 188
rect 33292 1996 33332 2036
rect 33196 1240 33236 1280
rect 33388 1912 33428 1952
rect 33580 2332 33620 2372
rect 33484 1072 33524 1112
rect 33292 736 33332 776
rect 34540 5692 34580 5732
rect 34156 4936 34196 4976
rect 34444 4768 34484 4808
rect 33928 4516 33968 4556
rect 34010 4516 34050 4556
rect 34092 4516 34132 4556
rect 34174 4516 34214 4556
rect 34256 4516 34296 4556
rect 34348 4348 34388 4388
rect 33928 3004 33968 3044
rect 34010 3004 34050 3044
rect 34092 3004 34132 3044
rect 34174 3004 34214 3044
rect 34256 3004 34296 3044
rect 34444 3760 34484 3800
rect 34444 3424 34484 3464
rect 34636 3508 34676 3548
rect 34540 3172 34580 3212
rect 34348 2836 34388 2876
rect 34252 2752 34292 2792
rect 34540 2752 34580 2792
rect 33772 1828 33812 1868
rect 35168 6784 35208 6824
rect 35250 6784 35290 6824
rect 35332 6784 35372 6824
rect 35414 6784 35454 6824
rect 35496 6784 35536 6824
rect 35020 5944 35060 5984
rect 35404 5944 35444 5984
rect 34828 5860 34868 5900
rect 35404 5608 35444 5648
rect 35692 6868 35732 6908
rect 35884 6868 35924 6908
rect 36172 7708 36212 7748
rect 36076 6112 36116 6152
rect 35980 5776 36020 5816
rect 35168 5272 35208 5312
rect 35250 5272 35290 5312
rect 35332 5272 35372 5312
rect 35414 5272 35454 5312
rect 35496 5272 35536 5312
rect 35788 5356 35828 5396
rect 35788 5104 35828 5144
rect 35020 4432 35060 4472
rect 34828 4096 34868 4136
rect 35596 4852 35636 4892
rect 35404 4180 35444 4220
rect 35168 3760 35208 3800
rect 35250 3760 35290 3800
rect 35332 3760 35372 3800
rect 35414 3760 35454 3800
rect 35496 3760 35536 3800
rect 35212 3004 35252 3044
rect 34732 2584 34772 2624
rect 35212 2584 35252 2624
rect 35692 3676 35732 3716
rect 36460 7708 36500 7748
rect 36364 6280 36404 6320
rect 36556 6364 36596 6404
rect 36844 7876 36884 7916
rect 37324 7960 37364 8000
rect 37036 7372 37076 7412
rect 36844 6364 36884 6404
rect 36748 5524 36788 5564
rect 35884 4180 35924 4220
rect 36268 4096 36308 4136
rect 35788 3424 35828 3464
rect 35884 3340 35924 3380
rect 35168 2248 35208 2288
rect 35250 2248 35290 2288
rect 35332 2248 35372 2288
rect 35414 2248 35454 2288
rect 35496 2248 35536 2288
rect 33928 1492 33968 1532
rect 34010 1492 34050 1532
rect 34092 1492 34132 1532
rect 34174 1492 34214 1532
rect 34256 1492 34296 1532
rect 35404 1912 35444 1952
rect 34828 1240 34868 1280
rect 35308 1240 35348 1280
rect 34636 1072 34676 1112
rect 35168 736 35208 776
rect 35250 736 35290 776
rect 35332 736 35372 776
rect 35414 736 35454 776
rect 35496 736 35536 776
rect 35020 652 35060 692
rect 35884 2668 35924 2708
rect 35788 2248 35828 2288
rect 36076 2584 36116 2624
rect 36940 4096 36980 4136
rect 37132 4096 37172 4136
rect 36364 3088 36404 3128
rect 36364 2752 36404 2792
rect 35692 1912 35732 1952
rect 36652 3928 36692 3968
rect 36748 3592 36788 3632
rect 36556 3340 36596 3380
rect 36556 2920 36596 2960
rect 36748 2752 36788 2792
rect 36556 2668 36596 2708
rect 36460 2584 36500 2624
rect 35884 1828 35924 1868
rect 36172 1828 36212 1868
rect 36460 1240 36500 1280
rect 36844 1240 36884 1280
rect 36268 1072 36308 1112
rect 37708 3459 37748 3464
rect 37708 3424 37748 3459
rect 37324 3340 37364 3380
rect 40012 9808 40052 9848
rect 40684 10480 40724 10520
rect 41452 10144 41492 10184
rect 41260 9640 41300 9680
rect 41068 9472 41108 9512
rect 38476 8716 38516 8756
rect 37900 7876 37940 7916
rect 38092 7960 38132 8000
rect 38092 7624 38132 7664
rect 38572 8044 38612 8084
rect 37996 6448 38036 6488
rect 37900 6364 37940 6404
rect 38092 6364 38132 6404
rect 38188 4012 38228 4052
rect 38572 7120 38612 7160
rect 38860 7120 38900 7160
rect 38476 4096 38516 4136
rect 38380 4012 38420 4052
rect 38284 3928 38324 3968
rect 38092 3676 38132 3716
rect 38284 3676 38324 3716
rect 37132 3004 37172 3044
rect 37612 2589 37652 2624
rect 37612 2584 37652 2589
rect 37036 2248 37076 2288
rect 38092 3256 38132 3296
rect 37900 1996 37940 2036
rect 36268 904 36308 944
rect 36940 904 36980 944
rect 36652 652 36692 692
rect 35596 400 35636 440
rect 37996 1576 38036 1616
rect 38668 3928 38708 3968
rect 38860 4264 38900 4304
rect 38860 4012 38900 4052
rect 39820 8716 39860 8756
rect 39244 6364 39284 6404
rect 39628 6280 39668 6320
rect 39052 5776 39092 5816
rect 39436 5608 39476 5648
rect 39148 4096 39188 4136
rect 38764 2080 38804 2120
rect 38956 2500 38996 2540
rect 40876 9388 40916 9428
rect 41452 9052 41492 9092
rect 41068 8800 41108 8840
rect 40492 8548 40532 8588
rect 40876 8380 40916 8420
rect 41452 8464 41492 8504
rect 41260 8212 41300 8252
rect 40684 8128 40724 8168
rect 40492 7876 40532 7916
rect 40684 7456 40724 7496
rect 40492 7372 40532 7412
rect 40684 6784 40724 6824
rect 41260 7876 41300 7916
rect 41068 7792 41108 7832
rect 40876 6700 40916 6740
rect 40780 6448 40820 6488
rect 40204 5188 40244 5228
rect 40684 5776 40724 5816
rect 40492 5692 40532 5732
rect 40876 5440 40916 5480
rect 40396 5104 40436 5144
rect 40684 5104 40724 5144
rect 39820 4348 39860 4388
rect 39532 3508 39572 3548
rect 40396 4936 40436 4976
rect 40300 4348 40340 4388
rect 40876 4852 40916 4892
rect 40492 4600 40532 4640
rect 40876 4180 40916 4220
rect 40108 4096 40148 4136
rect 40684 4096 40724 4136
rect 40108 3760 40148 3800
rect 40588 3760 40628 3800
rect 40492 3592 40532 3632
rect 39052 2332 39092 2372
rect 38956 2080 38996 2120
rect 39724 2164 39764 2204
rect 38956 1408 38996 1448
rect 38572 1156 38612 1196
rect 39532 1156 39572 1196
rect 39724 1072 39764 1112
rect 38284 904 38324 944
rect 37900 820 37940 860
rect 37516 316 37556 356
rect 34444 232 34484 272
rect 41068 7120 41108 7160
rect 41068 6448 41108 6488
rect 41164 6364 41204 6404
rect 41068 6112 41108 6152
rect 41068 5440 41108 5480
rect 41068 4432 41108 4472
rect 40972 3508 41012 3548
rect 41068 3424 41108 3464
rect 40876 3340 40916 3380
rect 41452 4768 41492 4808
rect 41260 4684 41300 4724
rect 41260 4012 41300 4052
rect 41452 3760 41492 3800
rect 40684 3172 40724 3212
rect 41260 3004 41300 3044
rect 40876 2836 40916 2876
rect 41068 2752 41108 2792
rect 41452 2416 41492 2456
rect 41548 2080 41588 2120
rect 41068 1744 41108 1784
rect 40876 1240 40916 1280
rect 41644 1240 41684 1280
rect 40492 1156 40532 1196
rect 40300 1072 40340 1112
rect 41260 1156 41300 1196
rect 40876 988 40916 1028
rect 40108 820 40148 860
rect 40300 736 40340 776
rect 40684 400 40724 440
rect 39724 64 39764 104
rect 41452 64 41492 104
<< metal3 >>
rect 17923 10648 17932 10688
rect 17972 10648 29260 10688
rect 29300 10648 29309 10688
rect 5251 10564 5260 10604
rect 5300 10564 11596 10604
rect 11636 10564 11645 10604
rect 0 10520 80 10540
rect 259 10520 317 10521
rect 42928 10520 43008 10540
rect 0 10480 268 10520
rect 308 10480 317 10520
rect 23683 10480 23692 10520
rect 23732 10480 29740 10520
rect 29780 10480 29789 10520
rect 40675 10480 40684 10520
rect 40724 10480 43008 10520
rect 0 10460 80 10480
rect 259 10479 317 10480
rect 42928 10460 43008 10480
rect 0 10184 80 10204
rect 42928 10184 43008 10204
rect 0 10144 556 10184
rect 596 10144 605 10184
rect 41443 10144 41452 10184
rect 41492 10144 43008 10184
rect 0 10124 80 10144
rect 42928 10124 43008 10144
rect 27139 10060 27148 10100
rect 27188 10060 32428 10100
rect 32468 10060 32477 10100
rect 24835 9976 24844 10016
rect 24884 9976 32044 10016
rect 32084 9976 32093 10016
rect 29443 9892 29452 9932
rect 29492 9892 32812 9932
rect 32852 9892 32861 9932
rect 0 9848 80 9868
rect 42928 9848 43008 9868
rect 0 9808 2540 9848
rect 4919 9808 4928 9848
rect 4968 9808 5010 9848
rect 5050 9808 5092 9848
rect 5132 9808 5174 9848
rect 5214 9808 5256 9848
rect 5296 9808 5305 9848
rect 20039 9808 20048 9848
rect 20088 9808 20130 9848
rect 20170 9808 20212 9848
rect 20252 9808 20294 9848
rect 20334 9808 20376 9848
rect 20416 9808 20425 9848
rect 35159 9808 35168 9848
rect 35208 9808 35250 9848
rect 35290 9808 35332 9848
rect 35372 9808 35414 9848
rect 35454 9808 35496 9848
rect 35536 9808 35545 9848
rect 40003 9808 40012 9848
rect 40052 9808 43008 9848
rect 0 9788 80 9808
rect 2500 9764 2540 9808
rect 42928 9788 43008 9808
rect 2500 9724 5932 9764
rect 5972 9724 5981 9764
rect 11683 9640 11692 9680
rect 11732 9640 12172 9680
rect 12212 9640 12221 9680
rect 24259 9640 24268 9680
rect 24308 9640 41260 9680
rect 41300 9640 41309 9680
rect 2947 9556 2956 9596
rect 2996 9556 3916 9596
rect 3956 9556 4204 9596
rect 4244 9556 4253 9596
rect 31660 9556 36556 9596
rect 36596 9556 36605 9596
rect 0 9512 80 9532
rect 1219 9512 1277 9513
rect 10051 9512 10109 9513
rect 31660 9512 31700 9556
rect 42928 9512 43008 9532
rect 0 9472 1228 9512
rect 1268 9472 1277 9512
rect 3619 9472 3628 9512
rect 3668 9472 4396 9512
rect 4436 9472 4445 9512
rect 10051 9472 10060 9512
rect 10100 9472 10252 9512
rect 10292 9472 10301 9512
rect 14659 9472 14668 9512
rect 14708 9472 24268 9512
rect 24308 9472 24317 9512
rect 29827 9472 29836 9512
rect 29876 9472 31660 9512
rect 31700 9472 31709 9512
rect 34531 9472 34540 9512
rect 34580 9472 35212 9512
rect 35252 9472 35261 9512
rect 36163 9472 36172 9512
rect 36212 9472 36844 9512
rect 36884 9472 36893 9512
rect 41059 9472 41068 9512
rect 41108 9472 43008 9512
rect 0 9452 80 9472
rect 1219 9471 1277 9472
rect 10051 9471 10109 9472
rect 42928 9452 43008 9472
rect 15235 9428 15293 9429
rect 15150 9388 15244 9428
rect 15284 9388 15293 9428
rect 15235 9387 15293 9388
rect 30787 9428 30845 9429
rect 30787 9388 30796 9428
rect 30836 9388 32236 9428
rect 32276 9388 32285 9428
rect 37780 9388 40876 9428
rect 40916 9388 40925 9428
rect 30787 9387 30845 9388
rect 4291 9344 4349 9345
rect 37780 9344 37820 9388
rect 3811 9304 3820 9344
rect 3860 9304 4300 9344
rect 4340 9304 4349 9344
rect 12547 9304 12556 9344
rect 12596 9304 37820 9344
rect 4291 9303 4349 9304
rect 34243 9220 34252 9260
rect 34292 9220 34868 9260
rect 0 9176 80 9196
rect 34828 9176 34868 9220
rect 42928 9176 43008 9196
rect 0 9136 1228 9176
rect 1268 9136 1277 9176
rect 34819 9136 34828 9176
rect 34868 9136 34877 9176
rect 41452 9136 43008 9176
rect 0 9116 80 9136
rect 41452 9092 41492 9136
rect 42928 9116 43008 9136
rect 3679 9052 3688 9092
rect 3728 9052 3770 9092
rect 3810 9052 3852 9092
rect 3892 9052 3934 9092
rect 3974 9052 4016 9092
rect 4056 9052 4065 9092
rect 18799 9052 18808 9092
rect 18848 9052 18890 9092
rect 18930 9052 18972 9092
rect 19012 9052 19054 9092
rect 19094 9052 19136 9092
rect 19176 9052 19185 9092
rect 25987 9052 25996 9092
rect 26036 9052 30604 9092
rect 30644 9052 30653 9092
rect 33919 9052 33928 9092
rect 33968 9052 34010 9092
rect 34050 9052 34092 9092
rect 34132 9052 34174 9092
rect 34214 9052 34256 9092
rect 34296 9052 34305 9092
rect 35875 9052 35884 9092
rect 35924 9052 36844 9092
rect 36884 9052 36893 9092
rect 41443 9052 41452 9092
rect 41492 9052 41501 9092
rect 31171 9008 31229 9009
rect 31171 8968 31180 9008
rect 31220 8968 32620 9008
rect 32660 8968 32669 9008
rect 31171 8967 31229 8968
rect 3427 8884 3436 8924
rect 3476 8884 4012 8924
rect 4052 8884 4061 8924
rect 14275 8884 14284 8924
rect 14324 8884 22060 8924
rect 22100 8884 22109 8924
rect 28291 8884 28300 8924
rect 28340 8884 31756 8924
rect 31796 8884 31805 8924
rect 0 8840 80 8860
rect 42928 8840 43008 8860
rect 0 8800 1804 8840
rect 1844 8800 9676 8840
rect 9716 8800 9725 8840
rect 11491 8800 11500 8840
rect 11540 8800 13132 8840
rect 13172 8800 13516 8840
rect 13556 8800 13708 8840
rect 13748 8800 15340 8840
rect 15380 8800 16492 8840
rect 16532 8800 17164 8840
rect 17204 8800 17213 8840
rect 19075 8800 19084 8840
rect 19124 8800 19372 8840
rect 19412 8800 19421 8840
rect 20140 8800 23020 8840
rect 23060 8800 23069 8840
rect 30883 8800 30892 8840
rect 30932 8800 32140 8840
rect 32180 8800 32189 8840
rect 35011 8800 35020 8840
rect 35060 8800 36172 8840
rect 36212 8800 36221 8840
rect 41059 8800 41068 8840
rect 41108 8800 43008 8840
rect 0 8780 80 8800
rect 12451 8756 12509 8757
rect 5347 8716 5356 8756
rect 5396 8716 6028 8756
rect 6068 8716 7220 8756
rect 12366 8716 12460 8756
rect 12500 8716 12509 8756
rect 6403 8672 6461 8673
rect 7180 8672 7220 8716
rect 12451 8715 12509 8716
rect 8035 8672 8093 8673
rect 15907 8672 15965 8673
rect 20140 8672 20180 8800
rect 42928 8780 43008 8800
rect 39811 8756 39869 8757
rect 22435 8716 22444 8756
rect 22484 8716 25516 8756
rect 25556 8716 38476 8756
rect 38516 8716 38525 8756
rect 39726 8716 39820 8756
rect 39860 8716 39869 8756
rect 2659 8632 2668 8672
rect 2708 8632 2860 8672
rect 2900 8632 2909 8672
rect 3331 8632 3340 8672
rect 3380 8632 3628 8672
rect 3668 8632 3677 8672
rect 6318 8632 6412 8672
rect 6452 8632 6461 8672
rect 7171 8632 7180 8672
rect 7220 8632 7660 8672
rect 7700 8632 7709 8672
rect 7950 8632 8044 8672
rect 8084 8632 8093 8672
rect 9667 8632 9676 8672
rect 9716 8632 15916 8672
rect 15956 8632 15965 8672
rect 16675 8632 16684 8672
rect 16724 8632 18220 8672
rect 18260 8632 18269 8672
rect 18691 8632 18700 8672
rect 18740 8632 20180 8672
rect 6403 8631 6461 8632
rect 8035 8631 8093 8632
rect 15907 8631 15965 8632
rect 6412 8588 6452 8631
rect 14083 8588 14141 8589
rect 22444 8588 22484 8716
rect 39811 8715 39869 8716
rect 30019 8672 30077 8673
rect 22531 8632 22540 8672
rect 22580 8632 25900 8672
rect 25940 8632 25949 8672
rect 26563 8632 26572 8672
rect 26612 8632 27532 8672
rect 27572 8632 27581 8672
rect 29934 8632 30028 8672
rect 30068 8632 30077 8672
rect 30019 8631 30077 8632
rect 24355 8588 24413 8589
rect 3043 8548 3052 8588
rect 3092 8548 4396 8588
rect 4436 8548 4445 8588
rect 6412 8548 8428 8588
rect 8468 8548 8477 8588
rect 13998 8548 14092 8588
rect 14132 8548 14141 8588
rect 14467 8548 14476 8588
rect 14516 8548 18124 8588
rect 18164 8548 22484 8588
rect 24270 8548 24364 8588
rect 24404 8548 24413 8588
rect 0 8504 80 8524
rect 4204 8504 4244 8548
rect 14083 8547 14141 8548
rect 24355 8547 24413 8548
rect 27811 8588 27869 8589
rect 27811 8548 27820 8588
rect 27860 8548 28780 8588
rect 28820 8548 40492 8588
rect 40532 8548 40541 8588
rect 27811 8547 27869 8548
rect 4771 8504 4829 8505
rect 22339 8504 22397 8505
rect 23779 8504 23837 8505
rect 25411 8504 25469 8505
rect 42928 8504 43008 8524
rect 0 8464 1708 8504
rect 1748 8464 1757 8504
rect 4195 8464 4204 8504
rect 4244 8464 4284 8504
rect 4686 8464 4780 8504
rect 4820 8464 12172 8504
rect 12212 8464 12556 8504
rect 12596 8464 12605 8504
rect 20227 8464 20236 8504
rect 20276 8464 20316 8504
rect 22254 8464 22348 8504
rect 22388 8464 23788 8504
rect 23828 8464 23837 8504
rect 0 8444 80 8464
rect 4771 8463 4829 8464
rect 20236 8420 20276 8464
rect 22339 8463 22397 8464
rect 23779 8463 23837 8464
rect 24076 8464 25324 8504
rect 25364 8464 25420 8504
rect 25460 8464 25488 8504
rect 31075 8464 31084 8504
rect 31124 8464 31564 8504
rect 31604 8464 31613 8504
rect 41443 8464 41452 8504
rect 41492 8464 43008 8504
rect 24076 8420 24116 8464
rect 25411 8463 25469 8464
rect 42928 8444 43008 8464
rect 3811 8380 3820 8420
rect 3860 8380 4396 8420
rect 4436 8380 4445 8420
rect 11875 8380 11884 8420
rect 11924 8380 20716 8420
rect 20756 8380 20765 8420
rect 21475 8380 21484 8420
rect 21524 8380 23308 8420
rect 23348 8380 24076 8420
rect 24116 8380 24125 8420
rect 24355 8380 24364 8420
rect 24404 8380 40876 8420
rect 40916 8380 40925 8420
rect 4919 8296 4928 8336
rect 4968 8296 5010 8336
rect 5050 8296 5092 8336
rect 5132 8296 5174 8336
rect 5214 8296 5256 8336
rect 5296 8296 5305 8336
rect 20039 8296 20048 8336
rect 20088 8296 20130 8336
rect 20170 8296 20212 8336
rect 20252 8296 20294 8336
rect 20334 8296 20376 8336
rect 20416 8296 20425 8336
rect 22531 8296 22540 8336
rect 22580 8296 22589 8336
rect 35159 8296 35168 8336
rect 35208 8296 35250 8336
rect 35290 8296 35332 8336
rect 35372 8296 35414 8336
rect 35454 8296 35496 8336
rect 35536 8296 35545 8336
rect 22540 8252 22580 8296
rect 2851 8212 2860 8252
rect 2900 8212 3340 8252
rect 3380 8212 3389 8252
rect 7171 8212 7180 8252
rect 7220 8212 10060 8252
rect 10100 8212 10109 8252
rect 17827 8212 17836 8252
rect 17876 8212 17885 8252
rect 18211 8212 18220 8252
rect 18260 8212 22580 8252
rect 22819 8212 22828 8252
rect 22868 8212 41260 8252
rect 41300 8212 41309 8252
rect 0 8168 80 8188
rect 17836 8168 17876 8212
rect 22828 8168 22868 8212
rect 42928 8168 43008 8188
rect 0 8128 1516 8168
rect 1556 8128 2540 8168
rect 2659 8128 2668 8168
rect 2708 8128 5356 8168
rect 5396 8128 5405 8168
rect 5923 8128 5932 8168
rect 5972 8128 8812 8168
rect 8852 8128 8861 8168
rect 10531 8128 10540 8168
rect 10580 8128 22868 8168
rect 33283 8128 33292 8168
rect 33332 8128 34348 8168
rect 34388 8128 34397 8168
rect 40675 8128 40684 8168
rect 40724 8128 43008 8168
rect 0 8108 80 8128
rect 2500 8084 2540 8128
rect 42928 8108 43008 8128
rect 2500 8044 16108 8084
rect 16148 8044 17836 8084
rect 17876 8044 17885 8084
rect 19075 8044 19084 8084
rect 19124 8044 21004 8084
rect 21044 8044 22348 8084
rect 22388 8044 22397 8084
rect 24931 8044 24940 8084
rect 24980 8044 26380 8084
rect 26420 8044 26429 8084
rect 28684 8044 29164 8084
rect 29204 8044 29213 8084
rect 31747 8044 31756 8084
rect 31796 8044 33004 8084
rect 33044 8044 33053 8084
rect 33667 8044 33676 8084
rect 33716 8044 38572 8084
rect 38612 8044 38621 8084
rect 9091 8000 9149 8001
rect 13795 8000 13853 8001
rect 17635 8000 17693 8001
rect 26380 8000 26420 8044
rect 28684 8000 28724 8044
rect 1219 7960 1228 8000
rect 1268 7960 4012 8000
rect 4052 7960 4061 8000
rect 7363 7960 7372 8000
rect 7412 7960 7948 8000
rect 7988 7960 7997 8000
rect 9006 7960 9100 8000
rect 9140 7960 9149 8000
rect 9283 7960 9292 8000
rect 9332 7960 10156 8000
rect 10196 7960 10676 8000
rect 10915 7960 10924 8000
rect 10964 7960 11116 8000
rect 11156 7960 11828 8000
rect 13710 7960 13804 8000
rect 13844 7960 13853 8000
rect 15043 7960 15052 8000
rect 15092 7960 17644 8000
rect 17684 7960 19852 8000
rect 19892 7960 19901 8000
rect 23011 7960 23020 8000
rect 23060 7960 25900 8000
rect 25940 7960 25949 8000
rect 26380 7960 28628 8000
rect 28675 7960 28684 8000
rect 28724 7960 28733 8000
rect 28960 7960 33580 8000
rect 33620 7960 33629 8000
rect 35299 7960 35308 8000
rect 35348 7960 37324 8000
rect 37364 7960 37373 8000
rect 38083 7960 38092 8000
rect 38132 7960 41300 8000
rect 4012 7916 4052 7960
rect 9091 7959 9149 7960
rect 10636 7916 10676 7960
rect 11788 7916 11828 7960
rect 13795 7959 13853 7960
rect 15052 7916 15092 7960
rect 17635 7959 17693 7960
rect 27715 7916 27773 7917
rect 28588 7916 28628 7960
rect 28960 7916 29000 7960
rect 33091 7916 33149 7917
rect 33292 7916 33332 7960
rect 41260 7916 41300 7960
rect 3139 7876 3148 7916
rect 3188 7876 3628 7916
rect 3668 7876 3677 7916
rect 4012 7876 10540 7916
rect 10580 7876 10589 7916
rect 10636 7876 11500 7916
rect 11540 7876 11549 7916
rect 11779 7876 11788 7916
rect 11828 7876 13420 7916
rect 13460 7876 15092 7916
rect 16003 7876 16012 7916
rect 16052 7876 17260 7916
rect 17300 7876 17309 7916
rect 17443 7876 17452 7916
rect 17492 7876 19084 7916
rect 19124 7876 19133 7916
rect 19363 7876 19372 7916
rect 19412 7876 21580 7916
rect 21620 7876 21629 7916
rect 24547 7876 24556 7916
rect 24596 7876 27148 7916
rect 27188 7876 27197 7916
rect 27630 7876 27724 7916
rect 27764 7876 28396 7916
rect 28436 7876 28445 7916
rect 28588 7876 29000 7916
rect 29251 7876 29260 7916
rect 29300 7876 31564 7916
rect 31604 7876 31613 7916
rect 32131 7876 32140 7916
rect 32180 7876 32524 7916
rect 32564 7876 32573 7916
rect 33006 7876 33100 7916
rect 33140 7876 33149 7916
rect 33283 7876 33292 7916
rect 33332 7876 33372 7916
rect 36835 7876 36844 7916
rect 36884 7876 37900 7916
rect 37940 7876 37949 7916
rect 40483 7876 40492 7916
rect 40532 7876 40541 7916
rect 41251 7876 41260 7916
rect 41300 7876 41309 7916
rect 27715 7875 27773 7876
rect 33091 7875 33149 7876
rect 0 7832 80 7852
rect 40492 7832 40532 7876
rect 42928 7832 43008 7852
rect 0 7792 1420 7832
rect 1460 7792 17356 7832
rect 17396 7792 17405 7832
rect 17827 7792 17836 7832
rect 17876 7792 33388 7832
rect 33428 7792 40532 7832
rect 41059 7792 41068 7832
rect 41108 7792 43008 7832
rect 0 7772 80 7792
rect 42928 7772 43008 7792
rect 4099 7708 4108 7748
rect 4148 7708 4492 7748
rect 4532 7708 4541 7748
rect 7555 7708 7564 7748
rect 7604 7708 9964 7748
rect 10004 7708 10013 7748
rect 11971 7708 11980 7748
rect 12020 7708 12844 7748
rect 12884 7708 12893 7748
rect 18604 7708 19564 7748
rect 19604 7708 19613 7748
rect 23875 7708 23884 7748
rect 23924 7708 24268 7748
rect 24308 7708 24317 7748
rect 26371 7708 26380 7748
rect 26420 7708 27052 7748
rect 27092 7708 27101 7748
rect 32515 7708 32524 7748
rect 32564 7708 36172 7748
rect 36212 7708 36460 7748
rect 36500 7708 36509 7748
rect 18604 7664 18644 7708
rect 547 7624 556 7664
rect 596 7624 7604 7664
rect 7843 7624 7852 7664
rect 7892 7624 9292 7664
rect 9332 7624 9341 7664
rect 10051 7624 10060 7664
rect 10100 7624 18644 7664
rect 18700 7624 19756 7664
rect 19796 7624 38092 7664
rect 38132 7624 38141 7664
rect 7564 7580 7604 7624
rect 9283 7580 9341 7581
rect 13795 7580 13853 7581
rect 18700 7580 18740 7624
rect 3679 7540 3688 7580
rect 3728 7540 3770 7580
rect 3810 7540 3852 7580
rect 3892 7540 3934 7580
rect 3974 7540 4016 7580
rect 4056 7540 4065 7580
rect 4291 7540 4300 7580
rect 4340 7540 6604 7580
rect 6644 7540 7508 7580
rect 7555 7540 7564 7580
rect 7604 7540 7613 7580
rect 8035 7540 8044 7580
rect 8084 7540 8620 7580
rect 8660 7540 8669 7580
rect 8803 7540 8812 7580
rect 8852 7540 9292 7580
rect 9332 7540 13132 7580
rect 13172 7540 13804 7580
rect 13844 7540 13853 7580
rect 14755 7540 14764 7580
rect 14804 7540 18740 7580
rect 18799 7540 18808 7580
rect 18848 7540 18890 7580
rect 18930 7540 18972 7580
rect 19012 7540 19054 7580
rect 19094 7540 19136 7580
rect 19176 7540 19185 7580
rect 26275 7540 26284 7580
rect 26324 7540 26860 7580
rect 26900 7540 26909 7580
rect 29155 7540 29164 7580
rect 29204 7540 31660 7580
rect 31700 7540 32428 7580
rect 32468 7540 32477 7580
rect 32611 7540 32620 7580
rect 32660 7540 33100 7580
rect 33140 7540 33149 7580
rect 33919 7540 33928 7580
rect 33968 7540 34010 7580
rect 34050 7540 34092 7580
rect 34132 7540 34174 7580
rect 34214 7540 34256 7580
rect 34296 7540 34305 7580
rect 0 7496 80 7516
rect 5347 7496 5405 7497
rect 7468 7496 7508 7540
rect 9283 7539 9341 7540
rect 13795 7539 13853 7540
rect 42928 7496 43008 7516
rect 0 7456 1612 7496
rect 1652 7456 2540 7496
rect 3427 7456 3436 7496
rect 3476 7456 5164 7496
rect 5204 7456 5213 7496
rect 5347 7456 5356 7496
rect 5396 7456 5452 7496
rect 5492 7456 5501 7496
rect 6019 7456 6028 7496
rect 6068 7456 6316 7496
rect 6356 7456 6365 7496
rect 7468 7456 7756 7496
rect 7796 7456 7805 7496
rect 16396 7456 28780 7496
rect 28820 7456 28829 7496
rect 40675 7456 40684 7496
rect 40724 7456 43008 7496
rect 0 7436 80 7456
rect 2500 7412 2540 7456
rect 4396 7412 4436 7456
rect 5347 7455 5405 7456
rect 2500 7372 3572 7412
rect 4387 7372 4396 7412
rect 4436 7372 4445 7412
rect 4492 7372 16300 7412
rect 16340 7372 16349 7412
rect 3532 7328 3572 7372
rect 4492 7328 4532 7372
rect 16396 7328 16436 7456
rect 42928 7436 43008 7456
rect 27715 7372 27724 7412
rect 27764 7372 37036 7412
rect 37076 7372 40492 7412
rect 40532 7372 40541 7412
rect 2947 7288 2956 7328
rect 2996 7288 3436 7328
rect 3476 7288 3485 7328
rect 3532 7288 4532 7328
rect 5347 7288 5356 7328
rect 5396 7288 6124 7328
rect 6164 7288 6173 7328
rect 6883 7288 6892 7328
rect 6932 7288 8332 7328
rect 8372 7288 8381 7328
rect 9667 7288 9676 7328
rect 9716 7288 9725 7328
rect 11884 7288 12556 7328
rect 12596 7288 16436 7328
rect 19843 7288 19852 7328
rect 19892 7288 29260 7328
rect 29300 7288 29309 7328
rect 5443 7244 5501 7245
rect 9676 7244 9716 7288
rect 5155 7204 5164 7244
rect 5204 7204 5452 7244
rect 5492 7204 6740 7244
rect 6787 7204 6796 7244
rect 6836 7204 7660 7244
rect 7700 7204 9716 7244
rect 5443 7203 5501 7204
rect 0 7160 80 7180
rect 6700 7160 6740 7204
rect 11884 7160 11924 7288
rect 28867 7244 28925 7245
rect 13411 7204 13420 7244
rect 13460 7204 14380 7244
rect 14420 7204 19508 7244
rect 19747 7204 19756 7244
rect 19796 7204 24596 7244
rect 28782 7204 28876 7244
rect 28916 7204 28925 7244
rect 16387 7160 16445 7161
rect 19363 7160 19421 7161
rect 0 7120 1900 7160
rect 1940 7120 1949 7160
rect 3235 7120 3244 7160
rect 3284 7120 4204 7160
rect 4244 7120 4253 7160
rect 5251 7120 5260 7160
rect 5300 7120 5309 7160
rect 5443 7120 5452 7160
rect 5492 7120 6220 7160
rect 6260 7120 6269 7160
rect 6700 7120 7852 7160
rect 7892 7120 8840 7160
rect 8995 7120 9004 7160
rect 9044 7120 9772 7160
rect 9812 7120 9821 7160
rect 11395 7120 11404 7160
rect 11444 7120 11692 7160
rect 11732 7120 11741 7160
rect 11875 7120 11884 7160
rect 11924 7120 11933 7160
rect 16291 7120 16300 7160
rect 16340 7120 16396 7160
rect 16436 7120 16445 7160
rect 19278 7120 19372 7160
rect 19412 7120 19421 7160
rect 19468 7160 19508 7204
rect 24163 7160 24221 7161
rect 19468 7120 21676 7160
rect 21716 7120 21725 7160
rect 24078 7120 24172 7160
rect 24212 7120 24221 7160
rect 0 7100 80 7120
rect 4387 7036 4396 7076
rect 4436 7036 4780 7076
rect 4820 7036 4829 7076
rect 5260 6992 5300 7120
rect 8800 7076 8840 7120
rect 11404 7076 11444 7120
rect 16387 7119 16445 7120
rect 19363 7119 19421 7120
rect 24163 7119 24221 7120
rect 24556 7076 24596 7204
rect 28867 7203 28925 7204
rect 25411 7160 25469 7161
rect 27619 7160 27677 7161
rect 42928 7160 43008 7180
rect 25326 7120 25420 7160
rect 25460 7120 25612 7160
rect 25652 7120 26476 7160
rect 26516 7120 26525 7160
rect 27619 7120 27628 7160
rect 27668 7120 27724 7160
rect 27764 7120 27773 7160
rect 28963 7120 28972 7160
rect 29012 7120 30124 7160
rect 30164 7120 30173 7160
rect 31363 7120 31372 7160
rect 31412 7120 32908 7160
rect 32948 7120 33772 7160
rect 33812 7120 34636 7160
rect 34676 7120 34685 7160
rect 37780 7120 38572 7160
rect 38612 7120 38860 7160
rect 38900 7120 38909 7160
rect 41059 7120 41068 7160
rect 41108 7120 43008 7160
rect 25411 7119 25469 7120
rect 27619 7119 27677 7120
rect 31651 7076 31709 7077
rect 7651 7036 7660 7076
rect 7700 7036 8236 7076
rect 8276 7036 8285 7076
rect 8800 7036 11444 7076
rect 14179 7036 14188 7076
rect 14228 7036 19756 7076
rect 19796 7036 19805 7076
rect 21091 7036 21100 7076
rect 21140 7036 21580 7076
rect 21620 7036 21629 7076
rect 24556 7036 29164 7076
rect 29204 7036 29213 7076
rect 31566 7036 31660 7076
rect 31700 7036 34348 7076
rect 34388 7036 34397 7076
rect 31651 7035 31709 7036
rect 12163 6992 12221 6993
rect 37780 6992 37820 7120
rect 42928 7100 43008 7120
rect 4867 6952 4876 6992
rect 4916 6952 4925 6992
rect 5260 6952 5452 6992
rect 5492 6952 5501 6992
rect 5923 6952 5932 6992
rect 5972 6952 6508 6992
rect 6548 6952 6557 6992
rect 6691 6952 6700 6992
rect 6740 6952 9196 6992
rect 9236 6952 9245 6992
rect 11587 6952 11596 6992
rect 11636 6952 12172 6992
rect 12212 6952 12221 6992
rect 13027 6952 13036 6992
rect 13076 6952 25900 6992
rect 25940 6952 25949 6992
rect 26275 6952 26284 6992
rect 26324 6952 37820 6992
rect 4195 6908 4253 6909
rect 4876 6908 4916 6952
rect 12163 6951 12221 6952
rect 3619 6868 3628 6908
rect 3668 6868 4204 6908
rect 4244 6868 8332 6908
rect 8372 6868 11884 6908
rect 11924 6868 11933 6908
rect 13891 6868 13900 6908
rect 13940 6868 21004 6908
rect 21044 6868 21053 6908
rect 25219 6868 25228 6908
rect 25268 6868 35692 6908
rect 35732 6868 35884 6908
rect 35924 6868 35933 6908
rect 4195 6867 4253 6868
rect 0 6824 80 6844
rect 42928 6824 43008 6844
rect 0 6784 1420 6824
rect 1460 6784 1469 6824
rect 4919 6784 4928 6824
rect 4968 6784 5010 6824
rect 5050 6784 5092 6824
rect 5132 6784 5174 6824
rect 5214 6784 5256 6824
rect 5296 6784 5305 6824
rect 5635 6784 5644 6824
rect 5684 6784 8140 6824
rect 8180 6784 11596 6824
rect 11636 6784 12364 6824
rect 12404 6784 12413 6824
rect 20039 6784 20048 6824
rect 20088 6784 20130 6824
rect 20170 6784 20212 6824
rect 20252 6784 20294 6824
rect 20334 6784 20376 6824
rect 20416 6784 20425 6824
rect 35159 6784 35168 6824
rect 35208 6784 35250 6824
rect 35290 6784 35332 6824
rect 35372 6784 35414 6824
rect 35454 6784 35496 6824
rect 35536 6784 35545 6824
rect 40675 6784 40684 6824
rect 40724 6784 43008 6824
rect 0 6764 80 6784
rect 42928 6764 43008 6784
rect 9283 6740 9341 6741
rect 9198 6700 9292 6740
rect 9332 6700 9341 6740
rect 9763 6700 9772 6740
rect 9812 6700 9821 6740
rect 9868 6700 14668 6740
rect 14708 6700 14717 6740
rect 17731 6700 17740 6740
rect 17780 6700 17932 6740
rect 17972 6700 17981 6740
rect 20140 6700 22060 6740
rect 22100 6700 25996 6740
rect 26036 6700 26284 6740
rect 26324 6700 26333 6740
rect 28963 6700 28972 6740
rect 29012 6700 30028 6740
rect 30068 6700 30077 6740
rect 32515 6700 32524 6740
rect 32564 6700 40876 6740
rect 40916 6700 40925 6740
rect 9283 6699 9341 6700
rect 5731 6656 5789 6657
rect 9772 6656 9812 6700
rect 3139 6616 3148 6656
rect 3188 6616 3197 6656
rect 5646 6616 5740 6656
rect 5780 6616 5789 6656
rect 8803 6616 8812 6656
rect 8852 6616 9812 6656
rect 3148 6572 3188 6616
rect 5731 6615 5789 6616
rect 9868 6572 9908 6700
rect 20140 6656 20180 6700
rect 14275 6616 14284 6656
rect 14324 6616 18412 6656
rect 18452 6616 20180 6656
rect 21283 6616 21292 6656
rect 21332 6616 21580 6656
rect 21620 6616 21629 6656
rect 24163 6616 24172 6656
rect 24212 6616 38036 6656
rect 19843 6572 19901 6573
rect 3148 6532 3340 6572
rect 3380 6532 3389 6572
rect 7555 6532 7564 6572
rect 7604 6532 9868 6572
rect 9908 6532 9917 6572
rect 11212 6532 19852 6572
rect 19892 6532 19901 6572
rect 20515 6532 20524 6572
rect 20564 6532 29740 6572
rect 29780 6532 30220 6572
rect 30260 6532 30269 6572
rect 30499 6532 30508 6572
rect 30548 6532 37820 6572
rect 0 6488 80 6508
rect 1699 6488 1757 6489
rect 4291 6488 4349 6489
rect 5347 6488 5405 6489
rect 0 6448 1516 6488
rect 1556 6448 1565 6488
rect 1699 6448 1708 6488
rect 1748 6448 1842 6488
rect 2659 6448 2668 6488
rect 2708 6448 2956 6488
rect 2996 6448 3005 6488
rect 3139 6448 3148 6488
rect 3188 6448 3916 6488
rect 3956 6448 3965 6488
rect 4206 6448 4300 6488
rect 4340 6448 4349 6488
rect 4579 6448 4588 6488
rect 4628 6448 5068 6488
rect 5108 6448 5117 6488
rect 5262 6448 5356 6488
rect 5396 6448 6220 6488
rect 6260 6448 7180 6488
rect 7220 6448 7229 6488
rect 9571 6448 9580 6488
rect 9620 6448 11116 6488
rect 11156 6448 11165 6488
rect 0 6428 80 6448
rect 1699 6447 1757 6448
rect 3916 6320 3956 6448
rect 4291 6447 4349 6448
rect 5347 6447 5405 6448
rect 11212 6404 11252 6532
rect 19843 6531 19901 6532
rect 14755 6488 14813 6489
rect 25315 6488 25373 6489
rect 14670 6448 14764 6488
rect 14804 6448 14813 6488
rect 17539 6448 17548 6488
rect 17588 6448 19756 6488
rect 19796 6448 19805 6488
rect 22060 6448 22636 6488
rect 22676 6448 25324 6488
rect 25364 6448 25373 6488
rect 14755 6447 14813 6448
rect 18691 6404 18749 6405
rect 22060 6404 22100 6448
rect 25315 6447 25373 6448
rect 27715 6488 27773 6489
rect 30508 6488 30548 6532
rect 27715 6448 27724 6488
rect 27764 6448 28300 6488
rect 28340 6448 30548 6488
rect 31459 6448 31468 6488
rect 31508 6448 31948 6488
rect 31988 6448 31997 6488
rect 27715 6447 27773 6448
rect 31747 6404 31805 6405
rect 4483 6364 4492 6404
rect 4532 6364 5780 6404
rect 7651 6364 7660 6404
rect 7700 6364 11252 6404
rect 11320 6364 12076 6404
rect 12116 6364 13900 6404
rect 13940 6364 13949 6404
rect 17443 6364 17452 6404
rect 17492 6364 18508 6404
rect 18548 6364 18557 6404
rect 18691 6364 18700 6404
rect 18740 6364 18988 6404
rect 19028 6364 22100 6404
rect 22147 6364 22156 6404
rect 22196 6364 25324 6404
rect 25364 6364 25373 6404
rect 28003 6364 28012 6404
rect 28052 6364 29548 6404
rect 29588 6364 31276 6404
rect 31316 6364 31325 6404
rect 31747 6364 31756 6404
rect 31796 6364 31890 6404
rect 32323 6364 32332 6404
rect 32372 6364 32812 6404
rect 32852 6364 32861 6404
rect 36547 6364 36556 6404
rect 36596 6364 36844 6404
rect 36884 6364 36893 6404
rect 5539 6320 5597 6321
rect 3916 6280 4300 6320
rect 4340 6280 5548 6320
rect 5588 6280 5597 6320
rect 5740 6320 5780 6364
rect 11320 6320 11360 6364
rect 17923 6320 17981 6321
rect 5740 6280 11360 6320
rect 17347 6280 17356 6320
rect 17396 6280 17932 6320
rect 17972 6280 17981 6320
rect 18508 6320 18548 6364
rect 18691 6363 18749 6364
rect 22156 6320 22196 6364
rect 31747 6363 31805 6364
rect 37780 6320 37820 6532
rect 37996 6488 38036 6616
rect 42928 6488 43008 6508
rect 37987 6448 37996 6488
rect 38036 6448 40780 6488
rect 40820 6448 40829 6488
rect 41059 6448 41068 6488
rect 41108 6448 43008 6488
rect 42928 6428 43008 6448
rect 37891 6364 37900 6404
rect 37940 6364 38092 6404
rect 38132 6364 39244 6404
rect 39284 6364 39293 6404
rect 39340 6364 41164 6404
rect 41204 6364 41213 6404
rect 39340 6320 39380 6364
rect 39619 6320 39677 6321
rect 18508 6280 22196 6320
rect 26947 6280 26956 6320
rect 26996 6280 36364 6320
rect 36404 6280 36413 6320
rect 37780 6280 39380 6320
rect 39534 6280 39628 6320
rect 39668 6280 39677 6320
rect 5539 6279 5597 6280
rect 17923 6279 17981 6280
rect 39619 6279 39677 6280
rect 4387 6236 4445 6237
rect 5731 6236 5789 6237
rect 4195 6196 4204 6236
rect 4244 6196 4396 6236
rect 4436 6196 4445 6236
rect 5347 6196 5356 6236
rect 5396 6196 5740 6236
rect 5780 6196 5789 6236
rect 11299 6196 11308 6236
rect 11348 6196 11596 6236
rect 11636 6196 11645 6236
rect 31747 6196 31756 6236
rect 31796 6196 32140 6236
rect 32180 6196 32189 6236
rect 33379 6196 33388 6236
rect 33428 6196 33964 6236
rect 34004 6196 34013 6236
rect 4387 6195 4445 6196
rect 5731 6195 5789 6196
rect 0 6152 80 6172
rect 5635 6152 5693 6153
rect 42928 6152 43008 6172
rect 0 6112 1324 6152
rect 1364 6112 1373 6152
rect 5550 6112 5644 6152
rect 5684 6112 5693 6152
rect 11203 6112 11212 6152
rect 11252 6112 18028 6152
rect 18068 6112 18077 6152
rect 30115 6112 30124 6152
rect 30164 6112 36076 6152
rect 36116 6112 36125 6152
rect 41059 6112 41068 6152
rect 41108 6112 43008 6152
rect 0 6092 80 6112
rect 5635 6111 5693 6112
rect 42928 6092 43008 6112
rect 21379 6068 21437 6069
rect 3679 6028 3688 6068
rect 3728 6028 3770 6068
rect 3810 6028 3852 6068
rect 3892 6028 3934 6068
rect 3974 6028 4016 6068
rect 4056 6028 4065 6068
rect 4867 6028 4876 6068
rect 4916 6028 6028 6068
rect 6068 6028 6077 6068
rect 6892 6028 11980 6068
rect 12020 6028 12029 6068
rect 18799 6028 18808 6068
rect 18848 6028 18890 6068
rect 18930 6028 18972 6068
rect 19012 6028 19054 6068
rect 19094 6028 19136 6068
rect 19176 6028 19185 6068
rect 21379 6028 21388 6068
rect 21428 6028 24460 6068
rect 24500 6028 33812 6068
rect 33919 6028 33928 6068
rect 33968 6028 34010 6068
rect 34050 6028 34092 6068
rect 34132 6028 34174 6068
rect 34214 6028 34256 6068
rect 34296 6028 34305 6068
rect 6892 5984 6932 6028
rect 21379 6027 21437 6028
rect 30115 5984 30173 5985
rect 31747 5984 31805 5985
rect 1219 5944 1228 5984
rect 1268 5944 6932 5984
rect 6988 5944 12460 5984
rect 12500 5944 12509 5984
rect 19555 5944 19564 5984
rect 19604 5944 30124 5984
rect 30164 5944 31756 5984
rect 31796 5944 31805 5984
rect 33772 5984 33812 6028
rect 33772 5944 35020 5984
rect 35060 5944 35404 5984
rect 35444 5944 35453 5984
rect 5539 5900 5597 5901
rect 4099 5860 4108 5900
rect 4148 5860 5260 5900
rect 5300 5860 5309 5900
rect 5539 5860 5548 5900
rect 5588 5860 5644 5900
rect 5684 5860 5693 5900
rect 5539 5859 5597 5860
rect 0 5816 80 5836
rect 6988 5816 7028 5944
rect 30115 5943 30173 5944
rect 31747 5943 31805 5944
rect 10243 5860 10252 5900
rect 10292 5860 17836 5900
rect 17876 5860 17885 5900
rect 26467 5860 26476 5900
rect 26516 5860 34828 5900
rect 34868 5860 34877 5900
rect 42928 5816 43008 5836
rect 0 5776 1036 5816
rect 1076 5776 1085 5816
rect 2467 5776 2476 5816
rect 2516 5776 7028 5816
rect 15811 5776 15820 5816
rect 15860 5776 25228 5816
rect 25268 5776 25277 5816
rect 28771 5776 28780 5816
rect 28820 5776 35980 5816
rect 36020 5776 39052 5816
rect 39092 5776 39101 5816
rect 40675 5776 40684 5816
rect 40724 5776 43008 5816
rect 0 5756 80 5776
rect 42928 5756 43008 5776
rect 19363 5732 19421 5733
rect 22051 5732 22109 5733
rect 5731 5692 5740 5732
rect 5780 5692 10540 5732
rect 10580 5692 10828 5732
rect 10868 5692 19372 5732
rect 19412 5692 19421 5732
rect 19651 5692 19660 5732
rect 19700 5692 20236 5732
rect 20276 5692 20285 5732
rect 21966 5692 22060 5732
rect 22100 5692 26476 5732
rect 26516 5692 26525 5732
rect 32899 5692 32908 5732
rect 32948 5692 33100 5732
rect 33140 5692 33292 5732
rect 33332 5692 33341 5732
rect 34531 5692 34540 5732
rect 34580 5692 40492 5732
rect 40532 5692 40541 5732
rect 19363 5691 19421 5692
rect 22051 5691 22109 5692
rect 8419 5648 8477 5649
rect 16387 5648 16445 5649
rect 3043 5608 3052 5648
rect 3092 5608 4108 5648
rect 4148 5608 4972 5648
rect 5012 5608 5356 5648
rect 5396 5608 5836 5648
rect 5876 5608 6988 5648
rect 7028 5608 7180 5648
rect 7220 5608 7229 5648
rect 8334 5608 8428 5648
rect 8468 5608 8477 5648
rect 13507 5608 13516 5648
rect 13556 5608 14380 5648
rect 14420 5608 16012 5648
rect 16052 5608 16061 5648
rect 16302 5608 16396 5648
rect 16436 5608 16445 5648
rect 17155 5608 17164 5648
rect 17204 5608 21676 5648
rect 21716 5608 29000 5648
rect 31939 5608 31948 5648
rect 31988 5608 32140 5648
rect 32180 5608 32189 5648
rect 33187 5608 33196 5648
rect 33236 5608 33772 5648
rect 33812 5608 33821 5648
rect 35395 5608 35404 5648
rect 35444 5608 39436 5648
rect 39476 5608 39485 5648
rect 8419 5607 8477 5608
rect 16387 5607 16445 5608
rect 4771 5564 4829 5565
rect 5347 5564 5405 5565
rect 28960 5564 29000 5608
rect 32611 5564 32669 5565
rect 4771 5524 4780 5564
rect 4820 5524 4876 5564
rect 4916 5524 4925 5564
rect 5156 5524 5165 5564
rect 5205 5524 5356 5564
rect 5396 5524 5405 5564
rect 6211 5524 6220 5564
rect 6260 5524 7468 5564
rect 7508 5524 11116 5564
rect 11156 5524 11165 5564
rect 15523 5524 15532 5564
rect 15572 5524 26860 5564
rect 26900 5524 26909 5564
rect 28960 5524 30164 5564
rect 31555 5524 31564 5564
rect 31604 5524 31852 5564
rect 31892 5524 31901 5564
rect 32611 5524 32620 5564
rect 32660 5524 36748 5564
rect 36788 5524 36797 5564
rect 4771 5523 4829 5524
rect 5347 5523 5405 5524
rect 0 5480 80 5500
rect 11779 5480 11837 5481
rect 30124 5480 30164 5524
rect 32611 5523 32669 5524
rect 42928 5480 43008 5500
rect 0 5440 7564 5480
rect 7604 5440 7613 5480
rect 11694 5440 11788 5480
rect 11828 5440 11837 5480
rect 14563 5440 14572 5480
rect 14612 5440 15436 5480
rect 15476 5440 15485 5480
rect 15532 5440 27724 5480
rect 27764 5440 27773 5480
rect 30115 5440 30124 5480
rect 30164 5440 40876 5480
rect 40916 5440 40925 5480
rect 41059 5440 41068 5480
rect 41108 5440 43008 5480
rect 0 5420 80 5440
rect 11779 5439 11837 5440
rect 10051 5396 10109 5397
rect 2275 5356 2284 5396
rect 2324 5356 10060 5396
rect 10100 5356 10109 5396
rect 10051 5355 10109 5356
rect 3523 5312 3581 5313
rect 5635 5312 5693 5313
rect 15532 5312 15572 5440
rect 27724 5396 27764 5440
rect 42928 5420 43008 5440
rect 20707 5356 20716 5396
rect 20756 5356 24748 5396
rect 24788 5356 24797 5396
rect 27724 5356 35788 5396
rect 35828 5356 35837 5396
rect 20611 5312 20669 5313
rect 30115 5312 30173 5313
rect 3523 5272 3532 5312
rect 3572 5272 4300 5312
rect 4340 5272 4349 5312
rect 4919 5272 4928 5312
rect 4968 5272 5010 5312
rect 5050 5272 5092 5312
rect 5132 5272 5174 5312
rect 5214 5272 5256 5312
rect 5296 5272 5305 5312
rect 5347 5272 5356 5312
rect 5396 5272 5644 5312
rect 5684 5272 5693 5312
rect 14851 5272 14860 5312
rect 14900 5272 15572 5312
rect 16003 5272 16012 5312
rect 16052 5272 17644 5312
rect 17684 5272 17693 5312
rect 17827 5272 17836 5312
rect 17876 5272 18124 5312
rect 18164 5272 18700 5312
rect 18740 5272 18749 5312
rect 20039 5272 20048 5312
rect 20088 5272 20130 5312
rect 20170 5272 20212 5312
rect 20252 5272 20294 5312
rect 20334 5272 20376 5312
rect 20416 5272 20425 5312
rect 20515 5272 20524 5312
rect 20564 5272 20620 5312
rect 20660 5272 20669 5312
rect 22915 5272 22924 5312
rect 22964 5272 23308 5312
rect 23348 5272 23357 5312
rect 30030 5272 30124 5312
rect 30164 5272 30173 5312
rect 33283 5272 33292 5312
rect 33332 5272 33676 5312
rect 33716 5272 33725 5312
rect 35159 5272 35168 5312
rect 35208 5272 35250 5312
rect 35290 5272 35332 5312
rect 35372 5272 35414 5312
rect 35454 5272 35496 5312
rect 35536 5272 35545 5312
rect 3523 5271 3581 5272
rect 5635 5271 5693 5272
rect 20611 5271 20669 5272
rect 30115 5271 30173 5272
rect 20995 5228 21053 5229
rect 1123 5188 1132 5228
rect 1172 5188 9100 5228
rect 9140 5188 9149 5228
rect 18403 5188 18412 5228
rect 18452 5188 20620 5228
rect 20660 5188 20669 5228
rect 20995 5188 21004 5228
rect 21044 5188 21196 5228
rect 21236 5188 21245 5228
rect 22147 5188 22156 5228
rect 22196 5188 28204 5228
rect 28244 5188 28253 5228
rect 32515 5188 32524 5228
rect 32564 5188 32573 5228
rect 33571 5188 33580 5228
rect 33620 5188 40204 5228
rect 40244 5188 40253 5228
rect 20995 5187 21053 5188
rect 0 5144 80 5164
rect 3715 5144 3773 5145
rect 4099 5144 4157 5145
rect 22156 5144 22196 5188
rect 0 5104 2668 5144
rect 2708 5104 3724 5144
rect 3764 5104 3773 5144
rect 3907 5104 3916 5144
rect 3956 5104 4108 5144
rect 4148 5104 4157 5144
rect 5251 5104 5260 5144
rect 5300 5104 5548 5144
rect 5588 5104 5597 5144
rect 6595 5104 6604 5144
rect 6644 5104 10252 5144
rect 10292 5104 10301 5144
rect 15715 5104 15724 5144
rect 15764 5104 18644 5144
rect 18691 5104 18700 5144
rect 18740 5104 22196 5144
rect 23491 5104 23500 5144
rect 23540 5104 23980 5144
rect 24020 5104 24029 5144
rect 25603 5104 25612 5144
rect 25652 5104 29548 5144
rect 29588 5104 29597 5144
rect 0 5084 80 5104
rect 3715 5103 3773 5104
rect 4099 5103 4157 5104
rect 18604 5060 18644 5104
rect 23971 5060 24029 5061
rect 32524 5060 32564 5188
rect 42928 5144 43008 5164
rect 35779 5104 35788 5144
rect 35828 5104 40396 5144
rect 40436 5104 40445 5144
rect 40675 5104 40684 5144
rect 40724 5104 43008 5144
rect 42928 5084 43008 5104
rect 1315 5020 1324 5060
rect 1364 5020 1708 5060
rect 1748 5020 17164 5060
rect 17204 5020 17213 5060
rect 18499 5020 18508 5060
rect 18548 5020 18557 5060
rect 18604 5020 23020 5060
rect 23060 5020 23069 5060
rect 23971 5020 23980 5060
rect 24020 5020 27052 5060
rect 27092 5020 27101 5060
rect 27148 5020 32564 5060
rect 1603 4976 1661 4977
rect 18508 4976 18548 5020
rect 23971 5019 24029 5020
rect 22627 4976 22685 4977
rect 26371 4976 26429 4977
rect 1518 4936 1612 4976
rect 1652 4936 1661 4976
rect 4099 4936 4108 4976
rect 4148 4936 4157 4976
rect 5059 4936 5068 4976
rect 5108 4936 5300 4976
rect 11107 4936 11116 4976
rect 11156 4936 12172 4976
rect 12212 4936 12221 4976
rect 16195 4936 16204 4976
rect 16244 4936 16780 4976
rect 16820 4936 16829 4976
rect 18508 4936 21140 4976
rect 1603 4935 1661 4936
rect 4108 4892 4148 4936
rect 3052 4852 4492 4892
rect 4532 4852 4541 4892
rect 0 4808 80 4828
rect 3052 4808 3092 4852
rect 5260 4808 5300 4936
rect 19267 4892 19325 4893
rect 21100 4892 21140 4936
rect 22627 4936 22636 4976
rect 22676 4936 22924 4976
rect 22964 4936 22973 4976
rect 23971 4936 23980 4976
rect 24020 4936 25900 4976
rect 25940 4936 25949 4976
rect 26286 4936 26380 4976
rect 26420 4936 26429 4976
rect 22627 4935 22685 4936
rect 26371 4935 26429 4936
rect 23875 4892 23933 4893
rect 27148 4892 27188 5020
rect 30211 4976 30269 4977
rect 29059 4936 29068 4976
rect 29108 4936 30220 4976
rect 30260 4936 30269 4976
rect 34147 4936 34156 4976
rect 34196 4936 40396 4976
rect 40436 4936 40445 4976
rect 30211 4935 30269 4936
rect 13603 4852 13612 4892
rect 13652 4852 16972 4892
rect 17012 4852 17260 4892
rect 17300 4852 17309 4892
rect 17635 4852 17644 4892
rect 17684 4852 18220 4892
rect 18260 4852 19084 4892
rect 19124 4852 19133 4892
rect 19182 4852 19276 4892
rect 19316 4852 19325 4892
rect 19267 4851 19325 4852
rect 20140 4852 20716 4892
rect 20756 4852 20765 4892
rect 21091 4852 21100 4892
rect 21140 4852 21149 4892
rect 23790 4852 23884 4892
rect 23924 4852 23933 4892
rect 24067 4852 24076 4892
rect 24116 4852 24460 4892
rect 24500 4852 24844 4892
rect 24884 4852 24893 4892
rect 25699 4852 25708 4892
rect 25748 4852 27188 4892
rect 27235 4892 27293 4893
rect 27235 4852 27244 4892
rect 27284 4852 32428 4892
rect 32468 4852 32477 4892
rect 32524 4852 35596 4892
rect 35636 4852 35645 4892
rect 37780 4852 40876 4892
rect 40916 4852 40925 4892
rect 20140 4808 20180 4852
rect 23875 4851 23933 4852
rect 27235 4851 27293 4852
rect 32524 4808 32564 4852
rect 37780 4808 37820 4852
rect 42928 4808 43008 4828
rect 0 4768 2380 4808
rect 2420 4768 2429 4808
rect 3043 4768 3052 4808
rect 3092 4768 3101 4808
rect 3331 4768 3340 4808
rect 3380 4768 3820 4808
rect 3860 4768 3869 4808
rect 5251 4768 5260 4808
rect 5300 4768 8524 4808
rect 8564 4768 10196 4808
rect 10531 4768 10540 4808
rect 10580 4768 12364 4808
rect 12404 4768 12413 4808
rect 15619 4768 15628 4808
rect 15668 4768 20180 4808
rect 21283 4768 21292 4808
rect 21332 4768 21484 4808
rect 21524 4768 21533 4808
rect 24259 4768 24268 4808
rect 24308 4768 24940 4808
rect 24980 4768 24989 4808
rect 31939 4768 31948 4808
rect 31988 4768 32236 4808
rect 32276 4768 32285 4808
rect 32515 4768 32524 4808
rect 32564 4768 32573 4808
rect 34435 4768 34444 4808
rect 34484 4768 37820 4808
rect 41443 4768 41452 4808
rect 41492 4768 43008 4808
rect 0 4748 80 4768
rect 5347 4724 5405 4725
rect 5155 4684 5164 4724
rect 5204 4684 5356 4724
rect 5396 4684 5405 4724
rect 5347 4683 5405 4684
rect 1987 4600 1996 4640
rect 2036 4600 8716 4640
rect 8756 4600 8765 4640
rect 3679 4516 3688 4556
rect 3728 4516 3770 4556
rect 3810 4516 3852 4556
rect 3892 4516 3934 4556
rect 3974 4516 4016 4556
rect 4056 4516 4065 4556
rect 0 4472 80 4492
rect 1219 4472 1277 4473
rect 5443 4472 5501 4473
rect 0 4432 1228 4472
rect 1268 4432 1277 4472
rect 3235 4432 3244 4472
rect 3284 4432 4300 4472
rect 4340 4432 4349 4472
rect 5155 4432 5164 4472
rect 5204 4432 5452 4472
rect 5492 4432 5501 4472
rect 8716 4472 8756 4600
rect 10156 4556 10196 4768
rect 42928 4748 43008 4768
rect 26371 4724 26429 4725
rect 10243 4684 10252 4724
rect 10292 4684 10636 4724
rect 10676 4684 13996 4724
rect 14036 4684 14045 4724
rect 14956 4684 18892 4724
rect 18932 4684 18941 4724
rect 19363 4684 19372 4724
rect 19412 4684 20044 4724
rect 20084 4684 24364 4724
rect 24404 4684 24413 4724
rect 26371 4684 26380 4724
rect 26420 4684 41260 4724
rect 41300 4684 41309 4724
rect 11587 4640 11645 4641
rect 14956 4640 14996 4684
rect 26371 4683 26429 4684
rect 11587 4600 11596 4640
rect 11636 4600 14996 4640
rect 17059 4600 17068 4640
rect 17108 4600 24172 4640
rect 24212 4600 24221 4640
rect 28291 4600 28300 4640
rect 28340 4600 40492 4640
rect 40532 4600 40541 4640
rect 11587 4599 11645 4600
rect 10156 4516 12748 4556
rect 12788 4516 13420 4556
rect 13460 4516 13469 4556
rect 18799 4516 18808 4556
rect 18848 4516 18890 4556
rect 18930 4516 18972 4556
rect 19012 4516 19054 4556
rect 19094 4516 19136 4556
rect 19176 4516 19185 4556
rect 21283 4516 21292 4556
rect 21332 4516 23692 4556
rect 23732 4516 30316 4556
rect 30356 4516 30365 4556
rect 33919 4516 33928 4556
rect 33968 4516 34010 4556
rect 34050 4516 34092 4556
rect 34132 4516 34174 4556
rect 34214 4516 34256 4556
rect 34296 4516 34305 4556
rect 42928 4472 43008 4492
rect 8716 4432 11360 4472
rect 11971 4432 11980 4472
rect 12020 4432 12268 4472
rect 12308 4432 14092 4472
rect 14132 4432 14141 4472
rect 20140 4432 24076 4472
rect 24116 4432 24125 4472
rect 28387 4432 28396 4472
rect 28436 4432 35020 4472
rect 35060 4432 35069 4472
rect 41059 4432 41068 4472
rect 41108 4432 43008 4472
rect 0 4412 80 4432
rect 1219 4431 1277 4432
rect 5443 4431 5501 4432
rect 4291 4388 4349 4389
rect 11320 4388 11360 4432
rect 20140 4388 20180 4432
rect 23779 4388 23837 4389
rect 34348 4388 34388 4432
rect 42928 4412 43008 4432
rect 3907 4348 3916 4388
rect 3956 4348 4300 4388
rect 4340 4348 8236 4388
rect 8276 4348 8285 4388
rect 8419 4348 8428 4388
rect 8468 4348 9484 4388
rect 9524 4348 9533 4388
rect 11320 4348 20180 4388
rect 22339 4348 22348 4388
rect 22388 4348 23596 4388
rect 23636 4348 23645 4388
rect 23779 4348 23788 4388
rect 23828 4348 29000 4388
rect 34339 4348 34348 4388
rect 34388 4348 34428 4388
rect 39811 4348 39820 4388
rect 39860 4348 40300 4388
rect 40340 4348 40349 4388
rect 4291 4347 4349 4348
rect 23779 4347 23837 4348
rect 28960 4304 29000 4348
rect 172 4264 12116 4304
rect 17347 4264 17356 4304
rect 17396 4264 17405 4304
rect 18595 4264 18604 4304
rect 18644 4264 19372 4304
rect 19412 4264 19564 4304
rect 19604 4264 19613 4304
rect 19939 4264 19948 4304
rect 19988 4264 23980 4304
rect 24020 4264 24029 4304
rect 28960 4264 38860 4304
rect 38900 4264 38909 4304
rect 0 4136 80 4156
rect 0 4076 116 4136
rect 76 4052 116 4076
rect 172 4052 212 4264
rect 2179 4180 2188 4220
rect 2228 4180 2380 4220
rect 2420 4180 8044 4220
rect 8084 4180 8093 4220
rect 8227 4180 8236 4220
rect 8276 4180 11980 4220
rect 12020 4180 12029 4220
rect 12076 4137 12116 4264
rect 17356 4220 17396 4264
rect 25699 4220 25757 4221
rect 16579 4180 16588 4220
rect 16628 4180 21716 4220
rect 24067 4180 24076 4220
rect 24116 4180 25132 4220
rect 25172 4180 25181 4220
rect 25614 4180 25708 4220
rect 25748 4180 25757 4220
rect 27523 4180 27532 4220
rect 27572 4180 27820 4220
rect 27860 4180 27869 4220
rect 32803 4180 32812 4220
rect 32852 4180 33676 4220
rect 33716 4180 33725 4220
rect 34636 4180 35404 4220
rect 35444 4180 35453 4220
rect 35875 4180 35884 4220
rect 35924 4180 40876 4220
rect 40916 4180 40925 4220
rect 4387 4136 4445 4137
rect 12067 4136 12125 4137
rect 19363 4136 19421 4137
rect 21676 4136 21716 4180
rect 25699 4179 25757 4180
rect 31747 4136 31805 4137
rect 34636 4136 34676 4180
rect 34819 4136 34877 4137
rect 3811 4096 3820 4136
rect 3860 4096 4396 4136
rect 4436 4096 5780 4136
rect 5827 4096 5836 4136
rect 5876 4096 6124 4136
rect 6164 4096 6173 4136
rect 9379 4096 9388 4136
rect 9428 4096 9964 4136
rect 10004 4096 11692 4136
rect 11732 4096 11741 4136
rect 11875 4096 11884 4136
rect 11924 4096 11933 4136
rect 12067 4096 12076 4136
rect 12116 4096 12210 4136
rect 12355 4096 12364 4136
rect 12404 4096 13324 4136
rect 13364 4096 15148 4136
rect 15188 4096 15916 4136
rect 15956 4096 15965 4136
rect 18211 4096 18220 4136
rect 18260 4096 18604 4136
rect 18644 4096 18653 4136
rect 19267 4096 19276 4136
rect 19316 4096 19372 4136
rect 19412 4096 19421 4136
rect 19555 4096 19564 4136
rect 19604 4096 20524 4136
rect 20564 4096 21292 4136
rect 21332 4096 21341 4136
rect 21667 4096 21676 4136
rect 21716 4096 28012 4136
rect 28052 4096 28061 4136
rect 31747 4096 31756 4136
rect 31796 4096 33580 4136
rect 33620 4096 34676 4136
rect 34734 4096 34828 4136
rect 34868 4096 34877 4136
rect 35404 4136 35444 4180
rect 42928 4136 43008 4156
rect 35404 4096 36268 4136
rect 36308 4096 36940 4136
rect 36980 4096 37132 4136
rect 37172 4096 38476 4136
rect 38516 4096 39148 4136
rect 39188 4096 40108 4136
rect 40148 4096 40157 4136
rect 40675 4096 40684 4136
rect 40724 4096 43008 4136
rect 4387 4095 4445 4096
rect 5740 4052 5780 4096
rect 10435 4052 10493 4053
rect 11884 4052 11924 4096
rect 12067 4095 12125 4096
rect 19363 4095 19421 4096
rect 31747 4095 31805 4096
rect 34819 4095 34877 4096
rect 42928 4076 43008 4096
rect 14179 4052 14237 4053
rect 15235 4052 15293 4053
rect 76 4012 212 4052
rect 2947 4012 2956 4052
rect 2996 4012 3148 4052
rect 3188 4012 3532 4052
rect 3572 4012 4684 4052
rect 4724 4012 4972 4052
rect 5012 4012 5644 4052
rect 5684 4012 5693 4052
rect 5740 4012 8840 4052
rect 10350 4012 10444 4052
rect 10484 4012 10493 4052
rect 3715 3928 3724 3968
rect 3764 3928 4492 3968
rect 4532 3928 4541 3968
rect 5251 3928 5260 3968
rect 5300 3928 5309 3968
rect 4099 3884 4157 3885
rect 5260 3884 5300 3928
rect 4003 3844 4012 3884
rect 4052 3844 4108 3884
rect 4148 3844 4157 3884
rect 4099 3843 4157 3844
rect 4780 3844 5300 3884
rect 0 3800 80 3820
rect 3235 3800 3293 3801
rect 4780 3800 4820 3844
rect 0 3760 2476 3800
rect 2516 3760 2525 3800
rect 3235 3760 3244 3800
rect 3284 3760 3340 3800
rect 3380 3760 3389 3800
rect 3436 3760 4820 3800
rect 4919 3760 4928 3800
rect 4968 3760 5010 3800
rect 5050 3760 5092 3800
rect 5132 3760 5174 3800
rect 5214 3760 5256 3800
rect 5296 3760 5305 3800
rect 0 3740 80 3760
rect 3235 3759 3293 3760
rect 0 3464 80 3484
rect 1603 3464 1661 3465
rect 3436 3464 3476 3760
rect 3619 3676 3628 3716
rect 3668 3676 4588 3716
rect 4628 3676 4637 3716
rect 5356 3632 5396 4012
rect 8800 3968 8840 4012
rect 10435 4011 10493 4012
rect 11320 4012 11980 4052
rect 12020 4012 13460 4052
rect 13507 4012 13516 4052
rect 13556 4012 13996 4052
rect 14036 4012 14045 4052
rect 14179 4012 14188 4052
rect 14228 4012 15244 4052
rect 15284 4012 15293 4052
rect 16963 4012 16972 4052
rect 17012 4012 21580 4052
rect 21620 4012 27628 4052
rect 27668 4012 38188 4052
rect 38228 4012 38380 4052
rect 38420 4012 38429 4052
rect 38851 4012 38860 4052
rect 38900 4012 41260 4052
rect 41300 4012 41309 4052
rect 11320 3968 11360 4012
rect 13420 3968 13460 4012
rect 14179 4011 14237 4012
rect 15235 4011 15293 4012
rect 7363 3928 7372 3968
rect 7412 3928 7756 3968
rect 7796 3928 7805 3968
rect 8800 3928 11360 3968
rect 11875 3928 11884 3968
rect 11924 3928 12460 3968
rect 12500 3928 12509 3968
rect 13420 3928 14092 3968
rect 14132 3928 14141 3968
rect 20035 3928 20044 3968
rect 20084 3928 21196 3968
rect 21236 3928 21245 3968
rect 23884 3928 26092 3968
rect 26132 3928 26141 3968
rect 29059 3928 29068 3968
rect 29108 3928 36652 3968
rect 36692 3928 36701 3968
rect 38275 3928 38284 3968
rect 38324 3928 38668 3968
rect 38708 3928 38717 3968
rect 19651 3884 19709 3885
rect 8035 3844 8044 3884
rect 8084 3844 19660 3884
rect 19700 3844 19709 3884
rect 19651 3843 19709 3844
rect 19660 3800 19700 3843
rect 21187 3800 21245 3801
rect 23884 3800 23924 3928
rect 23971 3844 23980 3884
rect 24020 3844 30412 3884
rect 30452 3844 30461 3884
rect 30979 3844 30988 3884
rect 31028 3844 31564 3884
rect 31604 3844 32428 3884
rect 32468 3844 32812 3884
rect 32852 3844 32861 3884
rect 42928 3800 43008 3820
rect 5923 3760 5932 3800
rect 5972 3760 6220 3800
rect 6260 3760 10252 3800
rect 10292 3760 10301 3800
rect 15043 3760 15052 3800
rect 15092 3760 16972 3800
rect 17012 3760 18220 3800
rect 18260 3760 18269 3800
rect 19651 3760 19660 3800
rect 19700 3760 19709 3800
rect 20039 3760 20048 3800
rect 20088 3760 20130 3800
rect 20170 3760 20212 3800
rect 20252 3760 20294 3800
rect 20334 3760 20376 3800
rect 20416 3760 20425 3800
rect 21187 3760 21196 3800
rect 21236 3760 21388 3800
rect 21428 3760 21437 3800
rect 21484 3760 23404 3800
rect 23444 3760 23453 3800
rect 23875 3760 23884 3800
rect 23924 3760 23933 3800
rect 24451 3760 24460 3800
rect 24500 3760 25844 3800
rect 26083 3760 26092 3800
rect 26132 3760 31756 3800
rect 31796 3760 31805 3800
rect 32035 3760 32044 3800
rect 32084 3760 34444 3800
rect 34484 3760 34493 3800
rect 35159 3760 35168 3800
rect 35208 3760 35250 3800
rect 35290 3760 35332 3800
rect 35372 3760 35414 3800
rect 35454 3760 35496 3800
rect 35536 3760 35545 3800
rect 40099 3760 40108 3800
rect 40148 3760 40588 3800
rect 40628 3760 40637 3800
rect 41443 3760 41452 3800
rect 41492 3760 43008 3800
rect 21187 3759 21245 3760
rect 21484 3716 21524 3760
rect 11299 3676 11308 3716
rect 11348 3676 16876 3716
rect 16916 3676 16925 3716
rect 20140 3676 21524 3716
rect 22627 3716 22685 3717
rect 24460 3716 24500 3760
rect 25804 3716 25844 3760
rect 42928 3740 43008 3760
rect 22627 3676 22636 3716
rect 22676 3676 24500 3716
rect 24739 3676 24748 3716
rect 24788 3676 25708 3716
rect 25748 3676 25757 3716
rect 25804 3676 26572 3716
rect 26612 3676 27532 3716
rect 27572 3676 27581 3716
rect 30787 3676 30796 3716
rect 30836 3676 31276 3716
rect 31316 3676 33100 3716
rect 33140 3676 35692 3716
rect 35732 3676 38092 3716
rect 38132 3676 38284 3716
rect 38324 3676 38333 3716
rect 11203 3632 11261 3633
rect 20140 3632 20180 3676
rect 22627 3675 22685 3676
rect 32707 3632 32765 3633
rect 3907 3592 3916 3632
rect 3956 3592 4780 3632
rect 4820 3592 4829 3632
rect 5155 3592 5164 3632
rect 5204 3592 5396 3632
rect 10147 3592 10156 3632
rect 10196 3592 10924 3632
rect 10964 3592 10973 3632
rect 11118 3592 11212 3632
rect 11252 3592 11261 3632
rect 11875 3592 11884 3632
rect 11924 3592 12076 3632
rect 12116 3592 12125 3632
rect 12835 3592 12844 3632
rect 12884 3592 20180 3632
rect 20899 3592 20908 3632
rect 20948 3592 21292 3632
rect 21332 3592 21341 3632
rect 22627 3592 22636 3632
rect 22676 3592 22828 3632
rect 22868 3592 22877 3632
rect 25507 3592 25516 3632
rect 25556 3592 25996 3632
rect 26036 3592 26045 3632
rect 28771 3592 28780 3632
rect 28820 3592 32044 3632
rect 32084 3592 32093 3632
rect 32707 3592 32716 3632
rect 32756 3592 36748 3632
rect 36788 3592 36797 3632
rect 36844 3592 40492 3632
rect 40532 3592 40541 3632
rect 11203 3591 11261 3592
rect 32707 3591 32765 3592
rect 12163 3548 12221 3549
rect 4012 3508 4396 3548
rect 4436 3508 5068 3548
rect 5108 3508 7084 3548
rect 7124 3508 7133 3548
rect 7267 3508 7276 3548
rect 7316 3508 7852 3548
rect 7892 3508 7901 3548
rect 10723 3508 10732 3548
rect 10772 3508 11116 3548
rect 11156 3508 11165 3548
rect 12078 3508 12172 3548
rect 12212 3508 17356 3548
rect 17396 3508 17405 3548
rect 18019 3508 18028 3548
rect 18068 3508 23308 3548
rect 23348 3508 23357 3548
rect 23491 3508 23500 3548
rect 23540 3508 23692 3548
rect 23732 3508 23741 3548
rect 25315 3508 25324 3548
rect 25364 3508 26668 3548
rect 26708 3508 26717 3548
rect 31459 3508 31468 3548
rect 31508 3508 31756 3548
rect 31796 3508 31805 3548
rect 33475 3508 33484 3548
rect 33524 3508 34636 3548
rect 34676 3508 34685 3548
rect 4012 3464 4052 3508
rect 12163 3507 12221 3508
rect 14179 3464 14237 3465
rect 14956 3464 14996 3508
rect 16387 3464 16445 3465
rect 20995 3464 21053 3465
rect 21475 3464 21533 3465
rect 22627 3464 22685 3465
rect 23779 3464 23837 3465
rect 24451 3464 24509 3465
rect 31843 3464 31901 3465
rect 34435 3464 34493 3465
rect 36844 3464 36884 3592
rect 39523 3548 39581 3549
rect 39438 3508 39532 3548
rect 39572 3508 40972 3548
rect 41012 3508 41021 3548
rect 39523 3507 39581 3508
rect 38083 3464 38141 3465
rect 42928 3464 43008 3484
rect 0 3424 1228 3464
rect 1268 3424 1277 3464
rect 1518 3424 1612 3464
rect 1652 3424 1900 3464
rect 1940 3424 1949 3464
rect 3427 3424 3436 3464
rect 3476 3424 3485 3464
rect 4003 3424 4012 3464
rect 4052 3424 4061 3464
rect 4483 3424 4492 3464
rect 4532 3424 4541 3464
rect 4675 3424 4684 3464
rect 4724 3424 4972 3464
rect 5012 3424 5021 3464
rect 5155 3424 5164 3464
rect 5204 3424 5548 3464
rect 5588 3424 5597 3464
rect 8131 3424 8140 3464
rect 8180 3424 8189 3464
rect 8611 3424 8620 3464
rect 8660 3424 9868 3464
rect 9908 3424 11212 3464
rect 11252 3424 13996 3464
rect 14036 3424 14045 3464
rect 14179 3424 14188 3464
rect 14228 3424 14322 3464
rect 14947 3424 14956 3464
rect 14996 3424 15005 3464
rect 16302 3424 16396 3464
rect 16436 3424 16445 3464
rect 20910 3424 21004 3464
rect 21044 3424 21053 3464
rect 21390 3424 21484 3464
rect 21524 3424 22444 3464
rect 22484 3424 22493 3464
rect 22627 3424 22636 3464
rect 22676 3424 22770 3464
rect 23203 3424 23212 3464
rect 23252 3424 23788 3464
rect 23828 3424 23837 3464
rect 24366 3424 24460 3464
rect 24500 3424 24509 3464
rect 25987 3424 25996 3464
rect 26036 3424 28588 3464
rect 28628 3424 28637 3464
rect 31758 3424 31852 3464
rect 31892 3424 31901 3464
rect 34350 3424 34444 3464
rect 34484 3424 35788 3464
rect 35828 3424 35837 3464
rect 35980 3424 36884 3464
rect 37699 3424 37708 3464
rect 37748 3424 38092 3464
rect 38132 3424 38141 3464
rect 41059 3424 41068 3464
rect 41108 3424 43008 3464
rect 0 3404 80 3424
rect 1603 3423 1661 3424
rect 2947 3340 2956 3380
rect 2996 3340 3628 3380
rect 3668 3340 3677 3380
rect 4492 3296 4532 3424
rect 8140 3380 8180 3424
rect 14179 3423 14237 3424
rect 16387 3423 16445 3424
rect 20995 3423 21053 3424
rect 21475 3423 21533 3424
rect 22627 3423 22685 3424
rect 23779 3423 23837 3424
rect 24451 3423 24509 3424
rect 31843 3423 31901 3424
rect 34435 3423 34493 3424
rect 12355 3380 12413 3381
rect 21955 3380 22013 3381
rect 22636 3380 22676 3423
rect 31852 3380 31892 3423
rect 4579 3340 4588 3380
rect 4628 3340 8180 3380
rect 8707 3340 8716 3380
rect 8756 3340 12364 3380
rect 12404 3340 12413 3380
rect 20899 3340 20908 3380
rect 20948 3340 21964 3380
rect 22004 3340 22676 3380
rect 24163 3340 24172 3380
rect 24212 3340 24652 3380
rect 24692 3340 24701 3380
rect 26851 3340 26860 3380
rect 26900 3340 27628 3380
rect 27668 3340 29356 3380
rect 29396 3340 29405 3380
rect 31852 3340 35884 3380
rect 35924 3340 35933 3380
rect 12355 3339 12413 3340
rect 21955 3339 22013 3340
rect 35980 3296 36020 3424
rect 38083 3423 38141 3424
rect 42928 3404 43008 3424
rect 36547 3340 36556 3380
rect 36596 3340 37324 3380
rect 37364 3340 40876 3380
rect 40916 3340 40925 3380
rect 38083 3296 38141 3297
rect 4099 3256 4108 3296
rect 4148 3256 4532 3296
rect 15139 3256 15148 3296
rect 15188 3256 15436 3296
rect 15476 3256 17644 3296
rect 17684 3256 17693 3296
rect 22435 3256 22444 3296
rect 22484 3256 28108 3296
rect 28148 3256 28300 3296
rect 28340 3256 28349 3296
rect 30019 3256 30028 3296
rect 30068 3256 36020 3296
rect 37998 3256 38092 3296
rect 38132 3256 38141 3296
rect 38083 3255 38141 3256
rect 18883 3212 18941 3213
rect 1027 3172 1036 3212
rect 1076 3172 5932 3212
rect 5972 3172 5981 3212
rect 13411 3172 13420 3212
rect 13460 3172 18892 3212
rect 18932 3172 18941 3212
rect 26275 3172 26284 3212
rect 26324 3172 32428 3212
rect 32468 3172 32477 3212
rect 32524 3172 34540 3212
rect 34580 3172 34589 3212
rect 40675 3172 40684 3212
rect 40724 3172 40733 3212
rect 18883 3171 18941 3172
rect 0 3128 80 3148
rect 27235 3128 27293 3129
rect 0 3088 2284 3128
rect 2324 3088 2333 3128
rect 2380 3088 8716 3128
rect 8756 3088 8765 3128
rect 14467 3088 14476 3128
rect 14516 3088 15244 3128
rect 15284 3088 27244 3128
rect 27284 3088 27293 3128
rect 0 3068 80 3088
rect 2380 3044 2420 3088
rect 27235 3087 27293 3088
rect 30211 3128 30269 3129
rect 32524 3128 32564 3172
rect 30211 3088 30220 3128
rect 30260 3088 30412 3128
rect 30452 3088 32564 3128
rect 32611 3128 32669 3129
rect 37315 3128 37373 3129
rect 40684 3128 40724 3172
rect 42928 3128 43008 3148
rect 32611 3088 32620 3128
rect 32660 3088 36364 3128
rect 36404 3088 36413 3128
rect 37315 3088 37324 3128
rect 37364 3088 37820 3128
rect 40684 3088 43008 3128
rect 30211 3087 30269 3088
rect 32611 3087 32669 3088
rect 37315 3087 37373 3088
rect 3235 3044 3293 3045
rect 20035 3044 20093 3045
rect 37780 3044 37820 3088
rect 42928 3068 43008 3088
rect 1507 3004 1516 3044
rect 1556 3004 2420 3044
rect 3150 3004 3244 3044
rect 3284 3004 3293 3044
rect 3523 3004 3532 3044
rect 3572 3004 3581 3044
rect 3679 3004 3688 3044
rect 3728 3004 3770 3044
rect 3810 3004 3852 3044
rect 3892 3004 3934 3044
rect 3974 3004 4016 3044
rect 4056 3004 4065 3044
rect 16675 3004 16684 3044
rect 16724 3004 16972 3044
rect 17012 3004 17021 3044
rect 18799 3004 18808 3044
rect 18848 3004 18890 3044
rect 18930 3004 18972 3044
rect 19012 3004 19054 3044
rect 19094 3004 19136 3044
rect 19176 3004 19185 3044
rect 19939 3004 19948 3044
rect 19988 3004 20044 3044
rect 20084 3004 20093 3044
rect 20227 3004 20236 3044
rect 20276 3004 23116 3044
rect 23156 3004 24076 3044
rect 24116 3004 24125 3044
rect 24172 3004 25804 3044
rect 25844 3004 25996 3044
rect 26036 3004 26045 3044
rect 26467 3004 26476 3044
rect 26516 3004 27148 3044
rect 27188 3004 27197 3044
rect 29347 3004 29356 3044
rect 29396 3004 30796 3044
rect 30836 3004 30845 3044
rect 33919 3004 33928 3044
rect 33968 3004 34010 3044
rect 34050 3004 34092 3044
rect 34132 3004 34174 3044
rect 34214 3004 34256 3044
rect 34296 3004 34305 3044
rect 35203 3004 35212 3044
rect 35252 3004 37132 3044
rect 37172 3004 37181 3044
rect 37780 3004 41260 3044
rect 41300 3004 41309 3044
rect 3235 3003 3293 3004
rect 3532 2876 3572 3004
rect 20035 3003 20093 3004
rect 24172 2960 24212 3004
rect 17347 2920 17356 2960
rect 17396 2920 20140 2960
rect 20180 2920 22580 2960
rect 23587 2920 23596 2960
rect 23636 2920 23788 2960
rect 23828 2920 23837 2960
rect 24163 2920 24172 2960
rect 24212 2920 24221 2960
rect 25699 2920 25708 2960
rect 25748 2920 36556 2960
rect 36596 2920 36605 2960
rect 4771 2876 4829 2877
rect 15427 2876 15485 2877
rect 22540 2876 22580 2920
rect 3532 2836 4012 2876
rect 4052 2836 4061 2876
rect 4771 2836 4780 2876
rect 4820 2836 4972 2876
rect 5012 2836 13132 2876
rect 13172 2836 14764 2876
rect 14804 2836 15436 2876
rect 15476 2836 15485 2876
rect 15619 2836 15628 2876
rect 15668 2836 21716 2876
rect 22540 2836 32756 2876
rect 32995 2836 33004 2876
rect 33044 2836 33484 2876
rect 33524 2836 33533 2876
rect 34339 2836 34348 2876
rect 34388 2836 40876 2876
rect 40916 2836 40925 2876
rect 4771 2835 4829 2836
rect 15427 2835 15485 2836
rect 0 2792 80 2812
rect 4195 2792 4253 2793
rect 18115 2792 18173 2793
rect 21676 2792 21716 2836
rect 0 2752 1132 2792
rect 1172 2752 1181 2792
rect 3331 2752 3340 2792
rect 3380 2752 3724 2792
rect 3764 2752 3773 2792
rect 4195 2752 4204 2792
rect 4244 2752 4300 2792
rect 4340 2752 4349 2792
rect 7555 2752 7564 2792
rect 7604 2752 17932 2792
rect 17972 2752 18124 2792
rect 18164 2752 18173 2792
rect 19747 2752 19756 2792
rect 19796 2752 21620 2792
rect 21676 2752 23212 2792
rect 23252 2752 23261 2792
rect 24076 2752 24748 2792
rect 24788 2752 25132 2792
rect 25172 2752 25181 2792
rect 27523 2752 27532 2792
rect 27572 2752 28972 2792
rect 29012 2752 29164 2792
rect 29204 2752 30220 2792
rect 30260 2752 30269 2792
rect 0 2732 80 2752
rect 4195 2751 4253 2752
rect 18115 2751 18173 2752
rect 3523 2708 3581 2709
rect 10435 2708 10493 2709
rect 21580 2708 21620 2752
rect 24076 2708 24116 2752
rect 32716 2708 32756 2836
rect 42928 2792 43008 2812
rect 32899 2752 32908 2792
rect 32948 2752 33292 2792
rect 33332 2752 33341 2792
rect 34243 2752 34252 2792
rect 34292 2752 34540 2792
rect 34580 2752 34589 2792
rect 36355 2752 36364 2792
rect 36404 2752 36748 2792
rect 36788 2752 36797 2792
rect 41059 2752 41068 2792
rect 41108 2752 43008 2792
rect 42928 2732 43008 2752
rect 3438 2668 3532 2708
rect 3572 2668 3581 2708
rect 3811 2668 3820 2708
rect 3860 2668 7468 2708
rect 7508 2668 7517 2708
rect 10435 2668 10444 2708
rect 10484 2668 11360 2708
rect 11971 2668 11980 2708
rect 12020 2668 12172 2708
rect 12212 2668 14476 2708
rect 14516 2668 15724 2708
rect 15764 2668 16780 2708
rect 16820 2668 16829 2708
rect 19267 2668 19276 2708
rect 19316 2668 20908 2708
rect 20948 2668 20957 2708
rect 21580 2668 24116 2708
rect 26179 2668 26188 2708
rect 26228 2668 28916 2708
rect 32716 2668 33044 2708
rect 35875 2668 35884 2708
rect 35924 2668 36556 2708
rect 36596 2668 36605 2708
rect 3523 2667 3581 2668
rect 10435 2667 10493 2668
rect 5923 2624 5981 2625
rect 11320 2624 11360 2668
rect 16099 2624 16157 2625
rect 20227 2624 20285 2625
rect 28675 2624 28733 2625
rect 28876 2624 28916 2668
rect 33004 2624 33044 2668
rect 3427 2584 3436 2624
rect 3476 2584 4148 2624
rect 4195 2584 4204 2624
rect 4244 2584 4253 2624
rect 5838 2584 5932 2624
rect 5972 2584 5981 2624
rect 7171 2584 7180 2624
rect 7220 2584 8812 2624
rect 8852 2584 8861 2624
rect 9091 2584 9100 2624
rect 9140 2584 9149 2624
rect 9667 2584 9676 2624
rect 9716 2584 10676 2624
rect 11320 2584 13420 2624
rect 13460 2584 13469 2624
rect 13699 2584 13708 2624
rect 13748 2584 15244 2624
rect 15284 2584 15293 2624
rect 15907 2584 15916 2624
rect 15956 2584 16108 2624
rect 16148 2584 16157 2624
rect 17155 2584 17164 2624
rect 17204 2584 17644 2624
rect 17684 2584 18604 2624
rect 18644 2584 18653 2624
rect 19372 2584 19564 2624
rect 19604 2584 19613 2624
rect 19747 2584 19756 2624
rect 19796 2584 20180 2624
rect 4108 2540 4148 2584
rect 4099 2500 4108 2540
rect 4148 2500 4157 2540
rect 0 2456 80 2476
rect 4204 2456 4244 2584
rect 5923 2583 5981 2584
rect 5124 2500 5164 2540
rect 5204 2500 5213 2540
rect 5164 2456 5204 2500
rect 7180 2456 7220 2584
rect 0 2416 2540 2456
rect 4204 2416 5204 2456
rect 5347 2416 5356 2456
rect 5396 2416 7220 2456
rect 9100 2456 9140 2584
rect 10636 2456 10676 2584
rect 16099 2583 16157 2584
rect 19372 2540 19412 2584
rect 20140 2540 20180 2584
rect 20227 2584 20236 2624
rect 20276 2584 20468 2624
rect 23491 2584 23500 2624
rect 23540 2584 24460 2624
rect 24500 2584 24509 2624
rect 28675 2584 28684 2624
rect 28724 2584 28780 2624
rect 28820 2584 28829 2624
rect 28876 2584 29644 2624
rect 29684 2584 29693 2624
rect 30115 2584 30124 2624
rect 30164 2584 31852 2624
rect 31892 2584 32236 2624
rect 32276 2584 32285 2624
rect 32332 2584 32524 2624
rect 32564 2584 32573 2624
rect 33004 2584 34732 2624
rect 34772 2584 35212 2624
rect 35252 2584 35261 2624
rect 36067 2584 36076 2624
rect 36116 2584 36460 2624
rect 36500 2584 36509 2624
rect 37603 2584 37612 2624
rect 37652 2584 38996 2624
rect 20227 2583 20285 2584
rect 11491 2500 11500 2540
rect 11540 2500 11692 2540
rect 11732 2500 11741 2540
rect 15108 2500 15148 2540
rect 15188 2500 15197 2540
rect 19363 2500 19372 2540
rect 19412 2500 19421 2540
rect 19756 2500 20084 2540
rect 20140 2500 20236 2540
rect 20276 2500 20285 2540
rect 15148 2456 15188 2500
rect 19756 2456 19796 2500
rect 9100 2416 10540 2456
rect 10580 2416 10589 2456
rect 10636 2416 11360 2456
rect 12643 2416 12652 2456
rect 12692 2416 13036 2456
rect 13076 2416 13085 2456
rect 14755 2416 14764 2456
rect 14804 2416 15188 2456
rect 15244 2416 19796 2456
rect 0 2396 80 2416
rect 2500 2372 2540 2416
rect 8035 2372 8093 2373
rect 11320 2372 11360 2416
rect 15139 2372 15197 2373
rect 2500 2332 8044 2372
rect 8084 2332 8093 2372
rect 10435 2332 10444 2372
rect 10484 2332 11212 2372
rect 11252 2332 11261 2372
rect 11320 2332 15148 2372
rect 15188 2332 15197 2372
rect 8035 2331 8093 2332
rect 15139 2331 15197 2332
rect 11587 2288 11645 2289
rect 15244 2288 15284 2416
rect 15331 2372 15389 2373
rect 20044 2372 20084 2500
rect 20323 2456 20381 2457
rect 20238 2416 20332 2456
rect 20372 2416 20381 2456
rect 20428 2456 20468 2584
rect 28675 2583 28733 2584
rect 30595 2540 30653 2541
rect 31084 2540 31124 2584
rect 27204 2500 27244 2540
rect 27284 2500 27293 2540
rect 30595 2500 30604 2540
rect 30644 2500 30892 2540
rect 30932 2500 30941 2540
rect 31075 2500 31084 2540
rect 31124 2500 31133 2540
rect 27244 2456 27284 2500
rect 30595 2499 30653 2500
rect 32332 2456 32372 2584
rect 38956 2540 38996 2584
rect 38947 2500 38956 2540
rect 38996 2500 39005 2540
rect 42928 2456 43008 2476
rect 20428 2416 20716 2456
rect 20756 2416 20765 2456
rect 27244 2416 27916 2456
rect 27956 2416 27965 2456
rect 28579 2416 28588 2456
rect 28628 2416 32372 2456
rect 41443 2416 41452 2456
rect 41492 2416 43008 2456
rect 20323 2415 20381 2416
rect 42928 2396 43008 2416
rect 15331 2332 15340 2372
rect 15380 2332 19948 2372
rect 19988 2332 19997 2372
rect 20044 2332 27820 2372
rect 27860 2332 27869 2372
rect 28003 2332 28012 2372
rect 28052 2332 28780 2372
rect 28820 2332 32332 2372
rect 32372 2332 32381 2372
rect 33571 2332 33580 2372
rect 33620 2332 39052 2372
rect 39092 2332 39101 2372
rect 15331 2331 15389 2332
rect 19939 2288 19997 2289
rect 23971 2288 24029 2289
rect 4919 2248 4928 2288
rect 4968 2248 5010 2288
rect 5050 2248 5092 2288
rect 5132 2248 5174 2288
rect 5214 2248 5256 2288
rect 5296 2248 5305 2288
rect 6595 2248 6604 2288
rect 6644 2248 8908 2288
rect 8948 2248 11596 2288
rect 11636 2248 11645 2288
rect 11779 2248 11788 2288
rect 11828 2248 15284 2288
rect 15340 2248 18892 2288
rect 18932 2248 18941 2288
rect 19843 2248 19852 2288
rect 19892 2248 19948 2288
rect 19988 2248 19997 2288
rect 20039 2248 20048 2288
rect 20088 2248 20130 2288
rect 20170 2248 20212 2288
rect 20252 2248 20294 2288
rect 20334 2248 20376 2288
rect 20416 2248 20425 2288
rect 23875 2248 23884 2288
rect 23924 2248 23980 2288
rect 24020 2248 24029 2288
rect 24547 2248 24556 2288
rect 24596 2248 24940 2288
rect 24980 2248 24989 2288
rect 29923 2248 29932 2288
rect 29972 2248 30412 2288
rect 30452 2248 30461 2288
rect 35159 2248 35168 2288
rect 35208 2248 35250 2288
rect 35290 2248 35332 2288
rect 35372 2248 35414 2288
rect 35454 2248 35496 2288
rect 35536 2248 35545 2288
rect 35779 2248 35788 2288
rect 35828 2248 37036 2288
rect 37076 2248 37085 2288
rect 11587 2247 11645 2248
rect 15340 2204 15380 2248
rect 19939 2247 19997 2248
rect 23971 2247 24029 2248
rect 5827 2164 5836 2204
rect 5876 2164 6028 2204
rect 6068 2164 8332 2204
rect 8372 2164 8381 2204
rect 9859 2164 9868 2204
rect 9908 2164 15380 2204
rect 15427 2204 15485 2205
rect 15427 2164 15436 2204
rect 15476 2164 20180 2204
rect 26083 2164 26092 2204
rect 26132 2164 26380 2204
rect 26420 2164 26429 2204
rect 28867 2164 28876 2204
rect 28916 2164 39724 2204
rect 39764 2164 39773 2204
rect 15427 2163 15485 2164
rect 0 2120 80 2140
rect 20140 2120 20180 2164
rect 42928 2120 43008 2140
rect 0 2080 7660 2120
rect 7700 2080 7709 2120
rect 8131 2080 8140 2120
rect 8180 2080 9484 2120
rect 9524 2080 10388 2120
rect 10627 2080 10636 2120
rect 10676 2080 12652 2120
rect 12692 2080 12701 2120
rect 13987 2080 13996 2120
rect 14036 2080 14668 2120
rect 14708 2080 14717 2120
rect 14851 2080 14860 2120
rect 14900 2080 15436 2120
rect 15476 2080 15485 2120
rect 17155 2080 17164 2120
rect 17204 2080 17452 2120
rect 17492 2080 17501 2120
rect 18883 2080 18892 2120
rect 18932 2080 19756 2120
rect 19796 2080 19805 2120
rect 20140 2080 20428 2120
rect 20468 2080 20477 2120
rect 23395 2080 23404 2120
rect 23444 2080 28396 2120
rect 28436 2080 28445 2120
rect 31267 2080 31276 2120
rect 31316 2080 32044 2120
rect 32084 2080 32093 2120
rect 38755 2080 38764 2120
rect 38804 2080 38956 2120
rect 38996 2080 39005 2120
rect 41539 2080 41548 2120
rect 41588 2080 43008 2120
rect 0 2060 80 2080
rect 7267 2036 7325 2037
rect 9571 2036 9629 2037
rect 5251 1996 5260 2036
rect 5300 1996 7084 2036
rect 7124 1996 7133 2036
rect 7267 1996 7276 2036
rect 7316 1996 7410 2036
rect 9486 1996 9580 2036
rect 9620 1996 9629 2036
rect 10348 2036 10388 2080
rect 42928 2060 43008 2080
rect 29827 2036 29885 2037
rect 10348 1996 11360 2036
rect 12835 1996 12844 2036
rect 12884 1996 21484 2036
rect 21524 1996 21533 2036
rect 25324 1996 28108 2036
rect 28148 1996 28157 2036
rect 29742 1996 29836 2036
rect 29876 1996 29885 2036
rect 33283 1996 33292 2036
rect 33332 1996 37900 2036
rect 37940 1996 37949 2036
rect 7267 1995 7325 1996
rect 9571 1995 9629 1996
rect 11203 1952 11261 1953
rect 2659 1912 2668 1952
rect 2708 1912 5548 1952
rect 5588 1912 5597 1952
rect 7363 1912 7372 1952
rect 7412 1912 7852 1952
rect 7892 1912 7901 1952
rect 8323 1912 8332 1952
rect 8372 1912 11212 1952
rect 11252 1912 11261 1952
rect 11320 1952 11360 1996
rect 25324 1953 25364 1996
rect 29827 1995 29885 1996
rect 14371 1952 14429 1953
rect 25315 1952 25373 1953
rect 11320 1912 14380 1952
rect 14420 1912 14429 1952
rect 14947 1912 14956 1952
rect 14996 1912 16204 1952
rect 16244 1912 16253 1952
rect 17539 1912 17548 1952
rect 17588 1912 17597 1952
rect 19363 1912 19372 1952
rect 19412 1912 20716 1952
rect 20756 1912 21388 1952
rect 21428 1912 21437 1952
rect 25230 1912 25324 1952
rect 25364 1912 25373 1952
rect 27331 1912 27340 1952
rect 27380 1912 27724 1952
rect 27764 1912 27773 1952
rect 28963 1912 28972 1952
rect 29012 1912 29260 1952
rect 29300 1912 29309 1952
rect 31555 1912 31564 1952
rect 31604 1912 32084 1952
rect 32995 1912 33004 1952
rect 33044 1912 33388 1952
rect 33428 1912 33437 1952
rect 35395 1912 35404 1952
rect 35444 1912 35692 1952
rect 35732 1912 35741 1952
rect 11203 1911 11261 1912
rect 14371 1911 14429 1912
rect 17548 1868 17588 1912
rect 25315 1911 25373 1912
rect 26467 1868 26525 1869
rect 30595 1868 30653 1869
rect 30979 1868 31037 1869
rect 5635 1828 5644 1868
rect 5684 1828 5932 1868
rect 5972 1828 5981 1868
rect 6115 1828 6124 1868
rect 6164 1828 6508 1868
rect 6548 1828 8428 1868
rect 8468 1828 8477 1868
rect 10339 1828 10348 1868
rect 10388 1828 17588 1868
rect 17731 1828 17740 1868
rect 17780 1828 17932 1868
rect 17972 1828 19412 1868
rect 20227 1828 20236 1868
rect 20276 1828 20908 1868
rect 20948 1828 21196 1868
rect 21236 1828 21245 1868
rect 26467 1828 26476 1868
rect 26516 1828 27244 1868
rect 27284 1828 27293 1868
rect 29443 1828 29452 1868
rect 29492 1828 30220 1868
rect 30260 1828 30269 1868
rect 30510 1828 30604 1868
rect 30644 1828 30653 1868
rect 30894 1828 30988 1868
rect 31028 1828 31037 1868
rect 0 1784 80 1804
rect 5932 1784 5972 1828
rect 18019 1784 18077 1785
rect 0 1744 2540 1784
rect 5932 1744 7948 1784
rect 7988 1744 10444 1784
rect 10484 1744 10493 1784
rect 14563 1744 14572 1784
rect 14612 1744 15628 1784
rect 15668 1744 16780 1784
rect 16820 1744 16829 1784
rect 17934 1744 18028 1784
rect 18068 1744 18077 1784
rect 0 1724 80 1744
rect 2500 1616 2540 1744
rect 18019 1743 18077 1744
rect 19372 1700 19412 1828
rect 26467 1827 26525 1828
rect 30595 1827 30653 1828
rect 30979 1827 31037 1828
rect 20323 1784 20381 1785
rect 32044 1784 32084 1912
rect 32611 1868 32669 1869
rect 33955 1868 34013 1869
rect 32515 1828 32524 1868
rect 32564 1828 32620 1868
rect 32660 1828 32669 1868
rect 32611 1827 32669 1828
rect 32740 1828 33772 1868
rect 33812 1828 33821 1868
rect 33955 1828 33964 1868
rect 34004 1828 35884 1868
rect 35924 1828 36172 1868
rect 36212 1828 36221 1868
rect 20323 1744 20332 1784
rect 20372 1744 28300 1784
rect 28340 1744 31756 1784
rect 31796 1744 31805 1784
rect 32044 1744 32332 1784
rect 32372 1744 32381 1784
rect 20323 1743 20381 1744
rect 20803 1700 20861 1701
rect 23971 1700 24029 1701
rect 32740 1700 32780 1828
rect 33955 1827 34013 1828
rect 42928 1784 43008 1804
rect 41059 1744 41068 1784
rect 41108 1744 43008 1784
rect 42928 1724 43008 1744
rect 3619 1660 3628 1700
rect 3668 1660 6796 1700
rect 6836 1660 6845 1700
rect 8332 1660 10156 1700
rect 10196 1660 10348 1700
rect 10388 1660 10397 1700
rect 10819 1660 10828 1700
rect 10868 1660 13036 1700
rect 13076 1660 13085 1700
rect 13219 1660 13228 1700
rect 13268 1660 19276 1700
rect 19316 1660 19325 1700
rect 19372 1660 19660 1700
rect 19700 1660 19709 1700
rect 20718 1660 20812 1700
rect 20852 1660 20861 1700
rect 23491 1660 23500 1700
rect 23540 1660 23692 1700
rect 23732 1660 23741 1700
rect 23875 1660 23884 1700
rect 23924 1660 23980 1700
rect 24020 1660 24029 1700
rect 25315 1660 25324 1700
rect 25364 1660 32428 1700
rect 32468 1660 32477 1700
rect 32611 1660 32620 1700
rect 32660 1660 32780 1700
rect 2500 1576 8140 1616
rect 8180 1576 8189 1616
rect 8332 1532 8372 1660
rect 20803 1659 20861 1660
rect 23971 1659 24029 1660
rect 10243 1576 10252 1616
rect 10292 1576 10540 1616
rect 10580 1576 10589 1616
rect 10723 1576 10732 1616
rect 10772 1576 11020 1616
rect 11060 1576 11069 1616
rect 11203 1576 11212 1616
rect 11252 1576 12940 1616
rect 12980 1576 12989 1616
rect 13315 1576 13324 1616
rect 13364 1576 17740 1616
rect 17780 1576 17789 1616
rect 17923 1576 17932 1616
rect 17972 1576 18508 1616
rect 18548 1576 20180 1616
rect 26755 1576 26764 1616
rect 26804 1576 37996 1616
rect 38036 1576 38045 1616
rect 20140 1532 20180 1576
rect 3679 1492 3688 1532
rect 3728 1492 3770 1532
rect 3810 1492 3852 1532
rect 3892 1492 3934 1532
rect 3974 1492 4016 1532
rect 4056 1492 4065 1532
rect 5443 1492 5452 1532
rect 5492 1492 8372 1532
rect 8419 1492 8428 1532
rect 8468 1492 10868 1532
rect 11683 1492 11692 1532
rect 11732 1492 17548 1532
rect 17588 1492 17597 1532
rect 18799 1492 18808 1532
rect 18848 1492 18890 1532
rect 18930 1492 18972 1532
rect 19012 1492 19054 1532
rect 19094 1492 19136 1532
rect 19176 1492 19185 1532
rect 20140 1492 28012 1532
rect 28052 1492 28061 1532
rect 28387 1492 28396 1532
rect 28436 1492 30028 1532
rect 30068 1492 30077 1532
rect 33919 1492 33928 1532
rect 33968 1492 34010 1532
rect 34050 1492 34092 1532
rect 34132 1492 34174 1532
rect 34214 1492 34256 1532
rect 34296 1492 34305 1532
rect 0 1448 80 1468
rect 10828 1448 10868 1492
rect 11203 1448 11261 1449
rect 14467 1448 14525 1449
rect 42928 1448 43008 1468
rect 0 1408 9140 1448
rect 10819 1408 10828 1448
rect 10868 1408 10877 1448
rect 11118 1408 11212 1448
rect 11252 1408 11261 1448
rect 11395 1408 11404 1448
rect 11444 1408 14476 1448
rect 14516 1408 14525 1448
rect 15715 1408 15724 1448
rect 15764 1408 18164 1448
rect 18595 1408 18604 1448
rect 18644 1408 20044 1448
rect 20084 1408 20093 1448
rect 20524 1408 27860 1448
rect 38947 1408 38956 1448
rect 38996 1408 43008 1448
rect 0 1388 80 1408
rect 9100 1281 9140 1408
rect 11203 1407 11261 1408
rect 14467 1407 14525 1408
rect 11587 1364 11645 1365
rect 18019 1364 18077 1365
rect 10531 1324 10540 1364
rect 10580 1324 11116 1364
rect 11156 1324 11165 1364
rect 11502 1324 11596 1364
rect 11636 1324 11645 1364
rect 11587 1323 11645 1324
rect 14668 1324 14996 1364
rect 16291 1324 16300 1364
rect 16340 1324 18028 1364
rect 18068 1324 18077 1364
rect 9091 1280 9149 1281
rect 14668 1280 14708 1324
rect 14851 1280 14909 1281
rect 9006 1240 9100 1280
rect 9140 1240 9149 1280
rect 10147 1240 10156 1280
rect 10196 1240 10924 1280
rect 10964 1240 11404 1280
rect 11444 1240 11453 1280
rect 12076 1240 14708 1280
rect 14766 1240 14860 1280
rect 14900 1240 14909 1280
rect 14956 1280 14996 1324
rect 18019 1323 18077 1324
rect 18124 1280 18164 1408
rect 18691 1364 18749 1365
rect 18691 1324 18700 1364
rect 18740 1324 18892 1364
rect 18932 1324 18941 1364
rect 19651 1324 19660 1364
rect 19700 1324 20180 1364
rect 18691 1323 18749 1324
rect 20140 1280 20180 1324
rect 20524 1280 20564 1408
rect 20611 1364 20669 1365
rect 20611 1324 20620 1364
rect 20660 1324 20812 1364
rect 20852 1324 20861 1364
rect 21004 1324 21332 1364
rect 21859 1324 21868 1364
rect 21908 1324 22156 1364
rect 22196 1324 22205 1364
rect 25603 1324 25612 1364
rect 25652 1324 26284 1364
rect 26324 1324 26333 1364
rect 26764 1324 26860 1364
rect 26900 1324 26909 1364
rect 20611 1323 20669 1324
rect 20707 1280 20765 1281
rect 14956 1240 15284 1280
rect 15331 1240 15340 1280
rect 15380 1240 16396 1280
rect 16436 1240 16445 1280
rect 18124 1240 19084 1280
rect 19124 1240 19133 1280
rect 20140 1240 20564 1280
rect 20622 1240 20716 1280
rect 20756 1240 20765 1280
rect 9091 1239 9149 1240
rect 12076 1196 12116 1240
rect 14851 1239 14909 1240
rect 15244 1196 15284 1240
rect 20707 1239 20765 1240
rect 16099 1196 16157 1197
rect 21004 1196 21044 1324
rect 21187 1280 21245 1281
rect 21102 1240 21196 1280
rect 21236 1240 21245 1280
rect 21292 1280 21332 1324
rect 26764 1280 26804 1324
rect 26947 1280 27005 1281
rect 21292 1240 23500 1280
rect 23540 1240 23549 1280
rect 23683 1240 23692 1280
rect 23732 1240 24076 1280
rect 24116 1240 24125 1280
rect 24259 1240 24268 1280
rect 24308 1240 25132 1280
rect 25172 1240 25181 1280
rect 25708 1240 26804 1280
rect 26862 1240 26956 1280
rect 26996 1240 27005 1280
rect 27820 1280 27860 1408
rect 42928 1388 43008 1408
rect 28195 1324 28204 1364
rect 28244 1324 31372 1364
rect 31412 1324 31421 1364
rect 32131 1324 32140 1364
rect 32180 1324 32620 1364
rect 32660 1324 32669 1364
rect 28204 1280 28244 1324
rect 27820 1240 28244 1280
rect 28960 1240 31660 1280
rect 31700 1240 31709 1280
rect 32035 1240 32044 1280
rect 32084 1240 33196 1280
rect 33236 1240 33245 1280
rect 34819 1240 34828 1280
rect 34868 1240 35308 1280
rect 35348 1240 35357 1280
rect 36451 1240 36460 1280
rect 36500 1240 36844 1280
rect 36884 1240 36893 1280
rect 40867 1240 40876 1280
rect 40916 1240 41644 1280
rect 41684 1240 41693 1280
rect 21187 1239 21245 1240
rect 4099 1156 4108 1196
rect 4148 1156 10732 1196
rect 10772 1156 10781 1196
rect 11320 1156 12116 1196
rect 12163 1156 12172 1196
rect 12212 1156 15148 1196
rect 15188 1156 15197 1196
rect 15244 1156 16108 1196
rect 16148 1156 16157 1196
rect 17731 1156 17740 1196
rect 17780 1156 20140 1196
rect 20180 1156 20189 1196
rect 20236 1156 21044 1196
rect 21091 1156 21100 1196
rect 21140 1156 21772 1196
rect 21812 1156 21821 1196
rect 22915 1156 22924 1196
rect 22964 1156 23308 1196
rect 23348 1156 23357 1196
rect 0 1112 80 1132
rect 1219 1112 1277 1113
rect 10732 1112 10772 1156
rect 11320 1112 11360 1156
rect 16099 1155 16157 1156
rect 12355 1112 12413 1113
rect 17347 1112 17405 1113
rect 20236 1112 20276 1156
rect 21955 1112 22013 1113
rect 0 1072 1228 1112
rect 1268 1072 1277 1112
rect 2563 1072 2572 1112
rect 2612 1072 3436 1112
rect 3476 1072 4300 1112
rect 4340 1072 5068 1112
rect 5108 1072 5117 1112
rect 6307 1072 6316 1112
rect 6356 1072 10156 1112
rect 10196 1072 10205 1112
rect 10732 1072 11360 1112
rect 12270 1072 12364 1112
rect 12404 1072 12413 1112
rect 15235 1072 15244 1112
rect 15284 1072 17356 1112
rect 17396 1072 17405 1112
rect 18979 1072 18988 1112
rect 19028 1072 20276 1112
rect 20323 1072 20332 1112
rect 20372 1072 21964 1112
rect 22004 1072 22013 1112
rect 23500 1112 23540 1240
rect 24451 1196 24509 1197
rect 25708 1196 25748 1240
rect 26947 1239 27005 1240
rect 24451 1156 24460 1196
rect 24500 1156 24748 1196
rect 24788 1156 25708 1196
rect 25748 1156 25757 1196
rect 26083 1156 26092 1196
rect 26132 1156 27340 1196
rect 27380 1156 27389 1196
rect 24451 1155 24509 1156
rect 28960 1112 29000 1240
rect 40291 1196 40349 1197
rect 41251 1196 41309 1197
rect 30700 1156 38572 1196
rect 38612 1156 39532 1196
rect 39572 1156 39581 1196
rect 40291 1156 40300 1196
rect 40340 1156 40492 1196
rect 40532 1156 40541 1196
rect 41166 1156 41260 1196
rect 41300 1156 41309 1196
rect 29155 1112 29213 1113
rect 30700 1112 30740 1156
rect 40291 1155 40349 1156
rect 41251 1155 41309 1156
rect 34627 1112 34685 1113
rect 42928 1112 43008 1132
rect 23500 1072 29000 1112
rect 29070 1072 29164 1112
rect 29204 1072 30740 1112
rect 32740 1072 33484 1112
rect 33524 1072 33533 1112
rect 34542 1072 34636 1112
rect 34676 1072 34685 1112
rect 36259 1072 36268 1112
rect 36308 1072 39724 1112
rect 39764 1072 39773 1112
rect 40291 1072 40300 1112
rect 40340 1072 43008 1112
rect 0 1052 80 1072
rect 1219 1071 1277 1072
rect 12355 1071 12413 1072
rect 15244 1028 15284 1072
rect 17347 1071 17405 1072
rect 21955 1071 22013 1072
rect 29155 1071 29213 1072
rect 4483 988 4492 1028
rect 4532 988 5260 1028
rect 5300 988 5309 1028
rect 6028 988 15284 1028
rect 18883 1028 18941 1029
rect 32740 1028 32780 1072
rect 34627 1071 34685 1072
rect 18883 988 18892 1028
rect 18932 988 21620 1028
rect 21667 988 21676 1028
rect 21716 988 22156 1028
rect 22196 988 22205 1028
rect 22924 988 28492 1028
rect 28532 988 28541 1028
rect 29347 988 29356 1028
rect 29396 988 30028 1028
rect 30068 988 30508 1028
rect 30548 988 30557 1028
rect 30892 988 32780 1028
rect 34636 1028 34676 1071
rect 42928 1052 43008 1072
rect 34636 988 40876 1028
rect 40916 988 40925 1028
rect 6028 944 6068 988
rect 18883 987 18941 988
rect 6979 944 7037 945
rect 15619 944 15677 945
rect 20515 944 20573 945
rect 1315 904 1324 944
rect 1364 904 6068 944
rect 6894 904 6988 944
rect 7028 904 7037 944
rect 10339 904 10348 944
rect 10388 904 13612 944
rect 13652 904 14668 944
rect 14708 904 14717 944
rect 15534 904 15628 944
rect 15668 904 15677 944
rect 18403 904 18412 944
rect 18452 904 18700 944
rect 18740 904 18749 944
rect 19267 904 19276 944
rect 19316 904 20524 944
rect 20564 904 20573 944
rect 21580 944 21620 988
rect 22924 944 22964 988
rect 30892 944 30932 988
rect 21580 904 22964 944
rect 23107 904 23116 944
rect 23156 904 23692 944
rect 23732 904 23741 944
rect 24547 904 24556 944
rect 24596 904 24844 944
rect 24884 904 24893 944
rect 27427 904 27436 944
rect 27476 904 27916 944
rect 27956 904 27965 944
rect 28675 904 28684 944
rect 28724 904 29260 944
rect 29300 904 29309 944
rect 29356 904 30932 944
rect 31276 904 36268 944
rect 36308 904 36317 944
rect 36931 904 36940 944
rect 36980 904 38284 944
rect 38324 904 38333 944
rect 6979 903 7037 904
rect 15619 903 15677 904
rect 20515 903 20573 904
rect 29356 860 29396 904
rect 13027 820 13036 860
rect 13076 820 19660 860
rect 19700 820 19709 860
rect 25027 820 25036 860
rect 25076 820 26668 860
rect 26708 820 26717 860
rect 28960 820 29396 860
rect 30691 820 30700 860
rect 30740 820 30988 860
rect 31028 820 31037 860
rect 0 776 80 796
rect 17635 776 17693 777
rect 20611 776 20669 777
rect 28960 776 29000 820
rect 30787 776 30845 777
rect 31171 776 31229 777
rect 0 736 212 776
rect 4919 736 4928 776
rect 4968 736 5010 776
rect 5050 736 5092 776
rect 5132 736 5174 776
rect 5214 736 5256 776
rect 5296 736 5305 776
rect 11875 736 11884 776
rect 11924 736 16492 776
rect 16532 736 17644 776
rect 17684 736 17693 776
rect 20039 736 20048 776
rect 20088 736 20130 776
rect 20170 736 20212 776
rect 20252 736 20294 776
rect 20334 736 20376 776
rect 20416 736 20425 776
rect 20526 736 20620 776
rect 20660 736 20669 776
rect 0 716 80 736
rect 172 608 212 736
rect 17635 735 17693 736
rect 20611 735 20669 736
rect 20716 736 25228 776
rect 25268 736 25277 776
rect 26563 736 26572 776
rect 26612 736 29000 776
rect 30702 736 30796 776
rect 30836 736 30845 776
rect 31086 736 31180 776
rect 31220 736 31229 776
rect 20716 692 20756 736
rect 30787 735 30845 736
rect 31171 735 31229 736
rect 31276 692 31316 904
rect 31651 820 31660 860
rect 31700 820 37900 860
rect 37940 820 40108 860
rect 40148 820 40157 860
rect 42928 776 43008 796
rect 32899 736 32908 776
rect 32948 736 33292 776
rect 33332 736 33341 776
rect 35159 736 35168 776
rect 35208 736 35250 776
rect 35290 736 35332 776
rect 35372 736 35414 776
rect 35454 736 35496 776
rect 35536 736 35545 776
rect 40291 736 40300 776
rect 40340 736 43008 776
rect 42928 716 43008 736
rect 33091 692 33149 693
rect 15811 652 15820 692
rect 15860 652 20756 692
rect 27043 652 27052 692
rect 27092 652 31316 692
rect 32323 652 32332 692
rect 32372 652 33100 692
rect 33140 652 33149 692
rect 35011 652 35020 692
rect 35060 652 36652 692
rect 36692 652 36701 692
rect 33091 651 33149 652
rect 172 568 18988 608
rect 19028 568 19037 608
rect 19843 568 19852 608
rect 19892 568 24172 608
rect 24212 568 24221 608
rect 31939 568 31948 608
rect 31988 568 32716 608
rect 32756 568 32765 608
rect 20707 524 20765 525
rect 20707 484 20716 524
rect 20756 484 27052 524
rect 27092 484 27101 524
rect 20707 483 20765 484
rect 0 440 80 460
rect 23875 440 23933 441
rect 42928 440 43008 460
rect 0 400 1324 440
rect 1364 400 1373 440
rect 16195 400 16204 440
rect 16244 400 23884 440
rect 23924 400 23933 440
rect 28099 400 28108 440
rect 28148 400 35596 440
rect 35636 400 35645 440
rect 40675 400 40684 440
rect 40724 400 43008 440
rect 0 380 80 400
rect 23875 399 23933 400
rect 42928 380 43008 400
rect 20803 356 20861 357
rect 14659 316 14668 356
rect 14708 316 20812 356
rect 20852 316 20861 356
rect 22531 316 22540 356
rect 22580 316 23980 356
rect 24020 316 24029 356
rect 28675 316 28684 356
rect 28724 316 37516 356
rect 37556 316 37565 356
rect 20803 315 20861 316
rect 14371 232 14380 272
rect 14420 232 16012 272
rect 16052 232 16061 272
rect 25603 232 25612 272
rect 25652 232 34444 272
rect 34484 232 34493 272
rect 32707 188 32765 189
rect 20227 148 20236 188
rect 20276 148 30892 188
rect 30932 148 30941 188
rect 32622 148 32716 188
rect 32756 148 32765 188
rect 32707 147 32765 148
rect 0 104 80 124
rect 19267 104 19325 105
rect 42928 104 43008 124
rect 0 64 4108 104
rect 4148 64 4157 104
rect 9475 64 9484 104
rect 9524 64 19276 104
rect 19316 64 19325 104
rect 28291 64 28300 104
rect 28340 64 39724 104
rect 39764 64 39773 104
rect 41443 64 41452 104
rect 41492 64 43008 104
rect 0 44 80 64
rect 19267 63 19325 64
rect 42928 44 43008 64
<< via3 >>
rect 268 10480 308 10520
rect 4928 9808 4968 9848
rect 5010 9808 5050 9848
rect 5092 9808 5132 9848
rect 5174 9808 5214 9848
rect 5256 9808 5296 9848
rect 20048 9808 20088 9848
rect 20130 9808 20170 9848
rect 20212 9808 20252 9848
rect 20294 9808 20334 9848
rect 20376 9808 20416 9848
rect 35168 9808 35208 9848
rect 35250 9808 35290 9848
rect 35332 9808 35372 9848
rect 35414 9808 35454 9848
rect 35496 9808 35536 9848
rect 1228 9472 1268 9512
rect 10060 9472 10100 9512
rect 15244 9388 15284 9428
rect 30796 9388 30836 9428
rect 4300 9304 4340 9344
rect 3688 9052 3728 9092
rect 3770 9052 3810 9092
rect 3852 9052 3892 9092
rect 3934 9052 3974 9092
rect 4016 9052 4056 9092
rect 18808 9052 18848 9092
rect 18890 9052 18930 9092
rect 18972 9052 19012 9092
rect 19054 9052 19094 9092
rect 19136 9052 19176 9092
rect 33928 9052 33968 9092
rect 34010 9052 34050 9092
rect 34092 9052 34132 9092
rect 34174 9052 34214 9092
rect 34256 9052 34296 9092
rect 31180 8968 31220 9008
rect 12460 8716 12500 8756
rect 39820 8716 39860 8756
rect 6412 8632 6452 8672
rect 8044 8632 8084 8672
rect 15916 8632 15956 8672
rect 30028 8632 30068 8672
rect 14092 8548 14132 8588
rect 24364 8548 24404 8588
rect 27820 8548 27860 8588
rect 4780 8464 4820 8504
rect 22348 8464 22388 8504
rect 23788 8464 23828 8504
rect 25420 8464 25460 8504
rect 4928 8296 4968 8336
rect 5010 8296 5050 8336
rect 5092 8296 5132 8336
rect 5174 8296 5214 8336
rect 5256 8296 5296 8336
rect 20048 8296 20088 8336
rect 20130 8296 20170 8336
rect 20212 8296 20252 8336
rect 20294 8296 20334 8336
rect 20376 8296 20416 8336
rect 35168 8296 35208 8336
rect 35250 8296 35290 8336
rect 35332 8296 35372 8336
rect 35414 8296 35454 8336
rect 35496 8296 35536 8336
rect 9100 7960 9140 8000
rect 13804 7960 13844 8000
rect 17644 7960 17684 8000
rect 27724 7876 27764 7916
rect 33100 7876 33140 7916
rect 3688 7540 3728 7580
rect 3770 7540 3810 7580
rect 3852 7540 3892 7580
rect 3934 7540 3974 7580
rect 4016 7540 4056 7580
rect 9292 7540 9332 7580
rect 13804 7540 13844 7580
rect 18808 7540 18848 7580
rect 18890 7540 18930 7580
rect 18972 7540 19012 7580
rect 19054 7540 19094 7580
rect 19136 7540 19176 7580
rect 33928 7540 33968 7580
rect 34010 7540 34050 7580
rect 34092 7540 34132 7580
rect 34174 7540 34214 7580
rect 34256 7540 34296 7580
rect 5356 7456 5396 7496
rect 5452 7204 5492 7244
rect 28876 7204 28916 7244
rect 16396 7120 16436 7160
rect 19372 7120 19412 7160
rect 24172 7120 24212 7160
rect 25420 7120 25460 7160
rect 27628 7120 27668 7160
rect 31660 7036 31700 7076
rect 12172 6952 12212 6992
rect 4204 6868 4244 6908
rect 4928 6784 4968 6824
rect 5010 6784 5050 6824
rect 5092 6784 5132 6824
rect 5174 6784 5214 6824
rect 5256 6784 5296 6824
rect 20048 6784 20088 6824
rect 20130 6784 20170 6824
rect 20212 6784 20252 6824
rect 20294 6784 20334 6824
rect 20376 6784 20416 6824
rect 35168 6784 35208 6824
rect 35250 6784 35290 6824
rect 35332 6784 35372 6824
rect 35414 6784 35454 6824
rect 35496 6784 35536 6824
rect 9292 6700 9332 6740
rect 5740 6616 5780 6656
rect 19852 6532 19892 6572
rect 1708 6448 1748 6488
rect 4300 6448 4340 6488
rect 5356 6448 5396 6488
rect 14764 6448 14804 6488
rect 25324 6448 25364 6488
rect 27724 6448 27764 6488
rect 18700 6364 18740 6404
rect 31756 6364 31796 6404
rect 5548 6280 5588 6320
rect 17932 6280 17972 6320
rect 39628 6280 39668 6320
rect 4396 6196 4436 6236
rect 5740 6196 5780 6236
rect 5644 6112 5684 6152
rect 3688 6028 3728 6068
rect 3770 6028 3810 6068
rect 3852 6028 3892 6068
rect 3934 6028 3974 6068
rect 4016 6028 4056 6068
rect 18808 6028 18848 6068
rect 18890 6028 18930 6068
rect 18972 6028 19012 6068
rect 19054 6028 19094 6068
rect 19136 6028 19176 6068
rect 21388 6028 21428 6068
rect 33928 6028 33968 6068
rect 34010 6028 34050 6068
rect 34092 6028 34132 6068
rect 34174 6028 34214 6068
rect 34256 6028 34296 6068
rect 30124 5944 30164 5984
rect 31756 5944 31796 5984
rect 5548 5860 5588 5900
rect 19372 5692 19412 5732
rect 22060 5692 22100 5732
rect 8428 5608 8468 5648
rect 16396 5608 16436 5648
rect 4780 5524 4820 5564
rect 5356 5524 5396 5564
rect 32620 5524 32660 5564
rect 11788 5440 11828 5480
rect 10060 5356 10100 5396
rect 3532 5272 3572 5312
rect 4928 5272 4968 5312
rect 5010 5272 5050 5312
rect 5092 5272 5132 5312
rect 5174 5272 5214 5312
rect 5256 5272 5296 5312
rect 5644 5272 5684 5312
rect 20048 5272 20088 5312
rect 20130 5272 20170 5312
rect 20212 5272 20252 5312
rect 20294 5272 20334 5312
rect 20376 5272 20416 5312
rect 20620 5272 20660 5312
rect 30124 5272 30164 5312
rect 35168 5272 35208 5312
rect 35250 5272 35290 5312
rect 35332 5272 35372 5312
rect 35414 5272 35454 5312
rect 35496 5272 35536 5312
rect 21004 5188 21044 5228
rect 3724 5104 3764 5144
rect 4108 5104 4148 5144
rect 23980 5020 24020 5060
rect 1612 4936 1652 4976
rect 22636 4936 22676 4976
rect 26380 4936 26420 4976
rect 30220 4936 30260 4976
rect 19276 4852 19316 4892
rect 23884 4852 23924 4892
rect 27244 4852 27284 4892
rect 5356 4684 5396 4724
rect 3688 4516 3728 4556
rect 3770 4516 3810 4556
rect 3852 4516 3892 4556
rect 3934 4516 3974 4556
rect 4016 4516 4056 4556
rect 1228 4432 1268 4472
rect 5452 4432 5492 4472
rect 26380 4684 26420 4724
rect 11596 4600 11636 4640
rect 18808 4516 18848 4556
rect 18890 4516 18930 4556
rect 18972 4516 19012 4556
rect 19054 4516 19094 4556
rect 19136 4516 19176 4556
rect 33928 4516 33968 4556
rect 34010 4516 34050 4556
rect 34092 4516 34132 4556
rect 34174 4516 34214 4556
rect 34256 4516 34296 4556
rect 4300 4348 4340 4388
rect 23788 4348 23828 4388
rect 25708 4180 25748 4220
rect 4396 4096 4436 4136
rect 12076 4096 12116 4136
rect 19372 4096 19412 4136
rect 31756 4096 31796 4136
rect 34828 4096 34868 4136
rect 10444 4012 10484 4052
rect 4108 3844 4148 3884
rect 3244 3760 3284 3800
rect 4928 3760 4968 3800
rect 5010 3760 5050 3800
rect 5092 3760 5132 3800
rect 5174 3760 5214 3800
rect 5256 3760 5296 3800
rect 14188 4012 14228 4052
rect 15244 4012 15284 4052
rect 19660 3844 19700 3884
rect 20048 3760 20088 3800
rect 20130 3760 20170 3800
rect 20212 3760 20252 3800
rect 20294 3760 20334 3800
rect 20376 3760 20416 3800
rect 21196 3760 21236 3800
rect 35168 3760 35208 3800
rect 35250 3760 35290 3800
rect 35332 3760 35372 3800
rect 35414 3760 35454 3800
rect 35496 3760 35536 3800
rect 22636 3676 22676 3716
rect 11212 3592 11252 3632
rect 32716 3592 32756 3632
rect 12172 3508 12212 3548
rect 39532 3508 39572 3548
rect 1612 3424 1652 3464
rect 14188 3424 14228 3464
rect 16396 3424 16436 3464
rect 21004 3424 21044 3464
rect 21484 3424 21524 3464
rect 22636 3424 22676 3464
rect 23788 3424 23828 3464
rect 24460 3424 24500 3464
rect 31852 3424 31892 3464
rect 34444 3424 34484 3464
rect 38092 3424 38132 3464
rect 12364 3340 12404 3380
rect 21964 3340 22004 3380
rect 38092 3256 38132 3296
rect 18892 3172 18932 3212
rect 27244 3088 27284 3128
rect 30220 3088 30260 3128
rect 32620 3088 32660 3128
rect 37324 3088 37364 3128
rect 3244 3004 3284 3044
rect 3688 3004 3728 3044
rect 3770 3004 3810 3044
rect 3852 3004 3892 3044
rect 3934 3004 3974 3044
rect 4016 3004 4056 3044
rect 18808 3004 18848 3044
rect 18890 3004 18930 3044
rect 18972 3004 19012 3044
rect 19054 3004 19094 3044
rect 19136 3004 19176 3044
rect 20044 3004 20084 3044
rect 33928 3004 33968 3044
rect 34010 3004 34050 3044
rect 34092 3004 34132 3044
rect 34174 3004 34214 3044
rect 34256 3004 34296 3044
rect 4780 2836 4820 2876
rect 15436 2836 15476 2876
rect 4204 2752 4244 2792
rect 18124 2752 18164 2792
rect 3532 2668 3572 2708
rect 10444 2668 10484 2708
rect 5932 2584 5972 2624
rect 16108 2584 16148 2624
rect 20236 2584 20276 2624
rect 28684 2584 28724 2624
rect 8044 2332 8084 2372
rect 15148 2332 15188 2372
rect 20332 2416 20372 2456
rect 30604 2500 30644 2540
rect 15340 2332 15380 2372
rect 4928 2248 4968 2288
rect 5010 2248 5050 2288
rect 5092 2248 5132 2288
rect 5174 2248 5214 2288
rect 5256 2248 5296 2288
rect 11596 2248 11636 2288
rect 19948 2248 19988 2288
rect 20048 2248 20088 2288
rect 20130 2248 20170 2288
rect 20212 2248 20252 2288
rect 20294 2248 20334 2288
rect 20376 2248 20416 2288
rect 23980 2248 24020 2288
rect 35168 2248 35208 2288
rect 35250 2248 35290 2288
rect 35332 2248 35372 2288
rect 35414 2248 35454 2288
rect 35496 2248 35536 2288
rect 15436 2164 15476 2204
rect 7276 1996 7316 2036
rect 9580 1996 9620 2036
rect 29836 1996 29876 2036
rect 11212 1912 11252 1952
rect 14380 1912 14420 1952
rect 25324 1912 25364 1952
rect 26476 1828 26516 1868
rect 30604 1828 30644 1868
rect 30988 1828 31028 1868
rect 18028 1744 18068 1784
rect 32620 1828 32660 1868
rect 33964 1828 34004 1868
rect 20332 1744 20372 1784
rect 20812 1660 20852 1700
rect 23980 1660 24020 1700
rect 3688 1492 3728 1532
rect 3770 1492 3810 1532
rect 3852 1492 3892 1532
rect 3934 1492 3974 1532
rect 4016 1492 4056 1532
rect 18808 1492 18848 1532
rect 18890 1492 18930 1532
rect 18972 1492 19012 1532
rect 19054 1492 19094 1532
rect 19136 1492 19176 1532
rect 33928 1492 33968 1532
rect 34010 1492 34050 1532
rect 34092 1492 34132 1532
rect 34174 1492 34214 1532
rect 34256 1492 34296 1532
rect 11212 1408 11252 1448
rect 14476 1408 14516 1448
rect 11596 1324 11636 1364
rect 18028 1324 18068 1364
rect 9100 1240 9140 1280
rect 14860 1240 14900 1280
rect 18700 1324 18740 1364
rect 20620 1324 20660 1364
rect 20716 1240 20756 1280
rect 21196 1240 21236 1280
rect 26956 1240 26996 1280
rect 16108 1156 16148 1196
rect 1228 1072 1268 1112
rect 12364 1072 12404 1112
rect 17356 1072 17396 1112
rect 21964 1072 22004 1112
rect 24460 1156 24500 1196
rect 40300 1156 40340 1196
rect 41260 1156 41300 1196
rect 29164 1072 29204 1112
rect 34636 1072 34676 1112
rect 18892 988 18932 1028
rect 6988 904 7028 944
rect 15628 904 15668 944
rect 20524 904 20564 944
rect 4928 736 4968 776
rect 5010 736 5050 776
rect 5092 736 5132 776
rect 5174 736 5214 776
rect 5256 736 5296 776
rect 17644 736 17684 776
rect 20048 736 20088 776
rect 20130 736 20170 776
rect 20212 736 20252 776
rect 20294 736 20334 776
rect 20376 736 20416 776
rect 20620 736 20660 776
rect 30796 736 30836 776
rect 31180 736 31220 776
rect 35168 736 35208 776
rect 35250 736 35290 776
rect 35332 736 35372 776
rect 35414 736 35454 776
rect 35496 736 35536 776
rect 33100 652 33140 692
rect 20716 484 20756 524
rect 23884 400 23924 440
rect 20812 316 20852 356
rect 32716 148 32756 188
rect 19276 64 19316 104
<< metal4 >>
rect 268 10520 308 10529
rect 268 8597 308 10480
rect 4928 9848 5296 9857
rect 4968 9808 5010 9848
rect 5050 9808 5092 9848
rect 5132 9808 5174 9848
rect 5214 9808 5256 9848
rect 4928 9799 5296 9808
rect 20048 9848 20416 9857
rect 20088 9808 20130 9848
rect 20170 9808 20212 9848
rect 20252 9808 20294 9848
rect 20334 9808 20376 9848
rect 20048 9799 20416 9808
rect 35168 9848 35536 9857
rect 35208 9808 35250 9848
rect 35290 9808 35332 9848
rect 35372 9808 35414 9848
rect 35454 9808 35496 9848
rect 35168 9799 35536 9808
rect 1228 9512 1268 9521
rect 1228 8681 1268 9472
rect 10060 9512 10100 9521
rect 4300 9344 4340 9353
rect 3688 9092 4056 9101
rect 3728 9052 3770 9092
rect 3810 9052 3852 9092
rect 3892 9052 3934 9092
rect 3974 9052 4016 9092
rect 3688 9043 4056 9052
rect 1227 8672 1269 8681
rect 1227 8632 1228 8672
rect 1268 8632 1269 8672
rect 1227 8623 1269 8632
rect 267 8588 309 8597
rect 267 8548 268 8588
rect 308 8548 309 8588
rect 267 8539 309 8548
rect 3688 7580 4056 7589
rect 3728 7540 3770 7580
rect 3810 7540 3852 7580
rect 3892 7540 3934 7580
rect 3974 7540 4016 7580
rect 3688 7531 4056 7540
rect 4204 6908 4244 6917
rect 1707 6488 1749 6497
rect 1707 6448 1708 6488
rect 1748 6448 1749 6488
rect 1707 6439 1749 6448
rect 1708 6354 1748 6439
rect 3688 6068 4056 6077
rect 3728 6028 3770 6068
rect 3810 6028 3852 6068
rect 3892 6028 3934 6068
rect 3974 6028 4016 6068
rect 3688 6019 4056 6028
rect 3532 5312 3572 5321
rect 1611 4976 1653 4985
rect 1611 4936 1612 4976
rect 1652 4936 1653 4976
rect 1611 4927 1653 4936
rect 1612 4842 1652 4927
rect 1228 4472 1268 4483
rect 1228 4397 1268 4432
rect 1227 4388 1269 4397
rect 1227 4348 1228 4388
rect 1268 4348 1269 4388
rect 1227 4339 1269 4348
rect 3244 3800 3284 3809
rect 1611 3464 1653 3473
rect 1611 3424 1612 3464
rect 1652 3424 1653 3464
rect 1611 3415 1653 3424
rect 1612 3330 1652 3415
rect 3244 3044 3284 3760
rect 3244 2995 3284 3004
rect 3532 2708 3572 5272
rect 3724 5144 3764 5155
rect 3724 5069 3764 5104
rect 4108 5144 4148 5153
rect 3723 5060 3765 5069
rect 3723 5020 3724 5060
rect 3764 5020 3765 5060
rect 3723 5011 3765 5020
rect 3688 4556 4056 4565
rect 3728 4516 3770 4556
rect 3810 4516 3852 4556
rect 3892 4516 3934 4556
rect 3974 4516 4016 4556
rect 3688 4507 4056 4516
rect 4108 3884 4148 5104
rect 4108 3835 4148 3844
rect 3688 3044 4056 3053
rect 3728 3004 3770 3044
rect 3810 3004 3852 3044
rect 3892 3004 3934 3044
rect 3974 3004 4016 3044
rect 3688 2995 4056 3004
rect 4204 2792 4244 6868
rect 4300 6488 4340 9304
rect 4779 8672 4821 8681
rect 4779 8632 4780 8672
rect 4820 8632 4821 8672
rect 4779 8623 4821 8632
rect 6412 8672 6452 8683
rect 4780 8504 4820 8623
rect 6412 8597 6452 8632
rect 8044 8672 8084 8681
rect 6411 8588 6453 8597
rect 6411 8548 6412 8588
rect 6452 8548 6453 8588
rect 6411 8539 6453 8548
rect 4780 8455 4820 8464
rect 4928 8336 5296 8345
rect 4968 8296 5010 8336
rect 5050 8296 5092 8336
rect 5132 8296 5174 8336
rect 5214 8296 5256 8336
rect 4928 8287 5296 8296
rect 5356 7496 5396 7505
rect 4928 6824 5296 6833
rect 4968 6784 5010 6824
rect 5050 6784 5092 6824
rect 5132 6784 5174 6824
rect 5214 6784 5256 6824
rect 4928 6775 5296 6784
rect 4300 4388 4340 6448
rect 5356 6488 5396 7456
rect 5356 6439 5396 6448
rect 5452 7244 5492 7253
rect 4300 4339 4340 4348
rect 4396 6236 4436 6245
rect 4396 4136 4436 6196
rect 4396 4087 4436 4096
rect 4780 5564 4820 5573
rect 4780 2876 4820 5524
rect 5356 5564 5396 5573
rect 4928 5312 5296 5321
rect 4968 5272 5010 5312
rect 5050 5272 5092 5312
rect 5132 5272 5174 5312
rect 5214 5272 5256 5312
rect 4928 5263 5296 5272
rect 5356 4724 5396 5524
rect 5356 4675 5396 4684
rect 5452 4472 5492 7204
rect 5740 6656 5780 6665
rect 5548 6320 5588 6329
rect 5548 5900 5588 6280
rect 5740 6236 5780 6616
rect 5740 6187 5780 6196
rect 5548 5851 5588 5860
rect 5644 6152 5684 6161
rect 5644 5312 5684 6112
rect 8044 5573 8084 8632
rect 9099 8000 9141 8009
rect 9099 7960 9100 8000
rect 9140 7960 9141 8000
rect 9099 7951 9141 7960
rect 9100 7866 9140 7951
rect 9292 7580 9332 7589
rect 9292 6740 9332 7540
rect 10060 7253 10100 9472
rect 15244 9428 15284 9437
rect 12459 8756 12501 8765
rect 12459 8716 12460 8756
rect 12500 8716 12501 8756
rect 12459 8707 12501 8716
rect 12460 8622 12500 8707
rect 15244 8681 15284 9388
rect 30796 9428 30836 9437
rect 18808 9092 19176 9101
rect 18848 9052 18890 9092
rect 18930 9052 18972 9092
rect 19012 9052 19054 9092
rect 19094 9052 19136 9092
rect 18808 9043 19176 9052
rect 22347 8756 22389 8765
rect 22347 8716 22348 8756
rect 22388 8716 22389 8756
rect 22347 8707 22389 8716
rect 15243 8672 15285 8681
rect 15243 8632 15244 8672
rect 15284 8632 15285 8672
rect 15243 8623 15285 8632
rect 15916 8672 15956 8683
rect 14092 8588 14132 8597
rect 13803 8000 13845 8009
rect 13803 7960 13804 8000
rect 13844 7960 13845 8000
rect 13803 7951 13845 7960
rect 13804 7580 13844 7951
rect 13804 7531 13844 7540
rect 10059 7244 10101 7253
rect 10059 7204 10060 7244
rect 10100 7204 10101 7244
rect 10059 7195 10101 7204
rect 9292 6691 9332 6700
rect 8427 5648 8469 5657
rect 8427 5608 8428 5648
rect 8468 5608 8469 5648
rect 8427 5599 8469 5608
rect 8043 5564 8085 5573
rect 8043 5524 8044 5564
rect 8084 5524 8085 5564
rect 8043 5515 8085 5524
rect 5644 5263 5684 5272
rect 5452 4423 5492 4432
rect 4928 3800 5296 3809
rect 4968 3760 5010 3800
rect 5050 3760 5092 3800
rect 5132 3760 5174 3800
rect 5214 3760 5256 3800
rect 4928 3751 5296 3760
rect 4780 2827 4820 2836
rect 4204 2743 4244 2752
rect 3532 2659 3572 2668
rect 5932 2633 5972 2718
rect 5931 2624 5973 2633
rect 5931 2584 5932 2624
rect 5972 2584 5973 2624
rect 5931 2575 5973 2584
rect 8044 2372 8084 5515
rect 8428 5514 8468 5599
rect 10060 5396 10100 7195
rect 14092 7085 14132 8548
rect 14091 7076 14133 7085
rect 14091 7036 14092 7076
rect 14132 7036 14133 7076
rect 14091 7027 14133 7036
rect 12172 6992 12212 7001
rect 11787 5480 11829 5489
rect 11787 5440 11788 5480
rect 11828 5440 11829 5480
rect 11787 5431 11829 5440
rect 10060 5347 10100 5356
rect 11788 5346 11828 5431
rect 11596 4640 11636 4649
rect 10444 4052 10484 4061
rect 10444 3473 10484 4012
rect 11212 3632 11252 3641
rect 10443 3464 10485 3473
rect 10443 3424 10444 3464
rect 10484 3424 10485 3464
rect 10443 3415 10485 3424
rect 10444 2708 10484 3415
rect 10444 2659 10484 2668
rect 8044 2323 8084 2332
rect 4928 2288 5296 2297
rect 4968 2248 5010 2288
rect 5050 2248 5092 2288
rect 5132 2248 5174 2288
rect 5214 2248 5256 2288
rect 4928 2239 5296 2248
rect 7275 2036 7317 2045
rect 7275 1996 7276 2036
rect 7316 1996 7317 2036
rect 7275 1987 7317 1996
rect 9579 2036 9621 2045
rect 9579 1996 9580 2036
rect 9620 1996 9621 2036
rect 9579 1987 9621 1996
rect 7276 1902 7316 1987
rect 9580 1902 9620 1987
rect 11212 1952 11252 3592
rect 3688 1532 4056 1541
rect 3728 1492 3770 1532
rect 3810 1492 3852 1532
rect 3892 1492 3934 1532
rect 3974 1492 4016 1532
rect 3688 1483 4056 1492
rect 11212 1448 11252 1912
rect 11212 1399 11252 1408
rect 11596 2288 11636 4600
rect 12075 4136 12117 4145
rect 12075 4096 12076 4136
rect 12116 4096 12117 4136
rect 12075 4087 12117 4096
rect 12076 4002 12116 4087
rect 12172 3548 12212 6952
rect 14092 4145 14132 7027
rect 14763 6488 14805 6497
rect 14763 6448 14764 6488
rect 14804 6448 14805 6488
rect 14763 6439 14805 6448
rect 14764 6354 14804 6439
rect 14187 4388 14229 4397
rect 14187 4348 14188 4388
rect 14228 4348 14229 4388
rect 14187 4339 14229 4348
rect 14091 4136 14133 4145
rect 14091 4096 14092 4136
rect 14132 4096 14133 4136
rect 14091 4087 14133 4096
rect 12172 3499 12212 3508
rect 14188 4052 14228 4339
rect 12363 3464 12405 3473
rect 12363 3424 12364 3464
rect 12404 3424 12405 3464
rect 12363 3415 12405 3424
rect 14188 3464 14228 4012
rect 15244 4052 15284 8623
rect 15916 8597 15956 8632
rect 15915 8588 15957 8597
rect 15915 8548 15916 8588
rect 15956 8548 15957 8588
rect 15915 8539 15957 8548
rect 22348 8504 22388 8707
rect 30027 8672 30069 8681
rect 30027 8632 30028 8672
rect 30068 8632 30069 8672
rect 30027 8623 30069 8632
rect 24363 8588 24405 8597
rect 24363 8548 24364 8588
rect 24404 8548 24405 8588
rect 24363 8539 24405 8548
rect 27820 8588 27860 8597
rect 22348 8455 22388 8464
rect 23788 8504 23828 8513
rect 20048 8336 20416 8345
rect 20088 8296 20130 8336
rect 20170 8296 20212 8336
rect 20252 8296 20294 8336
rect 20334 8296 20376 8336
rect 20048 8287 20416 8296
rect 17644 8000 17684 8009
rect 16396 7160 16436 7169
rect 16396 7001 16436 7120
rect 16395 6992 16437 7001
rect 16395 6952 16396 6992
rect 16436 6952 16437 6992
rect 16395 6943 16437 6952
rect 16395 5648 16437 5657
rect 16395 5608 16396 5648
rect 16436 5608 16437 5648
rect 16395 5599 16437 5608
rect 16396 5514 16436 5599
rect 15244 4003 15284 4012
rect 17644 3641 17684 7960
rect 18808 7580 19176 7589
rect 18848 7540 18890 7580
rect 18930 7540 18972 7580
rect 19012 7540 19054 7580
rect 19094 7540 19136 7580
rect 18808 7531 19176 7540
rect 17931 7160 17973 7169
rect 17931 7120 17932 7160
rect 17972 7120 17973 7160
rect 17931 7111 17973 7120
rect 19372 7160 19412 7169
rect 17932 6320 17972 7111
rect 17932 6271 17972 6280
rect 18700 6404 18740 6413
rect 17643 3632 17685 3641
rect 17643 3592 17644 3632
rect 17684 3592 17685 3632
rect 17643 3583 17685 3592
rect 16395 3548 16437 3557
rect 16395 3508 16396 3548
rect 16436 3508 16437 3548
rect 16395 3499 16437 3508
rect 14188 3415 14228 3424
rect 16396 3464 16436 3499
rect 11596 1364 11636 2248
rect 11596 1315 11636 1324
rect 12364 3380 12404 3415
rect 16396 3413 16436 3424
rect 9100 1280 9140 1289
rect 1228 1112 1268 1121
rect 1228 533 1268 1072
rect 9100 1037 9140 1240
rect 12364 1112 12404 3340
rect 14859 3296 14901 3305
rect 14859 3256 14860 3296
rect 14900 3256 14901 3296
rect 14859 3247 14901 3256
rect 14475 2120 14517 2129
rect 14475 2080 14476 2120
rect 14516 2080 14517 2120
rect 14475 2071 14517 2080
rect 12364 1063 12404 1072
rect 14380 1952 14420 1961
rect 9099 1028 9141 1037
rect 9099 988 9100 1028
rect 9140 988 9141 1028
rect 9099 979 9141 988
rect 14380 953 14420 1912
rect 14476 1448 14516 2071
rect 14476 1399 14516 1408
rect 14860 1280 14900 3247
rect 15436 2876 15476 2885
rect 15148 2372 15188 2381
rect 15340 2372 15380 2381
rect 15188 2332 15340 2372
rect 15148 2323 15188 2332
rect 15340 2323 15380 2332
rect 15436 2204 15476 2836
rect 15436 2155 15476 2164
rect 16108 2624 16148 2633
rect 15627 1868 15669 1877
rect 15627 1828 15628 1868
rect 15668 1828 15669 1868
rect 15627 1819 15669 1828
rect 14860 1231 14900 1240
rect 6988 944 7028 953
rect 4928 776 5296 785
rect 4968 736 5010 776
rect 5050 736 5092 776
rect 5132 736 5174 776
rect 5214 736 5256 776
rect 4928 727 5296 736
rect 6988 617 7028 904
rect 14379 944 14421 953
rect 14379 904 14380 944
rect 14420 904 14421 944
rect 14379 895 14421 904
rect 15628 944 15668 1819
rect 16108 1205 16148 2584
rect 16107 1196 16149 1205
rect 16107 1156 16108 1196
rect 16148 1156 16149 1196
rect 16107 1147 16149 1156
rect 16108 1062 16148 1147
rect 17355 1112 17397 1121
rect 17355 1072 17356 1112
rect 17396 1072 17397 1112
rect 17355 1063 17397 1072
rect 17356 978 17396 1063
rect 15628 895 15668 904
rect 17644 776 17684 3583
rect 18124 2792 18164 2801
rect 18124 2549 18164 2752
rect 18123 2540 18165 2549
rect 18123 2500 18124 2540
rect 18164 2500 18165 2540
rect 18123 2491 18165 2500
rect 18028 1784 18068 1795
rect 18028 1709 18068 1744
rect 18027 1700 18069 1709
rect 18027 1660 18028 1700
rect 18068 1660 18069 1700
rect 18027 1651 18069 1660
rect 18028 1364 18068 1651
rect 18028 1315 18068 1324
rect 18700 1364 18740 6364
rect 18808 6068 19176 6077
rect 18848 6028 18890 6068
rect 18930 6028 18972 6068
rect 19012 6028 19054 6068
rect 19094 6028 19136 6068
rect 18808 6019 19176 6028
rect 19372 5732 19412 7120
rect 20048 6824 20416 6833
rect 20088 6784 20130 6824
rect 20170 6784 20212 6824
rect 20252 6784 20294 6824
rect 20334 6784 20376 6824
rect 20048 6775 20416 6784
rect 19851 6572 19893 6581
rect 19851 6532 19852 6572
rect 19892 6532 19893 6572
rect 19851 6523 19893 6532
rect 19852 6438 19892 6523
rect 19372 5683 19412 5692
rect 21388 6068 21428 6077
rect 20048 5312 20416 5321
rect 20088 5272 20130 5312
rect 20170 5272 20212 5312
rect 20252 5272 20294 5312
rect 20334 5272 20376 5312
rect 20048 5263 20416 5272
rect 20620 5312 20660 5321
rect 19371 4976 19413 4985
rect 19371 4936 19372 4976
rect 19412 4936 19413 4976
rect 19371 4927 19413 4936
rect 19276 4892 19316 4901
rect 19276 4565 19316 4852
rect 18808 4556 19176 4565
rect 18848 4516 18890 4556
rect 18930 4516 18972 4556
rect 19012 4516 19054 4556
rect 19094 4516 19136 4556
rect 18808 4507 19176 4516
rect 19275 4556 19317 4565
rect 19275 4516 19276 4556
rect 19316 4516 19317 4556
rect 19275 4507 19317 4516
rect 19372 4145 19412 4927
rect 19659 4724 19701 4733
rect 19659 4684 19660 4724
rect 19700 4684 19701 4724
rect 19659 4675 19701 4684
rect 19371 4136 19413 4145
rect 19371 4096 19372 4136
rect 19412 4096 19413 4136
rect 19371 4087 19413 4096
rect 19372 4001 19412 4087
rect 19660 3884 19700 4675
rect 19660 3835 19700 3844
rect 20048 3800 20416 3809
rect 20088 3760 20130 3800
rect 20170 3760 20212 3800
rect 20252 3760 20294 3800
rect 20334 3760 20376 3800
rect 20048 3751 20416 3760
rect 18891 3380 18933 3389
rect 18891 3340 18892 3380
rect 18932 3340 18933 3380
rect 18891 3331 18933 3340
rect 18892 3212 18932 3331
rect 18892 3163 18932 3172
rect 18808 3044 19176 3053
rect 18848 3004 18890 3044
rect 18930 3004 18972 3044
rect 19012 3004 19054 3044
rect 19094 3004 19136 3044
rect 18808 2995 19176 3004
rect 20044 3044 20084 3053
rect 20044 2540 20084 3004
rect 20236 2624 20276 2633
rect 20236 2540 20276 2584
rect 20044 2500 20276 2540
rect 20332 2456 20372 2465
rect 19948 2416 20332 2456
rect 19948 2288 19988 2416
rect 20332 2407 20372 2416
rect 19948 2239 19988 2248
rect 20048 2288 20416 2297
rect 20088 2248 20130 2288
rect 20170 2248 20212 2288
rect 20252 2248 20294 2288
rect 20334 2248 20376 2288
rect 20048 2239 20416 2248
rect 19275 1784 19317 1793
rect 19275 1744 19276 1784
rect 19316 1744 19317 1784
rect 19275 1735 19317 1744
rect 20332 1784 20372 1793
rect 18808 1532 19176 1541
rect 18848 1492 18890 1532
rect 18930 1492 18972 1532
rect 19012 1492 19054 1532
rect 19094 1492 19136 1532
rect 18808 1483 19176 1492
rect 18700 1315 18740 1324
rect 17644 727 17684 736
rect 18892 1028 18932 1037
rect 18892 617 18932 988
rect 6987 608 7029 617
rect 6987 568 6988 608
rect 7028 568 7029 608
rect 6987 559 7029 568
rect 18891 608 18933 617
rect 18891 568 18892 608
rect 18932 568 18933 608
rect 18891 559 18933 568
rect 1227 524 1269 533
rect 1227 484 1228 524
rect 1268 484 1269 524
rect 1227 475 1269 484
rect 19276 104 19316 1735
rect 20235 1700 20277 1709
rect 20332 1700 20372 1744
rect 20235 1660 20236 1700
rect 20276 1660 20372 1700
rect 20235 1651 20277 1660
rect 20620 1364 20660 5272
rect 21004 5228 21044 5237
rect 20811 4556 20853 4565
rect 20811 4516 20812 4556
rect 20852 4516 20853 4556
rect 20811 4507 20853 4516
rect 20620 1315 20660 1324
rect 20812 1700 20852 4507
rect 21004 3464 21044 5188
rect 21388 4565 21428 6028
rect 22060 5732 22100 5741
rect 22060 5573 22100 5692
rect 22059 5564 22101 5573
rect 22059 5524 22060 5564
rect 22100 5524 22101 5564
rect 22059 5515 22101 5524
rect 21483 5060 21525 5069
rect 21483 5020 21484 5060
rect 21524 5020 21525 5060
rect 21483 5011 21525 5020
rect 21387 4556 21429 4565
rect 21387 4516 21388 4556
rect 21428 4516 21429 4556
rect 21387 4507 21429 4516
rect 21004 3415 21044 3424
rect 21196 3800 21236 3809
rect 20716 1280 20756 1289
rect 20524 944 20564 953
rect 20564 904 20660 944
rect 20524 895 20564 904
rect 20048 776 20416 785
rect 20088 736 20130 776
rect 20170 736 20212 776
rect 20252 736 20294 776
rect 20334 736 20376 776
rect 20048 727 20416 736
rect 20620 776 20660 904
rect 20620 727 20660 736
rect 20716 533 20756 1240
rect 20715 524 20757 533
rect 20715 484 20716 524
rect 20756 484 20757 524
rect 20715 475 20757 484
rect 20716 389 20756 475
rect 20812 356 20852 1660
rect 21196 1280 21236 3760
rect 21484 3464 21524 5011
rect 21484 3415 21524 3424
rect 22636 4976 22676 4985
rect 22636 3716 22676 4936
rect 22636 3464 22676 3676
rect 22636 3415 22676 3424
rect 23788 4388 23828 8464
rect 24364 8454 24404 8539
rect 25420 8504 25460 8513
rect 24171 7160 24213 7169
rect 24171 7120 24172 7160
rect 24212 7120 24213 7160
rect 24171 7111 24213 7120
rect 25420 7160 25460 8464
rect 27723 7916 27765 7925
rect 27723 7876 27724 7916
rect 27764 7876 27765 7916
rect 27723 7867 27765 7876
rect 27724 7782 27764 7867
rect 25420 7111 25460 7120
rect 27628 7160 27668 7169
rect 24172 7026 24212 7111
rect 27628 7001 27668 7120
rect 27627 6992 27669 7001
rect 27627 6952 27628 6992
rect 27668 6952 27669 6992
rect 27627 6943 27669 6952
rect 27723 6572 27765 6581
rect 27723 6532 27724 6572
rect 27764 6532 27765 6572
rect 27723 6523 27765 6532
rect 25324 6488 25364 6497
rect 23979 5480 24021 5489
rect 23979 5440 23980 5480
rect 24020 5440 24021 5480
rect 23979 5431 24021 5440
rect 23980 5060 24020 5431
rect 23980 5011 24020 5020
rect 23788 3464 23828 4348
rect 23788 3415 23828 3424
rect 23884 4892 23924 4901
rect 21196 1231 21236 1240
rect 21964 3380 22004 3389
rect 21964 1112 22004 3340
rect 21964 1063 22004 1072
rect 23884 440 23924 4852
rect 24459 3632 24501 3641
rect 24459 3592 24460 3632
rect 24500 3592 24501 3632
rect 24459 3583 24501 3592
rect 24460 3464 24500 3583
rect 23980 2288 24020 2297
rect 23980 1700 24020 2248
rect 23980 1651 24020 1660
rect 24460 1196 24500 3424
rect 25324 1952 25364 6448
rect 27724 6488 27764 6523
rect 27724 6437 27764 6448
rect 26955 5732 26997 5741
rect 26955 5692 26956 5732
rect 26996 5692 26997 5732
rect 26955 5683 26997 5692
rect 26380 4976 26420 4985
rect 26380 4733 26420 4936
rect 26379 4724 26421 4733
rect 26379 4684 26380 4724
rect 26420 4684 26421 4724
rect 26379 4675 26421 4684
rect 26380 4589 26420 4675
rect 25708 4220 25748 4231
rect 25708 4145 25748 4180
rect 25707 4136 25749 4145
rect 25707 4096 25708 4136
rect 25748 4096 25749 4136
rect 25707 4087 25749 4096
rect 25324 1903 25364 1912
rect 26379 1952 26421 1961
rect 26379 1912 26380 1952
rect 26420 1912 26516 1952
rect 26379 1903 26421 1912
rect 26476 1868 26516 1912
rect 26476 1819 26516 1828
rect 26956 1280 26996 5683
rect 27820 5657 27860 8548
rect 30028 8538 30068 8623
rect 28875 7244 28917 7253
rect 28875 7204 28876 7244
rect 28916 7204 28917 7244
rect 28875 7195 28917 7204
rect 28876 7110 28916 7195
rect 30124 5984 30164 5993
rect 27819 5648 27861 5657
rect 27819 5608 27820 5648
rect 27860 5608 27861 5648
rect 27819 5599 27861 5608
rect 30124 5312 30164 5944
rect 30124 5263 30164 5272
rect 30220 4976 30260 4985
rect 27244 4892 27284 4901
rect 27244 3128 27284 4852
rect 27244 3079 27284 3088
rect 30220 3128 30260 4936
rect 30220 2633 30260 3088
rect 28684 2624 28724 2633
rect 28684 2465 28724 2584
rect 30219 2624 30261 2633
rect 30219 2584 30220 2624
rect 30260 2584 30261 2624
rect 30219 2575 30261 2584
rect 30604 2540 30644 2549
rect 28683 2456 28725 2465
rect 28683 2416 28684 2456
rect 28724 2416 28725 2456
rect 28683 2407 28725 2416
rect 29835 2036 29877 2045
rect 29835 1996 29836 2036
rect 29876 1996 29877 2036
rect 29835 1987 29877 1996
rect 29836 1902 29876 1987
rect 30604 1868 30644 2500
rect 30604 1793 30644 1828
rect 30603 1784 30645 1793
rect 30603 1744 30604 1784
rect 30644 1744 30645 1784
rect 30603 1735 30645 1744
rect 26956 1231 26996 1240
rect 24460 1147 24500 1156
rect 29164 1112 29204 1123
rect 29164 1037 29204 1072
rect 29163 1028 29205 1037
rect 29163 988 29164 1028
rect 29204 988 29205 1028
rect 29163 979 29205 988
rect 30796 776 30836 9388
rect 33928 9092 34296 9101
rect 33968 9052 34010 9092
rect 34050 9052 34092 9092
rect 34132 9052 34174 9092
rect 34214 9052 34256 9092
rect 33928 9043 34296 9052
rect 31180 9008 31220 9017
rect 30987 1868 31029 1877
rect 30987 1828 30988 1868
rect 31028 1828 31029 1868
rect 30987 1819 31029 1828
rect 30988 1734 31028 1819
rect 30796 727 30836 736
rect 31180 776 31220 8968
rect 39820 8756 39860 8765
rect 35168 8336 35536 8345
rect 35208 8296 35250 8336
rect 35290 8296 35332 8336
rect 35372 8296 35414 8336
rect 35454 8296 35496 8336
rect 35168 8287 35536 8296
rect 39820 8009 39860 8716
rect 39819 8000 39861 8009
rect 39819 7960 39820 8000
rect 39860 7960 39861 8000
rect 39819 7951 39861 7960
rect 33100 7916 33140 7925
rect 31659 7076 31701 7085
rect 31659 7036 31660 7076
rect 31700 7036 31701 7076
rect 31659 7027 31701 7036
rect 31660 6942 31700 7027
rect 31756 6404 31796 6413
rect 31756 5984 31796 6364
rect 31756 4136 31796 5944
rect 31756 4087 31796 4096
rect 32620 5564 32660 5573
rect 31852 3464 31892 3473
rect 31852 3305 31892 3424
rect 32620 3380 32660 5524
rect 32716 3632 32756 3643
rect 32716 3557 32756 3592
rect 32715 3548 32757 3557
rect 32715 3508 32716 3548
rect 32756 3508 32757 3548
rect 32715 3499 32757 3508
rect 32620 3340 32756 3380
rect 31851 3296 31893 3305
rect 31851 3256 31852 3296
rect 31892 3256 31893 3296
rect 31851 3247 31893 3256
rect 32620 3128 32660 3137
rect 32620 1868 32660 3088
rect 32620 1819 32660 1828
rect 31180 727 31220 736
rect 23884 391 23924 400
rect 20812 307 20852 316
rect 32716 188 32756 3340
rect 33100 692 33140 7876
rect 33928 7580 34296 7589
rect 33968 7540 34010 7580
rect 34050 7540 34092 7580
rect 34132 7540 34174 7580
rect 34214 7540 34256 7580
rect 33928 7531 34296 7540
rect 35168 6824 35536 6833
rect 35208 6784 35250 6824
rect 35290 6784 35332 6824
rect 35372 6784 35414 6824
rect 35454 6784 35496 6824
rect 35168 6775 35536 6784
rect 39628 6320 39668 6329
rect 33928 6068 34296 6077
rect 33968 6028 34010 6068
rect 34050 6028 34092 6068
rect 34132 6028 34174 6068
rect 34214 6028 34256 6068
rect 33928 6019 34296 6028
rect 39628 5741 39668 6280
rect 39627 5732 39669 5741
rect 39627 5692 39628 5732
rect 39668 5692 39669 5732
rect 39627 5683 39669 5692
rect 35168 5312 35536 5321
rect 35208 5272 35250 5312
rect 35290 5272 35332 5312
rect 35372 5272 35414 5312
rect 35454 5272 35496 5312
rect 35168 5263 35536 5272
rect 33928 4556 34296 4565
rect 33968 4516 34010 4556
rect 34050 4516 34092 4556
rect 34132 4516 34174 4556
rect 34214 4516 34256 4556
rect 33928 4507 34296 4516
rect 34827 4136 34869 4145
rect 34827 4096 34828 4136
rect 34868 4096 34869 4136
rect 34827 4087 34869 4096
rect 37323 4136 37365 4145
rect 37323 4096 37324 4136
rect 37364 4096 37365 4136
rect 37323 4087 37365 4096
rect 34828 4002 34868 4087
rect 35168 3800 35536 3809
rect 35208 3760 35250 3800
rect 35290 3760 35332 3800
rect 35372 3760 35414 3800
rect 35454 3760 35496 3800
rect 35168 3751 35536 3760
rect 34443 3464 34485 3473
rect 34443 3424 34444 3464
rect 34484 3424 34485 3464
rect 34443 3415 34485 3424
rect 34444 3330 34484 3415
rect 37324 3128 37364 4087
rect 39532 3548 39572 3557
rect 38092 3464 38132 3473
rect 38092 3296 38132 3424
rect 39532 3389 39572 3508
rect 39531 3380 39573 3389
rect 39531 3340 39532 3380
rect 39572 3340 39573 3380
rect 39531 3331 39573 3340
rect 38092 3247 38132 3256
rect 37324 3079 37364 3088
rect 33928 3044 34296 3053
rect 33968 3004 34010 3044
rect 34050 3004 34092 3044
rect 34132 3004 34174 3044
rect 34214 3004 34256 3044
rect 33928 2995 34296 3004
rect 35168 2288 35536 2297
rect 35208 2248 35250 2288
rect 35290 2248 35332 2288
rect 35372 2248 35414 2288
rect 35454 2248 35496 2288
rect 35168 2239 35536 2248
rect 33963 2120 34005 2129
rect 33963 2080 33964 2120
rect 34004 2080 34005 2120
rect 33963 2071 34005 2080
rect 33964 1868 34004 2071
rect 33964 1819 34004 1828
rect 33928 1532 34296 1541
rect 33968 1492 34010 1532
rect 34050 1492 34092 1532
rect 34132 1492 34174 1532
rect 34214 1492 34256 1532
rect 33928 1483 34296 1492
rect 40300 1196 40340 1205
rect 34636 1112 34676 1121
rect 34636 953 34676 1072
rect 40203 1112 40245 1121
rect 40300 1112 40340 1156
rect 41259 1196 41301 1205
rect 41259 1156 41260 1196
rect 41300 1156 41301 1196
rect 41259 1147 41301 1156
rect 40203 1072 40204 1112
rect 40244 1072 40340 1112
rect 40203 1063 40245 1072
rect 41260 1062 41300 1147
rect 34635 944 34677 953
rect 34635 904 34636 944
rect 34676 904 34677 944
rect 34635 895 34677 904
rect 35168 776 35536 785
rect 35208 736 35250 776
rect 35290 736 35332 776
rect 35372 736 35414 776
rect 35454 736 35496 776
rect 35168 727 35536 736
rect 33100 643 33140 652
rect 32716 139 32756 148
rect 19276 55 19316 64
<< via4 >>
rect 4928 9808 4968 9848
rect 5010 9808 5050 9848
rect 5092 9808 5132 9848
rect 5174 9808 5214 9848
rect 5256 9808 5296 9848
rect 20048 9808 20088 9848
rect 20130 9808 20170 9848
rect 20212 9808 20252 9848
rect 20294 9808 20334 9848
rect 20376 9808 20416 9848
rect 35168 9808 35208 9848
rect 35250 9808 35290 9848
rect 35332 9808 35372 9848
rect 35414 9808 35454 9848
rect 35496 9808 35536 9848
rect 3688 9052 3728 9092
rect 3770 9052 3810 9092
rect 3852 9052 3892 9092
rect 3934 9052 3974 9092
rect 4016 9052 4056 9092
rect 1228 8632 1268 8672
rect 268 8548 308 8588
rect 3688 7540 3728 7580
rect 3770 7540 3810 7580
rect 3852 7540 3892 7580
rect 3934 7540 3974 7580
rect 4016 7540 4056 7580
rect 1708 6448 1748 6488
rect 3688 6028 3728 6068
rect 3770 6028 3810 6068
rect 3852 6028 3892 6068
rect 3934 6028 3974 6068
rect 4016 6028 4056 6068
rect 1612 4936 1652 4976
rect 1228 4348 1268 4388
rect 1612 3424 1652 3464
rect 3724 5020 3764 5060
rect 3688 4516 3728 4556
rect 3770 4516 3810 4556
rect 3852 4516 3892 4556
rect 3934 4516 3974 4556
rect 4016 4516 4056 4556
rect 3688 3004 3728 3044
rect 3770 3004 3810 3044
rect 3852 3004 3892 3044
rect 3934 3004 3974 3044
rect 4016 3004 4056 3044
rect 4780 8632 4820 8672
rect 6412 8548 6452 8588
rect 4928 8296 4968 8336
rect 5010 8296 5050 8336
rect 5092 8296 5132 8336
rect 5174 8296 5214 8336
rect 5256 8296 5296 8336
rect 4928 6784 4968 6824
rect 5010 6784 5050 6824
rect 5092 6784 5132 6824
rect 5174 6784 5214 6824
rect 5256 6784 5296 6824
rect 4928 5272 4968 5312
rect 5010 5272 5050 5312
rect 5092 5272 5132 5312
rect 5174 5272 5214 5312
rect 5256 5272 5296 5312
rect 9100 7960 9140 8000
rect 12460 8716 12500 8756
rect 18808 9052 18848 9092
rect 18890 9052 18930 9092
rect 18972 9052 19012 9092
rect 19054 9052 19094 9092
rect 19136 9052 19176 9092
rect 22348 8716 22388 8756
rect 15244 8632 15284 8672
rect 13804 7960 13844 8000
rect 10060 7204 10100 7244
rect 8428 5608 8468 5648
rect 8044 5524 8084 5564
rect 4928 3760 4968 3800
rect 5010 3760 5050 3800
rect 5092 3760 5132 3800
rect 5174 3760 5214 3800
rect 5256 3760 5296 3800
rect 5932 2584 5972 2624
rect 14092 7036 14132 7076
rect 11788 5440 11828 5480
rect 10444 3424 10484 3464
rect 4928 2248 4968 2288
rect 5010 2248 5050 2288
rect 5092 2248 5132 2288
rect 5174 2248 5214 2288
rect 5256 2248 5296 2288
rect 7276 1996 7316 2036
rect 9580 1996 9620 2036
rect 3688 1492 3728 1532
rect 3770 1492 3810 1532
rect 3852 1492 3892 1532
rect 3934 1492 3974 1532
rect 4016 1492 4056 1532
rect 12076 4096 12116 4136
rect 14764 6448 14804 6488
rect 14188 4348 14228 4388
rect 14092 4096 14132 4136
rect 12364 3424 12404 3464
rect 15916 8548 15956 8588
rect 30028 8632 30068 8672
rect 24364 8548 24404 8588
rect 20048 8296 20088 8336
rect 20130 8296 20170 8336
rect 20212 8296 20252 8336
rect 20294 8296 20334 8336
rect 20376 8296 20416 8336
rect 16396 6952 16436 6992
rect 16396 5608 16436 5648
rect 18808 7540 18848 7580
rect 18890 7540 18930 7580
rect 18972 7540 19012 7580
rect 19054 7540 19094 7580
rect 19136 7540 19176 7580
rect 17932 7120 17972 7160
rect 17644 3592 17684 3632
rect 16396 3508 16436 3548
rect 14860 3256 14900 3296
rect 14476 2080 14516 2120
rect 9100 988 9140 1028
rect 15628 1828 15668 1868
rect 4928 736 4968 776
rect 5010 736 5050 776
rect 5092 736 5132 776
rect 5174 736 5214 776
rect 5256 736 5296 776
rect 14380 904 14420 944
rect 16108 1156 16148 1196
rect 17356 1072 17396 1112
rect 18124 2500 18164 2540
rect 18028 1660 18068 1700
rect 18808 6028 18848 6068
rect 18890 6028 18930 6068
rect 18972 6028 19012 6068
rect 19054 6028 19094 6068
rect 19136 6028 19176 6068
rect 20048 6784 20088 6824
rect 20130 6784 20170 6824
rect 20212 6784 20252 6824
rect 20294 6784 20334 6824
rect 20376 6784 20416 6824
rect 19852 6532 19892 6572
rect 20048 5272 20088 5312
rect 20130 5272 20170 5312
rect 20212 5272 20252 5312
rect 20294 5272 20334 5312
rect 20376 5272 20416 5312
rect 19372 4936 19412 4976
rect 18808 4516 18848 4556
rect 18890 4516 18930 4556
rect 18972 4516 19012 4556
rect 19054 4516 19094 4556
rect 19136 4516 19176 4556
rect 19276 4516 19316 4556
rect 19660 4684 19700 4724
rect 19372 4096 19412 4136
rect 20048 3760 20088 3800
rect 20130 3760 20170 3800
rect 20212 3760 20252 3800
rect 20294 3760 20334 3800
rect 20376 3760 20416 3800
rect 18892 3340 18932 3380
rect 18808 3004 18848 3044
rect 18890 3004 18930 3044
rect 18972 3004 19012 3044
rect 19054 3004 19094 3044
rect 19136 3004 19176 3044
rect 20048 2248 20088 2288
rect 20130 2248 20170 2288
rect 20212 2248 20252 2288
rect 20294 2248 20334 2288
rect 20376 2248 20416 2288
rect 19276 1744 19316 1784
rect 18808 1492 18848 1532
rect 18890 1492 18930 1532
rect 18972 1492 19012 1532
rect 19054 1492 19094 1532
rect 19136 1492 19176 1532
rect 6988 568 7028 608
rect 18892 568 18932 608
rect 1228 484 1268 524
rect 20236 1660 20276 1700
rect 20812 4516 20852 4556
rect 22060 5524 22100 5564
rect 21484 5020 21524 5060
rect 21388 4516 21428 4556
rect 20048 736 20088 776
rect 20130 736 20170 776
rect 20212 736 20252 776
rect 20294 736 20334 776
rect 20376 736 20416 776
rect 20716 484 20756 524
rect 24172 7120 24212 7160
rect 27724 7876 27764 7916
rect 27628 6952 27668 6992
rect 27724 6532 27764 6572
rect 23980 5440 24020 5480
rect 24460 3592 24500 3632
rect 26956 5692 26996 5732
rect 26380 4684 26420 4724
rect 25708 4096 25748 4136
rect 26380 1912 26420 1952
rect 28876 7204 28916 7244
rect 27820 5608 27860 5648
rect 30220 2584 30260 2624
rect 28684 2416 28724 2456
rect 29836 1996 29876 2036
rect 30604 1744 30644 1784
rect 29164 988 29204 1028
rect 33928 9052 33968 9092
rect 34010 9052 34050 9092
rect 34092 9052 34132 9092
rect 34174 9052 34214 9092
rect 34256 9052 34296 9092
rect 30988 1828 31028 1868
rect 35168 8296 35208 8336
rect 35250 8296 35290 8336
rect 35332 8296 35372 8336
rect 35414 8296 35454 8336
rect 35496 8296 35536 8336
rect 39820 7960 39860 8000
rect 31660 7036 31700 7076
rect 32716 3508 32756 3548
rect 31852 3256 31892 3296
rect 33928 7540 33968 7580
rect 34010 7540 34050 7580
rect 34092 7540 34132 7580
rect 34174 7540 34214 7580
rect 34256 7540 34296 7580
rect 35168 6784 35208 6824
rect 35250 6784 35290 6824
rect 35332 6784 35372 6824
rect 35414 6784 35454 6824
rect 35496 6784 35536 6824
rect 33928 6028 33968 6068
rect 34010 6028 34050 6068
rect 34092 6028 34132 6068
rect 34174 6028 34214 6068
rect 34256 6028 34296 6068
rect 39628 5692 39668 5732
rect 35168 5272 35208 5312
rect 35250 5272 35290 5312
rect 35332 5272 35372 5312
rect 35414 5272 35454 5312
rect 35496 5272 35536 5312
rect 33928 4516 33968 4556
rect 34010 4516 34050 4556
rect 34092 4516 34132 4556
rect 34174 4516 34214 4556
rect 34256 4516 34296 4556
rect 34828 4096 34868 4136
rect 37324 4096 37364 4136
rect 35168 3760 35208 3800
rect 35250 3760 35290 3800
rect 35332 3760 35372 3800
rect 35414 3760 35454 3800
rect 35496 3760 35536 3800
rect 34444 3424 34484 3464
rect 39532 3340 39572 3380
rect 33928 3004 33968 3044
rect 34010 3004 34050 3044
rect 34092 3004 34132 3044
rect 34174 3004 34214 3044
rect 34256 3004 34296 3044
rect 35168 2248 35208 2288
rect 35250 2248 35290 2288
rect 35332 2248 35372 2288
rect 35414 2248 35454 2288
rect 35496 2248 35536 2288
rect 33964 2080 34004 2120
rect 33928 1492 33968 1532
rect 34010 1492 34050 1532
rect 34092 1492 34132 1532
rect 34174 1492 34214 1532
rect 34256 1492 34296 1532
rect 41260 1156 41300 1196
rect 40204 1072 40244 1112
rect 34636 904 34676 944
rect 35168 736 35208 776
rect 35250 736 35290 776
rect 35332 736 35372 776
rect 35414 736 35454 776
rect 35496 736 35536 776
<< metal5 >>
rect 4919 9871 5305 9890
rect 4919 9848 4985 9871
rect 5071 9848 5153 9871
rect 5239 9848 5305 9871
rect 4919 9808 4928 9848
rect 4968 9808 4985 9848
rect 5071 9808 5092 9848
rect 5132 9808 5153 9848
rect 5239 9808 5256 9848
rect 5296 9808 5305 9848
rect 4919 9785 4985 9808
rect 5071 9785 5153 9808
rect 5239 9785 5305 9808
rect 4919 9766 5305 9785
rect 20039 9871 20425 9890
rect 20039 9848 20105 9871
rect 20191 9848 20273 9871
rect 20359 9848 20425 9871
rect 20039 9808 20048 9848
rect 20088 9808 20105 9848
rect 20191 9808 20212 9848
rect 20252 9808 20273 9848
rect 20359 9808 20376 9848
rect 20416 9808 20425 9848
rect 20039 9785 20105 9808
rect 20191 9785 20273 9808
rect 20359 9785 20425 9808
rect 20039 9766 20425 9785
rect 35159 9871 35545 9890
rect 35159 9848 35225 9871
rect 35311 9848 35393 9871
rect 35479 9848 35545 9871
rect 35159 9808 35168 9848
rect 35208 9808 35225 9848
rect 35311 9808 35332 9848
rect 35372 9808 35393 9848
rect 35479 9808 35496 9848
rect 35536 9808 35545 9848
rect 35159 9785 35225 9808
rect 35311 9785 35393 9808
rect 35479 9785 35545 9808
rect 35159 9766 35545 9785
rect 3679 9115 4065 9134
rect 3679 9092 3745 9115
rect 3831 9092 3913 9115
rect 3999 9092 4065 9115
rect 3679 9052 3688 9092
rect 3728 9052 3745 9092
rect 3831 9052 3852 9092
rect 3892 9052 3913 9092
rect 3999 9052 4016 9092
rect 4056 9052 4065 9092
rect 3679 9029 3745 9052
rect 3831 9029 3913 9052
rect 3999 9029 4065 9052
rect 3679 9010 4065 9029
rect 18799 9115 19185 9134
rect 18799 9092 18865 9115
rect 18951 9092 19033 9115
rect 19119 9092 19185 9115
rect 18799 9052 18808 9092
rect 18848 9052 18865 9092
rect 18951 9052 18972 9092
rect 19012 9052 19033 9092
rect 19119 9052 19136 9092
rect 19176 9052 19185 9092
rect 18799 9029 18865 9052
rect 18951 9029 19033 9052
rect 19119 9029 19185 9052
rect 18799 9010 19185 9029
rect 33919 9115 34305 9134
rect 33919 9092 33985 9115
rect 34071 9092 34153 9115
rect 34239 9092 34305 9115
rect 33919 9052 33928 9092
rect 33968 9052 33985 9092
rect 34071 9052 34092 9092
rect 34132 9052 34153 9092
rect 34239 9052 34256 9092
rect 34296 9052 34305 9092
rect 33919 9029 33985 9052
rect 34071 9029 34153 9052
rect 34239 9029 34305 9052
rect 33919 9010 34305 9029
rect 12451 8716 12460 8756
rect 12500 8716 22348 8756
rect 22388 8716 22397 8756
rect 1219 8632 1228 8672
rect 1268 8632 4780 8672
rect 4820 8632 4829 8672
rect 15235 8632 15244 8672
rect 15284 8632 30028 8672
rect 30068 8632 30077 8672
rect 259 8548 268 8588
rect 308 8548 6412 8588
rect 6452 8548 6461 8588
rect 15907 8548 15916 8588
rect 15956 8548 24364 8588
rect 24404 8548 24413 8588
rect 4919 8359 5305 8378
rect 4919 8336 4985 8359
rect 5071 8336 5153 8359
rect 5239 8336 5305 8359
rect 4919 8296 4928 8336
rect 4968 8296 4985 8336
rect 5071 8296 5092 8336
rect 5132 8296 5153 8336
rect 5239 8296 5256 8336
rect 5296 8296 5305 8336
rect 4919 8273 4985 8296
rect 5071 8273 5153 8296
rect 5239 8273 5305 8296
rect 4919 8254 5305 8273
rect 20039 8359 20425 8378
rect 20039 8336 20105 8359
rect 20191 8336 20273 8359
rect 20359 8336 20425 8359
rect 20039 8296 20048 8336
rect 20088 8296 20105 8336
rect 20191 8296 20212 8336
rect 20252 8296 20273 8336
rect 20359 8296 20376 8336
rect 20416 8296 20425 8336
rect 20039 8273 20105 8296
rect 20191 8273 20273 8296
rect 20359 8273 20425 8296
rect 20039 8254 20425 8273
rect 35159 8359 35545 8378
rect 35159 8336 35225 8359
rect 35311 8336 35393 8359
rect 35479 8336 35545 8359
rect 35159 8296 35168 8336
rect 35208 8296 35225 8336
rect 35311 8296 35332 8336
rect 35372 8296 35393 8336
rect 35479 8296 35496 8336
rect 35536 8296 35545 8336
rect 35159 8273 35225 8296
rect 35311 8273 35393 8296
rect 35479 8273 35545 8296
rect 35159 8254 35545 8273
rect 9091 7960 9100 8000
rect 9140 7960 11360 8000
rect 13795 7960 13804 8000
rect 13844 7960 39820 8000
rect 39860 7960 39869 8000
rect 11320 7916 11360 7960
rect 11320 7876 27724 7916
rect 27764 7876 27773 7916
rect 3679 7603 4065 7622
rect 3679 7580 3745 7603
rect 3831 7580 3913 7603
rect 3999 7580 4065 7603
rect 3679 7540 3688 7580
rect 3728 7540 3745 7580
rect 3831 7540 3852 7580
rect 3892 7540 3913 7580
rect 3999 7540 4016 7580
rect 4056 7540 4065 7580
rect 3679 7517 3745 7540
rect 3831 7517 3913 7540
rect 3999 7517 4065 7540
rect 3679 7498 4065 7517
rect 18799 7603 19185 7622
rect 18799 7580 18865 7603
rect 18951 7580 19033 7603
rect 19119 7580 19185 7603
rect 18799 7540 18808 7580
rect 18848 7540 18865 7580
rect 18951 7540 18972 7580
rect 19012 7540 19033 7580
rect 19119 7540 19136 7580
rect 19176 7540 19185 7580
rect 18799 7517 18865 7540
rect 18951 7517 19033 7540
rect 19119 7517 19185 7540
rect 18799 7498 19185 7517
rect 33919 7603 34305 7622
rect 33919 7580 33985 7603
rect 34071 7580 34153 7603
rect 34239 7580 34305 7603
rect 33919 7540 33928 7580
rect 33968 7540 33985 7580
rect 34071 7540 34092 7580
rect 34132 7540 34153 7580
rect 34239 7540 34256 7580
rect 34296 7540 34305 7580
rect 33919 7517 33985 7540
rect 34071 7517 34153 7540
rect 34239 7517 34305 7540
rect 33919 7498 34305 7517
rect 10051 7204 10060 7244
rect 10100 7204 28876 7244
rect 28916 7204 28925 7244
rect 17923 7120 17932 7160
rect 17972 7120 24172 7160
rect 24212 7120 24221 7160
rect 14083 7036 14092 7076
rect 14132 7036 31660 7076
rect 31700 7036 31709 7076
rect 16387 6952 16396 6992
rect 16436 6952 27628 6992
rect 27668 6952 27677 6992
rect 4919 6847 5305 6866
rect 4919 6824 4985 6847
rect 5071 6824 5153 6847
rect 5239 6824 5305 6847
rect 4919 6784 4928 6824
rect 4968 6784 4985 6824
rect 5071 6784 5092 6824
rect 5132 6784 5153 6824
rect 5239 6784 5256 6824
rect 5296 6784 5305 6824
rect 4919 6761 4985 6784
rect 5071 6761 5153 6784
rect 5239 6761 5305 6784
rect 4919 6742 5305 6761
rect 20039 6847 20425 6866
rect 20039 6824 20105 6847
rect 20191 6824 20273 6847
rect 20359 6824 20425 6847
rect 20039 6784 20048 6824
rect 20088 6784 20105 6824
rect 20191 6784 20212 6824
rect 20252 6784 20273 6824
rect 20359 6784 20376 6824
rect 20416 6784 20425 6824
rect 20039 6761 20105 6784
rect 20191 6761 20273 6784
rect 20359 6761 20425 6784
rect 20039 6742 20425 6761
rect 35159 6847 35545 6866
rect 35159 6824 35225 6847
rect 35311 6824 35393 6847
rect 35479 6824 35545 6847
rect 35159 6784 35168 6824
rect 35208 6784 35225 6824
rect 35311 6784 35332 6824
rect 35372 6784 35393 6824
rect 35479 6784 35496 6824
rect 35536 6784 35545 6824
rect 35159 6761 35225 6784
rect 35311 6761 35393 6784
rect 35479 6761 35545 6784
rect 35159 6742 35545 6761
rect 19843 6532 19852 6572
rect 19892 6532 27724 6572
rect 27764 6532 27773 6572
rect 1699 6448 1708 6488
rect 1748 6448 14764 6488
rect 14804 6448 14813 6488
rect 3679 6091 4065 6110
rect 3679 6068 3745 6091
rect 3831 6068 3913 6091
rect 3999 6068 4065 6091
rect 3679 6028 3688 6068
rect 3728 6028 3745 6068
rect 3831 6028 3852 6068
rect 3892 6028 3913 6068
rect 3999 6028 4016 6068
rect 4056 6028 4065 6068
rect 3679 6005 3745 6028
rect 3831 6005 3913 6028
rect 3999 6005 4065 6028
rect 3679 5986 4065 6005
rect 18799 6091 19185 6110
rect 18799 6068 18865 6091
rect 18951 6068 19033 6091
rect 19119 6068 19185 6091
rect 18799 6028 18808 6068
rect 18848 6028 18865 6068
rect 18951 6028 18972 6068
rect 19012 6028 19033 6068
rect 19119 6028 19136 6068
rect 19176 6028 19185 6068
rect 18799 6005 18865 6028
rect 18951 6005 19033 6028
rect 19119 6005 19185 6028
rect 18799 5986 19185 6005
rect 33919 6091 34305 6110
rect 33919 6068 33985 6091
rect 34071 6068 34153 6091
rect 34239 6068 34305 6091
rect 33919 6028 33928 6068
rect 33968 6028 33985 6068
rect 34071 6028 34092 6068
rect 34132 6028 34153 6068
rect 34239 6028 34256 6068
rect 34296 6028 34305 6068
rect 33919 6005 33985 6028
rect 34071 6005 34153 6028
rect 34239 6005 34305 6028
rect 33919 5986 34305 6005
rect 26947 5692 26956 5732
rect 26996 5692 39628 5732
rect 39668 5692 39677 5732
rect 8419 5608 8428 5648
rect 8468 5608 16396 5648
rect 16436 5608 27820 5648
rect 27860 5608 27869 5648
rect 8035 5524 8044 5564
rect 8084 5524 22060 5564
rect 22100 5524 22109 5564
rect 11779 5440 11788 5480
rect 11828 5440 23980 5480
rect 24020 5440 24029 5480
rect 4919 5335 5305 5354
rect 4919 5312 4985 5335
rect 5071 5312 5153 5335
rect 5239 5312 5305 5335
rect 4919 5272 4928 5312
rect 4968 5272 4985 5312
rect 5071 5272 5092 5312
rect 5132 5272 5153 5312
rect 5239 5272 5256 5312
rect 5296 5272 5305 5312
rect 4919 5249 4985 5272
rect 5071 5249 5153 5272
rect 5239 5249 5305 5272
rect 4919 5230 5305 5249
rect 20039 5335 20425 5354
rect 20039 5312 20105 5335
rect 20191 5312 20273 5335
rect 20359 5312 20425 5335
rect 20039 5272 20048 5312
rect 20088 5272 20105 5312
rect 20191 5272 20212 5312
rect 20252 5272 20273 5312
rect 20359 5272 20376 5312
rect 20416 5272 20425 5312
rect 20039 5249 20105 5272
rect 20191 5249 20273 5272
rect 20359 5249 20425 5272
rect 20039 5230 20425 5249
rect 35159 5335 35545 5354
rect 35159 5312 35225 5335
rect 35311 5312 35393 5335
rect 35479 5312 35545 5335
rect 35159 5272 35168 5312
rect 35208 5272 35225 5312
rect 35311 5272 35332 5312
rect 35372 5272 35393 5312
rect 35479 5272 35496 5312
rect 35536 5272 35545 5312
rect 35159 5249 35225 5272
rect 35311 5249 35393 5272
rect 35479 5249 35545 5272
rect 35159 5230 35545 5249
rect 3715 5020 3724 5060
rect 3764 5020 21484 5060
rect 21524 5020 21533 5060
rect 1603 4936 1612 4976
rect 1652 4936 19372 4976
rect 19412 4936 19421 4976
rect 19651 4684 19660 4724
rect 19700 4684 26380 4724
rect 26420 4684 26429 4724
rect 3679 4579 4065 4598
rect 3679 4556 3745 4579
rect 3831 4556 3913 4579
rect 3999 4556 4065 4579
rect 3679 4516 3688 4556
rect 3728 4516 3745 4556
rect 3831 4516 3852 4556
rect 3892 4516 3913 4556
rect 3999 4516 4016 4556
rect 4056 4516 4065 4556
rect 3679 4493 3745 4516
rect 3831 4493 3913 4516
rect 3999 4493 4065 4516
rect 3679 4474 4065 4493
rect 18799 4579 19185 4598
rect 18799 4556 18865 4579
rect 18951 4556 19033 4579
rect 19119 4556 19185 4579
rect 33919 4579 34305 4598
rect 33919 4556 33985 4579
rect 34071 4556 34153 4579
rect 34239 4556 34305 4579
rect 18799 4516 18808 4556
rect 18848 4516 18865 4556
rect 18951 4516 18972 4556
rect 19012 4516 19033 4556
rect 19119 4516 19136 4556
rect 19176 4516 19185 4556
rect 19267 4516 19276 4556
rect 19316 4516 20812 4556
rect 20852 4516 21388 4556
rect 21428 4516 21437 4556
rect 33919 4516 33928 4556
rect 33968 4516 33985 4556
rect 34071 4516 34092 4556
rect 34132 4516 34153 4556
rect 34239 4516 34256 4556
rect 34296 4516 34305 4556
rect 18799 4493 18865 4516
rect 18951 4493 19033 4516
rect 19119 4493 19185 4516
rect 18799 4474 19185 4493
rect 33919 4493 33985 4516
rect 34071 4493 34153 4516
rect 34239 4493 34305 4516
rect 33919 4474 34305 4493
rect 1219 4348 1228 4388
rect 1268 4348 14188 4388
rect 14228 4348 14237 4388
rect 12067 4096 12076 4136
rect 12116 4096 14092 4136
rect 14132 4096 14141 4136
rect 19363 4096 19372 4136
rect 19412 4096 25708 4136
rect 25748 4096 25757 4136
rect 34819 4096 34828 4136
rect 34868 4096 37324 4136
rect 37364 4096 37373 4136
rect 4919 3823 5305 3842
rect 4919 3800 4985 3823
rect 5071 3800 5153 3823
rect 5239 3800 5305 3823
rect 4919 3760 4928 3800
rect 4968 3760 4985 3800
rect 5071 3760 5092 3800
rect 5132 3760 5153 3800
rect 5239 3760 5256 3800
rect 5296 3760 5305 3800
rect 4919 3737 4985 3760
rect 5071 3737 5153 3760
rect 5239 3737 5305 3760
rect 4919 3718 5305 3737
rect 20039 3823 20425 3842
rect 20039 3800 20105 3823
rect 20191 3800 20273 3823
rect 20359 3800 20425 3823
rect 20039 3760 20048 3800
rect 20088 3760 20105 3800
rect 20191 3760 20212 3800
rect 20252 3760 20273 3800
rect 20359 3760 20376 3800
rect 20416 3760 20425 3800
rect 20039 3737 20105 3760
rect 20191 3737 20273 3760
rect 20359 3737 20425 3760
rect 20039 3718 20425 3737
rect 35159 3823 35545 3842
rect 35159 3800 35225 3823
rect 35311 3800 35393 3823
rect 35479 3800 35545 3823
rect 35159 3760 35168 3800
rect 35208 3760 35225 3800
rect 35311 3760 35332 3800
rect 35372 3760 35393 3800
rect 35479 3760 35496 3800
rect 35536 3760 35545 3800
rect 35159 3737 35225 3760
rect 35311 3737 35393 3760
rect 35479 3737 35545 3760
rect 35159 3718 35545 3737
rect 17635 3592 17644 3632
rect 17684 3592 24460 3632
rect 24500 3592 24509 3632
rect 16387 3508 16396 3548
rect 16436 3508 32716 3548
rect 32756 3508 32765 3548
rect 1603 3424 1612 3464
rect 1652 3424 10444 3464
rect 10484 3424 10493 3464
rect 12355 3424 12364 3464
rect 12404 3424 34444 3464
rect 34484 3424 34493 3464
rect 18883 3340 18892 3380
rect 18932 3340 39532 3380
rect 39572 3340 39581 3380
rect 14851 3256 14860 3296
rect 14900 3256 31852 3296
rect 31892 3256 31901 3296
rect 3679 3067 4065 3086
rect 3679 3044 3745 3067
rect 3831 3044 3913 3067
rect 3999 3044 4065 3067
rect 3679 3004 3688 3044
rect 3728 3004 3745 3044
rect 3831 3004 3852 3044
rect 3892 3004 3913 3044
rect 3999 3004 4016 3044
rect 4056 3004 4065 3044
rect 3679 2981 3745 3004
rect 3831 2981 3913 3004
rect 3999 2981 4065 3004
rect 3679 2962 4065 2981
rect 18799 3067 19185 3086
rect 18799 3044 18865 3067
rect 18951 3044 19033 3067
rect 19119 3044 19185 3067
rect 18799 3004 18808 3044
rect 18848 3004 18865 3044
rect 18951 3004 18972 3044
rect 19012 3004 19033 3044
rect 19119 3004 19136 3044
rect 19176 3004 19185 3044
rect 18799 2981 18865 3004
rect 18951 2981 19033 3004
rect 19119 2981 19185 3004
rect 18799 2962 19185 2981
rect 33919 3067 34305 3086
rect 33919 3044 33985 3067
rect 34071 3044 34153 3067
rect 34239 3044 34305 3067
rect 33919 3004 33928 3044
rect 33968 3004 33985 3044
rect 34071 3004 34092 3044
rect 34132 3004 34153 3044
rect 34239 3004 34256 3044
rect 34296 3004 34305 3044
rect 33919 2981 33985 3004
rect 34071 2981 34153 3004
rect 34239 2981 34305 3004
rect 33919 2962 34305 2981
rect 5923 2584 5932 2624
rect 5972 2584 30220 2624
rect 30260 2584 30269 2624
rect 18092 2500 18124 2540
rect 18164 2500 18173 2540
rect 18092 2456 18132 2500
rect 18092 2416 28684 2456
rect 28724 2416 28733 2456
rect 4919 2311 5305 2330
rect 4919 2288 4985 2311
rect 5071 2288 5153 2311
rect 5239 2288 5305 2311
rect 4919 2248 4928 2288
rect 4968 2248 4985 2288
rect 5071 2248 5092 2288
rect 5132 2248 5153 2288
rect 5239 2248 5256 2288
rect 5296 2248 5305 2288
rect 4919 2225 4985 2248
rect 5071 2225 5153 2248
rect 5239 2225 5305 2248
rect 4919 2206 5305 2225
rect 20039 2311 20425 2330
rect 20039 2288 20105 2311
rect 20191 2288 20273 2311
rect 20359 2288 20425 2311
rect 20039 2248 20048 2288
rect 20088 2248 20105 2288
rect 20191 2248 20212 2288
rect 20252 2248 20273 2288
rect 20359 2248 20376 2288
rect 20416 2248 20425 2288
rect 20039 2225 20105 2248
rect 20191 2225 20273 2248
rect 20359 2225 20425 2248
rect 20039 2206 20425 2225
rect 35159 2311 35545 2330
rect 35159 2288 35225 2311
rect 35311 2288 35393 2311
rect 35479 2288 35545 2311
rect 35159 2248 35168 2288
rect 35208 2248 35225 2288
rect 35311 2248 35332 2288
rect 35372 2248 35393 2288
rect 35479 2248 35496 2288
rect 35536 2248 35545 2288
rect 35159 2225 35225 2248
rect 35311 2225 35393 2248
rect 35479 2225 35545 2248
rect 35159 2206 35545 2225
rect 14467 2080 14476 2120
rect 14516 2080 33964 2120
rect 34004 2080 34013 2120
rect 7267 1996 7276 2036
rect 7316 1996 9468 2036
rect 9571 1996 9580 2036
rect 9620 1996 29836 2036
rect 29876 1996 29885 2036
rect 9428 1952 9468 1996
rect 9428 1912 26380 1952
rect 26420 1912 26429 1952
rect 15619 1828 15628 1868
rect 15668 1828 30988 1868
rect 31028 1828 31037 1868
rect 19267 1744 19276 1784
rect 19316 1744 30604 1784
rect 30644 1744 30653 1784
rect 18019 1660 18028 1700
rect 18068 1660 20236 1700
rect 20276 1660 20285 1700
rect 3679 1555 4065 1574
rect 3679 1532 3745 1555
rect 3831 1532 3913 1555
rect 3999 1532 4065 1555
rect 3679 1492 3688 1532
rect 3728 1492 3745 1532
rect 3831 1492 3852 1532
rect 3892 1492 3913 1532
rect 3999 1492 4016 1532
rect 4056 1492 4065 1532
rect 3679 1469 3745 1492
rect 3831 1469 3913 1492
rect 3999 1469 4065 1492
rect 3679 1450 4065 1469
rect 18799 1555 19185 1574
rect 18799 1532 18865 1555
rect 18951 1532 19033 1555
rect 19119 1532 19185 1555
rect 18799 1492 18808 1532
rect 18848 1492 18865 1532
rect 18951 1492 18972 1532
rect 19012 1492 19033 1532
rect 19119 1492 19136 1532
rect 19176 1492 19185 1532
rect 18799 1469 18865 1492
rect 18951 1469 19033 1492
rect 19119 1469 19185 1492
rect 18799 1450 19185 1469
rect 33919 1555 34305 1574
rect 33919 1532 33985 1555
rect 34071 1532 34153 1555
rect 34239 1532 34305 1555
rect 33919 1492 33928 1532
rect 33968 1492 33985 1532
rect 34071 1492 34092 1532
rect 34132 1492 34153 1532
rect 34239 1492 34256 1532
rect 34296 1492 34305 1532
rect 33919 1469 33985 1492
rect 34071 1469 34153 1492
rect 34239 1469 34305 1492
rect 33919 1450 34305 1469
rect 16099 1156 16108 1196
rect 16148 1156 41260 1196
rect 41300 1156 41309 1196
rect 17347 1072 17356 1112
rect 17396 1072 40204 1112
rect 40244 1072 40253 1112
rect 9091 988 9100 1028
rect 9140 988 29164 1028
rect 29204 988 29213 1028
rect 14371 904 14380 944
rect 14420 904 34636 944
rect 34676 904 34685 944
rect 4919 799 5305 818
rect 4919 776 4985 799
rect 5071 776 5153 799
rect 5239 776 5305 799
rect 4919 736 4928 776
rect 4968 736 4985 776
rect 5071 736 5092 776
rect 5132 736 5153 776
rect 5239 736 5256 776
rect 5296 736 5305 776
rect 4919 713 4985 736
rect 5071 713 5153 736
rect 5239 713 5305 736
rect 4919 694 5305 713
rect 20039 799 20425 818
rect 20039 776 20105 799
rect 20191 776 20273 799
rect 20359 776 20425 799
rect 20039 736 20048 776
rect 20088 736 20105 776
rect 20191 736 20212 776
rect 20252 736 20273 776
rect 20359 736 20376 776
rect 20416 736 20425 776
rect 20039 713 20105 736
rect 20191 713 20273 736
rect 20359 713 20425 736
rect 20039 694 20425 713
rect 35159 799 35545 818
rect 35159 776 35225 799
rect 35311 776 35393 799
rect 35479 776 35545 799
rect 35159 736 35168 776
rect 35208 736 35225 776
rect 35311 736 35332 776
rect 35372 736 35393 776
rect 35479 736 35496 776
rect 35536 736 35545 776
rect 35159 713 35225 736
rect 35311 713 35393 736
rect 35479 713 35545 736
rect 35159 694 35545 713
rect 6979 568 6988 608
rect 7028 568 18892 608
rect 18932 568 18941 608
rect 1219 484 1228 524
rect 1268 484 20716 524
rect 20756 484 20765 524
<< via5 >>
rect 4985 9848 5071 9871
rect 5153 9848 5239 9871
rect 4985 9808 5010 9848
rect 5010 9808 5050 9848
rect 5050 9808 5071 9848
rect 5153 9808 5174 9848
rect 5174 9808 5214 9848
rect 5214 9808 5239 9848
rect 4985 9785 5071 9808
rect 5153 9785 5239 9808
rect 20105 9848 20191 9871
rect 20273 9848 20359 9871
rect 20105 9808 20130 9848
rect 20130 9808 20170 9848
rect 20170 9808 20191 9848
rect 20273 9808 20294 9848
rect 20294 9808 20334 9848
rect 20334 9808 20359 9848
rect 20105 9785 20191 9808
rect 20273 9785 20359 9808
rect 35225 9848 35311 9871
rect 35393 9848 35479 9871
rect 35225 9808 35250 9848
rect 35250 9808 35290 9848
rect 35290 9808 35311 9848
rect 35393 9808 35414 9848
rect 35414 9808 35454 9848
rect 35454 9808 35479 9848
rect 35225 9785 35311 9808
rect 35393 9785 35479 9808
rect 3745 9092 3831 9115
rect 3913 9092 3999 9115
rect 3745 9052 3770 9092
rect 3770 9052 3810 9092
rect 3810 9052 3831 9092
rect 3913 9052 3934 9092
rect 3934 9052 3974 9092
rect 3974 9052 3999 9092
rect 3745 9029 3831 9052
rect 3913 9029 3999 9052
rect 18865 9092 18951 9115
rect 19033 9092 19119 9115
rect 18865 9052 18890 9092
rect 18890 9052 18930 9092
rect 18930 9052 18951 9092
rect 19033 9052 19054 9092
rect 19054 9052 19094 9092
rect 19094 9052 19119 9092
rect 18865 9029 18951 9052
rect 19033 9029 19119 9052
rect 33985 9092 34071 9115
rect 34153 9092 34239 9115
rect 33985 9052 34010 9092
rect 34010 9052 34050 9092
rect 34050 9052 34071 9092
rect 34153 9052 34174 9092
rect 34174 9052 34214 9092
rect 34214 9052 34239 9092
rect 33985 9029 34071 9052
rect 34153 9029 34239 9052
rect 4985 8336 5071 8359
rect 5153 8336 5239 8359
rect 4985 8296 5010 8336
rect 5010 8296 5050 8336
rect 5050 8296 5071 8336
rect 5153 8296 5174 8336
rect 5174 8296 5214 8336
rect 5214 8296 5239 8336
rect 4985 8273 5071 8296
rect 5153 8273 5239 8296
rect 20105 8336 20191 8359
rect 20273 8336 20359 8359
rect 20105 8296 20130 8336
rect 20130 8296 20170 8336
rect 20170 8296 20191 8336
rect 20273 8296 20294 8336
rect 20294 8296 20334 8336
rect 20334 8296 20359 8336
rect 20105 8273 20191 8296
rect 20273 8273 20359 8296
rect 35225 8336 35311 8359
rect 35393 8336 35479 8359
rect 35225 8296 35250 8336
rect 35250 8296 35290 8336
rect 35290 8296 35311 8336
rect 35393 8296 35414 8336
rect 35414 8296 35454 8336
rect 35454 8296 35479 8336
rect 35225 8273 35311 8296
rect 35393 8273 35479 8296
rect 3745 7580 3831 7603
rect 3913 7580 3999 7603
rect 3745 7540 3770 7580
rect 3770 7540 3810 7580
rect 3810 7540 3831 7580
rect 3913 7540 3934 7580
rect 3934 7540 3974 7580
rect 3974 7540 3999 7580
rect 3745 7517 3831 7540
rect 3913 7517 3999 7540
rect 18865 7580 18951 7603
rect 19033 7580 19119 7603
rect 18865 7540 18890 7580
rect 18890 7540 18930 7580
rect 18930 7540 18951 7580
rect 19033 7540 19054 7580
rect 19054 7540 19094 7580
rect 19094 7540 19119 7580
rect 18865 7517 18951 7540
rect 19033 7517 19119 7540
rect 33985 7580 34071 7603
rect 34153 7580 34239 7603
rect 33985 7540 34010 7580
rect 34010 7540 34050 7580
rect 34050 7540 34071 7580
rect 34153 7540 34174 7580
rect 34174 7540 34214 7580
rect 34214 7540 34239 7580
rect 33985 7517 34071 7540
rect 34153 7517 34239 7540
rect 4985 6824 5071 6847
rect 5153 6824 5239 6847
rect 4985 6784 5010 6824
rect 5010 6784 5050 6824
rect 5050 6784 5071 6824
rect 5153 6784 5174 6824
rect 5174 6784 5214 6824
rect 5214 6784 5239 6824
rect 4985 6761 5071 6784
rect 5153 6761 5239 6784
rect 20105 6824 20191 6847
rect 20273 6824 20359 6847
rect 20105 6784 20130 6824
rect 20130 6784 20170 6824
rect 20170 6784 20191 6824
rect 20273 6784 20294 6824
rect 20294 6784 20334 6824
rect 20334 6784 20359 6824
rect 20105 6761 20191 6784
rect 20273 6761 20359 6784
rect 35225 6824 35311 6847
rect 35393 6824 35479 6847
rect 35225 6784 35250 6824
rect 35250 6784 35290 6824
rect 35290 6784 35311 6824
rect 35393 6784 35414 6824
rect 35414 6784 35454 6824
rect 35454 6784 35479 6824
rect 35225 6761 35311 6784
rect 35393 6761 35479 6784
rect 3745 6068 3831 6091
rect 3913 6068 3999 6091
rect 3745 6028 3770 6068
rect 3770 6028 3810 6068
rect 3810 6028 3831 6068
rect 3913 6028 3934 6068
rect 3934 6028 3974 6068
rect 3974 6028 3999 6068
rect 3745 6005 3831 6028
rect 3913 6005 3999 6028
rect 18865 6068 18951 6091
rect 19033 6068 19119 6091
rect 18865 6028 18890 6068
rect 18890 6028 18930 6068
rect 18930 6028 18951 6068
rect 19033 6028 19054 6068
rect 19054 6028 19094 6068
rect 19094 6028 19119 6068
rect 18865 6005 18951 6028
rect 19033 6005 19119 6028
rect 33985 6068 34071 6091
rect 34153 6068 34239 6091
rect 33985 6028 34010 6068
rect 34010 6028 34050 6068
rect 34050 6028 34071 6068
rect 34153 6028 34174 6068
rect 34174 6028 34214 6068
rect 34214 6028 34239 6068
rect 33985 6005 34071 6028
rect 34153 6005 34239 6028
rect 4985 5312 5071 5335
rect 5153 5312 5239 5335
rect 4985 5272 5010 5312
rect 5010 5272 5050 5312
rect 5050 5272 5071 5312
rect 5153 5272 5174 5312
rect 5174 5272 5214 5312
rect 5214 5272 5239 5312
rect 4985 5249 5071 5272
rect 5153 5249 5239 5272
rect 20105 5312 20191 5335
rect 20273 5312 20359 5335
rect 20105 5272 20130 5312
rect 20130 5272 20170 5312
rect 20170 5272 20191 5312
rect 20273 5272 20294 5312
rect 20294 5272 20334 5312
rect 20334 5272 20359 5312
rect 20105 5249 20191 5272
rect 20273 5249 20359 5272
rect 35225 5312 35311 5335
rect 35393 5312 35479 5335
rect 35225 5272 35250 5312
rect 35250 5272 35290 5312
rect 35290 5272 35311 5312
rect 35393 5272 35414 5312
rect 35414 5272 35454 5312
rect 35454 5272 35479 5312
rect 35225 5249 35311 5272
rect 35393 5249 35479 5272
rect 3745 4556 3831 4579
rect 3913 4556 3999 4579
rect 3745 4516 3770 4556
rect 3770 4516 3810 4556
rect 3810 4516 3831 4556
rect 3913 4516 3934 4556
rect 3934 4516 3974 4556
rect 3974 4516 3999 4556
rect 3745 4493 3831 4516
rect 3913 4493 3999 4516
rect 18865 4556 18951 4579
rect 19033 4556 19119 4579
rect 33985 4556 34071 4579
rect 34153 4556 34239 4579
rect 18865 4516 18890 4556
rect 18890 4516 18930 4556
rect 18930 4516 18951 4556
rect 19033 4516 19054 4556
rect 19054 4516 19094 4556
rect 19094 4516 19119 4556
rect 33985 4516 34010 4556
rect 34010 4516 34050 4556
rect 34050 4516 34071 4556
rect 34153 4516 34174 4556
rect 34174 4516 34214 4556
rect 34214 4516 34239 4556
rect 18865 4493 18951 4516
rect 19033 4493 19119 4516
rect 33985 4493 34071 4516
rect 34153 4493 34239 4516
rect 4985 3800 5071 3823
rect 5153 3800 5239 3823
rect 4985 3760 5010 3800
rect 5010 3760 5050 3800
rect 5050 3760 5071 3800
rect 5153 3760 5174 3800
rect 5174 3760 5214 3800
rect 5214 3760 5239 3800
rect 4985 3737 5071 3760
rect 5153 3737 5239 3760
rect 20105 3800 20191 3823
rect 20273 3800 20359 3823
rect 20105 3760 20130 3800
rect 20130 3760 20170 3800
rect 20170 3760 20191 3800
rect 20273 3760 20294 3800
rect 20294 3760 20334 3800
rect 20334 3760 20359 3800
rect 20105 3737 20191 3760
rect 20273 3737 20359 3760
rect 35225 3800 35311 3823
rect 35393 3800 35479 3823
rect 35225 3760 35250 3800
rect 35250 3760 35290 3800
rect 35290 3760 35311 3800
rect 35393 3760 35414 3800
rect 35414 3760 35454 3800
rect 35454 3760 35479 3800
rect 35225 3737 35311 3760
rect 35393 3737 35479 3760
rect 3745 3044 3831 3067
rect 3913 3044 3999 3067
rect 3745 3004 3770 3044
rect 3770 3004 3810 3044
rect 3810 3004 3831 3044
rect 3913 3004 3934 3044
rect 3934 3004 3974 3044
rect 3974 3004 3999 3044
rect 3745 2981 3831 3004
rect 3913 2981 3999 3004
rect 18865 3044 18951 3067
rect 19033 3044 19119 3067
rect 18865 3004 18890 3044
rect 18890 3004 18930 3044
rect 18930 3004 18951 3044
rect 19033 3004 19054 3044
rect 19054 3004 19094 3044
rect 19094 3004 19119 3044
rect 18865 2981 18951 3004
rect 19033 2981 19119 3004
rect 33985 3044 34071 3067
rect 34153 3044 34239 3067
rect 33985 3004 34010 3044
rect 34010 3004 34050 3044
rect 34050 3004 34071 3044
rect 34153 3004 34174 3044
rect 34174 3004 34214 3044
rect 34214 3004 34239 3044
rect 33985 2981 34071 3004
rect 34153 2981 34239 3004
rect 4985 2288 5071 2311
rect 5153 2288 5239 2311
rect 4985 2248 5010 2288
rect 5010 2248 5050 2288
rect 5050 2248 5071 2288
rect 5153 2248 5174 2288
rect 5174 2248 5214 2288
rect 5214 2248 5239 2288
rect 4985 2225 5071 2248
rect 5153 2225 5239 2248
rect 20105 2288 20191 2311
rect 20273 2288 20359 2311
rect 20105 2248 20130 2288
rect 20130 2248 20170 2288
rect 20170 2248 20191 2288
rect 20273 2248 20294 2288
rect 20294 2248 20334 2288
rect 20334 2248 20359 2288
rect 20105 2225 20191 2248
rect 20273 2225 20359 2248
rect 35225 2288 35311 2311
rect 35393 2288 35479 2311
rect 35225 2248 35250 2288
rect 35250 2248 35290 2288
rect 35290 2248 35311 2288
rect 35393 2248 35414 2288
rect 35414 2248 35454 2288
rect 35454 2248 35479 2288
rect 35225 2225 35311 2248
rect 35393 2225 35479 2248
rect 3745 1532 3831 1555
rect 3913 1532 3999 1555
rect 3745 1492 3770 1532
rect 3770 1492 3810 1532
rect 3810 1492 3831 1532
rect 3913 1492 3934 1532
rect 3934 1492 3974 1532
rect 3974 1492 3999 1532
rect 3745 1469 3831 1492
rect 3913 1469 3999 1492
rect 18865 1532 18951 1555
rect 19033 1532 19119 1555
rect 18865 1492 18890 1532
rect 18890 1492 18930 1532
rect 18930 1492 18951 1532
rect 19033 1492 19054 1532
rect 19054 1492 19094 1532
rect 19094 1492 19119 1532
rect 18865 1469 18951 1492
rect 19033 1469 19119 1492
rect 33985 1532 34071 1555
rect 34153 1532 34239 1555
rect 33985 1492 34010 1532
rect 34010 1492 34050 1532
rect 34050 1492 34071 1532
rect 34153 1492 34174 1532
rect 34174 1492 34214 1532
rect 34214 1492 34239 1532
rect 33985 1469 34071 1492
rect 34153 1469 34239 1492
rect 4985 776 5071 799
rect 5153 776 5239 799
rect 4985 736 5010 776
rect 5010 736 5050 776
rect 5050 736 5071 776
rect 5153 736 5174 776
rect 5174 736 5214 776
rect 5214 736 5239 776
rect 4985 713 5071 736
rect 5153 713 5239 736
rect 20105 776 20191 799
rect 20273 776 20359 799
rect 20105 736 20130 776
rect 20130 736 20170 776
rect 20170 736 20191 776
rect 20273 736 20294 776
rect 20294 736 20334 776
rect 20334 736 20359 776
rect 20105 713 20191 736
rect 20273 713 20359 736
rect 35225 776 35311 799
rect 35393 776 35479 799
rect 35225 736 35250 776
rect 35250 736 35290 776
rect 35290 736 35311 776
rect 35393 736 35414 776
rect 35414 736 35454 776
rect 35454 736 35479 776
rect 35225 713 35311 736
rect 35393 713 35479 736
<< metal6 >>
rect 3652 9115 4092 10752
rect 3652 9029 3745 9115
rect 3831 9029 3913 9115
rect 3999 9029 4092 9115
rect 3652 7603 4092 9029
rect 3652 7517 3745 7603
rect 3831 7517 3913 7603
rect 3999 7517 4092 7603
rect 3652 6091 4092 7517
rect 3652 6005 3745 6091
rect 3831 6005 3913 6091
rect 3999 6005 4092 6091
rect 3652 4579 4092 6005
rect 3652 4493 3745 4579
rect 3831 4493 3913 4579
rect 3999 4493 4092 4579
rect 3652 3067 4092 4493
rect 3652 2981 3745 3067
rect 3831 2981 3913 3067
rect 3999 2981 4092 3067
rect 3652 1555 4092 2981
rect 3652 1469 3745 1555
rect 3831 1469 3913 1555
rect 3999 1469 4092 1555
rect 3652 0 4092 1469
rect 4892 9871 5332 10752
rect 4892 9785 4985 9871
rect 5071 9785 5153 9871
rect 5239 9785 5332 9871
rect 4892 8359 5332 9785
rect 4892 8273 4985 8359
rect 5071 8273 5153 8359
rect 5239 8273 5332 8359
rect 4892 6847 5332 8273
rect 4892 6761 4985 6847
rect 5071 6761 5153 6847
rect 5239 6761 5332 6847
rect 4892 5335 5332 6761
rect 4892 5249 4985 5335
rect 5071 5249 5153 5335
rect 5239 5249 5332 5335
rect 4892 3823 5332 5249
rect 4892 3737 4985 3823
rect 5071 3737 5153 3823
rect 5239 3737 5332 3823
rect 4892 2311 5332 3737
rect 4892 2225 4985 2311
rect 5071 2225 5153 2311
rect 5239 2225 5332 2311
rect 4892 799 5332 2225
rect 4892 713 4985 799
rect 5071 713 5153 799
rect 5239 713 5332 799
rect 4892 0 5332 713
rect 18772 9115 19212 10752
rect 18772 9029 18865 9115
rect 18951 9029 19033 9115
rect 19119 9029 19212 9115
rect 18772 7603 19212 9029
rect 18772 7517 18865 7603
rect 18951 7517 19033 7603
rect 19119 7517 19212 7603
rect 18772 6091 19212 7517
rect 18772 6005 18865 6091
rect 18951 6005 19033 6091
rect 19119 6005 19212 6091
rect 18772 4579 19212 6005
rect 18772 4493 18865 4579
rect 18951 4493 19033 4579
rect 19119 4493 19212 4579
rect 18772 3067 19212 4493
rect 18772 2981 18865 3067
rect 18951 2981 19033 3067
rect 19119 2981 19212 3067
rect 18772 1555 19212 2981
rect 18772 1469 18865 1555
rect 18951 1469 19033 1555
rect 19119 1469 19212 1555
rect 18772 0 19212 1469
rect 20012 9871 20452 10752
rect 20012 9785 20105 9871
rect 20191 9785 20273 9871
rect 20359 9785 20452 9871
rect 20012 8359 20452 9785
rect 20012 8273 20105 8359
rect 20191 8273 20273 8359
rect 20359 8273 20452 8359
rect 20012 6847 20452 8273
rect 20012 6761 20105 6847
rect 20191 6761 20273 6847
rect 20359 6761 20452 6847
rect 20012 5335 20452 6761
rect 20012 5249 20105 5335
rect 20191 5249 20273 5335
rect 20359 5249 20452 5335
rect 20012 3823 20452 5249
rect 20012 3737 20105 3823
rect 20191 3737 20273 3823
rect 20359 3737 20452 3823
rect 20012 2311 20452 3737
rect 20012 2225 20105 2311
rect 20191 2225 20273 2311
rect 20359 2225 20452 2311
rect 20012 799 20452 2225
rect 20012 713 20105 799
rect 20191 713 20273 799
rect 20359 713 20452 799
rect 20012 0 20452 713
rect 33892 9115 34332 10752
rect 33892 9029 33985 9115
rect 34071 9029 34153 9115
rect 34239 9029 34332 9115
rect 33892 7603 34332 9029
rect 33892 7517 33985 7603
rect 34071 7517 34153 7603
rect 34239 7517 34332 7603
rect 33892 6091 34332 7517
rect 33892 6005 33985 6091
rect 34071 6005 34153 6091
rect 34239 6005 34332 6091
rect 33892 4579 34332 6005
rect 33892 4493 33985 4579
rect 34071 4493 34153 4579
rect 34239 4493 34332 4579
rect 33892 3067 34332 4493
rect 33892 2981 33985 3067
rect 34071 2981 34153 3067
rect 34239 2981 34332 3067
rect 33892 1555 34332 2981
rect 33892 1469 33985 1555
rect 34071 1469 34153 1555
rect 34239 1469 34332 1555
rect 33892 0 34332 1469
rect 35132 9871 35572 10752
rect 35132 9785 35225 9871
rect 35311 9785 35393 9871
rect 35479 9785 35572 9871
rect 35132 8359 35572 9785
rect 35132 8273 35225 8359
rect 35311 8273 35393 8359
rect 35479 8273 35572 8359
rect 35132 6847 35572 8273
rect 35132 6761 35225 6847
rect 35311 6761 35393 6847
rect 35479 6761 35572 6847
rect 35132 5335 35572 6761
rect 35132 5249 35225 5335
rect 35311 5249 35393 5335
rect 35479 5249 35572 5335
rect 35132 3823 35572 5249
rect 35132 3737 35225 3823
rect 35311 3737 35393 3823
rect 35479 3737 35572 3823
rect 35132 2311 35572 3737
rect 35132 2225 35225 2311
rect 35311 2225 35393 2311
rect 35479 2225 35572 2311
rect 35132 799 35572 2225
rect 35132 713 35225 799
rect 35311 713 35393 799
rect 35479 713 35572 799
rect 35132 0 35572 713
use sg13g2_mux4_1  _047_
timestamp 1677257233
transform 1 0 23232 0 -1 5292
box -48 -56 2064 834
use sg13g2_mux4_1  _048_
timestamp 1677257233
transform 1 0 27552 0 -1 2268
box -48 -56 2064 834
use sg13g2_mux4_1  _049_
timestamp 1677257233
transform 1 0 20928 0 1 3780
box -48 -56 2064 834
use sg13g2_mux4_1  _050_
timestamp 1677257233
transform 1 0 13824 0 1 3780
box -48 -56 2064 834
use sg13g2_mux4_1  _051_
timestamp 1677257233
transform 1 0 21792 0 1 8316
box -48 -56 2064 834
use sg13g2_mux4_1  _052_
timestamp 1677257233
transform 1 0 28512 0 -1 8316
box -48 -56 2064 834
use sg13g2_mux4_1  _053_
timestamp 1677257233
transform 1 0 21408 0 -1 6804
box -48 -56 2064 834
use sg13g2_mux4_1  _054_
timestamp 1677257233
transform 1 0 10944 0 -1 2268
box -48 -56 2064 834
use sg13g2_mux4_1  _055_
timestamp 1677257233
transform 1 0 20160 0 -1 2268
box -48 -56 2064 834
use sg13g2_mux4_1  _056_
timestamp 1677257233
transform 1 0 17280 0 -1 2268
box -48 -56 2064 834
use sg13g2_mux4_1  _057_
timestamp 1677257233
transform 1 0 16608 0 -1 5292
box -48 -56 2064 834
use sg13g2_mux4_1  _058_
timestamp 1677257233
transform 1 0 13728 0 -1 5292
box -48 -56 2064 834
use sg13g2_mux4_1  _059_
timestamp 1677257233
transform 1 0 17472 0 1 8316
box -48 -56 2064 834
use sg13g2_mux4_1  _060_
timestamp 1677257233
transform 1 0 19104 0 1 6804
box -48 -56 2064 834
use sg13g2_mux4_1  _061_
timestamp 1677257233
transform 1 0 17760 0 -1 6804
box -48 -56 2064 834
use sg13g2_mux4_1  _062_
timestamp 1677257233
transform 1 0 10752 0 1 2268
box -48 -56 2064 834
use sg13g2_mux4_1  _063_
timestamp 1677257233
transform 1 0 18624 0 -1 5292
box -48 -56 2064 834
use sg13g2_mux2_1  _064_
timestamp 1677247768
transform 1 0 30432 0 1 3780
box -48 -56 1008 834
use sg13g2_mux2_1  _065_
timestamp 1677247768
transform 1 0 19488 0 1 2268
box -48 -56 1008 834
use sg13g2_mux2_1  _066_
timestamp 1677247768
transform 1 0 23616 0 1 2268
box -48 -56 1008 834
use sg13g2_mux2_1  _067_
timestamp 1677247768
transform 1 0 8256 0 -1 5292
box -48 -56 1008 834
use sg13g2_nand2b_1  _068_
timestamp 1676567195
transform 1 0 3744 0 -1 9828
box -48 -56 528 834
use sg13g2_o21ai_1  _069_
timestamp 1685175443
transform -1 0 4416 0 1 8316
box -48 -56 538 834
use sg13g2_nand3_1  _070_
timestamp 1683988354
transform 1 0 3456 0 1 8316
box -48 -56 528 834
use sg13g2_o21ai_1  _071_
timestamp 1685175443
transform 1 0 3264 0 -1 9828
box -48 -56 538 834
use sg13g2_nand3b_1  _072_
timestamp 1676573470
transform 1 0 3264 0 -1 8316
box -48 -56 720 834
use sg13g2_o21ai_1  _073_
timestamp 1685175443
transform -1 0 3360 0 1 6804
box -48 -56 538 834
use sg13g2_nand2_1  _074_
timestamp 1676557249
transform 1 0 3360 0 -1 6804
box -48 -56 432 834
use sg13g2_nand4_1  _075_
timestamp 1685201930
transform 1 0 3360 0 1 6804
box -48 -56 624 834
use sg13g2_o21ai_1  _076_
timestamp 1685175443
transform 1 0 4224 0 -1 9828
box -48 -56 538 834
use sg13g2_nand2b_1  _077_
timestamp 1676567195
transform -1 0 8736 0 -1 8316
box -48 -56 528 834
use sg13g2_mux4_1  _078_
timestamp 1677257233
transform 1 0 7104 0 1 6804
box -48 -56 2064 834
use sg13g2_o21ai_1  _079_
timestamp 1685175443
transform -1 0 8256 0 -1 8316
box -48 -56 538 834
use sg13g2_o21ai_1  _080_
timestamp 1685175443
transform -1 0 7104 0 1 6804
box -48 -56 538 834
use sg13g2_nand2b_1  _081_
timestamp 1676567195
transform 1 0 9120 0 1 6804
box -48 -56 528 834
use sg13g2_o21ai_1  _082_
timestamp 1685175443
transform 1 0 9600 0 1 6804
box -48 -56 538 834
use sg13g2_inv_1  _083_
timestamp 1676382929
transform -1 0 4800 0 -1 5292
box -48 -56 336 834
use sg13g2_inv_1  _084_
timestamp 1676382929
transform 1 0 2976 0 -1 8316
box -48 -56 336 834
use sg13g2_mux2_1  _085_
timestamp 1677247768
transform 1 0 3744 0 -1 6804
box -48 -56 1008 834
use sg13g2_or2_1  _086_
timestamp 1684236171
transform 1 0 4224 0 1 6804
box -48 -56 528 834
use sg13g2_a21oi_1  _087_
timestamp 1683973020
transform 1 0 4032 0 1 5292
box -48 -56 528 834
use sg13g2_a221oi_1  _088_
timestamp 1685197497
transform -1 0 5472 0 -1 6804
box -48 -56 816 834
use sg13g2_nand2_1  _089_
timestamp 1676557249
transform 1 0 4992 0 -1 5292
box -48 -56 432 834
use sg13g2_nand2b_1  _090_
timestamp 1676567195
transform 1 0 4704 0 1 6804
box -48 -56 528 834
use sg13g2_a21oi_1  _091_
timestamp 1683973020
transform -1 0 5472 0 1 5292
box -48 -56 528 834
use sg13g2_nor2b_1  _092_
timestamp 1685181386
transform 1 0 4512 0 1 5292
box -54 -56 528 834
use sg13g2_o21ai_1  _093_
timestamp 1685175443
transform 1 0 5472 0 -1 6804
box -48 -56 538 834
use sg13g2_o21ai_1  _094_
timestamp 1685175443
transform 1 0 5952 0 -1 6804
box -48 -56 538 834
use sg13g2_o21ai_1  _095_
timestamp 1685175443
transform 1 0 5184 0 1 6804
box -48 -56 538 834
use sg13g2_mux4_1  _096_
timestamp 1677257233
transform 1 0 5472 0 1 5292
box -48 -56 2064 834
use sg13g2_mux4_1  _097_
timestamp 1677257233
transform 1 0 5376 0 -1 5292
box -48 -56 2064 834
use sg13g2_mux2_1  _098_
timestamp 1677247768
transform -1 0 7392 0 -1 6804
box -48 -56 1008 834
use sg13g2_nand2b_1  _099_
timestamp 1676567195
transform 1 0 6144 0 1 6804
box -48 -56 528 834
use sg13g2_o21ai_1  _100_
timestamp 1685175443
transform 1 0 5664 0 1 6804
box -48 -56 538 834
use sg13g2_mux2_1  _101_
timestamp 1677247768
transform 1 0 3360 0 1 3780
box -48 -56 1008 834
use sg13g2_or2_1  _102_
timestamp 1684236171
transform -1 0 5280 0 1 3780
box -48 -56 528 834
use sg13g2_a21oi_1  _103_
timestamp 1683973020
transform 1 0 4320 0 1 3780
box -48 -56 528 834
use sg13g2_a221oi_1  _104_
timestamp 1685197497
transform 1 0 3552 0 -1 3780
box -48 -56 816 834
use sg13g2_nand2_1  _105_
timestamp 1676557249
transform 1 0 3168 0 -1 3780
box -48 -56 432 834
use sg13g2_nand2b_1  _106_
timestamp 1676567195
transform 1 0 4128 0 1 2268
box -48 -56 528 834
use sg13g2_a21oi_1  _107_
timestamp 1683973020
transform 1 0 4032 0 -1 5292
box -48 -56 528 834
use sg13g2_nor2b_1  _108_
timestamp 1685181386
transform -1 0 5280 0 1 2268
box -54 -56 528 834
use sg13g2_o21ai_1  _109_
timestamp 1685175443
transform -1 0 5376 0 -1 3780
box -48 -56 538 834
use sg13g2_o21ai_1  _110_
timestamp 1685175443
transform -1 0 4896 0 -1 3780
box -48 -56 538 834
use sg13g2_o21ai_1  _111_
timestamp 1685175443
transform -1 0 3648 0 1 2268
box -48 -56 538 834
use sg13g2_mux4_1  _112_
timestamp 1677257233
transform 1 0 5376 0 -1 3780
box -48 -56 2064 834
use sg13g2_mux4_1  _113_
timestamp 1677257233
transform 1 0 5472 0 1 3780
box -48 -56 2064 834
use sg13g2_mux2_1  _114_
timestamp 1677247768
transform -1 0 8352 0 -1 3780
box -48 -56 1008 834
use sg13g2_nand2b_1  _115_
timestamp 1676567195
transform 1 0 3648 0 1 2268
box -48 -56 528 834
use sg13g2_o21ai_1  _116_
timestamp 1685175443
transform -1 0 4032 0 -1 5292
box -48 -56 538 834
use sg13g2_mux4_1  _117_
timestamp 1677257233
transform 1 0 7680 0 -1 2268
box -48 -56 2064 834
use sg13g2_mux4_1  _118_
timestamp 1677257233
transform 1 0 5088 0 1 756
box -48 -56 2064 834
use sg13g2_mux4_1  _119_
timestamp 1677257233
transform 1 0 35136 0 1 5292
box -48 -56 2064 834
use sg13g2_mux4_1  _120_
timestamp 1677257233
transform 1 0 38112 0 -1 5292
box -48 -56 2064 834
use sg13g2_mux4_1  _121_
timestamp 1677257233
transform 1 0 35904 0 1 2268
box -48 -56 2064 834
use sg13g2_mux4_1  _122_
timestamp 1677257233
transform 1 0 31776 0 -1 5292
box -48 -56 2064 834
use sg13g2_mux4_1  _123_
timestamp 1677257233
transform 1 0 38112 0 -1 2268
box -48 -56 2064 834
use sg13g2_mux4_1  _124_
timestamp 1677257233
transform 1 0 35136 0 -1 2268
box -48 -56 2064 834
use sg13g2_mux4_1  _125_
timestamp 1677257233
transform 1 0 5376 0 -1 2268
box -48 -56 2064 834
use sg13g2_mux4_1  _126_
timestamp 1677257233
transform 1 0 9888 0 1 5292
box -48 -56 2064 834
use sg13g2_mux4_1  _127_
timestamp 1677257233
transform 1 0 13632 0 1 6804
box -48 -56 2064 834
use sg13g2_mux4_1  _128_
timestamp 1677257233
transform 1 0 11136 0 1 6804
box -48 -56 2064 834
use sg13g2_mux4_1  _129_
timestamp 1677257233
transform 1 0 34944 0 1 6804
box -48 -56 2064 834
use sg13g2_mux4_1  _130_
timestamp 1677257233
transform 1 0 37824 0 1 6804
box -48 -56 2064 834
use sg13g2_mux4_1  _131_
timestamp 1677257233
transform 1 0 36000 0 -1 3780
box -48 -56 2064 834
use sg13g2_mux4_1  _132_
timestamp 1677257233
transform 1 0 31680 0 1 5292
box -48 -56 2064 834
use sg13g2_mux4_1  _133_
timestamp 1677257233
transform 1 0 31104 0 1 756
box -48 -56 2064 834
use sg13g2_mux4_1  _134_
timestamp 1677257233
transform 1 0 27360 0 1 3780
box -48 -56 2064 834
use sg13g2_mux4_1  _135_
timestamp 1677257233
transform 1 0 30912 0 -1 8316
box -48 -56 2064 834
use sg13g2_mux4_1  _136_
timestamp 1677257233
transform 1 0 24768 0 -1 3780
box -48 -56 2064 834
use sg13g2_mux4_1  _137_
timestamp 1677257233
transform 1 0 31584 0 -1 3780
box -48 -56 2064 834
use sg13g2_mux4_1  _138_
timestamp 1677257233
transform 1 0 27456 0 1 5292
box -48 -56 2064 834
use sg13g2_mux4_1  _139_
timestamp 1677257233
transform 1 0 30336 0 -1 2268
box -48 -56 2064 834
use sg13g2_mux4_1  _140_
timestamp 1677257233
transform 1 0 24576 0 -1 2268
box -48 -56 2064 834
use sg13g2_mux4_1  _141_
timestamp 1677257233
transform 1 0 14976 0 -1 2268
box -48 -56 2064 834
use sg13g2_mux4_1  _142_
timestamp 1677257233
transform 1 0 25248 0 1 8316
box -48 -56 2064 834
use sg13g2_mux4_1  _143_
timestamp 1677257233
transform 1 0 10944 0 -1 3780
box -48 -56 2064 834
use sg13g2_mux4_1  _144_
timestamp 1677257233
transform 1 0 23712 0 1 5292
box -48 -56 2064 834
use sg13g2_mux4_1  _145_
timestamp 1677257233
transform 1 0 16128 0 -1 3780
box -48 -56 2064 834
use sg13g2_mux4_1  _146_
timestamp 1677257233
transform 1 0 25152 0 -1 8316
box -48 -56 2064 834
use sg13g2_mux4_1  _147_
timestamp 1677257233
transform 1 0 13728 0 1 2268
box -48 -56 2064 834
use sg13g2_dlhq_1  _148_
timestamp 1678805552
transform 1 0 7680 0 -1 9828
box -50 -56 1692 834
use sg13g2_dlhq_1  _149_
timestamp 1678805552
transform 1 0 7968 0 1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _150_
timestamp 1678805552
transform 1 0 8832 0 -1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _151_
timestamp 1678805552
transform 1 0 10176 0 -1 9828
box -50 -56 1692 834
use sg13g2_dlhq_1  _152_
timestamp 1678805552
transform 1 0 11808 0 -1 9828
box -50 -56 1692 834
use sg13g2_dlhq_1  _153_
timestamp 1678805552
transform 1 0 12384 0 1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _154_
timestamp 1678805552
transform 1 0 14016 0 1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _155_
timestamp 1678805552
transform 1 0 15168 0 -1 9828
box -50 -56 1692 834
use sg13g2_dlhq_1  _156_
timestamp 1678805552
transform 1 0 7968 0 1 3780
box -50 -56 1692 834
use sg13g2_dlhq_1  _157_
timestamp 1678805552
transform 1 0 22368 0 -1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _158_
timestamp 1678805552
transform 1 0 17856 0 1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _159_
timestamp 1678805552
transform 1 0 28992 0 -1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _160_
timestamp 1678805552
transform 1 0 17280 0 1 3780
box -50 -56 1692 834
use sg13g2_dlhq_1  _161_
timestamp 1678805552
transform 1 0 19200 0 1 3780
box -50 -56 1692 834
use sg13g2_dlhq_1  _162_
timestamp 1678805552
transform 1 0 8640 0 -1 3780
box -50 -56 1692 834
use sg13g2_dlhq_1  _163_
timestamp 1678805552
transform 1 0 10368 0 1 3780
box -50 -56 1692 834
use sg13g2_dlhq_1  _164_
timestamp 1678805552
transform 1 0 16224 0 1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _165_
timestamp 1678805552
transform 1 0 17952 0 1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _166_
timestamp 1678805552
transform 1 0 17760 0 -1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _167_
timestamp 1678805552
transform 1 0 19680 0 -1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _168_
timestamp 1678805552
transform 1 0 15840 0 1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _169_
timestamp 1678805552
transform 1 0 17760 0 -1 9828
box -50 -56 1692 834
use sg13g2_dlhq_1  _170_
timestamp 1678805552
transform 1 0 12192 0 -1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _171_
timestamp 1678805552
transform 1 0 13056 0 1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _172_
timestamp 1678805552
transform 1 0 14688 0 1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _173_
timestamp 1678805552
transform 1 0 16320 0 1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _174_
timestamp 1678805552
transform 1 0 15840 0 1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _175_
timestamp 1678805552
transform 1 0 17280 0 1 756
box -50 -56 1692 834
use sg13g2_dlhq_1  _176_
timestamp 1678805552
transform 1 0 18912 0 1 756
box -50 -56 1692 834
use sg13g2_dlhq_1  _177_
timestamp 1678805552
transform 1 0 20640 0 1 756
box -50 -56 1692 834
use sg13g2_dlhq_1  _178_
timestamp 1678805552
transform 1 0 9024 0 1 756
box -50 -56 1692 834
use sg13g2_dlhq_1  _179_
timestamp 1678805552
transform 1 0 9120 0 1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _180_
timestamp 1678805552
transform 1 0 19776 0 -1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _181_
timestamp 1678805552
transform 1 0 21984 0 1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _182_
timestamp 1678805552
transform 1 0 27648 0 -1 9828
box -50 -56 1692 834
use sg13g2_dlhq_1  _183_
timestamp 1678805552
transform 1 0 28800 0 1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _184_
timestamp 1678805552
transform 1 0 20160 0 1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _185_
timestamp 1678805552
transform 1 0 22368 0 -1 9828
box -50 -56 1692 834
use sg13g2_dlhq_1  _186_
timestamp 1678805552
transform 1 0 12000 0 1 3780
box -50 -56 1692 834
use sg13g2_dlhq_1  _187_
timestamp 1678805552
transform 1 0 14112 0 -1 3780
box -50 -56 1692 834
use sg13g2_dlhq_1  _188_
timestamp 1678805552
transform 1 0 19584 0 -1 3780
box -50 -56 1692 834
use sg13g2_dlhq_1  _189_
timestamp 1678805552
transform 1 0 21312 0 -1 3780
box -50 -56 1692 834
use sg13g2_dlhq_1  _190_
timestamp 1678805552
transform -1 0 28896 0 1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _191_
timestamp 1678805552
transform -1 0 30528 0 1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _192_
timestamp 1678805552
transform 1 0 21600 0 -1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _193_
timestamp 1678805552
transform -1 0 25824 0 1 3780
box -50 -56 1692 834
use sg13g2_dlhq_1  _194_
timestamp 1678805552
transform 1 0 12288 0 1 756
box -50 -56 1692 834
use sg13g2_dlhq_1  _195_
timestamp 1678805552
transform 1 0 13344 0 -1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _196_
timestamp 1678805552
transform -1 0 27840 0 1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _197_
timestamp 1678805552
transform 1 0 24096 0 1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _198_
timestamp 1678805552
transform 1 0 16032 0 -1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _199_
timestamp 1678805552
transform 1 0 14688 0 -1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _200_
timestamp 1678805552
transform 1 0 24288 0 -1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _201_
timestamp 1678805552
transform 1 0 22752 0 -1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _202_
timestamp 1678805552
transform 1 0 11040 0 -1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _203_
timestamp 1678805552
transform 1 0 9216 0 -1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _204_
timestamp 1678805552
transform 1 0 24192 0 -1 9828
box -50 -56 1692 834
use sg13g2_dlhq_1  _205_
timestamp 1678805552
transform -1 0 28896 0 1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _206_
timestamp 1678805552
transform 1 0 10656 0 1 756
box -50 -56 1692 834
use sg13g2_dlhq_1  _207_
timestamp 1678805552
transform 1 0 15168 0 1 756
box -50 -56 1692 834
use sg13g2_dlhq_1  _208_
timestamp 1678805552
transform 1 0 23424 0 1 756
box -50 -56 1692 834
use sg13g2_dlhq_1  _209_
timestamp 1678805552
transform -1 0 27168 0 1 756
box -50 -56 1692 834
use sg13g2_dlhq_1  _210_
timestamp 1678805552
transform 1 0 29088 0 1 756
box -50 -56 1692 834
use sg13g2_dlhq_1  _211_
timestamp 1678805552
transform -1 0 34752 0 1 756
box -50 -56 1692 834
use sg13g2_dlhq_1  _212_
timestamp 1678805552
transform 1 0 28224 0 -1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _213_
timestamp 1678805552
transform 1 0 26400 0 -1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _214_
timestamp 1678805552
transform -1 0 34464 0 1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _215_
timestamp 1678805552
transform 1 0 29952 0 -1 3780
box -50 -56 1692 834
use sg13g2_dlhq_1  _216_
timestamp 1678805552
transform 1 0 25632 0 1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _217_
timestamp 1678805552
transform 1 0 23136 0 -1 3780
box -50 -56 1692 834
use sg13g2_dlhq_1  _218_
timestamp 1678805552
transform 1 0 31584 0 1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _219_
timestamp 1678805552
transform 1 0 30048 0 1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _220_
timestamp 1678805552
transform 1 0 26304 0 -1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _221_
timestamp 1678805552
transform 1 0 28032 0 -1 3780
box -50 -56 1692 834
use sg13g2_dlhq_1  _222_
timestamp 1678805552
transform -1 0 32160 0 1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _223_
timestamp 1678805552
transform -1 0 34368 0 -1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _224_
timestamp 1678805552
transform 1 0 30048 0 1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _225_
timestamp 1678805552
transform 1 0 32448 0 -1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _226_
timestamp 1678805552
transform 1 0 34368 0 -1 3780
box -50 -56 1692 834
use sg13g2_dlhq_1  _227_
timestamp 1678805552
transform -1 0 39648 0 -1 3780
box -50 -56 1692 834
use sg13g2_dlhq_1  _228_
timestamp 1678805552
transform 1 0 36864 0 1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _229_
timestamp 1678805552
transform 1 0 37920 0 -1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _230_
timestamp 1678805552
transform 1 0 33312 0 1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _231_
timestamp 1678805552
transform -1 0 38208 0 -1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _232_
timestamp 1678805552
transform 1 0 9600 0 1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _233_
timestamp 1678805552
transform 1 0 10464 0 -1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _234_
timestamp 1678805552
transform 1 0 12096 0 -1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _235_
timestamp 1678805552
transform 1 0 13728 0 -1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _236_
timestamp 1678805552
transform 1 0 9792 0 -1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _237_
timestamp 1678805552
transform 1 0 8256 0 1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _238_
timestamp 1678805552
transform 1 0 3744 0 -1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _239_
timestamp 1678805552
transform 1 0 1248 0 1 756
box -50 -56 1692 834
use sg13g2_dlhq_1  _240_
timestamp 1678805552
transform -1 0 38016 0 1 756
box -50 -56 1692 834
use sg13g2_dlhq_1  _241_
timestamp 1678805552
transform -1 0 36384 0 1 756
box -50 -56 1692 834
use sg13g2_dlhq_1  _242_
timestamp 1678805552
transform -1 0 39648 0 1 756
box -50 -56 1692 834
use sg13g2_dlhq_1  _243_
timestamp 1678805552
transform -1 0 41760 0 -1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _244_
timestamp 1678805552
transform 1 0 30432 0 -1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _245_
timestamp 1678805552
transform -1 0 34944 0 1 3780
box -50 -56 1692 834
use sg13g2_dlhq_1  _246_
timestamp 1678805552
transform 1 0 34944 0 1 3780
box -50 -56 1692 834
use sg13g2_dlhq_1  _247_
timestamp 1678805552
transform -1 0 40512 0 1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _248_
timestamp 1678805552
transform 1 0 37152 0 1 3780
box -50 -56 1692 834
use sg13g2_dlhq_1  _249_
timestamp 1678805552
transform 1 0 38784 0 1 3780
box -50 -56 1692 834
use sg13g2_dlhq_1  _250_
timestamp 1678805552
transform 1 0 34080 0 -1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _251_
timestamp 1678805552
transform 1 0 35808 0 -1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _252_
timestamp 1678805552
transform 1 0 2112 0 -1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _253_
timestamp 1678805552
transform 1 0 2976 0 1 756
box -50 -56 1692 834
use sg13g2_dlhq_1  _254_
timestamp 1678805552
transform 1 0 7488 0 1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _255_
timestamp 1678805552
transform 1 0 5856 0 1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _256_
timestamp 1678805552
transform 1 0 1440 0 1 3780
box -50 -56 1692 834
use sg13g2_dlhq_1  _257_
timestamp 1678805552
transform 1 0 1536 0 -1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _258_
timestamp 1678805552
transform 1 0 1440 0 1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _259_
timestamp 1678805552
transform 1 0 1536 0 -1 3780
box -50 -56 1692 834
use sg13g2_dlhq_1  _260_
timestamp 1678805552
transform 1 0 1536 0 1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _261_
timestamp 1678805552
transform 1 0 1344 0 -1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _262_
timestamp 1678805552
transform 1 0 1440 0 -1 9828
box -50 -56 1692 834
use sg13g2_dlhq_1  _263_
timestamp 1678805552
transform 1 0 1632 0 -1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _264_
timestamp 1678805552
transform 1 0 1536 0 1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _265_
timestamp 1678805552
transform 1 0 3936 0 -1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _266_
timestamp 1678805552
transform 1 0 4704 0 1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _267_
timestamp 1678805552
transform 1 0 5856 0 -1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _268_
timestamp 1678805552
transform 1 0 7488 0 -1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _269_
timestamp 1678805552
transform 1 0 6336 0 1 8316
box -50 -56 1692 834
use sg13g2_dfrbpq_1  _270_
timestamp 1746535128
transform 1 0 33504 0 1 8316
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _271_
timestamp 1746535128
transform 1 0 33984 0 -1 8316
box -48 -56 2640 834
use sg13g2_tiehi  _272_
timestamp 1680000651
transform 1 0 33120 0 -1 9828
box -48 -56 432 834
use sg13g2_tiehi  _273_
timestamp 1680000651
transform -1 0 35136 0 -1 9828
box -48 -56 432 834
use sg13g2_buf_1  _274_
timestamp 1676381911
transform 1 0 41184 0 1 756
box -48 -56 432 834
use sg13g2_buf_1  _275_
timestamp 1676381911
transform 1 0 40416 0 1 756
box -48 -56 432 834
use sg13g2_buf_1  _276_
timestamp 1676381911
transform 1 0 40032 0 1 756
box -48 -56 432 834
use sg13g2_buf_1  _277_
timestamp 1676381911
transform 1 0 40032 0 -1 3780
box -48 -56 432 834
use sg13g2_buf_1  _278_
timestamp 1676381911
transform 1 0 38496 0 1 2268
box -48 -56 432 834
use sg13g2_buf_1  _279_
timestamp 1676381911
transform 1 0 40800 0 1 756
box -48 -56 432 834
use sg13g2_buf_1  _280_
timestamp 1676381911
transform 1 0 41184 0 -1 3780
box -48 -56 432 834
use sg13g2_buf_1  _281_
timestamp 1676381911
transform 1 0 41184 0 1 2268
box -48 -56 432 834
use sg13g2_buf_1  _282_
timestamp 1676381911
transform 1 0 40800 0 1 2268
box -48 -56 432 834
use sg13g2_buf_1  _283_
timestamp 1676381911
transform 1 0 40416 0 -1 3780
box -48 -56 432 834
use sg13g2_buf_1  _284_
timestamp 1676381911
transform 1 0 40800 0 -1 3780
box -48 -56 432 834
use sg13g2_buf_1  _285_
timestamp 1676381911
transform 1 0 41184 0 1 3780
box -48 -56 432 834
use sg13g2_buf_1  _286_
timestamp 1676381911
transform 1 0 40416 0 1 3780
box -48 -56 432 834
use sg13g2_buf_1  _287_
timestamp 1676381911
transform 1 0 40800 0 1 3780
box -48 -56 432 834
use sg13g2_buf_1  _288_
timestamp 1676381911
transform 1 0 41184 0 -1 5292
box -48 -56 432 834
use sg13g2_buf_1  _289_
timestamp 1676381911
transform 1 0 40416 0 -1 5292
box -48 -56 432 834
use sg13g2_buf_1  _290_
timestamp 1676381911
transform 1 0 40800 0 -1 5292
box -48 -56 432 834
use sg13g2_buf_1  _291_
timestamp 1676381911
transform 1 0 40416 0 1 5292
box -48 -56 432 834
use sg13g2_buf_1  _292_
timestamp 1676381911
transform 1 0 40800 0 1 5292
box -48 -56 432 834
use sg13g2_buf_1  _293_
timestamp 1676381911
transform 1 0 40800 0 -1 6804
box -48 -56 432 834
use sg13g2_buf_1  _294_
timestamp 1676381911
transform 1 0 40416 0 -1 6804
box -48 -56 432 834
use sg13g2_buf_1  _295_
timestamp 1676381911
transform 1 0 40800 0 1 6804
box -48 -56 432 834
use sg13g2_buf_1  _296_
timestamp 1676381911
transform 1 0 40416 0 1 6804
box -48 -56 432 834
use sg13g2_buf_1  _297_
timestamp 1676381911
transform 1 0 40800 0 -1 8316
box -48 -56 432 834
use sg13g2_buf_1  _298_
timestamp 1676381911
transform 1 0 40416 0 -1 8316
box -48 -56 432 834
use sg13g2_buf_1  _299_
timestamp 1676381911
transform 1 0 41184 0 -1 8316
box -48 -56 432 834
use sg13g2_buf_1  _300_
timestamp 1676381911
transform 1 0 40800 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  _301_
timestamp 1676381911
transform 1 0 41184 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  _302_
timestamp 1676381911
transform 1 0 40800 0 -1 9828
box -48 -56 432 834
use sg13g2_buf_1  _303_
timestamp 1676381911
transform 1 0 39744 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  _304_
timestamp 1676381911
transform 1 0 41184 0 -1 9828
box -48 -56 432 834
use sg13g2_buf_1  _305_
timestamp 1676381911
transform 1 0 40416 0 -1 9828
box -48 -56 432 834
use sg13g2_buf_1  _306_
timestamp 1676381911
transform -1 0 19776 0 -1 9828
box -48 -56 432 834
use sg13g2_buf_1  _307_
timestamp 1676381911
transform 1 0 19776 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  _308_
timestamp 1676381911
transform 1 0 21120 0 -1 9828
box -48 -56 432 834
use sg13g2_buf_1  _309_
timestamp 1676381911
transform 1 0 22272 0 -1 8316
box -48 -56 432 834
use sg13g2_buf_1  _310_
timestamp 1676381911
transform -1 0 30048 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  _311_
timestamp 1676381911
transform -1 0 32352 0 -1 9828
box -48 -56 432 834
use sg13g2_buf_1  _312_
timestamp 1676381911
transform -1 0 30912 0 -1 8316
box -48 -56 432 834
use sg13g2_buf_1  _313_
timestamp 1676381911
transform -1 0 32736 0 -1 9828
box -48 -56 432 834
use sg13g2_buf_1  _314_
timestamp 1676381911
transform -1 0 32064 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  _315_
timestamp 1676381911
transform -1 0 33120 0 -1 9828
box -48 -56 432 834
use sg13g2_buf_1  _316_
timestamp 1676381911
transform -1 0 32448 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  _317_
timestamp 1676381911
transform -1 0 32832 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  _318_
timestamp 1676381911
transform -1 0 33216 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  _319_
timestamp 1676381911
transform 1 0 33024 0 -1 8316
box -48 -56 432 834
use sg13g2_buf_1  _320_
timestamp 1676381911
transform -1 0 36480 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  _321_
timestamp 1676381911
transform -1 0 36864 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  _322_
timestamp 1676381911
transform -1 0 38016 0 -1 9828
box -48 -56 432 834
use sg13g2_buf_1  _323_
timestamp 1676381911
transform 1 0 38496 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  _324_
timestamp 1676381911
transform 1 0 38880 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  _325_
timestamp 1676381911
transform 1 0 40128 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  _326_
timestamp 1676381911
transform 1 0 10560 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _327_
timestamp 1676381911
transform -1 0 24384 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _328_
timestamp 1676381911
transform 1 0 19776 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _329_
timestamp 1676381911
transform -1 0 31104 0 1 756
box -48 -56 432 834
use sg13g2_buf_1  _330_
timestamp 1676381911
transform -1 0 20832 0 1 2268
box -48 -56 432 834
use sg13g2_buf_1  _331_
timestamp 1676381911
transform 1 0 12960 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _332_
timestamp 1676381911
transform 1 0 20160 0 1 5292
box -48 -56 432 834
use sg13g2_buf_1  _333_
timestamp 1676381911
transform -1 0 21504 0 1 6804
box -48 -56 432 834
use sg13g2_buf_1  _334_
timestamp 1676381911
transform -1 0 21696 0 -1 8316
box -48 -56 432 834
use sg13g2_buf_1  _335_
timestamp 1676381911
transform 1 0 20640 0 -1 5292
box -48 -56 432 834
use sg13g2_buf_1  _336_
timestamp 1676381911
transform 1 0 21024 0 -1 5292
box -48 -56 432 834
use sg13g2_buf_1  _337_
timestamp 1676381911
transform 1 0 20832 0 1 2268
box -48 -56 432 834
use sg13g2_buf_1  _338_
timestamp 1676381911
transform -1 0 22272 0 1 2268
box -48 -56 432 834
use sg13g2_buf_1  _339_
timestamp 1676381911
transform 1 0 21408 0 1 2268
box -48 -56 432 834
use sg13g2_buf_1  _340_
timestamp 1676381911
transform -1 0 23808 0 -1 6804
box -48 -56 432 834
use sg13g2_buf_1  _341_
timestamp 1676381911
transform -1 0 30816 0 1 6804
box -48 -56 432 834
use sg13g2_buf_1  _342_
timestamp 1676381911
transform -1 0 23520 0 1 6804
box -48 -56 432 834
use sg13g2_buf_1  _343_
timestamp 1676381911
transform -1 0 23328 0 1 3780
box -48 -56 432 834
use sg13g2_buf_1  _344_
timestamp 1676381911
transform 1 0 22848 0 1 2268
box -48 -56 432 834
use sg13g2_buf_1  _345_
timestamp 1676381911
transform -1 0 30336 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _346_
timestamp 1676381911
transform -1 0 24192 0 1 3780
box -48 -56 432 834
use sg13g2_buf_1  _347_
timestamp 1676381911
transform 1 0 22848 0 1 756
box -48 -56 432 834
use sg13g2_buf_1  _348_
timestamp 1676381911
transform -1 0 26400 0 -1 6804
box -48 -56 432 834
use sg13g2_buf_1  _349_
timestamp 1676381911
transform 1 0 23232 0 1 2268
box -48 -56 432 834
use sg13g2_buf_1  _350_
timestamp 1676381911
transform -1 0 25632 0 -1 5292
box -48 -56 432 834
use sg13g2_buf_1  _351_
timestamp 1676381911
transform 1 0 23424 0 1 3780
box -48 -56 432 834
use sg13g2_buf_1  _352_
timestamp 1676381911
transform -1 0 27552 0 -1 8316
box -48 -56 432 834
use sg13g2_buf_1  _353_
timestamp 1676381911
transform 1 0 24576 0 1 2268
box -48 -56 432 834
use sg13g2_buf_1  _354_
timestamp 1676381911
transform -1 0 26976 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _355_
timestamp 1676381911
transform -1 0 32736 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _356_
timestamp 1676381911
transform -1 0 29856 0 1 5292
box -48 -56 432 834
use sg13g2_buf_1  _357_
timestamp 1676381911
transform -1 0 34752 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _358_
timestamp 1676381911
transform 1 0 25248 0 1 2268
box -48 -56 432 834
use sg13g2_buf_1  _359_
timestamp 1676381911
transform -1 0 32448 0 -1 6804
box -48 -56 432 834
use sg13g2_buf_1  _360_
timestamp 1676381911
transform -1 0 29760 0 1 3780
box -48 -56 432 834
use sg13g2_buf_1  _361_
timestamp 1676381911
transform -1 0 32832 0 1 2268
box -48 -56 432 834
use sg13g2_buf_1  _362_
timestamp 1676381911
transform -1 0 33312 0 1 3780
box -48 -56 432 834
use sg13g2_buf_1  _363_
timestamp 1676381911
transform -1 0 38304 0 1 2268
box -48 -56 432 834
use sg13g2_buf_1  _364_
timestamp 1676381911
transform -1 0 39936 0 -1 6804
box -48 -56 432 834
use sg13g2_buf_1  _365_
timestamp 1676381911
transform -1 0 36672 0 -1 6804
box -48 -56 432 834
use sg13g2_buf_1  _366_
timestamp 1676381911
transform 1 0 25824 0 1 6804
box -48 -56 432 834
use sg13g2_buf_1  _367_
timestamp 1676381911
transform 1 0 26784 0 1 5292
box -48 -56 432 834
use sg13g2_buf_1  _368_
timestamp 1676381911
transform 1 0 26976 0 1 3780
box -48 -56 432 834
use sg13g2_buf_1  _369_
timestamp 1676381911
transform 1 0 27168 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _370_
timestamp 1676381911
transform -1 0 35904 0 1 2268
box -48 -56 432 834
use sg13g2_buf_1  _371_
timestamp 1676381911
transform -1 0 40032 0 1 756
box -48 -56 432 834
use sg13g2_buf_1  _372_
timestamp 1676381911
transform -1 0 32928 0 1 3780
box -48 -56 432 834
use sg13g2_buf_1  _373_
timestamp 1676381911
transform -1 0 37824 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _374_
timestamp 1676381911
transform -1 0 40032 0 -1 3780
box -48 -56 432 834
use sg13g2_buf_1  _375_
timestamp 1676381911
transform -1 0 36960 0 1 3780
box -48 -56 432 834
use sg13g2_buf_1  _376_
timestamp 1676381911
transform 1 0 28416 0 1 756
box -48 -56 432 834
use sg13g2_buf_1  _377_
timestamp 1676381911
transform -1 0 29952 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _378_
timestamp 1676381911
transform -1 0 29568 0 1 8316
box -48 -56 432 834
use sg13g2_buf_8  clkbuf_0_UserCLK_regs
timestamp 1676451365
transform -1 0 36384 0 -1 9828
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_0_UserCLK
timestamp 1676451365
transform -1 0 31968 0 -1 9828
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_1_0__f_UserCLK
timestamp 1676451365
transform -1 0 30720 0 -1 9828
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_1_0__f_UserCLK_regs
timestamp 1676451365
transform 1 0 36672 0 -1 6804
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_1_1__f_UserCLK_regs
timestamp 1676451365
transform -1 0 34752 0 -1 9828
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_regs_0_UserCLK
timestamp 1676451365
transform 1 0 36384 0 -1 9828
box -48 -56 1296 834
use sg13g2_fill_1  FILLER_0_0
timestamp 1677579658
transform 1 0 1152 0 1 756
box -48 -56 144 834
use sg13g2_fill_1  FILLER_0_18
timestamp 1677579658
transform 1 0 2880 0 1 756
box -48 -56 144 834
use sg13g2_decap_4  FILLER_0_36
timestamp 1679577901
transform 1 0 4608 0 1 756
box -48 -56 432 834
use sg13g2_fill_1  FILLER_0_40
timestamp 1677579658
transform 1 0 4992 0 1 756
box -48 -56 144 834
use sg13g2_decap_8  FILLER_0_62
timestamp 1679581782
transform 1 0 7104 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_69
timestamp 1679581782
transform 1 0 7776 0 1 756
box -48 -56 720 834
use sg13g2_decap_4  FILLER_0_76
timestamp 1679577901
transform 1 0 8448 0 1 756
box -48 -56 432 834
use sg13g2_fill_2  FILLER_0_80
timestamp 1677580104
transform 1 0 8832 0 1 756
box -48 -56 240 834
use sg13g2_decap_8  FILLER_0_133
timestamp 1679581782
transform 1 0 13920 0 1 756
box -48 -56 720 834
use sg13g2_decap_4  FILLER_0_140
timestamp 1679577901
transform 1 0 14592 0 1 756
box -48 -56 432 834
use sg13g2_fill_2  FILLER_0_144
timestamp 1677580104
transform 1 0 14976 0 1 756
box -48 -56 240 834
use sg13g2_decap_4  FILLER_0_163
timestamp 1679577901
transform 1 0 16800 0 1 756
box -48 -56 432 834
use sg13g2_fill_1  FILLER_0_167
timestamp 1677579658
transform 1 0 17184 0 1 756
box -48 -56 144 834
use sg13g2_fill_1  FILLER_0_202
timestamp 1677579658
transform 1 0 20544 0 1 756
box -48 -56 144 834
use sg13g2_decap_4  FILLER_0_220
timestamp 1679577901
transform 1 0 22272 0 1 756
box -48 -56 432 834
use sg13g2_fill_2  FILLER_0_224
timestamp 1677580104
transform 1 0 22656 0 1 756
box -48 -56 240 834
use sg13g2_fill_2  FILLER_0_230
timestamp 1677580104
transform 1 0 23232 0 1 756
box -48 -56 240 834
use sg13g2_decap_4  FILLER_0_249
timestamp 1679577901
transform 1 0 25056 0 1 756
box -48 -56 432 834
use sg13g2_fill_1  FILLER_0_253
timestamp 1677579658
transform 1 0 25440 0 1 756
box -48 -56 144 834
use sg13g2_decap_8  FILLER_0_271
timestamp 1679581782
transform 1 0 27168 0 1 756
box -48 -56 720 834
use sg13g2_decap_4  FILLER_0_278
timestamp 1679577901
transform 1 0 27840 0 1 756
box -48 -56 432 834
use sg13g2_fill_2  FILLER_0_282
timestamp 1677580104
transform 1 0 28224 0 1 756
box -48 -56 240 834
use sg13g2_fill_2  FILLER_0_288
timestamp 1677580104
transform 1 0 28800 0 1 756
box -48 -56 240 834
use sg13g2_fill_1  FILLER_0_290
timestamp 1677579658
transform 1 0 28992 0 1 756
box -48 -56 144 834
use sg13g2_fill_2  FILLER_0_421
timestamp 1677580104
transform 1 0 41568 0 1 756
box -48 -56 240 834
use sg13g2_fill_1  FILLER_0_423
timestamp 1677579658
transform 1 0 41760 0 1 756
box -48 -56 144 834
use sg13g2_decap_8  FILLER_1_0
timestamp 1679581782
transform 1 0 1152 0 -1 2268
box -48 -56 720 834
use sg13g2_fill_2  FILLER_1_7
timestamp 1677580104
transform 1 0 1824 0 -1 2268
box -48 -56 240 834
use sg13g2_fill_1  FILLER_1_9
timestamp 1677579658
transform 1 0 2016 0 -1 2268
box -48 -56 144 834
use sg13g2_fill_2  FILLER_1_65
timestamp 1677580104
transform 1 0 7392 0 -1 2268
box -48 -56 240 834
use sg13g2_fill_1  FILLER_1_67
timestamp 1677579658
transform 1 0 7584 0 -1 2268
box -48 -56 144 834
use sg13g2_decap_8  FILLER_1_89
timestamp 1679581782
transform 1 0 9696 0 -1 2268
box -48 -56 720 834
use sg13g2_fill_2  FILLER_1_96
timestamp 1677580104
transform 1 0 10368 0 -1 2268
box -48 -56 240 834
use sg13g2_fill_2  FILLER_1_165
timestamp 1677580104
transform 1 0 16992 0 -1 2268
box -48 -56 240 834
use sg13g2_fill_1  FILLER_1_167
timestamp 1677579658
transform 1 0 17184 0 -1 2268
box -48 -56 144 834
use sg13g2_decap_4  FILLER_1_189
timestamp 1679577901
transform 1 0 19296 0 -1 2268
box -48 -56 432 834
use sg13g2_fill_1  FILLER_1_193
timestamp 1677579658
transform 1 0 19680 0 -1 2268
box -48 -56 144 834
use sg13g2_fill_2  FILLER_1_219
timestamp 1677580104
transform 1 0 22176 0 -1 2268
box -48 -56 240 834
use sg13g2_fill_2  FILLER_1_242
timestamp 1677580104
transform 1 0 24384 0 -1 2268
box -48 -56 240 834
use sg13g2_fill_2  FILLER_1_269
timestamp 1677580104
transform 1 0 26976 0 -1 2268
box -48 -56 240 834
use sg13g2_decap_4  FILLER_1_350
timestamp 1679577901
transform 1 0 34752 0 -1 2268
box -48 -56 432 834
use sg13g2_fill_2  FILLER_1_375
timestamp 1677580104
transform 1 0 37152 0 -1 2268
box -48 -56 240 834
use sg13g2_fill_1  FILLER_1_377
timestamp 1677579658
transform 1 0 37344 0 -1 2268
box -48 -56 144 834
use sg13g2_fill_2  FILLER_1_382
timestamp 1677580104
transform 1 0 37824 0 -1 2268
box -48 -56 240 834
use sg13g2_fill_1  FILLER_1_384
timestamp 1677579658
transform 1 0 38016 0 -1 2268
box -48 -56 144 834
use sg13g2_fill_1  FILLER_1_423
timestamp 1677579658
transform 1 0 41760 0 -1 2268
box -48 -56 144 834
use sg13g2_fill_2  FILLER_2_0
timestamp 1677580104
transform 1 0 1152 0 1 2268
box -48 -56 240 834
use sg13g2_fill_1  FILLER_2_2
timestamp 1677579658
transform 1 0 1344 0 1 2268
box -48 -56 144 834
use sg13g2_fill_1  FILLER_2_20
timestamp 1677579658
transform 1 0 3072 0 1 2268
box -48 -56 144 834
use sg13g2_fill_2  FILLER_2_36
timestamp 1677580104
transform 1 0 4608 0 1 2268
box -48 -56 240 834
use sg13g2_decap_4  FILLER_2_43
timestamp 1679577901
transform 1 0 5280 0 1 2268
box -48 -56 432 834
use sg13g2_fill_2  FILLER_2_47
timestamp 1677580104
transform 1 0 5664 0 1 2268
box -48 -56 240 834
use sg13g2_decap_8  FILLER_2_121
timestamp 1679581782
transform 1 0 12768 0 1 2268
box -48 -56 720 834
use sg13g2_fill_2  FILLER_2_128
timestamp 1677580104
transform 1 0 13440 0 1 2268
box -48 -56 240 834
use sg13g2_fill_1  FILLER_2_130
timestamp 1677579658
transform 1 0 13632 0 1 2268
box -48 -56 144 834
use sg13g2_fill_1  FILLER_2_152
timestamp 1677579658
transform 1 0 15744 0 1 2268
box -48 -56 144 834
use sg13g2_decap_4  FILLER_2_170
timestamp 1679577901
transform 1 0 17472 0 1 2268
box -48 -56 432 834
use sg13g2_fill_2  FILLER_2_209
timestamp 1677580104
transform 1 0 21216 0 1 2268
box -48 -56 240 834
use sg13g2_fill_1  FILLER_2_215
timestamp 1677579658
transform 1 0 21792 0 1 2268
box -48 -56 144 834
use sg13g2_decap_4  FILLER_2_220
timestamp 1679577901
transform 1 0 22272 0 1 2268
box -48 -56 432 834
use sg13g2_fill_2  FILLER_2_224
timestamp 1677580104
transform 1 0 22656 0 1 2268
box -48 -56 240 834
use sg13g2_fill_2  FILLER_2_248
timestamp 1677580104
transform 1 0 24960 0 1 2268
box -48 -56 240 834
use sg13g2_fill_1  FILLER_2_250
timestamp 1677579658
transform 1 0 25152 0 1 2268
box -48 -56 144 834
use sg13g2_fill_2  FILLER_2_323
timestamp 1677580104
transform 1 0 32160 0 1 2268
box -48 -56 240 834
use sg13g2_fill_1  FILLER_2_325
timestamp 1677579658
transform 1 0 32352 0 1 2268
box -48 -56 144 834
use sg13g2_decap_8  FILLER_2_347
timestamp 1679581782
transform 1 0 34464 0 1 2268
box -48 -56 720 834
use sg13g2_decap_4  FILLER_2_354
timestamp 1679577901
transform 1 0 35136 0 1 2268
box -48 -56 432 834
use sg13g2_fill_2  FILLER_2_387
timestamp 1677580104
transform 1 0 38304 0 1 2268
box -48 -56 240 834
use sg13g2_fill_2  FILLER_2_410
timestamp 1677580104
transform 1 0 40512 0 1 2268
box -48 -56 240 834
use sg13g2_fill_1  FILLER_2_412
timestamp 1677579658
transform 1 0 40704 0 1 2268
box -48 -56 144 834
use sg13g2_fill_2  FILLER_2_421
timestamp 1677580104
transform 1 0 41568 0 1 2268
box -48 -56 240 834
use sg13g2_fill_1  FILLER_2_423
timestamp 1677579658
transform 1 0 41760 0 1 2268
box -48 -56 144 834
use sg13g2_decap_4  FILLER_3_0
timestamp 1679577901
transform 1 0 1152 0 -1 3780
box -48 -56 432 834
use sg13g2_fill_1  FILLER_3_33
timestamp 1677579658
transform 1 0 4320 0 -1 3780
box -48 -56 144 834
use sg13g2_fill_2  FILLER_3_75
timestamp 1677580104
transform 1 0 8352 0 -1 3780
box -48 -56 240 834
use sg13g2_fill_1  FILLER_3_77
timestamp 1677579658
transform 1 0 8544 0 -1 3780
box -48 -56 144 834
use sg13g2_decap_8  FILLER_3_95
timestamp 1679581782
transform 1 0 10272 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_123
timestamp 1679581782
transform 1 0 12960 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_4  FILLER_3_130
timestamp 1679577901
transform 1 0 13632 0 -1 3780
box -48 -56 432 834
use sg13g2_fill_1  FILLER_3_134
timestamp 1677579658
transform 1 0 14016 0 -1 3780
box -48 -56 144 834
use sg13g2_decap_4  FILLER_3_152
timestamp 1679577901
transform 1 0 15744 0 -1 3780
box -48 -56 432 834
use sg13g2_decap_8  FILLER_3_177
timestamp 1679581782
transform 1 0 18144 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_184
timestamp 1679581782
transform 1 0 18816 0 -1 3780
box -48 -56 720 834
use sg13g2_fill_1  FILLER_3_191
timestamp 1677579658
transform 1 0 19488 0 -1 3780
box -48 -56 144 834
use sg13g2_fill_1  FILLER_3_209
timestamp 1677579658
transform 1 0 21216 0 -1 3780
box -48 -56 144 834
use sg13g2_fill_2  FILLER_3_227
timestamp 1677580104
transform 1 0 22944 0 -1 3780
box -48 -56 240 834
use sg13g2_decap_8  FILLER_3_267
timestamp 1679581782
transform 1 0 26784 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_4  FILLER_3_274
timestamp 1679577901
transform 1 0 27456 0 -1 3780
box -48 -56 432 834
use sg13g2_fill_2  FILLER_3_278
timestamp 1677580104
transform 1 0 27840 0 -1 3780
box -48 -56 240 834
use sg13g2_fill_2  FILLER_3_297
timestamp 1677580104
transform 1 0 29664 0 -1 3780
box -48 -56 240 834
use sg13g2_fill_1  FILLER_3_299
timestamp 1677579658
transform 1 0 29856 0 -1 3780
box -48 -56 144 834
use sg13g2_decap_8  FILLER_3_338
timestamp 1679581782
transform 1 0 33600 0 -1 3780
box -48 -56 720 834
use sg13g2_fill_1  FILLER_3_345
timestamp 1677579658
transform 1 0 34272 0 -1 3780
box -48 -56 144 834
use sg13g2_fill_2  FILLER_3_421
timestamp 1677580104
transform 1 0 41568 0 -1 3780
box -48 -56 240 834
use sg13g2_fill_1  FILLER_3_423
timestamp 1677579658
transform 1 0 41760 0 -1 3780
box -48 -56 144 834
use sg13g2_fill_2  FILLER_4_0
timestamp 1677580104
transform 1 0 1152 0 1 3780
box -48 -56 240 834
use sg13g2_fill_1  FILLER_4_2
timestamp 1677579658
transform 1 0 1344 0 1 3780
box -48 -56 144 834
use sg13g2_fill_2  FILLER_4_20
timestamp 1677580104
transform 1 0 3072 0 1 3780
box -48 -56 240 834
use sg13g2_fill_1  FILLER_4_22
timestamp 1677579658
transform 1 0 3264 0 1 3780
box -48 -56 144 834
use sg13g2_fill_2  FILLER_4_43
timestamp 1677580104
transform 1 0 5280 0 1 3780
box -48 -56 240 834
use sg13g2_decap_4  FILLER_4_66
timestamp 1679577901
transform 1 0 7488 0 1 3780
box -48 -56 432 834
use sg13g2_fill_1  FILLER_4_70
timestamp 1677579658
transform 1 0 7872 0 1 3780
box -48 -56 144 834
use sg13g2_decap_8  FILLER_4_88
timestamp 1679581782
transform 1 0 9600 0 1 3780
box -48 -56 720 834
use sg13g2_fill_1  FILLER_4_95
timestamp 1677579658
transform 1 0 10272 0 1 3780
box -48 -56 144 834
use sg13g2_fill_2  FILLER_4_130
timestamp 1677580104
transform 1 0 13632 0 1 3780
box -48 -56 240 834
use sg13g2_decap_8  FILLER_4_153
timestamp 1679581782
transform 1 0 15840 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_160
timestamp 1679581782
transform 1 0 16512 0 1 3780
box -48 -56 720 834
use sg13g2_fill_1  FILLER_4_167
timestamp 1677579658
transform 1 0 17184 0 1 3780
box -48 -56 144 834
use sg13g2_fill_2  FILLER_4_185
timestamp 1677580104
transform 1 0 18912 0 1 3780
box -48 -56 240 834
use sg13g2_fill_1  FILLER_4_187
timestamp 1677579658
transform 1 0 19104 0 1 3780
box -48 -56 144 834
use sg13g2_fill_1  FILLER_4_205
timestamp 1677579658
transform 1 0 20832 0 1 3780
box -48 -56 144 834
use sg13g2_fill_1  FILLER_4_231
timestamp 1677579658
transform 1 0 23328 0 1 3780
box -48 -56 144 834
use sg13g2_decap_8  FILLER_4_257
timestamp 1679581782
transform 1 0 25824 0 1 3780
box -48 -56 720 834
use sg13g2_decap_4  FILLER_4_264
timestamp 1679577901
transform 1 0 26496 0 1 3780
box -48 -56 432 834
use sg13g2_fill_1  FILLER_4_268
timestamp 1677579658
transform 1 0 26880 0 1 3780
box -48 -56 144 834
use sg13g2_decap_8  FILLER_4_298
timestamp 1679581782
transform 1 0 29760 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_315
timestamp 1679581782
transform 1 0 31392 0 1 3780
box -48 -56 720 834
use sg13g2_decap_4  FILLER_4_322
timestamp 1679577901
transform 1 0 32064 0 1 3780
box -48 -56 432 834
use sg13g2_fill_1  FILLER_4_326
timestamp 1677579658
transform 1 0 32448 0 1 3780
box -48 -56 144 834
use sg13g2_fill_2  FILLER_4_373
timestamp 1677580104
transform 1 0 36960 0 1 3780
box -48 -56 240 834
use sg13g2_fill_2  FILLER_4_421
timestamp 1677580104
transform 1 0 41568 0 1 3780
box -48 -56 240 834
use sg13g2_fill_1  FILLER_4_423
timestamp 1677579658
transform 1 0 41760 0 1 3780
box -48 -56 144 834
use sg13g2_decap_4  FILLER_5_0
timestamp 1679577901
transform 1 0 1152 0 -1 5292
box -48 -56 432 834
use sg13g2_decap_4  FILLER_5_21
timestamp 1679577901
transform 1 0 3168 0 -1 5292
box -48 -56 432 834
use sg13g2_fill_2  FILLER_5_38
timestamp 1677580104
transform 1 0 4800 0 -1 5292
box -48 -56 240 834
use sg13g2_decap_8  FILLER_5_65
timestamp 1679581782
transform 1 0 7392 0 -1 5292
box -48 -56 720 834
use sg13g2_fill_2  FILLER_5_72
timestamp 1677580104
transform 1 0 8064 0 -1 5292
box -48 -56 240 834
use sg13g2_fill_2  FILLER_5_101
timestamp 1677580104
transform 1 0 10848 0 -1 5292
box -48 -56 240 834
use sg13g2_decap_8  FILLER_5_120
timestamp 1679581782
transform 1 0 12672 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_4  FILLER_5_127
timestamp 1679577901
transform 1 0 13344 0 -1 5292
box -48 -56 432 834
use sg13g2_decap_8  FILLER_5_152
timestamp 1679581782
transform 1 0 15744 0 -1 5292
box -48 -56 720 834
use sg13g2_fill_2  FILLER_5_159
timestamp 1677580104
transform 1 0 16416 0 -1 5292
box -48 -56 240 834
use sg13g2_fill_2  FILLER_5_211
timestamp 1677580104
transform 1 0 21408 0 -1 5292
box -48 -56 240 834
use sg13g2_decap_8  FILLER_5_255
timestamp 1679581782
transform 1 0 25632 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_279
timestamp 1679581782
transform 1 0 27936 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_4  FILLER_5_286
timestamp 1679577901
transform 1 0 28608 0 -1 5292
box -48 -56 432 834
use sg13g2_decap_8  FILLER_5_307
timestamp 1679581782
transform 1 0 30624 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_4  FILLER_5_314
timestamp 1679577901
transform 1 0 31296 0 -1 5292
box -48 -56 432 834
use sg13g2_fill_1  FILLER_5_318
timestamp 1677579658
transform 1 0 31680 0 -1 5292
box -48 -56 144 834
use sg13g2_fill_2  FILLER_5_340
timestamp 1677580104
transform 1 0 33792 0 -1 5292
box -48 -56 240 834
use sg13g2_fill_1  FILLER_5_342
timestamp 1677579658
transform 1 0 33984 0 -1 5292
box -48 -56 144 834
use sg13g2_fill_1  FILLER_5_360
timestamp 1677579658
transform 1 0 35712 0 -1 5292
box -48 -56 144 834
use sg13g2_decap_8  FILLER_5_378
timestamp 1679581782
transform 1 0 37440 0 -1 5292
box -48 -56 720 834
use sg13g2_fill_2  FILLER_5_406
timestamp 1677580104
transform 1 0 40128 0 -1 5292
box -48 -56 240 834
use sg13g2_fill_1  FILLER_5_408
timestamp 1677579658
transform 1 0 40320 0 -1 5292
box -48 -56 144 834
use sg13g2_fill_2  FILLER_5_421
timestamp 1677580104
transform 1 0 41568 0 -1 5292
box -48 -56 240 834
use sg13g2_fill_1  FILLER_5_423
timestamp 1677579658
transform 1 0 41760 0 -1 5292
box -48 -56 144 834
use sg13g2_decap_4  FILLER_6_0
timestamp 1679577901
transform 1 0 1152 0 1 5292
box -48 -56 432 834
use sg13g2_decap_8  FILLER_6_21
timestamp 1679581782
transform 1 0 3168 0 1 5292
box -48 -56 720 834
use sg13g2_fill_2  FILLER_6_28
timestamp 1677580104
transform 1 0 3840 0 1 5292
box -48 -56 240 834
use sg13g2_decap_8  FILLER_6_66
timestamp 1679581782
transform 1 0 7488 0 1 5292
box -48 -56 720 834
use sg13g2_fill_1  FILLER_6_73
timestamp 1677579658
transform 1 0 8160 0 1 5292
box -48 -56 144 834
use sg13g2_decap_8  FILLER_6_112
timestamp 1679581782
transform 1 0 11904 0 1 5292
box -48 -56 720 834
use sg13g2_decap_4  FILLER_6_119
timestamp 1679577901
transform 1 0 12576 0 1 5292
box -48 -56 432 834
use sg13g2_fill_1  FILLER_6_123
timestamp 1677579658
transform 1 0 12960 0 1 5292
box -48 -56 144 834
use sg13g2_decap_4  FILLER_6_192
timestamp 1679577901
transform 1 0 19584 0 1 5292
box -48 -56 432 834
use sg13g2_fill_2  FILLER_6_196
timestamp 1677580104
transform 1 0 19968 0 1 5292
box -48 -56 240 834
use sg13g2_decap_8  FILLER_6_202
timestamp 1679581782
transform 1 0 20544 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_209
timestamp 1679581782
transform 1 0 21216 0 1 5292
box -48 -56 720 834
use sg13g2_fill_1  FILLER_6_216
timestamp 1677579658
transform 1 0 21888 0 1 5292
box -48 -56 144 834
use sg13g2_fill_1  FILLER_6_234
timestamp 1677579658
transform 1 0 23616 0 1 5292
box -48 -56 144 834
use sg13g2_decap_8  FILLER_6_256
timestamp 1679581782
transform 1 0 25728 0 1 5292
box -48 -56 720 834
use sg13g2_decap_4  FILLER_6_263
timestamp 1679577901
transform 1 0 26400 0 1 5292
box -48 -56 432 834
use sg13g2_fill_2  FILLER_6_271
timestamp 1677580104
transform 1 0 27168 0 1 5292
box -48 -56 240 834
use sg13g2_fill_1  FILLER_6_273
timestamp 1677579658
transform 1 0 27360 0 1 5292
box -48 -56 144 834
use sg13g2_fill_2  FILLER_6_299
timestamp 1677580104
transform 1 0 29856 0 1 5292
box -48 -56 240 834
use sg13g2_decap_8  FILLER_6_339
timestamp 1679581782
transform 1 0 33696 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_346
timestamp 1679581782
transform 1 0 34368 0 1 5292
box -48 -56 720 834
use sg13g2_fill_1  FILLER_6_353
timestamp 1677579658
transform 1 0 35040 0 1 5292
box -48 -56 144 834
use sg13g2_decap_8  FILLER_6_375
timestamp 1679581782
transform 1 0 37152 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_382
timestamp 1679581782
transform 1 0 37824 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_389
timestamp 1679581782
transform 1 0 38496 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_396
timestamp 1679581782
transform 1 0 39168 0 1 5292
box -48 -56 720 834
use sg13g2_decap_4  FILLER_6_403
timestamp 1679577901
transform 1 0 39840 0 1 5292
box -48 -56 432 834
use sg13g2_fill_2  FILLER_6_407
timestamp 1677580104
transform 1 0 40224 0 1 5292
box -48 -56 240 834
use sg13g2_decap_8  FILLER_6_417
timestamp 1679581782
transform 1 0 41184 0 1 5292
box -48 -56 720 834
use sg13g2_decap_4  FILLER_7_0
timestamp 1679577901
transform 1 0 1152 0 -1 6804
box -48 -56 432 834
use sg13g2_fill_1  FILLER_7_4
timestamp 1677579658
transform 1 0 1536 0 -1 6804
box -48 -56 144 834
use sg13g2_fill_1  FILLER_7_22
timestamp 1677579658
transform 1 0 3264 0 -1 6804
box -48 -56 144 834
use sg13g2_fill_1  FILLER_7_65
timestamp 1677579658
transform 1 0 7392 0 -1 6804
box -48 -56 144 834
use sg13g2_decap_8  FILLER_7_83
timestamp 1679581782
transform 1 0 9120 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_107
timestamp 1679581782
transform 1 0 11424 0 -1 6804
box -48 -56 720 834
use sg13g2_fill_1  FILLER_7_114
timestamp 1677579658
transform 1 0 12096 0 -1 6804
box -48 -56 144 834
use sg13g2_decap_8  FILLER_7_132
timestamp 1679581782
transform 1 0 13824 0 -1 6804
box -48 -56 720 834
use sg13g2_fill_2  FILLER_7_139
timestamp 1677580104
transform 1 0 14496 0 -1 6804
box -48 -56 240 834
use sg13g2_decap_8  FILLER_7_158
timestamp 1679581782
transform 1 0 16320 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_165
timestamp 1679581782
transform 1 0 16992 0 -1 6804
box -48 -56 720 834
use sg13g2_fill_1  FILLER_7_172
timestamp 1677579658
transform 1 0 17664 0 -1 6804
box -48 -56 144 834
use sg13g2_decap_4  FILLER_7_236
timestamp 1679577901
transform 1 0 23808 0 -1 6804
box -48 -56 432 834
use sg13g2_fill_1  FILLER_7_240
timestamp 1677579658
transform 1 0 24192 0 -1 6804
box -48 -56 144 834
use sg13g2_fill_1  FILLER_7_258
timestamp 1677579658
transform 1 0 25920 0 -1 6804
box -48 -56 144 834
use sg13g2_fill_2  FILLER_7_280
timestamp 1677580104
transform 1 0 28032 0 -1 6804
box -48 -56 240 834
use sg13g2_decap_4  FILLER_7_299
timestamp 1679577901
transform 1 0 29856 0 -1 6804
box -48 -56 432 834
use sg13g2_fill_2  FILLER_7_303
timestamp 1677580104
transform 1 0 30240 0 -1 6804
box -48 -56 240 834
use sg13g2_decap_8  FILLER_7_343
timestamp 1679581782
transform 1 0 34080 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_350
timestamp 1679581782
transform 1 0 34752 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_357
timestamp 1679581782
transform 1 0 35424 0 -1 6804
box -48 -56 720 834
use sg13g2_fill_2  FILLER_7_364
timestamp 1677580104
transform 1 0 36096 0 -1 6804
box -48 -56 240 834
use sg13g2_decap_4  FILLER_7_404
timestamp 1679577901
transform 1 0 39936 0 -1 6804
box -48 -56 432 834
use sg13g2_fill_1  FILLER_7_408
timestamp 1677579658
transform 1 0 40320 0 -1 6804
box -48 -56 144 834
use sg13g2_decap_8  FILLER_7_417
timestamp 1679581782
transform 1 0 41184 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_0
timestamp 1679581782
transform 1 0 1152 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_7
timestamp 1679581782
transform 1 0 1824 0 1 6804
box -48 -56 720 834
use sg13g2_decap_4  FILLER_8_14
timestamp 1679577901
transform 1 0 2496 0 1 6804
box -48 -56 432 834
use sg13g2_fill_2  FILLER_8_29
timestamp 1677580104
transform 1 0 3936 0 1 6804
box -48 -56 240 834
use sg13g2_fill_1  FILLER_8_31
timestamp 1677579658
transform 1 0 4128 0 1 6804
box -48 -56 144 834
use sg13g2_decap_8  FILLER_8_93
timestamp 1679581782
transform 1 0 10080 0 1 6804
box -48 -56 720 834
use sg13g2_decap_4  FILLER_8_100
timestamp 1679577901
transform 1 0 10752 0 1 6804
box -48 -56 432 834
use sg13g2_decap_4  FILLER_8_125
timestamp 1679577901
transform 1 0 13152 0 1 6804
box -48 -56 432 834
use sg13g2_fill_1  FILLER_8_129
timestamp 1677579658
transform 1 0 13536 0 1 6804
box -48 -56 144 834
use sg13g2_decap_4  FILLER_8_151
timestamp 1679577901
transform 1 0 15648 0 1 6804
box -48 -56 432 834
use sg13g2_fill_2  FILLER_8_155
timestamp 1677580104
transform 1 0 16032 0 1 6804
box -48 -56 240 834
use sg13g2_decap_8  FILLER_8_174
timestamp 1679581782
transform 1 0 17856 0 1 6804
box -48 -56 720 834
use sg13g2_decap_4  FILLER_8_181
timestamp 1679577901
transform 1 0 18528 0 1 6804
box -48 -56 432 834
use sg13g2_fill_2  FILLER_8_185
timestamp 1677580104
transform 1 0 18912 0 1 6804
box -48 -56 240 834
use sg13g2_decap_8  FILLER_8_212
timestamp 1679581782
transform 1 0 21504 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_219
timestamp 1679581782
transform 1 0 22176 0 1 6804
box -48 -56 720 834
use sg13g2_fill_2  FILLER_8_226
timestamp 1677580104
transform 1 0 22848 0 1 6804
box -48 -56 240 834
use sg13g2_fill_1  FILLER_8_228
timestamp 1677579658
transform 1 0 23040 0 1 6804
box -48 -56 144 834
use sg13g2_decap_4  FILLER_8_233
timestamp 1679577901
transform 1 0 23520 0 1 6804
box -48 -56 432 834
use sg13g2_fill_2  FILLER_8_237
timestamp 1677580104
transform 1 0 23904 0 1 6804
box -48 -56 240 834
use sg13g2_fill_1  FILLER_8_256
timestamp 1677579658
transform 1 0 25728 0 1 6804
box -48 -56 144 834
use sg13g2_decap_8  FILLER_8_278
timestamp 1679581782
transform 1 0 27840 0 1 6804
box -48 -56 720 834
use sg13g2_fill_2  FILLER_8_285
timestamp 1677580104
transform 1 0 28512 0 1 6804
box -48 -56 240 834
use sg13g2_fill_1  FILLER_8_287
timestamp 1677579658
transform 1 0 28704 0 1 6804
box -48 -56 144 834
use sg13g2_decap_8  FILLER_8_309
timestamp 1679581782
transform 1 0 30816 0 1 6804
box -48 -56 720 834
use sg13g2_fill_1  FILLER_8_316
timestamp 1677579658
transform 1 0 31488 0 1 6804
box -48 -56 144 834
use sg13g2_fill_1  FILLER_8_334
timestamp 1677579658
transform 1 0 33216 0 1 6804
box -48 -56 144 834
use sg13g2_decap_8  FILLER_8_373
timestamp 1679581782
transform 1 0 36960 0 1 6804
box -48 -56 720 834
use sg13g2_fill_2  FILLER_8_380
timestamp 1677580104
transform 1 0 37632 0 1 6804
box -48 -56 240 834
use sg13g2_decap_4  FILLER_8_403
timestamp 1679577901
transform 1 0 39840 0 1 6804
box -48 -56 432 834
use sg13g2_fill_2  FILLER_8_407
timestamp 1677580104
transform 1 0 40224 0 1 6804
box -48 -56 240 834
use sg13g2_decap_8  FILLER_8_417
timestamp 1679581782
transform 1 0 41184 0 1 6804
box -48 -56 720 834
use sg13g2_fill_2  FILLER_9_0
timestamp 1677580104
transform 1 0 1152 0 -1 8316
box -48 -56 240 834
use sg13g2_fill_2  FILLER_9_46
timestamp 1677580104
transform 1 0 5568 0 -1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_9_48
timestamp 1677579658
transform 1 0 5760 0 -1 8316
box -48 -56 144 834
use sg13g2_fill_2  FILLER_9_66
timestamp 1677580104
transform 1 0 7488 0 -1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_9_68
timestamp 1677579658
transform 1 0 7680 0 -1 8316
box -48 -56 144 834
use sg13g2_fill_1  FILLER_9_79
timestamp 1677579658
transform 1 0 8736 0 -1 8316
box -48 -56 144 834
use sg13g2_decap_8  FILLER_9_148
timestamp 1679581782
transform 1 0 15360 0 -1 8316
box -48 -56 720 834
use sg13g2_fill_1  FILLER_9_172
timestamp 1677579658
transform 1 0 17664 0 -1 8316
box -48 -56 144 834
use sg13g2_fill_2  FILLER_9_190
timestamp 1677580104
transform 1 0 19392 0 -1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_9_192
timestamp 1677579658
transform 1 0 19584 0 -1 8316
box -48 -56 144 834
use sg13g2_decap_4  FILLER_9_214
timestamp 1679577901
transform 1 0 21696 0 -1 8316
box -48 -56 432 834
use sg13g2_fill_2  FILLER_9_218
timestamp 1677580104
transform 1 0 22080 0 -1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_9_224
timestamp 1677579658
transform 1 0 22656 0 -1 8316
box -48 -56 144 834
use sg13g2_decap_8  FILLER_9_242
timestamp 1679581782
transform 1 0 24384 0 -1 8316
box -48 -56 720 834
use sg13g2_fill_1  FILLER_9_249
timestamp 1677579658
transform 1 0 25056 0 -1 8316
box -48 -56 144 834
use sg13g2_decap_8  FILLER_9_275
timestamp 1679581782
transform 1 0 27552 0 -1 8316
box -48 -56 720 834
use sg13g2_fill_2  FILLER_9_282
timestamp 1677580104
transform 1 0 28224 0 -1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_9_284
timestamp 1677579658
transform 1 0 28416 0 -1 8316
box -48 -56 144 834
use sg13g2_fill_1  FILLER_9_331
timestamp 1677579658
transform 1 0 32928 0 -1 8316
box -48 -56 144 834
use sg13g2_decap_4  FILLER_9_336
timestamp 1679577901
transform 1 0 33408 0 -1 8316
box -48 -56 432 834
use sg13g2_fill_2  FILLER_9_340
timestamp 1677580104
transform 1 0 33792 0 -1 8316
box -48 -56 240 834
use sg13g2_decap_8  FILLER_9_386
timestamp 1679581782
transform 1 0 38208 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_393
timestamp 1679581782
transform 1 0 38880 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_400
timestamp 1679581782
transform 1 0 39552 0 -1 8316
box -48 -56 720 834
use sg13g2_fill_2  FILLER_9_407
timestamp 1677580104
transform 1 0 40224 0 -1 8316
box -48 -56 240 834
use sg13g2_fill_2  FILLER_9_421
timestamp 1677580104
transform 1 0 41568 0 -1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_9_423
timestamp 1677579658
transform 1 0 41760 0 -1 8316
box -48 -56 144 834
use sg13g2_decap_4  FILLER_10_0
timestamp 1679577901
transform 1 0 1152 0 1 8316
box -48 -56 432 834
use sg13g2_fill_2  FILLER_10_21
timestamp 1677580104
transform 1 0 3168 0 1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_10_23
timestamp 1677579658
transform 1 0 3360 0 1 8316
box -48 -56 144 834
use sg13g2_fill_2  FILLER_10_34
timestamp 1677580104
transform 1 0 4416 0 1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_10_36
timestamp 1677579658
transform 1 0 4608 0 1 8316
box -48 -56 144 834
use sg13g2_decap_8  FILLER_10_105
timestamp 1679581782
transform 1 0 11232 0 1 8316
box -48 -56 720 834
use sg13g2_decap_4  FILLER_10_112
timestamp 1679577901
transform 1 0 11904 0 1 8316
box -48 -56 432 834
use sg13g2_fill_1  FILLER_10_116
timestamp 1677579658
transform 1 0 12288 0 1 8316
box -48 -56 144 834
use sg13g2_fill_2  FILLER_10_151
timestamp 1677580104
transform 1 0 15648 0 1 8316
box -48 -56 240 834
use sg13g2_fill_2  FILLER_10_191
timestamp 1677580104
transform 1 0 19488 0 1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_10_193
timestamp 1677579658
transform 1 0 19680 0 1 8316
box -48 -56 144 834
use sg13g2_decap_8  FILLER_10_236
timestamp 1679581782
transform 1 0 23808 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_243
timestamp 1679581782
transform 1 0 24480 0 1 8316
box -48 -56 720 834
use sg13g2_fill_1  FILLER_10_250
timestamp 1677579658
transform 1 0 25152 0 1 8316
box -48 -56 144 834
use sg13g2_fill_2  FILLER_10_289
timestamp 1677580104
transform 1 0 28896 0 1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_10_291
timestamp 1677579658
transform 1 0 29088 0 1 8316
box -48 -56 144 834
use sg13g2_fill_1  FILLER_10_296
timestamp 1677579658
transform 1 0 29568 0 1 8316
box -48 -56 144 834
use sg13g2_fill_2  FILLER_10_334
timestamp 1677580104
transform 1 0 33216 0 1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_10_336
timestamp 1677579658
transform 1 0 33408 0 1 8316
box -48 -56 144 834
use sg13g2_decap_4  FILLER_10_397
timestamp 1679577901
transform 1 0 39264 0 1 8316
box -48 -56 432 834
use sg13g2_fill_1  FILLER_10_401
timestamp 1677579658
transform 1 0 39648 0 1 8316
box -48 -56 144 834
use sg13g2_fill_2  FILLER_10_410
timestamp 1677580104
transform 1 0 40512 0 1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_10_412
timestamp 1677579658
transform 1 0 40704 0 1 8316
box -48 -56 144 834
use sg13g2_fill_2  FILLER_10_421
timestamp 1677580104
transform 1 0 41568 0 1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_10_423
timestamp 1677579658
transform 1 0 41760 0 1 8316
box -48 -56 144 834
use sg13g2_fill_2  FILLER_11_0
timestamp 1677580104
transform 1 0 1152 0 -1 9828
box -48 -56 240 834
use sg13g2_fill_1  FILLER_11_2
timestamp 1677579658
transform 1 0 1344 0 -1 9828
box -48 -56 144 834
use sg13g2_fill_2  FILLER_11_20
timestamp 1677580104
transform 1 0 3072 0 -1 9828
box -48 -56 240 834
use sg13g2_decap_8  FILLER_11_37
timestamp 1679581782
transform 1 0 4704 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_44
timestamp 1679581782
transform 1 0 5376 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_51
timestamp 1679581782
transform 1 0 6048 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_58
timestamp 1679581782
transform 1 0 6720 0 -1 9828
box -48 -56 720 834
use sg13g2_fill_2  FILLER_11_65
timestamp 1677580104
transform 1 0 7392 0 -1 9828
box -48 -56 240 834
use sg13g2_fill_1  FILLER_11_67
timestamp 1677579658
transform 1 0 7584 0 -1 9828
box -48 -56 144 834
use sg13g2_decap_8  FILLER_11_85
timestamp 1679581782
transform 1 0 9312 0 -1 9828
box -48 -56 720 834
use sg13g2_fill_2  FILLER_11_92
timestamp 1677580104
transform 1 0 9984 0 -1 9828
box -48 -56 240 834
use sg13g2_decap_8  FILLER_11_128
timestamp 1679581782
transform 1 0 13440 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_135
timestamp 1679581782
transform 1 0 14112 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_4  FILLER_11_142
timestamp 1679577901
transform 1 0 14784 0 -1 9828
box -48 -56 432 834
use sg13g2_decap_8  FILLER_11_163
timestamp 1679581782
transform 1 0 16800 0 -1 9828
box -48 -56 720 834
use sg13g2_fill_2  FILLER_11_170
timestamp 1677580104
transform 1 0 17472 0 -1 9828
box -48 -56 240 834
use sg13g2_fill_1  FILLER_11_172
timestamp 1677579658
transform 1 0 17664 0 -1 9828
box -48 -56 144 834
use sg13g2_decap_8  FILLER_11_194
timestamp 1679581782
transform 1 0 19776 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_201
timestamp 1679581782
transform 1 0 20448 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_212
timestamp 1679581782
transform 1 0 21504 0 -1 9828
box -48 -56 720 834
use sg13g2_fill_2  FILLER_11_219
timestamp 1677580104
transform 1 0 22176 0 -1 9828
box -48 -56 240 834
use sg13g2_fill_2  FILLER_11_238
timestamp 1677580104
transform 1 0 24000 0 -1 9828
box -48 -56 240 834
use sg13g2_decap_8  FILLER_11_257
timestamp 1679581782
transform 1 0 25824 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_264
timestamp 1679581782
transform 1 0 26496 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_4  FILLER_11_271
timestamp 1679577901
transform 1 0 27168 0 -1 9828
box -48 -56 432 834
use sg13g2_fill_1  FILLER_11_275
timestamp 1677579658
transform 1 0 27552 0 -1 9828
box -48 -56 144 834
use sg13g2_fill_2  FILLER_11_293
timestamp 1677580104
transform 1 0 29280 0 -1 9828
box -48 -56 240 834
use sg13g2_decap_8  FILLER_11_384
timestamp 1679581782
transform 1 0 38016 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_391
timestamp 1679581782
transform 1 0 38688 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_398
timestamp 1679581782
transform 1 0 39360 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_4  FILLER_11_405
timestamp 1679577901
transform 1 0 40032 0 -1 9828
box -48 -56 432 834
use sg13g2_fill_2  FILLER_11_421
timestamp 1677580104
transform 1 0 41568 0 -1 9828
box -48 -56 240 834
use sg13g2_fill_1  FILLER_11_423
timestamp 1677579658
transform 1 0 41760 0 -1 9828
box -48 -56 144 834
<< labels >>
flabel metal2 s 2936 10672 3016 10752 0 FreeSans 320 0 0 0 A_I_top
port 0 nsew signal output
flabel metal2 s 1784 10672 1864 10752 0 FreeSans 320 0 0 0 A_O_top
port 1 nsew signal input
flabel metal2 s 4088 10672 4168 10752 0 FreeSans 320 0 0 0 A_T_top
port 2 nsew signal output
flabel metal2 s 8696 10672 8776 10752 0 FreeSans 320 0 0 0 A_config_C_bit0
port 3 nsew signal output
flabel metal2 s 9848 10672 9928 10752 0 FreeSans 320 0 0 0 A_config_C_bit1
port 4 nsew signal output
flabel metal2 s 11000 10672 11080 10752 0 FreeSans 320 0 0 0 A_config_C_bit2
port 5 nsew signal output
flabel metal2 s 12152 10672 12232 10752 0 FreeSans 320 0 0 0 A_config_C_bit3
port 6 nsew signal output
flabel metal2 s 6392 10672 6472 10752 0 FreeSans 320 0 0 0 B_I_top
port 7 nsew signal output
flabel metal2 s 5240 10672 5320 10752 0 FreeSans 320 0 0 0 B_O_top
port 8 nsew signal input
flabel metal2 s 7544 10672 7624 10752 0 FreeSans 320 0 0 0 B_T_top
port 9 nsew signal output
flabel metal2 s 13304 10672 13384 10752 0 FreeSans 320 0 0 0 B_config_C_bit0
port 10 nsew signal output
flabel metal2 s 14456 10672 14536 10752 0 FreeSans 320 0 0 0 B_config_C_bit1
port 11 nsew signal output
flabel metal2 s 15608 10672 15688 10752 0 FreeSans 320 0 0 0 B_config_C_bit2
port 12 nsew signal output
flabel metal2 s 16760 10672 16840 10752 0 FreeSans 320 0 0 0 B_config_C_bit3
port 13 nsew signal output
flabel metal2 s 19448 0 19528 80 0 FreeSans 320 0 0 0 Ci
port 14 nsew signal input
flabel metal3 s 0 44 80 124 0 FreeSans 320 0 0 0 FrameData[0]
port 15 nsew signal input
flabel metal3 s 0 3404 80 3484 0 FreeSans 320 0 0 0 FrameData[10]
port 16 nsew signal input
flabel metal3 s 0 3740 80 3820 0 FreeSans 320 0 0 0 FrameData[11]
port 17 nsew signal input
flabel metal3 s 0 4076 80 4156 0 FreeSans 320 0 0 0 FrameData[12]
port 18 nsew signal input
flabel metal3 s 0 4412 80 4492 0 FreeSans 320 0 0 0 FrameData[13]
port 19 nsew signal input
flabel metal3 s 0 4748 80 4828 0 FreeSans 320 0 0 0 FrameData[14]
port 20 nsew signal input
flabel metal3 s 0 5084 80 5164 0 FreeSans 320 0 0 0 FrameData[15]
port 21 nsew signal input
flabel metal3 s 0 5420 80 5500 0 FreeSans 320 0 0 0 FrameData[16]
port 22 nsew signal input
flabel metal3 s 0 5756 80 5836 0 FreeSans 320 0 0 0 FrameData[17]
port 23 nsew signal input
flabel metal3 s 0 6092 80 6172 0 FreeSans 320 0 0 0 FrameData[18]
port 24 nsew signal input
flabel metal3 s 0 6428 80 6508 0 FreeSans 320 0 0 0 FrameData[19]
port 25 nsew signal input
flabel metal3 s 0 380 80 460 0 FreeSans 320 0 0 0 FrameData[1]
port 26 nsew signal input
flabel metal3 s 0 6764 80 6844 0 FreeSans 320 0 0 0 FrameData[20]
port 27 nsew signal input
flabel metal3 s 0 7100 80 7180 0 FreeSans 320 0 0 0 FrameData[21]
port 28 nsew signal input
flabel metal3 s 0 7436 80 7516 0 FreeSans 320 0 0 0 FrameData[22]
port 29 nsew signal input
flabel metal3 s 0 7772 80 7852 0 FreeSans 320 0 0 0 FrameData[23]
port 30 nsew signal input
flabel metal3 s 0 8108 80 8188 0 FreeSans 320 0 0 0 FrameData[24]
port 31 nsew signal input
flabel metal3 s 0 8444 80 8524 0 FreeSans 320 0 0 0 FrameData[25]
port 32 nsew signal input
flabel metal3 s 0 8780 80 8860 0 FreeSans 320 0 0 0 FrameData[26]
port 33 nsew signal input
flabel metal3 s 0 9116 80 9196 0 FreeSans 320 0 0 0 FrameData[27]
port 34 nsew signal input
flabel metal3 s 0 9452 80 9532 0 FreeSans 320 0 0 0 FrameData[28]
port 35 nsew signal input
flabel metal3 s 0 9788 80 9868 0 FreeSans 320 0 0 0 FrameData[29]
port 36 nsew signal input
flabel metal3 s 0 716 80 796 0 FreeSans 320 0 0 0 FrameData[2]
port 37 nsew signal input
flabel metal3 s 0 10124 80 10204 0 FreeSans 320 0 0 0 FrameData[30]
port 38 nsew signal input
flabel metal3 s 0 10460 80 10540 0 FreeSans 320 0 0 0 FrameData[31]
port 39 nsew signal input
flabel metal3 s 0 1052 80 1132 0 FreeSans 320 0 0 0 FrameData[3]
port 40 nsew signal input
flabel metal3 s 0 1388 80 1468 0 FreeSans 320 0 0 0 FrameData[4]
port 41 nsew signal input
flabel metal3 s 0 1724 80 1804 0 FreeSans 320 0 0 0 FrameData[5]
port 42 nsew signal input
flabel metal3 s 0 2060 80 2140 0 FreeSans 320 0 0 0 FrameData[6]
port 43 nsew signal input
flabel metal3 s 0 2396 80 2476 0 FreeSans 320 0 0 0 FrameData[7]
port 44 nsew signal input
flabel metal3 s 0 2732 80 2812 0 FreeSans 320 0 0 0 FrameData[8]
port 45 nsew signal input
flabel metal3 s 0 3068 80 3148 0 FreeSans 320 0 0 0 FrameData[9]
port 46 nsew signal input
flabel metal3 s 42928 44 43008 124 0 FreeSans 320 0 0 0 FrameData_O[0]
port 47 nsew signal output
flabel metal3 s 42928 3404 43008 3484 0 FreeSans 320 0 0 0 FrameData_O[10]
port 48 nsew signal output
flabel metal3 s 42928 3740 43008 3820 0 FreeSans 320 0 0 0 FrameData_O[11]
port 49 nsew signal output
flabel metal3 s 42928 4076 43008 4156 0 FreeSans 320 0 0 0 FrameData_O[12]
port 50 nsew signal output
flabel metal3 s 42928 4412 43008 4492 0 FreeSans 320 0 0 0 FrameData_O[13]
port 51 nsew signal output
flabel metal3 s 42928 4748 43008 4828 0 FreeSans 320 0 0 0 FrameData_O[14]
port 52 nsew signal output
flabel metal3 s 42928 5084 43008 5164 0 FreeSans 320 0 0 0 FrameData_O[15]
port 53 nsew signal output
flabel metal3 s 42928 5420 43008 5500 0 FreeSans 320 0 0 0 FrameData_O[16]
port 54 nsew signal output
flabel metal3 s 42928 5756 43008 5836 0 FreeSans 320 0 0 0 FrameData_O[17]
port 55 nsew signal output
flabel metal3 s 42928 6092 43008 6172 0 FreeSans 320 0 0 0 FrameData_O[18]
port 56 nsew signal output
flabel metal3 s 42928 6428 43008 6508 0 FreeSans 320 0 0 0 FrameData_O[19]
port 57 nsew signal output
flabel metal3 s 42928 380 43008 460 0 FreeSans 320 0 0 0 FrameData_O[1]
port 58 nsew signal output
flabel metal3 s 42928 6764 43008 6844 0 FreeSans 320 0 0 0 FrameData_O[20]
port 59 nsew signal output
flabel metal3 s 42928 7100 43008 7180 0 FreeSans 320 0 0 0 FrameData_O[21]
port 60 nsew signal output
flabel metal3 s 42928 7436 43008 7516 0 FreeSans 320 0 0 0 FrameData_O[22]
port 61 nsew signal output
flabel metal3 s 42928 7772 43008 7852 0 FreeSans 320 0 0 0 FrameData_O[23]
port 62 nsew signal output
flabel metal3 s 42928 8108 43008 8188 0 FreeSans 320 0 0 0 FrameData_O[24]
port 63 nsew signal output
flabel metal3 s 42928 8444 43008 8524 0 FreeSans 320 0 0 0 FrameData_O[25]
port 64 nsew signal output
flabel metal3 s 42928 8780 43008 8860 0 FreeSans 320 0 0 0 FrameData_O[26]
port 65 nsew signal output
flabel metal3 s 42928 9116 43008 9196 0 FreeSans 320 0 0 0 FrameData_O[27]
port 66 nsew signal output
flabel metal3 s 42928 9452 43008 9532 0 FreeSans 320 0 0 0 FrameData_O[28]
port 67 nsew signal output
flabel metal3 s 42928 9788 43008 9868 0 FreeSans 320 0 0 0 FrameData_O[29]
port 68 nsew signal output
flabel metal3 s 42928 716 43008 796 0 FreeSans 320 0 0 0 FrameData_O[2]
port 69 nsew signal output
flabel metal3 s 42928 10124 43008 10204 0 FreeSans 320 0 0 0 FrameData_O[30]
port 70 nsew signal output
flabel metal3 s 42928 10460 43008 10540 0 FreeSans 320 0 0 0 FrameData_O[31]
port 71 nsew signal output
flabel metal3 s 42928 1052 43008 1132 0 FreeSans 320 0 0 0 FrameData_O[3]
port 72 nsew signal output
flabel metal3 s 42928 1388 43008 1468 0 FreeSans 320 0 0 0 FrameData_O[4]
port 73 nsew signal output
flabel metal3 s 42928 1724 43008 1804 0 FreeSans 320 0 0 0 FrameData_O[5]
port 74 nsew signal output
flabel metal3 s 42928 2060 43008 2140 0 FreeSans 320 0 0 0 FrameData_O[6]
port 75 nsew signal output
flabel metal3 s 42928 2396 43008 2476 0 FreeSans 320 0 0 0 FrameData_O[7]
port 76 nsew signal output
flabel metal3 s 42928 2732 43008 2812 0 FreeSans 320 0 0 0 FrameData_O[8]
port 77 nsew signal output
flabel metal3 s 42928 3068 43008 3148 0 FreeSans 320 0 0 0 FrameData_O[9]
port 78 nsew signal output
flabel metal2 s 29816 0 29896 80 0 FreeSans 320 0 0 0 FrameStrobe[0]
port 79 nsew signal input
flabel metal2 s 31736 0 31816 80 0 FreeSans 320 0 0 0 FrameStrobe[10]
port 80 nsew signal input
flabel metal2 s 31928 0 32008 80 0 FreeSans 320 0 0 0 FrameStrobe[11]
port 81 nsew signal input
flabel metal2 s 32120 0 32200 80 0 FreeSans 320 0 0 0 FrameStrobe[12]
port 82 nsew signal input
flabel metal2 s 32312 0 32392 80 0 FreeSans 320 0 0 0 FrameStrobe[13]
port 83 nsew signal input
flabel metal2 s 32504 0 32584 80 0 FreeSans 320 0 0 0 FrameStrobe[14]
port 84 nsew signal input
flabel metal2 s 32696 0 32776 80 0 FreeSans 320 0 0 0 FrameStrobe[15]
port 85 nsew signal input
flabel metal2 s 32888 0 32968 80 0 FreeSans 320 0 0 0 FrameStrobe[16]
port 86 nsew signal input
flabel metal2 s 33080 0 33160 80 0 FreeSans 320 0 0 0 FrameStrobe[17]
port 87 nsew signal input
flabel metal2 s 33272 0 33352 80 0 FreeSans 320 0 0 0 FrameStrobe[18]
port 88 nsew signal input
flabel metal2 s 33464 0 33544 80 0 FreeSans 320 0 0 0 FrameStrobe[19]
port 89 nsew signal input
flabel metal2 s 30008 0 30088 80 0 FreeSans 320 0 0 0 FrameStrobe[1]
port 90 nsew signal input
flabel metal2 s 30200 0 30280 80 0 FreeSans 320 0 0 0 FrameStrobe[2]
port 91 nsew signal input
flabel metal2 s 30392 0 30472 80 0 FreeSans 320 0 0 0 FrameStrobe[3]
port 92 nsew signal input
flabel metal2 s 30584 0 30664 80 0 FreeSans 320 0 0 0 FrameStrobe[4]
port 93 nsew signal input
flabel metal2 s 30776 0 30856 80 0 FreeSans 320 0 0 0 FrameStrobe[5]
port 94 nsew signal input
flabel metal2 s 30968 0 31048 80 0 FreeSans 320 0 0 0 FrameStrobe[6]
port 95 nsew signal input
flabel metal2 s 31160 0 31240 80 0 FreeSans 320 0 0 0 FrameStrobe[7]
port 96 nsew signal input
flabel metal2 s 31352 0 31432 80 0 FreeSans 320 0 0 0 FrameStrobe[8]
port 97 nsew signal input
flabel metal2 s 31544 0 31624 80 0 FreeSans 320 0 0 0 FrameStrobe[9]
port 98 nsew signal input
flabel metal2 s 19064 10672 19144 10752 0 FreeSans 320 0 0 0 FrameStrobe_O[0]
port 99 nsew signal output
flabel metal2 s 30584 10672 30664 10752 0 FreeSans 320 0 0 0 FrameStrobe_O[10]
port 100 nsew signal output
flabel metal2 s 31736 10672 31816 10752 0 FreeSans 320 0 0 0 FrameStrobe_O[11]
port 101 nsew signal output
flabel metal2 s 32888 10672 32968 10752 0 FreeSans 320 0 0 0 FrameStrobe_O[12]
port 102 nsew signal output
flabel metal2 s 34040 10672 34120 10752 0 FreeSans 320 0 0 0 FrameStrobe_O[13]
port 103 nsew signal output
flabel metal2 s 35192 10672 35272 10752 0 FreeSans 320 0 0 0 FrameStrobe_O[14]
port 104 nsew signal output
flabel metal2 s 36344 10672 36424 10752 0 FreeSans 320 0 0 0 FrameStrobe_O[15]
port 105 nsew signal output
flabel metal2 s 37496 10672 37576 10752 0 FreeSans 320 0 0 0 FrameStrobe_O[16]
port 106 nsew signal output
flabel metal2 s 38648 10672 38728 10752 0 FreeSans 320 0 0 0 FrameStrobe_O[17]
port 107 nsew signal output
flabel metal2 s 39800 10672 39880 10752 0 FreeSans 320 0 0 0 FrameStrobe_O[18]
port 108 nsew signal output
flabel metal2 s 40952 10672 41032 10752 0 FreeSans 320 0 0 0 FrameStrobe_O[19]
port 109 nsew signal output
flabel metal2 s 20216 10672 20296 10752 0 FreeSans 320 0 0 0 FrameStrobe_O[1]
port 110 nsew signal output
flabel metal2 s 21368 10672 21448 10752 0 FreeSans 320 0 0 0 FrameStrobe_O[2]
port 111 nsew signal output
flabel metal2 s 22520 10672 22600 10752 0 FreeSans 320 0 0 0 FrameStrobe_O[3]
port 112 nsew signal output
flabel metal2 s 23672 10672 23752 10752 0 FreeSans 320 0 0 0 FrameStrobe_O[4]
port 113 nsew signal output
flabel metal2 s 24824 10672 24904 10752 0 FreeSans 320 0 0 0 FrameStrobe_O[5]
port 114 nsew signal output
flabel metal2 s 25976 10672 26056 10752 0 FreeSans 320 0 0 0 FrameStrobe_O[6]
port 115 nsew signal output
flabel metal2 s 27128 10672 27208 10752 0 FreeSans 320 0 0 0 FrameStrobe_O[7]
port 116 nsew signal output
flabel metal2 s 28280 10672 28360 10752 0 FreeSans 320 0 0 0 FrameStrobe_O[8]
port 117 nsew signal output
flabel metal2 s 29432 10672 29512 10752 0 FreeSans 320 0 0 0 FrameStrobe_O[9]
port 118 nsew signal output
flabel metal2 s 9464 0 9544 80 0 FreeSans 320 0 0 0 N1END[0]
port 119 nsew signal input
flabel metal2 s 9656 0 9736 80 0 FreeSans 320 0 0 0 N1END[1]
port 120 nsew signal input
flabel metal2 s 9848 0 9928 80 0 FreeSans 320 0 0 0 N1END[2]
port 121 nsew signal input
flabel metal2 s 10040 0 10120 80 0 FreeSans 320 0 0 0 N1END[3]
port 122 nsew signal input
flabel metal2 s 11768 0 11848 80 0 FreeSans 320 0 0 0 N2END[0]
port 123 nsew signal input
flabel metal2 s 11960 0 12040 80 0 FreeSans 320 0 0 0 N2END[1]
port 124 nsew signal input
flabel metal2 s 12152 0 12232 80 0 FreeSans 320 0 0 0 N2END[2]
port 125 nsew signal input
flabel metal2 s 12344 0 12424 80 0 FreeSans 320 0 0 0 N2END[3]
port 126 nsew signal input
flabel metal2 s 12536 0 12616 80 0 FreeSans 320 0 0 0 N2END[4]
port 127 nsew signal input
flabel metal2 s 12728 0 12808 80 0 FreeSans 320 0 0 0 N2END[5]
port 128 nsew signal input
flabel metal2 s 12920 0 13000 80 0 FreeSans 320 0 0 0 N2END[6]
port 129 nsew signal input
flabel metal2 s 13112 0 13192 80 0 FreeSans 320 0 0 0 N2END[7]
port 130 nsew signal input
flabel metal2 s 10232 0 10312 80 0 FreeSans 320 0 0 0 N2MID[0]
port 131 nsew signal input
flabel metal2 s 10424 0 10504 80 0 FreeSans 320 0 0 0 N2MID[1]
port 132 nsew signal input
flabel metal2 s 10616 0 10696 80 0 FreeSans 320 0 0 0 N2MID[2]
port 133 nsew signal input
flabel metal2 s 10808 0 10888 80 0 FreeSans 320 0 0 0 N2MID[3]
port 134 nsew signal input
flabel metal2 s 11000 0 11080 80 0 FreeSans 320 0 0 0 N2MID[4]
port 135 nsew signal input
flabel metal2 s 11192 0 11272 80 0 FreeSans 320 0 0 0 N2MID[5]
port 136 nsew signal input
flabel metal2 s 11384 0 11464 80 0 FreeSans 320 0 0 0 N2MID[6]
port 137 nsew signal input
flabel metal2 s 11576 0 11656 80 0 FreeSans 320 0 0 0 N2MID[7]
port 138 nsew signal input
flabel metal2 s 13304 0 13384 80 0 FreeSans 320 0 0 0 N4END[0]
port 139 nsew signal input
flabel metal2 s 15224 0 15304 80 0 FreeSans 320 0 0 0 N4END[10]
port 140 nsew signal input
flabel metal2 s 15416 0 15496 80 0 FreeSans 320 0 0 0 N4END[11]
port 141 nsew signal input
flabel metal2 s 15608 0 15688 80 0 FreeSans 320 0 0 0 N4END[12]
port 142 nsew signal input
flabel metal2 s 15800 0 15880 80 0 FreeSans 320 0 0 0 N4END[13]
port 143 nsew signal input
flabel metal2 s 15992 0 16072 80 0 FreeSans 320 0 0 0 N4END[14]
port 144 nsew signal input
flabel metal2 s 16184 0 16264 80 0 FreeSans 320 0 0 0 N4END[15]
port 145 nsew signal input
flabel metal2 s 13496 0 13576 80 0 FreeSans 320 0 0 0 N4END[1]
port 146 nsew signal input
flabel metal2 s 13688 0 13768 80 0 FreeSans 320 0 0 0 N4END[2]
port 147 nsew signal input
flabel metal2 s 13880 0 13960 80 0 FreeSans 320 0 0 0 N4END[3]
port 148 nsew signal input
flabel metal2 s 14072 0 14152 80 0 FreeSans 320 0 0 0 N4END[4]
port 149 nsew signal input
flabel metal2 s 14264 0 14344 80 0 FreeSans 320 0 0 0 N4END[5]
port 150 nsew signal input
flabel metal2 s 14456 0 14536 80 0 FreeSans 320 0 0 0 N4END[6]
port 151 nsew signal input
flabel metal2 s 14648 0 14728 80 0 FreeSans 320 0 0 0 N4END[7]
port 152 nsew signal input
flabel metal2 s 14840 0 14920 80 0 FreeSans 320 0 0 0 N4END[8]
port 153 nsew signal input
flabel metal2 s 15032 0 15112 80 0 FreeSans 320 0 0 0 N4END[9]
port 154 nsew signal input
flabel metal2 s 16376 0 16456 80 0 FreeSans 320 0 0 0 NN4END[0]
port 155 nsew signal input
flabel metal2 s 18296 0 18376 80 0 FreeSans 320 0 0 0 NN4END[10]
port 156 nsew signal input
flabel metal2 s 18488 0 18568 80 0 FreeSans 320 0 0 0 NN4END[11]
port 157 nsew signal input
flabel metal2 s 18680 0 18760 80 0 FreeSans 320 0 0 0 NN4END[12]
port 158 nsew signal input
flabel metal2 s 18872 0 18952 80 0 FreeSans 320 0 0 0 NN4END[13]
port 159 nsew signal input
flabel metal2 s 19064 0 19144 80 0 FreeSans 320 0 0 0 NN4END[14]
port 160 nsew signal input
flabel metal2 s 19256 0 19336 80 0 FreeSans 320 0 0 0 NN4END[15]
port 161 nsew signal input
flabel metal2 s 16568 0 16648 80 0 FreeSans 320 0 0 0 NN4END[1]
port 162 nsew signal input
flabel metal2 s 16760 0 16840 80 0 FreeSans 320 0 0 0 NN4END[2]
port 163 nsew signal input
flabel metal2 s 16952 0 17032 80 0 FreeSans 320 0 0 0 NN4END[3]
port 164 nsew signal input
flabel metal2 s 17144 0 17224 80 0 FreeSans 320 0 0 0 NN4END[4]
port 165 nsew signal input
flabel metal2 s 17336 0 17416 80 0 FreeSans 320 0 0 0 NN4END[5]
port 166 nsew signal input
flabel metal2 s 17528 0 17608 80 0 FreeSans 320 0 0 0 NN4END[6]
port 167 nsew signal input
flabel metal2 s 17720 0 17800 80 0 FreeSans 320 0 0 0 NN4END[7]
port 168 nsew signal input
flabel metal2 s 17912 0 17992 80 0 FreeSans 320 0 0 0 NN4END[8]
port 169 nsew signal input
flabel metal2 s 18104 0 18184 80 0 FreeSans 320 0 0 0 NN4END[9]
port 170 nsew signal input
flabel metal2 s 19640 0 19720 80 0 FreeSans 320 0 0 0 S1BEG[0]
port 171 nsew signal output
flabel metal2 s 19832 0 19912 80 0 FreeSans 320 0 0 0 S1BEG[1]
port 172 nsew signal output
flabel metal2 s 20024 0 20104 80 0 FreeSans 320 0 0 0 S1BEG[2]
port 173 nsew signal output
flabel metal2 s 20216 0 20296 80 0 FreeSans 320 0 0 0 S1BEG[3]
port 174 nsew signal output
flabel metal2 s 20408 0 20488 80 0 FreeSans 320 0 0 0 S2BEG[0]
port 175 nsew signal output
flabel metal2 s 20600 0 20680 80 0 FreeSans 320 0 0 0 S2BEG[1]
port 176 nsew signal output
flabel metal2 s 20792 0 20872 80 0 FreeSans 320 0 0 0 S2BEG[2]
port 177 nsew signal output
flabel metal2 s 20984 0 21064 80 0 FreeSans 320 0 0 0 S2BEG[3]
port 178 nsew signal output
flabel metal2 s 21176 0 21256 80 0 FreeSans 320 0 0 0 S2BEG[4]
port 179 nsew signal output
flabel metal2 s 21368 0 21448 80 0 FreeSans 320 0 0 0 S2BEG[5]
port 180 nsew signal output
flabel metal2 s 21560 0 21640 80 0 FreeSans 320 0 0 0 S2BEG[6]
port 181 nsew signal output
flabel metal2 s 21752 0 21832 80 0 FreeSans 320 0 0 0 S2BEG[7]
port 182 nsew signal output
flabel metal2 s 21944 0 22024 80 0 FreeSans 320 0 0 0 S2BEGb[0]
port 183 nsew signal output
flabel metal2 s 22136 0 22216 80 0 FreeSans 320 0 0 0 S2BEGb[1]
port 184 nsew signal output
flabel metal2 s 22328 0 22408 80 0 FreeSans 320 0 0 0 S2BEGb[2]
port 185 nsew signal output
flabel metal2 s 22520 0 22600 80 0 FreeSans 320 0 0 0 S2BEGb[3]
port 186 nsew signal output
flabel metal2 s 22712 0 22792 80 0 FreeSans 320 0 0 0 S2BEGb[4]
port 187 nsew signal output
flabel metal2 s 22904 0 22984 80 0 FreeSans 320 0 0 0 S2BEGb[5]
port 188 nsew signal output
flabel metal2 s 23096 0 23176 80 0 FreeSans 320 0 0 0 S2BEGb[6]
port 189 nsew signal output
flabel metal2 s 23288 0 23368 80 0 FreeSans 320 0 0 0 S2BEGb[7]
port 190 nsew signal output
flabel metal2 s 23480 0 23560 80 0 FreeSans 320 0 0 0 S4BEG[0]
port 191 nsew signal output
flabel metal2 s 25400 0 25480 80 0 FreeSans 320 0 0 0 S4BEG[10]
port 192 nsew signal output
flabel metal2 s 25592 0 25672 80 0 FreeSans 320 0 0 0 S4BEG[11]
port 193 nsew signal output
flabel metal2 s 25784 0 25864 80 0 FreeSans 320 0 0 0 S4BEG[12]
port 194 nsew signal output
flabel metal2 s 25976 0 26056 80 0 FreeSans 320 0 0 0 S4BEG[13]
port 195 nsew signal output
flabel metal2 s 26168 0 26248 80 0 FreeSans 320 0 0 0 S4BEG[14]
port 196 nsew signal output
flabel metal2 s 26360 0 26440 80 0 FreeSans 320 0 0 0 S4BEG[15]
port 197 nsew signal output
flabel metal2 s 23672 0 23752 80 0 FreeSans 320 0 0 0 S4BEG[1]
port 198 nsew signal output
flabel metal2 s 23864 0 23944 80 0 FreeSans 320 0 0 0 S4BEG[2]
port 199 nsew signal output
flabel metal2 s 24056 0 24136 80 0 FreeSans 320 0 0 0 S4BEG[3]
port 200 nsew signal output
flabel metal2 s 24248 0 24328 80 0 FreeSans 320 0 0 0 S4BEG[4]
port 201 nsew signal output
flabel metal2 s 24440 0 24520 80 0 FreeSans 320 0 0 0 S4BEG[5]
port 202 nsew signal output
flabel metal2 s 24632 0 24712 80 0 FreeSans 320 0 0 0 S4BEG[6]
port 203 nsew signal output
flabel metal2 s 24824 0 24904 80 0 FreeSans 320 0 0 0 S4BEG[7]
port 204 nsew signal output
flabel metal2 s 25016 0 25096 80 0 FreeSans 320 0 0 0 S4BEG[8]
port 205 nsew signal output
flabel metal2 s 25208 0 25288 80 0 FreeSans 320 0 0 0 S4BEG[9]
port 206 nsew signal output
flabel metal2 s 26552 0 26632 80 0 FreeSans 320 0 0 0 SS4BEG[0]
port 207 nsew signal output
flabel metal2 s 28472 0 28552 80 0 FreeSans 320 0 0 0 SS4BEG[10]
port 208 nsew signal output
flabel metal2 s 28664 0 28744 80 0 FreeSans 320 0 0 0 SS4BEG[11]
port 209 nsew signal output
flabel metal2 s 28856 0 28936 80 0 FreeSans 320 0 0 0 SS4BEG[12]
port 210 nsew signal output
flabel metal2 s 29048 0 29128 80 0 FreeSans 320 0 0 0 SS4BEG[13]
port 211 nsew signal output
flabel metal2 s 29240 0 29320 80 0 FreeSans 320 0 0 0 SS4BEG[14]
port 212 nsew signal output
flabel metal2 s 29432 0 29512 80 0 FreeSans 320 0 0 0 SS4BEG[15]
port 213 nsew signal output
flabel metal2 s 26744 0 26824 80 0 FreeSans 320 0 0 0 SS4BEG[1]
port 214 nsew signal output
flabel metal2 s 26936 0 27016 80 0 FreeSans 320 0 0 0 SS4BEG[2]
port 215 nsew signal output
flabel metal2 s 27128 0 27208 80 0 FreeSans 320 0 0 0 SS4BEG[3]
port 216 nsew signal output
flabel metal2 s 27320 0 27400 80 0 FreeSans 320 0 0 0 SS4BEG[4]
port 217 nsew signal output
flabel metal2 s 27512 0 27592 80 0 FreeSans 320 0 0 0 SS4BEG[5]
port 218 nsew signal output
flabel metal2 s 27704 0 27784 80 0 FreeSans 320 0 0 0 SS4BEG[6]
port 219 nsew signal output
flabel metal2 s 27896 0 27976 80 0 FreeSans 320 0 0 0 SS4BEG[7]
port 220 nsew signal output
flabel metal2 s 28088 0 28168 80 0 FreeSans 320 0 0 0 SS4BEG[8]
port 221 nsew signal output
flabel metal2 s 28280 0 28360 80 0 FreeSans 320 0 0 0 SS4BEG[9]
port 222 nsew signal output
flabel metal2 s 29624 0 29704 80 0 FreeSans 320 0 0 0 UserCLK
port 223 nsew signal input
flabel metal2 s 17912 10672 17992 10752 0 FreeSans 320 0 0 0 UserCLKo
port 224 nsew signal output
flabel metal6 s 4892 0 5332 10752 0 FreeSans 2624 90 0 0 VGND
port 225 nsew ground bidirectional
flabel metal6 s 4892 0 5332 328 0 FreeSans 2624 0 0 0 VGND
port 225 nsew ground bidirectional
flabel metal6 s 4892 10424 5332 10752 0 FreeSans 2624 0 0 0 VGND
port 225 nsew ground bidirectional
flabel metal6 s 20012 0 20452 10752 0 FreeSans 2624 90 0 0 VGND
port 225 nsew ground bidirectional
flabel metal6 s 20012 0 20452 328 0 FreeSans 2624 0 0 0 VGND
port 225 nsew ground bidirectional
flabel metal6 s 20012 10424 20452 10752 0 FreeSans 2624 0 0 0 VGND
port 225 nsew ground bidirectional
flabel metal6 s 35132 0 35572 10752 0 FreeSans 2624 90 0 0 VGND
port 225 nsew ground bidirectional
flabel metal6 s 35132 0 35572 328 0 FreeSans 2624 0 0 0 VGND
port 225 nsew ground bidirectional
flabel metal6 s 35132 10424 35572 10752 0 FreeSans 2624 0 0 0 VGND
port 225 nsew ground bidirectional
flabel metal6 s 3652 0 4092 10752 0 FreeSans 2624 90 0 0 VPWR
port 226 nsew power bidirectional
flabel metal6 s 3652 0 4092 328 0 FreeSans 2624 0 0 0 VPWR
port 226 nsew power bidirectional
flabel metal6 s 3652 10424 4092 10752 0 FreeSans 2624 0 0 0 VPWR
port 226 nsew power bidirectional
flabel metal6 s 18772 0 19212 10752 0 FreeSans 2624 90 0 0 VPWR
port 226 nsew power bidirectional
flabel metal6 s 18772 0 19212 328 0 FreeSans 2624 0 0 0 VPWR
port 226 nsew power bidirectional
flabel metal6 s 18772 10424 19212 10752 0 FreeSans 2624 0 0 0 VPWR
port 226 nsew power bidirectional
flabel metal6 s 33892 0 34332 10752 0 FreeSans 2624 90 0 0 VPWR
port 226 nsew power bidirectional
flabel metal6 s 33892 0 34332 328 0 FreeSans 2624 0 0 0 VPWR
port 226 nsew power bidirectional
flabel metal6 s 33892 10424 34332 10752 0 FreeSans 2624 0 0 0 VPWR
port 226 nsew power bidirectional
rlabel metal1 21504 9828 21504 9828 0 VGND
rlabel metal1 21504 9072 21504 9072 0 VPWR
rlabel metal2 3648 5460 3648 5460 0 A_I_top
rlabel metal2 1824 10638 1824 10638 0 A_O_top
rlabel metal2 4608 10186 4608 10186 0 A_T_top
rlabel metal2 9216 10186 9216 10186 0 A_config_C_bit0
rlabel metal2 9504 9766 9504 9766 0 A_config_C_bit1
rlabel metal2 10368 9430 10368 9430 0 A_config_C_bit2
rlabel metal3 11952 9660 11952 9660 0 A_config_C_bit3
rlabel metal2 6048 7308 6048 7308 0 B_I_top
rlabel metal2 20064 2562 20064 2562 0 B_O_top
rlabel metal2 9984 7434 9984 7434 0 B_T_top
rlabel metal2 13344 10176 13344 10176 0 B_config_C_bit0
rlabel metal2 13920 9240 13920 9240 0 B_config_C_bit1
rlabel metal2 15600 8820 15600 8820 0 B_config_C_bit2
rlabel metal2 16752 9660 16752 9660 0 B_config_C_bit3
rlabel metal3 15696 1176 15696 1176 0 FrameData[0]
rlabel metal3 654 3444 654 3444 0 FrameData[10]
rlabel metal3 1278 3780 1278 3780 0 FrameData[11]
rlabel metal3 78 4116 78 4116 0 FrameData[12]
rlabel metal3 654 4452 654 4452 0 FrameData[13]
rlabel metal3 1230 4788 1230 4788 0 FrameData[14]
rlabel metal2 2928 1092 2928 1092 0 FrameData[15]
rlabel metal5 18112 2478 18112 2478 0 FrameData[16]
rlabel metal2 1056 4494 1056 4494 0 FrameData[17]
rlabel metal2 1632 4116 1632 4116 0 FrameData[18]
rlabel metal2 1584 4956 1584 4956 0 FrameData[19]
rlabel metal2 1344 1008 1344 1008 0 FrameData[1]
rlabel metal2 1536 2814 1536 2814 0 FrameData[20]
rlabel metal3 1776 3444 1776 3444 0 FrameData[21]
rlabel metal2 1632 8064 1632 8064 0 FrameData[22]
rlabel metal2 1440 7896 1440 7896 0 FrameData[23]
rlabel metal2 1536 8820 1536 8820 0 FrameData[24]
rlabel metal3 894 8484 894 8484 0 FrameData[25]
rlabel metal2 1728 5628 1728 5628 0 FrameData[26]
rlabel metal2 1248 8568 1248 8568 0 FrameData[27]
rlabel metal4 1248 9072 1248 9072 0 FrameData[28]
rlabel metal4 13824 7770 13824 7770 0 FrameData[29]
rlabel metal3 126 756 126 756 0 FrameData[2]
rlabel metal3 318 10164 318 10164 0 FrameData[30]
rlabel metal3 174 10500 174 10500 0 FrameData[31]
rlabel metal3 654 1092 654 1092 0 FrameData[3]
rlabel metal2 39552 1134 39552 1134 0 FrameData[4]
rlabel metal4 34656 1008 34656 1008 0 FrameData[5]
rlabel metal2 19872 6510 19872 6510 0 FrameData[6]
rlabel metal2 34848 4998 34848 4998 0 FrameData[7]
rlabel metal3 606 2772 606 2772 0 FrameData[8]
rlabel metal3 1182 3108 1182 3108 0 FrameData[9]
rlabel metal2 41472 504 41472 504 0 FrameData_O[0]
rlabel metal3 42018 3444 42018 3444 0 FrameData_O[10]
rlabel metal3 42210 3780 42210 3780 0 FrameData_O[11]
rlabel metal3 41826 4116 41826 4116 0 FrameData_O[12]
rlabel metal2 41088 4410 41088 4410 0 FrameData_O[13]
rlabel metal3 42210 4788 42210 4788 0 FrameData_O[14]
rlabel metal2 40704 4956 40704 4956 0 FrameData_O[15]
rlabel metal2 41088 5124 41088 5124 0 FrameData_O[16]
rlabel metal3 41826 5796 41826 5796 0 FrameData_O[17]
rlabel metal2 41088 6006 41088 6006 0 FrameData_O[18]
rlabel metal3 42018 6468 42018 6468 0 FrameData_O[19]
rlabel metal2 40704 672 40704 672 0 FrameData_O[1]
rlabel metal2 40704 6720 40704 6720 0 FrameData_O[20]
rlabel metal3 42018 7140 42018 7140 0 FrameData_O[21]
rlabel metal2 40704 7434 40704 7434 0 FrameData_O[22]
rlabel metal3 42018 7812 42018 7812 0 FrameData_O[23]
rlabel metal3 41826 8148 41826 8148 0 FrameData_O[24]
rlabel metal2 41472 8316 41472 8316 0 FrameData_O[25]
rlabel metal3 42018 8820 42018 8820 0 FrameData_O[26]
rlabel metal2 41472 8946 41472 8946 0 FrameData_O[27]
rlabel metal3 42018 9492 42018 9492 0 FrameData_O[28]
rlabel metal2 40032 9324 40032 9324 0 FrameData_O[29]
rlabel metal2 40320 840 40320 840 0 FrameData_O[2]
rlabel metal2 41472 9912 41472 9912 0 FrameData_O[30]
rlabel metal2 40704 10080 40704 10080 0 FrameData_O[31]
rlabel metal3 41634 1092 41634 1092 0 FrameData_O[3]
rlabel metal2 38976 1764 38976 1764 0 FrameData_O[4]
rlabel metal2 41088 1512 41088 1512 0 FrameData_O[5]
rlabel metal3 42258 2100 42258 2100 0 FrameData_O[6]
rlabel metal3 42210 2436 42210 2436 0 FrameData_O[7]
rlabel metal3 42018 2772 42018 2772 0 FrameData_O[8]
rlabel metal3 41826 3108 41826 3108 0 FrameData_O[9]
rlabel metal2 40416 2184 40416 2184 0 FrameStrobe[0]
rlabel metal2 31776 534 31776 534 0 FrameStrobe[10]
rlabel metal2 31968 324 31968 324 0 FrameStrobe[11]
rlabel metal3 33276 1848 33276 1848 0 FrameStrobe[12]
rlabel metal2 32352 366 32352 366 0 FrameStrobe[13]
rlabel metal2 32544 954 32544 954 0 FrameStrobe[14]
rlabel metal2 32736 114 32736 114 0 FrameStrobe[15]
rlabel metal2 32928 408 32928 408 0 FrameStrobe[16]
rlabel metal2 33120 1248 33120 1248 0 FrameStrobe[17]
rlabel metal2 33312 324 33312 324 0 FrameStrobe[18]
rlabel metal2 33504 72 33504 72 0 FrameStrobe[19]
rlabel metal2 33408 1512 33408 1512 0 FrameStrobe[1]
rlabel metal2 30192 2016 30192 2016 0 FrameStrobe[2]
rlabel metal2 30432 492 30432 492 0 FrameStrobe[3]
rlabel metal2 30624 618 30624 618 0 FrameStrobe[4]
rlabel metal2 30816 408 30816 408 0 FrameStrobe[5]
rlabel metal2 31008 450 31008 450 0 FrameStrobe[6]
rlabel metal2 31200 408 31200 408 0 FrameStrobe[7]
rlabel metal2 31392 492 31392 492 0 FrameStrobe[8]
rlabel metal2 31584 912 31584 912 0 FrameStrobe[9]
rlabel metal2 19488 10186 19488 10186 0 FrameStrobe_O[0]
rlabel metal3 31536 8820 31536 8820 0 FrameStrobe_O[10]
rlabel metal2 32544 9766 32544 9766 0 FrameStrobe_O[11]
rlabel metal2 32928 9756 32928 9756 0 FrameStrobe_O[12]
rlabel metal3 33840 8148 33840 8148 0 FrameStrobe_O[13]
rlabel metal3 35616 8820 35616 8820 0 FrameStrobe_O[14]
rlabel metal2 36528 8820 36528 8820 0 FrameStrobe_O[15]
rlabel metal2 37728 9828 37728 9828 0 FrameStrobe_O[16]
rlabel metal2 38736 8820 38736 8820 0 FrameStrobe_O[17]
rlabel metal2 39168 9198 39168 9198 0 FrameStrobe_O[18]
rlabel metal2 40416 9766 40416 9766 0 FrameStrobe_O[19]
rlabel metal2 20016 8820 20016 8820 0 FrameStrobe_O[1]
rlabel metal2 21408 10176 21408 10176 0 FrameStrobe_O[2]
rlabel metal2 22608 8148 22608 8148 0 FrameStrobe_O[3]
rlabel metal2 29760 9660 29760 9660 0 FrameStrobe_O[4]
rlabel metal2 32064 9828 32064 9828 0 FrameStrobe_O[5]
rlabel metal2 30624 8442 30624 8442 0 FrameStrobe_O[6]
rlabel metal2 32448 9870 32448 9870 0 FrameStrobe_O[7]
rlabel metal2 31776 8862 31776 8862 0 FrameStrobe_O[8]
rlabel metal2 32832 9786 32832 9786 0 FrameStrobe_O[9]
rlabel metal2 36000 7140 36000 7140 0 Inst_A_IO_1_bidirectional_frame_config_pass.Q
rlabel metal2 32352 1428 32352 1428 0 Inst_B_IO_1_bidirectional_frame_config_pass.Q
rlabel metal2 7104 1971 7104 1971 0 Inst_N_IO_ConfigMem.Inst_frame0_bit0.Q
rlabel metal2 2736 924 2736 924 0 Inst_N_IO_ConfigMem.Inst_frame0_bit1.Q
rlabel metal3 38496 3948 38496 3948 0 Inst_N_IO_ConfigMem.Inst_frame0_bit10.Q
rlabel metal3 40080 4368 40080 4368 0 Inst_N_IO_ConfigMem.Inst_frame0_bit11.Q
rlabel metal2 35616 5292 35616 5292 0 Inst_N_IO_ConfigMem.Inst_frame0_bit12.Q
rlabel metal2 37344 5376 37344 5376 0 Inst_N_IO_ConfigMem.Inst_frame0_bit13.Q
rlabel metal2 6816 1393 6816 1393 0 Inst_N_IO_ConfigMem.Inst_frame0_bit14.Q
rlabel metal2 5280 1050 5280 1050 0 Inst_N_IO_ConfigMem.Inst_frame0_bit15.Q
rlabel metal2 9408 2181 9408 2181 0 Inst_N_IO_ConfigMem.Inst_frame0_bit16.Q
rlabel metal3 7632 1932 7632 1932 0 Inst_N_IO_ConfigMem.Inst_frame0_bit17.Q
rlabel metal3 4704 2436 4704 2436 0 Inst_N_IO_ConfigMem.Inst_frame0_bit18.Q
rlabel metal3 4128 4914 4128 4914 0 Inst_N_IO_ConfigMem.Inst_frame0_bit19.Q
rlabel metal3 36672 1260 36672 1260 0 Inst_N_IO_ConfigMem.Inst_frame0_bit2.Q
rlabel metal2 4608 3402 4608 3402 0 Inst_N_IO_ConfigMem.Inst_frame0_bit20.Q
rlabel metal2 3360 2940 3360 2940 0 Inst_N_IO_ConfigMem.Inst_frame0_bit21.Q
rlabel metal3 3744 8568 3744 8568 0 Inst_N_IO_ConfigMem.Inst_frame0_bit22.Q
rlabel metal3 3504 8652 3504 8652 0 Inst_N_IO_ConfigMem.Inst_frame0_bit23.Q
rlabel metal2 3936 9534 3936 9534 0 Inst_N_IO_ConfigMem.Inst_frame0_bit24.Q
rlabel metal3 3552 6468 3552 6468 0 Inst_N_IO_ConfigMem.Inst_frame0_bit25.Q
rlabel via2 7200 5630 7200 5630 0 Inst_N_IO_ConfigMem.Inst_frame0_bit26.Q
rlabel metal4 5376 6972 5376 6972 0 Inst_N_IO_ConfigMem.Inst_frame0_bit27.Q
rlabel metal2 6240 7812 6240 7812 0 Inst_N_IO_ConfigMem.Inst_frame0_bit28.Q
rlabel metal2 7392 8022 7392 8022 0 Inst_N_IO_ConfigMem.Inst_frame0_bit29.Q
rlabel metal3 35088 1260 35088 1260 0 Inst_N_IO_ConfigMem.Inst_frame0_bit3.Q
rlabel via1 8880 7144 8880 7144 0 Inst_N_IO_ConfigMem.Inst_frame0_bit30.Q
rlabel metal2 6816 7182 6816 7182 0 Inst_N_IO_ConfigMem.Inst_frame0_bit31.Q
rlabel metal2 38208 1344 38208 1344 0 Inst_N_IO_ConfigMem.Inst_frame0_bit4.Q
rlabel via1 39840 1927 39840 1927 0 Inst_N_IO_ConfigMem.Inst_frame0_bit5.Q
rlabel metal2 31968 5208 31968 5208 0 Inst_N_IO_ConfigMem.Inst_frame0_bit6.Q
rlabel metal2 33456 4368 33456 4368 0 Inst_N_IO_ConfigMem.Inst_frame0_bit7.Q
rlabel metal3 36288 2604 36288 2604 0 Inst_N_IO_ConfigMem.Inst_frame0_bit8.Q
rlabel via2 37632 2606 37632 2606 0 Inst_N_IO_ConfigMem.Inst_frame0_bit9.Q
rlabel metal2 12192 1218 12192 1218 0 Inst_N_IO_ConfigMem.Inst_frame1_bit0.Q
rlabel metal2 16704 1631 16704 1631 0 Inst_N_IO_ConfigMem.Inst_frame1_bit1.Q
rlabel metal2 27168 2940 27168 2940 0 Inst_N_IO_ConfigMem.Inst_frame1_bit10.Q
rlabel metal2 24960 3486 24960 3486 0 Inst_N_IO_ConfigMem.Inst_frame1_bit11.Q
rlabel metal2 33120 7476 33120 7476 0 Inst_N_IO_ConfigMem.Inst_frame1_bit12.Q
rlabel metal2 31104 8232 31104 8232 0 Inst_N_IO_ConfigMem.Inst_frame1_bit13.Q
rlabel metal2 27552 4158 27552 4158 0 Inst_N_IO_ConfigMem.Inst_frame1_bit14.Q
rlabel metal2 29376 3612 29376 3612 0 Inst_N_IO_ConfigMem.Inst_frame1_bit15.Q
rlabel metal2 31296 1050 31296 1050 0 Inst_N_IO_ConfigMem.Inst_frame1_bit16.Q
rlabel metal2 32832 1393 32832 1393 0 Inst_N_IO_ConfigMem.Inst_frame1_bit17.Q
rlabel metal2 31872 5586 31872 5586 0 Inst_N_IO_ConfigMem.Inst_frame1_bit18.Q
rlabel metal2 33408 5929 33408 5929 0 Inst_N_IO_ConfigMem.Inst_frame1_bit19.Q
rlabel metal2 24960 1512 24960 1512 0 Inst_N_IO_ConfigMem.Inst_frame1_bit2.Q
rlabel metal2 36192 3486 36192 3486 0 Inst_N_IO_ConfigMem.Inst_frame1_bit20.Q
rlabel via2 37728 3441 37728 3441 0 Inst_N_IO_ConfigMem.Inst_frame1_bit21.Q
rlabel metal2 38016 7812 38016 7812 0 Inst_N_IO_ConfigMem.Inst_frame1_bit22.Q
rlabel metal2 39504 6636 39504 6636 0 Inst_N_IO_ConfigMem.Inst_frame1_bit23.Q
rlabel metal2 35136 7098 35136 7098 0 Inst_N_IO_ConfigMem.Inst_frame1_bit24.Q
rlabel metal2 36672 7441 36672 7441 0 Inst_N_IO_ConfigMem.Inst_frame1_bit25.Q
rlabel metal2 11328 7812 11328 7812 0 Inst_N_IO_ConfigMem.Inst_frame1_bit26.Q
rlabel metal2 12864 7441 12864 7441 0 Inst_N_IO_ConfigMem.Inst_frame1_bit27.Q
rlabel metal2 13824 7434 13824 7434 0 Inst_N_IO_ConfigMem.Inst_frame1_bit28.Q
rlabel metal2 15360 7441 15360 7441 0 Inst_N_IO_ConfigMem.Inst_frame1_bit29.Q
rlabel metal3 25968 1344 25968 1344 0 Inst_N_IO_ConfigMem.Inst_frame1_bit3.Q
rlabel metal2 11616 5929 11616 5929 0 Inst_N_IO_ConfigMem.Inst_frame1_bit30.Q
rlabel metal2 10080 5586 10080 5586 0 Inst_N_IO_ConfigMem.Inst_frame1_bit31.Q
rlabel metal2 30576 1344 30576 1344 0 Inst_N_IO_ConfigMem.Inst_frame1_bit4.Q
rlabel metal2 32064 1589 32064 1589 0 Inst_N_IO_ConfigMem.Inst_frame1_bit5.Q
rlabel metal2 29232 5691 29232 5691 0 Inst_N_IO_ConfigMem.Inst_frame1_bit6.Q
rlabel metal2 27648 5964 27648 5964 0 Inst_N_IO_ConfigMem.Inst_frame1_bit7.Q
rlabel metal3 33120 2772 33120 2772 0 Inst_N_IO_ConfigMem.Inst_frame1_bit8.Q
rlabel metal2 31776 3486 31776 3486 0 Inst_N_IO_ConfigMem.Inst_frame1_bit9.Q
rlabel metal2 17424 1932 17424 1932 0 Inst_N_IO_ConfigMem.Inst_frame2_bit0.Q
rlabel metal2 18768 1260 18768 1260 0 Inst_N_IO_ConfigMem.Inst_frame2_bit1.Q
rlabel metal2 21984 8610 21984 8610 0 Inst_N_IO_ConfigMem.Inst_frame2_bit10.Q
rlabel via1 23568 8656 23568 8656 0 Inst_N_IO_ConfigMem.Inst_frame2_bit11.Q
rlabel metal2 14016 4074 14016 4074 0 Inst_N_IO_ConfigMem.Inst_frame2_bit12.Q
rlabel metal2 15648 3864 15648 3864 0 Inst_N_IO_ConfigMem.Inst_frame2_bit13.Q
rlabel metal2 21120 3864 21120 3864 0 Inst_N_IO_ConfigMem.Inst_frame2_bit14.Q
rlabel metal3 22752 3612 22752 3612 0 Inst_N_IO_ConfigMem.Inst_frame2_bit15.Q
rlabel metal3 27552 1932 27552 1932 0 Inst_N_IO_ConfigMem.Inst_frame2_bit16.Q
rlabel via2 29280 1929 29280 1929 0 Inst_N_IO_ConfigMem.Inst_frame2_bit17.Q
rlabel metal2 23424 4998 23424 4998 0 Inst_N_IO_ConfigMem.Inst_frame2_bit18.Q
rlabel metal2 24288 4578 24288 4578 0 Inst_N_IO_ConfigMem.Inst_frame2_bit19.Q
rlabel metal2 20400 1344 20400 1344 0 Inst_N_IO_ConfigMem.Inst_frame2_bit2.Q
rlabel metal2 13872 1260 13872 1260 0 Inst_N_IO_ConfigMem.Inst_frame2_bit20.Q
rlabel metal3 15168 2100 15168 2100 0 Inst_N_IO_ConfigMem.Inst_frame2_bit21.Q
rlabel metal2 26304 7476 26304 7476 0 Inst_N_IO_ConfigMem.Inst_frame2_bit22.Q
rlabel metal2 25632 7434 25632 7434 0 Inst_N_IO_ConfigMem.Inst_frame2_bit23.Q
rlabel metal2 17856 4113 17856 4113 0 Inst_N_IO_ConfigMem.Inst_frame2_bit24.Q
rlabel metal2 16320 4830 16320 4830 0 Inst_N_IO_ConfigMem.Inst_frame2_bit25.Q
rlabel metal2 25560 5670 25560 5670 0 Inst_N_IO_ConfigMem.Inst_frame2_bit26.Q
rlabel metal2 23904 6678 23904 6678 0 Inst_N_IO_ConfigMem.Inst_frame2_bit27.Q
rlabel metal2 12672 4071 12672 4071 0 Inst_N_IO_ConfigMem.Inst_frame2_bit28.Q
rlabel metal2 11136 3486 11136 3486 0 Inst_N_IO_ConfigMem.Inst_frame2_bit29.Q
rlabel metal3 22032 1344 22032 1344 0 Inst_N_IO_ConfigMem.Inst_frame2_bit3.Q
rlabel metal2 25440 8946 25440 8946 0 Inst_N_IO_ConfigMem.Inst_frame2_bit30.Q
rlabel via1 27024 8656 27024 8656 0 Inst_N_IO_ConfigMem.Inst_frame2_bit31.Q
rlabel metal3 10848 1344 10848 1344 0 Inst_N_IO_ConfigMem.Inst_frame2_bit4.Q
rlabel metal2 12672 2013 12672 2013 0 Inst_N_IO_ConfigMem.Inst_frame2_bit5.Q
rlabel metal2 21600 6552 21600 6552 0 Inst_N_IO_ConfigMem.Inst_frame2_bit6.Q
rlabel metal2 23472 5880 23472 5880 0 Inst_N_IO_ConfigMem.Inst_frame2_bit7.Q
rlabel metal2 29184 8652 29184 8652 0 Inst_N_IO_ConfigMem.Inst_frame2_bit8.Q
rlabel metal2 30336 7644 30336 7644 0 Inst_N_IO_ConfigMem.Inst_frame2_bit9.Q
rlabel metal2 18768 4368 18768 4368 0 Inst_N_IO_ConfigMem.Inst_frame3_bit18.Q
rlabel metal2 20688 4368 20688 4368 0 Inst_N_IO_ConfigMem.Inst_frame3_bit19.Q
rlabel metal2 10944 3108 10944 3108 0 Inst_N_IO_ConfigMem.Inst_frame3_bit20.Q
rlabel metal2 12480 3283 12480 3283 0 Inst_N_IO_ConfigMem.Inst_frame3_bit21.Q
rlabel metal2 17952 6594 17952 6594 0 Inst_N_IO_ConfigMem.Inst_frame3_bit22.Q
rlabel metal2 19488 6167 19488 6167 0 Inst_N_IO_ConfigMem.Inst_frame3_bit23.Q
rlabel metal2 19296 7434 19296 7434 0 Inst_N_IO_ConfigMem.Inst_frame3_bit24.Q
rlabel metal2 20880 7203 20880 7203 0 Inst_N_IO_ConfigMem.Inst_frame3_bit25.Q
rlabel metal2 17664 8610 17664 8610 0 Inst_N_IO_ConfigMem.Inst_frame3_bit26.Q
rlabel metal2 19248 8715 19248 8715 0 Inst_N_IO_ConfigMem.Inst_frame3_bit27.Q
rlabel metal2 13920 5586 13920 5586 0 Inst_N_IO_ConfigMem.Inst_frame3_bit28.Q
rlabel metal2 15456 5205 15456 5205 0 Inst_N_IO_ConfigMem.Inst_frame3_bit29.Q
rlabel metal3 16512 4956 16512 4956 0 Inst_N_IO_ConfigMem.Inst_frame3_bit30.Q
rlabel metal2 18336 5205 18336 5205 0 Inst_N_IO_ConfigMem.Inst_frame3_bit31.Q
rlabel metal3 8976 4368 8976 4368 0 Inst_N_IO_switch_matrix.DEBUG_select_S1BEG0[0]
rlabel metal2 23856 2016 23856 2016 0 Inst_N_IO_switch_matrix.DEBUG_select_S1BEG1[0]
rlabel metal2 19632 2604 19632 2604 0 Inst_N_IO_switch_matrix.DEBUG_select_S1BEG2[0]
rlabel metal2 30624 4410 30624 4410 0 Inst_N_IO_switch_matrix.DEBUG_select_S1BEG3[0]
rlabel metal3 9840 2436 9840 2436 0 Inst_N_IO_switch_matrix.S1BEG0
rlabel metal2 24384 2772 24384 2772 0 Inst_N_IO_switch_matrix.S1BEG1
rlabel metal4 19968 2352 19968 2352 0 Inst_N_IO_switch_matrix.S1BEG2
rlabel metal2 31104 1176 31104 1176 0 Inst_N_IO_switch_matrix.S1BEG3
rlabel metal2 20784 2688 20784 2688 0 Inst_N_IO_switch_matrix.S2BEG0
rlabel metal2 13056 2142 13056 2142 0 Inst_N_IO_switch_matrix.S2BEG1
rlabel metal2 19680 6132 19680 6132 0 Inst_N_IO_switch_matrix.S2BEG2
rlabel metal2 21408 7266 21408 7266 0 Inst_N_IO_switch_matrix.S2BEG3
rlabel metal2 19392 8190 19392 8190 0 Inst_N_IO_switch_matrix.S2BEG4
rlabel metal2 15648 4914 15648 4914 0 Inst_N_IO_switch_matrix.S2BEG5
rlabel metal3 18528 4998 18528 4998 0 Inst_N_IO_switch_matrix.S2BEG6
rlabel metal2 19248 2100 19248 2100 0 Inst_N_IO_switch_matrix.S2BEG7
rlabel metal2 22128 2100 22128 2100 0 Inst_N_IO_switch_matrix.S2BEGb0
rlabel metal3 17184 2016 17184 2016 0 Inst_N_IO_switch_matrix.S2BEGb1
rlabel metal2 23712 6468 23712 6468 0 Inst_N_IO_switch_matrix.S2BEGb2
rlabel metal2 30624 7224 30624 7224 0 Inst_N_IO_switch_matrix.S2BEGb3
rlabel metal2 23424 7854 23424 7854 0 Inst_N_IO_switch_matrix.S2BEGb4
rlabel metal3 18624 5082 18624 5082 0 Inst_N_IO_switch_matrix.S2BEGb5
rlabel metal2 22944 3318 22944 3318 0 Inst_N_IO_switch_matrix.S2BEGb6
rlabel metal3 29856 1848 29856 1848 0 Inst_N_IO_switch_matrix.S2BEGb7
rlabel metal3 24624 4200 24624 4200 0 Inst_N_IO_switch_matrix.S4BEG0
rlabel metal2 15648 2688 15648 2688 0 Inst_N_IO_switch_matrix.S4BEG1
rlabel metal2 29760 5670 29760 5670 0 Inst_N_IO_switch_matrix.S4BEG10
rlabel metal3 34080 3528 34080 3528 0 Inst_N_IO_switch_matrix.S4BEG11
rlabel metal2 25344 3108 25344 3108 0 Inst_N_IO_switch_matrix.S4BEG12
rlabel metal3 32592 6384 32592 6384 0 Inst_N_IO_switch_matrix.S4BEG13
rlabel metal2 29664 4158 29664 4158 0 Inst_N_IO_switch_matrix.S4BEG14
rlabel metal2 32784 2688 32784 2688 0 Inst_N_IO_switch_matrix.S4BEG15
rlabel metal2 26352 6384 26352 6384 0 Inst_N_IO_switch_matrix.S4BEG2
rlabel metal2 23328 3108 23328 3108 0 Inst_N_IO_switch_matrix.S4BEG3
rlabel metal2 25536 5166 25536 5166 0 Inst_N_IO_switch_matrix.S4BEG4
rlabel metal3 16512 3612 16512 3612 0 Inst_N_IO_switch_matrix.S4BEG5
rlabel metal2 27360 7896 27360 7896 0 Inst_N_IO_switch_matrix.S4BEG6
rlabel metal2 16992 3276 16992 3276 0 Inst_N_IO_switch_matrix.S4BEG7
rlabel metal2 26880 1932 26880 1932 0 Inst_N_IO_switch_matrix.S4BEG8
rlabel metal2 32640 1932 32640 1932 0 Inst_N_IO_switch_matrix.S4BEG9
rlabel metal2 33216 4830 33216 4830 0 Inst_N_IO_switch_matrix.SS4BEG0
rlabel metal2 38208 3108 38208 3108 0 Inst_N_IO_switch_matrix.SS4BEG1
rlabel metal3 33264 4200 33264 4200 0 Inst_N_IO_switch_matrix.SS4BEG10
rlabel metal2 37728 2184 37728 2184 0 Inst_N_IO_switch_matrix.SS4BEG11
rlabel metal2 39984 3360 39984 3360 0 Inst_N_IO_switch_matrix.SS4BEG12
rlabel metal2 36864 4830 36864 4830 0 Inst_N_IO_switch_matrix.SS4BEG13
rlabel metal4 18912 798 18912 798 0 Inst_N_IO_switch_matrix.SS4BEG14
rlabel metal2 29856 1938 29856 1938 0 Inst_N_IO_switch_matrix.SS4BEG15
rlabel metal2 39792 6384 39792 6384 0 Inst_N_IO_switch_matrix.SS4BEG2
rlabel metal3 36720 6384 36720 6384 0 Inst_N_IO_switch_matrix.SS4BEG3
rlabel metal2 25920 7098 25920 7098 0 Inst_N_IO_switch_matrix.SS4BEG4
rlabel metal2 15552 6258 15552 6258 0 Inst_N_IO_switch_matrix.SS4BEG5
rlabel metal4 24000 5250 24000 5250 0 Inst_N_IO_switch_matrix.SS4BEG6
rlabel metal5 9448 1974 9448 1974 0 Inst_N_IO_switch_matrix.SS4BEG7
rlabel metal2 37056 2184 37056 2184 0 Inst_N_IO_switch_matrix.SS4BEG8
rlabel metal2 39984 1176 39984 1176 0 Inst_N_IO_switch_matrix.SS4BEG9
rlabel metal2 30624 1880 30624 1880 0 N1END[0]
rlabel metal4 15264 2352 15264 2352 0 N1END[1]
rlabel metal3 15360 2226 15360 2226 0 N1END[2]
rlabel metal2 14016 3024 14016 3024 0 N1END[3]
rlabel metal3 19776 2478 19776 2478 0 N2END[0]
rlabel metal2 12000 492 12000 492 0 N2END[1]
rlabel metal2 12192 408 12192 408 0 N2END[2]
rlabel metal2 12384 450 12384 450 0 N2END[3]
rlabel metal3 11904 7224 11904 7224 0 N2END[4]
rlabel metal3 16944 7224 16944 7224 0 N2END[5]
rlabel metal2 12960 828 12960 828 0 N2END[6]
rlabel metal3 15120 2856 15120 2856 0 N2END[7]
rlabel metal3 17568 1890 17568 1890 0 N2MID[0]
rlabel metal2 16896 4326 16896 4326 0 N2MID[1]
rlabel metal2 14016 4830 14016 4830 0 N2MID[2]
rlabel metal2 17856 6510 17856 6510 0 N2MID[3]
rlabel metal4 19392 6426 19392 6426 0 N2MID[4]
rlabel metal2 18048 6300 18048 6300 0 N2MID[5]
rlabel metal2 11424 660 11424 660 0 N2MID[6]
rlabel metal4 11616 1806 11616 1806 0 N2MID[7]
rlabel metal2 31392 1218 31392 1218 0 N4END[0]
rlabel metal2 15264 450 15264 450 0 N4END[10]
rlabel metal2 15456 660 15456 660 0 N4END[11]
rlabel metal2 15648 492 15648 492 0 N4END[12]
rlabel metal2 15840 366 15840 366 0 N4END[13]
rlabel metal2 16032 156 16032 156 0 N4END[14]
rlabel metal2 16224 240 16224 240 0 N4END[15]
rlabel metal2 13536 1290 13536 1290 0 N4END[1]
rlabel metal3 14496 2604 14496 2604 0 N4END[2]
rlabel metal2 38736 1932 38736 1932 0 N4END[3]
rlabel metal3 35568 1932 35568 1932 0 N4END[4]
rlabel metal2 18432 6552 18432 6552 0 N4END[5]
rlabel metal3 34944 1848 34944 1848 0 N4END[6]
rlabel metal2 39312 1932 39312 1932 0 N4END[7]
rlabel metal2 35808 1974 35808 1974 0 N4END[8]
rlabel metal2 14976 3612 14976 3612 0 N4END[9]
rlabel metal2 31776 1470 31776 1470 0 NN4END[0]
rlabel metal2 18336 576 18336 576 0 NN4END[10]
rlabel metal2 18528 660 18528 660 0 NN4END[11]
rlabel metal2 18720 492 18720 492 0 NN4END[12]
rlabel metal2 28128 2268 28128 2268 0 NN4END[13]
rlabel metal2 15744 1638 15744 1638 0 NN4END[14]
rlabel metal2 19296 408 19296 408 0 NN4END[15]
rlabel metal2 17376 4578 17376 4578 0 NN4END[1]
rlabel metal2 15648 1806 15648 1806 0 NN4END[2]
rlabel metal3 17472 8652 17472 8652 0 NN4END[3]
rlabel metal2 17184 1080 17184 1080 0 NN4END[4]
rlabel metal2 17376 492 17376 492 0 NN4END[5]
rlabel metal2 11712 1680 11712 1680 0 NN4END[6]
rlabel metal2 17760 618 17760 618 0 NN4END[7]
rlabel metal2 18528 1764 18528 1764 0 NN4END[8]
rlabel metal2 17856 5124 17856 5124 0 NN4END[9]
rlabel metal2 19680 450 19680 450 0 S1BEG[0]
rlabel metal2 19872 324 19872 324 0 S1BEG[1]
rlabel metal2 20064 324 20064 324 0 S1BEG[2]
rlabel metal2 30912 546 30912 546 0 S1BEG[3]
rlabel metal2 20544 1512 20544 1512 0 S2BEG[0]
rlabel metal2 19296 1302 19296 1302 0 S2BEG[1]
rlabel metal2 20832 702 20832 702 0 S2BEG[2]
rlabel metal2 21024 1752 21024 1752 0 S2BEG[3]
rlabel metal2 21216 660 21216 660 0 S2BEG[4]
rlabel metal2 21408 660 21408 660 0 S2BEG[5]
rlabel metal2 21552 3612 21552 3612 0 S2BEG[6]
rlabel metal2 21120 1806 21120 1806 0 S2BEG[7]
rlabel metal2 21984 1890 21984 1890 0 S2BEGb[0]
rlabel metal2 21696 1722 21696 1722 0 S2BEGb[1]
rlabel metal3 22992 4368 22992 4368 0 S2BEGb[2]
rlabel metal2 30432 5418 30432 5418 0 S2BEGb[3]
rlabel metal2 22992 6972 22992 6972 0 S2BEGb[4]
rlabel metal2 22944 534 22944 534 0 S2BEGb[5]
rlabel metal2 23184 2436 23184 2436 0 S2BEGb[6]
rlabel metal2 30048 1596 30048 1596 0 S2BEGb[7]
rlabel metal2 23520 492 23520 492 0 S4BEG[0]
rlabel metal2 29568 5292 29568 5292 0 S4BEG[10]
rlabel metal2 34464 966 34464 966 0 S4BEG[11]
rlabel metal2 25536 1680 25536 1680 0 S4BEG[12]
rlabel metal2 31776 4998 31776 4998 0 S4BEG[13]
rlabel metal2 26208 1374 26208 1374 0 S4BEG[14]
rlabel metal2 32496 2436 32496 2436 0 S4BEG[15]
rlabel metal2 23712 492 23712 492 0 S4BEG[1]
rlabel metal2 23904 870 23904 870 0 S4BEG[2]
rlabel metal2 23520 2058 23520 2058 0 S4BEG[3]
rlabel metal2 24288 660 24288 660 0 S4BEG[4]
rlabel metal3 24000 2604 24000 2604 0 S4BEG[5]
rlabel metal2 24672 1290 24672 1290 0 S4BEG[6]
rlabel metal2 24912 2436 24912 2436 0 S4BEG[7]
rlabel metal2 25056 450 25056 450 0 S4BEG[8]
rlabel metal2 25248 324 25248 324 0 S4BEG[9]
rlabel metal3 33132 1092 33132 1092 0 SS4BEG[0]
rlabel metal3 32448 2604 32448 2604 0 SS4BEG[10]
rlabel metal2 37536 1008 37536 1008 0 SS4BEG[11]
rlabel metal2 28896 1122 28896 1122 0 SS4BEG[12]
rlabel metal3 32880 3948 32880 3948 0 SS4BEG[13]
rlabel metal2 29280 492 29280 492 0 SS4BEG[14]
rlabel metal2 29472 870 29472 870 0 SS4BEG[15]
rlabel metal2 38016 2016 38016 2016 0 SS4BEG[1]
rlabel metal2 26976 660 26976 660 0 SS4BEG[2]
rlabel metal2 27168 1290 27168 1290 0 SS4BEG[3]
rlabel metal2 27360 618 27360 618 0 SS4BEG[4]
rlabel metal2 27552 954 27552 954 0 SS4BEG[5]
rlabel metal2 27744 660 27744 660 0 SS4BEG[6]
rlabel metal2 27936 492 27936 492 0 SS4BEG[7]
rlabel metal2 35616 1428 35616 1428 0 SS4BEG[8]
rlabel metal2 39744 504 39744 504 0 SS4BEG[9]
rlabel metal2 29664 786 29664 786 0 UserCLK
rlabel metal3 36528 9492 36528 9492 0 UserCLK_regs
rlabel via2 17952 10680 17952 10680 0 UserCLKo
rlabel metal2 4560 5124 4560 5124 0 _000_
rlabel metal2 3648 7938 3648 7938 0 _001_
rlabel metal2 4891 6342 4891 6342 0 _002_
rlabel metal3 4848 6468 4848 6468 0 _003_
rlabel metal3 4704 5880 4704 5880 0 _004_
rlabel metal2 5760 6888 5760 6888 0 _005_
rlabel metal3 5280 4704 5280 4704 0 _006_
rlabel metal2 5088 5964 5088 5964 0 _007_
rlabel metal2 5376 5880 5376 5880 0 _008_
rlabel metal2 4896 5964 4896 5964 0 _009_
rlabel metal2 6144 6552 6144 6552 0 _010_
rlabel metal2 6336 6720 6336 6720 0 _011_
rlabel metal2 5568 7224 5568 7224 0 _012_
rlabel metal2 7392 6090 7392 6090 0 _013_
rlabel metal2 7200 5040 7200 5040 0 _014_
rlabel metal2 6384 7140 6384 7140 0 _015_
rlabel metal3 6240 6972 6240 6972 0 _016_
rlabel via1 4180 3444 4180 3444 0 _017_
rlabel metal2 3936 3528 3936 3528 0 _018_
rlabel metal2 3744 3696 3744 3696 0 _019_
rlabel metal2 4032 3738 4032 3738 0 _020_
rlabel metal2 3360 3570 3360 3570 0 _021_
rlabel metal2 4416 3276 4416 3276 0 _022_
rlabel metal2 3552 2646 3552 2646 0 _023_
rlabel metal2 4848 2856 4848 2856 0 _024_
rlabel metal3 4848 3444 4848 3444 0 _025_
rlabel metal3 3792 2604 3792 2604 0 _026_
rlabel metal2 3264 2814 3264 2814 0 _027_
rlabel metal2 7872 3486 7872 3486 0 _028_
rlabel metal2 7776 3738 7776 3738 0 _029_
rlabel metal2 3840 2646 3840 2646 0 _030_
rlabel metal3 3792 2856 3792 2856 0 _031_
rlabel metal2 4128 9156 4128 9156 0 _032_
rlabel metal2 4032 8778 4032 8778 0 _033_
rlabel metal2 3600 8904 3600 8904 0 _034_
rlabel metal3 4032 9492 4032 9492 0 _035_
rlabel metal2 3648 7224 3648 7224 0 _036_
rlabel metal2 2976 7224 2976 7224 0 _037_
rlabel metal2 3552 6594 3552 6594 0 _038_
rlabel metal2 3936 7392 3936 7392 0 _039_
rlabel metal2 6912 7224 6912 7224 0 _040_
rlabel metal2 9024 7098 9024 7098 0 _041_
rlabel metal2 9312 7392 9312 7392 0 _042_
rlabel metal3 7968 6972 7968 6972 0 _043_
rlabel metal2 9696 6972 9696 6972 0 _044_
rlabel metal2 33552 9324 33552 9324 0 _045_
rlabel metal2 34800 9324 34800 9324 0 _046_
rlabel metal2 30672 9492 30672 9492 0 clknet_0_UserCLK
rlabel metal2 35904 9156 35904 9156 0 clknet_0_UserCLK_regs
rlabel metal2 29472 9114 29472 9114 0 clknet_1_0__leaf_UserCLK
rlabel metal3 36336 7980 36336 7980 0 clknet_1_0__leaf_UserCLK_regs
rlabel metal2 34848 8904 34848 8904 0 clknet_1_1__leaf_UserCLK_regs
<< properties >>
string FIXED_BBOX 0 0 43008 10752
<< end >>
