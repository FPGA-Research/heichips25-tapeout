* NGSPICE file created from eFPGA.ext - technology: ihp-sg13g2

* Black-box entry subcircuit for LUT4AB abstract view
.subckt LUT4AB Ci Co E1BEG[0] E1BEG[1] E1BEG[2] E1BEG[3] E1END[0] E1END[1] E1END[2]
+ E1END[3] E2BEG[0] E2BEG[1] E2BEG[2] E2BEG[3] E2BEG[4] E2BEG[5] E2BEG[6] E2BEG[7]
+ E2BEGb[0] E2BEGb[1] E2BEGb[2] E2BEGb[3] E2BEGb[4] E2BEGb[5] E2BEGb[6] E2BEGb[7]
+ E2END[0] E2END[1] E2END[2] E2END[3] E2END[4] E2END[5] E2END[6] E2END[7] E2MID[0]
+ E2MID[1] E2MID[2] E2MID[3] E2MID[4] E2MID[5] E2MID[6] E2MID[7] E6BEG[0] E6BEG[10]
+ E6BEG[11] E6BEG[1] E6BEG[2] E6BEG[3] E6BEG[4] E6BEG[5] E6BEG[6] E6BEG[7] E6BEG[8]
+ E6BEG[9] E6END[0] E6END[10] E6END[11] E6END[1] E6END[2] E6END[3] E6END[4] E6END[5]
+ E6END[6] E6END[7] E6END[8] E6END[9] EE4BEG[0] EE4BEG[10] EE4BEG[11] EE4BEG[12] EE4BEG[13]
+ EE4BEG[14] EE4BEG[15] EE4BEG[1] EE4BEG[2] EE4BEG[3] EE4BEG[4] EE4BEG[5] EE4BEG[6]
+ EE4BEG[7] EE4BEG[8] EE4BEG[9] EE4END[0] EE4END[10] EE4END[11] EE4END[12] EE4END[13]
+ EE4END[14] EE4END[15] EE4END[1] EE4END[2] EE4END[3] EE4END[4] EE4END[5] EE4END[6]
+ EE4END[7] EE4END[8] EE4END[9] FrameData[0] FrameData[10] FrameData[11] FrameData[12]
+ FrameData[13] FrameData[14] FrameData[15] FrameData[16] FrameData[17] FrameData[18]
+ FrameData[19] FrameData[1] FrameData[20] FrameData[21] FrameData[22] FrameData[23]
+ FrameData[24] FrameData[25] FrameData[26] FrameData[27] FrameData[28] FrameData[29]
+ FrameData[2] FrameData[30] FrameData[31] FrameData[3] FrameData[4] FrameData[5]
+ FrameData[6] FrameData[7] FrameData[8] FrameData[9] FrameData_O[0] FrameData_O[10]
+ FrameData_O[11] FrameData_O[12] FrameData_O[13] FrameData_O[14] FrameData_O[15]
+ FrameData_O[16] FrameData_O[17] FrameData_O[18] FrameData_O[19] FrameData_O[1] FrameData_O[20]
+ FrameData_O[21] FrameData_O[22] FrameData_O[23] FrameData_O[24] FrameData_O[25]
+ FrameData_O[26] FrameData_O[27] FrameData_O[28] FrameData_O[29] FrameData_O[2] FrameData_O[30]
+ FrameData_O[31] FrameData_O[3] FrameData_O[4] FrameData_O[5] FrameData_O[6] FrameData_O[7]
+ FrameData_O[8] FrameData_O[9] FrameStrobe[0] FrameStrobe[10] FrameStrobe[11] FrameStrobe[12]
+ FrameStrobe[13] FrameStrobe[14] FrameStrobe[15] FrameStrobe[16] FrameStrobe[17]
+ FrameStrobe[18] FrameStrobe[19] FrameStrobe[1] FrameStrobe[2] FrameStrobe[3] FrameStrobe[4]
+ FrameStrobe[5] FrameStrobe[6] FrameStrobe[7] FrameStrobe[8] FrameStrobe[9] FrameStrobe_O[0]
+ FrameStrobe_O[10] FrameStrobe_O[11] FrameStrobe_O[12] FrameStrobe_O[13] FrameStrobe_O[14]
+ FrameStrobe_O[15] FrameStrobe_O[16] FrameStrobe_O[17] FrameStrobe_O[18] FrameStrobe_O[19]
+ FrameStrobe_O[1] FrameStrobe_O[2] FrameStrobe_O[3] FrameStrobe_O[4] FrameStrobe_O[5]
+ FrameStrobe_O[6] FrameStrobe_O[7] FrameStrobe_O[8] FrameStrobe_O[9] N1BEG[0] N1BEG[1]
+ N1BEG[2] N1BEG[3] N1END[0] N1END[1] N1END[2] N1END[3] N2BEG[0] N2BEG[1] N2BEG[2]
+ N2BEG[3] N2BEG[4] N2BEG[5] N2BEG[6] N2BEG[7] N2BEGb[0] N2BEGb[1] N2BEGb[2] N2BEGb[3]
+ N2BEGb[4] N2BEGb[5] N2BEGb[6] N2BEGb[7] N2END[0] N2END[1] N2END[2] N2END[3] N2END[4]
+ N2END[5] N2END[6] N2END[7] N2MID[0] N2MID[1] N2MID[2] N2MID[3] N2MID[4] N2MID[5]
+ N2MID[6] N2MID[7] N4BEG[0] N4BEG[10] N4BEG[11] N4BEG[12] N4BEG[13] N4BEG[14] N4BEG[15]
+ N4BEG[1] N4BEG[2] N4BEG[3] N4BEG[4] N4BEG[5] N4BEG[6] N4BEG[7] N4BEG[8] N4BEG[9]
+ N4END[0] N4END[10] N4END[11] N4END[12] N4END[13] N4END[14] N4END[15] N4END[1] N4END[2]
+ N4END[3] N4END[4] N4END[5] N4END[6] N4END[7] N4END[8] N4END[9] NN4BEG[0] NN4BEG[10]
+ NN4BEG[11] NN4BEG[12] NN4BEG[13] NN4BEG[14] NN4BEG[15] NN4BEG[1] NN4BEG[2] NN4BEG[3]
+ NN4BEG[4] NN4BEG[5] NN4BEG[6] NN4BEG[7] NN4BEG[8] NN4BEG[9] NN4END[0] NN4END[10]
+ NN4END[11] NN4END[12] NN4END[13] NN4END[14] NN4END[15] NN4END[1] NN4END[2] NN4END[3]
+ NN4END[4] NN4END[5] NN4END[6] NN4END[7] NN4END[8] NN4END[9] S1BEG[0] S1BEG[1] S1BEG[2]
+ S1BEG[3] S1END[0] S1END[1] S1END[2] S1END[3] S2BEG[0] S2BEG[1] S2BEG[2] S2BEG[3]
+ S2BEG[4] S2BEG[5] S2BEG[6] S2BEG[7] S2BEGb[0] S2BEGb[1] S2BEGb[2] S2BEGb[3] S2BEGb[4]
+ S2BEGb[5] S2BEGb[6] S2BEGb[7] S2END[0] S2END[1] S2END[2] S2END[3] S2END[4] S2END[5]
+ S2END[6] S2END[7] S2MID[0] S2MID[1] S2MID[2] S2MID[3] S2MID[4] S2MID[5] S2MID[6]
+ S2MID[7] S4BEG[0] S4BEG[10] S4BEG[11] S4BEG[12] S4BEG[13] S4BEG[14] S4BEG[15] S4BEG[1]
+ S4BEG[2] S4BEG[3] S4BEG[4] S4BEG[5] S4BEG[6] S4BEG[7] S4BEG[8] S4BEG[9] S4END[0]
+ S4END[10] S4END[11] S4END[12] S4END[13] S4END[14] S4END[15] S4END[1] S4END[2] S4END[3]
+ S4END[4] S4END[5] S4END[6] S4END[7] S4END[8] S4END[9] SS4BEG[0] SS4BEG[10] SS4BEG[11]
+ SS4BEG[12] SS4BEG[13] SS4BEG[14] SS4BEG[15] SS4BEG[1] SS4BEG[2] SS4BEG[3] SS4BEG[4]
+ SS4BEG[5] SS4BEG[6] SS4BEG[7] SS4BEG[8] SS4BEG[9] SS4END[0] SS4END[10] SS4END[11]
+ SS4END[12] SS4END[13] SS4END[14] SS4END[15] SS4END[1] SS4END[2] SS4END[3] SS4END[4]
+ SS4END[5] SS4END[6] SS4END[7] SS4END[8] SS4END[9] UserCLK UserCLKo VGND VPWR W1BEG[0]
+ W1BEG[1] W1BEG[2] W1BEG[3] W1END[0] W1END[1] W1END[2] W1END[3] W2BEG[0] W2BEG[1]
+ W2BEG[2] W2BEG[3] W2BEG[4] W2BEG[5] W2BEG[6] W2BEG[7] W2BEGb[0] W2BEGb[1] W2BEGb[2]
+ W2BEGb[3] W2BEGb[4] W2BEGb[5] W2BEGb[6] W2BEGb[7] W2END[0] W2END[1] W2END[2] W2END[3]
+ W2END[4] W2END[5] W2END[6] W2END[7] W2MID[0] W2MID[1] W2MID[2] W2MID[3] W2MID[4]
+ W2MID[5] W2MID[6] W2MID[7] W6BEG[0] W6BEG[10] W6BEG[11] W6BEG[1] W6BEG[2] W6BEG[3]
+ W6BEG[4] W6BEG[5] W6BEG[6] W6BEG[7] W6BEG[8] W6BEG[9] W6END[0] W6END[10] W6END[11]
+ W6END[1] W6END[2] W6END[3] W6END[4] W6END[5] W6END[6] W6END[7] W6END[8] W6END[9]
+ WW4BEG[0] WW4BEG[10] WW4BEG[11] WW4BEG[12] WW4BEG[13] WW4BEG[14] WW4BEG[15] WW4BEG[1]
+ WW4BEG[2] WW4BEG[3] WW4BEG[4] WW4BEG[5] WW4BEG[6] WW4BEG[7] WW4BEG[8] WW4BEG[9]
+ WW4END[0] WW4END[10] WW4END[11] WW4END[12] WW4END[13] WW4END[14] WW4END[15] WW4END[1]
+ WW4END[2] WW4END[3] WW4END[4] WW4END[5] WW4END[6] WW4END[7] WW4END[8] WW4END[9]
.ends

* Black-box entry subcircuit for W_TT_IF abstract view
.subckt W_TT_IF CLK_TT_PROJECT E1BEG[0] E1BEG[1] E1BEG[2] E1BEG[3] E2BEG[0] E2BEG[1]
+ E2BEG[2] E2BEG[3] E2BEG[4] E2BEG[5] E2BEG[6] E2BEG[7] E2BEGb[0] E2BEGb[1] E2BEGb[2]
+ E2BEGb[3] E2BEGb[4] E2BEGb[5] E2BEGb[6] E2BEGb[7] E6BEG[0] E6BEG[10] E6BEG[11] E6BEG[1]
+ E6BEG[2] E6BEG[3] E6BEG[4] E6BEG[5] E6BEG[6] E6BEG[7] E6BEG[8] E6BEG[9] EE4BEG[0]
+ EE4BEG[10] EE4BEG[11] EE4BEG[12] EE4BEG[13] EE4BEG[14] EE4BEG[15] EE4BEG[1] EE4BEG[2]
+ EE4BEG[3] EE4BEG[4] EE4BEG[5] EE4BEG[6] EE4BEG[7] EE4BEG[8] EE4BEG[9] ENA_TT_PROJECT
+ FrameData[0] FrameData[10] FrameData[11] FrameData[12] FrameData[13] FrameData[14]
+ FrameData[15] FrameData[16] FrameData[17] FrameData[18] FrameData[19] FrameData[1]
+ FrameData[20] FrameData[21] FrameData[22] FrameData[23] FrameData[24] FrameData[25]
+ FrameData[26] FrameData[27] FrameData[28] FrameData[29] FrameData[2] FrameData[30]
+ FrameData[31] FrameData[3] FrameData[4] FrameData[5] FrameData[6] FrameData[7] FrameData[8]
+ FrameData[9] FrameData_O[0] FrameData_O[10] FrameData_O[11] FrameData_O[12] FrameData_O[13]
+ FrameData_O[14] FrameData_O[15] FrameData_O[16] FrameData_O[17] FrameData_O[18]
+ FrameData_O[19] FrameData_O[1] FrameData_O[20] FrameData_O[21] FrameData_O[22] FrameData_O[23]
+ FrameData_O[24] FrameData_O[25] FrameData_O[26] FrameData_O[27] FrameData_O[28]
+ FrameData_O[29] FrameData_O[2] FrameData_O[30] FrameData_O[31] FrameData_O[3] FrameData_O[4]
+ FrameData_O[5] FrameData_O[6] FrameData_O[7] FrameData_O[8] FrameData_O[9] FrameStrobe[0]
+ FrameStrobe[10] FrameStrobe[11] FrameStrobe[12] FrameStrobe[13] FrameStrobe[14]
+ FrameStrobe[15] FrameStrobe[16] FrameStrobe[17] FrameStrobe[18] FrameStrobe[19]
+ FrameStrobe[1] FrameStrobe[2] FrameStrobe[3] FrameStrobe[4] FrameStrobe[5] FrameStrobe[6]
+ FrameStrobe[7] FrameStrobe[8] FrameStrobe[9] FrameStrobe_O[0] FrameStrobe_O[10]
+ FrameStrobe_O[11] FrameStrobe_O[12] FrameStrobe_O[13] FrameStrobe_O[14] FrameStrobe_O[15]
+ FrameStrobe_O[16] FrameStrobe_O[17] FrameStrobe_O[18] FrameStrobe_O[19] FrameStrobe_O[1]
+ FrameStrobe_O[2] FrameStrobe_O[3] FrameStrobe_O[4] FrameStrobe_O[5] FrameStrobe_O[6]
+ FrameStrobe_O[7] FrameStrobe_O[8] FrameStrobe_O[9] N1BEG[0] N1BEG[1] N1BEG[2] N1BEG[3]
+ N1END[0] N1END[1] N1END[2] N1END[3] N2BEG[0] N2BEG[1] N2BEG[2] N2BEG[3] N2BEG[4]
+ N2BEG[5] N2BEG[6] N2BEG[7] N2BEGb[0] N2BEGb[1] N2BEGb[2] N2BEGb[3] N2BEGb[4] N2BEGb[5]
+ N2BEGb[6] N2BEGb[7] N2END[0] N2END[1] N2END[2] N2END[3] N2END[4] N2END[5] N2END[6]
+ N2END[7] N2MID[0] N2MID[1] N2MID[2] N2MID[3] N2MID[4] N2MID[5] N2MID[6] N2MID[7]
+ N4BEG[0] N4BEG[10] N4BEG[11] N4BEG[12] N4BEG[13] N4BEG[14] N4BEG[15] N4BEG[1] N4BEG[2]
+ N4BEG[3] N4BEG[4] N4BEG[5] N4BEG[6] N4BEG[7] N4BEG[8] N4BEG[9] N4END[0] N4END[10]
+ N4END[11] N4END[12] N4END[13] N4END[14] N4END[15] N4END[1] N4END[2] N4END[3] N4END[4]
+ N4END[5] N4END[6] N4END[7] N4END[8] N4END[9] RST_N_TT_PROJECT S1BEG[0] S1BEG[1]
+ S1BEG[2] S1BEG[3] S1END[0] S1END[1] S1END[2] S1END[3] S2BEG[0] S2BEG[1] S2BEG[2]
+ S2BEG[3] S2BEG[4] S2BEG[5] S2BEG[6] S2BEG[7] S2BEGb[0] S2BEGb[1] S2BEGb[2] S2BEGb[3]
+ S2BEGb[4] S2BEGb[5] S2BEGb[6] S2BEGb[7] S2END[0] S2END[1] S2END[2] S2END[3] S2END[4]
+ S2END[5] S2END[6] S2END[7] S2MID[0] S2MID[1] S2MID[2] S2MID[3] S2MID[4] S2MID[5]
+ S2MID[6] S2MID[7] S4BEG[0] S4BEG[10] S4BEG[11] S4BEG[12] S4BEG[13] S4BEG[14] S4BEG[15]
+ S4BEG[1] S4BEG[2] S4BEG[3] S4BEG[4] S4BEG[5] S4BEG[6] S4BEG[7] S4BEG[8] S4BEG[9]
+ S4END[0] S4END[10] S4END[11] S4END[12] S4END[13] S4END[14] S4END[15] S4END[1] S4END[2]
+ S4END[3] S4END[4] S4END[5] S4END[6] S4END[7] S4END[8] S4END[9] UIO_IN_TT_PROJECT0
+ UIO_IN_TT_PROJECT1 UIO_IN_TT_PROJECT2 UIO_IN_TT_PROJECT3 UIO_IN_TT_PROJECT4 UIO_IN_TT_PROJECT5
+ UIO_IN_TT_PROJECT6 UIO_IN_TT_PROJECT7 UIO_OE_TT_PROJECT0 UIO_OE_TT_PROJECT1 UIO_OE_TT_PROJECT2
+ UIO_OE_TT_PROJECT3 UIO_OE_TT_PROJECT4 UIO_OE_TT_PROJECT5 UIO_OE_TT_PROJECT6 UIO_OE_TT_PROJECT7
+ UIO_OUT_TT_PROJECT0 UIO_OUT_TT_PROJECT1 UIO_OUT_TT_PROJECT2 UIO_OUT_TT_PROJECT3
+ UIO_OUT_TT_PROJECT4 UIO_OUT_TT_PROJECT5 UIO_OUT_TT_PROJECT6 UIO_OUT_TT_PROJECT7
+ UI_IN_TT_PROJECT0 UI_IN_TT_PROJECT1 UI_IN_TT_PROJECT2 UI_IN_TT_PROJECT3 UI_IN_TT_PROJECT4
+ UI_IN_TT_PROJECT5 UI_IN_TT_PROJECT6 UI_IN_TT_PROJECT7 UO_OUT_TT_PROJECT0 UO_OUT_TT_PROJECT1
+ UO_OUT_TT_PROJECT2 UO_OUT_TT_PROJECT3 UO_OUT_TT_PROJECT4 UO_OUT_TT_PROJECT5 UO_OUT_TT_PROJECT6
+ UO_OUT_TT_PROJECT7 UserCLK UserCLKo VGND VPWR W1END[0] W1END[1] W1END[2] W1END[3]
+ W2END[0] W2END[1] W2END[2] W2END[3] W2END[4] W2END[5] W2END[6] W2END[7] W2MID[0]
+ W2MID[1] W2MID[2] W2MID[3] W2MID[4] W2MID[5] W2MID[6] W2MID[7] W6END[0] W6END[10]
+ W6END[11] W6END[1] W6END[2] W6END[3] W6END[4] W6END[5] W6END[6] W6END[7] W6END[8]
+ W6END[9] WW4END[0] WW4END[10] WW4END[11] WW4END[12] WW4END[13] WW4END[14] WW4END[15]
+ WW4END[1] WW4END[2] WW4END[3] WW4END[4] WW4END[5] WW4END[6] WW4END[7] WW4END[8]
+ WW4END[9]
.ends

* Black-box entry subcircuit for SW_term abstract view
.subckt SW_term FrameData[0] FrameData[10] FrameData[11] FrameData[12] FrameData[13]
+ FrameData[14] FrameData[15] FrameData[16] FrameData[17] FrameData[18] FrameData[19]
+ FrameData[1] FrameData[20] FrameData[21] FrameData[22] FrameData[23] FrameData[24]
+ FrameData[25] FrameData[26] FrameData[27] FrameData[28] FrameData[29] FrameData[2]
+ FrameData[30] FrameData[31] FrameData[3] FrameData[4] FrameData[5] FrameData[6]
+ FrameData[7] FrameData[8] FrameData[9] FrameData_O[0] FrameData_O[10] FrameData_O[11]
+ FrameData_O[12] FrameData_O[13] FrameData_O[14] FrameData_O[15] FrameData_O[16]
+ FrameData_O[17] FrameData_O[18] FrameData_O[19] FrameData_O[1] FrameData_O[20] FrameData_O[21]
+ FrameData_O[22] FrameData_O[23] FrameData_O[24] FrameData_O[25] FrameData_O[26]
+ FrameData_O[27] FrameData_O[28] FrameData_O[29] FrameData_O[2] FrameData_O[30] FrameData_O[31]
+ FrameData_O[3] FrameData_O[4] FrameData_O[5] FrameData_O[6] FrameData_O[7] FrameData_O[8]
+ FrameData_O[9] FrameStrobe[0] FrameStrobe[10] FrameStrobe[11] FrameStrobe[12] FrameStrobe[13]
+ FrameStrobe[14] FrameStrobe[15] FrameStrobe[16] FrameStrobe[17] FrameStrobe[18]
+ FrameStrobe[19] FrameStrobe[1] FrameStrobe[2] FrameStrobe[3] FrameStrobe[4] FrameStrobe[5]
+ FrameStrobe[6] FrameStrobe[7] FrameStrobe[8] FrameStrobe[9] FrameStrobe_O[0] FrameStrobe_O[10]
+ FrameStrobe_O[11] FrameStrobe_O[12] FrameStrobe_O[13] FrameStrobe_O[14] FrameStrobe_O[15]
+ FrameStrobe_O[16] FrameStrobe_O[17] FrameStrobe_O[18] FrameStrobe_O[19] FrameStrobe_O[1]
+ FrameStrobe_O[2] FrameStrobe_O[3] FrameStrobe_O[4] FrameStrobe_O[5] FrameStrobe_O[6]
+ FrameStrobe_O[7] FrameStrobe_O[8] FrameStrobe_O[9] N1BEG[0] N1BEG[1] N1BEG[2] N1BEG[3]
+ N2BEG[0] N2BEG[1] N2BEG[2] N2BEG[3] N2BEG[4] N2BEG[5] N2BEG[6] N2BEG[7] N2BEGb[0]
+ N2BEGb[1] N2BEGb[2] N2BEGb[3] N2BEGb[4] N2BEGb[5] N2BEGb[6] N2BEGb[7] N4BEG[0] N4BEG[10]
+ N4BEG[11] N4BEG[12] N4BEG[13] N4BEG[14] N4BEG[15] N4BEG[1] N4BEG[2] N4BEG[3] N4BEG[4]
+ N4BEG[5] N4BEG[6] N4BEG[7] N4BEG[8] N4BEG[9] S1END[0] S1END[1] S1END[2] S1END[3]
+ S2END[0] S2END[1] S2END[2] S2END[3] S2END[4] S2END[5] S2END[6] S2END[7] S2MID[0]
+ S2MID[1] S2MID[2] S2MID[3] S2MID[4] S2MID[5] S2MID[6] S2MID[7] S4END[0] S4END[10]
+ S4END[11] S4END[12] S4END[13] S4END[14] S4END[15] S4END[1] S4END[2] S4END[3] S4END[4]
+ S4END[5] S4END[6] S4END[7] S4END[8] S4END[9] UserCLK UserCLKo VGND VPWR
.ends

* Black-box entry subcircuit for S_IO4 abstract view
.subckt S_IO4 A_I_top A_O_top A_T_top B_I_top B_O_top B_T_top C_I_top C_O_top C_T_top
+ Co D_I_top D_O_top D_T_top FrameData[0] FrameData[10] FrameData[11] FrameData[12]
+ FrameData[13] FrameData[14] FrameData[15] FrameData[16] FrameData[17] FrameData[18]
+ FrameData[19] FrameData[1] FrameData[20] FrameData[21] FrameData[22] FrameData[23]
+ FrameData[24] FrameData[25] FrameData[26] FrameData[27] FrameData[28] FrameData[29]
+ FrameData[2] FrameData[30] FrameData[31] FrameData[3] FrameData[4] FrameData[5]
+ FrameData[6] FrameData[7] FrameData[8] FrameData[9] FrameData_O[0] FrameData_O[10]
+ FrameData_O[11] FrameData_O[12] FrameData_O[13] FrameData_O[14] FrameData_O[15]
+ FrameData_O[16] FrameData_O[17] FrameData_O[18] FrameData_O[19] FrameData_O[1] FrameData_O[20]
+ FrameData_O[21] FrameData_O[22] FrameData_O[23] FrameData_O[24] FrameData_O[25]
+ FrameData_O[26] FrameData_O[27] FrameData_O[28] FrameData_O[29] FrameData_O[2] FrameData_O[30]
+ FrameData_O[31] FrameData_O[3] FrameData_O[4] FrameData_O[5] FrameData_O[6] FrameData_O[7]
+ FrameData_O[8] FrameData_O[9] FrameStrobe[0] FrameStrobe[10] FrameStrobe[11] FrameStrobe[12]
+ FrameStrobe[13] FrameStrobe[14] FrameStrobe[15] FrameStrobe[16] FrameStrobe[17]
+ FrameStrobe[18] FrameStrobe[19] FrameStrobe[1] FrameStrobe[2] FrameStrobe[3] FrameStrobe[4]
+ FrameStrobe[5] FrameStrobe[6] FrameStrobe[7] FrameStrobe[8] FrameStrobe[9] FrameStrobe_O[0]
+ FrameStrobe_O[10] FrameStrobe_O[11] FrameStrobe_O[12] FrameStrobe_O[13] FrameStrobe_O[14]
+ FrameStrobe_O[15] FrameStrobe_O[16] FrameStrobe_O[17] FrameStrobe_O[18] FrameStrobe_O[19]
+ FrameStrobe_O[1] FrameStrobe_O[2] FrameStrobe_O[3] FrameStrobe_O[4] FrameStrobe_O[5]
+ FrameStrobe_O[6] FrameStrobe_O[7] FrameStrobe_O[8] FrameStrobe_O[9] N1BEG[0] N1BEG[1]
+ N1BEG[2] N1BEG[3] N2BEG[0] N2BEG[1] N2BEG[2] N2BEG[3] N2BEG[4] N2BEG[5] N2BEG[6]
+ N2BEG[7] N2BEGb[0] N2BEGb[1] N2BEGb[2] N2BEGb[3] N2BEGb[4] N2BEGb[5] N2BEGb[6] N2BEGb[7]
+ N4BEG[0] N4BEG[10] N4BEG[11] N4BEG[12] N4BEG[13] N4BEG[14] N4BEG[15] N4BEG[1] N4BEG[2]
+ N4BEG[3] N4BEG[4] N4BEG[5] N4BEG[6] N4BEG[7] N4BEG[8] N4BEG[9] NN4BEG[0] NN4BEG[10]
+ NN4BEG[11] NN4BEG[12] NN4BEG[13] NN4BEG[14] NN4BEG[15] NN4BEG[1] NN4BEG[2] NN4BEG[3]
+ NN4BEG[4] NN4BEG[5] NN4BEG[6] NN4BEG[7] NN4BEG[8] NN4BEG[9] S1END[0] S1END[1] S1END[2]
+ S1END[3] S2END[0] S2END[1] S2END[2] S2END[3] S2END[4] S2END[5] S2END[6] S2END[7]
+ S2MID[0] S2MID[1] S2MID[2] S2MID[3] S2MID[4] S2MID[5] S2MID[6] S2MID[7] S4END[0]
+ S4END[10] S4END[11] S4END[12] S4END[13] S4END[14] S4END[15] S4END[1] S4END[2] S4END[3]
+ S4END[4] S4END[5] S4END[6] S4END[7] S4END[8] S4END[9] SS4END[0] SS4END[10] SS4END[11]
+ SS4END[12] SS4END[13] SS4END[14] SS4END[15] SS4END[1] SS4END[2] SS4END[3] SS4END[4]
+ SS4END[5] SS4END[6] SS4END[7] SS4END[8] SS4END[9] UserCLK UserCLKo VGND VPWR
.ends

* Black-box entry subcircuit for E_TT_IF abstract view
.subckt E_TT_IF CLK_TT_PROJECT E1END[0] E1END[1] E1END[2] E1END[3] E2END[0] E2END[1]
+ E2END[2] E2END[3] E2END[4] E2END[5] E2END[6] E2END[7] E2MID[0] E2MID[1] E2MID[2]
+ E2MID[3] E2MID[4] E2MID[5] E2MID[6] E2MID[7] E6END[0] E6END[10] E6END[11] E6END[1]
+ E6END[2] E6END[3] E6END[4] E6END[5] E6END[6] E6END[7] E6END[8] E6END[9] EE4END[0]
+ EE4END[10] EE4END[11] EE4END[12] EE4END[13] EE4END[14] EE4END[15] EE4END[1] EE4END[2]
+ EE4END[3] EE4END[4] EE4END[5] EE4END[6] EE4END[7] EE4END[8] EE4END[9] ENA_TT_PROJECT
+ FrameData[0] FrameData[10] FrameData[11] FrameData[12] FrameData[13] FrameData[14]
+ FrameData[15] FrameData[16] FrameData[17] FrameData[18] FrameData[19] FrameData[1]
+ FrameData[20] FrameData[21] FrameData[22] FrameData[23] FrameData[24] FrameData[25]
+ FrameData[26] FrameData[27] FrameData[28] FrameData[29] FrameData[2] FrameData[30]
+ FrameData[31] FrameData[3] FrameData[4] FrameData[5] FrameData[6] FrameData[7] FrameData[8]
+ FrameData[9] FrameData_O[0] FrameData_O[10] FrameData_O[11] FrameData_O[12] FrameData_O[13]
+ FrameData_O[14] FrameData_O[15] FrameData_O[16] FrameData_O[17] FrameData_O[18]
+ FrameData_O[19] FrameData_O[1] FrameData_O[20] FrameData_O[21] FrameData_O[22] FrameData_O[23]
+ FrameData_O[24] FrameData_O[25] FrameData_O[26] FrameData_O[27] FrameData_O[28]
+ FrameData_O[29] FrameData_O[2] FrameData_O[30] FrameData_O[31] FrameData_O[3] FrameData_O[4]
+ FrameData_O[5] FrameData_O[6] FrameData_O[7] FrameData_O[8] FrameData_O[9] FrameStrobe[0]
+ FrameStrobe[10] FrameStrobe[11] FrameStrobe[12] FrameStrobe[13] FrameStrobe[14]
+ FrameStrobe[15] FrameStrobe[16] FrameStrobe[17] FrameStrobe[18] FrameStrobe[19]
+ FrameStrobe[1] FrameStrobe[2] FrameStrobe[3] FrameStrobe[4] FrameStrobe[5] FrameStrobe[6]
+ FrameStrobe[7] FrameStrobe[8] FrameStrobe[9] FrameStrobe_O[0] FrameStrobe_O[10]
+ FrameStrobe_O[11] FrameStrobe_O[12] FrameStrobe_O[13] FrameStrobe_O[14] FrameStrobe_O[15]
+ FrameStrobe_O[16] FrameStrobe_O[17] FrameStrobe_O[18] FrameStrobe_O[19] FrameStrobe_O[1]
+ FrameStrobe_O[2] FrameStrobe_O[3] FrameStrobe_O[4] FrameStrobe_O[5] FrameStrobe_O[6]
+ FrameStrobe_O[7] FrameStrobe_O[8] FrameStrobe_O[9] N1BEG[0] N1BEG[1] N1BEG[2] N1BEG[3]
+ N1END[0] N1END[1] N1END[2] N1END[3] N2BEG[0] N2BEG[1] N2BEG[2] N2BEG[3] N2BEG[4]
+ N2BEG[5] N2BEG[6] N2BEG[7] N2BEGb[0] N2BEGb[1] N2BEGb[2] N2BEGb[3] N2BEGb[4] N2BEGb[5]
+ N2BEGb[6] N2BEGb[7] N2END[0] N2END[1] N2END[2] N2END[3] N2END[4] N2END[5] N2END[6]
+ N2END[7] N2MID[0] N2MID[1] N2MID[2] N2MID[3] N2MID[4] N2MID[5] N2MID[6] N2MID[7]
+ N4BEG[0] N4BEG[10] N4BEG[11] N4BEG[12] N4BEG[13] N4BEG[14] N4BEG[15] N4BEG[1] N4BEG[2]
+ N4BEG[3] N4BEG[4] N4BEG[5] N4BEG[6] N4BEG[7] N4BEG[8] N4BEG[9] N4END[0] N4END[10]
+ N4END[11] N4END[12] N4END[13] N4END[14] N4END[15] N4END[1] N4END[2] N4END[3] N4END[4]
+ N4END[5] N4END[6] N4END[7] N4END[8] N4END[9] RST_N_TT_PROJECT S1BEG[0] S1BEG[1]
+ S1BEG[2] S1BEG[3] S1END[0] S1END[1] S1END[2] S1END[3] S2BEG[0] S2BEG[1] S2BEG[2]
+ S2BEG[3] S2BEG[4] S2BEG[5] S2BEG[6] S2BEG[7] S2BEGb[0] S2BEGb[1] S2BEGb[2] S2BEGb[3]
+ S2BEGb[4] S2BEGb[5] S2BEGb[6] S2BEGb[7] S2END[0] S2END[1] S2END[2] S2END[3] S2END[4]
+ S2END[5] S2END[6] S2END[7] S2MID[0] S2MID[1] S2MID[2] S2MID[3] S2MID[4] S2MID[5]
+ S2MID[6] S2MID[7] S4BEG[0] S4BEG[10] S4BEG[11] S4BEG[12] S4BEG[13] S4BEG[14] S4BEG[15]
+ S4BEG[1] S4BEG[2] S4BEG[3] S4BEG[4] S4BEG[5] S4BEG[6] S4BEG[7] S4BEG[8] S4BEG[9]
+ S4END[0] S4END[10] S4END[11] S4END[12] S4END[13] S4END[14] S4END[15] S4END[1] S4END[2]
+ S4END[3] S4END[4] S4END[5] S4END[6] S4END[7] S4END[8] S4END[9] UIO_IN_TT_PROJECT0
+ UIO_IN_TT_PROJECT1 UIO_IN_TT_PROJECT2 UIO_IN_TT_PROJECT3 UIO_IN_TT_PROJECT4 UIO_IN_TT_PROJECT5
+ UIO_IN_TT_PROJECT6 UIO_IN_TT_PROJECT7 UIO_OE_TT_PROJECT0 UIO_OE_TT_PROJECT1 UIO_OE_TT_PROJECT2
+ UIO_OE_TT_PROJECT3 UIO_OE_TT_PROJECT4 UIO_OE_TT_PROJECT5 UIO_OE_TT_PROJECT6 UIO_OE_TT_PROJECT7
+ UIO_OUT_TT_PROJECT0 UIO_OUT_TT_PROJECT1 UIO_OUT_TT_PROJECT2 UIO_OUT_TT_PROJECT3
+ UIO_OUT_TT_PROJECT4 UIO_OUT_TT_PROJECT5 UIO_OUT_TT_PROJECT6 UIO_OUT_TT_PROJECT7
+ UI_IN_TT_PROJECT0 UI_IN_TT_PROJECT1 UI_IN_TT_PROJECT2 UI_IN_TT_PROJECT3 UI_IN_TT_PROJECT4
+ UI_IN_TT_PROJECT5 UI_IN_TT_PROJECT6 UI_IN_TT_PROJECT7 UO_OUT_TT_PROJECT0 UO_OUT_TT_PROJECT1
+ UO_OUT_TT_PROJECT2 UO_OUT_TT_PROJECT3 UO_OUT_TT_PROJECT4 UO_OUT_TT_PROJECT5 UO_OUT_TT_PROJECT6
+ UO_OUT_TT_PROJECT7 UserCLK UserCLKo VGND VPWR W1BEG[0] W1BEG[1] W1BEG[2] W1BEG[3]
+ W2BEG[0] W2BEG[1] W2BEG[2] W2BEG[3] W2BEG[4] W2BEG[5] W2BEG[6] W2BEG[7] W2BEGb[0]
+ W2BEGb[1] W2BEGb[2] W2BEGb[3] W2BEGb[4] W2BEGb[5] W2BEGb[6] W2BEGb[7] W6BEG[0] W6BEG[10]
+ W6BEG[11] W6BEG[1] W6BEG[2] W6BEG[3] W6BEG[4] W6BEG[5] W6BEG[6] W6BEG[7] W6BEG[8]
+ W6BEG[9] WW4BEG[0] WW4BEG[10] WW4BEG[11] WW4BEG[12] WW4BEG[13] WW4BEG[14] WW4BEG[15]
+ WW4BEG[1] WW4BEG[2] WW4BEG[3] WW4BEG[4] WW4BEG[5] WW4BEG[6] WW4BEG[7] WW4BEG[8]
+ WW4BEG[9]
.ends

* Black-box entry subcircuit for N_IO4 abstract view
.subckt N_IO4 A_I_top A_O_top A_T_top B_I_top B_O_top B_T_top C_I_top C_O_top C_T_top
+ Ci D_I_top D_O_top D_T_top FrameData[0] FrameData[10] FrameData[11] FrameData[12]
+ FrameData[13] FrameData[14] FrameData[15] FrameData[16] FrameData[17] FrameData[18]
+ FrameData[19] FrameData[1] FrameData[20] FrameData[21] FrameData[22] FrameData[23]
+ FrameData[24] FrameData[25] FrameData[26] FrameData[27] FrameData[28] FrameData[29]
+ FrameData[2] FrameData[30] FrameData[31] FrameData[3] FrameData[4] FrameData[5]
+ FrameData[6] FrameData[7] FrameData[8] FrameData[9] FrameData_O[0] FrameData_O[10]
+ FrameData_O[11] FrameData_O[12] FrameData_O[13] FrameData_O[14] FrameData_O[15]
+ FrameData_O[16] FrameData_O[17] FrameData_O[18] FrameData_O[19] FrameData_O[1] FrameData_O[20]
+ FrameData_O[21] FrameData_O[22] FrameData_O[23] FrameData_O[24] FrameData_O[25]
+ FrameData_O[26] FrameData_O[27] FrameData_O[28] FrameData_O[29] FrameData_O[2] FrameData_O[30]
+ FrameData_O[31] FrameData_O[3] FrameData_O[4] FrameData_O[5] FrameData_O[6] FrameData_O[7]
+ FrameData_O[8] FrameData_O[9] FrameStrobe[0] FrameStrobe[10] FrameStrobe[11] FrameStrobe[12]
+ FrameStrobe[13] FrameStrobe[14] FrameStrobe[15] FrameStrobe[16] FrameStrobe[17]
+ FrameStrobe[18] FrameStrobe[19] FrameStrobe[1] FrameStrobe[2] FrameStrobe[3] FrameStrobe[4]
+ FrameStrobe[5] FrameStrobe[6] FrameStrobe[7] FrameStrobe[8] FrameStrobe[9] FrameStrobe_O[0]
+ FrameStrobe_O[10] FrameStrobe_O[11] FrameStrobe_O[12] FrameStrobe_O[13] FrameStrobe_O[14]
+ FrameStrobe_O[15] FrameStrobe_O[16] FrameStrobe_O[17] FrameStrobe_O[18] FrameStrobe_O[19]
+ FrameStrobe_O[1] FrameStrobe_O[2] FrameStrobe_O[3] FrameStrobe_O[4] FrameStrobe_O[5]
+ FrameStrobe_O[6] FrameStrobe_O[7] FrameStrobe_O[8] FrameStrobe_O[9] N1END[0] N1END[1]
+ N1END[2] N1END[3] N2END[0] N2END[1] N2END[2] N2END[3] N2END[4] N2END[5] N2END[6]
+ N2END[7] N2MID[0] N2MID[1] N2MID[2] N2MID[3] N2MID[4] N2MID[5] N2MID[6] N2MID[7]
+ N4END[0] N4END[10] N4END[11] N4END[12] N4END[13] N4END[14] N4END[15] N4END[1] N4END[2]
+ N4END[3] N4END[4] N4END[5] N4END[6] N4END[7] N4END[8] N4END[9] NN4END[0] NN4END[10]
+ NN4END[11] NN4END[12] NN4END[13] NN4END[14] NN4END[15] NN4END[1] NN4END[2] NN4END[3]
+ NN4END[4] NN4END[5] NN4END[6] NN4END[7] NN4END[8] NN4END[9] S1BEG[0] S1BEG[1] S1BEG[2]
+ S1BEG[3] S2BEG[0] S2BEG[1] S2BEG[2] S2BEG[3] S2BEG[4] S2BEG[5] S2BEG[6] S2BEG[7]
+ S2BEGb[0] S2BEGb[1] S2BEGb[2] S2BEGb[3] S2BEGb[4] S2BEGb[5] S2BEGb[6] S2BEGb[7]
+ S4BEG[0] S4BEG[10] S4BEG[11] S4BEG[12] S4BEG[13] S4BEG[14] S4BEG[15] S4BEG[1] S4BEG[2]
+ S4BEG[3] S4BEG[4] S4BEG[5] S4BEG[6] S4BEG[7] S4BEG[8] S4BEG[9] SS4BEG[0] SS4BEG[10]
+ SS4BEG[11] SS4BEG[12] SS4BEG[13] SS4BEG[14] SS4BEG[15] SS4BEG[1] SS4BEG[2] SS4BEG[3]
+ SS4BEG[4] SS4BEG[5] SS4BEG[6] SS4BEG[7] SS4BEG[8] SS4BEG[9] UserCLK UserCLKo VGND
+ VPWR
.ends

* Black-box entry subcircuit for IHP_SRAM abstract view
.subckt IHP_SRAM ADDR_SRAM0 ADDR_SRAM1 ADDR_SRAM2 ADDR_SRAM3 ADDR_SRAM4 ADDR_SRAM5
+ ADDR_SRAM6 ADDR_SRAM7 ADDR_SRAM8 ADDR_SRAM9 BM_SRAM0 BM_SRAM1 BM_SRAM10 BM_SRAM11
+ BM_SRAM12 BM_SRAM13 BM_SRAM14 BM_SRAM15 BM_SRAM16 BM_SRAM17 BM_SRAM18 BM_SRAM19
+ BM_SRAM2 BM_SRAM20 BM_SRAM21 BM_SRAM22 BM_SRAM23 BM_SRAM24 BM_SRAM25 BM_SRAM26 BM_SRAM27
+ BM_SRAM28 BM_SRAM29 BM_SRAM3 BM_SRAM30 BM_SRAM31 BM_SRAM4 BM_SRAM5 BM_SRAM6 BM_SRAM7
+ BM_SRAM8 BM_SRAM9 CLK_SRAM CONFIGURED_top DIN_SRAM0 DIN_SRAM1 DIN_SRAM10 DIN_SRAM11
+ DIN_SRAM12 DIN_SRAM13 DIN_SRAM14 DIN_SRAM15 DIN_SRAM16 DIN_SRAM17 DIN_SRAM18 DIN_SRAM19
+ DIN_SRAM2 DIN_SRAM20 DIN_SRAM21 DIN_SRAM22 DIN_SRAM23 DIN_SRAM24 DIN_SRAM25 DIN_SRAM26
+ DIN_SRAM27 DIN_SRAM28 DIN_SRAM29 DIN_SRAM3 DIN_SRAM30 DIN_SRAM31 DIN_SRAM4 DIN_SRAM5
+ DIN_SRAM6 DIN_SRAM7 DIN_SRAM8 DIN_SRAM9 DOUT_SRAM0 DOUT_SRAM1 DOUT_SRAM10 DOUT_SRAM11
+ DOUT_SRAM12 DOUT_SRAM13 DOUT_SRAM14 DOUT_SRAM15 DOUT_SRAM16 DOUT_SRAM17 DOUT_SRAM18
+ DOUT_SRAM19 DOUT_SRAM2 DOUT_SRAM20 DOUT_SRAM21 DOUT_SRAM22 DOUT_SRAM23 DOUT_SRAM24
+ DOUT_SRAM25 DOUT_SRAM26 DOUT_SRAM27 DOUT_SRAM28 DOUT_SRAM29 DOUT_SRAM3 DOUT_SRAM30
+ DOUT_SRAM31 DOUT_SRAM4 DOUT_SRAM5 DOUT_SRAM6 DOUT_SRAM7 DOUT_SRAM8 DOUT_SRAM9 MEN_SRAM
+ REN_SRAM TIE_HIGH_SRAM TIE_LOW_SRAM Tile_X0Y0_E1END[0] Tile_X0Y0_E1END[1] Tile_X0Y0_E1END[2]
+ Tile_X0Y0_E1END[3] Tile_X0Y0_E2END[0] Tile_X0Y0_E2END[1] Tile_X0Y0_E2END[2] Tile_X0Y0_E2END[3]
+ Tile_X0Y0_E2END[4] Tile_X0Y0_E2END[5] Tile_X0Y0_E2END[6] Tile_X0Y0_E2END[7] Tile_X0Y0_E2MID[0]
+ Tile_X0Y0_E2MID[1] Tile_X0Y0_E2MID[2] Tile_X0Y0_E2MID[3] Tile_X0Y0_E2MID[4] Tile_X0Y0_E2MID[5]
+ Tile_X0Y0_E2MID[6] Tile_X0Y0_E2MID[7] Tile_X0Y0_E6END[0] Tile_X0Y0_E6END[10] Tile_X0Y0_E6END[11]
+ Tile_X0Y0_E6END[1] Tile_X0Y0_E6END[2] Tile_X0Y0_E6END[3] Tile_X0Y0_E6END[4] Tile_X0Y0_E6END[5]
+ Tile_X0Y0_E6END[6] Tile_X0Y0_E6END[7] Tile_X0Y0_E6END[8] Tile_X0Y0_E6END[9] Tile_X0Y0_EE4END[0]
+ Tile_X0Y0_EE4END[10] Tile_X0Y0_EE4END[11] Tile_X0Y0_EE4END[12] Tile_X0Y0_EE4END[13]
+ Tile_X0Y0_EE4END[14] Tile_X0Y0_EE4END[15] Tile_X0Y0_EE4END[1] Tile_X0Y0_EE4END[2]
+ Tile_X0Y0_EE4END[3] Tile_X0Y0_EE4END[4] Tile_X0Y0_EE4END[5] Tile_X0Y0_EE4END[6]
+ Tile_X0Y0_EE4END[7] Tile_X0Y0_EE4END[8] Tile_X0Y0_EE4END[9] Tile_X0Y0_FrameData[0]
+ Tile_X0Y0_FrameData[10] Tile_X0Y0_FrameData[11] Tile_X0Y0_FrameData[12] Tile_X0Y0_FrameData[13]
+ Tile_X0Y0_FrameData[14] Tile_X0Y0_FrameData[15] Tile_X0Y0_FrameData[16] Tile_X0Y0_FrameData[17]
+ Tile_X0Y0_FrameData[18] Tile_X0Y0_FrameData[19] Tile_X0Y0_FrameData[1] Tile_X0Y0_FrameData[20]
+ Tile_X0Y0_FrameData[21] Tile_X0Y0_FrameData[22] Tile_X0Y0_FrameData[23] Tile_X0Y0_FrameData[24]
+ Tile_X0Y0_FrameData[25] Tile_X0Y0_FrameData[26] Tile_X0Y0_FrameData[27] Tile_X0Y0_FrameData[28]
+ Tile_X0Y0_FrameData[29] Tile_X0Y0_FrameData[2] Tile_X0Y0_FrameData[30] Tile_X0Y0_FrameData[31]
+ Tile_X0Y0_FrameData[3] Tile_X0Y0_FrameData[4] Tile_X0Y0_FrameData[5] Tile_X0Y0_FrameData[6]
+ Tile_X0Y0_FrameData[7] Tile_X0Y0_FrameData[8] Tile_X0Y0_FrameData[9] Tile_X0Y0_FrameData_O[0]
+ Tile_X0Y0_FrameData_O[10] Tile_X0Y0_FrameData_O[11] Tile_X0Y0_FrameData_O[12] Tile_X0Y0_FrameData_O[13]
+ Tile_X0Y0_FrameData_O[14] Tile_X0Y0_FrameData_O[15] Tile_X0Y0_FrameData_O[16] Tile_X0Y0_FrameData_O[17]
+ Tile_X0Y0_FrameData_O[18] Tile_X0Y0_FrameData_O[19] Tile_X0Y0_FrameData_O[1] Tile_X0Y0_FrameData_O[20]
+ Tile_X0Y0_FrameData_O[21] Tile_X0Y0_FrameData_O[22] Tile_X0Y0_FrameData_O[23] Tile_X0Y0_FrameData_O[24]
+ Tile_X0Y0_FrameData_O[25] Tile_X0Y0_FrameData_O[26] Tile_X0Y0_FrameData_O[27] Tile_X0Y0_FrameData_O[28]
+ Tile_X0Y0_FrameData_O[29] Tile_X0Y0_FrameData_O[2] Tile_X0Y0_FrameData_O[30] Tile_X0Y0_FrameData_O[31]
+ Tile_X0Y0_FrameData_O[3] Tile_X0Y0_FrameData_O[4] Tile_X0Y0_FrameData_O[5] Tile_X0Y0_FrameData_O[6]
+ Tile_X0Y0_FrameData_O[7] Tile_X0Y0_FrameData_O[8] Tile_X0Y0_FrameData_O[9] Tile_X0Y0_FrameStrobe_O[0]
+ Tile_X0Y0_FrameStrobe_O[10] Tile_X0Y0_FrameStrobe_O[11] Tile_X0Y0_FrameStrobe_O[12]
+ Tile_X0Y0_FrameStrobe_O[13] Tile_X0Y0_FrameStrobe_O[14] Tile_X0Y0_FrameStrobe_O[15]
+ Tile_X0Y0_FrameStrobe_O[16] Tile_X0Y0_FrameStrobe_O[17] Tile_X0Y0_FrameStrobe_O[18]
+ Tile_X0Y0_FrameStrobe_O[19] Tile_X0Y0_FrameStrobe_O[1] Tile_X0Y0_FrameStrobe_O[2]
+ Tile_X0Y0_FrameStrobe_O[3] Tile_X0Y0_FrameStrobe_O[4] Tile_X0Y0_FrameStrobe_O[5]
+ Tile_X0Y0_FrameStrobe_O[6] Tile_X0Y0_FrameStrobe_O[7] Tile_X0Y0_FrameStrobe_O[8]
+ Tile_X0Y0_FrameStrobe_O[9] Tile_X0Y0_N1BEG[0] Tile_X0Y0_N1BEG[1] Tile_X0Y0_N1BEG[2]
+ Tile_X0Y0_N1BEG[3] Tile_X0Y0_N2BEG[0] Tile_X0Y0_N2BEG[1] Tile_X0Y0_N2BEG[2] Tile_X0Y0_N2BEG[3]
+ Tile_X0Y0_N2BEG[4] Tile_X0Y0_N2BEG[5] Tile_X0Y0_N2BEG[6] Tile_X0Y0_N2BEG[7] Tile_X0Y0_N2BEGb[0]
+ Tile_X0Y0_N2BEGb[1] Tile_X0Y0_N2BEGb[2] Tile_X0Y0_N2BEGb[3] Tile_X0Y0_N2BEGb[4]
+ Tile_X0Y0_N2BEGb[5] Tile_X0Y0_N2BEGb[6] Tile_X0Y0_N2BEGb[7] Tile_X0Y0_N4BEG[0] Tile_X0Y0_N4BEG[10]
+ Tile_X0Y0_N4BEG[11] Tile_X0Y0_N4BEG[12] Tile_X0Y0_N4BEG[13] Tile_X0Y0_N4BEG[14]
+ Tile_X0Y0_N4BEG[15] Tile_X0Y0_N4BEG[1] Tile_X0Y0_N4BEG[2] Tile_X0Y0_N4BEG[3] Tile_X0Y0_N4BEG[4]
+ Tile_X0Y0_N4BEG[5] Tile_X0Y0_N4BEG[6] Tile_X0Y0_N4BEG[7] Tile_X0Y0_N4BEG[8] Tile_X0Y0_N4BEG[9]
+ Tile_X0Y0_S1END[0] Tile_X0Y0_S1END[1] Tile_X0Y0_S1END[2] Tile_X0Y0_S1END[3] Tile_X0Y0_S2END[0]
+ Tile_X0Y0_S2END[1] Tile_X0Y0_S2END[2] Tile_X0Y0_S2END[3] Tile_X0Y0_S2END[4] Tile_X0Y0_S2END[5]
+ Tile_X0Y0_S2END[6] Tile_X0Y0_S2END[7] Tile_X0Y0_S2MID[0] Tile_X0Y0_S2MID[1] Tile_X0Y0_S2MID[2]
+ Tile_X0Y0_S2MID[3] Tile_X0Y0_S2MID[4] Tile_X0Y0_S2MID[5] Tile_X0Y0_S2MID[6] Tile_X0Y0_S2MID[7]
+ Tile_X0Y0_S4END[0] Tile_X0Y0_S4END[10] Tile_X0Y0_S4END[11] Tile_X0Y0_S4END[12] Tile_X0Y0_S4END[13]
+ Tile_X0Y0_S4END[14] Tile_X0Y0_S4END[15] Tile_X0Y0_S4END[1] Tile_X0Y0_S4END[2] Tile_X0Y0_S4END[3]
+ Tile_X0Y0_S4END[4] Tile_X0Y0_S4END[5] Tile_X0Y0_S4END[6] Tile_X0Y0_S4END[7] Tile_X0Y0_S4END[8]
+ Tile_X0Y0_S4END[9] Tile_X0Y0_UserCLKo Tile_X0Y0_W1BEG[0] Tile_X0Y0_W1BEG[1] Tile_X0Y0_W1BEG[2]
+ Tile_X0Y0_W1BEG[3] Tile_X0Y0_W2BEG[0] Tile_X0Y0_W2BEG[1] Tile_X0Y0_W2BEG[2] Tile_X0Y0_W2BEG[3]
+ Tile_X0Y0_W2BEG[4] Tile_X0Y0_W2BEG[5] Tile_X0Y0_W2BEG[6] Tile_X0Y0_W2BEG[7] Tile_X0Y0_W2BEGb[0]
+ Tile_X0Y0_W2BEGb[1] Tile_X0Y0_W2BEGb[2] Tile_X0Y0_W2BEGb[3] Tile_X0Y0_W2BEGb[4]
+ Tile_X0Y0_W2BEGb[5] Tile_X0Y0_W2BEGb[6] Tile_X0Y0_W2BEGb[7] Tile_X0Y0_W6BEG[0] Tile_X0Y0_W6BEG[10]
+ Tile_X0Y0_W6BEG[11] Tile_X0Y0_W6BEG[1] Tile_X0Y0_W6BEG[2] Tile_X0Y0_W6BEG[3] Tile_X0Y0_W6BEG[4]
+ Tile_X0Y0_W6BEG[5] Tile_X0Y0_W6BEG[6] Tile_X0Y0_W6BEG[7] Tile_X0Y0_W6BEG[8] Tile_X0Y0_W6BEG[9]
+ Tile_X0Y0_WW4BEG[0] Tile_X0Y0_WW4BEG[10] Tile_X0Y0_WW4BEG[11] Tile_X0Y0_WW4BEG[12]
+ Tile_X0Y0_WW4BEG[13] Tile_X0Y0_WW4BEG[14] Tile_X0Y0_WW4BEG[15] Tile_X0Y0_WW4BEG[1]
+ Tile_X0Y0_WW4BEG[2] Tile_X0Y0_WW4BEG[3] Tile_X0Y0_WW4BEG[4] Tile_X0Y0_WW4BEG[5]
+ Tile_X0Y0_WW4BEG[6] Tile_X0Y0_WW4BEG[7] Tile_X0Y0_WW4BEG[8] Tile_X0Y0_WW4BEG[9]
+ Tile_X0Y1_E1END[0] Tile_X0Y1_E1END[1] Tile_X0Y1_E1END[2] Tile_X0Y1_E1END[3] Tile_X0Y1_E2END[0]
+ Tile_X0Y1_E2END[1] Tile_X0Y1_E2END[2] Tile_X0Y1_E2END[3] Tile_X0Y1_E2END[4] Tile_X0Y1_E2END[5]
+ Tile_X0Y1_E2END[6] Tile_X0Y1_E2END[7] Tile_X0Y1_E2MID[0] Tile_X0Y1_E2MID[1] Tile_X0Y1_E2MID[2]
+ Tile_X0Y1_E2MID[3] Tile_X0Y1_E2MID[4] Tile_X0Y1_E2MID[5] Tile_X0Y1_E2MID[6] Tile_X0Y1_E2MID[7]
+ Tile_X0Y1_E6END[0] Tile_X0Y1_E6END[10] Tile_X0Y1_E6END[11] Tile_X0Y1_E6END[1] Tile_X0Y1_E6END[2]
+ Tile_X0Y1_E6END[3] Tile_X0Y1_E6END[4] Tile_X0Y1_E6END[5] Tile_X0Y1_E6END[6] Tile_X0Y1_E6END[7]
+ Tile_X0Y1_E6END[8] Tile_X0Y1_E6END[9] Tile_X0Y1_EE4END[0] Tile_X0Y1_EE4END[10] Tile_X0Y1_EE4END[11]
+ Tile_X0Y1_EE4END[12] Tile_X0Y1_EE4END[13] Tile_X0Y1_EE4END[14] Tile_X0Y1_EE4END[15]
+ Tile_X0Y1_EE4END[1] Tile_X0Y1_EE4END[2] Tile_X0Y1_EE4END[3] Tile_X0Y1_EE4END[4]
+ Tile_X0Y1_EE4END[5] Tile_X0Y1_EE4END[6] Tile_X0Y1_EE4END[7] Tile_X0Y1_EE4END[8]
+ Tile_X0Y1_EE4END[9] Tile_X0Y1_FrameData[0] Tile_X0Y1_FrameData[10] Tile_X0Y1_FrameData[11]
+ Tile_X0Y1_FrameData[12] Tile_X0Y1_FrameData[13] Tile_X0Y1_FrameData[14] Tile_X0Y1_FrameData[15]
+ Tile_X0Y1_FrameData[16] Tile_X0Y1_FrameData[17] Tile_X0Y1_FrameData[18] Tile_X0Y1_FrameData[19]
+ Tile_X0Y1_FrameData[1] Tile_X0Y1_FrameData[20] Tile_X0Y1_FrameData[21] Tile_X0Y1_FrameData[22]
+ Tile_X0Y1_FrameData[23] Tile_X0Y1_FrameData[24] Tile_X0Y1_FrameData[25] Tile_X0Y1_FrameData[26]
+ Tile_X0Y1_FrameData[27] Tile_X0Y1_FrameData[28] Tile_X0Y1_FrameData[29] Tile_X0Y1_FrameData[2]
+ Tile_X0Y1_FrameData[30] Tile_X0Y1_FrameData[31] Tile_X0Y1_FrameData[3] Tile_X0Y1_FrameData[4]
+ Tile_X0Y1_FrameData[5] Tile_X0Y1_FrameData[6] Tile_X0Y1_FrameData[7] Tile_X0Y1_FrameData[8]
+ Tile_X0Y1_FrameData[9] Tile_X0Y1_FrameData_O[0] Tile_X0Y1_FrameData_O[10] Tile_X0Y1_FrameData_O[11]
+ Tile_X0Y1_FrameData_O[12] Tile_X0Y1_FrameData_O[13] Tile_X0Y1_FrameData_O[14] Tile_X0Y1_FrameData_O[15]
+ Tile_X0Y1_FrameData_O[16] Tile_X0Y1_FrameData_O[17] Tile_X0Y1_FrameData_O[18] Tile_X0Y1_FrameData_O[19]
+ Tile_X0Y1_FrameData_O[1] Tile_X0Y1_FrameData_O[20] Tile_X0Y1_FrameData_O[21] Tile_X0Y1_FrameData_O[22]
+ Tile_X0Y1_FrameData_O[23] Tile_X0Y1_FrameData_O[24] Tile_X0Y1_FrameData_O[25] Tile_X0Y1_FrameData_O[26]
+ Tile_X0Y1_FrameData_O[27] Tile_X0Y1_FrameData_O[28] Tile_X0Y1_FrameData_O[29] Tile_X0Y1_FrameData_O[2]
+ Tile_X0Y1_FrameData_O[30] Tile_X0Y1_FrameData_O[31] Tile_X0Y1_FrameData_O[3] Tile_X0Y1_FrameData_O[4]
+ Tile_X0Y1_FrameData_O[5] Tile_X0Y1_FrameData_O[6] Tile_X0Y1_FrameData_O[7] Tile_X0Y1_FrameData_O[8]
+ Tile_X0Y1_FrameData_O[9] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_FrameStrobe[10] Tile_X0Y1_FrameStrobe[11]
+ Tile_X0Y1_FrameStrobe[12] Tile_X0Y1_FrameStrobe[13] Tile_X0Y1_FrameStrobe[14] Tile_X0Y1_FrameStrobe[15]
+ Tile_X0Y1_FrameStrobe[16] Tile_X0Y1_FrameStrobe[17] Tile_X0Y1_FrameStrobe[18] Tile_X0Y1_FrameStrobe[19]
+ Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_FrameStrobe[4]
+ Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_FrameStrobe[8]
+ Tile_X0Y1_FrameStrobe[9] Tile_X0Y1_N1END[0] Tile_X0Y1_N1END[1] Tile_X0Y1_N1END[2]
+ Tile_X0Y1_N1END[3] Tile_X0Y1_N2END[0] Tile_X0Y1_N2END[1] Tile_X0Y1_N2END[2] Tile_X0Y1_N2END[3]
+ Tile_X0Y1_N2END[4] Tile_X0Y1_N2END[5] Tile_X0Y1_N2END[6] Tile_X0Y1_N2END[7] Tile_X0Y1_N2MID[0]
+ Tile_X0Y1_N2MID[1] Tile_X0Y1_N2MID[2] Tile_X0Y1_N2MID[3] Tile_X0Y1_N2MID[4] Tile_X0Y1_N2MID[5]
+ Tile_X0Y1_N2MID[6] Tile_X0Y1_N2MID[7] Tile_X0Y1_N4END[0] Tile_X0Y1_N4END[10] Tile_X0Y1_N4END[11]
+ Tile_X0Y1_N4END[12] Tile_X0Y1_N4END[13] Tile_X0Y1_N4END[14] Tile_X0Y1_N4END[15]
+ Tile_X0Y1_N4END[1] Tile_X0Y1_N4END[2] Tile_X0Y1_N4END[3] Tile_X0Y1_N4END[4] Tile_X0Y1_N4END[5]
+ Tile_X0Y1_N4END[6] Tile_X0Y1_N4END[7] Tile_X0Y1_N4END[8] Tile_X0Y1_N4END[9] Tile_X0Y1_S1BEG[0]
+ Tile_X0Y1_S1BEG[1] Tile_X0Y1_S1BEG[2] Tile_X0Y1_S1BEG[3] Tile_X0Y1_S2BEG[0] Tile_X0Y1_S2BEG[1]
+ Tile_X0Y1_S2BEG[2] Tile_X0Y1_S2BEG[3] Tile_X0Y1_S2BEG[4] Tile_X0Y1_S2BEG[5] Tile_X0Y1_S2BEG[6]
+ Tile_X0Y1_S2BEG[7] Tile_X0Y1_S2BEGb[0] Tile_X0Y1_S2BEGb[1] Tile_X0Y1_S2BEGb[2] Tile_X0Y1_S2BEGb[3]
+ Tile_X0Y1_S2BEGb[4] Tile_X0Y1_S2BEGb[5] Tile_X0Y1_S2BEGb[6] Tile_X0Y1_S2BEGb[7]
+ Tile_X0Y1_S4BEG[0] Tile_X0Y1_S4BEG[10] Tile_X0Y1_S4BEG[11] Tile_X0Y1_S4BEG[12] Tile_X0Y1_S4BEG[13]
+ Tile_X0Y1_S4BEG[14] Tile_X0Y1_S4BEG[15] Tile_X0Y1_S4BEG[1] Tile_X0Y1_S4BEG[2] Tile_X0Y1_S4BEG[3]
+ Tile_X0Y1_S4BEG[4] Tile_X0Y1_S4BEG[5] Tile_X0Y1_S4BEG[6] Tile_X0Y1_S4BEG[7] Tile_X0Y1_S4BEG[8]
+ Tile_X0Y1_S4BEG[9] Tile_X0Y1_UserCLK Tile_X0Y1_W1BEG[0] Tile_X0Y1_W1BEG[1] Tile_X0Y1_W1BEG[2]
+ Tile_X0Y1_W1BEG[3] Tile_X0Y1_W2BEG[0] Tile_X0Y1_W2BEG[1] Tile_X0Y1_W2BEG[2] Tile_X0Y1_W2BEG[3]
+ Tile_X0Y1_W2BEG[4] Tile_X0Y1_W2BEG[5] Tile_X0Y1_W2BEG[6] Tile_X0Y1_W2BEG[7] Tile_X0Y1_W2BEGb[0]
+ Tile_X0Y1_W2BEGb[1] Tile_X0Y1_W2BEGb[2] Tile_X0Y1_W2BEGb[3] Tile_X0Y1_W2BEGb[4]
+ Tile_X0Y1_W2BEGb[5] Tile_X0Y1_W2BEGb[6] Tile_X0Y1_W2BEGb[7] Tile_X0Y1_W6BEG[0] Tile_X0Y1_W6BEG[10]
+ Tile_X0Y1_W6BEG[11] Tile_X0Y1_W6BEG[1] Tile_X0Y1_W6BEG[2] Tile_X0Y1_W6BEG[3] Tile_X0Y1_W6BEG[4]
+ Tile_X0Y1_W6BEG[5] Tile_X0Y1_W6BEG[6] Tile_X0Y1_W6BEG[7] Tile_X0Y1_W6BEG[8] Tile_X0Y1_W6BEG[9]
+ Tile_X0Y1_WW4BEG[0] Tile_X0Y1_WW4BEG[10] Tile_X0Y1_WW4BEG[11] Tile_X0Y1_WW4BEG[12]
+ Tile_X0Y1_WW4BEG[13] Tile_X0Y1_WW4BEG[14] Tile_X0Y1_WW4BEG[15] Tile_X0Y1_WW4BEG[1]
+ Tile_X0Y1_WW4BEG[2] Tile_X0Y1_WW4BEG[3] Tile_X0Y1_WW4BEG[4] Tile_X0Y1_WW4BEG[5]
+ Tile_X0Y1_WW4BEG[6] Tile_X0Y1_WW4BEG[7] Tile_X0Y1_WW4BEG[8] Tile_X0Y1_WW4BEG[9]
+ VGND VPWR WEN_SRAM
.ends

* Black-box entry subcircuit for SE_term abstract view
.subckt SE_term FrameData[0] FrameData[10] FrameData[11] FrameData[12] FrameData[13]
+ FrameData[14] FrameData[15] FrameData[16] FrameData[17] FrameData[18] FrameData[19]
+ FrameData[1] FrameData[20] FrameData[21] FrameData[22] FrameData[23] FrameData[24]
+ FrameData[25] FrameData[26] FrameData[27] FrameData[28] FrameData[29] FrameData[2]
+ FrameData[30] FrameData[31] FrameData[3] FrameData[4] FrameData[5] FrameData[6]
+ FrameData[7] FrameData[8] FrameData[9] FrameData_O[0] FrameData_O[10] FrameData_O[11]
+ FrameData_O[12] FrameData_O[13] FrameData_O[14] FrameData_O[15] FrameData_O[16]
+ FrameData_O[17] FrameData_O[18] FrameData_O[19] FrameData_O[1] FrameData_O[20] FrameData_O[21]
+ FrameData_O[22] FrameData_O[23] FrameData_O[24] FrameData_O[25] FrameData_O[26]
+ FrameData_O[27] FrameData_O[28] FrameData_O[29] FrameData_O[2] FrameData_O[30] FrameData_O[31]
+ FrameData_O[3] FrameData_O[4] FrameData_O[5] FrameData_O[6] FrameData_O[7] FrameData_O[8]
+ FrameData_O[9] FrameStrobe[0] FrameStrobe[10] FrameStrobe[11] FrameStrobe[12] FrameStrobe[13]
+ FrameStrobe[14] FrameStrobe[15] FrameStrobe[16] FrameStrobe[17] FrameStrobe[18]
+ FrameStrobe[19] FrameStrobe[1] FrameStrobe[2] FrameStrobe[3] FrameStrobe[4] FrameStrobe[5]
+ FrameStrobe[6] FrameStrobe[7] FrameStrobe[8] FrameStrobe[9] FrameStrobe_O[0] FrameStrobe_O[10]
+ FrameStrobe_O[11] FrameStrobe_O[12] FrameStrobe_O[13] FrameStrobe_O[14] FrameStrobe_O[15]
+ FrameStrobe_O[16] FrameStrobe_O[17] FrameStrobe_O[18] FrameStrobe_O[19] FrameStrobe_O[1]
+ FrameStrobe_O[2] FrameStrobe_O[3] FrameStrobe_O[4] FrameStrobe_O[5] FrameStrobe_O[6]
+ FrameStrobe_O[7] FrameStrobe_O[8] FrameStrobe_O[9] N1BEG[0] N1BEG[1] N1BEG[2] N1BEG[3]
+ N2BEG[0] N2BEG[1] N2BEG[2] N2BEG[3] N2BEG[4] N2BEG[5] N2BEG[6] N2BEG[7] N2BEGb[0]
+ N2BEGb[1] N2BEGb[2] N2BEGb[3] N2BEGb[4] N2BEGb[5] N2BEGb[6] N2BEGb[7] N4BEG[0] N4BEG[10]
+ N4BEG[11] N4BEG[12] N4BEG[13] N4BEG[14] N4BEG[15] N4BEG[1] N4BEG[2] N4BEG[3] N4BEG[4]
+ N4BEG[5] N4BEG[6] N4BEG[7] N4BEG[8] N4BEG[9] S1END[0] S1END[1] S1END[2] S1END[3]
+ S2END[0] S2END[1] S2END[2] S2END[3] S2END[4] S2END[5] S2END[6] S2END[7] S2MID[0]
+ S2MID[1] S2MID[2] S2MID[3] S2MID[4] S2MID[5] S2MID[6] S2MID[7] S4END[0] S4END[10]
+ S4END[11] S4END[12] S4END[13] S4END[14] S4END[15] S4END[1] S4END[2] S4END[3] S4END[4]
+ S4END[5] S4END[6] S4END[7] S4END[8] S4END[9] UserCLK UserCLKo VGND VPWR
.ends

* Black-box entry subcircuit for NW_term abstract view
.subckt NW_term FrameData[0] FrameData[10] FrameData[11] FrameData[12] FrameData[13]
+ FrameData[14] FrameData[15] FrameData[16] FrameData[17] FrameData[18] FrameData[19]
+ FrameData[1] FrameData[20] FrameData[21] FrameData[22] FrameData[23] FrameData[24]
+ FrameData[25] FrameData[26] FrameData[27] FrameData[28] FrameData[29] FrameData[2]
+ FrameData[30] FrameData[31] FrameData[3] FrameData[4] FrameData[5] FrameData[6]
+ FrameData[7] FrameData[8] FrameData[9] FrameData_O[0] FrameData_O[10] FrameData_O[11]
+ FrameData_O[12] FrameData_O[13] FrameData_O[14] FrameData_O[15] FrameData_O[16]
+ FrameData_O[17] FrameData_O[18] FrameData_O[19] FrameData_O[1] FrameData_O[20] FrameData_O[21]
+ FrameData_O[22] FrameData_O[23] FrameData_O[24] FrameData_O[25] FrameData_O[26]
+ FrameData_O[27] FrameData_O[28] FrameData_O[29] FrameData_O[2] FrameData_O[30] FrameData_O[31]
+ FrameData_O[3] FrameData_O[4] FrameData_O[5] FrameData_O[6] FrameData_O[7] FrameData_O[8]
+ FrameData_O[9] FrameStrobe[0] FrameStrobe[10] FrameStrobe[11] FrameStrobe[12] FrameStrobe[13]
+ FrameStrobe[14] FrameStrobe[15] FrameStrobe[16] FrameStrobe[17] FrameStrobe[18]
+ FrameStrobe[19] FrameStrobe[1] FrameStrobe[2] FrameStrobe[3] FrameStrobe[4] FrameStrobe[5]
+ FrameStrobe[6] FrameStrobe[7] FrameStrobe[8] FrameStrobe[9] FrameStrobe_O[0] FrameStrobe_O[10]
+ FrameStrobe_O[11] FrameStrobe_O[12] FrameStrobe_O[13] FrameStrobe_O[14] FrameStrobe_O[15]
+ FrameStrobe_O[16] FrameStrobe_O[17] FrameStrobe_O[18] FrameStrobe_O[19] FrameStrobe_O[1]
+ FrameStrobe_O[2] FrameStrobe_O[3] FrameStrobe_O[4] FrameStrobe_O[5] FrameStrobe_O[6]
+ FrameStrobe_O[7] FrameStrobe_O[8] FrameStrobe_O[9] N1END[0] N1END[1] N1END[2] N1END[3]
+ N2END[0] N2END[1] N2END[2] N2END[3] N2END[4] N2END[5] N2END[6] N2END[7] N2MID[0]
+ N2MID[1] N2MID[2] N2MID[3] N2MID[4] N2MID[5] N2MID[6] N2MID[7] N4END[0] N4END[10]
+ N4END[11] N4END[12] N4END[13] N4END[14] N4END[15] N4END[1] N4END[2] N4END[3] N4END[4]
+ N4END[5] N4END[6] N4END[7] N4END[8] N4END[9] S1BEG[0] S1BEG[1] S1BEG[2] S1BEG[3]
+ S2BEG[0] S2BEG[1] S2BEG[2] S2BEG[3] S2BEG[4] S2BEG[5] S2BEG[6] S2BEG[7] S2BEGb[0]
+ S2BEGb[1] S2BEGb[2] S2BEGb[3] S2BEGb[4] S2BEGb[5] S2BEGb[6] S2BEGb[7] S4BEG[0] S4BEG[10]
+ S4BEG[11] S4BEG[12] S4BEG[13] S4BEG[14] S4BEG[15] S4BEG[1] S4BEG[2] S4BEG[3] S4BEG[4]
+ S4BEG[5] S4BEG[6] S4BEG[7] S4BEG[8] S4BEG[9] UserCLK UserCLKo VGND VPWR
.ends

* Black-box entry subcircuit for NE_term abstract view
.subckt NE_term FrameData[0] FrameData[10] FrameData[11] FrameData[12] FrameData[13]
+ FrameData[14] FrameData[15] FrameData[16] FrameData[17] FrameData[18] FrameData[19]
+ FrameData[1] FrameData[20] FrameData[21] FrameData[22] FrameData[23] FrameData[24]
+ FrameData[25] FrameData[26] FrameData[27] FrameData[28] FrameData[29] FrameData[2]
+ FrameData[30] FrameData[31] FrameData[3] FrameData[4] FrameData[5] FrameData[6]
+ FrameData[7] FrameData[8] FrameData[9] FrameData_O[0] FrameData_O[10] FrameData_O[11]
+ FrameData_O[12] FrameData_O[13] FrameData_O[14] FrameData_O[15] FrameData_O[16]
+ FrameData_O[17] FrameData_O[18] FrameData_O[19] FrameData_O[1] FrameData_O[20] FrameData_O[21]
+ FrameData_O[22] FrameData_O[23] FrameData_O[24] FrameData_O[25] FrameData_O[26]
+ FrameData_O[27] FrameData_O[28] FrameData_O[29] FrameData_O[2] FrameData_O[30] FrameData_O[31]
+ FrameData_O[3] FrameData_O[4] FrameData_O[5] FrameData_O[6] FrameData_O[7] FrameData_O[8]
+ FrameData_O[9] FrameStrobe[0] FrameStrobe[10] FrameStrobe[11] FrameStrobe[12] FrameStrobe[13]
+ FrameStrobe[14] FrameStrobe[15] FrameStrobe[16] FrameStrobe[17] FrameStrobe[18]
+ FrameStrobe[19] FrameStrobe[1] FrameStrobe[2] FrameStrobe[3] FrameStrobe[4] FrameStrobe[5]
+ FrameStrobe[6] FrameStrobe[7] FrameStrobe[8] FrameStrobe[9] FrameStrobe_O[0] FrameStrobe_O[10]
+ FrameStrobe_O[11] FrameStrobe_O[12] FrameStrobe_O[13] FrameStrobe_O[14] FrameStrobe_O[15]
+ FrameStrobe_O[16] FrameStrobe_O[17] FrameStrobe_O[18] FrameStrobe_O[19] FrameStrobe_O[1]
+ FrameStrobe_O[2] FrameStrobe_O[3] FrameStrobe_O[4] FrameStrobe_O[5] FrameStrobe_O[6]
+ FrameStrobe_O[7] FrameStrobe_O[8] FrameStrobe_O[9] N1END[0] N1END[1] N1END[2] N1END[3]
+ N2END[0] N2END[1] N2END[2] N2END[3] N2END[4] N2END[5] N2END[6] N2END[7] N2MID[0]
+ N2MID[1] N2MID[2] N2MID[3] N2MID[4] N2MID[5] N2MID[6] N2MID[7] N4END[0] N4END[10]
+ N4END[11] N4END[12] N4END[13] N4END[14] N4END[15] N4END[1] N4END[2] N4END[3] N4END[4]
+ N4END[5] N4END[6] N4END[7] N4END[8] N4END[9] S1BEG[0] S1BEG[1] S1BEG[2] S1BEG[3]
+ S2BEG[0] S2BEG[1] S2BEG[2] S2BEG[3] S2BEG[4] S2BEG[5] S2BEG[6] S2BEG[7] S2BEGb[0]
+ S2BEGb[1] S2BEGb[2] S2BEGb[3] S2BEGb[4] S2BEGb[5] S2BEGb[6] S2BEGb[7] S4BEG[0] S4BEG[10]
+ S4BEG[11] S4BEG[12] S4BEG[13] S4BEG[14] S4BEG[15] S4BEG[1] S4BEG[2] S4BEG[3] S4BEG[4]
+ S4BEG[5] S4BEG[6] S4BEG[7] S4BEG[8] S4BEG[9] UserCLK UserCLKo VGND VPWR
.ends

.subckt eFPGA FrameData[0] FrameData[100] FrameData[101] FrameData[102] FrameData[103]
+ FrameData[104] FrameData[105] FrameData[106] FrameData[107] FrameData[108] FrameData[109]
+ FrameData[10] FrameData[110] FrameData[111] FrameData[112] FrameData[113] FrameData[114]
+ FrameData[115] FrameData[116] FrameData[117] FrameData[118] FrameData[119] FrameData[11]
+ FrameData[120] FrameData[121] FrameData[122] FrameData[123] FrameData[124] FrameData[125]
+ FrameData[126] FrameData[127] FrameData[128] FrameData[129] FrameData[12] FrameData[130]
+ FrameData[131] FrameData[132] FrameData[133] FrameData[134] FrameData[135] FrameData[136]
+ FrameData[137] FrameData[138] FrameData[139] FrameData[13] FrameData[140] FrameData[141]
+ FrameData[142] FrameData[143] FrameData[144] FrameData[145] FrameData[146] FrameData[147]
+ FrameData[148] FrameData[149] FrameData[14] FrameData[150] FrameData[151] FrameData[152]
+ FrameData[153] FrameData[154] FrameData[155] FrameData[156] FrameData[157] FrameData[158]
+ FrameData[159] FrameData[15] FrameData[160] FrameData[161] FrameData[162] FrameData[163]
+ FrameData[164] FrameData[165] FrameData[166] FrameData[167] FrameData[168] FrameData[169]
+ FrameData[16] FrameData[170] FrameData[171] FrameData[172] FrameData[173] FrameData[174]
+ FrameData[175] FrameData[176] FrameData[177] FrameData[178] FrameData[179] FrameData[17]
+ FrameData[180] FrameData[181] FrameData[182] FrameData[183] FrameData[184] FrameData[185]
+ FrameData[186] FrameData[187] FrameData[188] FrameData[189] FrameData[18] FrameData[190]
+ FrameData[191] FrameData[192] FrameData[193] FrameData[194] FrameData[195] FrameData[196]
+ FrameData[197] FrameData[198] FrameData[199] FrameData[19] FrameData[1] FrameData[200]
+ FrameData[201] FrameData[202] FrameData[203] FrameData[204] FrameData[205] FrameData[206]
+ FrameData[207] FrameData[208] FrameData[209] FrameData[20] FrameData[210] FrameData[211]
+ FrameData[212] FrameData[213] FrameData[214] FrameData[215] FrameData[216] FrameData[217]
+ FrameData[218] FrameData[219] FrameData[21] FrameData[220] FrameData[221] FrameData[222]
+ FrameData[223] FrameData[224] FrameData[225] FrameData[226] FrameData[227] FrameData[228]
+ FrameData[229] FrameData[22] FrameData[230] FrameData[231] FrameData[232] FrameData[233]
+ FrameData[234] FrameData[235] FrameData[236] FrameData[237] FrameData[238] FrameData[239]
+ FrameData[23] FrameData[240] FrameData[241] FrameData[242] FrameData[243] FrameData[244]
+ FrameData[245] FrameData[246] FrameData[247] FrameData[248] FrameData[249] FrameData[24]
+ FrameData[250] FrameData[251] FrameData[252] FrameData[253] FrameData[254] FrameData[255]
+ FrameData[256] FrameData[257] FrameData[258] FrameData[259] FrameData[25] FrameData[260]
+ FrameData[261] FrameData[262] FrameData[263] FrameData[264] FrameData[265] FrameData[266]
+ FrameData[267] FrameData[268] FrameData[269] FrameData[26] FrameData[270] FrameData[271]
+ FrameData[272] FrameData[273] FrameData[274] FrameData[275] FrameData[276] FrameData[277]
+ FrameData[278] FrameData[279] FrameData[27] FrameData[280] FrameData[281] FrameData[282]
+ FrameData[283] FrameData[284] FrameData[285] FrameData[286] FrameData[287] FrameData[288]
+ FrameData[289] FrameData[28] FrameData[290] FrameData[291] FrameData[292] FrameData[293]
+ FrameData[294] FrameData[295] FrameData[296] FrameData[297] FrameData[298] FrameData[299]
+ FrameData[29] FrameData[2] FrameData[300] FrameData[301] FrameData[302] FrameData[303]
+ FrameData[304] FrameData[305] FrameData[306] FrameData[307] FrameData[308] FrameData[309]
+ FrameData[30] FrameData[310] FrameData[311] FrameData[312] FrameData[313] FrameData[314]
+ FrameData[315] FrameData[316] FrameData[317] FrameData[318] FrameData[319] FrameData[31]
+ FrameData[32] FrameData[33] FrameData[34] FrameData[35] FrameData[36] FrameData[37]
+ FrameData[38] FrameData[39] FrameData[3] FrameData[40] FrameData[41] FrameData[42]
+ FrameData[43] FrameData[44] FrameData[45] FrameData[46] FrameData[47] FrameData[48]
+ FrameData[49] FrameData[4] FrameData[50] FrameData[51] FrameData[52] FrameData[53]
+ FrameData[54] FrameData[55] FrameData[56] FrameData[57] FrameData[58] FrameData[59]
+ FrameData[5] FrameData[60] FrameData[61] FrameData[62] FrameData[63] FrameData[64]
+ FrameData[65] FrameData[66] FrameData[67] FrameData[68] FrameData[69] FrameData[6]
+ FrameData[70] FrameData[71] FrameData[72] FrameData[73] FrameData[74] FrameData[75]
+ FrameData[76] FrameData[77] FrameData[78] FrameData[79] FrameData[7] FrameData[80]
+ FrameData[81] FrameData[82] FrameData[83] FrameData[84] FrameData[85] FrameData[86]
+ FrameData[87] FrameData[88] FrameData[89] FrameData[8] FrameData[90] FrameData[91]
+ FrameData[92] FrameData[93] FrameData[94] FrameData[95] FrameData[96] FrameData[97]
+ FrameData[98] FrameData[99] FrameData[9] FrameStrobe[0] FrameStrobe[100] FrameStrobe[101]
+ FrameStrobe[102] FrameStrobe[103] FrameStrobe[104] FrameStrobe[105] FrameStrobe[106]
+ FrameStrobe[107] FrameStrobe[108] FrameStrobe[109] FrameStrobe[10] FrameStrobe[110]
+ FrameStrobe[111] FrameStrobe[112] FrameStrobe[113] FrameStrobe[114] FrameStrobe[115]
+ FrameStrobe[116] FrameStrobe[117] FrameStrobe[118] FrameStrobe[119] FrameStrobe[11]
+ FrameStrobe[12] FrameStrobe[13] FrameStrobe[14] FrameStrobe[15] FrameStrobe[16]
+ FrameStrobe[17] FrameStrobe[18] FrameStrobe[19] FrameStrobe[1] FrameStrobe[20] FrameStrobe[21]
+ FrameStrobe[22] FrameStrobe[23] FrameStrobe[24] FrameStrobe[25] FrameStrobe[26]
+ FrameStrobe[27] FrameStrobe[28] FrameStrobe[29] FrameStrobe[2] FrameStrobe[30] FrameStrobe[31]
+ FrameStrobe[32] FrameStrobe[33] FrameStrobe[34] FrameStrobe[35] FrameStrobe[36]
+ FrameStrobe[37] FrameStrobe[38] FrameStrobe[39] FrameStrobe[3] FrameStrobe[40] FrameStrobe[41]
+ FrameStrobe[42] FrameStrobe[43] FrameStrobe[44] FrameStrobe[45] FrameStrobe[46]
+ FrameStrobe[47] FrameStrobe[48] FrameStrobe[49] FrameStrobe[4] FrameStrobe[50] FrameStrobe[51]
+ FrameStrobe[52] FrameStrobe[53] FrameStrobe[54] FrameStrobe[55] FrameStrobe[56]
+ FrameStrobe[57] FrameStrobe[58] FrameStrobe[59] FrameStrobe[5] FrameStrobe[60] FrameStrobe[61]
+ FrameStrobe[62] FrameStrobe[63] FrameStrobe[64] FrameStrobe[65] FrameStrobe[66]
+ FrameStrobe[67] FrameStrobe[68] FrameStrobe[69] FrameStrobe[6] FrameStrobe[70] FrameStrobe[71]
+ FrameStrobe[72] FrameStrobe[73] FrameStrobe[74] FrameStrobe[75] FrameStrobe[76]
+ FrameStrobe[77] FrameStrobe[78] FrameStrobe[79] FrameStrobe[7] FrameStrobe[80] FrameStrobe[81]
+ FrameStrobe[82] FrameStrobe[83] FrameStrobe[84] FrameStrobe[85] FrameStrobe[86]
+ FrameStrobe[87] FrameStrobe[88] FrameStrobe[89] FrameStrobe[8] FrameStrobe[90] FrameStrobe[91]
+ FrameStrobe[92] FrameStrobe[93] FrameStrobe[94] FrameStrobe[95] FrameStrobe[96]
+ FrameStrobe[97] FrameStrobe[98] FrameStrobe[99] FrameStrobe[9] Tile_X0Y1_CLK_TT_PROJECT
+ Tile_X0Y1_ENA_TT_PROJECT Tile_X0Y1_RST_N_TT_PROJECT Tile_X0Y1_UIO_IN_TT_PROJECT0
+ Tile_X0Y1_UIO_IN_TT_PROJECT1 Tile_X0Y1_UIO_IN_TT_PROJECT2 Tile_X0Y1_UIO_IN_TT_PROJECT3
+ Tile_X0Y1_UIO_IN_TT_PROJECT4 Tile_X0Y1_UIO_IN_TT_PROJECT5 Tile_X0Y1_UIO_IN_TT_PROJECT6
+ Tile_X0Y1_UIO_IN_TT_PROJECT7 Tile_X0Y1_UIO_OE_TT_PROJECT0 Tile_X0Y1_UIO_OE_TT_PROJECT1
+ Tile_X0Y1_UIO_OE_TT_PROJECT2 Tile_X0Y1_UIO_OE_TT_PROJECT3 Tile_X0Y1_UIO_OE_TT_PROJECT4
+ Tile_X0Y1_UIO_OE_TT_PROJECT5 Tile_X0Y1_UIO_OE_TT_PROJECT6 Tile_X0Y1_UIO_OE_TT_PROJECT7
+ Tile_X0Y1_UIO_OUT_TT_PROJECT0 Tile_X0Y1_UIO_OUT_TT_PROJECT1 Tile_X0Y1_UIO_OUT_TT_PROJECT2
+ Tile_X0Y1_UIO_OUT_TT_PROJECT3 Tile_X0Y1_UIO_OUT_TT_PROJECT4 Tile_X0Y1_UIO_OUT_TT_PROJECT5
+ Tile_X0Y1_UIO_OUT_TT_PROJECT6 Tile_X0Y1_UIO_OUT_TT_PROJECT7 Tile_X0Y1_UI_IN_TT_PROJECT0
+ Tile_X0Y1_UI_IN_TT_PROJECT1 Tile_X0Y1_UI_IN_TT_PROJECT2 Tile_X0Y1_UI_IN_TT_PROJECT3
+ Tile_X0Y1_UI_IN_TT_PROJECT4 Tile_X0Y1_UI_IN_TT_PROJECT5 Tile_X0Y1_UI_IN_TT_PROJECT6
+ Tile_X0Y1_UI_IN_TT_PROJECT7 Tile_X0Y1_UO_OUT_TT_PROJECT0 Tile_X0Y1_UO_OUT_TT_PROJECT1
+ Tile_X0Y1_UO_OUT_TT_PROJECT2 Tile_X0Y1_UO_OUT_TT_PROJECT3 Tile_X0Y1_UO_OUT_TT_PROJECT4
+ Tile_X0Y1_UO_OUT_TT_PROJECT5 Tile_X0Y1_UO_OUT_TT_PROJECT6 Tile_X0Y1_UO_OUT_TT_PROJECT7
+ Tile_X0Y2_CLK_TT_PROJECT Tile_X0Y2_ENA_TT_PROJECT Tile_X0Y2_RST_N_TT_PROJECT Tile_X0Y2_UIO_IN_TT_PROJECT0
+ Tile_X0Y2_UIO_IN_TT_PROJECT1 Tile_X0Y2_UIO_IN_TT_PROJECT2 Tile_X0Y2_UIO_IN_TT_PROJECT3
+ Tile_X0Y2_UIO_IN_TT_PROJECT4 Tile_X0Y2_UIO_IN_TT_PROJECT5 Tile_X0Y2_UIO_IN_TT_PROJECT6
+ Tile_X0Y2_UIO_IN_TT_PROJECT7 Tile_X0Y2_UIO_OE_TT_PROJECT0 Tile_X0Y2_UIO_OE_TT_PROJECT1
+ Tile_X0Y2_UIO_OE_TT_PROJECT2 Tile_X0Y2_UIO_OE_TT_PROJECT3 Tile_X0Y2_UIO_OE_TT_PROJECT4
+ Tile_X0Y2_UIO_OE_TT_PROJECT5 Tile_X0Y2_UIO_OE_TT_PROJECT6 Tile_X0Y2_UIO_OE_TT_PROJECT7
+ Tile_X0Y2_UIO_OUT_TT_PROJECT0 Tile_X0Y2_UIO_OUT_TT_PROJECT1 Tile_X0Y2_UIO_OUT_TT_PROJECT2
+ Tile_X0Y2_UIO_OUT_TT_PROJECT3 Tile_X0Y2_UIO_OUT_TT_PROJECT4 Tile_X0Y2_UIO_OUT_TT_PROJECT5
+ Tile_X0Y2_UIO_OUT_TT_PROJECT6 Tile_X0Y2_UIO_OUT_TT_PROJECT7 Tile_X0Y2_UI_IN_TT_PROJECT0
+ Tile_X0Y2_UI_IN_TT_PROJECT1 Tile_X0Y2_UI_IN_TT_PROJECT2 Tile_X0Y2_UI_IN_TT_PROJECT3
+ Tile_X0Y2_UI_IN_TT_PROJECT4 Tile_X0Y2_UI_IN_TT_PROJECT5 Tile_X0Y2_UI_IN_TT_PROJECT6
+ Tile_X0Y2_UI_IN_TT_PROJECT7 Tile_X0Y2_UO_OUT_TT_PROJECT0 Tile_X0Y2_UO_OUT_TT_PROJECT1
+ Tile_X0Y2_UO_OUT_TT_PROJECT2 Tile_X0Y2_UO_OUT_TT_PROJECT3 Tile_X0Y2_UO_OUT_TT_PROJECT4
+ Tile_X0Y2_UO_OUT_TT_PROJECT5 Tile_X0Y2_UO_OUT_TT_PROJECT6 Tile_X0Y2_UO_OUT_TT_PROJECT7
+ Tile_X0Y3_CLK_TT_PROJECT Tile_X0Y3_ENA_TT_PROJECT Tile_X0Y3_RST_N_TT_PROJECT Tile_X0Y3_UIO_IN_TT_PROJECT0
+ Tile_X0Y3_UIO_IN_TT_PROJECT1 Tile_X0Y3_UIO_IN_TT_PROJECT2 Tile_X0Y3_UIO_IN_TT_PROJECT3
+ Tile_X0Y3_UIO_IN_TT_PROJECT4 Tile_X0Y3_UIO_IN_TT_PROJECT5 Tile_X0Y3_UIO_IN_TT_PROJECT6
+ Tile_X0Y3_UIO_IN_TT_PROJECT7 Tile_X0Y3_UIO_OE_TT_PROJECT0 Tile_X0Y3_UIO_OE_TT_PROJECT1
+ Tile_X0Y3_UIO_OE_TT_PROJECT2 Tile_X0Y3_UIO_OE_TT_PROJECT3 Tile_X0Y3_UIO_OE_TT_PROJECT4
+ Tile_X0Y3_UIO_OE_TT_PROJECT5 Tile_X0Y3_UIO_OE_TT_PROJECT6 Tile_X0Y3_UIO_OE_TT_PROJECT7
+ Tile_X0Y3_UIO_OUT_TT_PROJECT0 Tile_X0Y3_UIO_OUT_TT_PROJECT1 Tile_X0Y3_UIO_OUT_TT_PROJECT2
+ Tile_X0Y3_UIO_OUT_TT_PROJECT3 Tile_X0Y3_UIO_OUT_TT_PROJECT4 Tile_X0Y3_UIO_OUT_TT_PROJECT5
+ Tile_X0Y3_UIO_OUT_TT_PROJECT6 Tile_X0Y3_UIO_OUT_TT_PROJECT7 Tile_X0Y3_UI_IN_TT_PROJECT0
+ Tile_X0Y3_UI_IN_TT_PROJECT1 Tile_X0Y3_UI_IN_TT_PROJECT2 Tile_X0Y3_UI_IN_TT_PROJECT3
+ Tile_X0Y3_UI_IN_TT_PROJECT4 Tile_X0Y3_UI_IN_TT_PROJECT5 Tile_X0Y3_UI_IN_TT_PROJECT6
+ Tile_X0Y3_UI_IN_TT_PROJECT7 Tile_X0Y3_UO_OUT_TT_PROJECT0 Tile_X0Y3_UO_OUT_TT_PROJECT1
+ Tile_X0Y3_UO_OUT_TT_PROJECT2 Tile_X0Y3_UO_OUT_TT_PROJECT3 Tile_X0Y3_UO_OUT_TT_PROJECT4
+ Tile_X0Y3_UO_OUT_TT_PROJECT5 Tile_X0Y3_UO_OUT_TT_PROJECT6 Tile_X0Y3_UO_OUT_TT_PROJECT7
+ Tile_X0Y4_CLK_TT_PROJECT Tile_X0Y4_ENA_TT_PROJECT Tile_X0Y4_RST_N_TT_PROJECT Tile_X0Y4_UIO_IN_TT_PROJECT0
+ Tile_X0Y4_UIO_IN_TT_PROJECT1 Tile_X0Y4_UIO_IN_TT_PROJECT2 Tile_X0Y4_UIO_IN_TT_PROJECT3
+ Tile_X0Y4_UIO_IN_TT_PROJECT4 Tile_X0Y4_UIO_IN_TT_PROJECT5 Tile_X0Y4_UIO_IN_TT_PROJECT6
+ Tile_X0Y4_UIO_IN_TT_PROJECT7 Tile_X0Y4_UIO_OE_TT_PROJECT0 Tile_X0Y4_UIO_OE_TT_PROJECT1
+ Tile_X0Y4_UIO_OE_TT_PROJECT2 Tile_X0Y4_UIO_OE_TT_PROJECT3 Tile_X0Y4_UIO_OE_TT_PROJECT4
+ Tile_X0Y4_UIO_OE_TT_PROJECT5 Tile_X0Y4_UIO_OE_TT_PROJECT6 Tile_X0Y4_UIO_OE_TT_PROJECT7
+ Tile_X0Y4_UIO_OUT_TT_PROJECT0 Tile_X0Y4_UIO_OUT_TT_PROJECT1 Tile_X0Y4_UIO_OUT_TT_PROJECT2
+ Tile_X0Y4_UIO_OUT_TT_PROJECT3 Tile_X0Y4_UIO_OUT_TT_PROJECT4 Tile_X0Y4_UIO_OUT_TT_PROJECT5
+ Tile_X0Y4_UIO_OUT_TT_PROJECT6 Tile_X0Y4_UIO_OUT_TT_PROJECT7 Tile_X0Y4_UI_IN_TT_PROJECT0
+ Tile_X0Y4_UI_IN_TT_PROJECT1 Tile_X0Y4_UI_IN_TT_PROJECT2 Tile_X0Y4_UI_IN_TT_PROJECT3
+ Tile_X0Y4_UI_IN_TT_PROJECT4 Tile_X0Y4_UI_IN_TT_PROJECT5 Tile_X0Y4_UI_IN_TT_PROJECT6
+ Tile_X0Y4_UI_IN_TT_PROJECT7 Tile_X0Y4_UO_OUT_TT_PROJECT0 Tile_X0Y4_UO_OUT_TT_PROJECT1
+ Tile_X0Y4_UO_OUT_TT_PROJECT2 Tile_X0Y4_UO_OUT_TT_PROJECT3 Tile_X0Y4_UO_OUT_TT_PROJECT4
+ Tile_X0Y4_UO_OUT_TT_PROJECT5 Tile_X0Y4_UO_OUT_TT_PROJECT6 Tile_X0Y4_UO_OUT_TT_PROJECT7
+ Tile_X0Y5_CLK_TT_PROJECT Tile_X0Y5_ENA_TT_PROJECT Tile_X0Y5_RST_N_TT_PROJECT Tile_X0Y5_UIO_IN_TT_PROJECT0
+ Tile_X0Y5_UIO_IN_TT_PROJECT1 Tile_X0Y5_UIO_IN_TT_PROJECT2 Tile_X0Y5_UIO_IN_TT_PROJECT3
+ Tile_X0Y5_UIO_IN_TT_PROJECT4 Tile_X0Y5_UIO_IN_TT_PROJECT5 Tile_X0Y5_UIO_IN_TT_PROJECT6
+ Tile_X0Y5_UIO_IN_TT_PROJECT7 Tile_X0Y5_UIO_OE_TT_PROJECT0 Tile_X0Y5_UIO_OE_TT_PROJECT1
+ Tile_X0Y5_UIO_OE_TT_PROJECT2 Tile_X0Y5_UIO_OE_TT_PROJECT3 Tile_X0Y5_UIO_OE_TT_PROJECT4
+ Tile_X0Y5_UIO_OE_TT_PROJECT5 Tile_X0Y5_UIO_OE_TT_PROJECT6 Tile_X0Y5_UIO_OE_TT_PROJECT7
+ Tile_X0Y5_UIO_OUT_TT_PROJECT0 Tile_X0Y5_UIO_OUT_TT_PROJECT1 Tile_X0Y5_UIO_OUT_TT_PROJECT2
+ Tile_X0Y5_UIO_OUT_TT_PROJECT3 Tile_X0Y5_UIO_OUT_TT_PROJECT4 Tile_X0Y5_UIO_OUT_TT_PROJECT5
+ Tile_X0Y5_UIO_OUT_TT_PROJECT6 Tile_X0Y5_UIO_OUT_TT_PROJECT7 Tile_X0Y5_UI_IN_TT_PROJECT0
+ Tile_X0Y5_UI_IN_TT_PROJECT1 Tile_X0Y5_UI_IN_TT_PROJECT2 Tile_X0Y5_UI_IN_TT_PROJECT3
+ Tile_X0Y5_UI_IN_TT_PROJECT4 Tile_X0Y5_UI_IN_TT_PROJECT5 Tile_X0Y5_UI_IN_TT_PROJECT6
+ Tile_X0Y5_UI_IN_TT_PROJECT7 Tile_X0Y5_UO_OUT_TT_PROJECT0 Tile_X0Y5_UO_OUT_TT_PROJECT1
+ Tile_X0Y5_UO_OUT_TT_PROJECT2 Tile_X0Y5_UO_OUT_TT_PROJECT3 Tile_X0Y5_UO_OUT_TT_PROJECT4
+ Tile_X0Y5_UO_OUT_TT_PROJECT5 Tile_X0Y5_UO_OUT_TT_PROJECT6 Tile_X0Y5_UO_OUT_TT_PROJECT7
+ Tile_X0Y6_CLK_TT_PROJECT Tile_X0Y6_ENA_TT_PROJECT Tile_X0Y6_RST_N_TT_PROJECT Tile_X0Y6_UIO_IN_TT_PROJECT0
+ Tile_X0Y6_UIO_IN_TT_PROJECT1 Tile_X0Y6_UIO_IN_TT_PROJECT2 Tile_X0Y6_UIO_IN_TT_PROJECT3
+ Tile_X0Y6_UIO_IN_TT_PROJECT4 Tile_X0Y6_UIO_IN_TT_PROJECT5 Tile_X0Y6_UIO_IN_TT_PROJECT6
+ Tile_X0Y6_UIO_IN_TT_PROJECT7 Tile_X0Y6_UIO_OE_TT_PROJECT0 Tile_X0Y6_UIO_OE_TT_PROJECT1
+ Tile_X0Y6_UIO_OE_TT_PROJECT2 Tile_X0Y6_UIO_OE_TT_PROJECT3 Tile_X0Y6_UIO_OE_TT_PROJECT4
+ Tile_X0Y6_UIO_OE_TT_PROJECT5 Tile_X0Y6_UIO_OE_TT_PROJECT6 Tile_X0Y6_UIO_OE_TT_PROJECT7
+ Tile_X0Y6_UIO_OUT_TT_PROJECT0 Tile_X0Y6_UIO_OUT_TT_PROJECT1 Tile_X0Y6_UIO_OUT_TT_PROJECT2
+ Tile_X0Y6_UIO_OUT_TT_PROJECT3 Tile_X0Y6_UIO_OUT_TT_PROJECT4 Tile_X0Y6_UIO_OUT_TT_PROJECT5
+ Tile_X0Y6_UIO_OUT_TT_PROJECT6 Tile_X0Y6_UIO_OUT_TT_PROJECT7 Tile_X0Y6_UI_IN_TT_PROJECT0
+ Tile_X0Y6_UI_IN_TT_PROJECT1 Tile_X0Y6_UI_IN_TT_PROJECT2 Tile_X0Y6_UI_IN_TT_PROJECT3
+ Tile_X0Y6_UI_IN_TT_PROJECT4 Tile_X0Y6_UI_IN_TT_PROJECT5 Tile_X0Y6_UI_IN_TT_PROJECT6
+ Tile_X0Y6_UI_IN_TT_PROJECT7 Tile_X0Y6_UO_OUT_TT_PROJECT0 Tile_X0Y6_UO_OUT_TT_PROJECT1
+ Tile_X0Y6_UO_OUT_TT_PROJECT2 Tile_X0Y6_UO_OUT_TT_PROJECT3 Tile_X0Y6_UO_OUT_TT_PROJECT4
+ Tile_X0Y6_UO_OUT_TT_PROJECT5 Tile_X0Y6_UO_OUT_TT_PROJECT6 Tile_X0Y6_UO_OUT_TT_PROJECT7
+ Tile_X0Y7_CLK_TT_PROJECT Tile_X0Y7_ENA_TT_PROJECT Tile_X0Y7_RST_N_TT_PROJECT Tile_X0Y7_UIO_IN_TT_PROJECT0
+ Tile_X0Y7_UIO_IN_TT_PROJECT1 Tile_X0Y7_UIO_IN_TT_PROJECT2 Tile_X0Y7_UIO_IN_TT_PROJECT3
+ Tile_X0Y7_UIO_IN_TT_PROJECT4 Tile_X0Y7_UIO_IN_TT_PROJECT5 Tile_X0Y7_UIO_IN_TT_PROJECT6
+ Tile_X0Y7_UIO_IN_TT_PROJECT7 Tile_X0Y7_UIO_OE_TT_PROJECT0 Tile_X0Y7_UIO_OE_TT_PROJECT1
+ Tile_X0Y7_UIO_OE_TT_PROJECT2 Tile_X0Y7_UIO_OE_TT_PROJECT3 Tile_X0Y7_UIO_OE_TT_PROJECT4
+ Tile_X0Y7_UIO_OE_TT_PROJECT5 Tile_X0Y7_UIO_OE_TT_PROJECT6 Tile_X0Y7_UIO_OE_TT_PROJECT7
+ Tile_X0Y7_UIO_OUT_TT_PROJECT0 Tile_X0Y7_UIO_OUT_TT_PROJECT1 Tile_X0Y7_UIO_OUT_TT_PROJECT2
+ Tile_X0Y7_UIO_OUT_TT_PROJECT3 Tile_X0Y7_UIO_OUT_TT_PROJECT4 Tile_X0Y7_UIO_OUT_TT_PROJECT5
+ Tile_X0Y7_UIO_OUT_TT_PROJECT6 Tile_X0Y7_UIO_OUT_TT_PROJECT7 Tile_X0Y7_UI_IN_TT_PROJECT0
+ Tile_X0Y7_UI_IN_TT_PROJECT1 Tile_X0Y7_UI_IN_TT_PROJECT2 Tile_X0Y7_UI_IN_TT_PROJECT3
+ Tile_X0Y7_UI_IN_TT_PROJECT4 Tile_X0Y7_UI_IN_TT_PROJECT5 Tile_X0Y7_UI_IN_TT_PROJECT6
+ Tile_X0Y7_UI_IN_TT_PROJECT7 Tile_X0Y7_UO_OUT_TT_PROJECT0 Tile_X0Y7_UO_OUT_TT_PROJECT1
+ Tile_X0Y7_UO_OUT_TT_PROJECT2 Tile_X0Y7_UO_OUT_TT_PROJECT3 Tile_X0Y7_UO_OUT_TT_PROJECT4
+ Tile_X0Y7_UO_OUT_TT_PROJECT5 Tile_X0Y7_UO_OUT_TT_PROJECT6 Tile_X0Y7_UO_OUT_TT_PROJECT7
+ Tile_X0Y8_CLK_TT_PROJECT Tile_X0Y8_ENA_TT_PROJECT Tile_X0Y8_RST_N_TT_PROJECT Tile_X0Y8_UIO_IN_TT_PROJECT0
+ Tile_X0Y8_UIO_IN_TT_PROJECT1 Tile_X0Y8_UIO_IN_TT_PROJECT2 Tile_X0Y8_UIO_IN_TT_PROJECT3
+ Tile_X0Y8_UIO_IN_TT_PROJECT4 Tile_X0Y8_UIO_IN_TT_PROJECT5 Tile_X0Y8_UIO_IN_TT_PROJECT6
+ Tile_X0Y8_UIO_IN_TT_PROJECT7 Tile_X0Y8_UIO_OE_TT_PROJECT0 Tile_X0Y8_UIO_OE_TT_PROJECT1
+ Tile_X0Y8_UIO_OE_TT_PROJECT2 Tile_X0Y8_UIO_OE_TT_PROJECT3 Tile_X0Y8_UIO_OE_TT_PROJECT4
+ Tile_X0Y8_UIO_OE_TT_PROJECT5 Tile_X0Y8_UIO_OE_TT_PROJECT6 Tile_X0Y8_UIO_OE_TT_PROJECT7
+ Tile_X0Y8_UIO_OUT_TT_PROJECT0 Tile_X0Y8_UIO_OUT_TT_PROJECT1 Tile_X0Y8_UIO_OUT_TT_PROJECT2
+ Tile_X0Y8_UIO_OUT_TT_PROJECT3 Tile_X0Y8_UIO_OUT_TT_PROJECT4 Tile_X0Y8_UIO_OUT_TT_PROJECT5
+ Tile_X0Y8_UIO_OUT_TT_PROJECT6 Tile_X0Y8_UIO_OUT_TT_PROJECT7 Tile_X0Y8_UI_IN_TT_PROJECT0
+ Tile_X0Y8_UI_IN_TT_PROJECT1 Tile_X0Y8_UI_IN_TT_PROJECT2 Tile_X0Y8_UI_IN_TT_PROJECT3
+ Tile_X0Y8_UI_IN_TT_PROJECT4 Tile_X0Y8_UI_IN_TT_PROJECT5 Tile_X0Y8_UI_IN_TT_PROJECT6
+ Tile_X0Y8_UI_IN_TT_PROJECT7 Tile_X0Y8_UO_OUT_TT_PROJECT0 Tile_X0Y8_UO_OUT_TT_PROJECT1
+ Tile_X0Y8_UO_OUT_TT_PROJECT2 Tile_X0Y8_UO_OUT_TT_PROJECT3 Tile_X0Y8_UO_OUT_TT_PROJECT4
+ Tile_X0Y8_UO_OUT_TT_PROJECT5 Tile_X0Y8_UO_OUT_TT_PROJECT6 Tile_X0Y8_UO_OUT_TT_PROJECT7
+ Tile_X1Y0_A_I_top Tile_X1Y0_A_O_top Tile_X1Y0_A_T_top Tile_X1Y0_B_I_top Tile_X1Y0_B_O_top
+ Tile_X1Y0_B_T_top Tile_X1Y0_C_I_top Tile_X1Y0_C_O_top Tile_X1Y0_C_T_top Tile_X1Y0_D_I_top
+ Tile_X1Y0_D_O_top Tile_X1Y0_D_T_top Tile_X1Y9_A_I_top Tile_X1Y9_A_O_top Tile_X1Y9_A_T_top
+ Tile_X1Y9_B_I_top Tile_X1Y9_B_O_top Tile_X1Y9_B_T_top Tile_X1Y9_C_I_top Tile_X1Y9_C_O_top
+ Tile_X1Y9_C_T_top Tile_X1Y9_D_I_top Tile_X1Y9_D_O_top Tile_X1Y9_D_T_top Tile_X2Y0_A_I_top
+ Tile_X2Y0_A_O_top Tile_X2Y0_A_T_top Tile_X2Y0_B_I_top Tile_X2Y0_B_O_top Tile_X2Y0_B_T_top
+ Tile_X2Y0_C_I_top Tile_X2Y0_C_O_top Tile_X2Y0_C_T_top Tile_X2Y0_D_I_top Tile_X2Y0_D_O_top
+ Tile_X2Y0_D_T_top Tile_X2Y9_A_I_top Tile_X2Y9_A_O_top Tile_X2Y9_A_T_top Tile_X2Y9_B_I_top
+ Tile_X2Y9_B_O_top Tile_X2Y9_B_T_top Tile_X2Y9_C_I_top Tile_X2Y9_C_O_top Tile_X2Y9_C_T_top
+ Tile_X2Y9_D_I_top Tile_X2Y9_D_O_top Tile_X2Y9_D_T_top Tile_X3Y0_A_I_top Tile_X3Y0_A_O_top
+ Tile_X3Y0_A_T_top Tile_X3Y0_B_I_top Tile_X3Y0_B_O_top Tile_X3Y0_B_T_top Tile_X3Y0_C_I_top
+ Tile_X3Y0_C_O_top Tile_X3Y0_C_T_top Tile_X3Y0_D_I_top Tile_X3Y0_D_O_top Tile_X3Y0_D_T_top
+ Tile_X3Y9_A_I_top Tile_X3Y9_A_O_top Tile_X3Y9_A_T_top Tile_X3Y9_B_I_top Tile_X3Y9_B_O_top
+ Tile_X3Y9_B_T_top Tile_X3Y9_C_I_top Tile_X3Y9_C_O_top Tile_X3Y9_C_T_top Tile_X3Y9_D_I_top
+ Tile_X3Y9_D_O_top Tile_X3Y9_D_T_top Tile_X4Y0_A_I_top Tile_X4Y0_A_O_top Tile_X4Y0_A_T_top
+ Tile_X4Y0_B_I_top Tile_X4Y0_B_O_top Tile_X4Y0_B_T_top Tile_X4Y0_C_I_top Tile_X4Y0_C_O_top
+ Tile_X4Y0_C_T_top Tile_X4Y0_D_I_top Tile_X4Y0_D_O_top Tile_X4Y0_D_T_top Tile_X4Y9_A_I_top
+ Tile_X4Y9_A_O_top Tile_X4Y9_A_T_top Tile_X4Y9_B_I_top Tile_X4Y9_B_O_top Tile_X4Y9_B_T_top
+ Tile_X4Y9_C_I_top Tile_X4Y9_C_O_top Tile_X4Y9_C_T_top Tile_X4Y9_D_I_top Tile_X4Y9_D_O_top
+ Tile_X4Y9_D_T_top Tile_X5Y2_ADDR_SRAM0 Tile_X5Y2_ADDR_SRAM1 Tile_X5Y2_ADDR_SRAM2
+ Tile_X5Y2_ADDR_SRAM3 Tile_X5Y2_ADDR_SRAM4 Tile_X5Y2_ADDR_SRAM5 Tile_X5Y2_ADDR_SRAM6
+ Tile_X5Y2_ADDR_SRAM7 Tile_X5Y2_ADDR_SRAM8 Tile_X5Y2_ADDR_SRAM9 Tile_X5Y2_BM_SRAM0
+ Tile_X5Y2_BM_SRAM1 Tile_X5Y2_BM_SRAM10 Tile_X5Y2_BM_SRAM11 Tile_X5Y2_BM_SRAM12 Tile_X5Y2_BM_SRAM13
+ Tile_X5Y2_BM_SRAM14 Tile_X5Y2_BM_SRAM15 Tile_X5Y2_BM_SRAM16 Tile_X5Y2_BM_SRAM17
+ Tile_X5Y2_BM_SRAM18 Tile_X5Y2_BM_SRAM19 Tile_X5Y2_BM_SRAM2 Tile_X5Y2_BM_SRAM20 Tile_X5Y2_BM_SRAM21
+ Tile_X5Y2_BM_SRAM22 Tile_X5Y2_BM_SRAM23 Tile_X5Y2_BM_SRAM24 Tile_X5Y2_BM_SRAM25
+ Tile_X5Y2_BM_SRAM26 Tile_X5Y2_BM_SRAM27 Tile_X5Y2_BM_SRAM28 Tile_X5Y2_BM_SRAM29
+ Tile_X5Y2_BM_SRAM3 Tile_X5Y2_BM_SRAM30 Tile_X5Y2_BM_SRAM31 Tile_X5Y2_BM_SRAM4 Tile_X5Y2_BM_SRAM5
+ Tile_X5Y2_BM_SRAM6 Tile_X5Y2_BM_SRAM7 Tile_X5Y2_BM_SRAM8 Tile_X5Y2_BM_SRAM9 Tile_X5Y2_CLK_SRAM
+ Tile_X5Y2_CONFIGURED_top Tile_X5Y2_DIN_SRAM0 Tile_X5Y2_DIN_SRAM1 Tile_X5Y2_DIN_SRAM10
+ Tile_X5Y2_DIN_SRAM11 Tile_X5Y2_DIN_SRAM12 Tile_X5Y2_DIN_SRAM13 Tile_X5Y2_DIN_SRAM14
+ Tile_X5Y2_DIN_SRAM15 Tile_X5Y2_DIN_SRAM16 Tile_X5Y2_DIN_SRAM17 Tile_X5Y2_DIN_SRAM18
+ Tile_X5Y2_DIN_SRAM19 Tile_X5Y2_DIN_SRAM2 Tile_X5Y2_DIN_SRAM20 Tile_X5Y2_DIN_SRAM21
+ Tile_X5Y2_DIN_SRAM22 Tile_X5Y2_DIN_SRAM23 Tile_X5Y2_DIN_SRAM24 Tile_X5Y2_DIN_SRAM25
+ Tile_X5Y2_DIN_SRAM26 Tile_X5Y2_DIN_SRAM27 Tile_X5Y2_DIN_SRAM28 Tile_X5Y2_DIN_SRAM29
+ Tile_X5Y2_DIN_SRAM3 Tile_X5Y2_DIN_SRAM30 Tile_X5Y2_DIN_SRAM31 Tile_X5Y2_DIN_SRAM4
+ Tile_X5Y2_DIN_SRAM5 Tile_X5Y2_DIN_SRAM6 Tile_X5Y2_DIN_SRAM7 Tile_X5Y2_DIN_SRAM8
+ Tile_X5Y2_DIN_SRAM9 Tile_X5Y2_DOUT_SRAM0 Tile_X5Y2_DOUT_SRAM1 Tile_X5Y2_DOUT_SRAM10
+ Tile_X5Y2_DOUT_SRAM11 Tile_X5Y2_DOUT_SRAM12 Tile_X5Y2_DOUT_SRAM13 Tile_X5Y2_DOUT_SRAM14
+ Tile_X5Y2_DOUT_SRAM15 Tile_X5Y2_DOUT_SRAM16 Tile_X5Y2_DOUT_SRAM17 Tile_X5Y2_DOUT_SRAM18
+ Tile_X5Y2_DOUT_SRAM19 Tile_X5Y2_DOUT_SRAM2 Tile_X5Y2_DOUT_SRAM20 Tile_X5Y2_DOUT_SRAM21
+ Tile_X5Y2_DOUT_SRAM22 Tile_X5Y2_DOUT_SRAM23 Tile_X5Y2_DOUT_SRAM24 Tile_X5Y2_DOUT_SRAM25
+ Tile_X5Y2_DOUT_SRAM26 Tile_X5Y2_DOUT_SRAM27 Tile_X5Y2_DOUT_SRAM28 Tile_X5Y2_DOUT_SRAM29
+ Tile_X5Y2_DOUT_SRAM3 Tile_X5Y2_DOUT_SRAM30 Tile_X5Y2_DOUT_SRAM31 Tile_X5Y2_DOUT_SRAM4
+ Tile_X5Y2_DOUT_SRAM5 Tile_X5Y2_DOUT_SRAM6 Tile_X5Y2_DOUT_SRAM7 Tile_X5Y2_DOUT_SRAM8
+ Tile_X5Y2_DOUT_SRAM9 Tile_X5Y2_MEN_SRAM Tile_X5Y2_REN_SRAM Tile_X5Y2_TIE_HIGH_SRAM
+ Tile_X5Y2_TIE_LOW_SRAM Tile_X5Y2_WEN_SRAM Tile_X5Y3_CLK_TT_PROJECT Tile_X5Y3_ENA_TT_PROJECT
+ Tile_X5Y3_RST_N_TT_PROJECT Tile_X5Y3_UIO_IN_TT_PROJECT0 Tile_X5Y3_UIO_IN_TT_PROJECT1
+ Tile_X5Y3_UIO_IN_TT_PROJECT2 Tile_X5Y3_UIO_IN_TT_PROJECT3 Tile_X5Y3_UIO_IN_TT_PROJECT4
+ Tile_X5Y3_UIO_IN_TT_PROJECT5 Tile_X5Y3_UIO_IN_TT_PROJECT6 Tile_X5Y3_UIO_IN_TT_PROJECT7
+ Tile_X5Y3_UIO_OE_TT_PROJECT0 Tile_X5Y3_UIO_OE_TT_PROJECT1 Tile_X5Y3_UIO_OE_TT_PROJECT2
+ Tile_X5Y3_UIO_OE_TT_PROJECT3 Tile_X5Y3_UIO_OE_TT_PROJECT4 Tile_X5Y3_UIO_OE_TT_PROJECT5
+ Tile_X5Y3_UIO_OE_TT_PROJECT6 Tile_X5Y3_UIO_OE_TT_PROJECT7 Tile_X5Y3_UIO_OUT_TT_PROJECT0
+ Tile_X5Y3_UIO_OUT_TT_PROJECT1 Tile_X5Y3_UIO_OUT_TT_PROJECT2 Tile_X5Y3_UIO_OUT_TT_PROJECT3
+ Tile_X5Y3_UIO_OUT_TT_PROJECT4 Tile_X5Y3_UIO_OUT_TT_PROJECT5 Tile_X5Y3_UIO_OUT_TT_PROJECT6
+ Tile_X5Y3_UIO_OUT_TT_PROJECT7 Tile_X5Y3_UI_IN_TT_PROJECT0 Tile_X5Y3_UI_IN_TT_PROJECT1
+ Tile_X5Y3_UI_IN_TT_PROJECT2 Tile_X5Y3_UI_IN_TT_PROJECT3 Tile_X5Y3_UI_IN_TT_PROJECT4
+ Tile_X5Y3_UI_IN_TT_PROJECT5 Tile_X5Y3_UI_IN_TT_PROJECT6 Tile_X5Y3_UI_IN_TT_PROJECT7
+ Tile_X5Y3_UO_OUT_TT_PROJECT0 Tile_X5Y3_UO_OUT_TT_PROJECT1 Tile_X5Y3_UO_OUT_TT_PROJECT2
+ Tile_X5Y3_UO_OUT_TT_PROJECT3 Tile_X5Y3_UO_OUT_TT_PROJECT4 Tile_X5Y3_UO_OUT_TT_PROJECT5
+ Tile_X5Y3_UO_OUT_TT_PROJECT6 Tile_X5Y3_UO_OUT_TT_PROJECT7 Tile_X5Y4_CLK_TT_PROJECT
+ Tile_X5Y4_ENA_TT_PROJECT Tile_X5Y4_RST_N_TT_PROJECT Tile_X5Y4_UIO_IN_TT_PROJECT0
+ Tile_X5Y4_UIO_IN_TT_PROJECT1 Tile_X5Y4_UIO_IN_TT_PROJECT2 Tile_X5Y4_UIO_IN_TT_PROJECT3
+ Tile_X5Y4_UIO_IN_TT_PROJECT4 Tile_X5Y4_UIO_IN_TT_PROJECT5 Tile_X5Y4_UIO_IN_TT_PROJECT6
+ Tile_X5Y4_UIO_IN_TT_PROJECT7 Tile_X5Y4_UIO_OE_TT_PROJECT0 Tile_X5Y4_UIO_OE_TT_PROJECT1
+ Tile_X5Y4_UIO_OE_TT_PROJECT2 Tile_X5Y4_UIO_OE_TT_PROJECT3 Tile_X5Y4_UIO_OE_TT_PROJECT4
+ Tile_X5Y4_UIO_OE_TT_PROJECT5 Tile_X5Y4_UIO_OE_TT_PROJECT6 Tile_X5Y4_UIO_OE_TT_PROJECT7
+ Tile_X5Y4_UIO_OUT_TT_PROJECT0 Tile_X5Y4_UIO_OUT_TT_PROJECT1 Tile_X5Y4_UIO_OUT_TT_PROJECT2
+ Tile_X5Y4_UIO_OUT_TT_PROJECT3 Tile_X5Y4_UIO_OUT_TT_PROJECT4 Tile_X5Y4_UIO_OUT_TT_PROJECT5
+ Tile_X5Y4_UIO_OUT_TT_PROJECT6 Tile_X5Y4_UIO_OUT_TT_PROJECT7 Tile_X5Y4_UI_IN_TT_PROJECT0
+ Tile_X5Y4_UI_IN_TT_PROJECT1 Tile_X5Y4_UI_IN_TT_PROJECT2 Tile_X5Y4_UI_IN_TT_PROJECT3
+ Tile_X5Y4_UI_IN_TT_PROJECT4 Tile_X5Y4_UI_IN_TT_PROJECT5 Tile_X5Y4_UI_IN_TT_PROJECT6
+ Tile_X5Y4_UI_IN_TT_PROJECT7 Tile_X5Y4_UO_OUT_TT_PROJECT0 Tile_X5Y4_UO_OUT_TT_PROJECT1
+ Tile_X5Y4_UO_OUT_TT_PROJECT2 Tile_X5Y4_UO_OUT_TT_PROJECT3 Tile_X5Y4_UO_OUT_TT_PROJECT4
+ Tile_X5Y4_UO_OUT_TT_PROJECT5 Tile_X5Y4_UO_OUT_TT_PROJECT6 Tile_X5Y4_UO_OUT_TT_PROJECT7
+ Tile_X5Y5_CLK_TT_PROJECT Tile_X5Y5_ENA_TT_PROJECT Tile_X5Y5_RST_N_TT_PROJECT Tile_X5Y5_UIO_IN_TT_PROJECT0
+ Tile_X5Y5_UIO_IN_TT_PROJECT1 Tile_X5Y5_UIO_IN_TT_PROJECT2 Tile_X5Y5_UIO_IN_TT_PROJECT3
+ Tile_X5Y5_UIO_IN_TT_PROJECT4 Tile_X5Y5_UIO_IN_TT_PROJECT5 Tile_X5Y5_UIO_IN_TT_PROJECT6
+ Tile_X5Y5_UIO_IN_TT_PROJECT7 Tile_X5Y5_UIO_OE_TT_PROJECT0 Tile_X5Y5_UIO_OE_TT_PROJECT1
+ Tile_X5Y5_UIO_OE_TT_PROJECT2 Tile_X5Y5_UIO_OE_TT_PROJECT3 Tile_X5Y5_UIO_OE_TT_PROJECT4
+ Tile_X5Y5_UIO_OE_TT_PROJECT5 Tile_X5Y5_UIO_OE_TT_PROJECT6 Tile_X5Y5_UIO_OE_TT_PROJECT7
+ Tile_X5Y5_UIO_OUT_TT_PROJECT0 Tile_X5Y5_UIO_OUT_TT_PROJECT1 Tile_X5Y5_UIO_OUT_TT_PROJECT2
+ Tile_X5Y5_UIO_OUT_TT_PROJECT3 Tile_X5Y5_UIO_OUT_TT_PROJECT4 Tile_X5Y5_UIO_OUT_TT_PROJECT5
+ Tile_X5Y5_UIO_OUT_TT_PROJECT6 Tile_X5Y5_UIO_OUT_TT_PROJECT7 Tile_X5Y5_UI_IN_TT_PROJECT0
+ Tile_X5Y5_UI_IN_TT_PROJECT1 Tile_X5Y5_UI_IN_TT_PROJECT2 Tile_X5Y5_UI_IN_TT_PROJECT3
+ Tile_X5Y5_UI_IN_TT_PROJECT4 Tile_X5Y5_UI_IN_TT_PROJECT5 Tile_X5Y5_UI_IN_TT_PROJECT6
+ Tile_X5Y5_UI_IN_TT_PROJECT7 Tile_X5Y5_UO_OUT_TT_PROJECT0 Tile_X5Y5_UO_OUT_TT_PROJECT1
+ Tile_X5Y5_UO_OUT_TT_PROJECT2 Tile_X5Y5_UO_OUT_TT_PROJECT3 Tile_X5Y5_UO_OUT_TT_PROJECT4
+ Tile_X5Y5_UO_OUT_TT_PROJECT5 Tile_X5Y5_UO_OUT_TT_PROJECT6 Tile_X5Y5_UO_OUT_TT_PROJECT7
+ Tile_X5Y6_CLK_TT_PROJECT Tile_X5Y6_ENA_TT_PROJECT Tile_X5Y6_RST_N_TT_PROJECT Tile_X5Y6_UIO_IN_TT_PROJECT0
+ Tile_X5Y6_UIO_IN_TT_PROJECT1 Tile_X5Y6_UIO_IN_TT_PROJECT2 Tile_X5Y6_UIO_IN_TT_PROJECT3
+ Tile_X5Y6_UIO_IN_TT_PROJECT4 Tile_X5Y6_UIO_IN_TT_PROJECT5 Tile_X5Y6_UIO_IN_TT_PROJECT6
+ Tile_X5Y6_UIO_IN_TT_PROJECT7 Tile_X5Y6_UIO_OE_TT_PROJECT0 Tile_X5Y6_UIO_OE_TT_PROJECT1
+ Tile_X5Y6_UIO_OE_TT_PROJECT2 Tile_X5Y6_UIO_OE_TT_PROJECT3 Tile_X5Y6_UIO_OE_TT_PROJECT4
+ Tile_X5Y6_UIO_OE_TT_PROJECT5 Tile_X5Y6_UIO_OE_TT_PROJECT6 Tile_X5Y6_UIO_OE_TT_PROJECT7
+ Tile_X5Y6_UIO_OUT_TT_PROJECT0 Tile_X5Y6_UIO_OUT_TT_PROJECT1 Tile_X5Y6_UIO_OUT_TT_PROJECT2
+ Tile_X5Y6_UIO_OUT_TT_PROJECT3 Tile_X5Y6_UIO_OUT_TT_PROJECT4 Tile_X5Y6_UIO_OUT_TT_PROJECT5
+ Tile_X5Y6_UIO_OUT_TT_PROJECT6 Tile_X5Y6_UIO_OUT_TT_PROJECT7 Tile_X5Y6_UI_IN_TT_PROJECT0
+ Tile_X5Y6_UI_IN_TT_PROJECT1 Tile_X5Y6_UI_IN_TT_PROJECT2 Tile_X5Y6_UI_IN_TT_PROJECT3
+ Tile_X5Y6_UI_IN_TT_PROJECT4 Tile_X5Y6_UI_IN_TT_PROJECT5 Tile_X5Y6_UI_IN_TT_PROJECT6
+ Tile_X5Y6_UI_IN_TT_PROJECT7 Tile_X5Y6_UO_OUT_TT_PROJECT0 Tile_X5Y6_UO_OUT_TT_PROJECT1
+ Tile_X5Y6_UO_OUT_TT_PROJECT2 Tile_X5Y6_UO_OUT_TT_PROJECT3 Tile_X5Y6_UO_OUT_TT_PROJECT4
+ Tile_X5Y6_UO_OUT_TT_PROJECT5 Tile_X5Y6_UO_OUT_TT_PROJECT6 Tile_X5Y6_UO_OUT_TT_PROJECT7
+ Tile_X5Y7_CLK_TT_PROJECT Tile_X5Y7_ENA_TT_PROJECT Tile_X5Y7_RST_N_TT_PROJECT Tile_X5Y7_UIO_IN_TT_PROJECT0
+ Tile_X5Y7_UIO_IN_TT_PROJECT1 Tile_X5Y7_UIO_IN_TT_PROJECT2 Tile_X5Y7_UIO_IN_TT_PROJECT3
+ Tile_X5Y7_UIO_IN_TT_PROJECT4 Tile_X5Y7_UIO_IN_TT_PROJECT5 Tile_X5Y7_UIO_IN_TT_PROJECT6
+ Tile_X5Y7_UIO_IN_TT_PROJECT7 Tile_X5Y7_UIO_OE_TT_PROJECT0 Tile_X5Y7_UIO_OE_TT_PROJECT1
+ Tile_X5Y7_UIO_OE_TT_PROJECT2 Tile_X5Y7_UIO_OE_TT_PROJECT3 Tile_X5Y7_UIO_OE_TT_PROJECT4
+ Tile_X5Y7_UIO_OE_TT_PROJECT5 Tile_X5Y7_UIO_OE_TT_PROJECT6 Tile_X5Y7_UIO_OE_TT_PROJECT7
+ Tile_X5Y7_UIO_OUT_TT_PROJECT0 Tile_X5Y7_UIO_OUT_TT_PROJECT1 Tile_X5Y7_UIO_OUT_TT_PROJECT2
+ Tile_X5Y7_UIO_OUT_TT_PROJECT3 Tile_X5Y7_UIO_OUT_TT_PROJECT4 Tile_X5Y7_UIO_OUT_TT_PROJECT5
+ Tile_X5Y7_UIO_OUT_TT_PROJECT6 Tile_X5Y7_UIO_OUT_TT_PROJECT7 Tile_X5Y7_UI_IN_TT_PROJECT0
+ Tile_X5Y7_UI_IN_TT_PROJECT1 Tile_X5Y7_UI_IN_TT_PROJECT2 Tile_X5Y7_UI_IN_TT_PROJECT3
+ Tile_X5Y7_UI_IN_TT_PROJECT4 Tile_X5Y7_UI_IN_TT_PROJECT5 Tile_X5Y7_UI_IN_TT_PROJECT6
+ Tile_X5Y7_UI_IN_TT_PROJECT7 Tile_X5Y7_UO_OUT_TT_PROJECT0 Tile_X5Y7_UO_OUT_TT_PROJECT1
+ Tile_X5Y7_UO_OUT_TT_PROJECT2 Tile_X5Y7_UO_OUT_TT_PROJECT3 Tile_X5Y7_UO_OUT_TT_PROJECT4
+ Tile_X5Y7_UO_OUT_TT_PROJECT5 Tile_X5Y7_UO_OUT_TT_PROJECT6 Tile_X5Y7_UO_OUT_TT_PROJECT7
+ Tile_X5Y8_CLK_TT_PROJECT Tile_X5Y8_ENA_TT_PROJECT Tile_X5Y8_RST_N_TT_PROJECT Tile_X5Y8_UIO_IN_TT_PROJECT0
+ Tile_X5Y8_UIO_IN_TT_PROJECT1 Tile_X5Y8_UIO_IN_TT_PROJECT2 Tile_X5Y8_UIO_IN_TT_PROJECT3
+ Tile_X5Y8_UIO_IN_TT_PROJECT4 Tile_X5Y8_UIO_IN_TT_PROJECT5 Tile_X5Y8_UIO_IN_TT_PROJECT6
+ Tile_X5Y8_UIO_IN_TT_PROJECT7 Tile_X5Y8_UIO_OE_TT_PROJECT0 Tile_X5Y8_UIO_OE_TT_PROJECT1
+ Tile_X5Y8_UIO_OE_TT_PROJECT2 Tile_X5Y8_UIO_OE_TT_PROJECT3 Tile_X5Y8_UIO_OE_TT_PROJECT4
+ Tile_X5Y8_UIO_OE_TT_PROJECT5 Tile_X5Y8_UIO_OE_TT_PROJECT6 Tile_X5Y8_UIO_OE_TT_PROJECT7
+ Tile_X5Y8_UIO_OUT_TT_PROJECT0 Tile_X5Y8_UIO_OUT_TT_PROJECT1 Tile_X5Y8_UIO_OUT_TT_PROJECT2
+ Tile_X5Y8_UIO_OUT_TT_PROJECT3 Tile_X5Y8_UIO_OUT_TT_PROJECT4 Tile_X5Y8_UIO_OUT_TT_PROJECT5
+ Tile_X5Y8_UIO_OUT_TT_PROJECT6 Tile_X5Y8_UIO_OUT_TT_PROJECT7 Tile_X5Y8_UI_IN_TT_PROJECT0
+ Tile_X5Y8_UI_IN_TT_PROJECT1 Tile_X5Y8_UI_IN_TT_PROJECT2 Tile_X5Y8_UI_IN_TT_PROJECT3
+ Tile_X5Y8_UI_IN_TT_PROJECT4 Tile_X5Y8_UI_IN_TT_PROJECT5 Tile_X5Y8_UI_IN_TT_PROJECT6
+ Tile_X5Y8_UI_IN_TT_PROJECT7 Tile_X5Y8_UO_OUT_TT_PROJECT0 Tile_X5Y8_UO_OUT_TT_PROJECT1
+ Tile_X5Y8_UO_OUT_TT_PROJECT2 Tile_X5Y8_UO_OUT_TT_PROJECT3 Tile_X5Y8_UO_OUT_TT_PROJECT4
+ Tile_X5Y8_UO_OUT_TT_PROJECT5 Tile_X5Y8_UO_OUT_TT_PROJECT6 Tile_X5Y8_UO_OUT_TT_PROJECT7
+ UserCLK VGND VPWR
XTile_X3Y3_LUT4AB Tile_X3Y4_LUT4AB/Co Tile_X3Y3_LUT4AB/Co Tile_X4Y3_LUT4AB/E1END[0]
+ Tile_X4Y3_LUT4AB/E1END[1] Tile_X4Y3_LUT4AB/E1END[2] Tile_X4Y3_LUT4AB/E1END[3] Tile_X3Y3_LUT4AB/E1END[0]
+ Tile_X3Y3_LUT4AB/E1END[1] Tile_X3Y3_LUT4AB/E1END[2] Tile_X3Y3_LUT4AB/E1END[3] Tile_X4Y3_LUT4AB/E2MID[0]
+ Tile_X4Y3_LUT4AB/E2MID[1] Tile_X4Y3_LUT4AB/E2MID[2] Tile_X4Y3_LUT4AB/E2MID[3] Tile_X4Y3_LUT4AB/E2MID[4]
+ Tile_X4Y3_LUT4AB/E2MID[5] Tile_X4Y3_LUT4AB/E2MID[6] Tile_X4Y3_LUT4AB/E2MID[7] Tile_X4Y3_LUT4AB/E2END[0]
+ Tile_X4Y3_LUT4AB/E2END[1] Tile_X4Y3_LUT4AB/E2END[2] Tile_X4Y3_LUT4AB/E2END[3] Tile_X4Y3_LUT4AB/E2END[4]
+ Tile_X4Y3_LUT4AB/E2END[5] Tile_X4Y3_LUT4AB/E2END[6] Tile_X4Y3_LUT4AB/E2END[7] Tile_X3Y3_LUT4AB/E2END[0]
+ Tile_X3Y3_LUT4AB/E2END[1] Tile_X3Y3_LUT4AB/E2END[2] Tile_X3Y3_LUT4AB/E2END[3] Tile_X3Y3_LUT4AB/E2END[4]
+ Tile_X3Y3_LUT4AB/E2END[5] Tile_X3Y3_LUT4AB/E2END[6] Tile_X3Y3_LUT4AB/E2END[7] Tile_X3Y3_LUT4AB/E2MID[0]
+ Tile_X3Y3_LUT4AB/E2MID[1] Tile_X3Y3_LUT4AB/E2MID[2] Tile_X3Y3_LUT4AB/E2MID[3] Tile_X3Y3_LUT4AB/E2MID[4]
+ Tile_X3Y3_LUT4AB/E2MID[5] Tile_X3Y3_LUT4AB/E2MID[6] Tile_X3Y3_LUT4AB/E2MID[7] Tile_X4Y3_LUT4AB/E6END[0]
+ Tile_X4Y3_LUT4AB/E6END[10] Tile_X4Y3_LUT4AB/E6END[11] Tile_X4Y3_LUT4AB/E6END[1]
+ Tile_X4Y3_LUT4AB/E6END[2] Tile_X4Y3_LUT4AB/E6END[3] Tile_X4Y3_LUT4AB/E6END[4] Tile_X4Y3_LUT4AB/E6END[5]
+ Tile_X4Y3_LUT4AB/E6END[6] Tile_X4Y3_LUT4AB/E6END[7] Tile_X4Y3_LUT4AB/E6END[8] Tile_X4Y3_LUT4AB/E6END[9]
+ Tile_X3Y3_LUT4AB/E6END[0] Tile_X3Y3_LUT4AB/E6END[10] Tile_X3Y3_LUT4AB/E6END[11]
+ Tile_X3Y3_LUT4AB/E6END[1] Tile_X3Y3_LUT4AB/E6END[2] Tile_X3Y3_LUT4AB/E6END[3] Tile_X3Y3_LUT4AB/E6END[4]
+ Tile_X3Y3_LUT4AB/E6END[5] Tile_X3Y3_LUT4AB/E6END[6] Tile_X3Y3_LUT4AB/E6END[7] Tile_X3Y3_LUT4AB/E6END[8]
+ Tile_X3Y3_LUT4AB/E6END[9] Tile_X4Y3_LUT4AB/EE4END[0] Tile_X4Y3_LUT4AB/EE4END[10]
+ Tile_X4Y3_LUT4AB/EE4END[11] Tile_X4Y3_LUT4AB/EE4END[12] Tile_X4Y3_LUT4AB/EE4END[13]
+ Tile_X4Y3_LUT4AB/EE4END[14] Tile_X4Y3_LUT4AB/EE4END[15] Tile_X4Y3_LUT4AB/EE4END[1]
+ Tile_X4Y3_LUT4AB/EE4END[2] Tile_X4Y3_LUT4AB/EE4END[3] Tile_X4Y3_LUT4AB/EE4END[4]
+ Tile_X4Y3_LUT4AB/EE4END[5] Tile_X4Y3_LUT4AB/EE4END[6] Tile_X4Y3_LUT4AB/EE4END[7]
+ Tile_X4Y3_LUT4AB/EE4END[8] Tile_X4Y3_LUT4AB/EE4END[9] Tile_X3Y3_LUT4AB/EE4END[0]
+ Tile_X3Y3_LUT4AB/EE4END[10] Tile_X3Y3_LUT4AB/EE4END[11] Tile_X3Y3_LUT4AB/EE4END[12]
+ Tile_X3Y3_LUT4AB/EE4END[13] Tile_X3Y3_LUT4AB/EE4END[14] Tile_X3Y3_LUT4AB/EE4END[15]
+ Tile_X3Y3_LUT4AB/EE4END[1] Tile_X3Y3_LUT4AB/EE4END[2] Tile_X3Y3_LUT4AB/EE4END[3]
+ Tile_X3Y3_LUT4AB/EE4END[4] Tile_X3Y3_LUT4AB/EE4END[5] Tile_X3Y3_LUT4AB/EE4END[6]
+ Tile_X3Y3_LUT4AB/EE4END[7] Tile_X3Y3_LUT4AB/EE4END[8] Tile_X3Y3_LUT4AB/EE4END[9]
+ Tile_X3Y3_LUT4AB/FrameData[0] Tile_X3Y3_LUT4AB/FrameData[10] Tile_X3Y3_LUT4AB/FrameData[11]
+ Tile_X3Y3_LUT4AB/FrameData[12] Tile_X3Y3_LUT4AB/FrameData[13] Tile_X3Y3_LUT4AB/FrameData[14]
+ Tile_X3Y3_LUT4AB/FrameData[15] Tile_X3Y3_LUT4AB/FrameData[16] Tile_X3Y3_LUT4AB/FrameData[17]
+ Tile_X3Y3_LUT4AB/FrameData[18] Tile_X3Y3_LUT4AB/FrameData[19] Tile_X3Y3_LUT4AB/FrameData[1]
+ Tile_X3Y3_LUT4AB/FrameData[20] Tile_X3Y3_LUT4AB/FrameData[21] Tile_X3Y3_LUT4AB/FrameData[22]
+ Tile_X3Y3_LUT4AB/FrameData[23] Tile_X3Y3_LUT4AB/FrameData[24] Tile_X3Y3_LUT4AB/FrameData[25]
+ Tile_X3Y3_LUT4AB/FrameData[26] Tile_X3Y3_LUT4AB/FrameData[27] Tile_X3Y3_LUT4AB/FrameData[28]
+ Tile_X3Y3_LUT4AB/FrameData[29] Tile_X3Y3_LUT4AB/FrameData[2] Tile_X3Y3_LUT4AB/FrameData[30]
+ Tile_X3Y3_LUT4AB/FrameData[31] Tile_X3Y3_LUT4AB/FrameData[3] Tile_X3Y3_LUT4AB/FrameData[4]
+ Tile_X3Y3_LUT4AB/FrameData[5] Tile_X3Y3_LUT4AB/FrameData[6] Tile_X3Y3_LUT4AB/FrameData[7]
+ Tile_X3Y3_LUT4AB/FrameData[8] Tile_X3Y3_LUT4AB/FrameData[9] Tile_X4Y3_LUT4AB/FrameData[0]
+ Tile_X4Y3_LUT4AB/FrameData[10] Tile_X4Y3_LUT4AB/FrameData[11] Tile_X4Y3_LUT4AB/FrameData[12]
+ Tile_X4Y3_LUT4AB/FrameData[13] Tile_X4Y3_LUT4AB/FrameData[14] Tile_X4Y3_LUT4AB/FrameData[15]
+ Tile_X4Y3_LUT4AB/FrameData[16] Tile_X4Y3_LUT4AB/FrameData[17] Tile_X4Y3_LUT4AB/FrameData[18]
+ Tile_X4Y3_LUT4AB/FrameData[19] Tile_X4Y3_LUT4AB/FrameData[1] Tile_X4Y3_LUT4AB/FrameData[20]
+ Tile_X4Y3_LUT4AB/FrameData[21] Tile_X4Y3_LUT4AB/FrameData[22] Tile_X4Y3_LUT4AB/FrameData[23]
+ Tile_X4Y3_LUT4AB/FrameData[24] Tile_X4Y3_LUT4AB/FrameData[25] Tile_X4Y3_LUT4AB/FrameData[26]
+ Tile_X4Y3_LUT4AB/FrameData[27] Tile_X4Y3_LUT4AB/FrameData[28] Tile_X4Y3_LUT4AB/FrameData[29]
+ Tile_X4Y3_LUT4AB/FrameData[2] Tile_X4Y3_LUT4AB/FrameData[30] Tile_X4Y3_LUT4AB/FrameData[31]
+ Tile_X4Y3_LUT4AB/FrameData[3] Tile_X4Y3_LUT4AB/FrameData[4] Tile_X4Y3_LUT4AB/FrameData[5]
+ Tile_X4Y3_LUT4AB/FrameData[6] Tile_X4Y3_LUT4AB/FrameData[7] Tile_X4Y3_LUT4AB/FrameData[8]
+ Tile_X4Y3_LUT4AB/FrameData[9] Tile_X3Y3_LUT4AB/FrameStrobe[0] Tile_X3Y3_LUT4AB/FrameStrobe[10]
+ Tile_X3Y3_LUT4AB/FrameStrobe[11] Tile_X3Y3_LUT4AB/FrameStrobe[12] Tile_X3Y3_LUT4AB/FrameStrobe[13]
+ Tile_X3Y3_LUT4AB/FrameStrobe[14] Tile_X3Y3_LUT4AB/FrameStrobe[15] Tile_X3Y3_LUT4AB/FrameStrobe[16]
+ Tile_X3Y3_LUT4AB/FrameStrobe[17] Tile_X3Y3_LUT4AB/FrameStrobe[18] Tile_X3Y3_LUT4AB/FrameStrobe[19]
+ Tile_X3Y3_LUT4AB/FrameStrobe[1] Tile_X3Y3_LUT4AB/FrameStrobe[2] Tile_X3Y3_LUT4AB/FrameStrobe[3]
+ Tile_X3Y3_LUT4AB/FrameStrobe[4] Tile_X3Y3_LUT4AB/FrameStrobe[5] Tile_X3Y3_LUT4AB/FrameStrobe[6]
+ Tile_X3Y3_LUT4AB/FrameStrobe[7] Tile_X3Y3_LUT4AB/FrameStrobe[8] Tile_X3Y3_LUT4AB/FrameStrobe[9]
+ Tile_X3Y2_LUT4AB/FrameStrobe[0] Tile_X3Y2_LUT4AB/FrameStrobe[10] Tile_X3Y2_LUT4AB/FrameStrobe[11]
+ Tile_X3Y2_LUT4AB/FrameStrobe[12] Tile_X3Y2_LUT4AB/FrameStrobe[13] Tile_X3Y2_LUT4AB/FrameStrobe[14]
+ Tile_X3Y2_LUT4AB/FrameStrobe[15] Tile_X3Y2_LUT4AB/FrameStrobe[16] Tile_X3Y2_LUT4AB/FrameStrobe[17]
+ Tile_X3Y2_LUT4AB/FrameStrobe[18] Tile_X3Y2_LUT4AB/FrameStrobe[19] Tile_X3Y2_LUT4AB/FrameStrobe[1]
+ Tile_X3Y2_LUT4AB/FrameStrobe[2] Tile_X3Y2_LUT4AB/FrameStrobe[3] Tile_X3Y2_LUT4AB/FrameStrobe[4]
+ Tile_X3Y2_LUT4AB/FrameStrobe[5] Tile_X3Y2_LUT4AB/FrameStrobe[6] Tile_X3Y2_LUT4AB/FrameStrobe[7]
+ Tile_X3Y2_LUT4AB/FrameStrobe[8] Tile_X3Y2_LUT4AB/FrameStrobe[9] Tile_X3Y3_LUT4AB/N1BEG[0]
+ Tile_X3Y3_LUT4AB/N1BEG[1] Tile_X3Y3_LUT4AB/N1BEG[2] Tile_X3Y3_LUT4AB/N1BEG[3] Tile_X3Y4_LUT4AB/N1BEG[0]
+ Tile_X3Y4_LUT4AB/N1BEG[1] Tile_X3Y4_LUT4AB/N1BEG[2] Tile_X3Y4_LUT4AB/N1BEG[3] Tile_X3Y3_LUT4AB/N2BEG[0]
+ Tile_X3Y3_LUT4AB/N2BEG[1] Tile_X3Y3_LUT4AB/N2BEG[2] Tile_X3Y3_LUT4AB/N2BEG[3] Tile_X3Y3_LUT4AB/N2BEG[4]
+ Tile_X3Y3_LUT4AB/N2BEG[5] Tile_X3Y3_LUT4AB/N2BEG[6] Tile_X3Y3_LUT4AB/N2BEG[7] Tile_X3Y2_LUT4AB/N2END[0]
+ Tile_X3Y2_LUT4AB/N2END[1] Tile_X3Y2_LUT4AB/N2END[2] Tile_X3Y2_LUT4AB/N2END[3] Tile_X3Y2_LUT4AB/N2END[4]
+ Tile_X3Y2_LUT4AB/N2END[5] Tile_X3Y2_LUT4AB/N2END[6] Tile_X3Y2_LUT4AB/N2END[7] Tile_X3Y3_LUT4AB/N2END[0]
+ Tile_X3Y3_LUT4AB/N2END[1] Tile_X3Y3_LUT4AB/N2END[2] Tile_X3Y3_LUT4AB/N2END[3] Tile_X3Y3_LUT4AB/N2END[4]
+ Tile_X3Y3_LUT4AB/N2END[5] Tile_X3Y3_LUT4AB/N2END[6] Tile_X3Y3_LUT4AB/N2END[7] Tile_X3Y4_LUT4AB/N2BEG[0]
+ Tile_X3Y4_LUT4AB/N2BEG[1] Tile_X3Y4_LUT4AB/N2BEG[2] Tile_X3Y4_LUT4AB/N2BEG[3] Tile_X3Y4_LUT4AB/N2BEG[4]
+ Tile_X3Y4_LUT4AB/N2BEG[5] Tile_X3Y4_LUT4AB/N2BEG[6] Tile_X3Y4_LUT4AB/N2BEG[7] Tile_X3Y3_LUT4AB/N4BEG[0]
+ Tile_X3Y3_LUT4AB/N4BEG[10] Tile_X3Y3_LUT4AB/N4BEG[11] Tile_X3Y3_LUT4AB/N4BEG[12]
+ Tile_X3Y3_LUT4AB/N4BEG[13] Tile_X3Y3_LUT4AB/N4BEG[14] Tile_X3Y3_LUT4AB/N4BEG[15]
+ Tile_X3Y3_LUT4AB/N4BEG[1] Tile_X3Y3_LUT4AB/N4BEG[2] Tile_X3Y3_LUT4AB/N4BEG[3] Tile_X3Y3_LUT4AB/N4BEG[4]
+ Tile_X3Y3_LUT4AB/N4BEG[5] Tile_X3Y3_LUT4AB/N4BEG[6] Tile_X3Y3_LUT4AB/N4BEG[7] Tile_X3Y3_LUT4AB/N4BEG[8]
+ Tile_X3Y3_LUT4AB/N4BEG[9] Tile_X3Y4_LUT4AB/N4BEG[0] Tile_X3Y4_LUT4AB/N4BEG[10] Tile_X3Y4_LUT4AB/N4BEG[11]
+ Tile_X3Y4_LUT4AB/N4BEG[12] Tile_X3Y4_LUT4AB/N4BEG[13] Tile_X3Y4_LUT4AB/N4BEG[14]
+ Tile_X3Y4_LUT4AB/N4BEG[15] Tile_X3Y4_LUT4AB/N4BEG[1] Tile_X3Y4_LUT4AB/N4BEG[2] Tile_X3Y4_LUT4AB/N4BEG[3]
+ Tile_X3Y4_LUT4AB/N4BEG[4] Tile_X3Y4_LUT4AB/N4BEG[5] Tile_X3Y4_LUT4AB/N4BEG[6] Tile_X3Y4_LUT4AB/N4BEG[7]
+ Tile_X3Y4_LUT4AB/N4BEG[8] Tile_X3Y4_LUT4AB/N4BEG[9] Tile_X3Y3_LUT4AB/NN4BEG[0] Tile_X3Y3_LUT4AB/NN4BEG[10]
+ Tile_X3Y3_LUT4AB/NN4BEG[11] Tile_X3Y3_LUT4AB/NN4BEG[12] Tile_X3Y3_LUT4AB/NN4BEG[13]
+ Tile_X3Y3_LUT4AB/NN4BEG[14] Tile_X3Y3_LUT4AB/NN4BEG[15] Tile_X3Y3_LUT4AB/NN4BEG[1]
+ Tile_X3Y3_LUT4AB/NN4BEG[2] Tile_X3Y3_LUT4AB/NN4BEG[3] Tile_X3Y3_LUT4AB/NN4BEG[4]
+ Tile_X3Y3_LUT4AB/NN4BEG[5] Tile_X3Y3_LUT4AB/NN4BEG[6] Tile_X3Y3_LUT4AB/NN4BEG[7]
+ Tile_X3Y3_LUT4AB/NN4BEG[8] Tile_X3Y3_LUT4AB/NN4BEG[9] Tile_X3Y4_LUT4AB/NN4BEG[0]
+ Tile_X3Y4_LUT4AB/NN4BEG[10] Tile_X3Y4_LUT4AB/NN4BEG[11] Tile_X3Y4_LUT4AB/NN4BEG[12]
+ Tile_X3Y4_LUT4AB/NN4BEG[13] Tile_X3Y4_LUT4AB/NN4BEG[14] Tile_X3Y4_LUT4AB/NN4BEG[15]
+ Tile_X3Y4_LUT4AB/NN4BEG[1] Tile_X3Y4_LUT4AB/NN4BEG[2] Tile_X3Y4_LUT4AB/NN4BEG[3]
+ Tile_X3Y4_LUT4AB/NN4BEG[4] Tile_X3Y4_LUT4AB/NN4BEG[5] Tile_X3Y4_LUT4AB/NN4BEG[6]
+ Tile_X3Y4_LUT4AB/NN4BEG[7] Tile_X3Y4_LUT4AB/NN4BEG[8] Tile_X3Y4_LUT4AB/NN4BEG[9]
+ Tile_X3Y4_LUT4AB/S1END[0] Tile_X3Y4_LUT4AB/S1END[1] Tile_X3Y4_LUT4AB/S1END[2] Tile_X3Y4_LUT4AB/S1END[3]
+ Tile_X3Y3_LUT4AB/S1END[0] Tile_X3Y3_LUT4AB/S1END[1] Tile_X3Y3_LUT4AB/S1END[2] Tile_X3Y3_LUT4AB/S1END[3]
+ Tile_X3Y4_LUT4AB/S2MID[0] Tile_X3Y4_LUT4AB/S2MID[1] Tile_X3Y4_LUT4AB/S2MID[2] Tile_X3Y4_LUT4AB/S2MID[3]
+ Tile_X3Y4_LUT4AB/S2MID[4] Tile_X3Y4_LUT4AB/S2MID[5] Tile_X3Y4_LUT4AB/S2MID[6] Tile_X3Y4_LUT4AB/S2MID[7]
+ Tile_X3Y4_LUT4AB/S2END[0] Tile_X3Y4_LUT4AB/S2END[1] Tile_X3Y4_LUT4AB/S2END[2] Tile_X3Y4_LUT4AB/S2END[3]
+ Tile_X3Y4_LUT4AB/S2END[4] Tile_X3Y4_LUT4AB/S2END[5] Tile_X3Y4_LUT4AB/S2END[6] Tile_X3Y4_LUT4AB/S2END[7]
+ Tile_X3Y3_LUT4AB/S2END[0] Tile_X3Y3_LUT4AB/S2END[1] Tile_X3Y3_LUT4AB/S2END[2] Tile_X3Y3_LUT4AB/S2END[3]
+ Tile_X3Y3_LUT4AB/S2END[4] Tile_X3Y3_LUT4AB/S2END[5] Tile_X3Y3_LUT4AB/S2END[6] Tile_X3Y3_LUT4AB/S2END[7]
+ Tile_X3Y3_LUT4AB/S2MID[0] Tile_X3Y3_LUT4AB/S2MID[1] Tile_X3Y3_LUT4AB/S2MID[2] Tile_X3Y3_LUT4AB/S2MID[3]
+ Tile_X3Y3_LUT4AB/S2MID[4] Tile_X3Y3_LUT4AB/S2MID[5] Tile_X3Y3_LUT4AB/S2MID[6] Tile_X3Y3_LUT4AB/S2MID[7]
+ Tile_X3Y4_LUT4AB/S4END[0] Tile_X3Y4_LUT4AB/S4END[10] Tile_X3Y4_LUT4AB/S4END[11]
+ Tile_X3Y4_LUT4AB/S4END[12] Tile_X3Y4_LUT4AB/S4END[13] Tile_X3Y4_LUT4AB/S4END[14]
+ Tile_X3Y4_LUT4AB/S4END[15] Tile_X3Y4_LUT4AB/S4END[1] Tile_X3Y4_LUT4AB/S4END[2] Tile_X3Y4_LUT4AB/S4END[3]
+ Tile_X3Y4_LUT4AB/S4END[4] Tile_X3Y4_LUT4AB/S4END[5] Tile_X3Y4_LUT4AB/S4END[6] Tile_X3Y4_LUT4AB/S4END[7]
+ Tile_X3Y4_LUT4AB/S4END[8] Tile_X3Y4_LUT4AB/S4END[9] Tile_X3Y3_LUT4AB/S4END[0] Tile_X3Y3_LUT4AB/S4END[10]
+ Tile_X3Y3_LUT4AB/S4END[11] Tile_X3Y3_LUT4AB/S4END[12] Tile_X3Y3_LUT4AB/S4END[13]
+ Tile_X3Y3_LUT4AB/S4END[14] Tile_X3Y3_LUT4AB/S4END[15] Tile_X3Y3_LUT4AB/S4END[1]
+ Tile_X3Y3_LUT4AB/S4END[2] Tile_X3Y3_LUT4AB/S4END[3] Tile_X3Y3_LUT4AB/S4END[4] Tile_X3Y3_LUT4AB/S4END[5]
+ Tile_X3Y3_LUT4AB/S4END[6] Tile_X3Y3_LUT4AB/S4END[7] Tile_X3Y3_LUT4AB/S4END[8] Tile_X3Y3_LUT4AB/S4END[9]
+ Tile_X3Y4_LUT4AB/SS4END[0] Tile_X3Y4_LUT4AB/SS4END[10] Tile_X3Y4_LUT4AB/SS4END[11]
+ Tile_X3Y4_LUT4AB/SS4END[12] Tile_X3Y4_LUT4AB/SS4END[13] Tile_X3Y4_LUT4AB/SS4END[14]
+ Tile_X3Y4_LUT4AB/SS4END[15] Tile_X3Y4_LUT4AB/SS4END[1] Tile_X3Y4_LUT4AB/SS4END[2]
+ Tile_X3Y4_LUT4AB/SS4END[3] Tile_X3Y4_LUT4AB/SS4END[4] Tile_X3Y4_LUT4AB/SS4END[5]
+ Tile_X3Y4_LUT4AB/SS4END[6] Tile_X3Y4_LUT4AB/SS4END[7] Tile_X3Y4_LUT4AB/SS4END[8]
+ Tile_X3Y4_LUT4AB/SS4END[9] Tile_X3Y3_LUT4AB/SS4END[0] Tile_X3Y3_LUT4AB/SS4END[10]
+ Tile_X3Y3_LUT4AB/SS4END[11] Tile_X3Y3_LUT4AB/SS4END[12] Tile_X3Y3_LUT4AB/SS4END[13]
+ Tile_X3Y3_LUT4AB/SS4END[14] Tile_X3Y3_LUT4AB/SS4END[15] Tile_X3Y3_LUT4AB/SS4END[1]
+ Tile_X3Y3_LUT4AB/SS4END[2] Tile_X3Y3_LUT4AB/SS4END[3] Tile_X3Y3_LUT4AB/SS4END[4]
+ Tile_X3Y3_LUT4AB/SS4END[5] Tile_X3Y3_LUT4AB/SS4END[6] Tile_X3Y3_LUT4AB/SS4END[7]
+ Tile_X3Y3_LUT4AB/SS4END[8] Tile_X3Y3_LUT4AB/SS4END[9] Tile_X3Y3_LUT4AB/UserCLK Tile_X3Y2_LUT4AB/UserCLK
+ VGND VPWR Tile_X3Y3_LUT4AB/W1BEG[0] Tile_X3Y3_LUT4AB/W1BEG[1] Tile_X3Y3_LUT4AB/W1BEG[2]
+ Tile_X3Y3_LUT4AB/W1BEG[3] Tile_X4Y3_LUT4AB/W1BEG[0] Tile_X4Y3_LUT4AB/W1BEG[1] Tile_X4Y3_LUT4AB/W1BEG[2]
+ Tile_X4Y3_LUT4AB/W1BEG[3] Tile_X3Y3_LUT4AB/W2BEG[0] Tile_X3Y3_LUT4AB/W2BEG[1] Tile_X3Y3_LUT4AB/W2BEG[2]
+ Tile_X3Y3_LUT4AB/W2BEG[3] Tile_X3Y3_LUT4AB/W2BEG[4] Tile_X3Y3_LUT4AB/W2BEG[5] Tile_X3Y3_LUT4AB/W2BEG[6]
+ Tile_X3Y3_LUT4AB/W2BEG[7] Tile_X2Y3_LUT4AB/W2END[0] Tile_X2Y3_LUT4AB/W2END[1] Tile_X2Y3_LUT4AB/W2END[2]
+ Tile_X2Y3_LUT4AB/W2END[3] Tile_X2Y3_LUT4AB/W2END[4] Tile_X2Y3_LUT4AB/W2END[5] Tile_X2Y3_LUT4AB/W2END[6]
+ Tile_X2Y3_LUT4AB/W2END[7] Tile_X3Y3_LUT4AB/W2END[0] Tile_X3Y3_LUT4AB/W2END[1] Tile_X3Y3_LUT4AB/W2END[2]
+ Tile_X3Y3_LUT4AB/W2END[3] Tile_X3Y3_LUT4AB/W2END[4] Tile_X3Y3_LUT4AB/W2END[5] Tile_X3Y3_LUT4AB/W2END[6]
+ Tile_X3Y3_LUT4AB/W2END[7] Tile_X4Y3_LUT4AB/W2BEG[0] Tile_X4Y3_LUT4AB/W2BEG[1] Tile_X4Y3_LUT4AB/W2BEG[2]
+ Tile_X4Y3_LUT4AB/W2BEG[3] Tile_X4Y3_LUT4AB/W2BEG[4] Tile_X4Y3_LUT4AB/W2BEG[5] Tile_X4Y3_LUT4AB/W2BEG[6]
+ Tile_X4Y3_LUT4AB/W2BEG[7] Tile_X3Y3_LUT4AB/W6BEG[0] Tile_X3Y3_LUT4AB/W6BEG[10] Tile_X3Y3_LUT4AB/W6BEG[11]
+ Tile_X3Y3_LUT4AB/W6BEG[1] Tile_X3Y3_LUT4AB/W6BEG[2] Tile_X3Y3_LUT4AB/W6BEG[3] Tile_X3Y3_LUT4AB/W6BEG[4]
+ Tile_X3Y3_LUT4AB/W6BEG[5] Tile_X3Y3_LUT4AB/W6BEG[6] Tile_X3Y3_LUT4AB/W6BEG[7] Tile_X3Y3_LUT4AB/W6BEG[8]
+ Tile_X3Y3_LUT4AB/W6BEG[9] Tile_X4Y3_LUT4AB/W6BEG[0] Tile_X4Y3_LUT4AB/W6BEG[10] Tile_X4Y3_LUT4AB/W6BEG[11]
+ Tile_X4Y3_LUT4AB/W6BEG[1] Tile_X4Y3_LUT4AB/W6BEG[2] Tile_X4Y3_LUT4AB/W6BEG[3] Tile_X4Y3_LUT4AB/W6BEG[4]
+ Tile_X4Y3_LUT4AB/W6BEG[5] Tile_X4Y3_LUT4AB/W6BEG[6] Tile_X4Y3_LUT4AB/W6BEG[7] Tile_X4Y3_LUT4AB/W6BEG[8]
+ Tile_X4Y3_LUT4AB/W6BEG[9] Tile_X3Y3_LUT4AB/WW4BEG[0] Tile_X3Y3_LUT4AB/WW4BEG[10]
+ Tile_X3Y3_LUT4AB/WW4BEG[11] Tile_X3Y3_LUT4AB/WW4BEG[12] Tile_X3Y3_LUT4AB/WW4BEG[13]
+ Tile_X3Y3_LUT4AB/WW4BEG[14] Tile_X3Y3_LUT4AB/WW4BEG[15] Tile_X3Y3_LUT4AB/WW4BEG[1]
+ Tile_X3Y3_LUT4AB/WW4BEG[2] Tile_X3Y3_LUT4AB/WW4BEG[3] Tile_X3Y3_LUT4AB/WW4BEG[4]
+ Tile_X3Y3_LUT4AB/WW4BEG[5] Tile_X3Y3_LUT4AB/WW4BEG[6] Tile_X3Y3_LUT4AB/WW4BEG[7]
+ Tile_X3Y3_LUT4AB/WW4BEG[8] Tile_X3Y3_LUT4AB/WW4BEG[9] Tile_X4Y3_LUT4AB/WW4BEG[0]
+ Tile_X4Y3_LUT4AB/WW4BEG[10] Tile_X4Y3_LUT4AB/WW4BEG[11] Tile_X4Y3_LUT4AB/WW4BEG[12]
+ Tile_X4Y3_LUT4AB/WW4BEG[13] Tile_X4Y3_LUT4AB/WW4BEG[14] Tile_X4Y3_LUT4AB/WW4BEG[15]
+ Tile_X4Y3_LUT4AB/WW4BEG[1] Tile_X4Y3_LUT4AB/WW4BEG[2] Tile_X4Y3_LUT4AB/WW4BEG[3]
+ Tile_X4Y3_LUT4AB/WW4BEG[4] Tile_X4Y3_LUT4AB/WW4BEG[5] Tile_X4Y3_LUT4AB/WW4BEG[6]
+ Tile_X4Y3_LUT4AB/WW4BEG[7] Tile_X4Y3_LUT4AB/WW4BEG[8] Tile_X4Y3_LUT4AB/WW4BEG[9]
+ LUT4AB
XTile_X0Y6_W_TT_IF Tile_X0Y6_CLK_TT_PROJECT Tile_X1Y6_LUT4AB/E1END[0] Tile_X1Y6_LUT4AB/E1END[1]
+ Tile_X1Y6_LUT4AB/E1END[2] Tile_X1Y6_LUT4AB/E1END[3] Tile_X1Y6_LUT4AB/E2MID[0] Tile_X1Y6_LUT4AB/E2MID[1]
+ Tile_X1Y6_LUT4AB/E2MID[2] Tile_X1Y6_LUT4AB/E2MID[3] Tile_X1Y6_LUT4AB/E2MID[4] Tile_X1Y6_LUT4AB/E2MID[5]
+ Tile_X1Y6_LUT4AB/E2MID[6] Tile_X1Y6_LUT4AB/E2MID[7] Tile_X1Y6_LUT4AB/E2END[0] Tile_X1Y6_LUT4AB/E2END[1]
+ Tile_X1Y6_LUT4AB/E2END[2] Tile_X1Y6_LUT4AB/E2END[3] Tile_X1Y6_LUT4AB/E2END[4] Tile_X1Y6_LUT4AB/E2END[5]
+ Tile_X1Y6_LUT4AB/E2END[6] Tile_X1Y6_LUT4AB/E2END[7] Tile_X1Y6_LUT4AB/E6END[0] Tile_X1Y6_LUT4AB/E6END[10]
+ Tile_X1Y6_LUT4AB/E6END[11] Tile_X1Y6_LUT4AB/E6END[1] Tile_X1Y6_LUT4AB/E6END[2] Tile_X1Y6_LUT4AB/E6END[3]
+ Tile_X1Y6_LUT4AB/E6END[4] Tile_X1Y6_LUT4AB/E6END[5] Tile_X1Y6_LUT4AB/E6END[6] Tile_X1Y6_LUT4AB/E6END[7]
+ Tile_X1Y6_LUT4AB/E6END[8] Tile_X1Y6_LUT4AB/E6END[9] Tile_X1Y6_LUT4AB/EE4END[0] Tile_X1Y6_LUT4AB/EE4END[10]
+ Tile_X1Y6_LUT4AB/EE4END[11] Tile_X1Y6_LUT4AB/EE4END[12] Tile_X1Y6_LUT4AB/EE4END[13]
+ Tile_X1Y6_LUT4AB/EE4END[14] Tile_X1Y6_LUT4AB/EE4END[15] Tile_X1Y6_LUT4AB/EE4END[1]
+ Tile_X1Y6_LUT4AB/EE4END[2] Tile_X1Y6_LUT4AB/EE4END[3] Tile_X1Y6_LUT4AB/EE4END[4]
+ Tile_X1Y6_LUT4AB/EE4END[5] Tile_X1Y6_LUT4AB/EE4END[6] Tile_X1Y6_LUT4AB/EE4END[7]
+ Tile_X1Y6_LUT4AB/EE4END[8] Tile_X1Y6_LUT4AB/EE4END[9] Tile_X0Y6_ENA_TT_PROJECT FrameData[192]
+ FrameData[202] FrameData[203] FrameData[204] FrameData[205] FrameData[206] FrameData[207]
+ FrameData[208] FrameData[209] FrameData[210] FrameData[211] FrameData[193] FrameData[212]
+ FrameData[213] FrameData[214] FrameData[215] FrameData[216] FrameData[217] FrameData[218]
+ FrameData[219] FrameData[220] FrameData[221] FrameData[194] FrameData[222] FrameData[223]
+ FrameData[195] FrameData[196] FrameData[197] FrameData[198] FrameData[199] FrameData[200]
+ FrameData[201] Tile_X1Y6_LUT4AB/FrameData[0] Tile_X1Y6_LUT4AB/FrameData[10] Tile_X1Y6_LUT4AB/FrameData[11]
+ Tile_X1Y6_LUT4AB/FrameData[12] Tile_X1Y6_LUT4AB/FrameData[13] Tile_X1Y6_LUT4AB/FrameData[14]
+ Tile_X1Y6_LUT4AB/FrameData[15] Tile_X1Y6_LUT4AB/FrameData[16] Tile_X1Y6_LUT4AB/FrameData[17]
+ Tile_X1Y6_LUT4AB/FrameData[18] Tile_X1Y6_LUT4AB/FrameData[19] Tile_X1Y6_LUT4AB/FrameData[1]
+ Tile_X1Y6_LUT4AB/FrameData[20] Tile_X1Y6_LUT4AB/FrameData[21] Tile_X1Y6_LUT4AB/FrameData[22]
+ Tile_X1Y6_LUT4AB/FrameData[23] Tile_X1Y6_LUT4AB/FrameData[24] Tile_X1Y6_LUT4AB/FrameData[25]
+ Tile_X1Y6_LUT4AB/FrameData[26] Tile_X1Y6_LUT4AB/FrameData[27] Tile_X1Y6_LUT4AB/FrameData[28]
+ Tile_X1Y6_LUT4AB/FrameData[29] Tile_X1Y6_LUT4AB/FrameData[2] Tile_X1Y6_LUT4AB/FrameData[30]
+ Tile_X1Y6_LUT4AB/FrameData[31] Tile_X1Y6_LUT4AB/FrameData[3] Tile_X1Y6_LUT4AB/FrameData[4]
+ Tile_X1Y6_LUT4AB/FrameData[5] Tile_X1Y6_LUT4AB/FrameData[6] Tile_X1Y6_LUT4AB/FrameData[7]
+ Tile_X1Y6_LUT4AB/FrameData[8] Tile_X1Y6_LUT4AB/FrameData[9] Tile_X0Y6_W_TT_IF/FrameStrobe[0]
+ Tile_X0Y6_W_TT_IF/FrameStrobe[10] Tile_X0Y6_W_TT_IF/FrameStrobe[11] Tile_X0Y6_W_TT_IF/FrameStrobe[12]
+ Tile_X0Y6_W_TT_IF/FrameStrobe[13] Tile_X0Y6_W_TT_IF/FrameStrobe[14] Tile_X0Y6_W_TT_IF/FrameStrobe[15]
+ Tile_X0Y6_W_TT_IF/FrameStrobe[16] Tile_X0Y6_W_TT_IF/FrameStrobe[17] Tile_X0Y6_W_TT_IF/FrameStrobe[18]
+ Tile_X0Y6_W_TT_IF/FrameStrobe[19] Tile_X0Y6_W_TT_IF/FrameStrobe[1] Tile_X0Y6_W_TT_IF/FrameStrobe[2]
+ Tile_X0Y6_W_TT_IF/FrameStrobe[3] Tile_X0Y6_W_TT_IF/FrameStrobe[4] Tile_X0Y6_W_TT_IF/FrameStrobe[5]
+ Tile_X0Y6_W_TT_IF/FrameStrobe[6] Tile_X0Y6_W_TT_IF/FrameStrobe[7] Tile_X0Y6_W_TT_IF/FrameStrobe[8]
+ Tile_X0Y6_W_TT_IF/FrameStrobe[9] Tile_X0Y5_W_TT_IF/FrameStrobe[0] Tile_X0Y5_W_TT_IF/FrameStrobe[10]
+ Tile_X0Y5_W_TT_IF/FrameStrobe[11] Tile_X0Y5_W_TT_IF/FrameStrobe[12] Tile_X0Y5_W_TT_IF/FrameStrobe[13]
+ Tile_X0Y5_W_TT_IF/FrameStrobe[14] Tile_X0Y5_W_TT_IF/FrameStrobe[15] Tile_X0Y5_W_TT_IF/FrameStrobe[16]
+ Tile_X0Y5_W_TT_IF/FrameStrobe[17] Tile_X0Y5_W_TT_IF/FrameStrobe[18] Tile_X0Y5_W_TT_IF/FrameStrobe[19]
+ Tile_X0Y5_W_TT_IF/FrameStrobe[1] Tile_X0Y5_W_TT_IF/FrameStrobe[2] Tile_X0Y5_W_TT_IF/FrameStrobe[3]
+ Tile_X0Y5_W_TT_IF/FrameStrobe[4] Tile_X0Y5_W_TT_IF/FrameStrobe[5] Tile_X0Y5_W_TT_IF/FrameStrobe[6]
+ Tile_X0Y5_W_TT_IF/FrameStrobe[7] Tile_X0Y5_W_TT_IF/FrameStrobe[8] Tile_X0Y5_W_TT_IF/FrameStrobe[9]
+ Tile_X0Y6_W_TT_IF/N1BEG[0] Tile_X0Y6_W_TT_IF/N1BEG[1] Tile_X0Y6_W_TT_IF/N1BEG[2]
+ Tile_X0Y6_W_TT_IF/N1BEG[3] Tile_X0Y7_W_TT_IF/N1BEG[0] Tile_X0Y7_W_TT_IF/N1BEG[1]
+ Tile_X0Y7_W_TT_IF/N1BEG[2] Tile_X0Y7_W_TT_IF/N1BEG[3] Tile_X0Y6_W_TT_IF/N2BEG[0]
+ Tile_X0Y6_W_TT_IF/N2BEG[1] Tile_X0Y6_W_TT_IF/N2BEG[2] Tile_X0Y6_W_TT_IF/N2BEG[3]
+ Tile_X0Y6_W_TT_IF/N2BEG[4] Tile_X0Y6_W_TT_IF/N2BEG[5] Tile_X0Y6_W_TT_IF/N2BEG[6]
+ Tile_X0Y6_W_TT_IF/N2BEG[7] Tile_X0Y5_W_TT_IF/N2END[0] Tile_X0Y5_W_TT_IF/N2END[1]
+ Tile_X0Y5_W_TT_IF/N2END[2] Tile_X0Y5_W_TT_IF/N2END[3] Tile_X0Y5_W_TT_IF/N2END[4]
+ Tile_X0Y5_W_TT_IF/N2END[5] Tile_X0Y5_W_TT_IF/N2END[6] Tile_X0Y5_W_TT_IF/N2END[7]
+ Tile_X0Y6_W_TT_IF/N2END[0] Tile_X0Y6_W_TT_IF/N2END[1] Tile_X0Y6_W_TT_IF/N2END[2]
+ Tile_X0Y6_W_TT_IF/N2END[3] Tile_X0Y6_W_TT_IF/N2END[4] Tile_X0Y6_W_TT_IF/N2END[5]
+ Tile_X0Y6_W_TT_IF/N2END[6] Tile_X0Y6_W_TT_IF/N2END[7] Tile_X0Y7_W_TT_IF/N2BEG[0]
+ Tile_X0Y7_W_TT_IF/N2BEG[1] Tile_X0Y7_W_TT_IF/N2BEG[2] Tile_X0Y7_W_TT_IF/N2BEG[3]
+ Tile_X0Y7_W_TT_IF/N2BEG[4] Tile_X0Y7_W_TT_IF/N2BEG[5] Tile_X0Y7_W_TT_IF/N2BEG[6]
+ Tile_X0Y7_W_TT_IF/N2BEG[7] Tile_X0Y6_W_TT_IF/N4BEG[0] Tile_X0Y6_W_TT_IF/N4BEG[10]
+ Tile_X0Y6_W_TT_IF/N4BEG[11] Tile_X0Y6_W_TT_IF/N4BEG[12] Tile_X0Y6_W_TT_IF/N4BEG[13]
+ Tile_X0Y6_W_TT_IF/N4BEG[14] Tile_X0Y6_W_TT_IF/N4BEG[15] Tile_X0Y6_W_TT_IF/N4BEG[1]
+ Tile_X0Y6_W_TT_IF/N4BEG[2] Tile_X0Y6_W_TT_IF/N4BEG[3] Tile_X0Y6_W_TT_IF/N4BEG[4]
+ Tile_X0Y6_W_TT_IF/N4BEG[5] Tile_X0Y6_W_TT_IF/N4BEG[6] Tile_X0Y6_W_TT_IF/N4BEG[7]
+ Tile_X0Y6_W_TT_IF/N4BEG[8] Tile_X0Y6_W_TT_IF/N4BEG[9] Tile_X0Y7_W_TT_IF/N4BEG[0]
+ Tile_X0Y7_W_TT_IF/N4BEG[10] Tile_X0Y7_W_TT_IF/N4BEG[11] Tile_X0Y7_W_TT_IF/N4BEG[12]
+ Tile_X0Y7_W_TT_IF/N4BEG[13] Tile_X0Y7_W_TT_IF/N4BEG[14] Tile_X0Y7_W_TT_IF/N4BEG[15]
+ Tile_X0Y7_W_TT_IF/N4BEG[1] Tile_X0Y7_W_TT_IF/N4BEG[2] Tile_X0Y7_W_TT_IF/N4BEG[3]
+ Tile_X0Y7_W_TT_IF/N4BEG[4] Tile_X0Y7_W_TT_IF/N4BEG[5] Tile_X0Y7_W_TT_IF/N4BEG[6]
+ Tile_X0Y7_W_TT_IF/N4BEG[7] Tile_X0Y7_W_TT_IF/N4BEG[8] Tile_X0Y7_W_TT_IF/N4BEG[9]
+ Tile_X0Y6_RST_N_TT_PROJECT Tile_X0Y7_W_TT_IF/S1END[0] Tile_X0Y7_W_TT_IF/S1END[1]
+ Tile_X0Y7_W_TT_IF/S1END[2] Tile_X0Y7_W_TT_IF/S1END[3] Tile_X0Y6_W_TT_IF/S1END[0]
+ Tile_X0Y6_W_TT_IF/S1END[1] Tile_X0Y6_W_TT_IF/S1END[2] Tile_X0Y6_W_TT_IF/S1END[3]
+ Tile_X0Y7_W_TT_IF/S2MID[0] Tile_X0Y7_W_TT_IF/S2MID[1] Tile_X0Y7_W_TT_IF/S2MID[2]
+ Tile_X0Y7_W_TT_IF/S2MID[3] Tile_X0Y7_W_TT_IF/S2MID[4] Tile_X0Y7_W_TT_IF/S2MID[5]
+ Tile_X0Y7_W_TT_IF/S2MID[6] Tile_X0Y7_W_TT_IF/S2MID[7] Tile_X0Y7_W_TT_IF/S2END[0]
+ Tile_X0Y7_W_TT_IF/S2END[1] Tile_X0Y7_W_TT_IF/S2END[2] Tile_X0Y7_W_TT_IF/S2END[3]
+ Tile_X0Y7_W_TT_IF/S2END[4] Tile_X0Y7_W_TT_IF/S2END[5] Tile_X0Y7_W_TT_IF/S2END[6]
+ Tile_X0Y7_W_TT_IF/S2END[7] Tile_X0Y6_W_TT_IF/S2END[0] Tile_X0Y6_W_TT_IF/S2END[1]
+ Tile_X0Y6_W_TT_IF/S2END[2] Tile_X0Y6_W_TT_IF/S2END[3] Tile_X0Y6_W_TT_IF/S2END[4]
+ Tile_X0Y6_W_TT_IF/S2END[5] Tile_X0Y6_W_TT_IF/S2END[6] Tile_X0Y6_W_TT_IF/S2END[7]
+ Tile_X0Y6_W_TT_IF/S2MID[0] Tile_X0Y6_W_TT_IF/S2MID[1] Tile_X0Y6_W_TT_IF/S2MID[2]
+ Tile_X0Y6_W_TT_IF/S2MID[3] Tile_X0Y6_W_TT_IF/S2MID[4] Tile_X0Y6_W_TT_IF/S2MID[5]
+ Tile_X0Y6_W_TT_IF/S2MID[6] Tile_X0Y6_W_TT_IF/S2MID[7] Tile_X0Y7_W_TT_IF/S4END[0]
+ Tile_X0Y7_W_TT_IF/S4END[10] Tile_X0Y7_W_TT_IF/S4END[11] Tile_X0Y7_W_TT_IF/S4END[12]
+ Tile_X0Y7_W_TT_IF/S4END[13] Tile_X0Y7_W_TT_IF/S4END[14] Tile_X0Y7_W_TT_IF/S4END[15]
+ Tile_X0Y7_W_TT_IF/S4END[1] Tile_X0Y7_W_TT_IF/S4END[2] Tile_X0Y7_W_TT_IF/S4END[3]
+ Tile_X0Y7_W_TT_IF/S4END[4] Tile_X0Y7_W_TT_IF/S4END[5] Tile_X0Y7_W_TT_IF/S4END[6]
+ Tile_X0Y7_W_TT_IF/S4END[7] Tile_X0Y7_W_TT_IF/S4END[8] Tile_X0Y7_W_TT_IF/S4END[9]
+ Tile_X0Y6_W_TT_IF/S4END[0] Tile_X0Y6_W_TT_IF/S4END[10] Tile_X0Y6_W_TT_IF/S4END[11]
+ Tile_X0Y6_W_TT_IF/S4END[12] Tile_X0Y6_W_TT_IF/S4END[13] Tile_X0Y6_W_TT_IF/S4END[14]
+ Tile_X0Y6_W_TT_IF/S4END[15] Tile_X0Y6_W_TT_IF/S4END[1] Tile_X0Y6_W_TT_IF/S4END[2]
+ Tile_X0Y6_W_TT_IF/S4END[3] Tile_X0Y6_W_TT_IF/S4END[4] Tile_X0Y6_W_TT_IF/S4END[5]
+ Tile_X0Y6_W_TT_IF/S4END[6] Tile_X0Y6_W_TT_IF/S4END[7] Tile_X0Y6_W_TT_IF/S4END[8]
+ Tile_X0Y6_W_TT_IF/S4END[9] Tile_X0Y6_UIO_IN_TT_PROJECT0 Tile_X0Y6_UIO_IN_TT_PROJECT1
+ Tile_X0Y6_UIO_IN_TT_PROJECT2 Tile_X0Y6_UIO_IN_TT_PROJECT3 Tile_X0Y6_UIO_IN_TT_PROJECT4
+ Tile_X0Y6_UIO_IN_TT_PROJECT5 Tile_X0Y6_UIO_IN_TT_PROJECT6 Tile_X0Y6_UIO_IN_TT_PROJECT7
+ Tile_X0Y6_UIO_OE_TT_PROJECT0 Tile_X0Y6_UIO_OE_TT_PROJECT1 Tile_X0Y6_UIO_OE_TT_PROJECT2
+ Tile_X0Y6_UIO_OE_TT_PROJECT3 Tile_X0Y6_UIO_OE_TT_PROJECT4 Tile_X0Y6_UIO_OE_TT_PROJECT5
+ Tile_X0Y6_UIO_OE_TT_PROJECT6 Tile_X0Y6_UIO_OE_TT_PROJECT7 Tile_X0Y6_UIO_OUT_TT_PROJECT0
+ Tile_X0Y6_UIO_OUT_TT_PROJECT1 Tile_X0Y6_UIO_OUT_TT_PROJECT2 Tile_X0Y6_UIO_OUT_TT_PROJECT3
+ Tile_X0Y6_UIO_OUT_TT_PROJECT4 Tile_X0Y6_UIO_OUT_TT_PROJECT5 Tile_X0Y6_UIO_OUT_TT_PROJECT6
+ Tile_X0Y6_UIO_OUT_TT_PROJECT7 Tile_X0Y6_UI_IN_TT_PROJECT0 Tile_X0Y6_UI_IN_TT_PROJECT1
+ Tile_X0Y6_UI_IN_TT_PROJECT2 Tile_X0Y6_UI_IN_TT_PROJECT3 Tile_X0Y6_UI_IN_TT_PROJECT4
+ Tile_X0Y6_UI_IN_TT_PROJECT5 Tile_X0Y6_UI_IN_TT_PROJECT6 Tile_X0Y6_UI_IN_TT_PROJECT7
+ Tile_X0Y6_UO_OUT_TT_PROJECT0 Tile_X0Y6_UO_OUT_TT_PROJECT1 Tile_X0Y6_UO_OUT_TT_PROJECT2
+ Tile_X0Y6_UO_OUT_TT_PROJECT3 Tile_X0Y6_UO_OUT_TT_PROJECT4 Tile_X0Y6_UO_OUT_TT_PROJECT5
+ Tile_X0Y6_UO_OUT_TT_PROJECT6 Tile_X0Y6_UO_OUT_TT_PROJECT7 Tile_X0Y6_W_TT_IF/UserCLK
+ Tile_X0Y5_W_TT_IF/UserCLK VGND VPWR Tile_X1Y6_LUT4AB/W1BEG[0] Tile_X1Y6_LUT4AB/W1BEG[1]
+ Tile_X1Y6_LUT4AB/W1BEG[2] Tile_X1Y6_LUT4AB/W1BEG[3] Tile_X1Y6_LUT4AB/W2BEGb[0] Tile_X1Y6_LUT4AB/W2BEGb[1]
+ Tile_X1Y6_LUT4AB/W2BEGb[2] Tile_X1Y6_LUT4AB/W2BEGb[3] Tile_X1Y6_LUT4AB/W2BEGb[4]
+ Tile_X1Y6_LUT4AB/W2BEGb[5] Tile_X1Y6_LUT4AB/W2BEGb[6] Tile_X1Y6_LUT4AB/W2BEGb[7]
+ Tile_X1Y6_LUT4AB/W2BEG[0] Tile_X1Y6_LUT4AB/W2BEG[1] Tile_X1Y6_LUT4AB/W2BEG[2] Tile_X1Y6_LUT4AB/W2BEG[3]
+ Tile_X1Y6_LUT4AB/W2BEG[4] Tile_X1Y6_LUT4AB/W2BEG[5] Tile_X1Y6_LUT4AB/W2BEG[6] Tile_X1Y6_LUT4AB/W2BEG[7]
+ Tile_X1Y6_LUT4AB/W6BEG[0] Tile_X1Y6_LUT4AB/W6BEG[10] Tile_X1Y6_LUT4AB/W6BEG[11]
+ Tile_X1Y6_LUT4AB/W6BEG[1] Tile_X1Y6_LUT4AB/W6BEG[2] Tile_X1Y6_LUT4AB/W6BEG[3] Tile_X1Y6_LUT4AB/W6BEG[4]
+ Tile_X1Y6_LUT4AB/W6BEG[5] Tile_X1Y6_LUT4AB/W6BEG[6] Tile_X1Y6_LUT4AB/W6BEG[7] Tile_X1Y6_LUT4AB/W6BEG[8]
+ Tile_X1Y6_LUT4AB/W6BEG[9] Tile_X1Y6_LUT4AB/WW4BEG[0] Tile_X1Y6_LUT4AB/WW4BEG[10]
+ Tile_X1Y6_LUT4AB/WW4BEG[11] Tile_X1Y6_LUT4AB/WW4BEG[12] Tile_X1Y6_LUT4AB/WW4BEG[13]
+ Tile_X1Y6_LUT4AB/WW4BEG[14] Tile_X1Y6_LUT4AB/WW4BEG[15] Tile_X1Y6_LUT4AB/WW4BEG[1]
+ Tile_X1Y6_LUT4AB/WW4BEG[2] Tile_X1Y6_LUT4AB/WW4BEG[3] Tile_X1Y6_LUT4AB/WW4BEG[4]
+ Tile_X1Y6_LUT4AB/WW4BEG[5] Tile_X1Y6_LUT4AB/WW4BEG[6] Tile_X1Y6_LUT4AB/WW4BEG[7]
+ Tile_X1Y6_LUT4AB/WW4BEG[8] Tile_X1Y6_LUT4AB/WW4BEG[9] W_TT_IF
XTile_X2Y7_LUT4AB Tile_X2Y8_LUT4AB/Co Tile_X2Y7_LUT4AB/Co Tile_X3Y7_LUT4AB/E1END[0]
+ Tile_X3Y7_LUT4AB/E1END[1] Tile_X3Y7_LUT4AB/E1END[2] Tile_X3Y7_LUT4AB/E1END[3] Tile_X2Y7_LUT4AB/E1END[0]
+ Tile_X2Y7_LUT4AB/E1END[1] Tile_X2Y7_LUT4AB/E1END[2] Tile_X2Y7_LUT4AB/E1END[3] Tile_X3Y7_LUT4AB/E2MID[0]
+ Tile_X3Y7_LUT4AB/E2MID[1] Tile_X3Y7_LUT4AB/E2MID[2] Tile_X3Y7_LUT4AB/E2MID[3] Tile_X3Y7_LUT4AB/E2MID[4]
+ Tile_X3Y7_LUT4AB/E2MID[5] Tile_X3Y7_LUT4AB/E2MID[6] Tile_X3Y7_LUT4AB/E2MID[7] Tile_X3Y7_LUT4AB/E2END[0]
+ Tile_X3Y7_LUT4AB/E2END[1] Tile_X3Y7_LUT4AB/E2END[2] Tile_X3Y7_LUT4AB/E2END[3] Tile_X3Y7_LUT4AB/E2END[4]
+ Tile_X3Y7_LUT4AB/E2END[5] Tile_X3Y7_LUT4AB/E2END[6] Tile_X3Y7_LUT4AB/E2END[7] Tile_X2Y7_LUT4AB/E2END[0]
+ Tile_X2Y7_LUT4AB/E2END[1] Tile_X2Y7_LUT4AB/E2END[2] Tile_X2Y7_LUT4AB/E2END[3] Tile_X2Y7_LUT4AB/E2END[4]
+ Tile_X2Y7_LUT4AB/E2END[5] Tile_X2Y7_LUT4AB/E2END[6] Tile_X2Y7_LUT4AB/E2END[7] Tile_X2Y7_LUT4AB/E2MID[0]
+ Tile_X2Y7_LUT4AB/E2MID[1] Tile_X2Y7_LUT4AB/E2MID[2] Tile_X2Y7_LUT4AB/E2MID[3] Tile_X2Y7_LUT4AB/E2MID[4]
+ Tile_X2Y7_LUT4AB/E2MID[5] Tile_X2Y7_LUT4AB/E2MID[6] Tile_X2Y7_LUT4AB/E2MID[7] Tile_X3Y7_LUT4AB/E6END[0]
+ Tile_X3Y7_LUT4AB/E6END[10] Tile_X3Y7_LUT4AB/E6END[11] Tile_X3Y7_LUT4AB/E6END[1]
+ Tile_X3Y7_LUT4AB/E6END[2] Tile_X3Y7_LUT4AB/E6END[3] Tile_X3Y7_LUT4AB/E6END[4] Tile_X3Y7_LUT4AB/E6END[5]
+ Tile_X3Y7_LUT4AB/E6END[6] Tile_X3Y7_LUT4AB/E6END[7] Tile_X3Y7_LUT4AB/E6END[8] Tile_X3Y7_LUT4AB/E6END[9]
+ Tile_X2Y7_LUT4AB/E6END[0] Tile_X2Y7_LUT4AB/E6END[10] Tile_X2Y7_LUT4AB/E6END[11]
+ Tile_X2Y7_LUT4AB/E6END[1] Tile_X2Y7_LUT4AB/E6END[2] Tile_X2Y7_LUT4AB/E6END[3] Tile_X2Y7_LUT4AB/E6END[4]
+ Tile_X2Y7_LUT4AB/E6END[5] Tile_X2Y7_LUT4AB/E6END[6] Tile_X2Y7_LUT4AB/E6END[7] Tile_X2Y7_LUT4AB/E6END[8]
+ Tile_X2Y7_LUT4AB/E6END[9] Tile_X3Y7_LUT4AB/EE4END[0] Tile_X3Y7_LUT4AB/EE4END[10]
+ Tile_X3Y7_LUT4AB/EE4END[11] Tile_X3Y7_LUT4AB/EE4END[12] Tile_X3Y7_LUT4AB/EE4END[13]
+ Tile_X3Y7_LUT4AB/EE4END[14] Tile_X3Y7_LUT4AB/EE4END[15] Tile_X3Y7_LUT4AB/EE4END[1]
+ Tile_X3Y7_LUT4AB/EE4END[2] Tile_X3Y7_LUT4AB/EE4END[3] Tile_X3Y7_LUT4AB/EE4END[4]
+ Tile_X3Y7_LUT4AB/EE4END[5] Tile_X3Y7_LUT4AB/EE4END[6] Tile_X3Y7_LUT4AB/EE4END[7]
+ Tile_X3Y7_LUT4AB/EE4END[8] Tile_X3Y7_LUT4AB/EE4END[9] Tile_X2Y7_LUT4AB/EE4END[0]
+ Tile_X2Y7_LUT4AB/EE4END[10] Tile_X2Y7_LUT4AB/EE4END[11] Tile_X2Y7_LUT4AB/EE4END[12]
+ Tile_X2Y7_LUT4AB/EE4END[13] Tile_X2Y7_LUT4AB/EE4END[14] Tile_X2Y7_LUT4AB/EE4END[15]
+ Tile_X2Y7_LUT4AB/EE4END[1] Tile_X2Y7_LUT4AB/EE4END[2] Tile_X2Y7_LUT4AB/EE4END[3]
+ Tile_X2Y7_LUT4AB/EE4END[4] Tile_X2Y7_LUT4AB/EE4END[5] Tile_X2Y7_LUT4AB/EE4END[6]
+ Tile_X2Y7_LUT4AB/EE4END[7] Tile_X2Y7_LUT4AB/EE4END[8] Tile_X2Y7_LUT4AB/EE4END[9]
+ Tile_X2Y7_LUT4AB/FrameData[0] Tile_X2Y7_LUT4AB/FrameData[10] Tile_X2Y7_LUT4AB/FrameData[11]
+ Tile_X2Y7_LUT4AB/FrameData[12] Tile_X2Y7_LUT4AB/FrameData[13] Tile_X2Y7_LUT4AB/FrameData[14]
+ Tile_X2Y7_LUT4AB/FrameData[15] Tile_X2Y7_LUT4AB/FrameData[16] Tile_X2Y7_LUT4AB/FrameData[17]
+ Tile_X2Y7_LUT4AB/FrameData[18] Tile_X2Y7_LUT4AB/FrameData[19] Tile_X2Y7_LUT4AB/FrameData[1]
+ Tile_X2Y7_LUT4AB/FrameData[20] Tile_X2Y7_LUT4AB/FrameData[21] Tile_X2Y7_LUT4AB/FrameData[22]
+ Tile_X2Y7_LUT4AB/FrameData[23] Tile_X2Y7_LUT4AB/FrameData[24] Tile_X2Y7_LUT4AB/FrameData[25]
+ Tile_X2Y7_LUT4AB/FrameData[26] Tile_X2Y7_LUT4AB/FrameData[27] Tile_X2Y7_LUT4AB/FrameData[28]
+ Tile_X2Y7_LUT4AB/FrameData[29] Tile_X2Y7_LUT4AB/FrameData[2] Tile_X2Y7_LUT4AB/FrameData[30]
+ Tile_X2Y7_LUT4AB/FrameData[31] Tile_X2Y7_LUT4AB/FrameData[3] Tile_X2Y7_LUT4AB/FrameData[4]
+ Tile_X2Y7_LUT4AB/FrameData[5] Tile_X2Y7_LUT4AB/FrameData[6] Tile_X2Y7_LUT4AB/FrameData[7]
+ Tile_X2Y7_LUT4AB/FrameData[8] Tile_X2Y7_LUT4AB/FrameData[9] Tile_X3Y7_LUT4AB/FrameData[0]
+ Tile_X3Y7_LUT4AB/FrameData[10] Tile_X3Y7_LUT4AB/FrameData[11] Tile_X3Y7_LUT4AB/FrameData[12]
+ Tile_X3Y7_LUT4AB/FrameData[13] Tile_X3Y7_LUT4AB/FrameData[14] Tile_X3Y7_LUT4AB/FrameData[15]
+ Tile_X3Y7_LUT4AB/FrameData[16] Tile_X3Y7_LUT4AB/FrameData[17] Tile_X3Y7_LUT4AB/FrameData[18]
+ Tile_X3Y7_LUT4AB/FrameData[19] Tile_X3Y7_LUT4AB/FrameData[1] Tile_X3Y7_LUT4AB/FrameData[20]
+ Tile_X3Y7_LUT4AB/FrameData[21] Tile_X3Y7_LUT4AB/FrameData[22] Tile_X3Y7_LUT4AB/FrameData[23]
+ Tile_X3Y7_LUT4AB/FrameData[24] Tile_X3Y7_LUT4AB/FrameData[25] Tile_X3Y7_LUT4AB/FrameData[26]
+ Tile_X3Y7_LUT4AB/FrameData[27] Tile_X3Y7_LUT4AB/FrameData[28] Tile_X3Y7_LUT4AB/FrameData[29]
+ Tile_X3Y7_LUT4AB/FrameData[2] Tile_X3Y7_LUT4AB/FrameData[30] Tile_X3Y7_LUT4AB/FrameData[31]
+ Tile_X3Y7_LUT4AB/FrameData[3] Tile_X3Y7_LUT4AB/FrameData[4] Tile_X3Y7_LUT4AB/FrameData[5]
+ Tile_X3Y7_LUT4AB/FrameData[6] Tile_X3Y7_LUT4AB/FrameData[7] Tile_X3Y7_LUT4AB/FrameData[8]
+ Tile_X3Y7_LUT4AB/FrameData[9] Tile_X2Y7_LUT4AB/FrameStrobe[0] Tile_X2Y7_LUT4AB/FrameStrobe[10]
+ Tile_X2Y7_LUT4AB/FrameStrobe[11] Tile_X2Y7_LUT4AB/FrameStrobe[12] Tile_X2Y7_LUT4AB/FrameStrobe[13]
+ Tile_X2Y7_LUT4AB/FrameStrobe[14] Tile_X2Y7_LUT4AB/FrameStrobe[15] Tile_X2Y7_LUT4AB/FrameStrobe[16]
+ Tile_X2Y7_LUT4AB/FrameStrobe[17] Tile_X2Y7_LUT4AB/FrameStrobe[18] Tile_X2Y7_LUT4AB/FrameStrobe[19]
+ Tile_X2Y7_LUT4AB/FrameStrobe[1] Tile_X2Y7_LUT4AB/FrameStrobe[2] Tile_X2Y7_LUT4AB/FrameStrobe[3]
+ Tile_X2Y7_LUT4AB/FrameStrobe[4] Tile_X2Y7_LUT4AB/FrameStrobe[5] Tile_X2Y7_LUT4AB/FrameStrobe[6]
+ Tile_X2Y7_LUT4AB/FrameStrobe[7] Tile_X2Y7_LUT4AB/FrameStrobe[8] Tile_X2Y7_LUT4AB/FrameStrobe[9]
+ Tile_X2Y6_LUT4AB/FrameStrobe[0] Tile_X2Y6_LUT4AB/FrameStrobe[10] Tile_X2Y6_LUT4AB/FrameStrobe[11]
+ Tile_X2Y6_LUT4AB/FrameStrobe[12] Tile_X2Y6_LUT4AB/FrameStrobe[13] Tile_X2Y6_LUT4AB/FrameStrobe[14]
+ Tile_X2Y6_LUT4AB/FrameStrobe[15] Tile_X2Y6_LUT4AB/FrameStrobe[16] Tile_X2Y6_LUT4AB/FrameStrobe[17]
+ Tile_X2Y6_LUT4AB/FrameStrobe[18] Tile_X2Y6_LUT4AB/FrameStrobe[19] Tile_X2Y6_LUT4AB/FrameStrobe[1]
+ Tile_X2Y6_LUT4AB/FrameStrobe[2] Tile_X2Y6_LUT4AB/FrameStrobe[3] Tile_X2Y6_LUT4AB/FrameStrobe[4]
+ Tile_X2Y6_LUT4AB/FrameStrobe[5] Tile_X2Y6_LUT4AB/FrameStrobe[6] Tile_X2Y6_LUT4AB/FrameStrobe[7]
+ Tile_X2Y6_LUT4AB/FrameStrobe[8] Tile_X2Y6_LUT4AB/FrameStrobe[9] Tile_X2Y7_LUT4AB/N1BEG[0]
+ Tile_X2Y7_LUT4AB/N1BEG[1] Tile_X2Y7_LUT4AB/N1BEG[2] Tile_X2Y7_LUT4AB/N1BEG[3] Tile_X2Y8_LUT4AB/N1BEG[0]
+ Tile_X2Y8_LUT4AB/N1BEG[1] Tile_X2Y8_LUT4AB/N1BEG[2] Tile_X2Y8_LUT4AB/N1BEG[3] Tile_X2Y7_LUT4AB/N2BEG[0]
+ Tile_X2Y7_LUT4AB/N2BEG[1] Tile_X2Y7_LUT4AB/N2BEG[2] Tile_X2Y7_LUT4AB/N2BEG[3] Tile_X2Y7_LUT4AB/N2BEG[4]
+ Tile_X2Y7_LUT4AB/N2BEG[5] Tile_X2Y7_LUT4AB/N2BEG[6] Tile_X2Y7_LUT4AB/N2BEG[7] Tile_X2Y6_LUT4AB/N2END[0]
+ Tile_X2Y6_LUT4AB/N2END[1] Tile_X2Y6_LUT4AB/N2END[2] Tile_X2Y6_LUT4AB/N2END[3] Tile_X2Y6_LUT4AB/N2END[4]
+ Tile_X2Y6_LUT4AB/N2END[5] Tile_X2Y6_LUT4AB/N2END[6] Tile_X2Y6_LUT4AB/N2END[7] Tile_X2Y7_LUT4AB/N2END[0]
+ Tile_X2Y7_LUT4AB/N2END[1] Tile_X2Y7_LUT4AB/N2END[2] Tile_X2Y7_LUT4AB/N2END[3] Tile_X2Y7_LUT4AB/N2END[4]
+ Tile_X2Y7_LUT4AB/N2END[5] Tile_X2Y7_LUT4AB/N2END[6] Tile_X2Y7_LUT4AB/N2END[7] Tile_X2Y8_LUT4AB/N2BEG[0]
+ Tile_X2Y8_LUT4AB/N2BEG[1] Tile_X2Y8_LUT4AB/N2BEG[2] Tile_X2Y8_LUT4AB/N2BEG[3] Tile_X2Y8_LUT4AB/N2BEG[4]
+ Tile_X2Y8_LUT4AB/N2BEG[5] Tile_X2Y8_LUT4AB/N2BEG[6] Tile_X2Y8_LUT4AB/N2BEG[7] Tile_X2Y7_LUT4AB/N4BEG[0]
+ Tile_X2Y7_LUT4AB/N4BEG[10] Tile_X2Y7_LUT4AB/N4BEG[11] Tile_X2Y7_LUT4AB/N4BEG[12]
+ Tile_X2Y7_LUT4AB/N4BEG[13] Tile_X2Y7_LUT4AB/N4BEG[14] Tile_X2Y7_LUT4AB/N4BEG[15]
+ Tile_X2Y7_LUT4AB/N4BEG[1] Tile_X2Y7_LUT4AB/N4BEG[2] Tile_X2Y7_LUT4AB/N4BEG[3] Tile_X2Y7_LUT4AB/N4BEG[4]
+ Tile_X2Y7_LUT4AB/N4BEG[5] Tile_X2Y7_LUT4AB/N4BEG[6] Tile_X2Y7_LUT4AB/N4BEG[7] Tile_X2Y7_LUT4AB/N4BEG[8]
+ Tile_X2Y7_LUT4AB/N4BEG[9] Tile_X2Y8_LUT4AB/N4BEG[0] Tile_X2Y8_LUT4AB/N4BEG[10] Tile_X2Y8_LUT4AB/N4BEG[11]
+ Tile_X2Y8_LUT4AB/N4BEG[12] Tile_X2Y8_LUT4AB/N4BEG[13] Tile_X2Y8_LUT4AB/N4BEG[14]
+ Tile_X2Y8_LUT4AB/N4BEG[15] Tile_X2Y8_LUT4AB/N4BEG[1] Tile_X2Y8_LUT4AB/N4BEG[2] Tile_X2Y8_LUT4AB/N4BEG[3]
+ Tile_X2Y8_LUT4AB/N4BEG[4] Tile_X2Y8_LUT4AB/N4BEG[5] Tile_X2Y8_LUT4AB/N4BEG[6] Tile_X2Y8_LUT4AB/N4BEG[7]
+ Tile_X2Y8_LUT4AB/N4BEG[8] Tile_X2Y8_LUT4AB/N4BEG[9] Tile_X2Y7_LUT4AB/NN4BEG[0] Tile_X2Y7_LUT4AB/NN4BEG[10]
+ Tile_X2Y7_LUT4AB/NN4BEG[11] Tile_X2Y7_LUT4AB/NN4BEG[12] Tile_X2Y7_LUT4AB/NN4BEG[13]
+ Tile_X2Y7_LUT4AB/NN4BEG[14] Tile_X2Y7_LUT4AB/NN4BEG[15] Tile_X2Y7_LUT4AB/NN4BEG[1]
+ Tile_X2Y7_LUT4AB/NN4BEG[2] Tile_X2Y7_LUT4AB/NN4BEG[3] Tile_X2Y7_LUT4AB/NN4BEG[4]
+ Tile_X2Y7_LUT4AB/NN4BEG[5] Tile_X2Y7_LUT4AB/NN4BEG[6] Tile_X2Y7_LUT4AB/NN4BEG[7]
+ Tile_X2Y7_LUT4AB/NN4BEG[8] Tile_X2Y7_LUT4AB/NN4BEG[9] Tile_X2Y8_LUT4AB/NN4BEG[0]
+ Tile_X2Y8_LUT4AB/NN4BEG[10] Tile_X2Y8_LUT4AB/NN4BEG[11] Tile_X2Y8_LUT4AB/NN4BEG[12]
+ Tile_X2Y8_LUT4AB/NN4BEG[13] Tile_X2Y8_LUT4AB/NN4BEG[14] Tile_X2Y8_LUT4AB/NN4BEG[15]
+ Tile_X2Y8_LUT4AB/NN4BEG[1] Tile_X2Y8_LUT4AB/NN4BEG[2] Tile_X2Y8_LUT4AB/NN4BEG[3]
+ Tile_X2Y8_LUT4AB/NN4BEG[4] Tile_X2Y8_LUT4AB/NN4BEG[5] Tile_X2Y8_LUT4AB/NN4BEG[6]
+ Tile_X2Y8_LUT4AB/NN4BEG[7] Tile_X2Y8_LUT4AB/NN4BEG[8] Tile_X2Y8_LUT4AB/NN4BEG[9]
+ Tile_X2Y8_LUT4AB/S1END[0] Tile_X2Y8_LUT4AB/S1END[1] Tile_X2Y8_LUT4AB/S1END[2] Tile_X2Y8_LUT4AB/S1END[3]
+ Tile_X2Y7_LUT4AB/S1END[0] Tile_X2Y7_LUT4AB/S1END[1] Tile_X2Y7_LUT4AB/S1END[2] Tile_X2Y7_LUT4AB/S1END[3]
+ Tile_X2Y8_LUT4AB/S2MID[0] Tile_X2Y8_LUT4AB/S2MID[1] Tile_X2Y8_LUT4AB/S2MID[2] Tile_X2Y8_LUT4AB/S2MID[3]
+ Tile_X2Y8_LUT4AB/S2MID[4] Tile_X2Y8_LUT4AB/S2MID[5] Tile_X2Y8_LUT4AB/S2MID[6] Tile_X2Y8_LUT4AB/S2MID[7]
+ Tile_X2Y8_LUT4AB/S2END[0] Tile_X2Y8_LUT4AB/S2END[1] Tile_X2Y8_LUT4AB/S2END[2] Tile_X2Y8_LUT4AB/S2END[3]
+ Tile_X2Y8_LUT4AB/S2END[4] Tile_X2Y8_LUT4AB/S2END[5] Tile_X2Y8_LUT4AB/S2END[6] Tile_X2Y8_LUT4AB/S2END[7]
+ Tile_X2Y7_LUT4AB/S2END[0] Tile_X2Y7_LUT4AB/S2END[1] Tile_X2Y7_LUT4AB/S2END[2] Tile_X2Y7_LUT4AB/S2END[3]
+ Tile_X2Y7_LUT4AB/S2END[4] Tile_X2Y7_LUT4AB/S2END[5] Tile_X2Y7_LUT4AB/S2END[6] Tile_X2Y7_LUT4AB/S2END[7]
+ Tile_X2Y7_LUT4AB/S2MID[0] Tile_X2Y7_LUT4AB/S2MID[1] Tile_X2Y7_LUT4AB/S2MID[2] Tile_X2Y7_LUT4AB/S2MID[3]
+ Tile_X2Y7_LUT4AB/S2MID[4] Tile_X2Y7_LUT4AB/S2MID[5] Tile_X2Y7_LUT4AB/S2MID[6] Tile_X2Y7_LUT4AB/S2MID[7]
+ Tile_X2Y8_LUT4AB/S4END[0] Tile_X2Y8_LUT4AB/S4END[10] Tile_X2Y8_LUT4AB/S4END[11]
+ Tile_X2Y8_LUT4AB/S4END[12] Tile_X2Y8_LUT4AB/S4END[13] Tile_X2Y8_LUT4AB/S4END[14]
+ Tile_X2Y8_LUT4AB/S4END[15] Tile_X2Y8_LUT4AB/S4END[1] Tile_X2Y8_LUT4AB/S4END[2] Tile_X2Y8_LUT4AB/S4END[3]
+ Tile_X2Y8_LUT4AB/S4END[4] Tile_X2Y8_LUT4AB/S4END[5] Tile_X2Y8_LUT4AB/S4END[6] Tile_X2Y8_LUT4AB/S4END[7]
+ Tile_X2Y8_LUT4AB/S4END[8] Tile_X2Y8_LUT4AB/S4END[9] Tile_X2Y7_LUT4AB/S4END[0] Tile_X2Y7_LUT4AB/S4END[10]
+ Tile_X2Y7_LUT4AB/S4END[11] Tile_X2Y7_LUT4AB/S4END[12] Tile_X2Y7_LUT4AB/S4END[13]
+ Tile_X2Y7_LUT4AB/S4END[14] Tile_X2Y7_LUT4AB/S4END[15] Tile_X2Y7_LUT4AB/S4END[1]
+ Tile_X2Y7_LUT4AB/S4END[2] Tile_X2Y7_LUT4AB/S4END[3] Tile_X2Y7_LUT4AB/S4END[4] Tile_X2Y7_LUT4AB/S4END[5]
+ Tile_X2Y7_LUT4AB/S4END[6] Tile_X2Y7_LUT4AB/S4END[7] Tile_X2Y7_LUT4AB/S4END[8] Tile_X2Y7_LUT4AB/S4END[9]
+ Tile_X2Y8_LUT4AB/SS4END[0] Tile_X2Y8_LUT4AB/SS4END[10] Tile_X2Y8_LUT4AB/SS4END[11]
+ Tile_X2Y8_LUT4AB/SS4END[12] Tile_X2Y8_LUT4AB/SS4END[13] Tile_X2Y8_LUT4AB/SS4END[14]
+ Tile_X2Y8_LUT4AB/SS4END[15] Tile_X2Y8_LUT4AB/SS4END[1] Tile_X2Y8_LUT4AB/SS4END[2]
+ Tile_X2Y8_LUT4AB/SS4END[3] Tile_X2Y8_LUT4AB/SS4END[4] Tile_X2Y8_LUT4AB/SS4END[5]
+ Tile_X2Y8_LUT4AB/SS4END[6] Tile_X2Y8_LUT4AB/SS4END[7] Tile_X2Y8_LUT4AB/SS4END[8]
+ Tile_X2Y8_LUT4AB/SS4END[9] Tile_X2Y7_LUT4AB/SS4END[0] Tile_X2Y7_LUT4AB/SS4END[10]
+ Tile_X2Y7_LUT4AB/SS4END[11] Tile_X2Y7_LUT4AB/SS4END[12] Tile_X2Y7_LUT4AB/SS4END[13]
+ Tile_X2Y7_LUT4AB/SS4END[14] Tile_X2Y7_LUT4AB/SS4END[15] Tile_X2Y7_LUT4AB/SS4END[1]
+ Tile_X2Y7_LUT4AB/SS4END[2] Tile_X2Y7_LUT4AB/SS4END[3] Tile_X2Y7_LUT4AB/SS4END[4]
+ Tile_X2Y7_LUT4AB/SS4END[5] Tile_X2Y7_LUT4AB/SS4END[6] Tile_X2Y7_LUT4AB/SS4END[7]
+ Tile_X2Y7_LUT4AB/SS4END[8] Tile_X2Y7_LUT4AB/SS4END[9] Tile_X2Y7_LUT4AB/UserCLK Tile_X2Y6_LUT4AB/UserCLK
+ VGND VPWR Tile_X2Y7_LUT4AB/W1BEG[0] Tile_X2Y7_LUT4AB/W1BEG[1] Tile_X2Y7_LUT4AB/W1BEG[2]
+ Tile_X2Y7_LUT4AB/W1BEG[3] Tile_X3Y7_LUT4AB/W1BEG[0] Tile_X3Y7_LUT4AB/W1BEG[1] Tile_X3Y7_LUT4AB/W1BEG[2]
+ Tile_X3Y7_LUT4AB/W1BEG[3] Tile_X2Y7_LUT4AB/W2BEG[0] Tile_X2Y7_LUT4AB/W2BEG[1] Tile_X2Y7_LUT4AB/W2BEG[2]
+ Tile_X2Y7_LUT4AB/W2BEG[3] Tile_X2Y7_LUT4AB/W2BEG[4] Tile_X2Y7_LUT4AB/W2BEG[5] Tile_X2Y7_LUT4AB/W2BEG[6]
+ Tile_X2Y7_LUT4AB/W2BEG[7] Tile_X1Y7_LUT4AB/W2END[0] Tile_X1Y7_LUT4AB/W2END[1] Tile_X1Y7_LUT4AB/W2END[2]
+ Tile_X1Y7_LUT4AB/W2END[3] Tile_X1Y7_LUT4AB/W2END[4] Tile_X1Y7_LUT4AB/W2END[5] Tile_X1Y7_LUT4AB/W2END[6]
+ Tile_X1Y7_LUT4AB/W2END[7] Tile_X2Y7_LUT4AB/W2END[0] Tile_X2Y7_LUT4AB/W2END[1] Tile_X2Y7_LUT4AB/W2END[2]
+ Tile_X2Y7_LUT4AB/W2END[3] Tile_X2Y7_LUT4AB/W2END[4] Tile_X2Y7_LUT4AB/W2END[5] Tile_X2Y7_LUT4AB/W2END[6]
+ Tile_X2Y7_LUT4AB/W2END[7] Tile_X3Y7_LUT4AB/W2BEG[0] Tile_X3Y7_LUT4AB/W2BEG[1] Tile_X3Y7_LUT4AB/W2BEG[2]
+ Tile_X3Y7_LUT4AB/W2BEG[3] Tile_X3Y7_LUT4AB/W2BEG[4] Tile_X3Y7_LUT4AB/W2BEG[5] Tile_X3Y7_LUT4AB/W2BEG[6]
+ Tile_X3Y7_LUT4AB/W2BEG[7] Tile_X2Y7_LUT4AB/W6BEG[0] Tile_X2Y7_LUT4AB/W6BEG[10] Tile_X2Y7_LUT4AB/W6BEG[11]
+ Tile_X2Y7_LUT4AB/W6BEG[1] Tile_X2Y7_LUT4AB/W6BEG[2] Tile_X2Y7_LUT4AB/W6BEG[3] Tile_X2Y7_LUT4AB/W6BEG[4]
+ Tile_X2Y7_LUT4AB/W6BEG[5] Tile_X2Y7_LUT4AB/W6BEG[6] Tile_X2Y7_LUT4AB/W6BEG[7] Tile_X2Y7_LUT4AB/W6BEG[8]
+ Tile_X2Y7_LUT4AB/W6BEG[9] Tile_X3Y7_LUT4AB/W6BEG[0] Tile_X3Y7_LUT4AB/W6BEG[10] Tile_X3Y7_LUT4AB/W6BEG[11]
+ Tile_X3Y7_LUT4AB/W6BEG[1] Tile_X3Y7_LUT4AB/W6BEG[2] Tile_X3Y7_LUT4AB/W6BEG[3] Tile_X3Y7_LUT4AB/W6BEG[4]
+ Tile_X3Y7_LUT4AB/W6BEG[5] Tile_X3Y7_LUT4AB/W6BEG[6] Tile_X3Y7_LUT4AB/W6BEG[7] Tile_X3Y7_LUT4AB/W6BEG[8]
+ Tile_X3Y7_LUT4AB/W6BEG[9] Tile_X2Y7_LUT4AB/WW4BEG[0] Tile_X2Y7_LUT4AB/WW4BEG[10]
+ Tile_X2Y7_LUT4AB/WW4BEG[11] Tile_X2Y7_LUT4AB/WW4BEG[12] Tile_X2Y7_LUT4AB/WW4BEG[13]
+ Tile_X2Y7_LUT4AB/WW4BEG[14] Tile_X2Y7_LUT4AB/WW4BEG[15] Tile_X2Y7_LUT4AB/WW4BEG[1]
+ Tile_X2Y7_LUT4AB/WW4BEG[2] Tile_X2Y7_LUT4AB/WW4BEG[3] Tile_X2Y7_LUT4AB/WW4BEG[4]
+ Tile_X2Y7_LUT4AB/WW4BEG[5] Tile_X2Y7_LUT4AB/WW4BEG[6] Tile_X2Y7_LUT4AB/WW4BEG[7]
+ Tile_X2Y7_LUT4AB/WW4BEG[8] Tile_X2Y7_LUT4AB/WW4BEG[9] Tile_X3Y7_LUT4AB/WW4BEG[0]
+ Tile_X3Y7_LUT4AB/WW4BEG[10] Tile_X3Y7_LUT4AB/WW4BEG[11] Tile_X3Y7_LUT4AB/WW4BEG[12]
+ Tile_X3Y7_LUT4AB/WW4BEG[13] Tile_X3Y7_LUT4AB/WW4BEG[14] Tile_X3Y7_LUT4AB/WW4BEG[15]
+ Tile_X3Y7_LUT4AB/WW4BEG[1] Tile_X3Y7_LUT4AB/WW4BEG[2] Tile_X3Y7_LUT4AB/WW4BEG[3]
+ Tile_X3Y7_LUT4AB/WW4BEG[4] Tile_X3Y7_LUT4AB/WW4BEG[5] Tile_X3Y7_LUT4AB/WW4BEG[6]
+ Tile_X3Y7_LUT4AB/WW4BEG[7] Tile_X3Y7_LUT4AB/WW4BEG[8] Tile_X3Y7_LUT4AB/WW4BEG[9]
+ LUT4AB
XTile_X0Y2_W_TT_IF Tile_X0Y2_CLK_TT_PROJECT Tile_X1Y2_LUT4AB/E1END[0] Tile_X1Y2_LUT4AB/E1END[1]
+ Tile_X1Y2_LUT4AB/E1END[2] Tile_X1Y2_LUT4AB/E1END[3] Tile_X1Y2_LUT4AB/E2MID[0] Tile_X1Y2_LUT4AB/E2MID[1]
+ Tile_X1Y2_LUT4AB/E2MID[2] Tile_X1Y2_LUT4AB/E2MID[3] Tile_X1Y2_LUT4AB/E2MID[4] Tile_X1Y2_LUT4AB/E2MID[5]
+ Tile_X1Y2_LUT4AB/E2MID[6] Tile_X1Y2_LUT4AB/E2MID[7] Tile_X1Y2_LUT4AB/E2END[0] Tile_X1Y2_LUT4AB/E2END[1]
+ Tile_X1Y2_LUT4AB/E2END[2] Tile_X1Y2_LUT4AB/E2END[3] Tile_X1Y2_LUT4AB/E2END[4] Tile_X1Y2_LUT4AB/E2END[5]
+ Tile_X1Y2_LUT4AB/E2END[6] Tile_X1Y2_LUT4AB/E2END[7] Tile_X1Y2_LUT4AB/E6END[0] Tile_X1Y2_LUT4AB/E6END[10]
+ Tile_X1Y2_LUT4AB/E6END[11] Tile_X1Y2_LUT4AB/E6END[1] Tile_X1Y2_LUT4AB/E6END[2] Tile_X1Y2_LUT4AB/E6END[3]
+ Tile_X1Y2_LUT4AB/E6END[4] Tile_X1Y2_LUT4AB/E6END[5] Tile_X1Y2_LUT4AB/E6END[6] Tile_X1Y2_LUT4AB/E6END[7]
+ Tile_X1Y2_LUT4AB/E6END[8] Tile_X1Y2_LUT4AB/E6END[9] Tile_X1Y2_LUT4AB/EE4END[0] Tile_X1Y2_LUT4AB/EE4END[10]
+ Tile_X1Y2_LUT4AB/EE4END[11] Tile_X1Y2_LUT4AB/EE4END[12] Tile_X1Y2_LUT4AB/EE4END[13]
+ Tile_X1Y2_LUT4AB/EE4END[14] Tile_X1Y2_LUT4AB/EE4END[15] Tile_X1Y2_LUT4AB/EE4END[1]
+ Tile_X1Y2_LUT4AB/EE4END[2] Tile_X1Y2_LUT4AB/EE4END[3] Tile_X1Y2_LUT4AB/EE4END[4]
+ Tile_X1Y2_LUT4AB/EE4END[5] Tile_X1Y2_LUT4AB/EE4END[6] Tile_X1Y2_LUT4AB/EE4END[7]
+ Tile_X1Y2_LUT4AB/EE4END[8] Tile_X1Y2_LUT4AB/EE4END[9] Tile_X0Y2_ENA_TT_PROJECT FrameData[64]
+ FrameData[74] FrameData[75] FrameData[76] FrameData[77] FrameData[78] FrameData[79]
+ FrameData[80] FrameData[81] FrameData[82] FrameData[83] FrameData[65] FrameData[84]
+ FrameData[85] FrameData[86] FrameData[87] FrameData[88] FrameData[89] FrameData[90]
+ FrameData[91] FrameData[92] FrameData[93] FrameData[66] FrameData[94] FrameData[95]
+ FrameData[67] FrameData[68] FrameData[69] FrameData[70] FrameData[71] FrameData[72]
+ FrameData[73] Tile_X1Y2_LUT4AB/FrameData[0] Tile_X1Y2_LUT4AB/FrameData[10] Tile_X1Y2_LUT4AB/FrameData[11]
+ Tile_X1Y2_LUT4AB/FrameData[12] Tile_X1Y2_LUT4AB/FrameData[13] Tile_X1Y2_LUT4AB/FrameData[14]
+ Tile_X1Y2_LUT4AB/FrameData[15] Tile_X1Y2_LUT4AB/FrameData[16] Tile_X1Y2_LUT4AB/FrameData[17]
+ Tile_X1Y2_LUT4AB/FrameData[18] Tile_X1Y2_LUT4AB/FrameData[19] Tile_X1Y2_LUT4AB/FrameData[1]
+ Tile_X1Y2_LUT4AB/FrameData[20] Tile_X1Y2_LUT4AB/FrameData[21] Tile_X1Y2_LUT4AB/FrameData[22]
+ Tile_X1Y2_LUT4AB/FrameData[23] Tile_X1Y2_LUT4AB/FrameData[24] Tile_X1Y2_LUT4AB/FrameData[25]
+ Tile_X1Y2_LUT4AB/FrameData[26] Tile_X1Y2_LUT4AB/FrameData[27] Tile_X1Y2_LUT4AB/FrameData[28]
+ Tile_X1Y2_LUT4AB/FrameData[29] Tile_X1Y2_LUT4AB/FrameData[2] Tile_X1Y2_LUT4AB/FrameData[30]
+ Tile_X1Y2_LUT4AB/FrameData[31] Tile_X1Y2_LUT4AB/FrameData[3] Tile_X1Y2_LUT4AB/FrameData[4]
+ Tile_X1Y2_LUT4AB/FrameData[5] Tile_X1Y2_LUT4AB/FrameData[6] Tile_X1Y2_LUT4AB/FrameData[7]
+ Tile_X1Y2_LUT4AB/FrameData[8] Tile_X1Y2_LUT4AB/FrameData[9] Tile_X0Y2_W_TT_IF/FrameStrobe[0]
+ Tile_X0Y2_W_TT_IF/FrameStrobe[10] Tile_X0Y2_W_TT_IF/FrameStrobe[11] Tile_X0Y2_W_TT_IF/FrameStrobe[12]
+ Tile_X0Y2_W_TT_IF/FrameStrobe[13] Tile_X0Y2_W_TT_IF/FrameStrobe[14] Tile_X0Y2_W_TT_IF/FrameStrobe[15]
+ Tile_X0Y2_W_TT_IF/FrameStrobe[16] Tile_X0Y2_W_TT_IF/FrameStrobe[17] Tile_X0Y2_W_TT_IF/FrameStrobe[18]
+ Tile_X0Y2_W_TT_IF/FrameStrobe[19] Tile_X0Y2_W_TT_IF/FrameStrobe[1] Tile_X0Y2_W_TT_IF/FrameStrobe[2]
+ Tile_X0Y2_W_TT_IF/FrameStrobe[3] Tile_X0Y2_W_TT_IF/FrameStrobe[4] Tile_X0Y2_W_TT_IF/FrameStrobe[5]
+ Tile_X0Y2_W_TT_IF/FrameStrobe[6] Tile_X0Y2_W_TT_IF/FrameStrobe[7] Tile_X0Y2_W_TT_IF/FrameStrobe[8]
+ Tile_X0Y2_W_TT_IF/FrameStrobe[9] Tile_X0Y1_W_TT_IF/FrameStrobe[0] Tile_X0Y1_W_TT_IF/FrameStrobe[10]
+ Tile_X0Y1_W_TT_IF/FrameStrobe[11] Tile_X0Y1_W_TT_IF/FrameStrobe[12] Tile_X0Y1_W_TT_IF/FrameStrobe[13]
+ Tile_X0Y1_W_TT_IF/FrameStrobe[14] Tile_X0Y1_W_TT_IF/FrameStrobe[15] Tile_X0Y1_W_TT_IF/FrameStrobe[16]
+ Tile_X0Y1_W_TT_IF/FrameStrobe[17] Tile_X0Y1_W_TT_IF/FrameStrobe[18] Tile_X0Y1_W_TT_IF/FrameStrobe[19]
+ Tile_X0Y1_W_TT_IF/FrameStrobe[1] Tile_X0Y1_W_TT_IF/FrameStrobe[2] Tile_X0Y1_W_TT_IF/FrameStrobe[3]
+ Tile_X0Y1_W_TT_IF/FrameStrobe[4] Tile_X0Y1_W_TT_IF/FrameStrobe[5] Tile_X0Y1_W_TT_IF/FrameStrobe[6]
+ Tile_X0Y1_W_TT_IF/FrameStrobe[7] Tile_X0Y1_W_TT_IF/FrameStrobe[8] Tile_X0Y1_W_TT_IF/FrameStrobe[9]
+ Tile_X0Y2_W_TT_IF/N1BEG[0] Tile_X0Y2_W_TT_IF/N1BEG[1] Tile_X0Y2_W_TT_IF/N1BEG[2]
+ Tile_X0Y2_W_TT_IF/N1BEG[3] Tile_X0Y3_W_TT_IF/N1BEG[0] Tile_X0Y3_W_TT_IF/N1BEG[1]
+ Tile_X0Y3_W_TT_IF/N1BEG[2] Tile_X0Y3_W_TT_IF/N1BEG[3] Tile_X0Y2_W_TT_IF/N2BEG[0]
+ Tile_X0Y2_W_TT_IF/N2BEG[1] Tile_X0Y2_W_TT_IF/N2BEG[2] Tile_X0Y2_W_TT_IF/N2BEG[3]
+ Tile_X0Y2_W_TT_IF/N2BEG[4] Tile_X0Y2_W_TT_IF/N2BEG[5] Tile_X0Y2_W_TT_IF/N2BEG[6]
+ Tile_X0Y2_W_TT_IF/N2BEG[7] Tile_X0Y1_W_TT_IF/N2END[0] Tile_X0Y1_W_TT_IF/N2END[1]
+ Tile_X0Y1_W_TT_IF/N2END[2] Tile_X0Y1_W_TT_IF/N2END[3] Tile_X0Y1_W_TT_IF/N2END[4]
+ Tile_X0Y1_W_TT_IF/N2END[5] Tile_X0Y1_W_TT_IF/N2END[6] Tile_X0Y1_W_TT_IF/N2END[7]
+ Tile_X0Y2_W_TT_IF/N2END[0] Tile_X0Y2_W_TT_IF/N2END[1] Tile_X0Y2_W_TT_IF/N2END[2]
+ Tile_X0Y2_W_TT_IF/N2END[3] Tile_X0Y2_W_TT_IF/N2END[4] Tile_X0Y2_W_TT_IF/N2END[5]
+ Tile_X0Y2_W_TT_IF/N2END[6] Tile_X0Y2_W_TT_IF/N2END[7] Tile_X0Y3_W_TT_IF/N2BEG[0]
+ Tile_X0Y3_W_TT_IF/N2BEG[1] Tile_X0Y3_W_TT_IF/N2BEG[2] Tile_X0Y3_W_TT_IF/N2BEG[3]
+ Tile_X0Y3_W_TT_IF/N2BEG[4] Tile_X0Y3_W_TT_IF/N2BEG[5] Tile_X0Y3_W_TT_IF/N2BEG[6]
+ Tile_X0Y3_W_TT_IF/N2BEG[7] Tile_X0Y2_W_TT_IF/N4BEG[0] Tile_X0Y2_W_TT_IF/N4BEG[10]
+ Tile_X0Y2_W_TT_IF/N4BEG[11] Tile_X0Y2_W_TT_IF/N4BEG[12] Tile_X0Y2_W_TT_IF/N4BEG[13]
+ Tile_X0Y2_W_TT_IF/N4BEG[14] Tile_X0Y2_W_TT_IF/N4BEG[15] Tile_X0Y2_W_TT_IF/N4BEG[1]
+ Tile_X0Y2_W_TT_IF/N4BEG[2] Tile_X0Y2_W_TT_IF/N4BEG[3] Tile_X0Y2_W_TT_IF/N4BEG[4]
+ Tile_X0Y2_W_TT_IF/N4BEG[5] Tile_X0Y2_W_TT_IF/N4BEG[6] Tile_X0Y2_W_TT_IF/N4BEG[7]
+ Tile_X0Y2_W_TT_IF/N4BEG[8] Tile_X0Y2_W_TT_IF/N4BEG[9] Tile_X0Y3_W_TT_IF/N4BEG[0]
+ Tile_X0Y3_W_TT_IF/N4BEG[10] Tile_X0Y3_W_TT_IF/N4BEG[11] Tile_X0Y3_W_TT_IF/N4BEG[12]
+ Tile_X0Y3_W_TT_IF/N4BEG[13] Tile_X0Y3_W_TT_IF/N4BEG[14] Tile_X0Y3_W_TT_IF/N4BEG[15]
+ Tile_X0Y3_W_TT_IF/N4BEG[1] Tile_X0Y3_W_TT_IF/N4BEG[2] Tile_X0Y3_W_TT_IF/N4BEG[3]
+ Tile_X0Y3_W_TT_IF/N4BEG[4] Tile_X0Y3_W_TT_IF/N4BEG[5] Tile_X0Y3_W_TT_IF/N4BEG[6]
+ Tile_X0Y3_W_TT_IF/N4BEG[7] Tile_X0Y3_W_TT_IF/N4BEG[8] Tile_X0Y3_W_TT_IF/N4BEG[9]
+ Tile_X0Y2_RST_N_TT_PROJECT Tile_X0Y3_W_TT_IF/S1END[0] Tile_X0Y3_W_TT_IF/S1END[1]
+ Tile_X0Y3_W_TT_IF/S1END[2] Tile_X0Y3_W_TT_IF/S1END[3] Tile_X0Y2_W_TT_IF/S1END[0]
+ Tile_X0Y2_W_TT_IF/S1END[1] Tile_X0Y2_W_TT_IF/S1END[2] Tile_X0Y2_W_TT_IF/S1END[3]
+ Tile_X0Y3_W_TT_IF/S2MID[0] Tile_X0Y3_W_TT_IF/S2MID[1] Tile_X0Y3_W_TT_IF/S2MID[2]
+ Tile_X0Y3_W_TT_IF/S2MID[3] Tile_X0Y3_W_TT_IF/S2MID[4] Tile_X0Y3_W_TT_IF/S2MID[5]
+ Tile_X0Y3_W_TT_IF/S2MID[6] Tile_X0Y3_W_TT_IF/S2MID[7] Tile_X0Y3_W_TT_IF/S2END[0]
+ Tile_X0Y3_W_TT_IF/S2END[1] Tile_X0Y3_W_TT_IF/S2END[2] Tile_X0Y3_W_TT_IF/S2END[3]
+ Tile_X0Y3_W_TT_IF/S2END[4] Tile_X0Y3_W_TT_IF/S2END[5] Tile_X0Y3_W_TT_IF/S2END[6]
+ Tile_X0Y3_W_TT_IF/S2END[7] Tile_X0Y2_W_TT_IF/S2END[0] Tile_X0Y2_W_TT_IF/S2END[1]
+ Tile_X0Y2_W_TT_IF/S2END[2] Tile_X0Y2_W_TT_IF/S2END[3] Tile_X0Y2_W_TT_IF/S2END[4]
+ Tile_X0Y2_W_TT_IF/S2END[5] Tile_X0Y2_W_TT_IF/S2END[6] Tile_X0Y2_W_TT_IF/S2END[7]
+ Tile_X0Y2_W_TT_IF/S2MID[0] Tile_X0Y2_W_TT_IF/S2MID[1] Tile_X0Y2_W_TT_IF/S2MID[2]
+ Tile_X0Y2_W_TT_IF/S2MID[3] Tile_X0Y2_W_TT_IF/S2MID[4] Tile_X0Y2_W_TT_IF/S2MID[5]
+ Tile_X0Y2_W_TT_IF/S2MID[6] Tile_X0Y2_W_TT_IF/S2MID[7] Tile_X0Y3_W_TT_IF/S4END[0]
+ Tile_X0Y3_W_TT_IF/S4END[10] Tile_X0Y3_W_TT_IF/S4END[11] Tile_X0Y3_W_TT_IF/S4END[12]
+ Tile_X0Y3_W_TT_IF/S4END[13] Tile_X0Y3_W_TT_IF/S4END[14] Tile_X0Y3_W_TT_IF/S4END[15]
+ Tile_X0Y3_W_TT_IF/S4END[1] Tile_X0Y3_W_TT_IF/S4END[2] Tile_X0Y3_W_TT_IF/S4END[3]
+ Tile_X0Y3_W_TT_IF/S4END[4] Tile_X0Y3_W_TT_IF/S4END[5] Tile_X0Y3_W_TT_IF/S4END[6]
+ Tile_X0Y3_W_TT_IF/S4END[7] Tile_X0Y3_W_TT_IF/S4END[8] Tile_X0Y3_W_TT_IF/S4END[9]
+ Tile_X0Y2_W_TT_IF/S4END[0] Tile_X0Y2_W_TT_IF/S4END[10] Tile_X0Y2_W_TT_IF/S4END[11]
+ Tile_X0Y2_W_TT_IF/S4END[12] Tile_X0Y2_W_TT_IF/S4END[13] Tile_X0Y2_W_TT_IF/S4END[14]
+ Tile_X0Y2_W_TT_IF/S4END[15] Tile_X0Y2_W_TT_IF/S4END[1] Tile_X0Y2_W_TT_IF/S4END[2]
+ Tile_X0Y2_W_TT_IF/S4END[3] Tile_X0Y2_W_TT_IF/S4END[4] Tile_X0Y2_W_TT_IF/S4END[5]
+ Tile_X0Y2_W_TT_IF/S4END[6] Tile_X0Y2_W_TT_IF/S4END[7] Tile_X0Y2_W_TT_IF/S4END[8]
+ Tile_X0Y2_W_TT_IF/S4END[9] Tile_X0Y2_UIO_IN_TT_PROJECT0 Tile_X0Y2_UIO_IN_TT_PROJECT1
+ Tile_X0Y2_UIO_IN_TT_PROJECT2 Tile_X0Y2_UIO_IN_TT_PROJECT3 Tile_X0Y2_UIO_IN_TT_PROJECT4
+ Tile_X0Y2_UIO_IN_TT_PROJECT5 Tile_X0Y2_UIO_IN_TT_PROJECT6 Tile_X0Y2_UIO_IN_TT_PROJECT7
+ Tile_X0Y2_UIO_OE_TT_PROJECT0 Tile_X0Y2_UIO_OE_TT_PROJECT1 Tile_X0Y2_UIO_OE_TT_PROJECT2
+ Tile_X0Y2_UIO_OE_TT_PROJECT3 Tile_X0Y2_UIO_OE_TT_PROJECT4 Tile_X0Y2_UIO_OE_TT_PROJECT5
+ Tile_X0Y2_UIO_OE_TT_PROJECT6 Tile_X0Y2_UIO_OE_TT_PROJECT7 Tile_X0Y2_UIO_OUT_TT_PROJECT0
+ Tile_X0Y2_UIO_OUT_TT_PROJECT1 Tile_X0Y2_UIO_OUT_TT_PROJECT2 Tile_X0Y2_UIO_OUT_TT_PROJECT3
+ Tile_X0Y2_UIO_OUT_TT_PROJECT4 Tile_X0Y2_UIO_OUT_TT_PROJECT5 Tile_X0Y2_UIO_OUT_TT_PROJECT6
+ Tile_X0Y2_UIO_OUT_TT_PROJECT7 Tile_X0Y2_UI_IN_TT_PROJECT0 Tile_X0Y2_UI_IN_TT_PROJECT1
+ Tile_X0Y2_UI_IN_TT_PROJECT2 Tile_X0Y2_UI_IN_TT_PROJECT3 Tile_X0Y2_UI_IN_TT_PROJECT4
+ Tile_X0Y2_UI_IN_TT_PROJECT5 Tile_X0Y2_UI_IN_TT_PROJECT6 Tile_X0Y2_UI_IN_TT_PROJECT7
+ Tile_X0Y2_UO_OUT_TT_PROJECT0 Tile_X0Y2_UO_OUT_TT_PROJECT1 Tile_X0Y2_UO_OUT_TT_PROJECT2
+ Tile_X0Y2_UO_OUT_TT_PROJECT3 Tile_X0Y2_UO_OUT_TT_PROJECT4 Tile_X0Y2_UO_OUT_TT_PROJECT5
+ Tile_X0Y2_UO_OUT_TT_PROJECT6 Tile_X0Y2_UO_OUT_TT_PROJECT7 Tile_X0Y2_W_TT_IF/UserCLK
+ Tile_X0Y1_W_TT_IF/UserCLK VGND VPWR Tile_X1Y2_LUT4AB/W1BEG[0] Tile_X1Y2_LUT4AB/W1BEG[1]
+ Tile_X1Y2_LUT4AB/W1BEG[2] Tile_X1Y2_LUT4AB/W1BEG[3] Tile_X1Y2_LUT4AB/W2BEGb[0] Tile_X1Y2_LUT4AB/W2BEGb[1]
+ Tile_X1Y2_LUT4AB/W2BEGb[2] Tile_X1Y2_LUT4AB/W2BEGb[3] Tile_X1Y2_LUT4AB/W2BEGb[4]
+ Tile_X1Y2_LUT4AB/W2BEGb[5] Tile_X1Y2_LUT4AB/W2BEGb[6] Tile_X1Y2_LUT4AB/W2BEGb[7]
+ Tile_X1Y2_LUT4AB/W2BEG[0] Tile_X1Y2_LUT4AB/W2BEG[1] Tile_X1Y2_LUT4AB/W2BEG[2] Tile_X1Y2_LUT4AB/W2BEG[3]
+ Tile_X1Y2_LUT4AB/W2BEG[4] Tile_X1Y2_LUT4AB/W2BEG[5] Tile_X1Y2_LUT4AB/W2BEG[6] Tile_X1Y2_LUT4AB/W2BEG[7]
+ Tile_X1Y2_LUT4AB/W6BEG[0] Tile_X1Y2_LUT4AB/W6BEG[10] Tile_X1Y2_LUT4AB/W6BEG[11]
+ Tile_X1Y2_LUT4AB/W6BEG[1] Tile_X1Y2_LUT4AB/W6BEG[2] Tile_X1Y2_LUT4AB/W6BEG[3] Tile_X1Y2_LUT4AB/W6BEG[4]
+ Tile_X1Y2_LUT4AB/W6BEG[5] Tile_X1Y2_LUT4AB/W6BEG[6] Tile_X1Y2_LUT4AB/W6BEG[7] Tile_X1Y2_LUT4AB/W6BEG[8]
+ Tile_X1Y2_LUT4AB/W6BEG[9] Tile_X1Y2_LUT4AB/WW4BEG[0] Tile_X1Y2_LUT4AB/WW4BEG[10]
+ Tile_X1Y2_LUT4AB/WW4BEG[11] Tile_X1Y2_LUT4AB/WW4BEG[12] Tile_X1Y2_LUT4AB/WW4BEG[13]
+ Tile_X1Y2_LUT4AB/WW4BEG[14] Tile_X1Y2_LUT4AB/WW4BEG[15] Tile_X1Y2_LUT4AB/WW4BEG[1]
+ Tile_X1Y2_LUT4AB/WW4BEG[2] Tile_X1Y2_LUT4AB/WW4BEG[3] Tile_X1Y2_LUT4AB/WW4BEG[4]
+ Tile_X1Y2_LUT4AB/WW4BEG[5] Tile_X1Y2_LUT4AB/WW4BEG[6] Tile_X1Y2_LUT4AB/WW4BEG[7]
+ Tile_X1Y2_LUT4AB/WW4BEG[8] Tile_X1Y2_LUT4AB/WW4BEG[9] W_TT_IF
XTile_X4Y5_LUT4AB Tile_X4Y6_LUT4AB/Co Tile_X4Y5_LUT4AB/Co Tile_X4Y5_LUT4AB/E1BEG[0]
+ Tile_X4Y5_LUT4AB/E1BEG[1] Tile_X4Y5_LUT4AB/E1BEG[2] Tile_X4Y5_LUT4AB/E1BEG[3] Tile_X4Y5_LUT4AB/E1END[0]
+ Tile_X4Y5_LUT4AB/E1END[1] Tile_X4Y5_LUT4AB/E1END[2] Tile_X4Y5_LUT4AB/E1END[3] Tile_X4Y5_LUT4AB/E2BEG[0]
+ Tile_X4Y5_LUT4AB/E2BEG[1] Tile_X4Y5_LUT4AB/E2BEG[2] Tile_X4Y5_LUT4AB/E2BEG[3] Tile_X4Y5_LUT4AB/E2BEG[4]
+ Tile_X4Y5_LUT4AB/E2BEG[5] Tile_X4Y5_LUT4AB/E2BEG[6] Tile_X4Y5_LUT4AB/E2BEG[7] Tile_X5Y5_E_TT_IF/E2END[0]
+ Tile_X5Y5_E_TT_IF/E2END[1] Tile_X5Y5_E_TT_IF/E2END[2] Tile_X5Y5_E_TT_IF/E2END[3]
+ Tile_X5Y5_E_TT_IF/E2END[4] Tile_X5Y5_E_TT_IF/E2END[5] Tile_X5Y5_E_TT_IF/E2END[6]
+ Tile_X5Y5_E_TT_IF/E2END[7] Tile_X4Y5_LUT4AB/E2END[0] Tile_X4Y5_LUT4AB/E2END[1] Tile_X4Y5_LUT4AB/E2END[2]
+ Tile_X4Y5_LUT4AB/E2END[3] Tile_X4Y5_LUT4AB/E2END[4] Tile_X4Y5_LUT4AB/E2END[5] Tile_X4Y5_LUT4AB/E2END[6]
+ Tile_X4Y5_LUT4AB/E2END[7] Tile_X4Y5_LUT4AB/E2MID[0] Tile_X4Y5_LUT4AB/E2MID[1] Tile_X4Y5_LUT4AB/E2MID[2]
+ Tile_X4Y5_LUT4AB/E2MID[3] Tile_X4Y5_LUT4AB/E2MID[4] Tile_X4Y5_LUT4AB/E2MID[5] Tile_X4Y5_LUT4AB/E2MID[6]
+ Tile_X4Y5_LUT4AB/E2MID[7] Tile_X4Y5_LUT4AB/E6BEG[0] Tile_X4Y5_LUT4AB/E6BEG[10] Tile_X4Y5_LUT4AB/E6BEG[11]
+ Tile_X4Y5_LUT4AB/E6BEG[1] Tile_X4Y5_LUT4AB/E6BEG[2] Tile_X4Y5_LUT4AB/E6BEG[3] Tile_X4Y5_LUT4AB/E6BEG[4]
+ Tile_X4Y5_LUT4AB/E6BEG[5] Tile_X4Y5_LUT4AB/E6BEG[6] Tile_X4Y5_LUT4AB/E6BEG[7] Tile_X4Y5_LUT4AB/E6BEG[8]
+ Tile_X4Y5_LUT4AB/E6BEG[9] Tile_X4Y5_LUT4AB/E6END[0] Tile_X4Y5_LUT4AB/E6END[10] Tile_X4Y5_LUT4AB/E6END[11]
+ Tile_X4Y5_LUT4AB/E6END[1] Tile_X4Y5_LUT4AB/E6END[2] Tile_X4Y5_LUT4AB/E6END[3] Tile_X4Y5_LUT4AB/E6END[4]
+ Tile_X4Y5_LUT4AB/E6END[5] Tile_X4Y5_LUT4AB/E6END[6] Tile_X4Y5_LUT4AB/E6END[7] Tile_X4Y5_LUT4AB/E6END[8]
+ Tile_X4Y5_LUT4AB/E6END[9] Tile_X4Y5_LUT4AB/EE4BEG[0] Tile_X4Y5_LUT4AB/EE4BEG[10]
+ Tile_X4Y5_LUT4AB/EE4BEG[11] Tile_X4Y5_LUT4AB/EE4BEG[12] Tile_X4Y5_LUT4AB/EE4BEG[13]
+ Tile_X4Y5_LUT4AB/EE4BEG[14] Tile_X4Y5_LUT4AB/EE4BEG[15] Tile_X4Y5_LUT4AB/EE4BEG[1]
+ Tile_X4Y5_LUT4AB/EE4BEG[2] Tile_X4Y5_LUT4AB/EE4BEG[3] Tile_X4Y5_LUT4AB/EE4BEG[4]
+ Tile_X4Y5_LUT4AB/EE4BEG[5] Tile_X4Y5_LUT4AB/EE4BEG[6] Tile_X4Y5_LUT4AB/EE4BEG[7]
+ Tile_X4Y5_LUT4AB/EE4BEG[8] Tile_X4Y5_LUT4AB/EE4BEG[9] Tile_X4Y5_LUT4AB/EE4END[0]
+ Tile_X4Y5_LUT4AB/EE4END[10] Tile_X4Y5_LUT4AB/EE4END[11] Tile_X4Y5_LUT4AB/EE4END[12]
+ Tile_X4Y5_LUT4AB/EE4END[13] Tile_X4Y5_LUT4AB/EE4END[14] Tile_X4Y5_LUT4AB/EE4END[15]
+ Tile_X4Y5_LUT4AB/EE4END[1] Tile_X4Y5_LUT4AB/EE4END[2] Tile_X4Y5_LUT4AB/EE4END[3]
+ Tile_X4Y5_LUT4AB/EE4END[4] Tile_X4Y5_LUT4AB/EE4END[5] Tile_X4Y5_LUT4AB/EE4END[6]
+ Tile_X4Y5_LUT4AB/EE4END[7] Tile_X4Y5_LUT4AB/EE4END[8] Tile_X4Y5_LUT4AB/EE4END[9]
+ Tile_X4Y5_LUT4AB/FrameData[0] Tile_X4Y5_LUT4AB/FrameData[10] Tile_X4Y5_LUT4AB/FrameData[11]
+ Tile_X4Y5_LUT4AB/FrameData[12] Tile_X4Y5_LUT4AB/FrameData[13] Tile_X4Y5_LUT4AB/FrameData[14]
+ Tile_X4Y5_LUT4AB/FrameData[15] Tile_X4Y5_LUT4AB/FrameData[16] Tile_X4Y5_LUT4AB/FrameData[17]
+ Tile_X4Y5_LUT4AB/FrameData[18] Tile_X4Y5_LUT4AB/FrameData[19] Tile_X4Y5_LUT4AB/FrameData[1]
+ Tile_X4Y5_LUT4AB/FrameData[20] Tile_X4Y5_LUT4AB/FrameData[21] Tile_X4Y5_LUT4AB/FrameData[22]
+ Tile_X4Y5_LUT4AB/FrameData[23] Tile_X4Y5_LUT4AB/FrameData[24] Tile_X4Y5_LUT4AB/FrameData[25]
+ Tile_X4Y5_LUT4AB/FrameData[26] Tile_X4Y5_LUT4AB/FrameData[27] Tile_X4Y5_LUT4AB/FrameData[28]
+ Tile_X4Y5_LUT4AB/FrameData[29] Tile_X4Y5_LUT4AB/FrameData[2] Tile_X4Y5_LUT4AB/FrameData[30]
+ Tile_X4Y5_LUT4AB/FrameData[31] Tile_X4Y5_LUT4AB/FrameData[3] Tile_X4Y5_LUT4AB/FrameData[4]
+ Tile_X4Y5_LUT4AB/FrameData[5] Tile_X4Y5_LUT4AB/FrameData[6] Tile_X4Y5_LUT4AB/FrameData[7]
+ Tile_X4Y5_LUT4AB/FrameData[8] Tile_X4Y5_LUT4AB/FrameData[9] Tile_X5Y5_E_TT_IF/FrameData[0]
+ Tile_X5Y5_E_TT_IF/FrameData[10] Tile_X5Y5_E_TT_IF/FrameData[11] Tile_X5Y5_E_TT_IF/FrameData[12]
+ Tile_X5Y5_E_TT_IF/FrameData[13] Tile_X5Y5_E_TT_IF/FrameData[14] Tile_X5Y5_E_TT_IF/FrameData[15]
+ Tile_X5Y5_E_TT_IF/FrameData[16] Tile_X5Y5_E_TT_IF/FrameData[17] Tile_X5Y5_E_TT_IF/FrameData[18]
+ Tile_X5Y5_E_TT_IF/FrameData[19] Tile_X5Y5_E_TT_IF/FrameData[1] Tile_X5Y5_E_TT_IF/FrameData[20]
+ Tile_X5Y5_E_TT_IF/FrameData[21] Tile_X5Y5_E_TT_IF/FrameData[22] Tile_X5Y5_E_TT_IF/FrameData[23]
+ Tile_X5Y5_E_TT_IF/FrameData[24] Tile_X5Y5_E_TT_IF/FrameData[25] Tile_X5Y5_E_TT_IF/FrameData[26]
+ Tile_X5Y5_E_TT_IF/FrameData[27] Tile_X5Y5_E_TT_IF/FrameData[28] Tile_X5Y5_E_TT_IF/FrameData[29]
+ Tile_X5Y5_E_TT_IF/FrameData[2] Tile_X5Y5_E_TT_IF/FrameData[30] Tile_X5Y5_E_TT_IF/FrameData[31]
+ Tile_X5Y5_E_TT_IF/FrameData[3] Tile_X5Y5_E_TT_IF/FrameData[4] Tile_X5Y5_E_TT_IF/FrameData[5]
+ Tile_X5Y5_E_TT_IF/FrameData[6] Tile_X5Y5_E_TT_IF/FrameData[7] Tile_X5Y5_E_TT_IF/FrameData[8]
+ Tile_X5Y5_E_TT_IF/FrameData[9] Tile_X4Y5_LUT4AB/FrameStrobe[0] Tile_X4Y5_LUT4AB/FrameStrobe[10]
+ Tile_X4Y5_LUT4AB/FrameStrobe[11] Tile_X4Y5_LUT4AB/FrameStrobe[12] Tile_X4Y5_LUT4AB/FrameStrobe[13]
+ Tile_X4Y5_LUT4AB/FrameStrobe[14] Tile_X4Y5_LUT4AB/FrameStrobe[15] Tile_X4Y5_LUT4AB/FrameStrobe[16]
+ Tile_X4Y5_LUT4AB/FrameStrobe[17] Tile_X4Y5_LUT4AB/FrameStrobe[18] Tile_X4Y5_LUT4AB/FrameStrobe[19]
+ Tile_X4Y5_LUT4AB/FrameStrobe[1] Tile_X4Y5_LUT4AB/FrameStrobe[2] Tile_X4Y5_LUT4AB/FrameStrobe[3]
+ Tile_X4Y5_LUT4AB/FrameStrobe[4] Tile_X4Y5_LUT4AB/FrameStrobe[5] Tile_X4Y5_LUT4AB/FrameStrobe[6]
+ Tile_X4Y5_LUT4AB/FrameStrobe[7] Tile_X4Y5_LUT4AB/FrameStrobe[8] Tile_X4Y5_LUT4AB/FrameStrobe[9]
+ Tile_X4Y4_LUT4AB/FrameStrobe[0] Tile_X4Y4_LUT4AB/FrameStrobe[10] Tile_X4Y4_LUT4AB/FrameStrobe[11]
+ Tile_X4Y4_LUT4AB/FrameStrobe[12] Tile_X4Y4_LUT4AB/FrameStrobe[13] Tile_X4Y4_LUT4AB/FrameStrobe[14]
+ Tile_X4Y4_LUT4AB/FrameStrobe[15] Tile_X4Y4_LUT4AB/FrameStrobe[16] Tile_X4Y4_LUT4AB/FrameStrobe[17]
+ Tile_X4Y4_LUT4AB/FrameStrobe[18] Tile_X4Y4_LUT4AB/FrameStrobe[19] Tile_X4Y4_LUT4AB/FrameStrobe[1]
+ Tile_X4Y4_LUT4AB/FrameStrobe[2] Tile_X4Y4_LUT4AB/FrameStrobe[3] Tile_X4Y4_LUT4AB/FrameStrobe[4]
+ Tile_X4Y4_LUT4AB/FrameStrobe[5] Tile_X4Y4_LUT4AB/FrameStrobe[6] Tile_X4Y4_LUT4AB/FrameStrobe[7]
+ Tile_X4Y4_LUT4AB/FrameStrobe[8] Tile_X4Y4_LUT4AB/FrameStrobe[9] Tile_X4Y5_LUT4AB/N1BEG[0]
+ Tile_X4Y5_LUT4AB/N1BEG[1] Tile_X4Y5_LUT4AB/N1BEG[2] Tile_X4Y5_LUT4AB/N1BEG[3] Tile_X4Y6_LUT4AB/N1BEG[0]
+ Tile_X4Y6_LUT4AB/N1BEG[1] Tile_X4Y6_LUT4AB/N1BEG[2] Tile_X4Y6_LUT4AB/N1BEG[3] Tile_X4Y5_LUT4AB/N2BEG[0]
+ Tile_X4Y5_LUT4AB/N2BEG[1] Tile_X4Y5_LUT4AB/N2BEG[2] Tile_X4Y5_LUT4AB/N2BEG[3] Tile_X4Y5_LUT4AB/N2BEG[4]
+ Tile_X4Y5_LUT4AB/N2BEG[5] Tile_X4Y5_LUT4AB/N2BEG[6] Tile_X4Y5_LUT4AB/N2BEG[7] Tile_X4Y4_LUT4AB/N2END[0]
+ Tile_X4Y4_LUT4AB/N2END[1] Tile_X4Y4_LUT4AB/N2END[2] Tile_X4Y4_LUT4AB/N2END[3] Tile_X4Y4_LUT4AB/N2END[4]
+ Tile_X4Y4_LUT4AB/N2END[5] Tile_X4Y4_LUT4AB/N2END[6] Tile_X4Y4_LUT4AB/N2END[7] Tile_X4Y5_LUT4AB/N2END[0]
+ Tile_X4Y5_LUT4AB/N2END[1] Tile_X4Y5_LUT4AB/N2END[2] Tile_X4Y5_LUT4AB/N2END[3] Tile_X4Y5_LUT4AB/N2END[4]
+ Tile_X4Y5_LUT4AB/N2END[5] Tile_X4Y5_LUT4AB/N2END[6] Tile_X4Y5_LUT4AB/N2END[7] Tile_X4Y6_LUT4AB/N2BEG[0]
+ Tile_X4Y6_LUT4AB/N2BEG[1] Tile_X4Y6_LUT4AB/N2BEG[2] Tile_X4Y6_LUT4AB/N2BEG[3] Tile_X4Y6_LUT4AB/N2BEG[4]
+ Tile_X4Y6_LUT4AB/N2BEG[5] Tile_X4Y6_LUT4AB/N2BEG[6] Tile_X4Y6_LUT4AB/N2BEG[7] Tile_X4Y5_LUT4AB/N4BEG[0]
+ Tile_X4Y5_LUT4AB/N4BEG[10] Tile_X4Y5_LUT4AB/N4BEG[11] Tile_X4Y5_LUT4AB/N4BEG[12]
+ Tile_X4Y5_LUT4AB/N4BEG[13] Tile_X4Y5_LUT4AB/N4BEG[14] Tile_X4Y5_LUT4AB/N4BEG[15]
+ Tile_X4Y5_LUT4AB/N4BEG[1] Tile_X4Y5_LUT4AB/N4BEG[2] Tile_X4Y5_LUT4AB/N4BEG[3] Tile_X4Y5_LUT4AB/N4BEG[4]
+ Tile_X4Y5_LUT4AB/N4BEG[5] Tile_X4Y5_LUT4AB/N4BEG[6] Tile_X4Y5_LUT4AB/N4BEG[7] Tile_X4Y5_LUT4AB/N4BEG[8]
+ Tile_X4Y5_LUT4AB/N4BEG[9] Tile_X4Y6_LUT4AB/N4BEG[0] Tile_X4Y6_LUT4AB/N4BEG[10] Tile_X4Y6_LUT4AB/N4BEG[11]
+ Tile_X4Y6_LUT4AB/N4BEG[12] Tile_X4Y6_LUT4AB/N4BEG[13] Tile_X4Y6_LUT4AB/N4BEG[14]
+ Tile_X4Y6_LUT4AB/N4BEG[15] Tile_X4Y6_LUT4AB/N4BEG[1] Tile_X4Y6_LUT4AB/N4BEG[2] Tile_X4Y6_LUT4AB/N4BEG[3]
+ Tile_X4Y6_LUT4AB/N4BEG[4] Tile_X4Y6_LUT4AB/N4BEG[5] Tile_X4Y6_LUT4AB/N4BEG[6] Tile_X4Y6_LUT4AB/N4BEG[7]
+ Tile_X4Y6_LUT4AB/N4BEG[8] Tile_X4Y6_LUT4AB/N4BEG[9] Tile_X4Y5_LUT4AB/NN4BEG[0] Tile_X4Y5_LUT4AB/NN4BEG[10]
+ Tile_X4Y5_LUT4AB/NN4BEG[11] Tile_X4Y5_LUT4AB/NN4BEG[12] Tile_X4Y5_LUT4AB/NN4BEG[13]
+ Tile_X4Y5_LUT4AB/NN4BEG[14] Tile_X4Y5_LUT4AB/NN4BEG[15] Tile_X4Y5_LUT4AB/NN4BEG[1]
+ Tile_X4Y5_LUT4AB/NN4BEG[2] Tile_X4Y5_LUT4AB/NN4BEG[3] Tile_X4Y5_LUT4AB/NN4BEG[4]
+ Tile_X4Y5_LUT4AB/NN4BEG[5] Tile_X4Y5_LUT4AB/NN4BEG[6] Tile_X4Y5_LUT4AB/NN4BEG[7]
+ Tile_X4Y5_LUT4AB/NN4BEG[8] Tile_X4Y5_LUT4AB/NN4BEG[9] Tile_X4Y6_LUT4AB/NN4BEG[0]
+ Tile_X4Y6_LUT4AB/NN4BEG[10] Tile_X4Y6_LUT4AB/NN4BEG[11] Tile_X4Y6_LUT4AB/NN4BEG[12]
+ Tile_X4Y6_LUT4AB/NN4BEG[13] Tile_X4Y6_LUT4AB/NN4BEG[14] Tile_X4Y6_LUT4AB/NN4BEG[15]
+ Tile_X4Y6_LUT4AB/NN4BEG[1] Tile_X4Y6_LUT4AB/NN4BEG[2] Tile_X4Y6_LUT4AB/NN4BEG[3]
+ Tile_X4Y6_LUT4AB/NN4BEG[4] Tile_X4Y6_LUT4AB/NN4BEG[5] Tile_X4Y6_LUT4AB/NN4BEG[6]
+ Tile_X4Y6_LUT4AB/NN4BEG[7] Tile_X4Y6_LUT4AB/NN4BEG[8] Tile_X4Y6_LUT4AB/NN4BEG[9]
+ Tile_X4Y6_LUT4AB/S1END[0] Tile_X4Y6_LUT4AB/S1END[1] Tile_X4Y6_LUT4AB/S1END[2] Tile_X4Y6_LUT4AB/S1END[3]
+ Tile_X4Y5_LUT4AB/S1END[0] Tile_X4Y5_LUT4AB/S1END[1] Tile_X4Y5_LUT4AB/S1END[2] Tile_X4Y5_LUT4AB/S1END[3]
+ Tile_X4Y6_LUT4AB/S2MID[0] Tile_X4Y6_LUT4AB/S2MID[1] Tile_X4Y6_LUT4AB/S2MID[2] Tile_X4Y6_LUT4AB/S2MID[3]
+ Tile_X4Y6_LUT4AB/S2MID[4] Tile_X4Y6_LUT4AB/S2MID[5] Tile_X4Y6_LUT4AB/S2MID[6] Tile_X4Y6_LUT4AB/S2MID[7]
+ Tile_X4Y6_LUT4AB/S2END[0] Tile_X4Y6_LUT4AB/S2END[1] Tile_X4Y6_LUT4AB/S2END[2] Tile_X4Y6_LUT4AB/S2END[3]
+ Tile_X4Y6_LUT4AB/S2END[4] Tile_X4Y6_LUT4AB/S2END[5] Tile_X4Y6_LUT4AB/S2END[6] Tile_X4Y6_LUT4AB/S2END[7]
+ Tile_X4Y5_LUT4AB/S2END[0] Tile_X4Y5_LUT4AB/S2END[1] Tile_X4Y5_LUT4AB/S2END[2] Tile_X4Y5_LUT4AB/S2END[3]
+ Tile_X4Y5_LUT4AB/S2END[4] Tile_X4Y5_LUT4AB/S2END[5] Tile_X4Y5_LUT4AB/S2END[6] Tile_X4Y5_LUT4AB/S2END[7]
+ Tile_X4Y5_LUT4AB/S2MID[0] Tile_X4Y5_LUT4AB/S2MID[1] Tile_X4Y5_LUT4AB/S2MID[2] Tile_X4Y5_LUT4AB/S2MID[3]
+ Tile_X4Y5_LUT4AB/S2MID[4] Tile_X4Y5_LUT4AB/S2MID[5] Tile_X4Y5_LUT4AB/S2MID[6] Tile_X4Y5_LUT4AB/S2MID[7]
+ Tile_X4Y6_LUT4AB/S4END[0] Tile_X4Y6_LUT4AB/S4END[10] Tile_X4Y6_LUT4AB/S4END[11]
+ Tile_X4Y6_LUT4AB/S4END[12] Tile_X4Y6_LUT4AB/S4END[13] Tile_X4Y6_LUT4AB/S4END[14]
+ Tile_X4Y6_LUT4AB/S4END[15] Tile_X4Y6_LUT4AB/S4END[1] Tile_X4Y6_LUT4AB/S4END[2] Tile_X4Y6_LUT4AB/S4END[3]
+ Tile_X4Y6_LUT4AB/S4END[4] Tile_X4Y6_LUT4AB/S4END[5] Tile_X4Y6_LUT4AB/S4END[6] Tile_X4Y6_LUT4AB/S4END[7]
+ Tile_X4Y6_LUT4AB/S4END[8] Tile_X4Y6_LUT4AB/S4END[9] Tile_X4Y5_LUT4AB/S4END[0] Tile_X4Y5_LUT4AB/S4END[10]
+ Tile_X4Y5_LUT4AB/S4END[11] Tile_X4Y5_LUT4AB/S4END[12] Tile_X4Y5_LUT4AB/S4END[13]
+ Tile_X4Y5_LUT4AB/S4END[14] Tile_X4Y5_LUT4AB/S4END[15] Tile_X4Y5_LUT4AB/S4END[1]
+ Tile_X4Y5_LUT4AB/S4END[2] Tile_X4Y5_LUT4AB/S4END[3] Tile_X4Y5_LUT4AB/S4END[4] Tile_X4Y5_LUT4AB/S4END[5]
+ Tile_X4Y5_LUT4AB/S4END[6] Tile_X4Y5_LUT4AB/S4END[7] Tile_X4Y5_LUT4AB/S4END[8] Tile_X4Y5_LUT4AB/S4END[9]
+ Tile_X4Y6_LUT4AB/SS4END[0] Tile_X4Y6_LUT4AB/SS4END[10] Tile_X4Y6_LUT4AB/SS4END[11]
+ Tile_X4Y6_LUT4AB/SS4END[12] Tile_X4Y6_LUT4AB/SS4END[13] Tile_X4Y6_LUT4AB/SS4END[14]
+ Tile_X4Y6_LUT4AB/SS4END[15] Tile_X4Y6_LUT4AB/SS4END[1] Tile_X4Y6_LUT4AB/SS4END[2]
+ Tile_X4Y6_LUT4AB/SS4END[3] Tile_X4Y6_LUT4AB/SS4END[4] Tile_X4Y6_LUT4AB/SS4END[5]
+ Tile_X4Y6_LUT4AB/SS4END[6] Tile_X4Y6_LUT4AB/SS4END[7] Tile_X4Y6_LUT4AB/SS4END[8]
+ Tile_X4Y6_LUT4AB/SS4END[9] Tile_X4Y5_LUT4AB/SS4END[0] Tile_X4Y5_LUT4AB/SS4END[10]
+ Tile_X4Y5_LUT4AB/SS4END[11] Tile_X4Y5_LUT4AB/SS4END[12] Tile_X4Y5_LUT4AB/SS4END[13]
+ Tile_X4Y5_LUT4AB/SS4END[14] Tile_X4Y5_LUT4AB/SS4END[15] Tile_X4Y5_LUT4AB/SS4END[1]
+ Tile_X4Y5_LUT4AB/SS4END[2] Tile_X4Y5_LUT4AB/SS4END[3] Tile_X4Y5_LUT4AB/SS4END[4]
+ Tile_X4Y5_LUT4AB/SS4END[5] Tile_X4Y5_LUT4AB/SS4END[6] Tile_X4Y5_LUT4AB/SS4END[7]
+ Tile_X4Y5_LUT4AB/SS4END[8] Tile_X4Y5_LUT4AB/SS4END[9] Tile_X4Y5_LUT4AB/UserCLK Tile_X4Y4_LUT4AB/UserCLK
+ VGND VPWR Tile_X4Y5_LUT4AB/W1BEG[0] Tile_X4Y5_LUT4AB/W1BEG[1] Tile_X4Y5_LUT4AB/W1BEG[2]
+ Tile_X4Y5_LUT4AB/W1BEG[3] Tile_X4Y5_LUT4AB/W1END[0] Tile_X4Y5_LUT4AB/W1END[1] Tile_X4Y5_LUT4AB/W1END[2]
+ Tile_X4Y5_LUT4AB/W1END[3] Tile_X4Y5_LUT4AB/W2BEG[0] Tile_X4Y5_LUT4AB/W2BEG[1] Tile_X4Y5_LUT4AB/W2BEG[2]
+ Tile_X4Y5_LUT4AB/W2BEG[3] Tile_X4Y5_LUT4AB/W2BEG[4] Tile_X4Y5_LUT4AB/W2BEG[5] Tile_X4Y5_LUT4AB/W2BEG[6]
+ Tile_X4Y5_LUT4AB/W2BEG[7] Tile_X3Y5_LUT4AB/W2END[0] Tile_X3Y5_LUT4AB/W2END[1] Tile_X3Y5_LUT4AB/W2END[2]
+ Tile_X3Y5_LUT4AB/W2END[3] Tile_X3Y5_LUT4AB/W2END[4] Tile_X3Y5_LUT4AB/W2END[5] Tile_X3Y5_LUT4AB/W2END[6]
+ Tile_X3Y5_LUT4AB/W2END[7] Tile_X4Y5_LUT4AB/W2END[0] Tile_X4Y5_LUT4AB/W2END[1] Tile_X4Y5_LUT4AB/W2END[2]
+ Tile_X4Y5_LUT4AB/W2END[3] Tile_X4Y5_LUT4AB/W2END[4] Tile_X4Y5_LUT4AB/W2END[5] Tile_X4Y5_LUT4AB/W2END[6]
+ Tile_X4Y5_LUT4AB/W2END[7] Tile_X4Y5_LUT4AB/W2MID[0] Tile_X4Y5_LUT4AB/W2MID[1] Tile_X4Y5_LUT4AB/W2MID[2]
+ Tile_X4Y5_LUT4AB/W2MID[3] Tile_X4Y5_LUT4AB/W2MID[4] Tile_X4Y5_LUT4AB/W2MID[5] Tile_X4Y5_LUT4AB/W2MID[6]
+ Tile_X4Y5_LUT4AB/W2MID[7] Tile_X4Y5_LUT4AB/W6BEG[0] Tile_X4Y5_LUT4AB/W6BEG[10] Tile_X4Y5_LUT4AB/W6BEG[11]
+ Tile_X4Y5_LUT4AB/W6BEG[1] Tile_X4Y5_LUT4AB/W6BEG[2] Tile_X4Y5_LUT4AB/W6BEG[3] Tile_X4Y5_LUT4AB/W6BEG[4]
+ Tile_X4Y5_LUT4AB/W6BEG[5] Tile_X4Y5_LUT4AB/W6BEG[6] Tile_X4Y5_LUT4AB/W6BEG[7] Tile_X4Y5_LUT4AB/W6BEG[8]
+ Tile_X4Y5_LUT4AB/W6BEG[9] Tile_X4Y5_LUT4AB/W6END[0] Tile_X4Y5_LUT4AB/W6END[10] Tile_X4Y5_LUT4AB/W6END[11]
+ Tile_X4Y5_LUT4AB/W6END[1] Tile_X4Y5_LUT4AB/W6END[2] Tile_X4Y5_LUT4AB/W6END[3] Tile_X4Y5_LUT4AB/W6END[4]
+ Tile_X4Y5_LUT4AB/W6END[5] Tile_X4Y5_LUT4AB/W6END[6] Tile_X4Y5_LUT4AB/W6END[7] Tile_X4Y5_LUT4AB/W6END[8]
+ Tile_X4Y5_LUT4AB/W6END[9] Tile_X4Y5_LUT4AB/WW4BEG[0] Tile_X4Y5_LUT4AB/WW4BEG[10]
+ Tile_X4Y5_LUT4AB/WW4BEG[11] Tile_X4Y5_LUT4AB/WW4BEG[12] Tile_X4Y5_LUT4AB/WW4BEG[13]
+ Tile_X4Y5_LUT4AB/WW4BEG[14] Tile_X4Y5_LUT4AB/WW4BEG[15] Tile_X4Y5_LUT4AB/WW4BEG[1]
+ Tile_X4Y5_LUT4AB/WW4BEG[2] Tile_X4Y5_LUT4AB/WW4BEG[3] Tile_X4Y5_LUT4AB/WW4BEG[4]
+ Tile_X4Y5_LUT4AB/WW4BEG[5] Tile_X4Y5_LUT4AB/WW4BEG[6] Tile_X4Y5_LUT4AB/WW4BEG[7]
+ Tile_X4Y5_LUT4AB/WW4BEG[8] Tile_X4Y5_LUT4AB/WW4BEG[9] Tile_X4Y5_LUT4AB/WW4END[0]
+ Tile_X4Y5_LUT4AB/WW4END[10] Tile_X4Y5_LUT4AB/WW4END[11] Tile_X4Y5_LUT4AB/WW4END[12]
+ Tile_X4Y5_LUT4AB/WW4END[13] Tile_X4Y5_LUT4AB/WW4END[14] Tile_X4Y5_LUT4AB/WW4END[15]
+ Tile_X4Y5_LUT4AB/WW4END[1] Tile_X4Y5_LUT4AB/WW4END[2] Tile_X4Y5_LUT4AB/WW4END[3]
+ Tile_X4Y5_LUT4AB/WW4END[4] Tile_X4Y5_LUT4AB/WW4END[5] Tile_X4Y5_LUT4AB/WW4END[6]
+ Tile_X4Y5_LUT4AB/WW4END[7] Tile_X4Y5_LUT4AB/WW4END[8] Tile_X4Y5_LUT4AB/WW4END[9]
+ LUT4AB
XTile_X0Y9_SW_term FrameData[288] FrameData[298] FrameData[299] FrameData[300] FrameData[301]
+ FrameData[302] FrameData[303] FrameData[304] FrameData[305] FrameData[306] FrameData[307]
+ FrameData[289] FrameData[308] FrameData[309] FrameData[310] FrameData[311] FrameData[312]
+ FrameData[313] FrameData[314] FrameData[315] FrameData[316] FrameData[317] FrameData[290]
+ FrameData[318] FrameData[319] FrameData[291] FrameData[292] FrameData[293] FrameData[294]
+ FrameData[295] FrameData[296] FrameData[297] Tile_X1Y9_S_IO4/FrameData[0] Tile_X1Y9_S_IO4/FrameData[10]
+ Tile_X1Y9_S_IO4/FrameData[11] Tile_X1Y9_S_IO4/FrameData[12] Tile_X1Y9_S_IO4/FrameData[13]
+ Tile_X1Y9_S_IO4/FrameData[14] Tile_X1Y9_S_IO4/FrameData[15] Tile_X1Y9_S_IO4/FrameData[16]
+ Tile_X1Y9_S_IO4/FrameData[17] Tile_X1Y9_S_IO4/FrameData[18] Tile_X1Y9_S_IO4/FrameData[19]
+ Tile_X1Y9_S_IO4/FrameData[1] Tile_X1Y9_S_IO4/FrameData[20] Tile_X1Y9_S_IO4/FrameData[21]
+ Tile_X1Y9_S_IO4/FrameData[22] Tile_X1Y9_S_IO4/FrameData[23] Tile_X1Y9_S_IO4/FrameData[24]
+ Tile_X1Y9_S_IO4/FrameData[25] Tile_X1Y9_S_IO4/FrameData[26] Tile_X1Y9_S_IO4/FrameData[27]
+ Tile_X1Y9_S_IO4/FrameData[28] Tile_X1Y9_S_IO4/FrameData[29] Tile_X1Y9_S_IO4/FrameData[2]
+ Tile_X1Y9_S_IO4/FrameData[30] Tile_X1Y9_S_IO4/FrameData[31] Tile_X1Y9_S_IO4/FrameData[3]
+ Tile_X1Y9_S_IO4/FrameData[4] Tile_X1Y9_S_IO4/FrameData[5] Tile_X1Y9_S_IO4/FrameData[6]
+ Tile_X1Y9_S_IO4/FrameData[7] Tile_X1Y9_S_IO4/FrameData[8] Tile_X1Y9_S_IO4/FrameData[9]
+ FrameStrobe[0] FrameStrobe[10] FrameStrobe[11] FrameStrobe[12] FrameStrobe[13] FrameStrobe[14]
+ FrameStrobe[15] FrameStrobe[16] FrameStrobe[17] FrameStrobe[18] FrameStrobe[19]
+ FrameStrobe[1] FrameStrobe[2] FrameStrobe[3] FrameStrobe[4] FrameStrobe[5] FrameStrobe[6]
+ FrameStrobe[7] FrameStrobe[8] FrameStrobe[9] Tile_X0Y8_W_TT_IF/FrameStrobe[0] Tile_X0Y8_W_TT_IF/FrameStrobe[10]
+ Tile_X0Y8_W_TT_IF/FrameStrobe[11] Tile_X0Y8_W_TT_IF/FrameStrobe[12] Tile_X0Y8_W_TT_IF/FrameStrobe[13]
+ Tile_X0Y8_W_TT_IF/FrameStrobe[14] Tile_X0Y8_W_TT_IF/FrameStrobe[15] Tile_X0Y8_W_TT_IF/FrameStrobe[16]
+ Tile_X0Y8_W_TT_IF/FrameStrobe[17] Tile_X0Y8_W_TT_IF/FrameStrobe[18] Tile_X0Y8_W_TT_IF/FrameStrobe[19]
+ Tile_X0Y8_W_TT_IF/FrameStrobe[1] Tile_X0Y8_W_TT_IF/FrameStrobe[2] Tile_X0Y8_W_TT_IF/FrameStrobe[3]
+ Tile_X0Y8_W_TT_IF/FrameStrobe[4] Tile_X0Y8_W_TT_IF/FrameStrobe[5] Tile_X0Y8_W_TT_IF/FrameStrobe[6]
+ Tile_X0Y8_W_TT_IF/FrameStrobe[7] Tile_X0Y8_W_TT_IF/FrameStrobe[8] Tile_X0Y8_W_TT_IF/FrameStrobe[9]
+ Tile_X0Y9_SW_term/N1BEG[0] Tile_X0Y9_SW_term/N1BEG[1] Tile_X0Y9_SW_term/N1BEG[2]
+ Tile_X0Y9_SW_term/N1BEG[3] Tile_X0Y9_SW_term/N2BEG[0] Tile_X0Y9_SW_term/N2BEG[1]
+ Tile_X0Y9_SW_term/N2BEG[2] Tile_X0Y9_SW_term/N2BEG[3] Tile_X0Y9_SW_term/N2BEG[4]
+ Tile_X0Y9_SW_term/N2BEG[5] Tile_X0Y9_SW_term/N2BEG[6] Tile_X0Y9_SW_term/N2BEG[7]
+ Tile_X0Y8_W_TT_IF/N2END[0] Tile_X0Y8_W_TT_IF/N2END[1] Tile_X0Y8_W_TT_IF/N2END[2]
+ Tile_X0Y8_W_TT_IF/N2END[3] Tile_X0Y8_W_TT_IF/N2END[4] Tile_X0Y8_W_TT_IF/N2END[5]
+ Tile_X0Y8_W_TT_IF/N2END[6] Tile_X0Y8_W_TT_IF/N2END[7] Tile_X0Y9_SW_term/N4BEG[0]
+ Tile_X0Y9_SW_term/N4BEG[10] Tile_X0Y9_SW_term/N4BEG[11] Tile_X0Y9_SW_term/N4BEG[12]
+ Tile_X0Y9_SW_term/N4BEG[13] Tile_X0Y9_SW_term/N4BEG[14] Tile_X0Y9_SW_term/N4BEG[15]
+ Tile_X0Y9_SW_term/N4BEG[1] Tile_X0Y9_SW_term/N4BEG[2] Tile_X0Y9_SW_term/N4BEG[3]
+ Tile_X0Y9_SW_term/N4BEG[4] Tile_X0Y9_SW_term/N4BEG[5] Tile_X0Y9_SW_term/N4BEG[6]
+ Tile_X0Y9_SW_term/N4BEG[7] Tile_X0Y9_SW_term/N4BEG[8] Tile_X0Y9_SW_term/N4BEG[9]
+ Tile_X0Y9_SW_term/S1END[0] Tile_X0Y9_SW_term/S1END[1] Tile_X0Y9_SW_term/S1END[2]
+ Tile_X0Y9_SW_term/S1END[3] Tile_X0Y9_SW_term/S2END[0] Tile_X0Y9_SW_term/S2END[1]
+ Tile_X0Y9_SW_term/S2END[2] Tile_X0Y9_SW_term/S2END[3] Tile_X0Y9_SW_term/S2END[4]
+ Tile_X0Y9_SW_term/S2END[5] Tile_X0Y9_SW_term/S2END[6] Tile_X0Y9_SW_term/S2END[7]
+ Tile_X0Y9_SW_term/S2MID[0] Tile_X0Y9_SW_term/S2MID[1] Tile_X0Y9_SW_term/S2MID[2]
+ Tile_X0Y9_SW_term/S2MID[3] Tile_X0Y9_SW_term/S2MID[4] Tile_X0Y9_SW_term/S2MID[5]
+ Tile_X0Y9_SW_term/S2MID[6] Tile_X0Y9_SW_term/S2MID[7] Tile_X0Y9_SW_term/S4END[0]
+ Tile_X0Y9_SW_term/S4END[10] Tile_X0Y9_SW_term/S4END[11] Tile_X0Y9_SW_term/S4END[12]
+ Tile_X0Y9_SW_term/S4END[13] Tile_X0Y9_SW_term/S4END[14] Tile_X0Y9_SW_term/S4END[15]
+ Tile_X0Y9_SW_term/S4END[1] Tile_X0Y9_SW_term/S4END[2] Tile_X0Y9_SW_term/S4END[3]
+ Tile_X0Y9_SW_term/S4END[4] Tile_X0Y9_SW_term/S4END[5] Tile_X0Y9_SW_term/S4END[6]
+ Tile_X0Y9_SW_term/S4END[7] Tile_X0Y9_SW_term/S4END[8] Tile_X0Y9_SW_term/S4END[9]
+ UserCLK Tile_X0Y8_W_TT_IF/UserCLK VGND VPWR SW_term
XTile_X2Y2_LUT4AB Tile_X2Y3_LUT4AB/Co Tile_X2Y2_LUT4AB/Co Tile_X3Y2_LUT4AB/E1END[0]
+ Tile_X3Y2_LUT4AB/E1END[1] Tile_X3Y2_LUT4AB/E1END[2] Tile_X3Y2_LUT4AB/E1END[3] Tile_X2Y2_LUT4AB/E1END[0]
+ Tile_X2Y2_LUT4AB/E1END[1] Tile_X2Y2_LUT4AB/E1END[2] Tile_X2Y2_LUT4AB/E1END[3] Tile_X3Y2_LUT4AB/E2MID[0]
+ Tile_X3Y2_LUT4AB/E2MID[1] Tile_X3Y2_LUT4AB/E2MID[2] Tile_X3Y2_LUT4AB/E2MID[3] Tile_X3Y2_LUT4AB/E2MID[4]
+ Tile_X3Y2_LUT4AB/E2MID[5] Tile_X3Y2_LUT4AB/E2MID[6] Tile_X3Y2_LUT4AB/E2MID[7] Tile_X3Y2_LUT4AB/E2END[0]
+ Tile_X3Y2_LUT4AB/E2END[1] Tile_X3Y2_LUT4AB/E2END[2] Tile_X3Y2_LUT4AB/E2END[3] Tile_X3Y2_LUT4AB/E2END[4]
+ Tile_X3Y2_LUT4AB/E2END[5] Tile_X3Y2_LUT4AB/E2END[6] Tile_X3Y2_LUT4AB/E2END[7] Tile_X2Y2_LUT4AB/E2END[0]
+ Tile_X2Y2_LUT4AB/E2END[1] Tile_X2Y2_LUT4AB/E2END[2] Tile_X2Y2_LUT4AB/E2END[3] Tile_X2Y2_LUT4AB/E2END[4]
+ Tile_X2Y2_LUT4AB/E2END[5] Tile_X2Y2_LUT4AB/E2END[6] Tile_X2Y2_LUT4AB/E2END[7] Tile_X2Y2_LUT4AB/E2MID[0]
+ Tile_X2Y2_LUT4AB/E2MID[1] Tile_X2Y2_LUT4AB/E2MID[2] Tile_X2Y2_LUT4AB/E2MID[3] Tile_X2Y2_LUT4AB/E2MID[4]
+ Tile_X2Y2_LUT4AB/E2MID[5] Tile_X2Y2_LUT4AB/E2MID[6] Tile_X2Y2_LUT4AB/E2MID[7] Tile_X3Y2_LUT4AB/E6END[0]
+ Tile_X3Y2_LUT4AB/E6END[10] Tile_X3Y2_LUT4AB/E6END[11] Tile_X3Y2_LUT4AB/E6END[1]
+ Tile_X3Y2_LUT4AB/E6END[2] Tile_X3Y2_LUT4AB/E6END[3] Tile_X3Y2_LUT4AB/E6END[4] Tile_X3Y2_LUT4AB/E6END[5]
+ Tile_X3Y2_LUT4AB/E6END[6] Tile_X3Y2_LUT4AB/E6END[7] Tile_X3Y2_LUT4AB/E6END[8] Tile_X3Y2_LUT4AB/E6END[9]
+ Tile_X2Y2_LUT4AB/E6END[0] Tile_X2Y2_LUT4AB/E6END[10] Tile_X2Y2_LUT4AB/E6END[11]
+ Tile_X2Y2_LUT4AB/E6END[1] Tile_X2Y2_LUT4AB/E6END[2] Tile_X2Y2_LUT4AB/E6END[3] Tile_X2Y2_LUT4AB/E6END[4]
+ Tile_X2Y2_LUT4AB/E6END[5] Tile_X2Y2_LUT4AB/E6END[6] Tile_X2Y2_LUT4AB/E6END[7] Tile_X2Y2_LUT4AB/E6END[8]
+ Tile_X2Y2_LUT4AB/E6END[9] Tile_X3Y2_LUT4AB/EE4END[0] Tile_X3Y2_LUT4AB/EE4END[10]
+ Tile_X3Y2_LUT4AB/EE4END[11] Tile_X3Y2_LUT4AB/EE4END[12] Tile_X3Y2_LUT4AB/EE4END[13]
+ Tile_X3Y2_LUT4AB/EE4END[14] Tile_X3Y2_LUT4AB/EE4END[15] Tile_X3Y2_LUT4AB/EE4END[1]
+ Tile_X3Y2_LUT4AB/EE4END[2] Tile_X3Y2_LUT4AB/EE4END[3] Tile_X3Y2_LUT4AB/EE4END[4]
+ Tile_X3Y2_LUT4AB/EE4END[5] Tile_X3Y2_LUT4AB/EE4END[6] Tile_X3Y2_LUT4AB/EE4END[7]
+ Tile_X3Y2_LUT4AB/EE4END[8] Tile_X3Y2_LUT4AB/EE4END[9] Tile_X2Y2_LUT4AB/EE4END[0]
+ Tile_X2Y2_LUT4AB/EE4END[10] Tile_X2Y2_LUT4AB/EE4END[11] Tile_X2Y2_LUT4AB/EE4END[12]
+ Tile_X2Y2_LUT4AB/EE4END[13] Tile_X2Y2_LUT4AB/EE4END[14] Tile_X2Y2_LUT4AB/EE4END[15]
+ Tile_X2Y2_LUT4AB/EE4END[1] Tile_X2Y2_LUT4AB/EE4END[2] Tile_X2Y2_LUT4AB/EE4END[3]
+ Tile_X2Y2_LUT4AB/EE4END[4] Tile_X2Y2_LUT4AB/EE4END[5] Tile_X2Y2_LUT4AB/EE4END[6]
+ Tile_X2Y2_LUT4AB/EE4END[7] Tile_X2Y2_LUT4AB/EE4END[8] Tile_X2Y2_LUT4AB/EE4END[9]
+ Tile_X2Y2_LUT4AB/FrameData[0] Tile_X2Y2_LUT4AB/FrameData[10] Tile_X2Y2_LUT4AB/FrameData[11]
+ Tile_X2Y2_LUT4AB/FrameData[12] Tile_X2Y2_LUT4AB/FrameData[13] Tile_X2Y2_LUT4AB/FrameData[14]
+ Tile_X2Y2_LUT4AB/FrameData[15] Tile_X2Y2_LUT4AB/FrameData[16] Tile_X2Y2_LUT4AB/FrameData[17]
+ Tile_X2Y2_LUT4AB/FrameData[18] Tile_X2Y2_LUT4AB/FrameData[19] Tile_X2Y2_LUT4AB/FrameData[1]
+ Tile_X2Y2_LUT4AB/FrameData[20] Tile_X2Y2_LUT4AB/FrameData[21] Tile_X2Y2_LUT4AB/FrameData[22]
+ Tile_X2Y2_LUT4AB/FrameData[23] Tile_X2Y2_LUT4AB/FrameData[24] Tile_X2Y2_LUT4AB/FrameData[25]
+ Tile_X2Y2_LUT4AB/FrameData[26] Tile_X2Y2_LUT4AB/FrameData[27] Tile_X2Y2_LUT4AB/FrameData[28]
+ Tile_X2Y2_LUT4AB/FrameData[29] Tile_X2Y2_LUT4AB/FrameData[2] Tile_X2Y2_LUT4AB/FrameData[30]
+ Tile_X2Y2_LUT4AB/FrameData[31] Tile_X2Y2_LUT4AB/FrameData[3] Tile_X2Y2_LUT4AB/FrameData[4]
+ Tile_X2Y2_LUT4AB/FrameData[5] Tile_X2Y2_LUT4AB/FrameData[6] Tile_X2Y2_LUT4AB/FrameData[7]
+ Tile_X2Y2_LUT4AB/FrameData[8] Tile_X2Y2_LUT4AB/FrameData[9] Tile_X3Y2_LUT4AB/FrameData[0]
+ Tile_X3Y2_LUT4AB/FrameData[10] Tile_X3Y2_LUT4AB/FrameData[11] Tile_X3Y2_LUT4AB/FrameData[12]
+ Tile_X3Y2_LUT4AB/FrameData[13] Tile_X3Y2_LUT4AB/FrameData[14] Tile_X3Y2_LUT4AB/FrameData[15]
+ Tile_X3Y2_LUT4AB/FrameData[16] Tile_X3Y2_LUT4AB/FrameData[17] Tile_X3Y2_LUT4AB/FrameData[18]
+ Tile_X3Y2_LUT4AB/FrameData[19] Tile_X3Y2_LUT4AB/FrameData[1] Tile_X3Y2_LUT4AB/FrameData[20]
+ Tile_X3Y2_LUT4AB/FrameData[21] Tile_X3Y2_LUT4AB/FrameData[22] Tile_X3Y2_LUT4AB/FrameData[23]
+ Tile_X3Y2_LUT4AB/FrameData[24] Tile_X3Y2_LUT4AB/FrameData[25] Tile_X3Y2_LUT4AB/FrameData[26]
+ Tile_X3Y2_LUT4AB/FrameData[27] Tile_X3Y2_LUT4AB/FrameData[28] Tile_X3Y2_LUT4AB/FrameData[29]
+ Tile_X3Y2_LUT4AB/FrameData[2] Tile_X3Y2_LUT4AB/FrameData[30] Tile_X3Y2_LUT4AB/FrameData[31]
+ Tile_X3Y2_LUT4AB/FrameData[3] Tile_X3Y2_LUT4AB/FrameData[4] Tile_X3Y2_LUT4AB/FrameData[5]
+ Tile_X3Y2_LUT4AB/FrameData[6] Tile_X3Y2_LUT4AB/FrameData[7] Tile_X3Y2_LUT4AB/FrameData[8]
+ Tile_X3Y2_LUT4AB/FrameData[9] Tile_X2Y2_LUT4AB/FrameStrobe[0] Tile_X2Y2_LUT4AB/FrameStrobe[10]
+ Tile_X2Y2_LUT4AB/FrameStrobe[11] Tile_X2Y2_LUT4AB/FrameStrobe[12] Tile_X2Y2_LUT4AB/FrameStrobe[13]
+ Tile_X2Y2_LUT4AB/FrameStrobe[14] Tile_X2Y2_LUT4AB/FrameStrobe[15] Tile_X2Y2_LUT4AB/FrameStrobe[16]
+ Tile_X2Y2_LUT4AB/FrameStrobe[17] Tile_X2Y2_LUT4AB/FrameStrobe[18] Tile_X2Y2_LUT4AB/FrameStrobe[19]
+ Tile_X2Y2_LUT4AB/FrameStrobe[1] Tile_X2Y2_LUT4AB/FrameStrobe[2] Tile_X2Y2_LUT4AB/FrameStrobe[3]
+ Tile_X2Y2_LUT4AB/FrameStrobe[4] Tile_X2Y2_LUT4AB/FrameStrobe[5] Tile_X2Y2_LUT4AB/FrameStrobe[6]
+ Tile_X2Y2_LUT4AB/FrameStrobe[7] Tile_X2Y2_LUT4AB/FrameStrobe[8] Tile_X2Y2_LUT4AB/FrameStrobe[9]
+ Tile_X2Y1_LUT4AB/FrameStrobe[0] Tile_X2Y1_LUT4AB/FrameStrobe[10] Tile_X2Y1_LUT4AB/FrameStrobe[11]
+ Tile_X2Y1_LUT4AB/FrameStrobe[12] Tile_X2Y1_LUT4AB/FrameStrobe[13] Tile_X2Y1_LUT4AB/FrameStrobe[14]
+ Tile_X2Y1_LUT4AB/FrameStrobe[15] Tile_X2Y1_LUT4AB/FrameStrobe[16] Tile_X2Y1_LUT4AB/FrameStrobe[17]
+ Tile_X2Y1_LUT4AB/FrameStrobe[18] Tile_X2Y1_LUT4AB/FrameStrobe[19] Tile_X2Y1_LUT4AB/FrameStrobe[1]
+ Tile_X2Y1_LUT4AB/FrameStrobe[2] Tile_X2Y1_LUT4AB/FrameStrobe[3] Tile_X2Y1_LUT4AB/FrameStrobe[4]
+ Tile_X2Y1_LUT4AB/FrameStrobe[5] Tile_X2Y1_LUT4AB/FrameStrobe[6] Tile_X2Y1_LUT4AB/FrameStrobe[7]
+ Tile_X2Y1_LUT4AB/FrameStrobe[8] Tile_X2Y1_LUT4AB/FrameStrobe[9] Tile_X2Y2_LUT4AB/N1BEG[0]
+ Tile_X2Y2_LUT4AB/N1BEG[1] Tile_X2Y2_LUT4AB/N1BEG[2] Tile_X2Y2_LUT4AB/N1BEG[3] Tile_X2Y3_LUT4AB/N1BEG[0]
+ Tile_X2Y3_LUT4AB/N1BEG[1] Tile_X2Y3_LUT4AB/N1BEG[2] Tile_X2Y3_LUT4AB/N1BEG[3] Tile_X2Y2_LUT4AB/N2BEG[0]
+ Tile_X2Y2_LUT4AB/N2BEG[1] Tile_X2Y2_LUT4AB/N2BEG[2] Tile_X2Y2_LUT4AB/N2BEG[3] Tile_X2Y2_LUT4AB/N2BEG[4]
+ Tile_X2Y2_LUT4AB/N2BEG[5] Tile_X2Y2_LUT4AB/N2BEG[6] Tile_X2Y2_LUT4AB/N2BEG[7] Tile_X2Y1_LUT4AB/N2END[0]
+ Tile_X2Y1_LUT4AB/N2END[1] Tile_X2Y1_LUT4AB/N2END[2] Tile_X2Y1_LUT4AB/N2END[3] Tile_X2Y1_LUT4AB/N2END[4]
+ Tile_X2Y1_LUT4AB/N2END[5] Tile_X2Y1_LUT4AB/N2END[6] Tile_X2Y1_LUT4AB/N2END[7] Tile_X2Y2_LUT4AB/N2END[0]
+ Tile_X2Y2_LUT4AB/N2END[1] Tile_X2Y2_LUT4AB/N2END[2] Tile_X2Y2_LUT4AB/N2END[3] Tile_X2Y2_LUT4AB/N2END[4]
+ Tile_X2Y2_LUT4AB/N2END[5] Tile_X2Y2_LUT4AB/N2END[6] Tile_X2Y2_LUT4AB/N2END[7] Tile_X2Y3_LUT4AB/N2BEG[0]
+ Tile_X2Y3_LUT4AB/N2BEG[1] Tile_X2Y3_LUT4AB/N2BEG[2] Tile_X2Y3_LUT4AB/N2BEG[3] Tile_X2Y3_LUT4AB/N2BEG[4]
+ Tile_X2Y3_LUT4AB/N2BEG[5] Tile_X2Y3_LUT4AB/N2BEG[6] Tile_X2Y3_LUT4AB/N2BEG[7] Tile_X2Y2_LUT4AB/N4BEG[0]
+ Tile_X2Y2_LUT4AB/N4BEG[10] Tile_X2Y2_LUT4AB/N4BEG[11] Tile_X2Y2_LUT4AB/N4BEG[12]
+ Tile_X2Y2_LUT4AB/N4BEG[13] Tile_X2Y2_LUT4AB/N4BEG[14] Tile_X2Y2_LUT4AB/N4BEG[15]
+ Tile_X2Y2_LUT4AB/N4BEG[1] Tile_X2Y2_LUT4AB/N4BEG[2] Tile_X2Y2_LUT4AB/N4BEG[3] Tile_X2Y2_LUT4AB/N4BEG[4]
+ Tile_X2Y2_LUT4AB/N4BEG[5] Tile_X2Y2_LUT4AB/N4BEG[6] Tile_X2Y2_LUT4AB/N4BEG[7] Tile_X2Y2_LUT4AB/N4BEG[8]
+ Tile_X2Y2_LUT4AB/N4BEG[9] Tile_X2Y3_LUT4AB/N4BEG[0] Tile_X2Y3_LUT4AB/N4BEG[10] Tile_X2Y3_LUT4AB/N4BEG[11]
+ Tile_X2Y3_LUT4AB/N4BEG[12] Tile_X2Y3_LUT4AB/N4BEG[13] Tile_X2Y3_LUT4AB/N4BEG[14]
+ Tile_X2Y3_LUT4AB/N4BEG[15] Tile_X2Y3_LUT4AB/N4BEG[1] Tile_X2Y3_LUT4AB/N4BEG[2] Tile_X2Y3_LUT4AB/N4BEG[3]
+ Tile_X2Y3_LUT4AB/N4BEG[4] Tile_X2Y3_LUT4AB/N4BEG[5] Tile_X2Y3_LUT4AB/N4BEG[6] Tile_X2Y3_LUT4AB/N4BEG[7]
+ Tile_X2Y3_LUT4AB/N4BEG[8] Tile_X2Y3_LUT4AB/N4BEG[9] Tile_X2Y2_LUT4AB/NN4BEG[0] Tile_X2Y2_LUT4AB/NN4BEG[10]
+ Tile_X2Y2_LUT4AB/NN4BEG[11] Tile_X2Y2_LUT4AB/NN4BEG[12] Tile_X2Y2_LUT4AB/NN4BEG[13]
+ Tile_X2Y2_LUT4AB/NN4BEG[14] Tile_X2Y2_LUT4AB/NN4BEG[15] Tile_X2Y2_LUT4AB/NN4BEG[1]
+ Tile_X2Y2_LUT4AB/NN4BEG[2] Tile_X2Y2_LUT4AB/NN4BEG[3] Tile_X2Y2_LUT4AB/NN4BEG[4]
+ Tile_X2Y2_LUT4AB/NN4BEG[5] Tile_X2Y2_LUT4AB/NN4BEG[6] Tile_X2Y2_LUT4AB/NN4BEG[7]
+ Tile_X2Y2_LUT4AB/NN4BEG[8] Tile_X2Y2_LUT4AB/NN4BEG[9] Tile_X2Y3_LUT4AB/NN4BEG[0]
+ Tile_X2Y3_LUT4AB/NN4BEG[10] Tile_X2Y3_LUT4AB/NN4BEG[11] Tile_X2Y3_LUT4AB/NN4BEG[12]
+ Tile_X2Y3_LUT4AB/NN4BEG[13] Tile_X2Y3_LUT4AB/NN4BEG[14] Tile_X2Y3_LUT4AB/NN4BEG[15]
+ Tile_X2Y3_LUT4AB/NN4BEG[1] Tile_X2Y3_LUT4AB/NN4BEG[2] Tile_X2Y3_LUT4AB/NN4BEG[3]
+ Tile_X2Y3_LUT4AB/NN4BEG[4] Tile_X2Y3_LUT4AB/NN4BEG[5] Tile_X2Y3_LUT4AB/NN4BEG[6]
+ Tile_X2Y3_LUT4AB/NN4BEG[7] Tile_X2Y3_LUT4AB/NN4BEG[8] Tile_X2Y3_LUT4AB/NN4BEG[9]
+ Tile_X2Y3_LUT4AB/S1END[0] Tile_X2Y3_LUT4AB/S1END[1] Tile_X2Y3_LUT4AB/S1END[2] Tile_X2Y3_LUT4AB/S1END[3]
+ Tile_X2Y2_LUT4AB/S1END[0] Tile_X2Y2_LUT4AB/S1END[1] Tile_X2Y2_LUT4AB/S1END[2] Tile_X2Y2_LUT4AB/S1END[3]
+ Tile_X2Y3_LUT4AB/S2MID[0] Tile_X2Y3_LUT4AB/S2MID[1] Tile_X2Y3_LUT4AB/S2MID[2] Tile_X2Y3_LUT4AB/S2MID[3]
+ Tile_X2Y3_LUT4AB/S2MID[4] Tile_X2Y3_LUT4AB/S2MID[5] Tile_X2Y3_LUT4AB/S2MID[6] Tile_X2Y3_LUT4AB/S2MID[7]
+ Tile_X2Y3_LUT4AB/S2END[0] Tile_X2Y3_LUT4AB/S2END[1] Tile_X2Y3_LUT4AB/S2END[2] Tile_X2Y3_LUT4AB/S2END[3]
+ Tile_X2Y3_LUT4AB/S2END[4] Tile_X2Y3_LUT4AB/S2END[5] Tile_X2Y3_LUT4AB/S2END[6] Tile_X2Y3_LUT4AB/S2END[7]
+ Tile_X2Y2_LUT4AB/S2END[0] Tile_X2Y2_LUT4AB/S2END[1] Tile_X2Y2_LUT4AB/S2END[2] Tile_X2Y2_LUT4AB/S2END[3]
+ Tile_X2Y2_LUT4AB/S2END[4] Tile_X2Y2_LUT4AB/S2END[5] Tile_X2Y2_LUT4AB/S2END[6] Tile_X2Y2_LUT4AB/S2END[7]
+ Tile_X2Y2_LUT4AB/S2MID[0] Tile_X2Y2_LUT4AB/S2MID[1] Tile_X2Y2_LUT4AB/S2MID[2] Tile_X2Y2_LUT4AB/S2MID[3]
+ Tile_X2Y2_LUT4AB/S2MID[4] Tile_X2Y2_LUT4AB/S2MID[5] Tile_X2Y2_LUT4AB/S2MID[6] Tile_X2Y2_LUT4AB/S2MID[7]
+ Tile_X2Y3_LUT4AB/S4END[0] Tile_X2Y3_LUT4AB/S4END[10] Tile_X2Y3_LUT4AB/S4END[11]
+ Tile_X2Y3_LUT4AB/S4END[12] Tile_X2Y3_LUT4AB/S4END[13] Tile_X2Y3_LUT4AB/S4END[14]
+ Tile_X2Y3_LUT4AB/S4END[15] Tile_X2Y3_LUT4AB/S4END[1] Tile_X2Y3_LUT4AB/S4END[2] Tile_X2Y3_LUT4AB/S4END[3]
+ Tile_X2Y3_LUT4AB/S4END[4] Tile_X2Y3_LUT4AB/S4END[5] Tile_X2Y3_LUT4AB/S4END[6] Tile_X2Y3_LUT4AB/S4END[7]
+ Tile_X2Y3_LUT4AB/S4END[8] Tile_X2Y3_LUT4AB/S4END[9] Tile_X2Y2_LUT4AB/S4END[0] Tile_X2Y2_LUT4AB/S4END[10]
+ Tile_X2Y2_LUT4AB/S4END[11] Tile_X2Y2_LUT4AB/S4END[12] Tile_X2Y2_LUT4AB/S4END[13]
+ Tile_X2Y2_LUT4AB/S4END[14] Tile_X2Y2_LUT4AB/S4END[15] Tile_X2Y2_LUT4AB/S4END[1]
+ Tile_X2Y2_LUT4AB/S4END[2] Tile_X2Y2_LUT4AB/S4END[3] Tile_X2Y2_LUT4AB/S4END[4] Tile_X2Y2_LUT4AB/S4END[5]
+ Tile_X2Y2_LUT4AB/S4END[6] Tile_X2Y2_LUT4AB/S4END[7] Tile_X2Y2_LUT4AB/S4END[8] Tile_X2Y2_LUT4AB/S4END[9]
+ Tile_X2Y3_LUT4AB/SS4END[0] Tile_X2Y3_LUT4AB/SS4END[10] Tile_X2Y3_LUT4AB/SS4END[11]
+ Tile_X2Y3_LUT4AB/SS4END[12] Tile_X2Y3_LUT4AB/SS4END[13] Tile_X2Y3_LUT4AB/SS4END[14]
+ Tile_X2Y3_LUT4AB/SS4END[15] Tile_X2Y3_LUT4AB/SS4END[1] Tile_X2Y3_LUT4AB/SS4END[2]
+ Tile_X2Y3_LUT4AB/SS4END[3] Tile_X2Y3_LUT4AB/SS4END[4] Tile_X2Y3_LUT4AB/SS4END[5]
+ Tile_X2Y3_LUT4AB/SS4END[6] Tile_X2Y3_LUT4AB/SS4END[7] Tile_X2Y3_LUT4AB/SS4END[8]
+ Tile_X2Y3_LUT4AB/SS4END[9] Tile_X2Y2_LUT4AB/SS4END[0] Tile_X2Y2_LUT4AB/SS4END[10]
+ Tile_X2Y2_LUT4AB/SS4END[11] Tile_X2Y2_LUT4AB/SS4END[12] Tile_X2Y2_LUT4AB/SS4END[13]
+ Tile_X2Y2_LUT4AB/SS4END[14] Tile_X2Y2_LUT4AB/SS4END[15] Tile_X2Y2_LUT4AB/SS4END[1]
+ Tile_X2Y2_LUT4AB/SS4END[2] Tile_X2Y2_LUT4AB/SS4END[3] Tile_X2Y2_LUT4AB/SS4END[4]
+ Tile_X2Y2_LUT4AB/SS4END[5] Tile_X2Y2_LUT4AB/SS4END[6] Tile_X2Y2_LUT4AB/SS4END[7]
+ Tile_X2Y2_LUT4AB/SS4END[8] Tile_X2Y2_LUT4AB/SS4END[9] Tile_X2Y2_LUT4AB/UserCLK Tile_X2Y1_LUT4AB/UserCLK
+ VGND VPWR Tile_X2Y2_LUT4AB/W1BEG[0] Tile_X2Y2_LUT4AB/W1BEG[1] Tile_X2Y2_LUT4AB/W1BEG[2]
+ Tile_X2Y2_LUT4AB/W1BEG[3] Tile_X3Y2_LUT4AB/W1BEG[0] Tile_X3Y2_LUT4AB/W1BEG[1] Tile_X3Y2_LUT4AB/W1BEG[2]
+ Tile_X3Y2_LUT4AB/W1BEG[3] Tile_X2Y2_LUT4AB/W2BEG[0] Tile_X2Y2_LUT4AB/W2BEG[1] Tile_X2Y2_LUT4AB/W2BEG[2]
+ Tile_X2Y2_LUT4AB/W2BEG[3] Tile_X2Y2_LUT4AB/W2BEG[4] Tile_X2Y2_LUT4AB/W2BEG[5] Tile_X2Y2_LUT4AB/W2BEG[6]
+ Tile_X2Y2_LUT4AB/W2BEG[7] Tile_X1Y2_LUT4AB/W2END[0] Tile_X1Y2_LUT4AB/W2END[1] Tile_X1Y2_LUT4AB/W2END[2]
+ Tile_X1Y2_LUT4AB/W2END[3] Tile_X1Y2_LUT4AB/W2END[4] Tile_X1Y2_LUT4AB/W2END[5] Tile_X1Y2_LUT4AB/W2END[6]
+ Tile_X1Y2_LUT4AB/W2END[7] Tile_X2Y2_LUT4AB/W2END[0] Tile_X2Y2_LUT4AB/W2END[1] Tile_X2Y2_LUT4AB/W2END[2]
+ Tile_X2Y2_LUT4AB/W2END[3] Tile_X2Y2_LUT4AB/W2END[4] Tile_X2Y2_LUT4AB/W2END[5] Tile_X2Y2_LUT4AB/W2END[6]
+ Tile_X2Y2_LUT4AB/W2END[7] Tile_X3Y2_LUT4AB/W2BEG[0] Tile_X3Y2_LUT4AB/W2BEG[1] Tile_X3Y2_LUT4AB/W2BEG[2]
+ Tile_X3Y2_LUT4AB/W2BEG[3] Tile_X3Y2_LUT4AB/W2BEG[4] Tile_X3Y2_LUT4AB/W2BEG[5] Tile_X3Y2_LUT4AB/W2BEG[6]
+ Tile_X3Y2_LUT4AB/W2BEG[7] Tile_X2Y2_LUT4AB/W6BEG[0] Tile_X2Y2_LUT4AB/W6BEG[10] Tile_X2Y2_LUT4AB/W6BEG[11]
+ Tile_X2Y2_LUT4AB/W6BEG[1] Tile_X2Y2_LUT4AB/W6BEG[2] Tile_X2Y2_LUT4AB/W6BEG[3] Tile_X2Y2_LUT4AB/W6BEG[4]
+ Tile_X2Y2_LUT4AB/W6BEG[5] Tile_X2Y2_LUT4AB/W6BEG[6] Tile_X2Y2_LUT4AB/W6BEG[7] Tile_X2Y2_LUT4AB/W6BEG[8]
+ Tile_X2Y2_LUT4AB/W6BEG[9] Tile_X3Y2_LUT4AB/W6BEG[0] Tile_X3Y2_LUT4AB/W6BEG[10] Tile_X3Y2_LUT4AB/W6BEG[11]
+ Tile_X3Y2_LUT4AB/W6BEG[1] Tile_X3Y2_LUT4AB/W6BEG[2] Tile_X3Y2_LUT4AB/W6BEG[3] Tile_X3Y2_LUT4AB/W6BEG[4]
+ Tile_X3Y2_LUT4AB/W6BEG[5] Tile_X3Y2_LUT4AB/W6BEG[6] Tile_X3Y2_LUT4AB/W6BEG[7] Tile_X3Y2_LUT4AB/W6BEG[8]
+ Tile_X3Y2_LUT4AB/W6BEG[9] Tile_X2Y2_LUT4AB/WW4BEG[0] Tile_X2Y2_LUT4AB/WW4BEG[10]
+ Tile_X2Y2_LUT4AB/WW4BEG[11] Tile_X2Y2_LUT4AB/WW4BEG[12] Tile_X2Y2_LUT4AB/WW4BEG[13]
+ Tile_X2Y2_LUT4AB/WW4BEG[14] Tile_X2Y2_LUT4AB/WW4BEG[15] Tile_X2Y2_LUT4AB/WW4BEG[1]
+ Tile_X2Y2_LUT4AB/WW4BEG[2] Tile_X2Y2_LUT4AB/WW4BEG[3] Tile_X2Y2_LUT4AB/WW4BEG[4]
+ Tile_X2Y2_LUT4AB/WW4BEG[5] Tile_X2Y2_LUT4AB/WW4BEG[6] Tile_X2Y2_LUT4AB/WW4BEG[7]
+ Tile_X2Y2_LUT4AB/WW4BEG[8] Tile_X2Y2_LUT4AB/WW4BEG[9] Tile_X3Y2_LUT4AB/WW4BEG[0]
+ Tile_X3Y2_LUT4AB/WW4BEG[10] Tile_X3Y2_LUT4AB/WW4BEG[11] Tile_X3Y2_LUT4AB/WW4BEG[12]
+ Tile_X3Y2_LUT4AB/WW4BEG[13] Tile_X3Y2_LUT4AB/WW4BEG[14] Tile_X3Y2_LUT4AB/WW4BEG[15]
+ Tile_X3Y2_LUT4AB/WW4BEG[1] Tile_X3Y2_LUT4AB/WW4BEG[2] Tile_X3Y2_LUT4AB/WW4BEG[3]
+ Tile_X3Y2_LUT4AB/WW4BEG[4] Tile_X3Y2_LUT4AB/WW4BEG[5] Tile_X3Y2_LUT4AB/WW4BEG[6]
+ Tile_X3Y2_LUT4AB/WW4BEG[7] Tile_X3Y2_LUT4AB/WW4BEG[8] Tile_X3Y2_LUT4AB/WW4BEG[9]
+ LUT4AB
XTile_X3Y9_S_IO4 Tile_X3Y9_A_I_top Tile_X3Y9_A_O_top Tile_X3Y9_A_T_top Tile_X3Y9_B_I_top
+ Tile_X3Y9_B_O_top Tile_X3Y9_B_T_top Tile_X3Y9_C_I_top Tile_X3Y9_C_O_top Tile_X3Y9_C_T_top
+ Tile_X3Y9_S_IO4/Co Tile_X3Y9_D_I_top Tile_X3Y9_D_O_top Tile_X3Y9_D_T_top Tile_X3Y9_S_IO4/FrameData[0]
+ Tile_X3Y9_S_IO4/FrameData[10] Tile_X3Y9_S_IO4/FrameData[11] Tile_X3Y9_S_IO4/FrameData[12]
+ Tile_X3Y9_S_IO4/FrameData[13] Tile_X3Y9_S_IO4/FrameData[14] Tile_X3Y9_S_IO4/FrameData[15]
+ Tile_X3Y9_S_IO4/FrameData[16] Tile_X3Y9_S_IO4/FrameData[17] Tile_X3Y9_S_IO4/FrameData[18]
+ Tile_X3Y9_S_IO4/FrameData[19] Tile_X3Y9_S_IO4/FrameData[1] Tile_X3Y9_S_IO4/FrameData[20]
+ Tile_X3Y9_S_IO4/FrameData[21] Tile_X3Y9_S_IO4/FrameData[22] Tile_X3Y9_S_IO4/FrameData[23]
+ Tile_X3Y9_S_IO4/FrameData[24] Tile_X3Y9_S_IO4/FrameData[25] Tile_X3Y9_S_IO4/FrameData[26]
+ Tile_X3Y9_S_IO4/FrameData[27] Tile_X3Y9_S_IO4/FrameData[28] Tile_X3Y9_S_IO4/FrameData[29]
+ Tile_X3Y9_S_IO4/FrameData[2] Tile_X3Y9_S_IO4/FrameData[30] Tile_X3Y9_S_IO4/FrameData[31]
+ Tile_X3Y9_S_IO4/FrameData[3] Tile_X3Y9_S_IO4/FrameData[4] Tile_X3Y9_S_IO4/FrameData[5]
+ Tile_X3Y9_S_IO4/FrameData[6] Tile_X3Y9_S_IO4/FrameData[7] Tile_X3Y9_S_IO4/FrameData[8]
+ Tile_X3Y9_S_IO4/FrameData[9] Tile_X4Y9_S_IO4/FrameData[0] Tile_X4Y9_S_IO4/FrameData[10]
+ Tile_X4Y9_S_IO4/FrameData[11] Tile_X4Y9_S_IO4/FrameData[12] Tile_X4Y9_S_IO4/FrameData[13]
+ Tile_X4Y9_S_IO4/FrameData[14] Tile_X4Y9_S_IO4/FrameData[15] Tile_X4Y9_S_IO4/FrameData[16]
+ Tile_X4Y9_S_IO4/FrameData[17] Tile_X4Y9_S_IO4/FrameData[18] Tile_X4Y9_S_IO4/FrameData[19]
+ Tile_X4Y9_S_IO4/FrameData[1] Tile_X4Y9_S_IO4/FrameData[20] Tile_X4Y9_S_IO4/FrameData[21]
+ Tile_X4Y9_S_IO4/FrameData[22] Tile_X4Y9_S_IO4/FrameData[23] Tile_X4Y9_S_IO4/FrameData[24]
+ Tile_X4Y9_S_IO4/FrameData[25] Tile_X4Y9_S_IO4/FrameData[26] Tile_X4Y9_S_IO4/FrameData[27]
+ Tile_X4Y9_S_IO4/FrameData[28] Tile_X4Y9_S_IO4/FrameData[29] Tile_X4Y9_S_IO4/FrameData[2]
+ Tile_X4Y9_S_IO4/FrameData[30] Tile_X4Y9_S_IO4/FrameData[31] Tile_X4Y9_S_IO4/FrameData[3]
+ Tile_X4Y9_S_IO4/FrameData[4] Tile_X4Y9_S_IO4/FrameData[5] Tile_X4Y9_S_IO4/FrameData[6]
+ Tile_X4Y9_S_IO4/FrameData[7] Tile_X4Y9_S_IO4/FrameData[8] Tile_X4Y9_S_IO4/FrameData[9]
+ FrameStrobe[60] FrameStrobe[70] FrameStrobe[71] FrameStrobe[72] FrameStrobe[73]
+ FrameStrobe[74] FrameStrobe[75] FrameStrobe[76] FrameStrobe[77] FrameStrobe[78]
+ FrameStrobe[79] FrameStrobe[61] FrameStrobe[62] FrameStrobe[63] FrameStrobe[64]
+ FrameStrobe[65] FrameStrobe[66] FrameStrobe[67] FrameStrobe[68] FrameStrobe[69]
+ Tile_X3Y8_LUT4AB/FrameStrobe[0] Tile_X3Y8_LUT4AB/FrameStrobe[10] Tile_X3Y8_LUT4AB/FrameStrobe[11]
+ Tile_X3Y8_LUT4AB/FrameStrobe[12] Tile_X3Y8_LUT4AB/FrameStrobe[13] Tile_X3Y8_LUT4AB/FrameStrobe[14]
+ Tile_X3Y8_LUT4AB/FrameStrobe[15] Tile_X3Y8_LUT4AB/FrameStrobe[16] Tile_X3Y8_LUT4AB/FrameStrobe[17]
+ Tile_X3Y8_LUT4AB/FrameStrobe[18] Tile_X3Y8_LUT4AB/FrameStrobe[19] Tile_X3Y8_LUT4AB/FrameStrobe[1]
+ Tile_X3Y8_LUT4AB/FrameStrobe[2] Tile_X3Y8_LUT4AB/FrameStrobe[3] Tile_X3Y8_LUT4AB/FrameStrobe[4]
+ Tile_X3Y8_LUT4AB/FrameStrobe[5] Tile_X3Y8_LUT4AB/FrameStrobe[6] Tile_X3Y8_LUT4AB/FrameStrobe[7]
+ Tile_X3Y8_LUT4AB/FrameStrobe[8] Tile_X3Y8_LUT4AB/FrameStrobe[9] Tile_X3Y9_S_IO4/N1BEG[0]
+ Tile_X3Y9_S_IO4/N1BEG[1] Tile_X3Y9_S_IO4/N1BEG[2] Tile_X3Y9_S_IO4/N1BEG[3] Tile_X3Y9_S_IO4/N2BEG[0]
+ Tile_X3Y9_S_IO4/N2BEG[1] Tile_X3Y9_S_IO4/N2BEG[2] Tile_X3Y9_S_IO4/N2BEG[3] Tile_X3Y9_S_IO4/N2BEG[4]
+ Tile_X3Y9_S_IO4/N2BEG[5] Tile_X3Y9_S_IO4/N2BEG[6] Tile_X3Y9_S_IO4/N2BEG[7] Tile_X3Y9_S_IO4/N2BEGb[0]
+ Tile_X3Y9_S_IO4/N2BEGb[1] Tile_X3Y9_S_IO4/N2BEGb[2] Tile_X3Y9_S_IO4/N2BEGb[3] Tile_X3Y9_S_IO4/N2BEGb[4]
+ Tile_X3Y9_S_IO4/N2BEGb[5] Tile_X3Y9_S_IO4/N2BEGb[6] Tile_X3Y9_S_IO4/N2BEGb[7] Tile_X3Y9_S_IO4/N4BEG[0]
+ Tile_X3Y9_S_IO4/N4BEG[10] Tile_X3Y9_S_IO4/N4BEG[11] Tile_X3Y9_S_IO4/N4BEG[12] Tile_X3Y9_S_IO4/N4BEG[13]
+ Tile_X3Y9_S_IO4/N4BEG[14] Tile_X3Y9_S_IO4/N4BEG[15] Tile_X3Y9_S_IO4/N4BEG[1] Tile_X3Y9_S_IO4/N4BEG[2]
+ Tile_X3Y9_S_IO4/N4BEG[3] Tile_X3Y9_S_IO4/N4BEG[4] Tile_X3Y9_S_IO4/N4BEG[5] Tile_X3Y9_S_IO4/N4BEG[6]
+ Tile_X3Y9_S_IO4/N4BEG[7] Tile_X3Y9_S_IO4/N4BEG[8] Tile_X3Y9_S_IO4/N4BEG[9] Tile_X3Y9_S_IO4/NN4BEG[0]
+ Tile_X3Y9_S_IO4/NN4BEG[10] Tile_X3Y9_S_IO4/NN4BEG[11] Tile_X3Y9_S_IO4/NN4BEG[12]
+ Tile_X3Y9_S_IO4/NN4BEG[13] Tile_X3Y9_S_IO4/NN4BEG[14] Tile_X3Y9_S_IO4/NN4BEG[15]
+ Tile_X3Y9_S_IO4/NN4BEG[1] Tile_X3Y9_S_IO4/NN4BEG[2] Tile_X3Y9_S_IO4/NN4BEG[3] Tile_X3Y9_S_IO4/NN4BEG[4]
+ Tile_X3Y9_S_IO4/NN4BEG[5] Tile_X3Y9_S_IO4/NN4BEG[6] Tile_X3Y9_S_IO4/NN4BEG[7] Tile_X3Y9_S_IO4/NN4BEG[8]
+ Tile_X3Y9_S_IO4/NN4BEG[9] Tile_X3Y9_S_IO4/S1END[0] Tile_X3Y9_S_IO4/S1END[1] Tile_X3Y9_S_IO4/S1END[2]
+ Tile_X3Y9_S_IO4/S1END[3] Tile_X3Y9_S_IO4/S2END[0] Tile_X3Y9_S_IO4/S2END[1] Tile_X3Y9_S_IO4/S2END[2]
+ Tile_X3Y9_S_IO4/S2END[3] Tile_X3Y9_S_IO4/S2END[4] Tile_X3Y9_S_IO4/S2END[5] Tile_X3Y9_S_IO4/S2END[6]
+ Tile_X3Y9_S_IO4/S2END[7] Tile_X3Y9_S_IO4/S2MID[0] Tile_X3Y9_S_IO4/S2MID[1] Tile_X3Y9_S_IO4/S2MID[2]
+ Tile_X3Y9_S_IO4/S2MID[3] Tile_X3Y9_S_IO4/S2MID[4] Tile_X3Y9_S_IO4/S2MID[5] Tile_X3Y9_S_IO4/S2MID[6]
+ Tile_X3Y9_S_IO4/S2MID[7] Tile_X3Y9_S_IO4/S4END[0] Tile_X3Y9_S_IO4/S4END[10] Tile_X3Y9_S_IO4/S4END[11]
+ Tile_X3Y9_S_IO4/S4END[12] Tile_X3Y9_S_IO4/S4END[13] Tile_X3Y9_S_IO4/S4END[14] Tile_X3Y9_S_IO4/S4END[15]
+ Tile_X3Y9_S_IO4/S4END[1] Tile_X3Y9_S_IO4/S4END[2] Tile_X3Y9_S_IO4/S4END[3] Tile_X3Y9_S_IO4/S4END[4]
+ Tile_X3Y9_S_IO4/S4END[5] Tile_X3Y9_S_IO4/S4END[6] Tile_X3Y9_S_IO4/S4END[7] Tile_X3Y9_S_IO4/S4END[8]
+ Tile_X3Y9_S_IO4/S4END[9] Tile_X3Y9_S_IO4/SS4END[0] Tile_X3Y9_S_IO4/SS4END[10] Tile_X3Y9_S_IO4/SS4END[11]
+ Tile_X3Y9_S_IO4/SS4END[12] Tile_X3Y9_S_IO4/SS4END[13] Tile_X3Y9_S_IO4/SS4END[14]
+ Tile_X3Y9_S_IO4/SS4END[15] Tile_X3Y9_S_IO4/SS4END[1] Tile_X3Y9_S_IO4/SS4END[2] Tile_X3Y9_S_IO4/SS4END[3]
+ Tile_X3Y9_S_IO4/SS4END[4] Tile_X3Y9_S_IO4/SS4END[5] Tile_X3Y9_S_IO4/SS4END[6] Tile_X3Y9_S_IO4/SS4END[7]
+ Tile_X3Y9_S_IO4/SS4END[8] Tile_X3Y9_S_IO4/SS4END[9] UserCLK Tile_X3Y9_S_IO4/UserCLKo
+ VGND VPWR S_IO4
XTile_X1Y6_LUT4AB Tile_X1Y7_LUT4AB/Co Tile_X1Y6_LUT4AB/Co Tile_X2Y6_LUT4AB/E1END[0]
+ Tile_X2Y6_LUT4AB/E1END[1] Tile_X2Y6_LUT4AB/E1END[2] Tile_X2Y6_LUT4AB/E1END[3] Tile_X1Y6_LUT4AB/E1END[0]
+ Tile_X1Y6_LUT4AB/E1END[1] Tile_X1Y6_LUT4AB/E1END[2] Tile_X1Y6_LUT4AB/E1END[3] Tile_X2Y6_LUT4AB/E2MID[0]
+ Tile_X2Y6_LUT4AB/E2MID[1] Tile_X2Y6_LUT4AB/E2MID[2] Tile_X2Y6_LUT4AB/E2MID[3] Tile_X2Y6_LUT4AB/E2MID[4]
+ Tile_X2Y6_LUT4AB/E2MID[5] Tile_X2Y6_LUT4AB/E2MID[6] Tile_X2Y6_LUT4AB/E2MID[7] Tile_X2Y6_LUT4AB/E2END[0]
+ Tile_X2Y6_LUT4AB/E2END[1] Tile_X2Y6_LUT4AB/E2END[2] Tile_X2Y6_LUT4AB/E2END[3] Tile_X2Y6_LUT4AB/E2END[4]
+ Tile_X2Y6_LUT4AB/E2END[5] Tile_X2Y6_LUT4AB/E2END[6] Tile_X2Y6_LUT4AB/E2END[7] Tile_X1Y6_LUT4AB/E2END[0]
+ Tile_X1Y6_LUT4AB/E2END[1] Tile_X1Y6_LUT4AB/E2END[2] Tile_X1Y6_LUT4AB/E2END[3] Tile_X1Y6_LUT4AB/E2END[4]
+ Tile_X1Y6_LUT4AB/E2END[5] Tile_X1Y6_LUT4AB/E2END[6] Tile_X1Y6_LUT4AB/E2END[7] Tile_X1Y6_LUT4AB/E2MID[0]
+ Tile_X1Y6_LUT4AB/E2MID[1] Tile_X1Y6_LUT4AB/E2MID[2] Tile_X1Y6_LUT4AB/E2MID[3] Tile_X1Y6_LUT4AB/E2MID[4]
+ Tile_X1Y6_LUT4AB/E2MID[5] Tile_X1Y6_LUT4AB/E2MID[6] Tile_X1Y6_LUT4AB/E2MID[7] Tile_X2Y6_LUT4AB/E6END[0]
+ Tile_X2Y6_LUT4AB/E6END[10] Tile_X2Y6_LUT4AB/E6END[11] Tile_X2Y6_LUT4AB/E6END[1]
+ Tile_X2Y6_LUT4AB/E6END[2] Tile_X2Y6_LUT4AB/E6END[3] Tile_X2Y6_LUT4AB/E6END[4] Tile_X2Y6_LUT4AB/E6END[5]
+ Tile_X2Y6_LUT4AB/E6END[6] Tile_X2Y6_LUT4AB/E6END[7] Tile_X2Y6_LUT4AB/E6END[8] Tile_X2Y6_LUT4AB/E6END[9]
+ Tile_X1Y6_LUT4AB/E6END[0] Tile_X1Y6_LUT4AB/E6END[10] Tile_X1Y6_LUT4AB/E6END[11]
+ Tile_X1Y6_LUT4AB/E6END[1] Tile_X1Y6_LUT4AB/E6END[2] Tile_X1Y6_LUT4AB/E6END[3] Tile_X1Y6_LUT4AB/E6END[4]
+ Tile_X1Y6_LUT4AB/E6END[5] Tile_X1Y6_LUT4AB/E6END[6] Tile_X1Y6_LUT4AB/E6END[7] Tile_X1Y6_LUT4AB/E6END[8]
+ Tile_X1Y6_LUT4AB/E6END[9] Tile_X2Y6_LUT4AB/EE4END[0] Tile_X2Y6_LUT4AB/EE4END[10]
+ Tile_X2Y6_LUT4AB/EE4END[11] Tile_X2Y6_LUT4AB/EE4END[12] Tile_X2Y6_LUT4AB/EE4END[13]
+ Tile_X2Y6_LUT4AB/EE4END[14] Tile_X2Y6_LUT4AB/EE4END[15] Tile_X2Y6_LUT4AB/EE4END[1]
+ Tile_X2Y6_LUT4AB/EE4END[2] Tile_X2Y6_LUT4AB/EE4END[3] Tile_X2Y6_LUT4AB/EE4END[4]
+ Tile_X2Y6_LUT4AB/EE4END[5] Tile_X2Y6_LUT4AB/EE4END[6] Tile_X2Y6_LUT4AB/EE4END[7]
+ Tile_X2Y6_LUT4AB/EE4END[8] Tile_X2Y6_LUT4AB/EE4END[9] Tile_X1Y6_LUT4AB/EE4END[0]
+ Tile_X1Y6_LUT4AB/EE4END[10] Tile_X1Y6_LUT4AB/EE4END[11] Tile_X1Y6_LUT4AB/EE4END[12]
+ Tile_X1Y6_LUT4AB/EE4END[13] Tile_X1Y6_LUT4AB/EE4END[14] Tile_X1Y6_LUT4AB/EE4END[15]
+ Tile_X1Y6_LUT4AB/EE4END[1] Tile_X1Y6_LUT4AB/EE4END[2] Tile_X1Y6_LUT4AB/EE4END[3]
+ Tile_X1Y6_LUT4AB/EE4END[4] Tile_X1Y6_LUT4AB/EE4END[5] Tile_X1Y6_LUT4AB/EE4END[6]
+ Tile_X1Y6_LUT4AB/EE4END[7] Tile_X1Y6_LUT4AB/EE4END[8] Tile_X1Y6_LUT4AB/EE4END[9]
+ Tile_X1Y6_LUT4AB/FrameData[0] Tile_X1Y6_LUT4AB/FrameData[10] Tile_X1Y6_LUT4AB/FrameData[11]
+ Tile_X1Y6_LUT4AB/FrameData[12] Tile_X1Y6_LUT4AB/FrameData[13] Tile_X1Y6_LUT4AB/FrameData[14]
+ Tile_X1Y6_LUT4AB/FrameData[15] Tile_X1Y6_LUT4AB/FrameData[16] Tile_X1Y6_LUT4AB/FrameData[17]
+ Tile_X1Y6_LUT4AB/FrameData[18] Tile_X1Y6_LUT4AB/FrameData[19] Tile_X1Y6_LUT4AB/FrameData[1]
+ Tile_X1Y6_LUT4AB/FrameData[20] Tile_X1Y6_LUT4AB/FrameData[21] Tile_X1Y6_LUT4AB/FrameData[22]
+ Tile_X1Y6_LUT4AB/FrameData[23] Tile_X1Y6_LUT4AB/FrameData[24] Tile_X1Y6_LUT4AB/FrameData[25]
+ Tile_X1Y6_LUT4AB/FrameData[26] Tile_X1Y6_LUT4AB/FrameData[27] Tile_X1Y6_LUT4AB/FrameData[28]
+ Tile_X1Y6_LUT4AB/FrameData[29] Tile_X1Y6_LUT4AB/FrameData[2] Tile_X1Y6_LUT4AB/FrameData[30]
+ Tile_X1Y6_LUT4AB/FrameData[31] Tile_X1Y6_LUT4AB/FrameData[3] Tile_X1Y6_LUT4AB/FrameData[4]
+ Tile_X1Y6_LUT4AB/FrameData[5] Tile_X1Y6_LUT4AB/FrameData[6] Tile_X1Y6_LUT4AB/FrameData[7]
+ Tile_X1Y6_LUT4AB/FrameData[8] Tile_X1Y6_LUT4AB/FrameData[9] Tile_X2Y6_LUT4AB/FrameData[0]
+ Tile_X2Y6_LUT4AB/FrameData[10] Tile_X2Y6_LUT4AB/FrameData[11] Tile_X2Y6_LUT4AB/FrameData[12]
+ Tile_X2Y6_LUT4AB/FrameData[13] Tile_X2Y6_LUT4AB/FrameData[14] Tile_X2Y6_LUT4AB/FrameData[15]
+ Tile_X2Y6_LUT4AB/FrameData[16] Tile_X2Y6_LUT4AB/FrameData[17] Tile_X2Y6_LUT4AB/FrameData[18]
+ Tile_X2Y6_LUT4AB/FrameData[19] Tile_X2Y6_LUT4AB/FrameData[1] Tile_X2Y6_LUT4AB/FrameData[20]
+ Tile_X2Y6_LUT4AB/FrameData[21] Tile_X2Y6_LUT4AB/FrameData[22] Tile_X2Y6_LUT4AB/FrameData[23]
+ Tile_X2Y6_LUT4AB/FrameData[24] Tile_X2Y6_LUT4AB/FrameData[25] Tile_X2Y6_LUT4AB/FrameData[26]
+ Tile_X2Y6_LUT4AB/FrameData[27] Tile_X2Y6_LUT4AB/FrameData[28] Tile_X2Y6_LUT4AB/FrameData[29]
+ Tile_X2Y6_LUT4AB/FrameData[2] Tile_X2Y6_LUT4AB/FrameData[30] Tile_X2Y6_LUT4AB/FrameData[31]
+ Tile_X2Y6_LUT4AB/FrameData[3] Tile_X2Y6_LUT4AB/FrameData[4] Tile_X2Y6_LUT4AB/FrameData[5]
+ Tile_X2Y6_LUT4AB/FrameData[6] Tile_X2Y6_LUT4AB/FrameData[7] Tile_X2Y6_LUT4AB/FrameData[8]
+ Tile_X2Y6_LUT4AB/FrameData[9] Tile_X1Y6_LUT4AB/FrameStrobe[0] Tile_X1Y6_LUT4AB/FrameStrobe[10]
+ Tile_X1Y6_LUT4AB/FrameStrobe[11] Tile_X1Y6_LUT4AB/FrameStrobe[12] Tile_X1Y6_LUT4AB/FrameStrobe[13]
+ Tile_X1Y6_LUT4AB/FrameStrobe[14] Tile_X1Y6_LUT4AB/FrameStrobe[15] Tile_X1Y6_LUT4AB/FrameStrobe[16]
+ Tile_X1Y6_LUT4AB/FrameStrobe[17] Tile_X1Y6_LUT4AB/FrameStrobe[18] Tile_X1Y6_LUT4AB/FrameStrobe[19]
+ Tile_X1Y6_LUT4AB/FrameStrobe[1] Tile_X1Y6_LUT4AB/FrameStrobe[2] Tile_X1Y6_LUT4AB/FrameStrobe[3]
+ Tile_X1Y6_LUT4AB/FrameStrobe[4] Tile_X1Y6_LUT4AB/FrameStrobe[5] Tile_X1Y6_LUT4AB/FrameStrobe[6]
+ Tile_X1Y6_LUT4AB/FrameStrobe[7] Tile_X1Y6_LUT4AB/FrameStrobe[8] Tile_X1Y6_LUT4AB/FrameStrobe[9]
+ Tile_X1Y5_LUT4AB/FrameStrobe[0] Tile_X1Y5_LUT4AB/FrameStrobe[10] Tile_X1Y5_LUT4AB/FrameStrobe[11]
+ Tile_X1Y5_LUT4AB/FrameStrobe[12] Tile_X1Y5_LUT4AB/FrameStrobe[13] Tile_X1Y5_LUT4AB/FrameStrobe[14]
+ Tile_X1Y5_LUT4AB/FrameStrobe[15] Tile_X1Y5_LUT4AB/FrameStrobe[16] Tile_X1Y5_LUT4AB/FrameStrobe[17]
+ Tile_X1Y5_LUT4AB/FrameStrobe[18] Tile_X1Y5_LUT4AB/FrameStrobe[19] Tile_X1Y5_LUT4AB/FrameStrobe[1]
+ Tile_X1Y5_LUT4AB/FrameStrobe[2] Tile_X1Y5_LUT4AB/FrameStrobe[3] Tile_X1Y5_LUT4AB/FrameStrobe[4]
+ Tile_X1Y5_LUT4AB/FrameStrobe[5] Tile_X1Y5_LUT4AB/FrameStrobe[6] Tile_X1Y5_LUT4AB/FrameStrobe[7]
+ Tile_X1Y5_LUT4AB/FrameStrobe[8] Tile_X1Y5_LUT4AB/FrameStrobe[9] Tile_X1Y6_LUT4AB/N1BEG[0]
+ Tile_X1Y6_LUT4AB/N1BEG[1] Tile_X1Y6_LUT4AB/N1BEG[2] Tile_X1Y6_LUT4AB/N1BEG[3] Tile_X1Y7_LUT4AB/N1BEG[0]
+ Tile_X1Y7_LUT4AB/N1BEG[1] Tile_X1Y7_LUT4AB/N1BEG[2] Tile_X1Y7_LUT4AB/N1BEG[3] Tile_X1Y6_LUT4AB/N2BEG[0]
+ Tile_X1Y6_LUT4AB/N2BEG[1] Tile_X1Y6_LUT4AB/N2BEG[2] Tile_X1Y6_LUT4AB/N2BEG[3] Tile_X1Y6_LUT4AB/N2BEG[4]
+ Tile_X1Y6_LUT4AB/N2BEG[5] Tile_X1Y6_LUT4AB/N2BEG[6] Tile_X1Y6_LUT4AB/N2BEG[7] Tile_X1Y5_LUT4AB/N2END[0]
+ Tile_X1Y5_LUT4AB/N2END[1] Tile_X1Y5_LUT4AB/N2END[2] Tile_X1Y5_LUT4AB/N2END[3] Tile_X1Y5_LUT4AB/N2END[4]
+ Tile_X1Y5_LUT4AB/N2END[5] Tile_X1Y5_LUT4AB/N2END[6] Tile_X1Y5_LUT4AB/N2END[7] Tile_X1Y6_LUT4AB/N2END[0]
+ Tile_X1Y6_LUT4AB/N2END[1] Tile_X1Y6_LUT4AB/N2END[2] Tile_X1Y6_LUT4AB/N2END[3] Tile_X1Y6_LUT4AB/N2END[4]
+ Tile_X1Y6_LUT4AB/N2END[5] Tile_X1Y6_LUT4AB/N2END[6] Tile_X1Y6_LUT4AB/N2END[7] Tile_X1Y7_LUT4AB/N2BEG[0]
+ Tile_X1Y7_LUT4AB/N2BEG[1] Tile_X1Y7_LUT4AB/N2BEG[2] Tile_X1Y7_LUT4AB/N2BEG[3] Tile_X1Y7_LUT4AB/N2BEG[4]
+ Tile_X1Y7_LUT4AB/N2BEG[5] Tile_X1Y7_LUT4AB/N2BEG[6] Tile_X1Y7_LUT4AB/N2BEG[7] Tile_X1Y6_LUT4AB/N4BEG[0]
+ Tile_X1Y6_LUT4AB/N4BEG[10] Tile_X1Y6_LUT4AB/N4BEG[11] Tile_X1Y6_LUT4AB/N4BEG[12]
+ Tile_X1Y6_LUT4AB/N4BEG[13] Tile_X1Y6_LUT4AB/N4BEG[14] Tile_X1Y6_LUT4AB/N4BEG[15]
+ Tile_X1Y6_LUT4AB/N4BEG[1] Tile_X1Y6_LUT4AB/N4BEG[2] Tile_X1Y6_LUT4AB/N4BEG[3] Tile_X1Y6_LUT4AB/N4BEG[4]
+ Tile_X1Y6_LUT4AB/N4BEG[5] Tile_X1Y6_LUT4AB/N4BEG[6] Tile_X1Y6_LUT4AB/N4BEG[7] Tile_X1Y6_LUT4AB/N4BEG[8]
+ Tile_X1Y6_LUT4AB/N4BEG[9] Tile_X1Y7_LUT4AB/N4BEG[0] Tile_X1Y7_LUT4AB/N4BEG[10] Tile_X1Y7_LUT4AB/N4BEG[11]
+ Tile_X1Y7_LUT4AB/N4BEG[12] Tile_X1Y7_LUT4AB/N4BEG[13] Tile_X1Y7_LUT4AB/N4BEG[14]
+ Tile_X1Y7_LUT4AB/N4BEG[15] Tile_X1Y7_LUT4AB/N4BEG[1] Tile_X1Y7_LUT4AB/N4BEG[2] Tile_X1Y7_LUT4AB/N4BEG[3]
+ Tile_X1Y7_LUT4AB/N4BEG[4] Tile_X1Y7_LUT4AB/N4BEG[5] Tile_X1Y7_LUT4AB/N4BEG[6] Tile_X1Y7_LUT4AB/N4BEG[7]
+ Tile_X1Y7_LUT4AB/N4BEG[8] Tile_X1Y7_LUT4AB/N4BEG[9] Tile_X1Y6_LUT4AB/NN4BEG[0] Tile_X1Y6_LUT4AB/NN4BEG[10]
+ Tile_X1Y6_LUT4AB/NN4BEG[11] Tile_X1Y6_LUT4AB/NN4BEG[12] Tile_X1Y6_LUT4AB/NN4BEG[13]
+ Tile_X1Y6_LUT4AB/NN4BEG[14] Tile_X1Y6_LUT4AB/NN4BEG[15] Tile_X1Y6_LUT4AB/NN4BEG[1]
+ Tile_X1Y6_LUT4AB/NN4BEG[2] Tile_X1Y6_LUT4AB/NN4BEG[3] Tile_X1Y6_LUT4AB/NN4BEG[4]
+ Tile_X1Y6_LUT4AB/NN4BEG[5] Tile_X1Y6_LUT4AB/NN4BEG[6] Tile_X1Y6_LUT4AB/NN4BEG[7]
+ Tile_X1Y6_LUT4AB/NN4BEG[8] Tile_X1Y6_LUT4AB/NN4BEG[9] Tile_X1Y7_LUT4AB/NN4BEG[0]
+ Tile_X1Y7_LUT4AB/NN4BEG[10] Tile_X1Y7_LUT4AB/NN4BEG[11] Tile_X1Y7_LUT4AB/NN4BEG[12]
+ Tile_X1Y7_LUT4AB/NN4BEG[13] Tile_X1Y7_LUT4AB/NN4BEG[14] Tile_X1Y7_LUT4AB/NN4BEG[15]
+ Tile_X1Y7_LUT4AB/NN4BEG[1] Tile_X1Y7_LUT4AB/NN4BEG[2] Tile_X1Y7_LUT4AB/NN4BEG[3]
+ Tile_X1Y7_LUT4AB/NN4BEG[4] Tile_X1Y7_LUT4AB/NN4BEG[5] Tile_X1Y7_LUT4AB/NN4BEG[6]
+ Tile_X1Y7_LUT4AB/NN4BEG[7] Tile_X1Y7_LUT4AB/NN4BEG[8] Tile_X1Y7_LUT4AB/NN4BEG[9]
+ Tile_X1Y7_LUT4AB/S1END[0] Tile_X1Y7_LUT4AB/S1END[1] Tile_X1Y7_LUT4AB/S1END[2] Tile_X1Y7_LUT4AB/S1END[3]
+ Tile_X1Y6_LUT4AB/S1END[0] Tile_X1Y6_LUT4AB/S1END[1] Tile_X1Y6_LUT4AB/S1END[2] Tile_X1Y6_LUT4AB/S1END[3]
+ Tile_X1Y7_LUT4AB/S2MID[0] Tile_X1Y7_LUT4AB/S2MID[1] Tile_X1Y7_LUT4AB/S2MID[2] Tile_X1Y7_LUT4AB/S2MID[3]
+ Tile_X1Y7_LUT4AB/S2MID[4] Tile_X1Y7_LUT4AB/S2MID[5] Tile_X1Y7_LUT4AB/S2MID[6] Tile_X1Y7_LUT4AB/S2MID[7]
+ Tile_X1Y7_LUT4AB/S2END[0] Tile_X1Y7_LUT4AB/S2END[1] Tile_X1Y7_LUT4AB/S2END[2] Tile_X1Y7_LUT4AB/S2END[3]
+ Tile_X1Y7_LUT4AB/S2END[4] Tile_X1Y7_LUT4AB/S2END[5] Tile_X1Y7_LUT4AB/S2END[6] Tile_X1Y7_LUT4AB/S2END[7]
+ Tile_X1Y6_LUT4AB/S2END[0] Tile_X1Y6_LUT4AB/S2END[1] Tile_X1Y6_LUT4AB/S2END[2] Tile_X1Y6_LUT4AB/S2END[3]
+ Tile_X1Y6_LUT4AB/S2END[4] Tile_X1Y6_LUT4AB/S2END[5] Tile_X1Y6_LUT4AB/S2END[6] Tile_X1Y6_LUT4AB/S2END[7]
+ Tile_X1Y6_LUT4AB/S2MID[0] Tile_X1Y6_LUT4AB/S2MID[1] Tile_X1Y6_LUT4AB/S2MID[2] Tile_X1Y6_LUT4AB/S2MID[3]
+ Tile_X1Y6_LUT4AB/S2MID[4] Tile_X1Y6_LUT4AB/S2MID[5] Tile_X1Y6_LUT4AB/S2MID[6] Tile_X1Y6_LUT4AB/S2MID[7]
+ Tile_X1Y7_LUT4AB/S4END[0] Tile_X1Y7_LUT4AB/S4END[10] Tile_X1Y7_LUT4AB/S4END[11]
+ Tile_X1Y7_LUT4AB/S4END[12] Tile_X1Y7_LUT4AB/S4END[13] Tile_X1Y7_LUT4AB/S4END[14]
+ Tile_X1Y7_LUT4AB/S4END[15] Tile_X1Y7_LUT4AB/S4END[1] Tile_X1Y7_LUT4AB/S4END[2] Tile_X1Y7_LUT4AB/S4END[3]
+ Tile_X1Y7_LUT4AB/S4END[4] Tile_X1Y7_LUT4AB/S4END[5] Tile_X1Y7_LUT4AB/S4END[6] Tile_X1Y7_LUT4AB/S4END[7]
+ Tile_X1Y7_LUT4AB/S4END[8] Tile_X1Y7_LUT4AB/S4END[9] Tile_X1Y6_LUT4AB/S4END[0] Tile_X1Y6_LUT4AB/S4END[10]
+ Tile_X1Y6_LUT4AB/S4END[11] Tile_X1Y6_LUT4AB/S4END[12] Tile_X1Y6_LUT4AB/S4END[13]
+ Tile_X1Y6_LUT4AB/S4END[14] Tile_X1Y6_LUT4AB/S4END[15] Tile_X1Y6_LUT4AB/S4END[1]
+ Tile_X1Y6_LUT4AB/S4END[2] Tile_X1Y6_LUT4AB/S4END[3] Tile_X1Y6_LUT4AB/S4END[4] Tile_X1Y6_LUT4AB/S4END[5]
+ Tile_X1Y6_LUT4AB/S4END[6] Tile_X1Y6_LUT4AB/S4END[7] Tile_X1Y6_LUT4AB/S4END[8] Tile_X1Y6_LUT4AB/S4END[9]
+ Tile_X1Y7_LUT4AB/SS4END[0] Tile_X1Y7_LUT4AB/SS4END[10] Tile_X1Y7_LUT4AB/SS4END[11]
+ Tile_X1Y7_LUT4AB/SS4END[12] Tile_X1Y7_LUT4AB/SS4END[13] Tile_X1Y7_LUT4AB/SS4END[14]
+ Tile_X1Y7_LUT4AB/SS4END[15] Tile_X1Y7_LUT4AB/SS4END[1] Tile_X1Y7_LUT4AB/SS4END[2]
+ Tile_X1Y7_LUT4AB/SS4END[3] Tile_X1Y7_LUT4AB/SS4END[4] Tile_X1Y7_LUT4AB/SS4END[5]
+ Tile_X1Y7_LUT4AB/SS4END[6] Tile_X1Y7_LUT4AB/SS4END[7] Tile_X1Y7_LUT4AB/SS4END[8]
+ Tile_X1Y7_LUT4AB/SS4END[9] Tile_X1Y6_LUT4AB/SS4END[0] Tile_X1Y6_LUT4AB/SS4END[10]
+ Tile_X1Y6_LUT4AB/SS4END[11] Tile_X1Y6_LUT4AB/SS4END[12] Tile_X1Y6_LUT4AB/SS4END[13]
+ Tile_X1Y6_LUT4AB/SS4END[14] Tile_X1Y6_LUT4AB/SS4END[15] Tile_X1Y6_LUT4AB/SS4END[1]
+ Tile_X1Y6_LUT4AB/SS4END[2] Tile_X1Y6_LUT4AB/SS4END[3] Tile_X1Y6_LUT4AB/SS4END[4]
+ Tile_X1Y6_LUT4AB/SS4END[5] Tile_X1Y6_LUT4AB/SS4END[6] Tile_X1Y6_LUT4AB/SS4END[7]
+ Tile_X1Y6_LUT4AB/SS4END[8] Tile_X1Y6_LUT4AB/SS4END[9] Tile_X1Y6_LUT4AB/UserCLK Tile_X1Y5_LUT4AB/UserCLK
+ VGND VPWR Tile_X1Y6_LUT4AB/W1BEG[0] Tile_X1Y6_LUT4AB/W1BEG[1] Tile_X1Y6_LUT4AB/W1BEG[2]
+ Tile_X1Y6_LUT4AB/W1BEG[3] Tile_X2Y6_LUT4AB/W1BEG[0] Tile_X2Y6_LUT4AB/W1BEG[1] Tile_X2Y6_LUT4AB/W1BEG[2]
+ Tile_X2Y6_LUT4AB/W1BEG[3] Tile_X1Y6_LUT4AB/W2BEG[0] Tile_X1Y6_LUT4AB/W2BEG[1] Tile_X1Y6_LUT4AB/W2BEG[2]
+ Tile_X1Y6_LUT4AB/W2BEG[3] Tile_X1Y6_LUT4AB/W2BEG[4] Tile_X1Y6_LUT4AB/W2BEG[5] Tile_X1Y6_LUT4AB/W2BEG[6]
+ Tile_X1Y6_LUT4AB/W2BEG[7] Tile_X1Y6_LUT4AB/W2BEGb[0] Tile_X1Y6_LUT4AB/W2BEGb[1]
+ Tile_X1Y6_LUT4AB/W2BEGb[2] Tile_X1Y6_LUT4AB/W2BEGb[3] Tile_X1Y6_LUT4AB/W2BEGb[4]
+ Tile_X1Y6_LUT4AB/W2BEGb[5] Tile_X1Y6_LUT4AB/W2BEGb[6] Tile_X1Y6_LUT4AB/W2BEGb[7]
+ Tile_X1Y6_LUT4AB/W2END[0] Tile_X1Y6_LUT4AB/W2END[1] Tile_X1Y6_LUT4AB/W2END[2] Tile_X1Y6_LUT4AB/W2END[3]
+ Tile_X1Y6_LUT4AB/W2END[4] Tile_X1Y6_LUT4AB/W2END[5] Tile_X1Y6_LUT4AB/W2END[6] Tile_X1Y6_LUT4AB/W2END[7]
+ Tile_X2Y6_LUT4AB/W2BEG[0] Tile_X2Y6_LUT4AB/W2BEG[1] Tile_X2Y6_LUT4AB/W2BEG[2] Tile_X2Y6_LUT4AB/W2BEG[3]
+ Tile_X2Y6_LUT4AB/W2BEG[4] Tile_X2Y6_LUT4AB/W2BEG[5] Tile_X2Y6_LUT4AB/W2BEG[6] Tile_X2Y6_LUT4AB/W2BEG[7]
+ Tile_X1Y6_LUT4AB/W6BEG[0] Tile_X1Y6_LUT4AB/W6BEG[10] Tile_X1Y6_LUT4AB/W6BEG[11]
+ Tile_X1Y6_LUT4AB/W6BEG[1] Tile_X1Y6_LUT4AB/W6BEG[2] Tile_X1Y6_LUT4AB/W6BEG[3] Tile_X1Y6_LUT4AB/W6BEG[4]
+ Tile_X1Y6_LUT4AB/W6BEG[5] Tile_X1Y6_LUT4AB/W6BEG[6] Tile_X1Y6_LUT4AB/W6BEG[7] Tile_X1Y6_LUT4AB/W6BEG[8]
+ Tile_X1Y6_LUT4AB/W6BEG[9] Tile_X2Y6_LUT4AB/W6BEG[0] Tile_X2Y6_LUT4AB/W6BEG[10] Tile_X2Y6_LUT4AB/W6BEG[11]
+ Tile_X2Y6_LUT4AB/W6BEG[1] Tile_X2Y6_LUT4AB/W6BEG[2] Tile_X2Y6_LUT4AB/W6BEG[3] Tile_X2Y6_LUT4AB/W6BEG[4]
+ Tile_X2Y6_LUT4AB/W6BEG[5] Tile_X2Y6_LUT4AB/W6BEG[6] Tile_X2Y6_LUT4AB/W6BEG[7] Tile_X2Y6_LUT4AB/W6BEG[8]
+ Tile_X2Y6_LUT4AB/W6BEG[9] Tile_X1Y6_LUT4AB/WW4BEG[0] Tile_X1Y6_LUT4AB/WW4BEG[10]
+ Tile_X1Y6_LUT4AB/WW4BEG[11] Tile_X1Y6_LUT4AB/WW4BEG[12] Tile_X1Y6_LUT4AB/WW4BEG[13]
+ Tile_X1Y6_LUT4AB/WW4BEG[14] Tile_X1Y6_LUT4AB/WW4BEG[15] Tile_X1Y6_LUT4AB/WW4BEG[1]
+ Tile_X1Y6_LUT4AB/WW4BEG[2] Tile_X1Y6_LUT4AB/WW4BEG[3] Tile_X1Y6_LUT4AB/WW4BEG[4]
+ Tile_X1Y6_LUT4AB/WW4BEG[5] Tile_X1Y6_LUT4AB/WW4BEG[6] Tile_X1Y6_LUT4AB/WW4BEG[7]
+ Tile_X1Y6_LUT4AB/WW4BEG[8] Tile_X1Y6_LUT4AB/WW4BEG[9] Tile_X2Y6_LUT4AB/WW4BEG[0]
+ Tile_X2Y6_LUT4AB/WW4BEG[10] Tile_X2Y6_LUT4AB/WW4BEG[11] Tile_X2Y6_LUT4AB/WW4BEG[12]
+ Tile_X2Y6_LUT4AB/WW4BEG[13] Tile_X2Y6_LUT4AB/WW4BEG[14] Tile_X2Y6_LUT4AB/WW4BEG[15]
+ Tile_X2Y6_LUT4AB/WW4BEG[1] Tile_X2Y6_LUT4AB/WW4BEG[2] Tile_X2Y6_LUT4AB/WW4BEG[3]
+ Tile_X2Y6_LUT4AB/WW4BEG[4] Tile_X2Y6_LUT4AB/WW4BEG[5] Tile_X2Y6_LUT4AB/WW4BEG[6]
+ Tile_X2Y6_LUT4AB/WW4BEG[7] Tile_X2Y6_LUT4AB/WW4BEG[8] Tile_X2Y6_LUT4AB/WW4BEG[9]
+ LUT4AB
XTile_X3Y4_LUT4AB Tile_X3Y5_LUT4AB/Co Tile_X3Y4_LUT4AB/Co Tile_X4Y4_LUT4AB/E1END[0]
+ Tile_X4Y4_LUT4AB/E1END[1] Tile_X4Y4_LUT4AB/E1END[2] Tile_X4Y4_LUT4AB/E1END[3] Tile_X3Y4_LUT4AB/E1END[0]
+ Tile_X3Y4_LUT4AB/E1END[1] Tile_X3Y4_LUT4AB/E1END[2] Tile_X3Y4_LUT4AB/E1END[3] Tile_X4Y4_LUT4AB/E2MID[0]
+ Tile_X4Y4_LUT4AB/E2MID[1] Tile_X4Y4_LUT4AB/E2MID[2] Tile_X4Y4_LUT4AB/E2MID[3] Tile_X4Y4_LUT4AB/E2MID[4]
+ Tile_X4Y4_LUT4AB/E2MID[5] Tile_X4Y4_LUT4AB/E2MID[6] Tile_X4Y4_LUT4AB/E2MID[7] Tile_X4Y4_LUT4AB/E2END[0]
+ Tile_X4Y4_LUT4AB/E2END[1] Tile_X4Y4_LUT4AB/E2END[2] Tile_X4Y4_LUT4AB/E2END[3] Tile_X4Y4_LUT4AB/E2END[4]
+ Tile_X4Y4_LUT4AB/E2END[5] Tile_X4Y4_LUT4AB/E2END[6] Tile_X4Y4_LUT4AB/E2END[7] Tile_X3Y4_LUT4AB/E2END[0]
+ Tile_X3Y4_LUT4AB/E2END[1] Tile_X3Y4_LUT4AB/E2END[2] Tile_X3Y4_LUT4AB/E2END[3] Tile_X3Y4_LUT4AB/E2END[4]
+ Tile_X3Y4_LUT4AB/E2END[5] Tile_X3Y4_LUT4AB/E2END[6] Tile_X3Y4_LUT4AB/E2END[7] Tile_X3Y4_LUT4AB/E2MID[0]
+ Tile_X3Y4_LUT4AB/E2MID[1] Tile_X3Y4_LUT4AB/E2MID[2] Tile_X3Y4_LUT4AB/E2MID[3] Tile_X3Y4_LUT4AB/E2MID[4]
+ Tile_X3Y4_LUT4AB/E2MID[5] Tile_X3Y4_LUT4AB/E2MID[6] Tile_X3Y4_LUT4AB/E2MID[7] Tile_X4Y4_LUT4AB/E6END[0]
+ Tile_X4Y4_LUT4AB/E6END[10] Tile_X4Y4_LUT4AB/E6END[11] Tile_X4Y4_LUT4AB/E6END[1]
+ Tile_X4Y4_LUT4AB/E6END[2] Tile_X4Y4_LUT4AB/E6END[3] Tile_X4Y4_LUT4AB/E6END[4] Tile_X4Y4_LUT4AB/E6END[5]
+ Tile_X4Y4_LUT4AB/E6END[6] Tile_X4Y4_LUT4AB/E6END[7] Tile_X4Y4_LUT4AB/E6END[8] Tile_X4Y4_LUT4AB/E6END[9]
+ Tile_X3Y4_LUT4AB/E6END[0] Tile_X3Y4_LUT4AB/E6END[10] Tile_X3Y4_LUT4AB/E6END[11]
+ Tile_X3Y4_LUT4AB/E6END[1] Tile_X3Y4_LUT4AB/E6END[2] Tile_X3Y4_LUT4AB/E6END[3] Tile_X3Y4_LUT4AB/E6END[4]
+ Tile_X3Y4_LUT4AB/E6END[5] Tile_X3Y4_LUT4AB/E6END[6] Tile_X3Y4_LUT4AB/E6END[7] Tile_X3Y4_LUT4AB/E6END[8]
+ Tile_X3Y4_LUT4AB/E6END[9] Tile_X4Y4_LUT4AB/EE4END[0] Tile_X4Y4_LUT4AB/EE4END[10]
+ Tile_X4Y4_LUT4AB/EE4END[11] Tile_X4Y4_LUT4AB/EE4END[12] Tile_X4Y4_LUT4AB/EE4END[13]
+ Tile_X4Y4_LUT4AB/EE4END[14] Tile_X4Y4_LUT4AB/EE4END[15] Tile_X4Y4_LUT4AB/EE4END[1]
+ Tile_X4Y4_LUT4AB/EE4END[2] Tile_X4Y4_LUT4AB/EE4END[3] Tile_X4Y4_LUT4AB/EE4END[4]
+ Tile_X4Y4_LUT4AB/EE4END[5] Tile_X4Y4_LUT4AB/EE4END[6] Tile_X4Y4_LUT4AB/EE4END[7]
+ Tile_X4Y4_LUT4AB/EE4END[8] Tile_X4Y4_LUT4AB/EE4END[9] Tile_X3Y4_LUT4AB/EE4END[0]
+ Tile_X3Y4_LUT4AB/EE4END[10] Tile_X3Y4_LUT4AB/EE4END[11] Tile_X3Y4_LUT4AB/EE4END[12]
+ Tile_X3Y4_LUT4AB/EE4END[13] Tile_X3Y4_LUT4AB/EE4END[14] Tile_X3Y4_LUT4AB/EE4END[15]
+ Tile_X3Y4_LUT4AB/EE4END[1] Tile_X3Y4_LUT4AB/EE4END[2] Tile_X3Y4_LUT4AB/EE4END[3]
+ Tile_X3Y4_LUT4AB/EE4END[4] Tile_X3Y4_LUT4AB/EE4END[5] Tile_X3Y4_LUT4AB/EE4END[6]
+ Tile_X3Y4_LUT4AB/EE4END[7] Tile_X3Y4_LUT4AB/EE4END[8] Tile_X3Y4_LUT4AB/EE4END[9]
+ Tile_X3Y4_LUT4AB/FrameData[0] Tile_X3Y4_LUT4AB/FrameData[10] Tile_X3Y4_LUT4AB/FrameData[11]
+ Tile_X3Y4_LUT4AB/FrameData[12] Tile_X3Y4_LUT4AB/FrameData[13] Tile_X3Y4_LUT4AB/FrameData[14]
+ Tile_X3Y4_LUT4AB/FrameData[15] Tile_X3Y4_LUT4AB/FrameData[16] Tile_X3Y4_LUT4AB/FrameData[17]
+ Tile_X3Y4_LUT4AB/FrameData[18] Tile_X3Y4_LUT4AB/FrameData[19] Tile_X3Y4_LUT4AB/FrameData[1]
+ Tile_X3Y4_LUT4AB/FrameData[20] Tile_X3Y4_LUT4AB/FrameData[21] Tile_X3Y4_LUT4AB/FrameData[22]
+ Tile_X3Y4_LUT4AB/FrameData[23] Tile_X3Y4_LUT4AB/FrameData[24] Tile_X3Y4_LUT4AB/FrameData[25]
+ Tile_X3Y4_LUT4AB/FrameData[26] Tile_X3Y4_LUT4AB/FrameData[27] Tile_X3Y4_LUT4AB/FrameData[28]
+ Tile_X3Y4_LUT4AB/FrameData[29] Tile_X3Y4_LUT4AB/FrameData[2] Tile_X3Y4_LUT4AB/FrameData[30]
+ Tile_X3Y4_LUT4AB/FrameData[31] Tile_X3Y4_LUT4AB/FrameData[3] Tile_X3Y4_LUT4AB/FrameData[4]
+ Tile_X3Y4_LUT4AB/FrameData[5] Tile_X3Y4_LUT4AB/FrameData[6] Tile_X3Y4_LUT4AB/FrameData[7]
+ Tile_X3Y4_LUT4AB/FrameData[8] Tile_X3Y4_LUT4AB/FrameData[9] Tile_X4Y4_LUT4AB/FrameData[0]
+ Tile_X4Y4_LUT4AB/FrameData[10] Tile_X4Y4_LUT4AB/FrameData[11] Tile_X4Y4_LUT4AB/FrameData[12]
+ Tile_X4Y4_LUT4AB/FrameData[13] Tile_X4Y4_LUT4AB/FrameData[14] Tile_X4Y4_LUT4AB/FrameData[15]
+ Tile_X4Y4_LUT4AB/FrameData[16] Tile_X4Y4_LUT4AB/FrameData[17] Tile_X4Y4_LUT4AB/FrameData[18]
+ Tile_X4Y4_LUT4AB/FrameData[19] Tile_X4Y4_LUT4AB/FrameData[1] Tile_X4Y4_LUT4AB/FrameData[20]
+ Tile_X4Y4_LUT4AB/FrameData[21] Tile_X4Y4_LUT4AB/FrameData[22] Tile_X4Y4_LUT4AB/FrameData[23]
+ Tile_X4Y4_LUT4AB/FrameData[24] Tile_X4Y4_LUT4AB/FrameData[25] Tile_X4Y4_LUT4AB/FrameData[26]
+ Tile_X4Y4_LUT4AB/FrameData[27] Tile_X4Y4_LUT4AB/FrameData[28] Tile_X4Y4_LUT4AB/FrameData[29]
+ Tile_X4Y4_LUT4AB/FrameData[2] Tile_X4Y4_LUT4AB/FrameData[30] Tile_X4Y4_LUT4AB/FrameData[31]
+ Tile_X4Y4_LUT4AB/FrameData[3] Tile_X4Y4_LUT4AB/FrameData[4] Tile_X4Y4_LUT4AB/FrameData[5]
+ Tile_X4Y4_LUT4AB/FrameData[6] Tile_X4Y4_LUT4AB/FrameData[7] Tile_X4Y4_LUT4AB/FrameData[8]
+ Tile_X4Y4_LUT4AB/FrameData[9] Tile_X3Y4_LUT4AB/FrameStrobe[0] Tile_X3Y4_LUT4AB/FrameStrobe[10]
+ Tile_X3Y4_LUT4AB/FrameStrobe[11] Tile_X3Y4_LUT4AB/FrameStrobe[12] Tile_X3Y4_LUT4AB/FrameStrobe[13]
+ Tile_X3Y4_LUT4AB/FrameStrobe[14] Tile_X3Y4_LUT4AB/FrameStrobe[15] Tile_X3Y4_LUT4AB/FrameStrobe[16]
+ Tile_X3Y4_LUT4AB/FrameStrobe[17] Tile_X3Y4_LUT4AB/FrameStrobe[18] Tile_X3Y4_LUT4AB/FrameStrobe[19]
+ Tile_X3Y4_LUT4AB/FrameStrobe[1] Tile_X3Y4_LUT4AB/FrameStrobe[2] Tile_X3Y4_LUT4AB/FrameStrobe[3]
+ Tile_X3Y4_LUT4AB/FrameStrobe[4] Tile_X3Y4_LUT4AB/FrameStrobe[5] Tile_X3Y4_LUT4AB/FrameStrobe[6]
+ Tile_X3Y4_LUT4AB/FrameStrobe[7] Tile_X3Y4_LUT4AB/FrameStrobe[8] Tile_X3Y4_LUT4AB/FrameStrobe[9]
+ Tile_X3Y3_LUT4AB/FrameStrobe[0] Tile_X3Y3_LUT4AB/FrameStrobe[10] Tile_X3Y3_LUT4AB/FrameStrobe[11]
+ Tile_X3Y3_LUT4AB/FrameStrobe[12] Tile_X3Y3_LUT4AB/FrameStrobe[13] Tile_X3Y3_LUT4AB/FrameStrobe[14]
+ Tile_X3Y3_LUT4AB/FrameStrobe[15] Tile_X3Y3_LUT4AB/FrameStrobe[16] Tile_X3Y3_LUT4AB/FrameStrobe[17]
+ Tile_X3Y3_LUT4AB/FrameStrobe[18] Tile_X3Y3_LUT4AB/FrameStrobe[19] Tile_X3Y3_LUT4AB/FrameStrobe[1]
+ Tile_X3Y3_LUT4AB/FrameStrobe[2] Tile_X3Y3_LUT4AB/FrameStrobe[3] Tile_X3Y3_LUT4AB/FrameStrobe[4]
+ Tile_X3Y3_LUT4AB/FrameStrobe[5] Tile_X3Y3_LUT4AB/FrameStrobe[6] Tile_X3Y3_LUT4AB/FrameStrobe[7]
+ Tile_X3Y3_LUT4AB/FrameStrobe[8] Tile_X3Y3_LUT4AB/FrameStrobe[9] Tile_X3Y4_LUT4AB/N1BEG[0]
+ Tile_X3Y4_LUT4AB/N1BEG[1] Tile_X3Y4_LUT4AB/N1BEG[2] Tile_X3Y4_LUT4AB/N1BEG[3] Tile_X3Y5_LUT4AB/N1BEG[0]
+ Tile_X3Y5_LUT4AB/N1BEG[1] Tile_X3Y5_LUT4AB/N1BEG[2] Tile_X3Y5_LUT4AB/N1BEG[3] Tile_X3Y4_LUT4AB/N2BEG[0]
+ Tile_X3Y4_LUT4AB/N2BEG[1] Tile_X3Y4_LUT4AB/N2BEG[2] Tile_X3Y4_LUT4AB/N2BEG[3] Tile_X3Y4_LUT4AB/N2BEG[4]
+ Tile_X3Y4_LUT4AB/N2BEG[5] Tile_X3Y4_LUT4AB/N2BEG[6] Tile_X3Y4_LUT4AB/N2BEG[7] Tile_X3Y3_LUT4AB/N2END[0]
+ Tile_X3Y3_LUT4AB/N2END[1] Tile_X3Y3_LUT4AB/N2END[2] Tile_X3Y3_LUT4AB/N2END[3] Tile_X3Y3_LUT4AB/N2END[4]
+ Tile_X3Y3_LUT4AB/N2END[5] Tile_X3Y3_LUT4AB/N2END[6] Tile_X3Y3_LUT4AB/N2END[7] Tile_X3Y4_LUT4AB/N2END[0]
+ Tile_X3Y4_LUT4AB/N2END[1] Tile_X3Y4_LUT4AB/N2END[2] Tile_X3Y4_LUT4AB/N2END[3] Tile_X3Y4_LUT4AB/N2END[4]
+ Tile_X3Y4_LUT4AB/N2END[5] Tile_X3Y4_LUT4AB/N2END[6] Tile_X3Y4_LUT4AB/N2END[7] Tile_X3Y5_LUT4AB/N2BEG[0]
+ Tile_X3Y5_LUT4AB/N2BEG[1] Tile_X3Y5_LUT4AB/N2BEG[2] Tile_X3Y5_LUT4AB/N2BEG[3] Tile_X3Y5_LUT4AB/N2BEG[4]
+ Tile_X3Y5_LUT4AB/N2BEG[5] Tile_X3Y5_LUT4AB/N2BEG[6] Tile_X3Y5_LUT4AB/N2BEG[7] Tile_X3Y4_LUT4AB/N4BEG[0]
+ Tile_X3Y4_LUT4AB/N4BEG[10] Tile_X3Y4_LUT4AB/N4BEG[11] Tile_X3Y4_LUT4AB/N4BEG[12]
+ Tile_X3Y4_LUT4AB/N4BEG[13] Tile_X3Y4_LUT4AB/N4BEG[14] Tile_X3Y4_LUT4AB/N4BEG[15]
+ Tile_X3Y4_LUT4AB/N4BEG[1] Tile_X3Y4_LUT4AB/N4BEG[2] Tile_X3Y4_LUT4AB/N4BEG[3] Tile_X3Y4_LUT4AB/N4BEG[4]
+ Tile_X3Y4_LUT4AB/N4BEG[5] Tile_X3Y4_LUT4AB/N4BEG[6] Tile_X3Y4_LUT4AB/N4BEG[7] Tile_X3Y4_LUT4AB/N4BEG[8]
+ Tile_X3Y4_LUT4AB/N4BEG[9] Tile_X3Y5_LUT4AB/N4BEG[0] Tile_X3Y5_LUT4AB/N4BEG[10] Tile_X3Y5_LUT4AB/N4BEG[11]
+ Tile_X3Y5_LUT4AB/N4BEG[12] Tile_X3Y5_LUT4AB/N4BEG[13] Tile_X3Y5_LUT4AB/N4BEG[14]
+ Tile_X3Y5_LUT4AB/N4BEG[15] Tile_X3Y5_LUT4AB/N4BEG[1] Tile_X3Y5_LUT4AB/N4BEG[2] Tile_X3Y5_LUT4AB/N4BEG[3]
+ Tile_X3Y5_LUT4AB/N4BEG[4] Tile_X3Y5_LUT4AB/N4BEG[5] Tile_X3Y5_LUT4AB/N4BEG[6] Tile_X3Y5_LUT4AB/N4BEG[7]
+ Tile_X3Y5_LUT4AB/N4BEG[8] Tile_X3Y5_LUT4AB/N4BEG[9] Tile_X3Y4_LUT4AB/NN4BEG[0] Tile_X3Y4_LUT4AB/NN4BEG[10]
+ Tile_X3Y4_LUT4AB/NN4BEG[11] Tile_X3Y4_LUT4AB/NN4BEG[12] Tile_X3Y4_LUT4AB/NN4BEG[13]
+ Tile_X3Y4_LUT4AB/NN4BEG[14] Tile_X3Y4_LUT4AB/NN4BEG[15] Tile_X3Y4_LUT4AB/NN4BEG[1]
+ Tile_X3Y4_LUT4AB/NN4BEG[2] Tile_X3Y4_LUT4AB/NN4BEG[3] Tile_X3Y4_LUT4AB/NN4BEG[4]
+ Tile_X3Y4_LUT4AB/NN4BEG[5] Tile_X3Y4_LUT4AB/NN4BEG[6] Tile_X3Y4_LUT4AB/NN4BEG[7]
+ Tile_X3Y4_LUT4AB/NN4BEG[8] Tile_X3Y4_LUT4AB/NN4BEG[9] Tile_X3Y5_LUT4AB/NN4BEG[0]
+ Tile_X3Y5_LUT4AB/NN4BEG[10] Tile_X3Y5_LUT4AB/NN4BEG[11] Tile_X3Y5_LUT4AB/NN4BEG[12]
+ Tile_X3Y5_LUT4AB/NN4BEG[13] Tile_X3Y5_LUT4AB/NN4BEG[14] Tile_X3Y5_LUT4AB/NN4BEG[15]
+ Tile_X3Y5_LUT4AB/NN4BEG[1] Tile_X3Y5_LUT4AB/NN4BEG[2] Tile_X3Y5_LUT4AB/NN4BEG[3]
+ Tile_X3Y5_LUT4AB/NN4BEG[4] Tile_X3Y5_LUT4AB/NN4BEG[5] Tile_X3Y5_LUT4AB/NN4BEG[6]
+ Tile_X3Y5_LUT4AB/NN4BEG[7] Tile_X3Y5_LUT4AB/NN4BEG[8] Tile_X3Y5_LUT4AB/NN4BEG[9]
+ Tile_X3Y5_LUT4AB/S1END[0] Tile_X3Y5_LUT4AB/S1END[1] Tile_X3Y5_LUT4AB/S1END[2] Tile_X3Y5_LUT4AB/S1END[3]
+ Tile_X3Y4_LUT4AB/S1END[0] Tile_X3Y4_LUT4AB/S1END[1] Tile_X3Y4_LUT4AB/S1END[2] Tile_X3Y4_LUT4AB/S1END[3]
+ Tile_X3Y5_LUT4AB/S2MID[0] Tile_X3Y5_LUT4AB/S2MID[1] Tile_X3Y5_LUT4AB/S2MID[2] Tile_X3Y5_LUT4AB/S2MID[3]
+ Tile_X3Y5_LUT4AB/S2MID[4] Tile_X3Y5_LUT4AB/S2MID[5] Tile_X3Y5_LUT4AB/S2MID[6] Tile_X3Y5_LUT4AB/S2MID[7]
+ Tile_X3Y5_LUT4AB/S2END[0] Tile_X3Y5_LUT4AB/S2END[1] Tile_X3Y5_LUT4AB/S2END[2] Tile_X3Y5_LUT4AB/S2END[3]
+ Tile_X3Y5_LUT4AB/S2END[4] Tile_X3Y5_LUT4AB/S2END[5] Tile_X3Y5_LUT4AB/S2END[6] Tile_X3Y5_LUT4AB/S2END[7]
+ Tile_X3Y4_LUT4AB/S2END[0] Tile_X3Y4_LUT4AB/S2END[1] Tile_X3Y4_LUT4AB/S2END[2] Tile_X3Y4_LUT4AB/S2END[3]
+ Tile_X3Y4_LUT4AB/S2END[4] Tile_X3Y4_LUT4AB/S2END[5] Tile_X3Y4_LUT4AB/S2END[6] Tile_X3Y4_LUT4AB/S2END[7]
+ Tile_X3Y4_LUT4AB/S2MID[0] Tile_X3Y4_LUT4AB/S2MID[1] Tile_X3Y4_LUT4AB/S2MID[2] Tile_X3Y4_LUT4AB/S2MID[3]
+ Tile_X3Y4_LUT4AB/S2MID[4] Tile_X3Y4_LUT4AB/S2MID[5] Tile_X3Y4_LUT4AB/S2MID[6] Tile_X3Y4_LUT4AB/S2MID[7]
+ Tile_X3Y5_LUT4AB/S4END[0] Tile_X3Y5_LUT4AB/S4END[10] Tile_X3Y5_LUT4AB/S4END[11]
+ Tile_X3Y5_LUT4AB/S4END[12] Tile_X3Y5_LUT4AB/S4END[13] Tile_X3Y5_LUT4AB/S4END[14]
+ Tile_X3Y5_LUT4AB/S4END[15] Tile_X3Y5_LUT4AB/S4END[1] Tile_X3Y5_LUT4AB/S4END[2] Tile_X3Y5_LUT4AB/S4END[3]
+ Tile_X3Y5_LUT4AB/S4END[4] Tile_X3Y5_LUT4AB/S4END[5] Tile_X3Y5_LUT4AB/S4END[6] Tile_X3Y5_LUT4AB/S4END[7]
+ Tile_X3Y5_LUT4AB/S4END[8] Tile_X3Y5_LUT4AB/S4END[9] Tile_X3Y4_LUT4AB/S4END[0] Tile_X3Y4_LUT4AB/S4END[10]
+ Tile_X3Y4_LUT4AB/S4END[11] Tile_X3Y4_LUT4AB/S4END[12] Tile_X3Y4_LUT4AB/S4END[13]
+ Tile_X3Y4_LUT4AB/S4END[14] Tile_X3Y4_LUT4AB/S4END[15] Tile_X3Y4_LUT4AB/S4END[1]
+ Tile_X3Y4_LUT4AB/S4END[2] Tile_X3Y4_LUT4AB/S4END[3] Tile_X3Y4_LUT4AB/S4END[4] Tile_X3Y4_LUT4AB/S4END[5]
+ Tile_X3Y4_LUT4AB/S4END[6] Tile_X3Y4_LUT4AB/S4END[7] Tile_X3Y4_LUT4AB/S4END[8] Tile_X3Y4_LUT4AB/S4END[9]
+ Tile_X3Y5_LUT4AB/SS4END[0] Tile_X3Y5_LUT4AB/SS4END[10] Tile_X3Y5_LUT4AB/SS4END[11]
+ Tile_X3Y5_LUT4AB/SS4END[12] Tile_X3Y5_LUT4AB/SS4END[13] Tile_X3Y5_LUT4AB/SS4END[14]
+ Tile_X3Y5_LUT4AB/SS4END[15] Tile_X3Y5_LUT4AB/SS4END[1] Tile_X3Y5_LUT4AB/SS4END[2]
+ Tile_X3Y5_LUT4AB/SS4END[3] Tile_X3Y5_LUT4AB/SS4END[4] Tile_X3Y5_LUT4AB/SS4END[5]
+ Tile_X3Y5_LUT4AB/SS4END[6] Tile_X3Y5_LUT4AB/SS4END[7] Tile_X3Y5_LUT4AB/SS4END[8]
+ Tile_X3Y5_LUT4AB/SS4END[9] Tile_X3Y4_LUT4AB/SS4END[0] Tile_X3Y4_LUT4AB/SS4END[10]
+ Tile_X3Y4_LUT4AB/SS4END[11] Tile_X3Y4_LUT4AB/SS4END[12] Tile_X3Y4_LUT4AB/SS4END[13]
+ Tile_X3Y4_LUT4AB/SS4END[14] Tile_X3Y4_LUT4AB/SS4END[15] Tile_X3Y4_LUT4AB/SS4END[1]
+ Tile_X3Y4_LUT4AB/SS4END[2] Tile_X3Y4_LUT4AB/SS4END[3] Tile_X3Y4_LUT4AB/SS4END[4]
+ Tile_X3Y4_LUT4AB/SS4END[5] Tile_X3Y4_LUT4AB/SS4END[6] Tile_X3Y4_LUT4AB/SS4END[7]
+ Tile_X3Y4_LUT4AB/SS4END[8] Tile_X3Y4_LUT4AB/SS4END[9] Tile_X3Y4_LUT4AB/UserCLK Tile_X3Y3_LUT4AB/UserCLK
+ VGND VPWR Tile_X3Y4_LUT4AB/W1BEG[0] Tile_X3Y4_LUT4AB/W1BEG[1] Tile_X3Y4_LUT4AB/W1BEG[2]
+ Tile_X3Y4_LUT4AB/W1BEG[3] Tile_X4Y4_LUT4AB/W1BEG[0] Tile_X4Y4_LUT4AB/W1BEG[1] Tile_X4Y4_LUT4AB/W1BEG[2]
+ Tile_X4Y4_LUT4AB/W1BEG[3] Tile_X3Y4_LUT4AB/W2BEG[0] Tile_X3Y4_LUT4AB/W2BEG[1] Tile_X3Y4_LUT4AB/W2BEG[2]
+ Tile_X3Y4_LUT4AB/W2BEG[3] Tile_X3Y4_LUT4AB/W2BEG[4] Tile_X3Y4_LUT4AB/W2BEG[5] Tile_X3Y4_LUT4AB/W2BEG[6]
+ Tile_X3Y4_LUT4AB/W2BEG[7] Tile_X2Y4_LUT4AB/W2END[0] Tile_X2Y4_LUT4AB/W2END[1] Tile_X2Y4_LUT4AB/W2END[2]
+ Tile_X2Y4_LUT4AB/W2END[3] Tile_X2Y4_LUT4AB/W2END[4] Tile_X2Y4_LUT4AB/W2END[5] Tile_X2Y4_LUT4AB/W2END[6]
+ Tile_X2Y4_LUT4AB/W2END[7] Tile_X3Y4_LUT4AB/W2END[0] Tile_X3Y4_LUT4AB/W2END[1] Tile_X3Y4_LUT4AB/W2END[2]
+ Tile_X3Y4_LUT4AB/W2END[3] Tile_X3Y4_LUT4AB/W2END[4] Tile_X3Y4_LUT4AB/W2END[5] Tile_X3Y4_LUT4AB/W2END[6]
+ Tile_X3Y4_LUT4AB/W2END[7] Tile_X4Y4_LUT4AB/W2BEG[0] Tile_X4Y4_LUT4AB/W2BEG[1] Tile_X4Y4_LUT4AB/W2BEG[2]
+ Tile_X4Y4_LUT4AB/W2BEG[3] Tile_X4Y4_LUT4AB/W2BEG[4] Tile_X4Y4_LUT4AB/W2BEG[5] Tile_X4Y4_LUT4AB/W2BEG[6]
+ Tile_X4Y4_LUT4AB/W2BEG[7] Tile_X3Y4_LUT4AB/W6BEG[0] Tile_X3Y4_LUT4AB/W6BEG[10] Tile_X3Y4_LUT4AB/W6BEG[11]
+ Tile_X3Y4_LUT4AB/W6BEG[1] Tile_X3Y4_LUT4AB/W6BEG[2] Tile_X3Y4_LUT4AB/W6BEG[3] Tile_X3Y4_LUT4AB/W6BEG[4]
+ Tile_X3Y4_LUT4AB/W6BEG[5] Tile_X3Y4_LUT4AB/W6BEG[6] Tile_X3Y4_LUT4AB/W6BEG[7] Tile_X3Y4_LUT4AB/W6BEG[8]
+ Tile_X3Y4_LUT4AB/W6BEG[9] Tile_X4Y4_LUT4AB/W6BEG[0] Tile_X4Y4_LUT4AB/W6BEG[10] Tile_X4Y4_LUT4AB/W6BEG[11]
+ Tile_X4Y4_LUT4AB/W6BEG[1] Tile_X4Y4_LUT4AB/W6BEG[2] Tile_X4Y4_LUT4AB/W6BEG[3] Tile_X4Y4_LUT4AB/W6BEG[4]
+ Tile_X4Y4_LUT4AB/W6BEG[5] Tile_X4Y4_LUT4AB/W6BEG[6] Tile_X4Y4_LUT4AB/W6BEG[7] Tile_X4Y4_LUT4AB/W6BEG[8]
+ Tile_X4Y4_LUT4AB/W6BEG[9] Tile_X3Y4_LUT4AB/WW4BEG[0] Tile_X3Y4_LUT4AB/WW4BEG[10]
+ Tile_X3Y4_LUT4AB/WW4BEG[11] Tile_X3Y4_LUT4AB/WW4BEG[12] Tile_X3Y4_LUT4AB/WW4BEG[13]
+ Tile_X3Y4_LUT4AB/WW4BEG[14] Tile_X3Y4_LUT4AB/WW4BEG[15] Tile_X3Y4_LUT4AB/WW4BEG[1]
+ Tile_X3Y4_LUT4AB/WW4BEG[2] Tile_X3Y4_LUT4AB/WW4BEG[3] Tile_X3Y4_LUT4AB/WW4BEG[4]
+ Tile_X3Y4_LUT4AB/WW4BEG[5] Tile_X3Y4_LUT4AB/WW4BEG[6] Tile_X3Y4_LUT4AB/WW4BEG[7]
+ Tile_X3Y4_LUT4AB/WW4BEG[8] Tile_X3Y4_LUT4AB/WW4BEG[9] Tile_X4Y4_LUT4AB/WW4BEG[0]
+ Tile_X4Y4_LUT4AB/WW4BEG[10] Tile_X4Y4_LUT4AB/WW4BEG[11] Tile_X4Y4_LUT4AB/WW4BEG[12]
+ Tile_X4Y4_LUT4AB/WW4BEG[13] Tile_X4Y4_LUT4AB/WW4BEG[14] Tile_X4Y4_LUT4AB/WW4BEG[15]
+ Tile_X4Y4_LUT4AB/WW4BEG[1] Tile_X4Y4_LUT4AB/WW4BEG[2] Tile_X4Y4_LUT4AB/WW4BEG[3]
+ Tile_X4Y4_LUT4AB/WW4BEG[4] Tile_X4Y4_LUT4AB/WW4BEG[5] Tile_X4Y4_LUT4AB/WW4BEG[6]
+ Tile_X4Y4_LUT4AB/WW4BEG[7] Tile_X4Y4_LUT4AB/WW4BEG[8] Tile_X4Y4_LUT4AB/WW4BEG[9]
+ LUT4AB
XTile_X5Y7_E_TT_IF Tile_X5Y7_CLK_TT_PROJECT Tile_X4Y7_LUT4AB/E1BEG[0] Tile_X4Y7_LUT4AB/E1BEG[1]
+ Tile_X4Y7_LUT4AB/E1BEG[2] Tile_X4Y7_LUT4AB/E1BEG[3] Tile_X5Y7_E_TT_IF/E2END[0] Tile_X5Y7_E_TT_IF/E2END[1]
+ Tile_X5Y7_E_TT_IF/E2END[2] Tile_X5Y7_E_TT_IF/E2END[3] Tile_X5Y7_E_TT_IF/E2END[4]
+ Tile_X5Y7_E_TT_IF/E2END[5] Tile_X5Y7_E_TT_IF/E2END[6] Tile_X5Y7_E_TT_IF/E2END[7]
+ Tile_X4Y7_LUT4AB/E2BEG[0] Tile_X4Y7_LUT4AB/E2BEG[1] Tile_X4Y7_LUT4AB/E2BEG[2] Tile_X4Y7_LUT4AB/E2BEG[3]
+ Tile_X4Y7_LUT4AB/E2BEG[4] Tile_X4Y7_LUT4AB/E2BEG[5] Tile_X4Y7_LUT4AB/E2BEG[6] Tile_X4Y7_LUT4AB/E2BEG[7]
+ Tile_X4Y7_LUT4AB/E6BEG[0] Tile_X4Y7_LUT4AB/E6BEG[10] Tile_X4Y7_LUT4AB/E6BEG[11]
+ Tile_X4Y7_LUT4AB/E6BEG[1] Tile_X4Y7_LUT4AB/E6BEG[2] Tile_X4Y7_LUT4AB/E6BEG[3] Tile_X4Y7_LUT4AB/E6BEG[4]
+ Tile_X4Y7_LUT4AB/E6BEG[5] Tile_X4Y7_LUT4AB/E6BEG[6] Tile_X4Y7_LUT4AB/E6BEG[7] Tile_X4Y7_LUT4AB/E6BEG[8]
+ Tile_X4Y7_LUT4AB/E6BEG[9] Tile_X4Y7_LUT4AB/EE4BEG[0] Tile_X4Y7_LUT4AB/EE4BEG[10]
+ Tile_X4Y7_LUT4AB/EE4BEG[11] Tile_X4Y7_LUT4AB/EE4BEG[12] Tile_X4Y7_LUT4AB/EE4BEG[13]
+ Tile_X4Y7_LUT4AB/EE4BEG[14] Tile_X4Y7_LUT4AB/EE4BEG[15] Tile_X4Y7_LUT4AB/EE4BEG[1]
+ Tile_X4Y7_LUT4AB/EE4BEG[2] Tile_X4Y7_LUT4AB/EE4BEG[3] Tile_X4Y7_LUT4AB/EE4BEG[4]
+ Tile_X4Y7_LUT4AB/EE4BEG[5] Tile_X4Y7_LUT4AB/EE4BEG[6] Tile_X4Y7_LUT4AB/EE4BEG[7]
+ Tile_X4Y7_LUT4AB/EE4BEG[8] Tile_X4Y7_LUT4AB/EE4BEG[9] Tile_X5Y7_ENA_TT_PROJECT Tile_X5Y7_E_TT_IF/FrameData[0]
+ Tile_X5Y7_E_TT_IF/FrameData[10] Tile_X5Y7_E_TT_IF/FrameData[11] Tile_X5Y7_E_TT_IF/FrameData[12]
+ Tile_X5Y7_E_TT_IF/FrameData[13] Tile_X5Y7_E_TT_IF/FrameData[14] Tile_X5Y7_E_TT_IF/FrameData[15]
+ Tile_X5Y7_E_TT_IF/FrameData[16] Tile_X5Y7_E_TT_IF/FrameData[17] Tile_X5Y7_E_TT_IF/FrameData[18]
+ Tile_X5Y7_E_TT_IF/FrameData[19] Tile_X5Y7_E_TT_IF/FrameData[1] Tile_X5Y7_E_TT_IF/FrameData[20]
+ Tile_X5Y7_E_TT_IF/FrameData[21] Tile_X5Y7_E_TT_IF/FrameData[22] Tile_X5Y7_E_TT_IF/FrameData[23]
+ Tile_X5Y7_E_TT_IF/FrameData[24] Tile_X5Y7_E_TT_IF/FrameData[25] Tile_X5Y7_E_TT_IF/FrameData[26]
+ Tile_X5Y7_E_TT_IF/FrameData[27] Tile_X5Y7_E_TT_IF/FrameData[28] Tile_X5Y7_E_TT_IF/FrameData[29]
+ Tile_X5Y7_E_TT_IF/FrameData[2] Tile_X5Y7_E_TT_IF/FrameData[30] Tile_X5Y7_E_TT_IF/FrameData[31]
+ Tile_X5Y7_E_TT_IF/FrameData[3] Tile_X5Y7_E_TT_IF/FrameData[4] Tile_X5Y7_E_TT_IF/FrameData[5]
+ Tile_X5Y7_E_TT_IF/FrameData[6] Tile_X5Y7_E_TT_IF/FrameData[7] Tile_X5Y7_E_TT_IF/FrameData[8]
+ Tile_X5Y7_E_TT_IF/FrameData[9] Tile_X5Y7_E_TT_IF/FrameData_O[0] Tile_X5Y7_E_TT_IF/FrameData_O[10]
+ Tile_X5Y7_E_TT_IF/FrameData_O[11] Tile_X5Y7_E_TT_IF/FrameData_O[12] Tile_X5Y7_E_TT_IF/FrameData_O[13]
+ Tile_X5Y7_E_TT_IF/FrameData_O[14] Tile_X5Y7_E_TT_IF/FrameData_O[15] Tile_X5Y7_E_TT_IF/FrameData_O[16]
+ Tile_X5Y7_E_TT_IF/FrameData_O[17] Tile_X5Y7_E_TT_IF/FrameData_O[18] Tile_X5Y7_E_TT_IF/FrameData_O[19]
+ Tile_X5Y7_E_TT_IF/FrameData_O[1] Tile_X5Y7_E_TT_IF/FrameData_O[20] Tile_X5Y7_E_TT_IF/FrameData_O[21]
+ Tile_X5Y7_E_TT_IF/FrameData_O[22] Tile_X5Y7_E_TT_IF/FrameData_O[23] Tile_X5Y7_E_TT_IF/FrameData_O[24]
+ Tile_X5Y7_E_TT_IF/FrameData_O[25] Tile_X5Y7_E_TT_IF/FrameData_O[26] Tile_X5Y7_E_TT_IF/FrameData_O[27]
+ Tile_X5Y7_E_TT_IF/FrameData_O[28] Tile_X5Y7_E_TT_IF/FrameData_O[29] Tile_X5Y7_E_TT_IF/FrameData_O[2]
+ Tile_X5Y7_E_TT_IF/FrameData_O[30] Tile_X5Y7_E_TT_IF/FrameData_O[31] Tile_X5Y7_E_TT_IF/FrameData_O[3]
+ Tile_X5Y7_E_TT_IF/FrameData_O[4] Tile_X5Y7_E_TT_IF/FrameData_O[5] Tile_X5Y7_E_TT_IF/FrameData_O[6]
+ Tile_X5Y7_E_TT_IF/FrameData_O[7] Tile_X5Y7_E_TT_IF/FrameData_O[8] Tile_X5Y7_E_TT_IF/FrameData_O[9]
+ Tile_X5Y7_E_TT_IF/FrameStrobe[0] Tile_X5Y7_E_TT_IF/FrameStrobe[10] Tile_X5Y7_E_TT_IF/FrameStrobe[11]
+ Tile_X5Y7_E_TT_IF/FrameStrobe[12] Tile_X5Y7_E_TT_IF/FrameStrobe[13] Tile_X5Y7_E_TT_IF/FrameStrobe[14]
+ Tile_X5Y7_E_TT_IF/FrameStrobe[15] Tile_X5Y7_E_TT_IF/FrameStrobe[16] Tile_X5Y7_E_TT_IF/FrameStrobe[17]
+ Tile_X5Y7_E_TT_IF/FrameStrobe[18] Tile_X5Y7_E_TT_IF/FrameStrobe[19] Tile_X5Y7_E_TT_IF/FrameStrobe[1]
+ Tile_X5Y7_E_TT_IF/FrameStrobe[2] Tile_X5Y7_E_TT_IF/FrameStrobe[3] Tile_X5Y7_E_TT_IF/FrameStrobe[4]
+ Tile_X5Y7_E_TT_IF/FrameStrobe[5] Tile_X5Y7_E_TT_IF/FrameStrobe[6] Tile_X5Y7_E_TT_IF/FrameStrobe[7]
+ Tile_X5Y7_E_TT_IF/FrameStrobe[8] Tile_X5Y7_E_TT_IF/FrameStrobe[9] Tile_X5Y6_E_TT_IF/FrameStrobe[0]
+ Tile_X5Y6_E_TT_IF/FrameStrobe[10] Tile_X5Y6_E_TT_IF/FrameStrobe[11] Tile_X5Y6_E_TT_IF/FrameStrobe[12]
+ Tile_X5Y6_E_TT_IF/FrameStrobe[13] Tile_X5Y6_E_TT_IF/FrameStrobe[14] Tile_X5Y6_E_TT_IF/FrameStrobe[15]
+ Tile_X5Y6_E_TT_IF/FrameStrobe[16] Tile_X5Y6_E_TT_IF/FrameStrobe[17] Tile_X5Y6_E_TT_IF/FrameStrobe[18]
+ Tile_X5Y6_E_TT_IF/FrameStrobe[19] Tile_X5Y6_E_TT_IF/FrameStrobe[1] Tile_X5Y6_E_TT_IF/FrameStrobe[2]
+ Tile_X5Y6_E_TT_IF/FrameStrobe[3] Tile_X5Y6_E_TT_IF/FrameStrobe[4] Tile_X5Y6_E_TT_IF/FrameStrobe[5]
+ Tile_X5Y6_E_TT_IF/FrameStrobe[6] Tile_X5Y6_E_TT_IF/FrameStrobe[7] Tile_X5Y6_E_TT_IF/FrameStrobe[8]
+ Tile_X5Y6_E_TT_IF/FrameStrobe[9] Tile_X5Y7_E_TT_IF/N1BEG[0] Tile_X5Y7_E_TT_IF/N1BEG[1]
+ Tile_X5Y7_E_TT_IF/N1BEG[2] Tile_X5Y7_E_TT_IF/N1BEG[3] Tile_X5Y8_E_TT_IF/N1BEG[0]
+ Tile_X5Y8_E_TT_IF/N1BEG[1] Tile_X5Y8_E_TT_IF/N1BEG[2] Tile_X5Y8_E_TT_IF/N1BEG[3]
+ Tile_X5Y7_E_TT_IF/N2BEG[0] Tile_X5Y7_E_TT_IF/N2BEG[1] Tile_X5Y7_E_TT_IF/N2BEG[2]
+ Tile_X5Y7_E_TT_IF/N2BEG[3] Tile_X5Y7_E_TT_IF/N2BEG[4] Tile_X5Y7_E_TT_IF/N2BEG[5]
+ Tile_X5Y7_E_TT_IF/N2BEG[6] Tile_X5Y7_E_TT_IF/N2BEG[7] Tile_X5Y6_E_TT_IF/N2END[0]
+ Tile_X5Y6_E_TT_IF/N2END[1] Tile_X5Y6_E_TT_IF/N2END[2] Tile_X5Y6_E_TT_IF/N2END[3]
+ Tile_X5Y6_E_TT_IF/N2END[4] Tile_X5Y6_E_TT_IF/N2END[5] Tile_X5Y6_E_TT_IF/N2END[6]
+ Tile_X5Y6_E_TT_IF/N2END[7] Tile_X5Y7_E_TT_IF/N2END[0] Tile_X5Y7_E_TT_IF/N2END[1]
+ Tile_X5Y7_E_TT_IF/N2END[2] Tile_X5Y7_E_TT_IF/N2END[3] Tile_X5Y7_E_TT_IF/N2END[4]
+ Tile_X5Y7_E_TT_IF/N2END[5] Tile_X5Y7_E_TT_IF/N2END[6] Tile_X5Y7_E_TT_IF/N2END[7]
+ Tile_X5Y8_E_TT_IF/N2BEG[0] Tile_X5Y8_E_TT_IF/N2BEG[1] Tile_X5Y8_E_TT_IF/N2BEG[2]
+ Tile_X5Y8_E_TT_IF/N2BEG[3] Tile_X5Y8_E_TT_IF/N2BEG[4] Tile_X5Y8_E_TT_IF/N2BEG[5]
+ Tile_X5Y8_E_TT_IF/N2BEG[6] Tile_X5Y8_E_TT_IF/N2BEG[7] Tile_X5Y7_E_TT_IF/N4BEG[0]
+ Tile_X5Y7_E_TT_IF/N4BEG[10] Tile_X5Y7_E_TT_IF/N4BEG[11] Tile_X5Y7_E_TT_IF/N4BEG[12]
+ Tile_X5Y7_E_TT_IF/N4BEG[13] Tile_X5Y7_E_TT_IF/N4BEG[14] Tile_X5Y7_E_TT_IF/N4BEG[15]
+ Tile_X5Y7_E_TT_IF/N4BEG[1] Tile_X5Y7_E_TT_IF/N4BEG[2] Tile_X5Y7_E_TT_IF/N4BEG[3]
+ Tile_X5Y7_E_TT_IF/N4BEG[4] Tile_X5Y7_E_TT_IF/N4BEG[5] Tile_X5Y7_E_TT_IF/N4BEG[6]
+ Tile_X5Y7_E_TT_IF/N4BEG[7] Tile_X5Y7_E_TT_IF/N4BEG[8] Tile_X5Y7_E_TT_IF/N4BEG[9]
+ Tile_X5Y8_E_TT_IF/N4BEG[0] Tile_X5Y8_E_TT_IF/N4BEG[10] Tile_X5Y8_E_TT_IF/N4BEG[11]
+ Tile_X5Y8_E_TT_IF/N4BEG[12] Tile_X5Y8_E_TT_IF/N4BEG[13] Tile_X5Y8_E_TT_IF/N4BEG[14]
+ Tile_X5Y8_E_TT_IF/N4BEG[15] Tile_X5Y8_E_TT_IF/N4BEG[1] Tile_X5Y8_E_TT_IF/N4BEG[2]
+ Tile_X5Y8_E_TT_IF/N4BEG[3] Tile_X5Y8_E_TT_IF/N4BEG[4] Tile_X5Y8_E_TT_IF/N4BEG[5]
+ Tile_X5Y8_E_TT_IF/N4BEG[6] Tile_X5Y8_E_TT_IF/N4BEG[7] Tile_X5Y8_E_TT_IF/N4BEG[8]
+ Tile_X5Y8_E_TT_IF/N4BEG[9] Tile_X5Y7_RST_N_TT_PROJECT Tile_X5Y8_E_TT_IF/S1END[0]
+ Tile_X5Y8_E_TT_IF/S1END[1] Tile_X5Y8_E_TT_IF/S1END[2] Tile_X5Y8_E_TT_IF/S1END[3]
+ Tile_X5Y7_E_TT_IF/S1END[0] Tile_X5Y7_E_TT_IF/S1END[1] Tile_X5Y7_E_TT_IF/S1END[2]
+ Tile_X5Y7_E_TT_IF/S1END[3] Tile_X5Y8_E_TT_IF/S2MID[0] Tile_X5Y8_E_TT_IF/S2MID[1]
+ Tile_X5Y8_E_TT_IF/S2MID[2] Tile_X5Y8_E_TT_IF/S2MID[3] Tile_X5Y8_E_TT_IF/S2MID[4]
+ Tile_X5Y8_E_TT_IF/S2MID[5] Tile_X5Y8_E_TT_IF/S2MID[6] Tile_X5Y8_E_TT_IF/S2MID[7]
+ Tile_X5Y8_E_TT_IF/S2END[0] Tile_X5Y8_E_TT_IF/S2END[1] Tile_X5Y8_E_TT_IF/S2END[2]
+ Tile_X5Y8_E_TT_IF/S2END[3] Tile_X5Y8_E_TT_IF/S2END[4] Tile_X5Y8_E_TT_IF/S2END[5]
+ Tile_X5Y8_E_TT_IF/S2END[6] Tile_X5Y8_E_TT_IF/S2END[7] Tile_X5Y7_E_TT_IF/S2END[0]
+ Tile_X5Y7_E_TT_IF/S2END[1] Tile_X5Y7_E_TT_IF/S2END[2] Tile_X5Y7_E_TT_IF/S2END[3]
+ Tile_X5Y7_E_TT_IF/S2END[4] Tile_X5Y7_E_TT_IF/S2END[5] Tile_X5Y7_E_TT_IF/S2END[6]
+ Tile_X5Y7_E_TT_IF/S2END[7] Tile_X5Y7_E_TT_IF/S2MID[0] Tile_X5Y7_E_TT_IF/S2MID[1]
+ Tile_X5Y7_E_TT_IF/S2MID[2] Tile_X5Y7_E_TT_IF/S2MID[3] Tile_X5Y7_E_TT_IF/S2MID[4]
+ Tile_X5Y7_E_TT_IF/S2MID[5] Tile_X5Y7_E_TT_IF/S2MID[6] Tile_X5Y7_E_TT_IF/S2MID[7]
+ Tile_X5Y8_E_TT_IF/S4END[0] Tile_X5Y8_E_TT_IF/S4END[10] Tile_X5Y8_E_TT_IF/S4END[11]
+ Tile_X5Y8_E_TT_IF/S4END[12] Tile_X5Y8_E_TT_IF/S4END[13] Tile_X5Y8_E_TT_IF/S4END[14]
+ Tile_X5Y8_E_TT_IF/S4END[15] Tile_X5Y8_E_TT_IF/S4END[1] Tile_X5Y8_E_TT_IF/S4END[2]
+ Tile_X5Y8_E_TT_IF/S4END[3] Tile_X5Y8_E_TT_IF/S4END[4] Tile_X5Y8_E_TT_IF/S4END[5]
+ Tile_X5Y8_E_TT_IF/S4END[6] Tile_X5Y8_E_TT_IF/S4END[7] Tile_X5Y8_E_TT_IF/S4END[8]
+ Tile_X5Y8_E_TT_IF/S4END[9] Tile_X5Y7_E_TT_IF/S4END[0] Tile_X5Y7_E_TT_IF/S4END[10]
+ Tile_X5Y7_E_TT_IF/S4END[11] Tile_X5Y7_E_TT_IF/S4END[12] Tile_X5Y7_E_TT_IF/S4END[13]
+ Tile_X5Y7_E_TT_IF/S4END[14] Tile_X5Y7_E_TT_IF/S4END[15] Tile_X5Y7_E_TT_IF/S4END[1]
+ Tile_X5Y7_E_TT_IF/S4END[2] Tile_X5Y7_E_TT_IF/S4END[3] Tile_X5Y7_E_TT_IF/S4END[4]
+ Tile_X5Y7_E_TT_IF/S4END[5] Tile_X5Y7_E_TT_IF/S4END[6] Tile_X5Y7_E_TT_IF/S4END[7]
+ Tile_X5Y7_E_TT_IF/S4END[8] Tile_X5Y7_E_TT_IF/S4END[9] Tile_X5Y7_UIO_IN_TT_PROJECT0
+ Tile_X5Y7_UIO_IN_TT_PROJECT1 Tile_X5Y7_UIO_IN_TT_PROJECT2 Tile_X5Y7_UIO_IN_TT_PROJECT3
+ Tile_X5Y7_UIO_IN_TT_PROJECT4 Tile_X5Y7_UIO_IN_TT_PROJECT5 Tile_X5Y7_UIO_IN_TT_PROJECT6
+ Tile_X5Y7_UIO_IN_TT_PROJECT7 Tile_X5Y7_UIO_OE_TT_PROJECT0 Tile_X5Y7_UIO_OE_TT_PROJECT1
+ Tile_X5Y7_UIO_OE_TT_PROJECT2 Tile_X5Y7_UIO_OE_TT_PROJECT3 Tile_X5Y7_UIO_OE_TT_PROJECT4
+ Tile_X5Y7_UIO_OE_TT_PROJECT5 Tile_X5Y7_UIO_OE_TT_PROJECT6 Tile_X5Y7_UIO_OE_TT_PROJECT7
+ Tile_X5Y7_UIO_OUT_TT_PROJECT0 Tile_X5Y7_UIO_OUT_TT_PROJECT1 Tile_X5Y7_UIO_OUT_TT_PROJECT2
+ Tile_X5Y7_UIO_OUT_TT_PROJECT3 Tile_X5Y7_UIO_OUT_TT_PROJECT4 Tile_X5Y7_UIO_OUT_TT_PROJECT5
+ Tile_X5Y7_UIO_OUT_TT_PROJECT6 Tile_X5Y7_UIO_OUT_TT_PROJECT7 Tile_X5Y7_UI_IN_TT_PROJECT0
+ Tile_X5Y7_UI_IN_TT_PROJECT1 Tile_X5Y7_UI_IN_TT_PROJECT2 Tile_X5Y7_UI_IN_TT_PROJECT3
+ Tile_X5Y7_UI_IN_TT_PROJECT4 Tile_X5Y7_UI_IN_TT_PROJECT5 Tile_X5Y7_UI_IN_TT_PROJECT6
+ Tile_X5Y7_UI_IN_TT_PROJECT7 Tile_X5Y7_UO_OUT_TT_PROJECT0 Tile_X5Y7_UO_OUT_TT_PROJECT1
+ Tile_X5Y7_UO_OUT_TT_PROJECT2 Tile_X5Y7_UO_OUT_TT_PROJECT3 Tile_X5Y7_UO_OUT_TT_PROJECT4
+ Tile_X5Y7_UO_OUT_TT_PROJECT5 Tile_X5Y7_UO_OUT_TT_PROJECT6 Tile_X5Y7_UO_OUT_TT_PROJECT7
+ Tile_X5Y7_E_TT_IF/UserCLK Tile_X5Y6_E_TT_IF/UserCLK VGND VPWR Tile_X4Y7_LUT4AB/W1END[0]
+ Tile_X4Y7_LUT4AB/W1END[1] Tile_X4Y7_LUT4AB/W1END[2] Tile_X4Y7_LUT4AB/W1END[3] Tile_X4Y7_LUT4AB/W2MID[0]
+ Tile_X4Y7_LUT4AB/W2MID[1] Tile_X4Y7_LUT4AB/W2MID[2] Tile_X4Y7_LUT4AB/W2MID[3] Tile_X4Y7_LUT4AB/W2MID[4]
+ Tile_X4Y7_LUT4AB/W2MID[5] Tile_X4Y7_LUT4AB/W2MID[6] Tile_X4Y7_LUT4AB/W2MID[7] Tile_X4Y7_LUT4AB/W2END[0]
+ Tile_X4Y7_LUT4AB/W2END[1] Tile_X4Y7_LUT4AB/W2END[2] Tile_X4Y7_LUT4AB/W2END[3] Tile_X4Y7_LUT4AB/W2END[4]
+ Tile_X4Y7_LUT4AB/W2END[5] Tile_X4Y7_LUT4AB/W2END[6] Tile_X4Y7_LUT4AB/W2END[7] Tile_X4Y7_LUT4AB/W6END[0]
+ Tile_X4Y7_LUT4AB/W6END[10] Tile_X4Y7_LUT4AB/W6END[11] Tile_X4Y7_LUT4AB/W6END[1]
+ Tile_X4Y7_LUT4AB/W6END[2] Tile_X4Y7_LUT4AB/W6END[3] Tile_X4Y7_LUT4AB/W6END[4] Tile_X4Y7_LUT4AB/W6END[5]
+ Tile_X4Y7_LUT4AB/W6END[6] Tile_X4Y7_LUT4AB/W6END[7] Tile_X4Y7_LUT4AB/W6END[8] Tile_X4Y7_LUT4AB/W6END[9]
+ Tile_X4Y7_LUT4AB/WW4END[0] Tile_X4Y7_LUT4AB/WW4END[10] Tile_X4Y7_LUT4AB/WW4END[11]
+ Tile_X4Y7_LUT4AB/WW4END[12] Tile_X4Y7_LUT4AB/WW4END[13] Tile_X4Y7_LUT4AB/WW4END[14]
+ Tile_X4Y7_LUT4AB/WW4END[15] Tile_X4Y7_LUT4AB/WW4END[1] Tile_X4Y7_LUT4AB/WW4END[2]
+ Tile_X4Y7_LUT4AB/WW4END[3] Tile_X4Y7_LUT4AB/WW4END[4] Tile_X4Y7_LUT4AB/WW4END[5]
+ Tile_X4Y7_LUT4AB/WW4END[6] Tile_X4Y7_LUT4AB/WW4END[7] Tile_X4Y7_LUT4AB/WW4END[8]
+ Tile_X4Y7_LUT4AB/WW4END[9] E_TT_IF
XTile_X2Y8_LUT4AB Tile_X2Y9_S_IO4/Co Tile_X2Y8_LUT4AB/Co Tile_X3Y8_LUT4AB/E1END[0]
+ Tile_X3Y8_LUT4AB/E1END[1] Tile_X3Y8_LUT4AB/E1END[2] Tile_X3Y8_LUT4AB/E1END[3] Tile_X2Y8_LUT4AB/E1END[0]
+ Tile_X2Y8_LUT4AB/E1END[1] Tile_X2Y8_LUT4AB/E1END[2] Tile_X2Y8_LUT4AB/E1END[3] Tile_X3Y8_LUT4AB/E2MID[0]
+ Tile_X3Y8_LUT4AB/E2MID[1] Tile_X3Y8_LUT4AB/E2MID[2] Tile_X3Y8_LUT4AB/E2MID[3] Tile_X3Y8_LUT4AB/E2MID[4]
+ Tile_X3Y8_LUT4AB/E2MID[5] Tile_X3Y8_LUT4AB/E2MID[6] Tile_X3Y8_LUT4AB/E2MID[7] Tile_X3Y8_LUT4AB/E2END[0]
+ Tile_X3Y8_LUT4AB/E2END[1] Tile_X3Y8_LUT4AB/E2END[2] Tile_X3Y8_LUT4AB/E2END[3] Tile_X3Y8_LUT4AB/E2END[4]
+ Tile_X3Y8_LUT4AB/E2END[5] Tile_X3Y8_LUT4AB/E2END[6] Tile_X3Y8_LUT4AB/E2END[7] Tile_X2Y8_LUT4AB/E2END[0]
+ Tile_X2Y8_LUT4AB/E2END[1] Tile_X2Y8_LUT4AB/E2END[2] Tile_X2Y8_LUT4AB/E2END[3] Tile_X2Y8_LUT4AB/E2END[4]
+ Tile_X2Y8_LUT4AB/E2END[5] Tile_X2Y8_LUT4AB/E2END[6] Tile_X2Y8_LUT4AB/E2END[7] Tile_X2Y8_LUT4AB/E2MID[0]
+ Tile_X2Y8_LUT4AB/E2MID[1] Tile_X2Y8_LUT4AB/E2MID[2] Tile_X2Y8_LUT4AB/E2MID[3] Tile_X2Y8_LUT4AB/E2MID[4]
+ Tile_X2Y8_LUT4AB/E2MID[5] Tile_X2Y8_LUT4AB/E2MID[6] Tile_X2Y8_LUT4AB/E2MID[7] Tile_X3Y8_LUT4AB/E6END[0]
+ Tile_X3Y8_LUT4AB/E6END[10] Tile_X3Y8_LUT4AB/E6END[11] Tile_X3Y8_LUT4AB/E6END[1]
+ Tile_X3Y8_LUT4AB/E6END[2] Tile_X3Y8_LUT4AB/E6END[3] Tile_X3Y8_LUT4AB/E6END[4] Tile_X3Y8_LUT4AB/E6END[5]
+ Tile_X3Y8_LUT4AB/E6END[6] Tile_X3Y8_LUT4AB/E6END[7] Tile_X3Y8_LUT4AB/E6END[8] Tile_X3Y8_LUT4AB/E6END[9]
+ Tile_X2Y8_LUT4AB/E6END[0] Tile_X2Y8_LUT4AB/E6END[10] Tile_X2Y8_LUT4AB/E6END[11]
+ Tile_X2Y8_LUT4AB/E6END[1] Tile_X2Y8_LUT4AB/E6END[2] Tile_X2Y8_LUT4AB/E6END[3] Tile_X2Y8_LUT4AB/E6END[4]
+ Tile_X2Y8_LUT4AB/E6END[5] Tile_X2Y8_LUT4AB/E6END[6] Tile_X2Y8_LUT4AB/E6END[7] Tile_X2Y8_LUT4AB/E6END[8]
+ Tile_X2Y8_LUT4AB/E6END[9] Tile_X3Y8_LUT4AB/EE4END[0] Tile_X3Y8_LUT4AB/EE4END[10]
+ Tile_X3Y8_LUT4AB/EE4END[11] Tile_X3Y8_LUT4AB/EE4END[12] Tile_X3Y8_LUT4AB/EE4END[13]
+ Tile_X3Y8_LUT4AB/EE4END[14] Tile_X3Y8_LUT4AB/EE4END[15] Tile_X3Y8_LUT4AB/EE4END[1]
+ Tile_X3Y8_LUT4AB/EE4END[2] Tile_X3Y8_LUT4AB/EE4END[3] Tile_X3Y8_LUT4AB/EE4END[4]
+ Tile_X3Y8_LUT4AB/EE4END[5] Tile_X3Y8_LUT4AB/EE4END[6] Tile_X3Y8_LUT4AB/EE4END[7]
+ Tile_X3Y8_LUT4AB/EE4END[8] Tile_X3Y8_LUT4AB/EE4END[9] Tile_X2Y8_LUT4AB/EE4END[0]
+ Tile_X2Y8_LUT4AB/EE4END[10] Tile_X2Y8_LUT4AB/EE4END[11] Tile_X2Y8_LUT4AB/EE4END[12]
+ Tile_X2Y8_LUT4AB/EE4END[13] Tile_X2Y8_LUT4AB/EE4END[14] Tile_X2Y8_LUT4AB/EE4END[15]
+ Tile_X2Y8_LUT4AB/EE4END[1] Tile_X2Y8_LUT4AB/EE4END[2] Tile_X2Y8_LUT4AB/EE4END[3]
+ Tile_X2Y8_LUT4AB/EE4END[4] Tile_X2Y8_LUT4AB/EE4END[5] Tile_X2Y8_LUT4AB/EE4END[6]
+ Tile_X2Y8_LUT4AB/EE4END[7] Tile_X2Y8_LUT4AB/EE4END[8] Tile_X2Y8_LUT4AB/EE4END[9]
+ Tile_X2Y8_LUT4AB/FrameData[0] Tile_X2Y8_LUT4AB/FrameData[10] Tile_X2Y8_LUT4AB/FrameData[11]
+ Tile_X2Y8_LUT4AB/FrameData[12] Tile_X2Y8_LUT4AB/FrameData[13] Tile_X2Y8_LUT4AB/FrameData[14]
+ Tile_X2Y8_LUT4AB/FrameData[15] Tile_X2Y8_LUT4AB/FrameData[16] Tile_X2Y8_LUT4AB/FrameData[17]
+ Tile_X2Y8_LUT4AB/FrameData[18] Tile_X2Y8_LUT4AB/FrameData[19] Tile_X2Y8_LUT4AB/FrameData[1]
+ Tile_X2Y8_LUT4AB/FrameData[20] Tile_X2Y8_LUT4AB/FrameData[21] Tile_X2Y8_LUT4AB/FrameData[22]
+ Tile_X2Y8_LUT4AB/FrameData[23] Tile_X2Y8_LUT4AB/FrameData[24] Tile_X2Y8_LUT4AB/FrameData[25]
+ Tile_X2Y8_LUT4AB/FrameData[26] Tile_X2Y8_LUT4AB/FrameData[27] Tile_X2Y8_LUT4AB/FrameData[28]
+ Tile_X2Y8_LUT4AB/FrameData[29] Tile_X2Y8_LUT4AB/FrameData[2] Tile_X2Y8_LUT4AB/FrameData[30]
+ Tile_X2Y8_LUT4AB/FrameData[31] Tile_X2Y8_LUT4AB/FrameData[3] Tile_X2Y8_LUT4AB/FrameData[4]
+ Tile_X2Y8_LUT4AB/FrameData[5] Tile_X2Y8_LUT4AB/FrameData[6] Tile_X2Y8_LUT4AB/FrameData[7]
+ Tile_X2Y8_LUT4AB/FrameData[8] Tile_X2Y8_LUT4AB/FrameData[9] Tile_X3Y8_LUT4AB/FrameData[0]
+ Tile_X3Y8_LUT4AB/FrameData[10] Tile_X3Y8_LUT4AB/FrameData[11] Tile_X3Y8_LUT4AB/FrameData[12]
+ Tile_X3Y8_LUT4AB/FrameData[13] Tile_X3Y8_LUT4AB/FrameData[14] Tile_X3Y8_LUT4AB/FrameData[15]
+ Tile_X3Y8_LUT4AB/FrameData[16] Tile_X3Y8_LUT4AB/FrameData[17] Tile_X3Y8_LUT4AB/FrameData[18]
+ Tile_X3Y8_LUT4AB/FrameData[19] Tile_X3Y8_LUT4AB/FrameData[1] Tile_X3Y8_LUT4AB/FrameData[20]
+ Tile_X3Y8_LUT4AB/FrameData[21] Tile_X3Y8_LUT4AB/FrameData[22] Tile_X3Y8_LUT4AB/FrameData[23]
+ Tile_X3Y8_LUT4AB/FrameData[24] Tile_X3Y8_LUT4AB/FrameData[25] Tile_X3Y8_LUT4AB/FrameData[26]
+ Tile_X3Y8_LUT4AB/FrameData[27] Tile_X3Y8_LUT4AB/FrameData[28] Tile_X3Y8_LUT4AB/FrameData[29]
+ Tile_X3Y8_LUT4AB/FrameData[2] Tile_X3Y8_LUT4AB/FrameData[30] Tile_X3Y8_LUT4AB/FrameData[31]
+ Tile_X3Y8_LUT4AB/FrameData[3] Tile_X3Y8_LUT4AB/FrameData[4] Tile_X3Y8_LUT4AB/FrameData[5]
+ Tile_X3Y8_LUT4AB/FrameData[6] Tile_X3Y8_LUT4AB/FrameData[7] Tile_X3Y8_LUT4AB/FrameData[8]
+ Tile_X3Y8_LUT4AB/FrameData[9] Tile_X2Y8_LUT4AB/FrameStrobe[0] Tile_X2Y8_LUT4AB/FrameStrobe[10]
+ Tile_X2Y8_LUT4AB/FrameStrobe[11] Tile_X2Y8_LUT4AB/FrameStrobe[12] Tile_X2Y8_LUT4AB/FrameStrobe[13]
+ Tile_X2Y8_LUT4AB/FrameStrobe[14] Tile_X2Y8_LUT4AB/FrameStrobe[15] Tile_X2Y8_LUT4AB/FrameStrobe[16]
+ Tile_X2Y8_LUT4AB/FrameStrobe[17] Tile_X2Y8_LUT4AB/FrameStrobe[18] Tile_X2Y8_LUT4AB/FrameStrobe[19]
+ Tile_X2Y8_LUT4AB/FrameStrobe[1] Tile_X2Y8_LUT4AB/FrameStrobe[2] Tile_X2Y8_LUT4AB/FrameStrobe[3]
+ Tile_X2Y8_LUT4AB/FrameStrobe[4] Tile_X2Y8_LUT4AB/FrameStrobe[5] Tile_X2Y8_LUT4AB/FrameStrobe[6]
+ Tile_X2Y8_LUT4AB/FrameStrobe[7] Tile_X2Y8_LUT4AB/FrameStrobe[8] Tile_X2Y8_LUT4AB/FrameStrobe[9]
+ Tile_X2Y7_LUT4AB/FrameStrobe[0] Tile_X2Y7_LUT4AB/FrameStrobe[10] Tile_X2Y7_LUT4AB/FrameStrobe[11]
+ Tile_X2Y7_LUT4AB/FrameStrobe[12] Tile_X2Y7_LUT4AB/FrameStrobe[13] Tile_X2Y7_LUT4AB/FrameStrobe[14]
+ Tile_X2Y7_LUT4AB/FrameStrobe[15] Tile_X2Y7_LUT4AB/FrameStrobe[16] Tile_X2Y7_LUT4AB/FrameStrobe[17]
+ Tile_X2Y7_LUT4AB/FrameStrobe[18] Tile_X2Y7_LUT4AB/FrameStrobe[19] Tile_X2Y7_LUT4AB/FrameStrobe[1]
+ Tile_X2Y7_LUT4AB/FrameStrobe[2] Tile_X2Y7_LUT4AB/FrameStrobe[3] Tile_X2Y7_LUT4AB/FrameStrobe[4]
+ Tile_X2Y7_LUT4AB/FrameStrobe[5] Tile_X2Y7_LUT4AB/FrameStrobe[6] Tile_X2Y7_LUT4AB/FrameStrobe[7]
+ Tile_X2Y7_LUT4AB/FrameStrobe[8] Tile_X2Y7_LUT4AB/FrameStrobe[9] Tile_X2Y8_LUT4AB/N1BEG[0]
+ Tile_X2Y8_LUT4AB/N1BEG[1] Tile_X2Y8_LUT4AB/N1BEG[2] Tile_X2Y8_LUT4AB/N1BEG[3] Tile_X2Y9_S_IO4/N1BEG[0]
+ Tile_X2Y9_S_IO4/N1BEG[1] Tile_X2Y9_S_IO4/N1BEG[2] Tile_X2Y9_S_IO4/N1BEG[3] Tile_X2Y8_LUT4AB/N2BEG[0]
+ Tile_X2Y8_LUT4AB/N2BEG[1] Tile_X2Y8_LUT4AB/N2BEG[2] Tile_X2Y8_LUT4AB/N2BEG[3] Tile_X2Y8_LUT4AB/N2BEG[4]
+ Tile_X2Y8_LUT4AB/N2BEG[5] Tile_X2Y8_LUT4AB/N2BEG[6] Tile_X2Y8_LUT4AB/N2BEG[7] Tile_X2Y7_LUT4AB/N2END[0]
+ Tile_X2Y7_LUT4AB/N2END[1] Tile_X2Y7_LUT4AB/N2END[2] Tile_X2Y7_LUT4AB/N2END[3] Tile_X2Y7_LUT4AB/N2END[4]
+ Tile_X2Y7_LUT4AB/N2END[5] Tile_X2Y7_LUT4AB/N2END[6] Tile_X2Y7_LUT4AB/N2END[7] Tile_X2Y9_S_IO4/N2BEGb[0]
+ Tile_X2Y9_S_IO4/N2BEGb[1] Tile_X2Y9_S_IO4/N2BEGb[2] Tile_X2Y9_S_IO4/N2BEGb[3] Tile_X2Y9_S_IO4/N2BEGb[4]
+ Tile_X2Y9_S_IO4/N2BEGb[5] Tile_X2Y9_S_IO4/N2BEGb[6] Tile_X2Y9_S_IO4/N2BEGb[7] Tile_X2Y9_S_IO4/N2BEG[0]
+ Tile_X2Y9_S_IO4/N2BEG[1] Tile_X2Y9_S_IO4/N2BEG[2] Tile_X2Y9_S_IO4/N2BEG[3] Tile_X2Y9_S_IO4/N2BEG[4]
+ Tile_X2Y9_S_IO4/N2BEG[5] Tile_X2Y9_S_IO4/N2BEG[6] Tile_X2Y9_S_IO4/N2BEG[7] Tile_X2Y8_LUT4AB/N4BEG[0]
+ Tile_X2Y8_LUT4AB/N4BEG[10] Tile_X2Y8_LUT4AB/N4BEG[11] Tile_X2Y8_LUT4AB/N4BEG[12]
+ Tile_X2Y8_LUT4AB/N4BEG[13] Tile_X2Y8_LUT4AB/N4BEG[14] Tile_X2Y8_LUT4AB/N4BEG[15]
+ Tile_X2Y8_LUT4AB/N4BEG[1] Tile_X2Y8_LUT4AB/N4BEG[2] Tile_X2Y8_LUT4AB/N4BEG[3] Tile_X2Y8_LUT4AB/N4BEG[4]
+ Tile_X2Y8_LUT4AB/N4BEG[5] Tile_X2Y8_LUT4AB/N4BEG[6] Tile_X2Y8_LUT4AB/N4BEG[7] Tile_X2Y8_LUT4AB/N4BEG[8]
+ Tile_X2Y8_LUT4AB/N4BEG[9] Tile_X2Y9_S_IO4/N4BEG[0] Tile_X2Y9_S_IO4/N4BEG[10] Tile_X2Y9_S_IO4/N4BEG[11]
+ Tile_X2Y9_S_IO4/N4BEG[12] Tile_X2Y9_S_IO4/N4BEG[13] Tile_X2Y9_S_IO4/N4BEG[14] Tile_X2Y9_S_IO4/N4BEG[15]
+ Tile_X2Y9_S_IO4/N4BEG[1] Tile_X2Y9_S_IO4/N4BEG[2] Tile_X2Y9_S_IO4/N4BEG[3] Tile_X2Y9_S_IO4/N4BEG[4]
+ Tile_X2Y9_S_IO4/N4BEG[5] Tile_X2Y9_S_IO4/N4BEG[6] Tile_X2Y9_S_IO4/N4BEG[7] Tile_X2Y9_S_IO4/N4BEG[8]
+ Tile_X2Y9_S_IO4/N4BEG[9] Tile_X2Y8_LUT4AB/NN4BEG[0] Tile_X2Y8_LUT4AB/NN4BEG[10]
+ Tile_X2Y8_LUT4AB/NN4BEG[11] Tile_X2Y8_LUT4AB/NN4BEG[12] Tile_X2Y8_LUT4AB/NN4BEG[13]
+ Tile_X2Y8_LUT4AB/NN4BEG[14] Tile_X2Y8_LUT4AB/NN4BEG[15] Tile_X2Y8_LUT4AB/NN4BEG[1]
+ Tile_X2Y8_LUT4AB/NN4BEG[2] Tile_X2Y8_LUT4AB/NN4BEG[3] Tile_X2Y8_LUT4AB/NN4BEG[4]
+ Tile_X2Y8_LUT4AB/NN4BEG[5] Tile_X2Y8_LUT4AB/NN4BEG[6] Tile_X2Y8_LUT4AB/NN4BEG[7]
+ Tile_X2Y8_LUT4AB/NN4BEG[8] Tile_X2Y8_LUT4AB/NN4BEG[9] Tile_X2Y9_S_IO4/NN4BEG[0]
+ Tile_X2Y9_S_IO4/NN4BEG[10] Tile_X2Y9_S_IO4/NN4BEG[11] Tile_X2Y9_S_IO4/NN4BEG[12]
+ Tile_X2Y9_S_IO4/NN4BEG[13] Tile_X2Y9_S_IO4/NN4BEG[14] Tile_X2Y9_S_IO4/NN4BEG[15]
+ Tile_X2Y9_S_IO4/NN4BEG[1] Tile_X2Y9_S_IO4/NN4BEG[2] Tile_X2Y9_S_IO4/NN4BEG[3] Tile_X2Y9_S_IO4/NN4BEG[4]
+ Tile_X2Y9_S_IO4/NN4BEG[5] Tile_X2Y9_S_IO4/NN4BEG[6] Tile_X2Y9_S_IO4/NN4BEG[7] Tile_X2Y9_S_IO4/NN4BEG[8]
+ Tile_X2Y9_S_IO4/NN4BEG[9] Tile_X2Y9_S_IO4/S1END[0] Tile_X2Y9_S_IO4/S1END[1] Tile_X2Y9_S_IO4/S1END[2]
+ Tile_X2Y9_S_IO4/S1END[3] Tile_X2Y8_LUT4AB/S1END[0] Tile_X2Y8_LUT4AB/S1END[1] Tile_X2Y8_LUT4AB/S1END[2]
+ Tile_X2Y8_LUT4AB/S1END[3] Tile_X2Y9_S_IO4/S2MID[0] Tile_X2Y9_S_IO4/S2MID[1] Tile_X2Y9_S_IO4/S2MID[2]
+ Tile_X2Y9_S_IO4/S2MID[3] Tile_X2Y9_S_IO4/S2MID[4] Tile_X2Y9_S_IO4/S2MID[5] Tile_X2Y9_S_IO4/S2MID[6]
+ Tile_X2Y9_S_IO4/S2MID[7] Tile_X2Y9_S_IO4/S2END[0] Tile_X2Y9_S_IO4/S2END[1] Tile_X2Y9_S_IO4/S2END[2]
+ Tile_X2Y9_S_IO4/S2END[3] Tile_X2Y9_S_IO4/S2END[4] Tile_X2Y9_S_IO4/S2END[5] Tile_X2Y9_S_IO4/S2END[6]
+ Tile_X2Y9_S_IO4/S2END[7] Tile_X2Y8_LUT4AB/S2END[0] Tile_X2Y8_LUT4AB/S2END[1] Tile_X2Y8_LUT4AB/S2END[2]
+ Tile_X2Y8_LUT4AB/S2END[3] Tile_X2Y8_LUT4AB/S2END[4] Tile_X2Y8_LUT4AB/S2END[5] Tile_X2Y8_LUT4AB/S2END[6]
+ Tile_X2Y8_LUT4AB/S2END[7] Tile_X2Y8_LUT4AB/S2MID[0] Tile_X2Y8_LUT4AB/S2MID[1] Tile_X2Y8_LUT4AB/S2MID[2]
+ Tile_X2Y8_LUT4AB/S2MID[3] Tile_X2Y8_LUT4AB/S2MID[4] Tile_X2Y8_LUT4AB/S2MID[5] Tile_X2Y8_LUT4AB/S2MID[6]
+ Tile_X2Y8_LUT4AB/S2MID[7] Tile_X2Y9_S_IO4/S4END[0] Tile_X2Y9_S_IO4/S4END[10] Tile_X2Y9_S_IO4/S4END[11]
+ Tile_X2Y9_S_IO4/S4END[12] Tile_X2Y9_S_IO4/S4END[13] Tile_X2Y9_S_IO4/S4END[14] Tile_X2Y9_S_IO4/S4END[15]
+ Tile_X2Y9_S_IO4/S4END[1] Tile_X2Y9_S_IO4/S4END[2] Tile_X2Y9_S_IO4/S4END[3] Tile_X2Y9_S_IO4/S4END[4]
+ Tile_X2Y9_S_IO4/S4END[5] Tile_X2Y9_S_IO4/S4END[6] Tile_X2Y9_S_IO4/S4END[7] Tile_X2Y9_S_IO4/S4END[8]
+ Tile_X2Y9_S_IO4/S4END[9] Tile_X2Y8_LUT4AB/S4END[0] Tile_X2Y8_LUT4AB/S4END[10] Tile_X2Y8_LUT4AB/S4END[11]
+ Tile_X2Y8_LUT4AB/S4END[12] Tile_X2Y8_LUT4AB/S4END[13] Tile_X2Y8_LUT4AB/S4END[14]
+ Tile_X2Y8_LUT4AB/S4END[15] Tile_X2Y8_LUT4AB/S4END[1] Tile_X2Y8_LUT4AB/S4END[2] Tile_X2Y8_LUT4AB/S4END[3]
+ Tile_X2Y8_LUT4AB/S4END[4] Tile_X2Y8_LUT4AB/S4END[5] Tile_X2Y8_LUT4AB/S4END[6] Tile_X2Y8_LUT4AB/S4END[7]
+ Tile_X2Y8_LUT4AB/S4END[8] Tile_X2Y8_LUT4AB/S4END[9] Tile_X2Y9_S_IO4/SS4END[0] Tile_X2Y9_S_IO4/SS4END[10]
+ Tile_X2Y9_S_IO4/SS4END[11] Tile_X2Y9_S_IO4/SS4END[12] Tile_X2Y9_S_IO4/SS4END[13]
+ Tile_X2Y9_S_IO4/SS4END[14] Tile_X2Y9_S_IO4/SS4END[15] Tile_X2Y9_S_IO4/SS4END[1]
+ Tile_X2Y9_S_IO4/SS4END[2] Tile_X2Y9_S_IO4/SS4END[3] Tile_X2Y9_S_IO4/SS4END[4] Tile_X2Y9_S_IO4/SS4END[5]
+ Tile_X2Y9_S_IO4/SS4END[6] Tile_X2Y9_S_IO4/SS4END[7] Tile_X2Y9_S_IO4/SS4END[8] Tile_X2Y9_S_IO4/SS4END[9]
+ Tile_X2Y8_LUT4AB/SS4END[0] Tile_X2Y8_LUT4AB/SS4END[10] Tile_X2Y8_LUT4AB/SS4END[11]
+ Tile_X2Y8_LUT4AB/SS4END[12] Tile_X2Y8_LUT4AB/SS4END[13] Tile_X2Y8_LUT4AB/SS4END[14]
+ Tile_X2Y8_LUT4AB/SS4END[15] Tile_X2Y8_LUT4AB/SS4END[1] Tile_X2Y8_LUT4AB/SS4END[2]
+ Tile_X2Y8_LUT4AB/SS4END[3] Tile_X2Y8_LUT4AB/SS4END[4] Tile_X2Y8_LUT4AB/SS4END[5]
+ Tile_X2Y8_LUT4AB/SS4END[6] Tile_X2Y8_LUT4AB/SS4END[7] Tile_X2Y8_LUT4AB/SS4END[8]
+ Tile_X2Y8_LUT4AB/SS4END[9] Tile_X2Y9_S_IO4/UserCLKo Tile_X2Y7_LUT4AB/UserCLK VGND
+ VPWR Tile_X2Y8_LUT4AB/W1BEG[0] Tile_X2Y8_LUT4AB/W1BEG[1] Tile_X2Y8_LUT4AB/W1BEG[2]
+ Tile_X2Y8_LUT4AB/W1BEG[3] Tile_X3Y8_LUT4AB/W1BEG[0] Tile_X3Y8_LUT4AB/W1BEG[1] Tile_X3Y8_LUT4AB/W1BEG[2]
+ Tile_X3Y8_LUT4AB/W1BEG[3] Tile_X2Y8_LUT4AB/W2BEG[0] Tile_X2Y8_LUT4AB/W2BEG[1] Tile_X2Y8_LUT4AB/W2BEG[2]
+ Tile_X2Y8_LUT4AB/W2BEG[3] Tile_X2Y8_LUT4AB/W2BEG[4] Tile_X2Y8_LUT4AB/W2BEG[5] Tile_X2Y8_LUT4AB/W2BEG[6]
+ Tile_X2Y8_LUT4AB/W2BEG[7] Tile_X1Y8_LUT4AB/W2END[0] Tile_X1Y8_LUT4AB/W2END[1] Tile_X1Y8_LUT4AB/W2END[2]
+ Tile_X1Y8_LUT4AB/W2END[3] Tile_X1Y8_LUT4AB/W2END[4] Tile_X1Y8_LUT4AB/W2END[5] Tile_X1Y8_LUT4AB/W2END[6]
+ Tile_X1Y8_LUT4AB/W2END[7] Tile_X2Y8_LUT4AB/W2END[0] Tile_X2Y8_LUT4AB/W2END[1] Tile_X2Y8_LUT4AB/W2END[2]
+ Tile_X2Y8_LUT4AB/W2END[3] Tile_X2Y8_LUT4AB/W2END[4] Tile_X2Y8_LUT4AB/W2END[5] Tile_X2Y8_LUT4AB/W2END[6]
+ Tile_X2Y8_LUT4AB/W2END[7] Tile_X3Y8_LUT4AB/W2BEG[0] Tile_X3Y8_LUT4AB/W2BEG[1] Tile_X3Y8_LUT4AB/W2BEG[2]
+ Tile_X3Y8_LUT4AB/W2BEG[3] Tile_X3Y8_LUT4AB/W2BEG[4] Tile_X3Y8_LUT4AB/W2BEG[5] Tile_X3Y8_LUT4AB/W2BEG[6]
+ Tile_X3Y8_LUT4AB/W2BEG[7] Tile_X2Y8_LUT4AB/W6BEG[0] Tile_X2Y8_LUT4AB/W6BEG[10] Tile_X2Y8_LUT4AB/W6BEG[11]
+ Tile_X2Y8_LUT4AB/W6BEG[1] Tile_X2Y8_LUT4AB/W6BEG[2] Tile_X2Y8_LUT4AB/W6BEG[3] Tile_X2Y8_LUT4AB/W6BEG[4]
+ Tile_X2Y8_LUT4AB/W6BEG[5] Tile_X2Y8_LUT4AB/W6BEG[6] Tile_X2Y8_LUT4AB/W6BEG[7] Tile_X2Y8_LUT4AB/W6BEG[8]
+ Tile_X2Y8_LUT4AB/W6BEG[9] Tile_X3Y8_LUT4AB/W6BEG[0] Tile_X3Y8_LUT4AB/W6BEG[10] Tile_X3Y8_LUT4AB/W6BEG[11]
+ Tile_X3Y8_LUT4AB/W6BEG[1] Tile_X3Y8_LUT4AB/W6BEG[2] Tile_X3Y8_LUT4AB/W6BEG[3] Tile_X3Y8_LUT4AB/W6BEG[4]
+ Tile_X3Y8_LUT4AB/W6BEG[5] Tile_X3Y8_LUT4AB/W6BEG[6] Tile_X3Y8_LUT4AB/W6BEG[7] Tile_X3Y8_LUT4AB/W6BEG[8]
+ Tile_X3Y8_LUT4AB/W6BEG[9] Tile_X2Y8_LUT4AB/WW4BEG[0] Tile_X2Y8_LUT4AB/WW4BEG[10]
+ Tile_X2Y8_LUT4AB/WW4BEG[11] Tile_X2Y8_LUT4AB/WW4BEG[12] Tile_X2Y8_LUT4AB/WW4BEG[13]
+ Tile_X2Y8_LUT4AB/WW4BEG[14] Tile_X2Y8_LUT4AB/WW4BEG[15] Tile_X2Y8_LUT4AB/WW4BEG[1]
+ Tile_X2Y8_LUT4AB/WW4BEG[2] Tile_X2Y8_LUT4AB/WW4BEG[3] Tile_X2Y8_LUT4AB/WW4BEG[4]
+ Tile_X2Y8_LUT4AB/WW4BEG[5] Tile_X2Y8_LUT4AB/WW4BEG[6] Tile_X2Y8_LUT4AB/WW4BEG[7]
+ Tile_X2Y8_LUT4AB/WW4BEG[8] Tile_X2Y8_LUT4AB/WW4BEG[9] Tile_X3Y8_LUT4AB/WW4BEG[0]
+ Tile_X3Y8_LUT4AB/WW4BEG[10] Tile_X3Y8_LUT4AB/WW4BEG[11] Tile_X3Y8_LUT4AB/WW4BEG[12]
+ Tile_X3Y8_LUT4AB/WW4BEG[13] Tile_X3Y8_LUT4AB/WW4BEG[14] Tile_X3Y8_LUT4AB/WW4BEG[15]
+ Tile_X3Y8_LUT4AB/WW4BEG[1] Tile_X3Y8_LUT4AB/WW4BEG[2] Tile_X3Y8_LUT4AB/WW4BEG[3]
+ Tile_X3Y8_LUT4AB/WW4BEG[4] Tile_X3Y8_LUT4AB/WW4BEG[5] Tile_X3Y8_LUT4AB/WW4BEG[6]
+ Tile_X3Y8_LUT4AB/WW4BEG[7] Tile_X3Y8_LUT4AB/WW4BEG[8] Tile_X3Y8_LUT4AB/WW4BEG[9]
+ LUT4AB
XTile_X2Y0_N_IO4 Tile_X2Y0_A_I_top Tile_X2Y0_A_O_top Tile_X2Y0_A_T_top Tile_X2Y0_B_I_top
+ Tile_X2Y0_B_O_top Tile_X2Y0_B_T_top Tile_X2Y0_C_I_top Tile_X2Y0_C_O_top Tile_X2Y0_C_T_top
+ Tile_X2Y0_N_IO4/Ci Tile_X2Y0_D_I_top Tile_X2Y0_D_O_top Tile_X2Y0_D_T_top Tile_X2Y0_N_IO4/FrameData[0]
+ Tile_X2Y0_N_IO4/FrameData[10] Tile_X2Y0_N_IO4/FrameData[11] Tile_X2Y0_N_IO4/FrameData[12]
+ Tile_X2Y0_N_IO4/FrameData[13] Tile_X2Y0_N_IO4/FrameData[14] Tile_X2Y0_N_IO4/FrameData[15]
+ Tile_X2Y0_N_IO4/FrameData[16] Tile_X2Y0_N_IO4/FrameData[17] Tile_X2Y0_N_IO4/FrameData[18]
+ Tile_X2Y0_N_IO4/FrameData[19] Tile_X2Y0_N_IO4/FrameData[1] Tile_X2Y0_N_IO4/FrameData[20]
+ Tile_X2Y0_N_IO4/FrameData[21] Tile_X2Y0_N_IO4/FrameData[22] Tile_X2Y0_N_IO4/FrameData[23]
+ Tile_X2Y0_N_IO4/FrameData[24] Tile_X2Y0_N_IO4/FrameData[25] Tile_X2Y0_N_IO4/FrameData[26]
+ Tile_X2Y0_N_IO4/FrameData[27] Tile_X2Y0_N_IO4/FrameData[28] Tile_X2Y0_N_IO4/FrameData[29]
+ Tile_X2Y0_N_IO4/FrameData[2] Tile_X2Y0_N_IO4/FrameData[30] Tile_X2Y0_N_IO4/FrameData[31]
+ Tile_X2Y0_N_IO4/FrameData[3] Tile_X2Y0_N_IO4/FrameData[4] Tile_X2Y0_N_IO4/FrameData[5]
+ Tile_X2Y0_N_IO4/FrameData[6] Tile_X2Y0_N_IO4/FrameData[7] Tile_X2Y0_N_IO4/FrameData[8]
+ Tile_X2Y0_N_IO4/FrameData[9] Tile_X3Y0_N_IO4/FrameData[0] Tile_X3Y0_N_IO4/FrameData[10]
+ Tile_X3Y0_N_IO4/FrameData[11] Tile_X3Y0_N_IO4/FrameData[12] Tile_X3Y0_N_IO4/FrameData[13]
+ Tile_X3Y0_N_IO4/FrameData[14] Tile_X3Y0_N_IO4/FrameData[15] Tile_X3Y0_N_IO4/FrameData[16]
+ Tile_X3Y0_N_IO4/FrameData[17] Tile_X3Y0_N_IO4/FrameData[18] Tile_X3Y0_N_IO4/FrameData[19]
+ Tile_X3Y0_N_IO4/FrameData[1] Tile_X3Y0_N_IO4/FrameData[20] Tile_X3Y0_N_IO4/FrameData[21]
+ Tile_X3Y0_N_IO4/FrameData[22] Tile_X3Y0_N_IO4/FrameData[23] Tile_X3Y0_N_IO4/FrameData[24]
+ Tile_X3Y0_N_IO4/FrameData[25] Tile_X3Y0_N_IO4/FrameData[26] Tile_X3Y0_N_IO4/FrameData[27]
+ Tile_X3Y0_N_IO4/FrameData[28] Tile_X3Y0_N_IO4/FrameData[29] Tile_X3Y0_N_IO4/FrameData[2]
+ Tile_X3Y0_N_IO4/FrameData[30] Tile_X3Y0_N_IO4/FrameData[31] Tile_X3Y0_N_IO4/FrameData[3]
+ Tile_X3Y0_N_IO4/FrameData[4] Tile_X3Y0_N_IO4/FrameData[5] Tile_X3Y0_N_IO4/FrameData[6]
+ Tile_X3Y0_N_IO4/FrameData[7] Tile_X3Y0_N_IO4/FrameData[8] Tile_X3Y0_N_IO4/FrameData[9]
+ Tile_X2Y0_N_IO4/FrameStrobe[0] Tile_X2Y0_N_IO4/FrameStrobe[10] Tile_X2Y0_N_IO4/FrameStrobe[11]
+ Tile_X2Y0_N_IO4/FrameStrobe[12] Tile_X2Y0_N_IO4/FrameStrobe[13] Tile_X2Y0_N_IO4/FrameStrobe[14]
+ Tile_X2Y0_N_IO4/FrameStrobe[15] Tile_X2Y0_N_IO4/FrameStrobe[16] Tile_X2Y0_N_IO4/FrameStrobe[17]
+ Tile_X2Y0_N_IO4/FrameStrobe[18] Tile_X2Y0_N_IO4/FrameStrobe[19] Tile_X2Y0_N_IO4/FrameStrobe[1]
+ Tile_X2Y0_N_IO4/FrameStrobe[2] Tile_X2Y0_N_IO4/FrameStrobe[3] Tile_X2Y0_N_IO4/FrameStrobe[4]
+ Tile_X2Y0_N_IO4/FrameStrobe[5] Tile_X2Y0_N_IO4/FrameStrobe[6] Tile_X2Y0_N_IO4/FrameStrobe[7]
+ Tile_X2Y0_N_IO4/FrameStrobe[8] Tile_X2Y0_N_IO4/FrameStrobe[9] Tile_X2Y0_N_IO4/FrameStrobe_O[0]
+ Tile_X2Y0_N_IO4/FrameStrobe_O[10] Tile_X2Y0_N_IO4/FrameStrobe_O[11] Tile_X2Y0_N_IO4/FrameStrobe_O[12]
+ Tile_X2Y0_N_IO4/FrameStrobe_O[13] Tile_X2Y0_N_IO4/FrameStrobe_O[14] Tile_X2Y0_N_IO4/FrameStrobe_O[15]
+ Tile_X2Y0_N_IO4/FrameStrobe_O[16] Tile_X2Y0_N_IO4/FrameStrobe_O[17] Tile_X2Y0_N_IO4/FrameStrobe_O[18]
+ Tile_X2Y0_N_IO4/FrameStrobe_O[19] Tile_X2Y0_N_IO4/FrameStrobe_O[1] Tile_X2Y0_N_IO4/FrameStrobe_O[2]
+ Tile_X2Y0_N_IO4/FrameStrobe_O[3] Tile_X2Y0_N_IO4/FrameStrobe_O[4] Tile_X2Y0_N_IO4/FrameStrobe_O[5]
+ Tile_X2Y0_N_IO4/FrameStrobe_O[6] Tile_X2Y0_N_IO4/FrameStrobe_O[7] Tile_X2Y0_N_IO4/FrameStrobe_O[8]
+ Tile_X2Y0_N_IO4/FrameStrobe_O[9] Tile_X2Y0_N_IO4/N1END[0] Tile_X2Y0_N_IO4/N1END[1]
+ Tile_X2Y0_N_IO4/N1END[2] Tile_X2Y0_N_IO4/N1END[3] Tile_X2Y0_N_IO4/N2END[0] Tile_X2Y0_N_IO4/N2END[1]
+ Tile_X2Y0_N_IO4/N2END[2] Tile_X2Y0_N_IO4/N2END[3] Tile_X2Y0_N_IO4/N2END[4] Tile_X2Y0_N_IO4/N2END[5]
+ Tile_X2Y0_N_IO4/N2END[6] Tile_X2Y0_N_IO4/N2END[7] Tile_X2Y0_N_IO4/N2MID[0] Tile_X2Y0_N_IO4/N2MID[1]
+ Tile_X2Y0_N_IO4/N2MID[2] Tile_X2Y0_N_IO4/N2MID[3] Tile_X2Y0_N_IO4/N2MID[4] Tile_X2Y0_N_IO4/N2MID[5]
+ Tile_X2Y0_N_IO4/N2MID[6] Tile_X2Y0_N_IO4/N2MID[7] Tile_X2Y0_N_IO4/N4END[0] Tile_X2Y0_N_IO4/N4END[10]
+ Tile_X2Y0_N_IO4/N4END[11] Tile_X2Y0_N_IO4/N4END[12] Tile_X2Y0_N_IO4/N4END[13] Tile_X2Y0_N_IO4/N4END[14]
+ Tile_X2Y0_N_IO4/N4END[15] Tile_X2Y0_N_IO4/N4END[1] Tile_X2Y0_N_IO4/N4END[2] Tile_X2Y0_N_IO4/N4END[3]
+ Tile_X2Y0_N_IO4/N4END[4] Tile_X2Y0_N_IO4/N4END[5] Tile_X2Y0_N_IO4/N4END[6] Tile_X2Y0_N_IO4/N4END[7]
+ Tile_X2Y0_N_IO4/N4END[8] Tile_X2Y0_N_IO4/N4END[9] Tile_X2Y0_N_IO4/NN4END[0] Tile_X2Y0_N_IO4/NN4END[10]
+ Tile_X2Y0_N_IO4/NN4END[11] Tile_X2Y0_N_IO4/NN4END[12] Tile_X2Y0_N_IO4/NN4END[13]
+ Tile_X2Y0_N_IO4/NN4END[14] Tile_X2Y0_N_IO4/NN4END[15] Tile_X2Y0_N_IO4/NN4END[1]
+ Tile_X2Y0_N_IO4/NN4END[2] Tile_X2Y0_N_IO4/NN4END[3] Tile_X2Y0_N_IO4/NN4END[4] Tile_X2Y0_N_IO4/NN4END[5]
+ Tile_X2Y0_N_IO4/NN4END[6] Tile_X2Y0_N_IO4/NN4END[7] Tile_X2Y0_N_IO4/NN4END[8] Tile_X2Y0_N_IO4/NN4END[9]
+ Tile_X2Y0_N_IO4/S1BEG[0] Tile_X2Y0_N_IO4/S1BEG[1] Tile_X2Y0_N_IO4/S1BEG[2] Tile_X2Y0_N_IO4/S1BEG[3]
+ Tile_X2Y0_N_IO4/S2BEG[0] Tile_X2Y0_N_IO4/S2BEG[1] Tile_X2Y0_N_IO4/S2BEG[2] Tile_X2Y0_N_IO4/S2BEG[3]
+ Tile_X2Y0_N_IO4/S2BEG[4] Tile_X2Y0_N_IO4/S2BEG[5] Tile_X2Y0_N_IO4/S2BEG[6] Tile_X2Y0_N_IO4/S2BEG[7]
+ Tile_X2Y1_LUT4AB/S2END[0] Tile_X2Y1_LUT4AB/S2END[1] Tile_X2Y1_LUT4AB/S2END[2] Tile_X2Y1_LUT4AB/S2END[3]
+ Tile_X2Y1_LUT4AB/S2END[4] Tile_X2Y1_LUT4AB/S2END[5] Tile_X2Y1_LUT4AB/S2END[6] Tile_X2Y1_LUT4AB/S2END[7]
+ Tile_X2Y0_N_IO4/S4BEG[0] Tile_X2Y0_N_IO4/S4BEG[10] Tile_X2Y0_N_IO4/S4BEG[11] Tile_X2Y0_N_IO4/S4BEG[12]
+ Tile_X2Y0_N_IO4/S4BEG[13] Tile_X2Y0_N_IO4/S4BEG[14] Tile_X2Y0_N_IO4/S4BEG[15] Tile_X2Y0_N_IO4/S4BEG[1]
+ Tile_X2Y0_N_IO4/S4BEG[2] Tile_X2Y0_N_IO4/S4BEG[3] Tile_X2Y0_N_IO4/S4BEG[4] Tile_X2Y0_N_IO4/S4BEG[5]
+ Tile_X2Y0_N_IO4/S4BEG[6] Tile_X2Y0_N_IO4/S4BEG[7] Tile_X2Y0_N_IO4/S4BEG[8] Tile_X2Y0_N_IO4/S4BEG[9]
+ Tile_X2Y0_N_IO4/SS4BEG[0] Tile_X2Y0_N_IO4/SS4BEG[10] Tile_X2Y0_N_IO4/SS4BEG[11]
+ Tile_X2Y0_N_IO4/SS4BEG[12] Tile_X2Y0_N_IO4/SS4BEG[13] Tile_X2Y0_N_IO4/SS4BEG[14]
+ Tile_X2Y0_N_IO4/SS4BEG[15] Tile_X2Y0_N_IO4/SS4BEG[1] Tile_X2Y0_N_IO4/SS4BEG[2] Tile_X2Y0_N_IO4/SS4BEG[3]
+ Tile_X2Y0_N_IO4/SS4BEG[4] Tile_X2Y0_N_IO4/SS4BEG[5] Tile_X2Y0_N_IO4/SS4BEG[6] Tile_X2Y0_N_IO4/SS4BEG[7]
+ Tile_X2Y0_N_IO4/SS4BEG[8] Tile_X2Y0_N_IO4/SS4BEG[9] Tile_X2Y0_N_IO4/UserCLK Tile_X2Y0_N_IO4/UserCLKo
+ VGND VPWR N_IO4
XTile_X1Y1_LUT4AB Tile_X1Y2_LUT4AB/Co Tile_X1Y0_N_IO4/Ci Tile_X2Y1_LUT4AB/E1END[0]
+ Tile_X2Y1_LUT4AB/E1END[1] Tile_X2Y1_LUT4AB/E1END[2] Tile_X2Y1_LUT4AB/E1END[3] Tile_X1Y1_LUT4AB/E1END[0]
+ Tile_X1Y1_LUT4AB/E1END[1] Tile_X1Y1_LUT4AB/E1END[2] Tile_X1Y1_LUT4AB/E1END[3] Tile_X2Y1_LUT4AB/E2MID[0]
+ Tile_X2Y1_LUT4AB/E2MID[1] Tile_X2Y1_LUT4AB/E2MID[2] Tile_X2Y1_LUT4AB/E2MID[3] Tile_X2Y1_LUT4AB/E2MID[4]
+ Tile_X2Y1_LUT4AB/E2MID[5] Tile_X2Y1_LUT4AB/E2MID[6] Tile_X2Y1_LUT4AB/E2MID[7] Tile_X2Y1_LUT4AB/E2END[0]
+ Tile_X2Y1_LUT4AB/E2END[1] Tile_X2Y1_LUT4AB/E2END[2] Tile_X2Y1_LUT4AB/E2END[3] Tile_X2Y1_LUT4AB/E2END[4]
+ Tile_X2Y1_LUT4AB/E2END[5] Tile_X2Y1_LUT4AB/E2END[6] Tile_X2Y1_LUT4AB/E2END[7] Tile_X1Y1_LUT4AB/E2END[0]
+ Tile_X1Y1_LUT4AB/E2END[1] Tile_X1Y1_LUT4AB/E2END[2] Tile_X1Y1_LUT4AB/E2END[3] Tile_X1Y1_LUT4AB/E2END[4]
+ Tile_X1Y1_LUT4AB/E2END[5] Tile_X1Y1_LUT4AB/E2END[6] Tile_X1Y1_LUT4AB/E2END[7] Tile_X1Y1_LUT4AB/E2MID[0]
+ Tile_X1Y1_LUT4AB/E2MID[1] Tile_X1Y1_LUT4AB/E2MID[2] Tile_X1Y1_LUT4AB/E2MID[3] Tile_X1Y1_LUT4AB/E2MID[4]
+ Tile_X1Y1_LUT4AB/E2MID[5] Tile_X1Y1_LUT4AB/E2MID[6] Tile_X1Y1_LUT4AB/E2MID[7] Tile_X2Y1_LUT4AB/E6END[0]
+ Tile_X2Y1_LUT4AB/E6END[10] Tile_X2Y1_LUT4AB/E6END[11] Tile_X2Y1_LUT4AB/E6END[1]
+ Tile_X2Y1_LUT4AB/E6END[2] Tile_X2Y1_LUT4AB/E6END[3] Tile_X2Y1_LUT4AB/E6END[4] Tile_X2Y1_LUT4AB/E6END[5]
+ Tile_X2Y1_LUT4AB/E6END[6] Tile_X2Y1_LUT4AB/E6END[7] Tile_X2Y1_LUT4AB/E6END[8] Tile_X2Y1_LUT4AB/E6END[9]
+ Tile_X1Y1_LUT4AB/E6END[0] Tile_X1Y1_LUT4AB/E6END[10] Tile_X1Y1_LUT4AB/E6END[11]
+ Tile_X1Y1_LUT4AB/E6END[1] Tile_X1Y1_LUT4AB/E6END[2] Tile_X1Y1_LUT4AB/E6END[3] Tile_X1Y1_LUT4AB/E6END[4]
+ Tile_X1Y1_LUT4AB/E6END[5] Tile_X1Y1_LUT4AB/E6END[6] Tile_X1Y1_LUT4AB/E6END[7] Tile_X1Y1_LUT4AB/E6END[8]
+ Tile_X1Y1_LUT4AB/E6END[9] Tile_X2Y1_LUT4AB/EE4END[0] Tile_X2Y1_LUT4AB/EE4END[10]
+ Tile_X2Y1_LUT4AB/EE4END[11] Tile_X2Y1_LUT4AB/EE4END[12] Tile_X2Y1_LUT4AB/EE4END[13]
+ Tile_X2Y1_LUT4AB/EE4END[14] Tile_X2Y1_LUT4AB/EE4END[15] Tile_X2Y1_LUT4AB/EE4END[1]
+ Tile_X2Y1_LUT4AB/EE4END[2] Tile_X2Y1_LUT4AB/EE4END[3] Tile_X2Y1_LUT4AB/EE4END[4]
+ Tile_X2Y1_LUT4AB/EE4END[5] Tile_X2Y1_LUT4AB/EE4END[6] Tile_X2Y1_LUT4AB/EE4END[7]
+ Tile_X2Y1_LUT4AB/EE4END[8] Tile_X2Y1_LUT4AB/EE4END[9] Tile_X1Y1_LUT4AB/EE4END[0]
+ Tile_X1Y1_LUT4AB/EE4END[10] Tile_X1Y1_LUT4AB/EE4END[11] Tile_X1Y1_LUT4AB/EE4END[12]
+ Tile_X1Y1_LUT4AB/EE4END[13] Tile_X1Y1_LUT4AB/EE4END[14] Tile_X1Y1_LUT4AB/EE4END[15]
+ Tile_X1Y1_LUT4AB/EE4END[1] Tile_X1Y1_LUT4AB/EE4END[2] Tile_X1Y1_LUT4AB/EE4END[3]
+ Tile_X1Y1_LUT4AB/EE4END[4] Tile_X1Y1_LUT4AB/EE4END[5] Tile_X1Y1_LUT4AB/EE4END[6]
+ Tile_X1Y1_LUT4AB/EE4END[7] Tile_X1Y1_LUT4AB/EE4END[8] Tile_X1Y1_LUT4AB/EE4END[9]
+ Tile_X1Y1_LUT4AB/FrameData[0] Tile_X1Y1_LUT4AB/FrameData[10] Tile_X1Y1_LUT4AB/FrameData[11]
+ Tile_X1Y1_LUT4AB/FrameData[12] Tile_X1Y1_LUT4AB/FrameData[13] Tile_X1Y1_LUT4AB/FrameData[14]
+ Tile_X1Y1_LUT4AB/FrameData[15] Tile_X1Y1_LUT4AB/FrameData[16] Tile_X1Y1_LUT4AB/FrameData[17]
+ Tile_X1Y1_LUT4AB/FrameData[18] Tile_X1Y1_LUT4AB/FrameData[19] Tile_X1Y1_LUT4AB/FrameData[1]
+ Tile_X1Y1_LUT4AB/FrameData[20] Tile_X1Y1_LUT4AB/FrameData[21] Tile_X1Y1_LUT4AB/FrameData[22]
+ Tile_X1Y1_LUT4AB/FrameData[23] Tile_X1Y1_LUT4AB/FrameData[24] Tile_X1Y1_LUT4AB/FrameData[25]
+ Tile_X1Y1_LUT4AB/FrameData[26] Tile_X1Y1_LUT4AB/FrameData[27] Tile_X1Y1_LUT4AB/FrameData[28]
+ Tile_X1Y1_LUT4AB/FrameData[29] Tile_X1Y1_LUT4AB/FrameData[2] Tile_X1Y1_LUT4AB/FrameData[30]
+ Tile_X1Y1_LUT4AB/FrameData[31] Tile_X1Y1_LUT4AB/FrameData[3] Tile_X1Y1_LUT4AB/FrameData[4]
+ Tile_X1Y1_LUT4AB/FrameData[5] Tile_X1Y1_LUT4AB/FrameData[6] Tile_X1Y1_LUT4AB/FrameData[7]
+ Tile_X1Y1_LUT4AB/FrameData[8] Tile_X1Y1_LUT4AB/FrameData[9] Tile_X2Y1_LUT4AB/FrameData[0]
+ Tile_X2Y1_LUT4AB/FrameData[10] Tile_X2Y1_LUT4AB/FrameData[11] Tile_X2Y1_LUT4AB/FrameData[12]
+ Tile_X2Y1_LUT4AB/FrameData[13] Tile_X2Y1_LUT4AB/FrameData[14] Tile_X2Y1_LUT4AB/FrameData[15]
+ Tile_X2Y1_LUT4AB/FrameData[16] Tile_X2Y1_LUT4AB/FrameData[17] Tile_X2Y1_LUT4AB/FrameData[18]
+ Tile_X2Y1_LUT4AB/FrameData[19] Tile_X2Y1_LUT4AB/FrameData[1] Tile_X2Y1_LUT4AB/FrameData[20]
+ Tile_X2Y1_LUT4AB/FrameData[21] Tile_X2Y1_LUT4AB/FrameData[22] Tile_X2Y1_LUT4AB/FrameData[23]
+ Tile_X2Y1_LUT4AB/FrameData[24] Tile_X2Y1_LUT4AB/FrameData[25] Tile_X2Y1_LUT4AB/FrameData[26]
+ Tile_X2Y1_LUT4AB/FrameData[27] Tile_X2Y1_LUT4AB/FrameData[28] Tile_X2Y1_LUT4AB/FrameData[29]
+ Tile_X2Y1_LUT4AB/FrameData[2] Tile_X2Y1_LUT4AB/FrameData[30] Tile_X2Y1_LUT4AB/FrameData[31]
+ Tile_X2Y1_LUT4AB/FrameData[3] Tile_X2Y1_LUT4AB/FrameData[4] Tile_X2Y1_LUT4AB/FrameData[5]
+ Tile_X2Y1_LUT4AB/FrameData[6] Tile_X2Y1_LUT4AB/FrameData[7] Tile_X2Y1_LUT4AB/FrameData[8]
+ Tile_X2Y1_LUT4AB/FrameData[9] Tile_X1Y1_LUT4AB/FrameStrobe[0] Tile_X1Y1_LUT4AB/FrameStrobe[10]
+ Tile_X1Y1_LUT4AB/FrameStrobe[11] Tile_X1Y1_LUT4AB/FrameStrobe[12] Tile_X1Y1_LUT4AB/FrameStrobe[13]
+ Tile_X1Y1_LUT4AB/FrameStrobe[14] Tile_X1Y1_LUT4AB/FrameStrobe[15] Tile_X1Y1_LUT4AB/FrameStrobe[16]
+ Tile_X1Y1_LUT4AB/FrameStrobe[17] Tile_X1Y1_LUT4AB/FrameStrobe[18] Tile_X1Y1_LUT4AB/FrameStrobe[19]
+ Tile_X1Y1_LUT4AB/FrameStrobe[1] Tile_X1Y1_LUT4AB/FrameStrobe[2] Tile_X1Y1_LUT4AB/FrameStrobe[3]
+ Tile_X1Y1_LUT4AB/FrameStrobe[4] Tile_X1Y1_LUT4AB/FrameStrobe[5] Tile_X1Y1_LUT4AB/FrameStrobe[6]
+ Tile_X1Y1_LUT4AB/FrameStrobe[7] Tile_X1Y1_LUT4AB/FrameStrobe[8] Tile_X1Y1_LUT4AB/FrameStrobe[9]
+ Tile_X1Y0_N_IO4/FrameStrobe[0] Tile_X1Y0_N_IO4/FrameStrobe[10] Tile_X1Y0_N_IO4/FrameStrobe[11]
+ Tile_X1Y0_N_IO4/FrameStrobe[12] Tile_X1Y0_N_IO4/FrameStrobe[13] Tile_X1Y0_N_IO4/FrameStrobe[14]
+ Tile_X1Y0_N_IO4/FrameStrobe[15] Tile_X1Y0_N_IO4/FrameStrobe[16] Tile_X1Y0_N_IO4/FrameStrobe[17]
+ Tile_X1Y0_N_IO4/FrameStrobe[18] Tile_X1Y0_N_IO4/FrameStrobe[19] Tile_X1Y0_N_IO4/FrameStrobe[1]
+ Tile_X1Y0_N_IO4/FrameStrobe[2] Tile_X1Y0_N_IO4/FrameStrobe[3] Tile_X1Y0_N_IO4/FrameStrobe[4]
+ Tile_X1Y0_N_IO4/FrameStrobe[5] Tile_X1Y0_N_IO4/FrameStrobe[6] Tile_X1Y0_N_IO4/FrameStrobe[7]
+ Tile_X1Y0_N_IO4/FrameStrobe[8] Tile_X1Y0_N_IO4/FrameStrobe[9] Tile_X1Y0_N_IO4/N1END[0]
+ Tile_X1Y0_N_IO4/N1END[1] Tile_X1Y0_N_IO4/N1END[2] Tile_X1Y0_N_IO4/N1END[3] Tile_X1Y2_LUT4AB/N1BEG[0]
+ Tile_X1Y2_LUT4AB/N1BEG[1] Tile_X1Y2_LUT4AB/N1BEG[2] Tile_X1Y2_LUT4AB/N1BEG[3] Tile_X1Y0_N_IO4/N2MID[0]
+ Tile_X1Y0_N_IO4/N2MID[1] Tile_X1Y0_N_IO4/N2MID[2] Tile_X1Y0_N_IO4/N2MID[3] Tile_X1Y0_N_IO4/N2MID[4]
+ Tile_X1Y0_N_IO4/N2MID[5] Tile_X1Y0_N_IO4/N2MID[6] Tile_X1Y0_N_IO4/N2MID[7] Tile_X1Y0_N_IO4/N2END[0]
+ Tile_X1Y0_N_IO4/N2END[1] Tile_X1Y0_N_IO4/N2END[2] Tile_X1Y0_N_IO4/N2END[3] Tile_X1Y0_N_IO4/N2END[4]
+ Tile_X1Y0_N_IO4/N2END[5] Tile_X1Y0_N_IO4/N2END[6] Tile_X1Y0_N_IO4/N2END[7] Tile_X1Y1_LUT4AB/N2END[0]
+ Tile_X1Y1_LUT4AB/N2END[1] Tile_X1Y1_LUT4AB/N2END[2] Tile_X1Y1_LUT4AB/N2END[3] Tile_X1Y1_LUT4AB/N2END[4]
+ Tile_X1Y1_LUT4AB/N2END[5] Tile_X1Y1_LUT4AB/N2END[6] Tile_X1Y1_LUT4AB/N2END[7] Tile_X1Y2_LUT4AB/N2BEG[0]
+ Tile_X1Y2_LUT4AB/N2BEG[1] Tile_X1Y2_LUT4AB/N2BEG[2] Tile_X1Y2_LUT4AB/N2BEG[3] Tile_X1Y2_LUT4AB/N2BEG[4]
+ Tile_X1Y2_LUT4AB/N2BEG[5] Tile_X1Y2_LUT4AB/N2BEG[6] Tile_X1Y2_LUT4AB/N2BEG[7] Tile_X1Y0_N_IO4/N4END[0]
+ Tile_X1Y0_N_IO4/N4END[10] Tile_X1Y0_N_IO4/N4END[11] Tile_X1Y0_N_IO4/N4END[12] Tile_X1Y0_N_IO4/N4END[13]
+ Tile_X1Y0_N_IO4/N4END[14] Tile_X1Y0_N_IO4/N4END[15] Tile_X1Y0_N_IO4/N4END[1] Tile_X1Y0_N_IO4/N4END[2]
+ Tile_X1Y0_N_IO4/N4END[3] Tile_X1Y0_N_IO4/N4END[4] Tile_X1Y0_N_IO4/N4END[5] Tile_X1Y0_N_IO4/N4END[6]
+ Tile_X1Y0_N_IO4/N4END[7] Tile_X1Y0_N_IO4/N4END[8] Tile_X1Y0_N_IO4/N4END[9] Tile_X1Y2_LUT4AB/N4BEG[0]
+ Tile_X1Y2_LUT4AB/N4BEG[10] Tile_X1Y2_LUT4AB/N4BEG[11] Tile_X1Y2_LUT4AB/N4BEG[12]
+ Tile_X1Y2_LUT4AB/N4BEG[13] Tile_X1Y2_LUT4AB/N4BEG[14] Tile_X1Y2_LUT4AB/N4BEG[15]
+ Tile_X1Y2_LUT4AB/N4BEG[1] Tile_X1Y2_LUT4AB/N4BEG[2] Tile_X1Y2_LUT4AB/N4BEG[3] Tile_X1Y2_LUT4AB/N4BEG[4]
+ Tile_X1Y2_LUT4AB/N4BEG[5] Tile_X1Y2_LUT4AB/N4BEG[6] Tile_X1Y2_LUT4AB/N4BEG[7] Tile_X1Y2_LUT4AB/N4BEG[8]
+ Tile_X1Y2_LUT4AB/N4BEG[9] Tile_X1Y0_N_IO4/NN4END[0] Tile_X1Y0_N_IO4/NN4END[10] Tile_X1Y0_N_IO4/NN4END[11]
+ Tile_X1Y0_N_IO4/NN4END[12] Tile_X1Y0_N_IO4/NN4END[13] Tile_X1Y0_N_IO4/NN4END[14]
+ Tile_X1Y0_N_IO4/NN4END[15] Tile_X1Y0_N_IO4/NN4END[1] Tile_X1Y0_N_IO4/NN4END[2] Tile_X1Y0_N_IO4/NN4END[3]
+ Tile_X1Y0_N_IO4/NN4END[4] Tile_X1Y0_N_IO4/NN4END[5] Tile_X1Y0_N_IO4/NN4END[6] Tile_X1Y0_N_IO4/NN4END[7]
+ Tile_X1Y0_N_IO4/NN4END[8] Tile_X1Y0_N_IO4/NN4END[9] Tile_X1Y2_LUT4AB/NN4BEG[0] Tile_X1Y2_LUT4AB/NN4BEG[10]
+ Tile_X1Y2_LUT4AB/NN4BEG[11] Tile_X1Y2_LUT4AB/NN4BEG[12] Tile_X1Y2_LUT4AB/NN4BEG[13]
+ Tile_X1Y2_LUT4AB/NN4BEG[14] Tile_X1Y2_LUT4AB/NN4BEG[15] Tile_X1Y2_LUT4AB/NN4BEG[1]
+ Tile_X1Y2_LUT4AB/NN4BEG[2] Tile_X1Y2_LUT4AB/NN4BEG[3] Tile_X1Y2_LUT4AB/NN4BEG[4]
+ Tile_X1Y2_LUT4AB/NN4BEG[5] Tile_X1Y2_LUT4AB/NN4BEG[6] Tile_X1Y2_LUT4AB/NN4BEG[7]
+ Tile_X1Y2_LUT4AB/NN4BEG[8] Tile_X1Y2_LUT4AB/NN4BEG[9] Tile_X1Y2_LUT4AB/S1END[0]
+ Tile_X1Y2_LUT4AB/S1END[1] Tile_X1Y2_LUT4AB/S1END[2] Tile_X1Y2_LUT4AB/S1END[3] Tile_X1Y0_N_IO4/S1BEG[0]
+ Tile_X1Y0_N_IO4/S1BEG[1] Tile_X1Y0_N_IO4/S1BEG[2] Tile_X1Y0_N_IO4/S1BEG[3] Tile_X1Y2_LUT4AB/S2MID[0]
+ Tile_X1Y2_LUT4AB/S2MID[1] Tile_X1Y2_LUT4AB/S2MID[2] Tile_X1Y2_LUT4AB/S2MID[3] Tile_X1Y2_LUT4AB/S2MID[4]
+ Tile_X1Y2_LUT4AB/S2MID[5] Tile_X1Y2_LUT4AB/S2MID[6] Tile_X1Y2_LUT4AB/S2MID[7] Tile_X1Y2_LUT4AB/S2END[0]
+ Tile_X1Y2_LUT4AB/S2END[1] Tile_X1Y2_LUT4AB/S2END[2] Tile_X1Y2_LUT4AB/S2END[3] Tile_X1Y2_LUT4AB/S2END[4]
+ Tile_X1Y2_LUT4AB/S2END[5] Tile_X1Y2_LUT4AB/S2END[6] Tile_X1Y2_LUT4AB/S2END[7] Tile_X1Y1_LUT4AB/S2END[0]
+ Tile_X1Y1_LUT4AB/S2END[1] Tile_X1Y1_LUT4AB/S2END[2] Tile_X1Y1_LUT4AB/S2END[3] Tile_X1Y1_LUT4AB/S2END[4]
+ Tile_X1Y1_LUT4AB/S2END[5] Tile_X1Y1_LUT4AB/S2END[6] Tile_X1Y1_LUT4AB/S2END[7] Tile_X1Y0_N_IO4/S2BEG[0]
+ Tile_X1Y0_N_IO4/S2BEG[1] Tile_X1Y0_N_IO4/S2BEG[2] Tile_X1Y0_N_IO4/S2BEG[3] Tile_X1Y0_N_IO4/S2BEG[4]
+ Tile_X1Y0_N_IO4/S2BEG[5] Tile_X1Y0_N_IO4/S2BEG[6] Tile_X1Y0_N_IO4/S2BEG[7] Tile_X1Y2_LUT4AB/S4END[0]
+ Tile_X1Y2_LUT4AB/S4END[10] Tile_X1Y2_LUT4AB/S4END[11] Tile_X1Y2_LUT4AB/S4END[12]
+ Tile_X1Y2_LUT4AB/S4END[13] Tile_X1Y2_LUT4AB/S4END[14] Tile_X1Y2_LUT4AB/S4END[15]
+ Tile_X1Y2_LUT4AB/S4END[1] Tile_X1Y2_LUT4AB/S4END[2] Tile_X1Y2_LUT4AB/S4END[3] Tile_X1Y2_LUT4AB/S4END[4]
+ Tile_X1Y2_LUT4AB/S4END[5] Tile_X1Y2_LUT4AB/S4END[6] Tile_X1Y2_LUT4AB/S4END[7] Tile_X1Y2_LUT4AB/S4END[8]
+ Tile_X1Y2_LUT4AB/S4END[9] Tile_X1Y0_N_IO4/S4BEG[0] Tile_X1Y0_N_IO4/S4BEG[10] Tile_X1Y0_N_IO4/S4BEG[11]
+ Tile_X1Y0_N_IO4/S4BEG[12] Tile_X1Y0_N_IO4/S4BEG[13] Tile_X1Y0_N_IO4/S4BEG[14] Tile_X1Y0_N_IO4/S4BEG[15]
+ Tile_X1Y0_N_IO4/S4BEG[1] Tile_X1Y0_N_IO4/S4BEG[2] Tile_X1Y0_N_IO4/S4BEG[3] Tile_X1Y0_N_IO4/S4BEG[4]
+ Tile_X1Y0_N_IO4/S4BEG[5] Tile_X1Y0_N_IO4/S4BEG[6] Tile_X1Y0_N_IO4/S4BEG[7] Tile_X1Y0_N_IO4/S4BEG[8]
+ Tile_X1Y0_N_IO4/S4BEG[9] Tile_X1Y2_LUT4AB/SS4END[0] Tile_X1Y2_LUT4AB/SS4END[10]
+ Tile_X1Y2_LUT4AB/SS4END[11] Tile_X1Y2_LUT4AB/SS4END[12] Tile_X1Y2_LUT4AB/SS4END[13]
+ Tile_X1Y2_LUT4AB/SS4END[14] Tile_X1Y2_LUT4AB/SS4END[15] Tile_X1Y2_LUT4AB/SS4END[1]
+ Tile_X1Y2_LUT4AB/SS4END[2] Tile_X1Y2_LUT4AB/SS4END[3] Tile_X1Y2_LUT4AB/SS4END[4]
+ Tile_X1Y2_LUT4AB/SS4END[5] Tile_X1Y2_LUT4AB/SS4END[6] Tile_X1Y2_LUT4AB/SS4END[7]
+ Tile_X1Y2_LUT4AB/SS4END[8] Tile_X1Y2_LUT4AB/SS4END[9] Tile_X1Y0_N_IO4/SS4BEG[0]
+ Tile_X1Y0_N_IO4/SS4BEG[10] Tile_X1Y0_N_IO4/SS4BEG[11] Tile_X1Y0_N_IO4/SS4BEG[12]
+ Tile_X1Y0_N_IO4/SS4BEG[13] Tile_X1Y0_N_IO4/SS4BEG[14] Tile_X1Y0_N_IO4/SS4BEG[15]
+ Tile_X1Y0_N_IO4/SS4BEG[1] Tile_X1Y0_N_IO4/SS4BEG[2] Tile_X1Y0_N_IO4/SS4BEG[3] Tile_X1Y0_N_IO4/SS4BEG[4]
+ Tile_X1Y0_N_IO4/SS4BEG[5] Tile_X1Y0_N_IO4/SS4BEG[6] Tile_X1Y0_N_IO4/SS4BEG[7] Tile_X1Y0_N_IO4/SS4BEG[8]
+ Tile_X1Y0_N_IO4/SS4BEG[9] Tile_X1Y1_LUT4AB/UserCLK Tile_X1Y0_N_IO4/UserCLK VGND
+ VPWR Tile_X1Y1_LUT4AB/W1BEG[0] Tile_X1Y1_LUT4AB/W1BEG[1] Tile_X1Y1_LUT4AB/W1BEG[2]
+ Tile_X1Y1_LUT4AB/W1BEG[3] Tile_X2Y1_LUT4AB/W1BEG[0] Tile_X2Y1_LUT4AB/W1BEG[1] Tile_X2Y1_LUT4AB/W1BEG[2]
+ Tile_X2Y1_LUT4AB/W1BEG[3] Tile_X1Y1_LUT4AB/W2BEG[0] Tile_X1Y1_LUT4AB/W2BEG[1] Tile_X1Y1_LUT4AB/W2BEG[2]
+ Tile_X1Y1_LUT4AB/W2BEG[3] Tile_X1Y1_LUT4AB/W2BEG[4] Tile_X1Y1_LUT4AB/W2BEG[5] Tile_X1Y1_LUT4AB/W2BEG[6]
+ Tile_X1Y1_LUT4AB/W2BEG[7] Tile_X1Y1_LUT4AB/W2BEGb[0] Tile_X1Y1_LUT4AB/W2BEGb[1]
+ Tile_X1Y1_LUT4AB/W2BEGb[2] Tile_X1Y1_LUT4AB/W2BEGb[3] Tile_X1Y1_LUT4AB/W2BEGb[4]
+ Tile_X1Y1_LUT4AB/W2BEGb[5] Tile_X1Y1_LUT4AB/W2BEGb[6] Tile_X1Y1_LUT4AB/W2BEGb[7]
+ Tile_X1Y1_LUT4AB/W2END[0] Tile_X1Y1_LUT4AB/W2END[1] Tile_X1Y1_LUT4AB/W2END[2] Tile_X1Y1_LUT4AB/W2END[3]
+ Tile_X1Y1_LUT4AB/W2END[4] Tile_X1Y1_LUT4AB/W2END[5] Tile_X1Y1_LUT4AB/W2END[6] Tile_X1Y1_LUT4AB/W2END[7]
+ Tile_X2Y1_LUT4AB/W2BEG[0] Tile_X2Y1_LUT4AB/W2BEG[1] Tile_X2Y1_LUT4AB/W2BEG[2] Tile_X2Y1_LUT4AB/W2BEG[3]
+ Tile_X2Y1_LUT4AB/W2BEG[4] Tile_X2Y1_LUT4AB/W2BEG[5] Tile_X2Y1_LUT4AB/W2BEG[6] Tile_X2Y1_LUT4AB/W2BEG[7]
+ Tile_X1Y1_LUT4AB/W6BEG[0] Tile_X1Y1_LUT4AB/W6BEG[10] Tile_X1Y1_LUT4AB/W6BEG[11]
+ Tile_X1Y1_LUT4AB/W6BEG[1] Tile_X1Y1_LUT4AB/W6BEG[2] Tile_X1Y1_LUT4AB/W6BEG[3] Tile_X1Y1_LUT4AB/W6BEG[4]
+ Tile_X1Y1_LUT4AB/W6BEG[5] Tile_X1Y1_LUT4AB/W6BEG[6] Tile_X1Y1_LUT4AB/W6BEG[7] Tile_X1Y1_LUT4AB/W6BEG[8]
+ Tile_X1Y1_LUT4AB/W6BEG[9] Tile_X2Y1_LUT4AB/W6BEG[0] Tile_X2Y1_LUT4AB/W6BEG[10] Tile_X2Y1_LUT4AB/W6BEG[11]
+ Tile_X2Y1_LUT4AB/W6BEG[1] Tile_X2Y1_LUT4AB/W6BEG[2] Tile_X2Y1_LUT4AB/W6BEG[3] Tile_X2Y1_LUT4AB/W6BEG[4]
+ Tile_X2Y1_LUT4AB/W6BEG[5] Tile_X2Y1_LUT4AB/W6BEG[6] Tile_X2Y1_LUT4AB/W6BEG[7] Tile_X2Y1_LUT4AB/W6BEG[8]
+ Tile_X2Y1_LUT4AB/W6BEG[9] Tile_X1Y1_LUT4AB/WW4BEG[0] Tile_X1Y1_LUT4AB/WW4BEG[10]
+ Tile_X1Y1_LUT4AB/WW4BEG[11] Tile_X1Y1_LUT4AB/WW4BEG[12] Tile_X1Y1_LUT4AB/WW4BEG[13]
+ Tile_X1Y1_LUT4AB/WW4BEG[14] Tile_X1Y1_LUT4AB/WW4BEG[15] Tile_X1Y1_LUT4AB/WW4BEG[1]
+ Tile_X1Y1_LUT4AB/WW4BEG[2] Tile_X1Y1_LUT4AB/WW4BEG[3] Tile_X1Y1_LUT4AB/WW4BEG[4]
+ Tile_X1Y1_LUT4AB/WW4BEG[5] Tile_X1Y1_LUT4AB/WW4BEG[6] Tile_X1Y1_LUT4AB/WW4BEG[7]
+ Tile_X1Y1_LUT4AB/WW4BEG[8] Tile_X1Y1_LUT4AB/WW4BEG[9] Tile_X2Y1_LUT4AB/WW4BEG[0]
+ Tile_X2Y1_LUT4AB/WW4BEG[10] Tile_X2Y1_LUT4AB/WW4BEG[11] Tile_X2Y1_LUT4AB/WW4BEG[12]
+ Tile_X2Y1_LUT4AB/WW4BEG[13] Tile_X2Y1_LUT4AB/WW4BEG[14] Tile_X2Y1_LUT4AB/WW4BEG[15]
+ Tile_X2Y1_LUT4AB/WW4BEG[1] Tile_X2Y1_LUT4AB/WW4BEG[2] Tile_X2Y1_LUT4AB/WW4BEG[3]
+ Tile_X2Y1_LUT4AB/WW4BEG[4] Tile_X2Y1_LUT4AB/WW4BEG[5] Tile_X2Y1_LUT4AB/WW4BEG[6]
+ Tile_X2Y1_LUT4AB/WW4BEG[7] Tile_X2Y1_LUT4AB/WW4BEG[8] Tile_X2Y1_LUT4AB/WW4BEG[9]
+ LUT4AB
XTile_X5Y3_E_TT_IF Tile_X5Y3_CLK_TT_PROJECT Tile_X4Y3_LUT4AB/E1BEG[0] Tile_X4Y3_LUT4AB/E1BEG[1]
+ Tile_X4Y3_LUT4AB/E1BEG[2] Tile_X4Y3_LUT4AB/E1BEG[3] Tile_X5Y3_E_TT_IF/E2END[0] Tile_X5Y3_E_TT_IF/E2END[1]
+ Tile_X5Y3_E_TT_IF/E2END[2] Tile_X5Y3_E_TT_IF/E2END[3] Tile_X5Y3_E_TT_IF/E2END[4]
+ Tile_X5Y3_E_TT_IF/E2END[5] Tile_X5Y3_E_TT_IF/E2END[6] Tile_X5Y3_E_TT_IF/E2END[7]
+ Tile_X4Y3_LUT4AB/E2BEG[0] Tile_X4Y3_LUT4AB/E2BEG[1] Tile_X4Y3_LUT4AB/E2BEG[2] Tile_X4Y3_LUT4AB/E2BEG[3]
+ Tile_X4Y3_LUT4AB/E2BEG[4] Tile_X4Y3_LUT4AB/E2BEG[5] Tile_X4Y3_LUT4AB/E2BEG[6] Tile_X4Y3_LUT4AB/E2BEG[7]
+ Tile_X4Y3_LUT4AB/E6BEG[0] Tile_X4Y3_LUT4AB/E6BEG[10] Tile_X4Y3_LUT4AB/E6BEG[11]
+ Tile_X4Y3_LUT4AB/E6BEG[1] Tile_X4Y3_LUT4AB/E6BEG[2] Tile_X4Y3_LUT4AB/E6BEG[3] Tile_X4Y3_LUT4AB/E6BEG[4]
+ Tile_X4Y3_LUT4AB/E6BEG[5] Tile_X4Y3_LUT4AB/E6BEG[6] Tile_X4Y3_LUT4AB/E6BEG[7] Tile_X4Y3_LUT4AB/E6BEG[8]
+ Tile_X4Y3_LUT4AB/E6BEG[9] Tile_X4Y3_LUT4AB/EE4BEG[0] Tile_X4Y3_LUT4AB/EE4BEG[10]
+ Tile_X4Y3_LUT4AB/EE4BEG[11] Tile_X4Y3_LUT4AB/EE4BEG[12] Tile_X4Y3_LUT4AB/EE4BEG[13]
+ Tile_X4Y3_LUT4AB/EE4BEG[14] Tile_X4Y3_LUT4AB/EE4BEG[15] Tile_X4Y3_LUT4AB/EE4BEG[1]
+ Tile_X4Y3_LUT4AB/EE4BEG[2] Tile_X4Y3_LUT4AB/EE4BEG[3] Tile_X4Y3_LUT4AB/EE4BEG[4]
+ Tile_X4Y3_LUT4AB/EE4BEG[5] Tile_X4Y3_LUT4AB/EE4BEG[6] Tile_X4Y3_LUT4AB/EE4BEG[7]
+ Tile_X4Y3_LUT4AB/EE4BEG[8] Tile_X4Y3_LUT4AB/EE4BEG[9] Tile_X5Y3_ENA_TT_PROJECT Tile_X5Y3_E_TT_IF/FrameData[0]
+ Tile_X5Y3_E_TT_IF/FrameData[10] Tile_X5Y3_E_TT_IF/FrameData[11] Tile_X5Y3_E_TT_IF/FrameData[12]
+ Tile_X5Y3_E_TT_IF/FrameData[13] Tile_X5Y3_E_TT_IF/FrameData[14] Tile_X5Y3_E_TT_IF/FrameData[15]
+ Tile_X5Y3_E_TT_IF/FrameData[16] Tile_X5Y3_E_TT_IF/FrameData[17] Tile_X5Y3_E_TT_IF/FrameData[18]
+ Tile_X5Y3_E_TT_IF/FrameData[19] Tile_X5Y3_E_TT_IF/FrameData[1] Tile_X5Y3_E_TT_IF/FrameData[20]
+ Tile_X5Y3_E_TT_IF/FrameData[21] Tile_X5Y3_E_TT_IF/FrameData[22] Tile_X5Y3_E_TT_IF/FrameData[23]
+ Tile_X5Y3_E_TT_IF/FrameData[24] Tile_X5Y3_E_TT_IF/FrameData[25] Tile_X5Y3_E_TT_IF/FrameData[26]
+ Tile_X5Y3_E_TT_IF/FrameData[27] Tile_X5Y3_E_TT_IF/FrameData[28] Tile_X5Y3_E_TT_IF/FrameData[29]
+ Tile_X5Y3_E_TT_IF/FrameData[2] Tile_X5Y3_E_TT_IF/FrameData[30] Tile_X5Y3_E_TT_IF/FrameData[31]
+ Tile_X5Y3_E_TT_IF/FrameData[3] Tile_X5Y3_E_TT_IF/FrameData[4] Tile_X5Y3_E_TT_IF/FrameData[5]
+ Tile_X5Y3_E_TT_IF/FrameData[6] Tile_X5Y3_E_TT_IF/FrameData[7] Tile_X5Y3_E_TT_IF/FrameData[8]
+ Tile_X5Y3_E_TT_IF/FrameData[9] Tile_X5Y3_E_TT_IF/FrameData_O[0] Tile_X5Y3_E_TT_IF/FrameData_O[10]
+ Tile_X5Y3_E_TT_IF/FrameData_O[11] Tile_X5Y3_E_TT_IF/FrameData_O[12] Tile_X5Y3_E_TT_IF/FrameData_O[13]
+ Tile_X5Y3_E_TT_IF/FrameData_O[14] Tile_X5Y3_E_TT_IF/FrameData_O[15] Tile_X5Y3_E_TT_IF/FrameData_O[16]
+ Tile_X5Y3_E_TT_IF/FrameData_O[17] Tile_X5Y3_E_TT_IF/FrameData_O[18] Tile_X5Y3_E_TT_IF/FrameData_O[19]
+ Tile_X5Y3_E_TT_IF/FrameData_O[1] Tile_X5Y3_E_TT_IF/FrameData_O[20] Tile_X5Y3_E_TT_IF/FrameData_O[21]
+ Tile_X5Y3_E_TT_IF/FrameData_O[22] Tile_X5Y3_E_TT_IF/FrameData_O[23] Tile_X5Y3_E_TT_IF/FrameData_O[24]
+ Tile_X5Y3_E_TT_IF/FrameData_O[25] Tile_X5Y3_E_TT_IF/FrameData_O[26] Tile_X5Y3_E_TT_IF/FrameData_O[27]
+ Tile_X5Y3_E_TT_IF/FrameData_O[28] Tile_X5Y3_E_TT_IF/FrameData_O[29] Tile_X5Y3_E_TT_IF/FrameData_O[2]
+ Tile_X5Y3_E_TT_IF/FrameData_O[30] Tile_X5Y3_E_TT_IF/FrameData_O[31] Tile_X5Y3_E_TT_IF/FrameData_O[3]
+ Tile_X5Y3_E_TT_IF/FrameData_O[4] Tile_X5Y3_E_TT_IF/FrameData_O[5] Tile_X5Y3_E_TT_IF/FrameData_O[6]
+ Tile_X5Y3_E_TT_IF/FrameData_O[7] Tile_X5Y3_E_TT_IF/FrameData_O[8] Tile_X5Y3_E_TT_IF/FrameData_O[9]
+ Tile_X5Y3_E_TT_IF/FrameStrobe[0] Tile_X5Y3_E_TT_IF/FrameStrobe[10] Tile_X5Y3_E_TT_IF/FrameStrobe[11]
+ Tile_X5Y3_E_TT_IF/FrameStrobe[12] Tile_X5Y3_E_TT_IF/FrameStrobe[13] Tile_X5Y3_E_TT_IF/FrameStrobe[14]
+ Tile_X5Y3_E_TT_IF/FrameStrobe[15] Tile_X5Y3_E_TT_IF/FrameStrobe[16] Tile_X5Y3_E_TT_IF/FrameStrobe[17]
+ Tile_X5Y3_E_TT_IF/FrameStrobe[18] Tile_X5Y3_E_TT_IF/FrameStrobe[19] Tile_X5Y3_E_TT_IF/FrameStrobe[1]
+ Tile_X5Y3_E_TT_IF/FrameStrobe[2] Tile_X5Y3_E_TT_IF/FrameStrobe[3] Tile_X5Y3_E_TT_IF/FrameStrobe[4]
+ Tile_X5Y3_E_TT_IF/FrameStrobe[5] Tile_X5Y3_E_TT_IF/FrameStrobe[6] Tile_X5Y3_E_TT_IF/FrameStrobe[7]
+ Tile_X5Y3_E_TT_IF/FrameStrobe[8] Tile_X5Y3_E_TT_IF/FrameStrobe[9] Tile_X5Y3_E_TT_IF/FrameStrobe_O[0]
+ Tile_X5Y3_E_TT_IF/FrameStrobe_O[10] Tile_X5Y3_E_TT_IF/FrameStrobe_O[11] Tile_X5Y3_E_TT_IF/FrameStrobe_O[12]
+ Tile_X5Y3_E_TT_IF/FrameStrobe_O[13] Tile_X5Y3_E_TT_IF/FrameStrobe_O[14] Tile_X5Y3_E_TT_IF/FrameStrobe_O[15]
+ Tile_X5Y3_E_TT_IF/FrameStrobe_O[16] Tile_X5Y3_E_TT_IF/FrameStrobe_O[17] Tile_X5Y3_E_TT_IF/FrameStrobe_O[18]
+ Tile_X5Y3_E_TT_IF/FrameStrobe_O[19] Tile_X5Y3_E_TT_IF/FrameStrobe_O[1] Tile_X5Y3_E_TT_IF/FrameStrobe_O[2]
+ Tile_X5Y3_E_TT_IF/FrameStrobe_O[3] Tile_X5Y3_E_TT_IF/FrameStrobe_O[4] Tile_X5Y3_E_TT_IF/FrameStrobe_O[5]
+ Tile_X5Y3_E_TT_IF/FrameStrobe_O[6] Tile_X5Y3_E_TT_IF/FrameStrobe_O[7] Tile_X5Y3_E_TT_IF/FrameStrobe_O[8]
+ Tile_X5Y3_E_TT_IF/FrameStrobe_O[9] Tile_X5Y3_E_TT_IF/N1BEG[0] Tile_X5Y3_E_TT_IF/N1BEG[1]
+ Tile_X5Y3_E_TT_IF/N1BEG[2] Tile_X5Y3_E_TT_IF/N1BEG[3] Tile_X5Y4_E_TT_IF/N1BEG[0]
+ Tile_X5Y4_E_TT_IF/N1BEG[1] Tile_X5Y4_E_TT_IF/N1BEG[2] Tile_X5Y4_E_TT_IF/N1BEG[3]
+ Tile_X5Y3_E_TT_IF/N2BEG[0] Tile_X5Y3_E_TT_IF/N2BEG[1] Tile_X5Y3_E_TT_IF/N2BEG[2]
+ Tile_X5Y3_E_TT_IF/N2BEG[3] Tile_X5Y3_E_TT_IF/N2BEG[4] Tile_X5Y3_E_TT_IF/N2BEG[5]
+ Tile_X5Y3_E_TT_IF/N2BEG[6] Tile_X5Y3_E_TT_IF/N2BEG[7] Tile_X5Y3_E_TT_IF/N2BEGb[0]
+ Tile_X5Y3_E_TT_IF/N2BEGb[1] Tile_X5Y3_E_TT_IF/N2BEGb[2] Tile_X5Y3_E_TT_IF/N2BEGb[3]
+ Tile_X5Y3_E_TT_IF/N2BEGb[4] Tile_X5Y3_E_TT_IF/N2BEGb[5] Tile_X5Y3_E_TT_IF/N2BEGb[6]
+ Tile_X5Y3_E_TT_IF/N2BEGb[7] Tile_X5Y3_E_TT_IF/N2END[0] Tile_X5Y3_E_TT_IF/N2END[1]
+ Tile_X5Y3_E_TT_IF/N2END[2] Tile_X5Y3_E_TT_IF/N2END[3] Tile_X5Y3_E_TT_IF/N2END[4]
+ Tile_X5Y3_E_TT_IF/N2END[5] Tile_X5Y3_E_TT_IF/N2END[6] Tile_X5Y3_E_TT_IF/N2END[7]
+ Tile_X5Y4_E_TT_IF/N2BEG[0] Tile_X5Y4_E_TT_IF/N2BEG[1] Tile_X5Y4_E_TT_IF/N2BEG[2]
+ Tile_X5Y4_E_TT_IF/N2BEG[3] Tile_X5Y4_E_TT_IF/N2BEG[4] Tile_X5Y4_E_TT_IF/N2BEG[5]
+ Tile_X5Y4_E_TT_IF/N2BEG[6] Tile_X5Y4_E_TT_IF/N2BEG[7] Tile_X5Y3_E_TT_IF/N4BEG[0]
+ Tile_X5Y3_E_TT_IF/N4BEG[10] Tile_X5Y3_E_TT_IF/N4BEG[11] Tile_X5Y3_E_TT_IF/N4BEG[12]
+ Tile_X5Y3_E_TT_IF/N4BEG[13] Tile_X5Y3_E_TT_IF/N4BEG[14] Tile_X5Y3_E_TT_IF/N4BEG[15]
+ Tile_X5Y3_E_TT_IF/N4BEG[1] Tile_X5Y3_E_TT_IF/N4BEG[2] Tile_X5Y3_E_TT_IF/N4BEG[3]
+ Tile_X5Y3_E_TT_IF/N4BEG[4] Tile_X5Y3_E_TT_IF/N4BEG[5] Tile_X5Y3_E_TT_IF/N4BEG[6]
+ Tile_X5Y3_E_TT_IF/N4BEG[7] Tile_X5Y3_E_TT_IF/N4BEG[8] Tile_X5Y3_E_TT_IF/N4BEG[9]
+ Tile_X5Y4_E_TT_IF/N4BEG[0] Tile_X5Y4_E_TT_IF/N4BEG[10] Tile_X5Y4_E_TT_IF/N4BEG[11]
+ Tile_X5Y4_E_TT_IF/N4BEG[12] Tile_X5Y4_E_TT_IF/N4BEG[13] Tile_X5Y4_E_TT_IF/N4BEG[14]
+ Tile_X5Y4_E_TT_IF/N4BEG[15] Tile_X5Y4_E_TT_IF/N4BEG[1] Tile_X5Y4_E_TT_IF/N4BEG[2]
+ Tile_X5Y4_E_TT_IF/N4BEG[3] Tile_X5Y4_E_TT_IF/N4BEG[4] Tile_X5Y4_E_TT_IF/N4BEG[5]
+ Tile_X5Y4_E_TT_IF/N4BEG[6] Tile_X5Y4_E_TT_IF/N4BEG[7] Tile_X5Y4_E_TT_IF/N4BEG[8]
+ Tile_X5Y4_E_TT_IF/N4BEG[9] Tile_X5Y3_RST_N_TT_PROJECT Tile_X5Y4_E_TT_IF/S1END[0]
+ Tile_X5Y4_E_TT_IF/S1END[1] Tile_X5Y4_E_TT_IF/S1END[2] Tile_X5Y4_E_TT_IF/S1END[3]
+ Tile_X5Y3_E_TT_IF/S1END[0] Tile_X5Y3_E_TT_IF/S1END[1] Tile_X5Y3_E_TT_IF/S1END[2]
+ Tile_X5Y3_E_TT_IF/S1END[3] Tile_X5Y4_E_TT_IF/S2MID[0] Tile_X5Y4_E_TT_IF/S2MID[1]
+ Tile_X5Y4_E_TT_IF/S2MID[2] Tile_X5Y4_E_TT_IF/S2MID[3] Tile_X5Y4_E_TT_IF/S2MID[4]
+ Tile_X5Y4_E_TT_IF/S2MID[5] Tile_X5Y4_E_TT_IF/S2MID[6] Tile_X5Y4_E_TT_IF/S2MID[7]
+ Tile_X5Y4_E_TT_IF/S2END[0] Tile_X5Y4_E_TT_IF/S2END[1] Tile_X5Y4_E_TT_IF/S2END[2]
+ Tile_X5Y4_E_TT_IF/S2END[3] Tile_X5Y4_E_TT_IF/S2END[4] Tile_X5Y4_E_TT_IF/S2END[5]
+ Tile_X5Y4_E_TT_IF/S2END[6] Tile_X5Y4_E_TT_IF/S2END[7] Tile_X5Y3_E_TT_IF/S2END[0]
+ Tile_X5Y3_E_TT_IF/S2END[1] Tile_X5Y3_E_TT_IF/S2END[2] Tile_X5Y3_E_TT_IF/S2END[3]
+ Tile_X5Y3_E_TT_IF/S2END[4] Tile_X5Y3_E_TT_IF/S2END[5] Tile_X5Y3_E_TT_IF/S2END[6]
+ Tile_X5Y3_E_TT_IF/S2END[7] Tile_X5Y3_E_TT_IF/S2MID[0] Tile_X5Y3_E_TT_IF/S2MID[1]
+ Tile_X5Y3_E_TT_IF/S2MID[2] Tile_X5Y3_E_TT_IF/S2MID[3] Tile_X5Y3_E_TT_IF/S2MID[4]
+ Tile_X5Y3_E_TT_IF/S2MID[5] Tile_X5Y3_E_TT_IF/S2MID[6] Tile_X5Y3_E_TT_IF/S2MID[7]
+ Tile_X5Y4_E_TT_IF/S4END[0] Tile_X5Y4_E_TT_IF/S4END[10] Tile_X5Y4_E_TT_IF/S4END[11]
+ Tile_X5Y4_E_TT_IF/S4END[12] Tile_X5Y4_E_TT_IF/S4END[13] Tile_X5Y4_E_TT_IF/S4END[14]
+ Tile_X5Y4_E_TT_IF/S4END[15] Tile_X5Y4_E_TT_IF/S4END[1] Tile_X5Y4_E_TT_IF/S4END[2]
+ Tile_X5Y4_E_TT_IF/S4END[3] Tile_X5Y4_E_TT_IF/S4END[4] Tile_X5Y4_E_TT_IF/S4END[5]
+ Tile_X5Y4_E_TT_IF/S4END[6] Tile_X5Y4_E_TT_IF/S4END[7] Tile_X5Y4_E_TT_IF/S4END[8]
+ Tile_X5Y4_E_TT_IF/S4END[9] Tile_X5Y3_E_TT_IF/S4END[0] Tile_X5Y3_E_TT_IF/S4END[10]
+ Tile_X5Y3_E_TT_IF/S4END[11] Tile_X5Y3_E_TT_IF/S4END[12] Tile_X5Y3_E_TT_IF/S4END[13]
+ Tile_X5Y3_E_TT_IF/S4END[14] Tile_X5Y3_E_TT_IF/S4END[15] Tile_X5Y3_E_TT_IF/S4END[1]
+ Tile_X5Y3_E_TT_IF/S4END[2] Tile_X5Y3_E_TT_IF/S4END[3] Tile_X5Y3_E_TT_IF/S4END[4]
+ Tile_X5Y3_E_TT_IF/S4END[5] Tile_X5Y3_E_TT_IF/S4END[6] Tile_X5Y3_E_TT_IF/S4END[7]
+ Tile_X5Y3_E_TT_IF/S4END[8] Tile_X5Y3_E_TT_IF/S4END[9] Tile_X5Y3_UIO_IN_TT_PROJECT0
+ Tile_X5Y3_UIO_IN_TT_PROJECT1 Tile_X5Y3_UIO_IN_TT_PROJECT2 Tile_X5Y3_UIO_IN_TT_PROJECT3
+ Tile_X5Y3_UIO_IN_TT_PROJECT4 Tile_X5Y3_UIO_IN_TT_PROJECT5 Tile_X5Y3_UIO_IN_TT_PROJECT6
+ Tile_X5Y3_UIO_IN_TT_PROJECT7 Tile_X5Y3_UIO_OE_TT_PROJECT0 Tile_X5Y3_UIO_OE_TT_PROJECT1
+ Tile_X5Y3_UIO_OE_TT_PROJECT2 Tile_X5Y3_UIO_OE_TT_PROJECT3 Tile_X5Y3_UIO_OE_TT_PROJECT4
+ Tile_X5Y3_UIO_OE_TT_PROJECT5 Tile_X5Y3_UIO_OE_TT_PROJECT6 Tile_X5Y3_UIO_OE_TT_PROJECT7
+ Tile_X5Y3_UIO_OUT_TT_PROJECT0 Tile_X5Y3_UIO_OUT_TT_PROJECT1 Tile_X5Y3_UIO_OUT_TT_PROJECT2
+ Tile_X5Y3_UIO_OUT_TT_PROJECT3 Tile_X5Y3_UIO_OUT_TT_PROJECT4 Tile_X5Y3_UIO_OUT_TT_PROJECT5
+ Tile_X5Y3_UIO_OUT_TT_PROJECT6 Tile_X5Y3_UIO_OUT_TT_PROJECT7 Tile_X5Y3_UI_IN_TT_PROJECT0
+ Tile_X5Y3_UI_IN_TT_PROJECT1 Tile_X5Y3_UI_IN_TT_PROJECT2 Tile_X5Y3_UI_IN_TT_PROJECT3
+ Tile_X5Y3_UI_IN_TT_PROJECT4 Tile_X5Y3_UI_IN_TT_PROJECT5 Tile_X5Y3_UI_IN_TT_PROJECT6
+ Tile_X5Y3_UI_IN_TT_PROJECT7 Tile_X5Y3_UO_OUT_TT_PROJECT0 Tile_X5Y3_UO_OUT_TT_PROJECT1
+ Tile_X5Y3_UO_OUT_TT_PROJECT2 Tile_X5Y3_UO_OUT_TT_PROJECT3 Tile_X5Y3_UO_OUT_TT_PROJECT4
+ Tile_X5Y3_UO_OUT_TT_PROJECT5 Tile_X5Y3_UO_OUT_TT_PROJECT6 Tile_X5Y3_UO_OUT_TT_PROJECT7
+ Tile_X5Y3_E_TT_IF/UserCLK Tile_X5Y3_E_TT_IF/UserCLKo VGND VPWR Tile_X4Y3_LUT4AB/W1END[0]
+ Tile_X4Y3_LUT4AB/W1END[1] Tile_X4Y3_LUT4AB/W1END[2] Tile_X4Y3_LUT4AB/W1END[3] Tile_X4Y3_LUT4AB/W2MID[0]
+ Tile_X4Y3_LUT4AB/W2MID[1] Tile_X4Y3_LUT4AB/W2MID[2] Tile_X4Y3_LUT4AB/W2MID[3] Tile_X4Y3_LUT4AB/W2MID[4]
+ Tile_X4Y3_LUT4AB/W2MID[5] Tile_X4Y3_LUT4AB/W2MID[6] Tile_X4Y3_LUT4AB/W2MID[7] Tile_X4Y3_LUT4AB/W2END[0]
+ Tile_X4Y3_LUT4AB/W2END[1] Tile_X4Y3_LUT4AB/W2END[2] Tile_X4Y3_LUT4AB/W2END[3] Tile_X4Y3_LUT4AB/W2END[4]
+ Tile_X4Y3_LUT4AB/W2END[5] Tile_X4Y3_LUT4AB/W2END[6] Tile_X4Y3_LUT4AB/W2END[7] Tile_X4Y3_LUT4AB/W6END[0]
+ Tile_X4Y3_LUT4AB/W6END[10] Tile_X4Y3_LUT4AB/W6END[11] Tile_X4Y3_LUT4AB/W6END[1]
+ Tile_X4Y3_LUT4AB/W6END[2] Tile_X4Y3_LUT4AB/W6END[3] Tile_X4Y3_LUT4AB/W6END[4] Tile_X4Y3_LUT4AB/W6END[5]
+ Tile_X4Y3_LUT4AB/W6END[6] Tile_X4Y3_LUT4AB/W6END[7] Tile_X4Y3_LUT4AB/W6END[8] Tile_X4Y3_LUT4AB/W6END[9]
+ Tile_X4Y3_LUT4AB/WW4END[0] Tile_X4Y3_LUT4AB/WW4END[10] Tile_X4Y3_LUT4AB/WW4END[11]
+ Tile_X4Y3_LUT4AB/WW4END[12] Tile_X4Y3_LUT4AB/WW4END[13] Tile_X4Y3_LUT4AB/WW4END[14]
+ Tile_X4Y3_LUT4AB/WW4END[15] Tile_X4Y3_LUT4AB/WW4END[1] Tile_X4Y3_LUT4AB/WW4END[2]
+ Tile_X4Y3_LUT4AB/WW4END[3] Tile_X4Y3_LUT4AB/WW4END[4] Tile_X4Y3_LUT4AB/WW4END[5]
+ Tile_X4Y3_LUT4AB/WW4END[6] Tile_X4Y3_LUT4AB/WW4END[7] Tile_X4Y3_LUT4AB/WW4END[8]
+ Tile_X4Y3_LUT4AB/WW4END[9] E_TT_IF
XTile_X4Y6_LUT4AB Tile_X4Y7_LUT4AB/Co Tile_X4Y6_LUT4AB/Co Tile_X4Y6_LUT4AB/E1BEG[0]
+ Tile_X4Y6_LUT4AB/E1BEG[1] Tile_X4Y6_LUT4AB/E1BEG[2] Tile_X4Y6_LUT4AB/E1BEG[3] Tile_X4Y6_LUT4AB/E1END[0]
+ Tile_X4Y6_LUT4AB/E1END[1] Tile_X4Y6_LUT4AB/E1END[2] Tile_X4Y6_LUT4AB/E1END[3] Tile_X4Y6_LUT4AB/E2BEG[0]
+ Tile_X4Y6_LUT4AB/E2BEG[1] Tile_X4Y6_LUT4AB/E2BEG[2] Tile_X4Y6_LUT4AB/E2BEG[3] Tile_X4Y6_LUT4AB/E2BEG[4]
+ Tile_X4Y6_LUT4AB/E2BEG[5] Tile_X4Y6_LUT4AB/E2BEG[6] Tile_X4Y6_LUT4AB/E2BEG[7] Tile_X5Y6_E_TT_IF/E2END[0]
+ Tile_X5Y6_E_TT_IF/E2END[1] Tile_X5Y6_E_TT_IF/E2END[2] Tile_X5Y6_E_TT_IF/E2END[3]
+ Tile_X5Y6_E_TT_IF/E2END[4] Tile_X5Y6_E_TT_IF/E2END[5] Tile_X5Y6_E_TT_IF/E2END[6]
+ Tile_X5Y6_E_TT_IF/E2END[7] Tile_X4Y6_LUT4AB/E2END[0] Tile_X4Y6_LUT4AB/E2END[1] Tile_X4Y6_LUT4AB/E2END[2]
+ Tile_X4Y6_LUT4AB/E2END[3] Tile_X4Y6_LUT4AB/E2END[4] Tile_X4Y6_LUT4AB/E2END[5] Tile_X4Y6_LUT4AB/E2END[6]
+ Tile_X4Y6_LUT4AB/E2END[7] Tile_X4Y6_LUT4AB/E2MID[0] Tile_X4Y6_LUT4AB/E2MID[1] Tile_X4Y6_LUT4AB/E2MID[2]
+ Tile_X4Y6_LUT4AB/E2MID[3] Tile_X4Y6_LUT4AB/E2MID[4] Tile_X4Y6_LUT4AB/E2MID[5] Tile_X4Y6_LUT4AB/E2MID[6]
+ Tile_X4Y6_LUT4AB/E2MID[7] Tile_X4Y6_LUT4AB/E6BEG[0] Tile_X4Y6_LUT4AB/E6BEG[10] Tile_X4Y6_LUT4AB/E6BEG[11]
+ Tile_X4Y6_LUT4AB/E6BEG[1] Tile_X4Y6_LUT4AB/E6BEG[2] Tile_X4Y6_LUT4AB/E6BEG[3] Tile_X4Y6_LUT4AB/E6BEG[4]
+ Tile_X4Y6_LUT4AB/E6BEG[5] Tile_X4Y6_LUT4AB/E6BEG[6] Tile_X4Y6_LUT4AB/E6BEG[7] Tile_X4Y6_LUT4AB/E6BEG[8]
+ Tile_X4Y6_LUT4AB/E6BEG[9] Tile_X4Y6_LUT4AB/E6END[0] Tile_X4Y6_LUT4AB/E6END[10] Tile_X4Y6_LUT4AB/E6END[11]
+ Tile_X4Y6_LUT4AB/E6END[1] Tile_X4Y6_LUT4AB/E6END[2] Tile_X4Y6_LUT4AB/E6END[3] Tile_X4Y6_LUT4AB/E6END[4]
+ Tile_X4Y6_LUT4AB/E6END[5] Tile_X4Y6_LUT4AB/E6END[6] Tile_X4Y6_LUT4AB/E6END[7] Tile_X4Y6_LUT4AB/E6END[8]
+ Tile_X4Y6_LUT4AB/E6END[9] Tile_X4Y6_LUT4AB/EE4BEG[0] Tile_X4Y6_LUT4AB/EE4BEG[10]
+ Tile_X4Y6_LUT4AB/EE4BEG[11] Tile_X4Y6_LUT4AB/EE4BEG[12] Tile_X4Y6_LUT4AB/EE4BEG[13]
+ Tile_X4Y6_LUT4AB/EE4BEG[14] Tile_X4Y6_LUT4AB/EE4BEG[15] Tile_X4Y6_LUT4AB/EE4BEG[1]
+ Tile_X4Y6_LUT4AB/EE4BEG[2] Tile_X4Y6_LUT4AB/EE4BEG[3] Tile_X4Y6_LUT4AB/EE4BEG[4]
+ Tile_X4Y6_LUT4AB/EE4BEG[5] Tile_X4Y6_LUT4AB/EE4BEG[6] Tile_X4Y6_LUT4AB/EE4BEG[7]
+ Tile_X4Y6_LUT4AB/EE4BEG[8] Tile_X4Y6_LUT4AB/EE4BEG[9] Tile_X4Y6_LUT4AB/EE4END[0]
+ Tile_X4Y6_LUT4AB/EE4END[10] Tile_X4Y6_LUT4AB/EE4END[11] Tile_X4Y6_LUT4AB/EE4END[12]
+ Tile_X4Y6_LUT4AB/EE4END[13] Tile_X4Y6_LUT4AB/EE4END[14] Tile_X4Y6_LUT4AB/EE4END[15]
+ Tile_X4Y6_LUT4AB/EE4END[1] Tile_X4Y6_LUT4AB/EE4END[2] Tile_X4Y6_LUT4AB/EE4END[3]
+ Tile_X4Y6_LUT4AB/EE4END[4] Tile_X4Y6_LUT4AB/EE4END[5] Tile_X4Y6_LUT4AB/EE4END[6]
+ Tile_X4Y6_LUT4AB/EE4END[7] Tile_X4Y6_LUT4AB/EE4END[8] Tile_X4Y6_LUT4AB/EE4END[9]
+ Tile_X4Y6_LUT4AB/FrameData[0] Tile_X4Y6_LUT4AB/FrameData[10] Tile_X4Y6_LUT4AB/FrameData[11]
+ Tile_X4Y6_LUT4AB/FrameData[12] Tile_X4Y6_LUT4AB/FrameData[13] Tile_X4Y6_LUT4AB/FrameData[14]
+ Tile_X4Y6_LUT4AB/FrameData[15] Tile_X4Y6_LUT4AB/FrameData[16] Tile_X4Y6_LUT4AB/FrameData[17]
+ Tile_X4Y6_LUT4AB/FrameData[18] Tile_X4Y6_LUT4AB/FrameData[19] Tile_X4Y6_LUT4AB/FrameData[1]
+ Tile_X4Y6_LUT4AB/FrameData[20] Tile_X4Y6_LUT4AB/FrameData[21] Tile_X4Y6_LUT4AB/FrameData[22]
+ Tile_X4Y6_LUT4AB/FrameData[23] Tile_X4Y6_LUT4AB/FrameData[24] Tile_X4Y6_LUT4AB/FrameData[25]
+ Tile_X4Y6_LUT4AB/FrameData[26] Tile_X4Y6_LUT4AB/FrameData[27] Tile_X4Y6_LUT4AB/FrameData[28]
+ Tile_X4Y6_LUT4AB/FrameData[29] Tile_X4Y6_LUT4AB/FrameData[2] Tile_X4Y6_LUT4AB/FrameData[30]
+ Tile_X4Y6_LUT4AB/FrameData[31] Tile_X4Y6_LUT4AB/FrameData[3] Tile_X4Y6_LUT4AB/FrameData[4]
+ Tile_X4Y6_LUT4AB/FrameData[5] Tile_X4Y6_LUT4AB/FrameData[6] Tile_X4Y6_LUT4AB/FrameData[7]
+ Tile_X4Y6_LUT4AB/FrameData[8] Tile_X4Y6_LUT4AB/FrameData[9] Tile_X5Y6_E_TT_IF/FrameData[0]
+ Tile_X5Y6_E_TT_IF/FrameData[10] Tile_X5Y6_E_TT_IF/FrameData[11] Tile_X5Y6_E_TT_IF/FrameData[12]
+ Tile_X5Y6_E_TT_IF/FrameData[13] Tile_X5Y6_E_TT_IF/FrameData[14] Tile_X5Y6_E_TT_IF/FrameData[15]
+ Tile_X5Y6_E_TT_IF/FrameData[16] Tile_X5Y6_E_TT_IF/FrameData[17] Tile_X5Y6_E_TT_IF/FrameData[18]
+ Tile_X5Y6_E_TT_IF/FrameData[19] Tile_X5Y6_E_TT_IF/FrameData[1] Tile_X5Y6_E_TT_IF/FrameData[20]
+ Tile_X5Y6_E_TT_IF/FrameData[21] Tile_X5Y6_E_TT_IF/FrameData[22] Tile_X5Y6_E_TT_IF/FrameData[23]
+ Tile_X5Y6_E_TT_IF/FrameData[24] Tile_X5Y6_E_TT_IF/FrameData[25] Tile_X5Y6_E_TT_IF/FrameData[26]
+ Tile_X5Y6_E_TT_IF/FrameData[27] Tile_X5Y6_E_TT_IF/FrameData[28] Tile_X5Y6_E_TT_IF/FrameData[29]
+ Tile_X5Y6_E_TT_IF/FrameData[2] Tile_X5Y6_E_TT_IF/FrameData[30] Tile_X5Y6_E_TT_IF/FrameData[31]
+ Tile_X5Y6_E_TT_IF/FrameData[3] Tile_X5Y6_E_TT_IF/FrameData[4] Tile_X5Y6_E_TT_IF/FrameData[5]
+ Tile_X5Y6_E_TT_IF/FrameData[6] Tile_X5Y6_E_TT_IF/FrameData[7] Tile_X5Y6_E_TT_IF/FrameData[8]
+ Tile_X5Y6_E_TT_IF/FrameData[9] Tile_X4Y6_LUT4AB/FrameStrobe[0] Tile_X4Y6_LUT4AB/FrameStrobe[10]
+ Tile_X4Y6_LUT4AB/FrameStrobe[11] Tile_X4Y6_LUT4AB/FrameStrobe[12] Tile_X4Y6_LUT4AB/FrameStrobe[13]
+ Tile_X4Y6_LUT4AB/FrameStrobe[14] Tile_X4Y6_LUT4AB/FrameStrobe[15] Tile_X4Y6_LUT4AB/FrameStrobe[16]
+ Tile_X4Y6_LUT4AB/FrameStrobe[17] Tile_X4Y6_LUT4AB/FrameStrobe[18] Tile_X4Y6_LUT4AB/FrameStrobe[19]
+ Tile_X4Y6_LUT4AB/FrameStrobe[1] Tile_X4Y6_LUT4AB/FrameStrobe[2] Tile_X4Y6_LUT4AB/FrameStrobe[3]
+ Tile_X4Y6_LUT4AB/FrameStrobe[4] Tile_X4Y6_LUT4AB/FrameStrobe[5] Tile_X4Y6_LUT4AB/FrameStrobe[6]
+ Tile_X4Y6_LUT4AB/FrameStrobe[7] Tile_X4Y6_LUT4AB/FrameStrobe[8] Tile_X4Y6_LUT4AB/FrameStrobe[9]
+ Tile_X4Y5_LUT4AB/FrameStrobe[0] Tile_X4Y5_LUT4AB/FrameStrobe[10] Tile_X4Y5_LUT4AB/FrameStrobe[11]
+ Tile_X4Y5_LUT4AB/FrameStrobe[12] Tile_X4Y5_LUT4AB/FrameStrobe[13] Tile_X4Y5_LUT4AB/FrameStrobe[14]
+ Tile_X4Y5_LUT4AB/FrameStrobe[15] Tile_X4Y5_LUT4AB/FrameStrobe[16] Tile_X4Y5_LUT4AB/FrameStrobe[17]
+ Tile_X4Y5_LUT4AB/FrameStrobe[18] Tile_X4Y5_LUT4AB/FrameStrobe[19] Tile_X4Y5_LUT4AB/FrameStrobe[1]
+ Tile_X4Y5_LUT4AB/FrameStrobe[2] Tile_X4Y5_LUT4AB/FrameStrobe[3] Tile_X4Y5_LUT4AB/FrameStrobe[4]
+ Tile_X4Y5_LUT4AB/FrameStrobe[5] Tile_X4Y5_LUT4AB/FrameStrobe[6] Tile_X4Y5_LUT4AB/FrameStrobe[7]
+ Tile_X4Y5_LUT4AB/FrameStrobe[8] Tile_X4Y5_LUT4AB/FrameStrobe[9] Tile_X4Y6_LUT4AB/N1BEG[0]
+ Tile_X4Y6_LUT4AB/N1BEG[1] Tile_X4Y6_LUT4AB/N1BEG[2] Tile_X4Y6_LUT4AB/N1BEG[3] Tile_X4Y7_LUT4AB/N1BEG[0]
+ Tile_X4Y7_LUT4AB/N1BEG[1] Tile_X4Y7_LUT4AB/N1BEG[2] Tile_X4Y7_LUT4AB/N1BEG[3] Tile_X4Y6_LUT4AB/N2BEG[0]
+ Tile_X4Y6_LUT4AB/N2BEG[1] Tile_X4Y6_LUT4AB/N2BEG[2] Tile_X4Y6_LUT4AB/N2BEG[3] Tile_X4Y6_LUT4AB/N2BEG[4]
+ Tile_X4Y6_LUT4AB/N2BEG[5] Tile_X4Y6_LUT4AB/N2BEG[6] Tile_X4Y6_LUT4AB/N2BEG[7] Tile_X4Y5_LUT4AB/N2END[0]
+ Tile_X4Y5_LUT4AB/N2END[1] Tile_X4Y5_LUT4AB/N2END[2] Tile_X4Y5_LUT4AB/N2END[3] Tile_X4Y5_LUT4AB/N2END[4]
+ Tile_X4Y5_LUT4AB/N2END[5] Tile_X4Y5_LUT4AB/N2END[6] Tile_X4Y5_LUT4AB/N2END[7] Tile_X4Y6_LUT4AB/N2END[0]
+ Tile_X4Y6_LUT4AB/N2END[1] Tile_X4Y6_LUT4AB/N2END[2] Tile_X4Y6_LUT4AB/N2END[3] Tile_X4Y6_LUT4AB/N2END[4]
+ Tile_X4Y6_LUT4AB/N2END[5] Tile_X4Y6_LUT4AB/N2END[6] Tile_X4Y6_LUT4AB/N2END[7] Tile_X4Y7_LUT4AB/N2BEG[0]
+ Tile_X4Y7_LUT4AB/N2BEG[1] Tile_X4Y7_LUT4AB/N2BEG[2] Tile_X4Y7_LUT4AB/N2BEG[3] Tile_X4Y7_LUT4AB/N2BEG[4]
+ Tile_X4Y7_LUT4AB/N2BEG[5] Tile_X4Y7_LUT4AB/N2BEG[6] Tile_X4Y7_LUT4AB/N2BEG[7] Tile_X4Y6_LUT4AB/N4BEG[0]
+ Tile_X4Y6_LUT4AB/N4BEG[10] Tile_X4Y6_LUT4AB/N4BEG[11] Tile_X4Y6_LUT4AB/N4BEG[12]
+ Tile_X4Y6_LUT4AB/N4BEG[13] Tile_X4Y6_LUT4AB/N4BEG[14] Tile_X4Y6_LUT4AB/N4BEG[15]
+ Tile_X4Y6_LUT4AB/N4BEG[1] Tile_X4Y6_LUT4AB/N4BEG[2] Tile_X4Y6_LUT4AB/N4BEG[3] Tile_X4Y6_LUT4AB/N4BEG[4]
+ Tile_X4Y6_LUT4AB/N4BEG[5] Tile_X4Y6_LUT4AB/N4BEG[6] Tile_X4Y6_LUT4AB/N4BEG[7] Tile_X4Y6_LUT4AB/N4BEG[8]
+ Tile_X4Y6_LUT4AB/N4BEG[9] Tile_X4Y7_LUT4AB/N4BEG[0] Tile_X4Y7_LUT4AB/N4BEG[10] Tile_X4Y7_LUT4AB/N4BEG[11]
+ Tile_X4Y7_LUT4AB/N4BEG[12] Tile_X4Y7_LUT4AB/N4BEG[13] Tile_X4Y7_LUT4AB/N4BEG[14]
+ Tile_X4Y7_LUT4AB/N4BEG[15] Tile_X4Y7_LUT4AB/N4BEG[1] Tile_X4Y7_LUT4AB/N4BEG[2] Tile_X4Y7_LUT4AB/N4BEG[3]
+ Tile_X4Y7_LUT4AB/N4BEG[4] Tile_X4Y7_LUT4AB/N4BEG[5] Tile_X4Y7_LUT4AB/N4BEG[6] Tile_X4Y7_LUT4AB/N4BEG[7]
+ Tile_X4Y7_LUT4AB/N4BEG[8] Tile_X4Y7_LUT4AB/N4BEG[9] Tile_X4Y6_LUT4AB/NN4BEG[0] Tile_X4Y6_LUT4AB/NN4BEG[10]
+ Tile_X4Y6_LUT4AB/NN4BEG[11] Tile_X4Y6_LUT4AB/NN4BEG[12] Tile_X4Y6_LUT4AB/NN4BEG[13]
+ Tile_X4Y6_LUT4AB/NN4BEG[14] Tile_X4Y6_LUT4AB/NN4BEG[15] Tile_X4Y6_LUT4AB/NN4BEG[1]
+ Tile_X4Y6_LUT4AB/NN4BEG[2] Tile_X4Y6_LUT4AB/NN4BEG[3] Tile_X4Y6_LUT4AB/NN4BEG[4]
+ Tile_X4Y6_LUT4AB/NN4BEG[5] Tile_X4Y6_LUT4AB/NN4BEG[6] Tile_X4Y6_LUT4AB/NN4BEG[7]
+ Tile_X4Y6_LUT4AB/NN4BEG[8] Tile_X4Y6_LUT4AB/NN4BEG[9] Tile_X4Y7_LUT4AB/NN4BEG[0]
+ Tile_X4Y7_LUT4AB/NN4BEG[10] Tile_X4Y7_LUT4AB/NN4BEG[11] Tile_X4Y7_LUT4AB/NN4BEG[12]
+ Tile_X4Y7_LUT4AB/NN4BEG[13] Tile_X4Y7_LUT4AB/NN4BEG[14] Tile_X4Y7_LUT4AB/NN4BEG[15]
+ Tile_X4Y7_LUT4AB/NN4BEG[1] Tile_X4Y7_LUT4AB/NN4BEG[2] Tile_X4Y7_LUT4AB/NN4BEG[3]
+ Tile_X4Y7_LUT4AB/NN4BEG[4] Tile_X4Y7_LUT4AB/NN4BEG[5] Tile_X4Y7_LUT4AB/NN4BEG[6]
+ Tile_X4Y7_LUT4AB/NN4BEG[7] Tile_X4Y7_LUT4AB/NN4BEG[8] Tile_X4Y7_LUT4AB/NN4BEG[9]
+ Tile_X4Y7_LUT4AB/S1END[0] Tile_X4Y7_LUT4AB/S1END[1] Tile_X4Y7_LUT4AB/S1END[2] Tile_X4Y7_LUT4AB/S1END[3]
+ Tile_X4Y6_LUT4AB/S1END[0] Tile_X4Y6_LUT4AB/S1END[1] Tile_X4Y6_LUT4AB/S1END[2] Tile_X4Y6_LUT4AB/S1END[3]
+ Tile_X4Y7_LUT4AB/S2MID[0] Tile_X4Y7_LUT4AB/S2MID[1] Tile_X4Y7_LUT4AB/S2MID[2] Tile_X4Y7_LUT4AB/S2MID[3]
+ Tile_X4Y7_LUT4AB/S2MID[4] Tile_X4Y7_LUT4AB/S2MID[5] Tile_X4Y7_LUT4AB/S2MID[6] Tile_X4Y7_LUT4AB/S2MID[7]
+ Tile_X4Y7_LUT4AB/S2END[0] Tile_X4Y7_LUT4AB/S2END[1] Tile_X4Y7_LUT4AB/S2END[2] Tile_X4Y7_LUT4AB/S2END[3]
+ Tile_X4Y7_LUT4AB/S2END[4] Tile_X4Y7_LUT4AB/S2END[5] Tile_X4Y7_LUT4AB/S2END[6] Tile_X4Y7_LUT4AB/S2END[7]
+ Tile_X4Y6_LUT4AB/S2END[0] Tile_X4Y6_LUT4AB/S2END[1] Tile_X4Y6_LUT4AB/S2END[2] Tile_X4Y6_LUT4AB/S2END[3]
+ Tile_X4Y6_LUT4AB/S2END[4] Tile_X4Y6_LUT4AB/S2END[5] Tile_X4Y6_LUT4AB/S2END[6] Tile_X4Y6_LUT4AB/S2END[7]
+ Tile_X4Y6_LUT4AB/S2MID[0] Tile_X4Y6_LUT4AB/S2MID[1] Tile_X4Y6_LUT4AB/S2MID[2] Tile_X4Y6_LUT4AB/S2MID[3]
+ Tile_X4Y6_LUT4AB/S2MID[4] Tile_X4Y6_LUT4AB/S2MID[5] Tile_X4Y6_LUT4AB/S2MID[6] Tile_X4Y6_LUT4AB/S2MID[7]
+ Tile_X4Y7_LUT4AB/S4END[0] Tile_X4Y7_LUT4AB/S4END[10] Tile_X4Y7_LUT4AB/S4END[11]
+ Tile_X4Y7_LUT4AB/S4END[12] Tile_X4Y7_LUT4AB/S4END[13] Tile_X4Y7_LUT4AB/S4END[14]
+ Tile_X4Y7_LUT4AB/S4END[15] Tile_X4Y7_LUT4AB/S4END[1] Tile_X4Y7_LUT4AB/S4END[2] Tile_X4Y7_LUT4AB/S4END[3]
+ Tile_X4Y7_LUT4AB/S4END[4] Tile_X4Y7_LUT4AB/S4END[5] Tile_X4Y7_LUT4AB/S4END[6] Tile_X4Y7_LUT4AB/S4END[7]
+ Tile_X4Y7_LUT4AB/S4END[8] Tile_X4Y7_LUT4AB/S4END[9] Tile_X4Y6_LUT4AB/S4END[0] Tile_X4Y6_LUT4AB/S4END[10]
+ Tile_X4Y6_LUT4AB/S4END[11] Tile_X4Y6_LUT4AB/S4END[12] Tile_X4Y6_LUT4AB/S4END[13]
+ Tile_X4Y6_LUT4AB/S4END[14] Tile_X4Y6_LUT4AB/S4END[15] Tile_X4Y6_LUT4AB/S4END[1]
+ Tile_X4Y6_LUT4AB/S4END[2] Tile_X4Y6_LUT4AB/S4END[3] Tile_X4Y6_LUT4AB/S4END[4] Tile_X4Y6_LUT4AB/S4END[5]
+ Tile_X4Y6_LUT4AB/S4END[6] Tile_X4Y6_LUT4AB/S4END[7] Tile_X4Y6_LUT4AB/S4END[8] Tile_X4Y6_LUT4AB/S4END[9]
+ Tile_X4Y7_LUT4AB/SS4END[0] Tile_X4Y7_LUT4AB/SS4END[10] Tile_X4Y7_LUT4AB/SS4END[11]
+ Tile_X4Y7_LUT4AB/SS4END[12] Tile_X4Y7_LUT4AB/SS4END[13] Tile_X4Y7_LUT4AB/SS4END[14]
+ Tile_X4Y7_LUT4AB/SS4END[15] Tile_X4Y7_LUT4AB/SS4END[1] Tile_X4Y7_LUT4AB/SS4END[2]
+ Tile_X4Y7_LUT4AB/SS4END[3] Tile_X4Y7_LUT4AB/SS4END[4] Tile_X4Y7_LUT4AB/SS4END[5]
+ Tile_X4Y7_LUT4AB/SS4END[6] Tile_X4Y7_LUT4AB/SS4END[7] Tile_X4Y7_LUT4AB/SS4END[8]
+ Tile_X4Y7_LUT4AB/SS4END[9] Tile_X4Y6_LUT4AB/SS4END[0] Tile_X4Y6_LUT4AB/SS4END[10]
+ Tile_X4Y6_LUT4AB/SS4END[11] Tile_X4Y6_LUT4AB/SS4END[12] Tile_X4Y6_LUT4AB/SS4END[13]
+ Tile_X4Y6_LUT4AB/SS4END[14] Tile_X4Y6_LUT4AB/SS4END[15] Tile_X4Y6_LUT4AB/SS4END[1]
+ Tile_X4Y6_LUT4AB/SS4END[2] Tile_X4Y6_LUT4AB/SS4END[3] Tile_X4Y6_LUT4AB/SS4END[4]
+ Tile_X4Y6_LUT4AB/SS4END[5] Tile_X4Y6_LUT4AB/SS4END[6] Tile_X4Y6_LUT4AB/SS4END[7]
+ Tile_X4Y6_LUT4AB/SS4END[8] Tile_X4Y6_LUT4AB/SS4END[9] Tile_X4Y6_LUT4AB/UserCLK Tile_X4Y5_LUT4AB/UserCLK
+ VGND VPWR Tile_X4Y6_LUT4AB/W1BEG[0] Tile_X4Y6_LUT4AB/W1BEG[1] Tile_X4Y6_LUT4AB/W1BEG[2]
+ Tile_X4Y6_LUT4AB/W1BEG[3] Tile_X4Y6_LUT4AB/W1END[0] Tile_X4Y6_LUT4AB/W1END[1] Tile_X4Y6_LUT4AB/W1END[2]
+ Tile_X4Y6_LUT4AB/W1END[3] Tile_X4Y6_LUT4AB/W2BEG[0] Tile_X4Y6_LUT4AB/W2BEG[1] Tile_X4Y6_LUT4AB/W2BEG[2]
+ Tile_X4Y6_LUT4AB/W2BEG[3] Tile_X4Y6_LUT4AB/W2BEG[4] Tile_X4Y6_LUT4AB/W2BEG[5] Tile_X4Y6_LUT4AB/W2BEG[6]
+ Tile_X4Y6_LUT4AB/W2BEG[7] Tile_X3Y6_LUT4AB/W2END[0] Tile_X3Y6_LUT4AB/W2END[1] Tile_X3Y6_LUT4AB/W2END[2]
+ Tile_X3Y6_LUT4AB/W2END[3] Tile_X3Y6_LUT4AB/W2END[4] Tile_X3Y6_LUT4AB/W2END[5] Tile_X3Y6_LUT4AB/W2END[6]
+ Tile_X3Y6_LUT4AB/W2END[7] Tile_X4Y6_LUT4AB/W2END[0] Tile_X4Y6_LUT4AB/W2END[1] Tile_X4Y6_LUT4AB/W2END[2]
+ Tile_X4Y6_LUT4AB/W2END[3] Tile_X4Y6_LUT4AB/W2END[4] Tile_X4Y6_LUT4AB/W2END[5] Tile_X4Y6_LUT4AB/W2END[6]
+ Tile_X4Y6_LUT4AB/W2END[7] Tile_X4Y6_LUT4AB/W2MID[0] Tile_X4Y6_LUT4AB/W2MID[1] Tile_X4Y6_LUT4AB/W2MID[2]
+ Tile_X4Y6_LUT4AB/W2MID[3] Tile_X4Y6_LUT4AB/W2MID[4] Tile_X4Y6_LUT4AB/W2MID[5] Tile_X4Y6_LUT4AB/W2MID[6]
+ Tile_X4Y6_LUT4AB/W2MID[7] Tile_X4Y6_LUT4AB/W6BEG[0] Tile_X4Y6_LUT4AB/W6BEG[10] Tile_X4Y6_LUT4AB/W6BEG[11]
+ Tile_X4Y6_LUT4AB/W6BEG[1] Tile_X4Y6_LUT4AB/W6BEG[2] Tile_X4Y6_LUT4AB/W6BEG[3] Tile_X4Y6_LUT4AB/W6BEG[4]
+ Tile_X4Y6_LUT4AB/W6BEG[5] Tile_X4Y6_LUT4AB/W6BEG[6] Tile_X4Y6_LUT4AB/W6BEG[7] Tile_X4Y6_LUT4AB/W6BEG[8]
+ Tile_X4Y6_LUT4AB/W6BEG[9] Tile_X4Y6_LUT4AB/W6END[0] Tile_X4Y6_LUT4AB/W6END[10] Tile_X4Y6_LUT4AB/W6END[11]
+ Tile_X4Y6_LUT4AB/W6END[1] Tile_X4Y6_LUT4AB/W6END[2] Tile_X4Y6_LUT4AB/W6END[3] Tile_X4Y6_LUT4AB/W6END[4]
+ Tile_X4Y6_LUT4AB/W6END[5] Tile_X4Y6_LUT4AB/W6END[6] Tile_X4Y6_LUT4AB/W6END[7] Tile_X4Y6_LUT4AB/W6END[8]
+ Tile_X4Y6_LUT4AB/W6END[9] Tile_X4Y6_LUT4AB/WW4BEG[0] Tile_X4Y6_LUT4AB/WW4BEG[10]
+ Tile_X4Y6_LUT4AB/WW4BEG[11] Tile_X4Y6_LUT4AB/WW4BEG[12] Tile_X4Y6_LUT4AB/WW4BEG[13]
+ Tile_X4Y6_LUT4AB/WW4BEG[14] Tile_X4Y6_LUT4AB/WW4BEG[15] Tile_X4Y6_LUT4AB/WW4BEG[1]
+ Tile_X4Y6_LUT4AB/WW4BEG[2] Tile_X4Y6_LUT4AB/WW4BEG[3] Tile_X4Y6_LUT4AB/WW4BEG[4]
+ Tile_X4Y6_LUT4AB/WW4BEG[5] Tile_X4Y6_LUT4AB/WW4BEG[6] Tile_X4Y6_LUT4AB/WW4BEG[7]
+ Tile_X4Y6_LUT4AB/WW4BEG[8] Tile_X4Y6_LUT4AB/WW4BEG[9] Tile_X4Y6_LUT4AB/WW4END[0]
+ Tile_X4Y6_LUT4AB/WW4END[10] Tile_X4Y6_LUT4AB/WW4END[11] Tile_X4Y6_LUT4AB/WW4END[12]
+ Tile_X4Y6_LUT4AB/WW4END[13] Tile_X4Y6_LUT4AB/WW4END[14] Tile_X4Y6_LUT4AB/WW4END[15]
+ Tile_X4Y6_LUT4AB/WW4END[1] Tile_X4Y6_LUT4AB/WW4END[2] Tile_X4Y6_LUT4AB/WW4END[3]
+ Tile_X4Y6_LUT4AB/WW4END[4] Tile_X4Y6_LUT4AB/WW4END[5] Tile_X4Y6_LUT4AB/WW4END[6]
+ Tile_X4Y6_LUT4AB/WW4END[7] Tile_X4Y6_LUT4AB/WW4END[8] Tile_X4Y6_LUT4AB/WW4END[9]
+ LUT4AB
XTile_X5Y1_IHP_SRAM Tile_X5Y2_ADDR_SRAM0 Tile_X5Y2_ADDR_SRAM1 Tile_X5Y2_ADDR_SRAM2
+ Tile_X5Y2_ADDR_SRAM3 Tile_X5Y2_ADDR_SRAM4 Tile_X5Y2_ADDR_SRAM5 Tile_X5Y2_ADDR_SRAM6
+ Tile_X5Y2_ADDR_SRAM7 Tile_X5Y2_ADDR_SRAM8 Tile_X5Y2_ADDR_SRAM9 Tile_X5Y2_BM_SRAM0
+ Tile_X5Y2_BM_SRAM1 Tile_X5Y2_BM_SRAM10 Tile_X5Y2_BM_SRAM11 Tile_X5Y2_BM_SRAM12 Tile_X5Y2_BM_SRAM13
+ Tile_X5Y2_BM_SRAM14 Tile_X5Y2_BM_SRAM15 Tile_X5Y2_BM_SRAM16 Tile_X5Y2_BM_SRAM17
+ Tile_X5Y2_BM_SRAM18 Tile_X5Y2_BM_SRAM19 Tile_X5Y2_BM_SRAM2 Tile_X5Y2_BM_SRAM20 Tile_X5Y2_BM_SRAM21
+ Tile_X5Y2_BM_SRAM22 Tile_X5Y2_BM_SRAM23 Tile_X5Y2_BM_SRAM24 Tile_X5Y2_BM_SRAM25
+ Tile_X5Y2_BM_SRAM26 Tile_X5Y2_BM_SRAM27 Tile_X5Y2_BM_SRAM28 Tile_X5Y2_BM_SRAM29
+ Tile_X5Y2_BM_SRAM3 Tile_X5Y2_BM_SRAM30 Tile_X5Y2_BM_SRAM31 Tile_X5Y2_BM_SRAM4 Tile_X5Y2_BM_SRAM5
+ Tile_X5Y2_BM_SRAM6 Tile_X5Y2_BM_SRAM7 Tile_X5Y2_BM_SRAM8 Tile_X5Y2_BM_SRAM9 Tile_X5Y2_CLK_SRAM
+ Tile_X5Y2_CONFIGURED_top Tile_X5Y2_DIN_SRAM0 Tile_X5Y2_DIN_SRAM1 Tile_X5Y2_DIN_SRAM10
+ Tile_X5Y2_DIN_SRAM11 Tile_X5Y2_DIN_SRAM12 Tile_X5Y2_DIN_SRAM13 Tile_X5Y2_DIN_SRAM14
+ Tile_X5Y2_DIN_SRAM15 Tile_X5Y2_DIN_SRAM16 Tile_X5Y2_DIN_SRAM17 Tile_X5Y2_DIN_SRAM18
+ Tile_X5Y2_DIN_SRAM19 Tile_X5Y2_DIN_SRAM2 Tile_X5Y2_DIN_SRAM20 Tile_X5Y2_DIN_SRAM21
+ Tile_X5Y2_DIN_SRAM22 Tile_X5Y2_DIN_SRAM23 Tile_X5Y2_DIN_SRAM24 Tile_X5Y2_DIN_SRAM25
+ Tile_X5Y2_DIN_SRAM26 Tile_X5Y2_DIN_SRAM27 Tile_X5Y2_DIN_SRAM28 Tile_X5Y2_DIN_SRAM29
+ Tile_X5Y2_DIN_SRAM3 Tile_X5Y2_DIN_SRAM30 Tile_X5Y2_DIN_SRAM31 Tile_X5Y2_DIN_SRAM4
+ Tile_X5Y2_DIN_SRAM5 Tile_X5Y2_DIN_SRAM6 Tile_X5Y2_DIN_SRAM7 Tile_X5Y2_DIN_SRAM8
+ Tile_X5Y2_DIN_SRAM9 Tile_X5Y2_DOUT_SRAM0 Tile_X5Y2_DOUT_SRAM1 Tile_X5Y2_DOUT_SRAM10
+ Tile_X5Y2_DOUT_SRAM11 Tile_X5Y2_DOUT_SRAM12 Tile_X5Y2_DOUT_SRAM13 Tile_X5Y2_DOUT_SRAM14
+ Tile_X5Y2_DOUT_SRAM15 Tile_X5Y2_DOUT_SRAM16 Tile_X5Y2_DOUT_SRAM17 Tile_X5Y2_DOUT_SRAM18
+ Tile_X5Y2_DOUT_SRAM19 Tile_X5Y2_DOUT_SRAM2 Tile_X5Y2_DOUT_SRAM20 Tile_X5Y2_DOUT_SRAM21
+ Tile_X5Y2_DOUT_SRAM22 Tile_X5Y2_DOUT_SRAM23 Tile_X5Y2_DOUT_SRAM24 Tile_X5Y2_DOUT_SRAM25
+ Tile_X5Y2_DOUT_SRAM26 Tile_X5Y2_DOUT_SRAM27 Tile_X5Y2_DOUT_SRAM28 Tile_X5Y2_DOUT_SRAM29
+ Tile_X5Y2_DOUT_SRAM3 Tile_X5Y2_DOUT_SRAM30 Tile_X5Y2_DOUT_SRAM31 Tile_X5Y2_DOUT_SRAM4
+ Tile_X5Y2_DOUT_SRAM5 Tile_X5Y2_DOUT_SRAM6 Tile_X5Y2_DOUT_SRAM7 Tile_X5Y2_DOUT_SRAM8
+ Tile_X5Y2_DOUT_SRAM9 Tile_X5Y2_MEN_SRAM Tile_X5Y2_REN_SRAM Tile_X5Y2_TIE_HIGH_SRAM
+ Tile_X5Y2_TIE_LOW_SRAM Tile_X4Y1_LUT4AB/E1BEG[0] Tile_X4Y1_LUT4AB/E1BEG[1] Tile_X4Y1_LUT4AB/E1BEG[2]
+ Tile_X4Y1_LUT4AB/E1BEG[3] Tile_X4Y1_LUT4AB/E2BEGb[0] Tile_X4Y1_LUT4AB/E2BEGb[1]
+ Tile_X4Y1_LUT4AB/E2BEGb[2] Tile_X4Y1_LUT4AB/E2BEGb[3] Tile_X4Y1_LUT4AB/E2BEGb[4]
+ Tile_X4Y1_LUT4AB/E2BEGb[5] Tile_X4Y1_LUT4AB/E2BEGb[6] Tile_X4Y1_LUT4AB/E2BEGb[7]
+ Tile_X4Y1_LUT4AB/E2BEG[0] Tile_X4Y1_LUT4AB/E2BEG[1] Tile_X4Y1_LUT4AB/E2BEG[2] Tile_X4Y1_LUT4AB/E2BEG[3]
+ Tile_X4Y1_LUT4AB/E2BEG[4] Tile_X4Y1_LUT4AB/E2BEG[5] Tile_X4Y1_LUT4AB/E2BEG[6] Tile_X4Y1_LUT4AB/E2BEG[7]
+ Tile_X4Y1_LUT4AB/E6BEG[0] Tile_X4Y1_LUT4AB/E6BEG[10] Tile_X4Y1_LUT4AB/E6BEG[11]
+ Tile_X4Y1_LUT4AB/E6BEG[1] Tile_X4Y1_LUT4AB/E6BEG[2] Tile_X4Y1_LUT4AB/E6BEG[3] Tile_X4Y1_LUT4AB/E6BEG[4]
+ Tile_X4Y1_LUT4AB/E6BEG[5] Tile_X4Y1_LUT4AB/E6BEG[6] Tile_X4Y1_LUT4AB/E6BEG[7] Tile_X4Y1_LUT4AB/E6BEG[8]
+ Tile_X4Y1_LUT4AB/E6BEG[9] Tile_X4Y1_LUT4AB/EE4BEG[0] Tile_X4Y1_LUT4AB/EE4BEG[10]
+ Tile_X4Y1_LUT4AB/EE4BEG[11] Tile_X4Y1_LUT4AB/EE4BEG[12] Tile_X4Y1_LUT4AB/EE4BEG[13]
+ Tile_X4Y1_LUT4AB/EE4BEG[14] Tile_X4Y1_LUT4AB/EE4BEG[15] Tile_X4Y1_LUT4AB/EE4BEG[1]
+ Tile_X4Y1_LUT4AB/EE4BEG[2] Tile_X4Y1_LUT4AB/EE4BEG[3] Tile_X4Y1_LUT4AB/EE4BEG[4]
+ Tile_X4Y1_LUT4AB/EE4BEG[5] Tile_X4Y1_LUT4AB/EE4BEG[6] Tile_X4Y1_LUT4AB/EE4BEG[7]
+ Tile_X4Y1_LUT4AB/EE4BEG[8] Tile_X4Y1_LUT4AB/EE4BEG[9] Tile_X4Y1_LUT4AB/FrameData_O[0]
+ Tile_X4Y1_LUT4AB/FrameData_O[10] Tile_X4Y1_LUT4AB/FrameData_O[11] Tile_X4Y1_LUT4AB/FrameData_O[12]
+ Tile_X4Y1_LUT4AB/FrameData_O[13] Tile_X4Y1_LUT4AB/FrameData_O[14] Tile_X4Y1_LUT4AB/FrameData_O[15]
+ Tile_X4Y1_LUT4AB/FrameData_O[16] Tile_X4Y1_LUT4AB/FrameData_O[17] Tile_X4Y1_LUT4AB/FrameData_O[18]
+ Tile_X4Y1_LUT4AB/FrameData_O[19] Tile_X4Y1_LUT4AB/FrameData_O[1] Tile_X4Y1_LUT4AB/FrameData_O[20]
+ Tile_X4Y1_LUT4AB/FrameData_O[21] Tile_X4Y1_LUT4AB/FrameData_O[22] Tile_X4Y1_LUT4AB/FrameData_O[23]
+ Tile_X4Y1_LUT4AB/FrameData_O[24] Tile_X4Y1_LUT4AB/FrameData_O[25] Tile_X4Y1_LUT4AB/FrameData_O[26]
+ Tile_X4Y1_LUT4AB/FrameData_O[27] Tile_X4Y1_LUT4AB/FrameData_O[28] Tile_X4Y1_LUT4AB/FrameData_O[29]
+ Tile_X4Y1_LUT4AB/FrameData_O[2] Tile_X4Y1_LUT4AB/FrameData_O[30] Tile_X4Y1_LUT4AB/FrameData_O[31]
+ Tile_X4Y1_LUT4AB/FrameData_O[3] Tile_X4Y1_LUT4AB/FrameData_O[4] Tile_X4Y1_LUT4AB/FrameData_O[5]
+ Tile_X4Y1_LUT4AB/FrameData_O[6] Tile_X4Y1_LUT4AB/FrameData_O[7] Tile_X4Y1_LUT4AB/FrameData_O[8]
+ Tile_X4Y1_LUT4AB/FrameData_O[9] Tile_X5Y1_IHP_SRAM/Tile_X0Y0_FrameData_O[0] Tile_X5Y1_IHP_SRAM/Tile_X0Y0_FrameData_O[10]
+ Tile_X5Y1_IHP_SRAM/Tile_X0Y0_FrameData_O[11] Tile_X5Y1_IHP_SRAM/Tile_X0Y0_FrameData_O[12]
+ Tile_X5Y1_IHP_SRAM/Tile_X0Y0_FrameData_O[13] Tile_X5Y1_IHP_SRAM/Tile_X0Y0_FrameData_O[14]
+ Tile_X5Y1_IHP_SRAM/Tile_X0Y0_FrameData_O[15] Tile_X5Y1_IHP_SRAM/Tile_X0Y0_FrameData_O[16]
+ Tile_X5Y1_IHP_SRAM/Tile_X0Y0_FrameData_O[17] Tile_X5Y1_IHP_SRAM/Tile_X0Y0_FrameData_O[18]
+ Tile_X5Y1_IHP_SRAM/Tile_X0Y0_FrameData_O[19] Tile_X5Y1_IHP_SRAM/Tile_X0Y0_FrameData_O[1]
+ Tile_X5Y1_IHP_SRAM/Tile_X0Y0_FrameData_O[20] Tile_X5Y1_IHP_SRAM/Tile_X0Y0_FrameData_O[21]
+ Tile_X5Y1_IHP_SRAM/Tile_X0Y0_FrameData_O[22] Tile_X5Y1_IHP_SRAM/Tile_X0Y0_FrameData_O[23]
+ Tile_X5Y1_IHP_SRAM/Tile_X0Y0_FrameData_O[24] Tile_X5Y1_IHP_SRAM/Tile_X0Y0_FrameData_O[25]
+ Tile_X5Y1_IHP_SRAM/Tile_X0Y0_FrameData_O[26] Tile_X5Y1_IHP_SRAM/Tile_X0Y0_FrameData_O[27]
+ Tile_X5Y1_IHP_SRAM/Tile_X0Y0_FrameData_O[28] Tile_X5Y1_IHP_SRAM/Tile_X0Y0_FrameData_O[29]
+ Tile_X5Y1_IHP_SRAM/Tile_X0Y0_FrameData_O[2] Tile_X5Y1_IHP_SRAM/Tile_X0Y0_FrameData_O[30]
+ Tile_X5Y1_IHP_SRAM/Tile_X0Y0_FrameData_O[31] Tile_X5Y1_IHP_SRAM/Tile_X0Y0_FrameData_O[3]
+ Tile_X5Y1_IHP_SRAM/Tile_X0Y0_FrameData_O[4] Tile_X5Y1_IHP_SRAM/Tile_X0Y0_FrameData_O[5]
+ Tile_X5Y1_IHP_SRAM/Tile_X0Y0_FrameData_O[6] Tile_X5Y1_IHP_SRAM/Tile_X0Y0_FrameData_O[7]
+ Tile_X5Y1_IHP_SRAM/Tile_X0Y0_FrameData_O[8] Tile_X5Y1_IHP_SRAM/Tile_X0Y0_FrameData_O[9]
+ Tile_X5Y0_NE_term/FrameStrobe[0] Tile_X5Y0_NE_term/FrameStrobe[10] Tile_X5Y0_NE_term/FrameStrobe[11]
+ Tile_X5Y0_NE_term/FrameStrobe[12] Tile_X5Y0_NE_term/FrameStrobe[13] Tile_X5Y0_NE_term/FrameStrobe[14]
+ Tile_X5Y0_NE_term/FrameStrobe[15] Tile_X5Y0_NE_term/FrameStrobe[16] Tile_X5Y0_NE_term/FrameStrobe[17]
+ Tile_X5Y0_NE_term/FrameStrobe[18] Tile_X5Y0_NE_term/FrameStrobe[19] Tile_X5Y0_NE_term/FrameStrobe[1]
+ Tile_X5Y0_NE_term/FrameStrobe[2] Tile_X5Y0_NE_term/FrameStrobe[3] Tile_X5Y0_NE_term/FrameStrobe[4]
+ Tile_X5Y0_NE_term/FrameStrobe[5] Tile_X5Y0_NE_term/FrameStrobe[6] Tile_X5Y0_NE_term/FrameStrobe[7]
+ Tile_X5Y0_NE_term/FrameStrobe[8] Tile_X5Y0_NE_term/FrameStrobe[9] Tile_X5Y0_NE_term/N1END[0]
+ Tile_X5Y0_NE_term/N1END[1] Tile_X5Y0_NE_term/N1END[2] Tile_X5Y0_NE_term/N1END[3]
+ Tile_X5Y0_NE_term/N2MID[0] Tile_X5Y0_NE_term/N2MID[1] Tile_X5Y0_NE_term/N2MID[2]
+ Tile_X5Y0_NE_term/N2MID[3] Tile_X5Y0_NE_term/N2MID[4] Tile_X5Y0_NE_term/N2MID[5]
+ Tile_X5Y0_NE_term/N2MID[6] Tile_X5Y0_NE_term/N2MID[7] Tile_X5Y0_NE_term/N2END[0]
+ Tile_X5Y0_NE_term/N2END[1] Tile_X5Y0_NE_term/N2END[2] Tile_X5Y0_NE_term/N2END[3]
+ Tile_X5Y0_NE_term/N2END[4] Tile_X5Y0_NE_term/N2END[5] Tile_X5Y0_NE_term/N2END[6]
+ Tile_X5Y0_NE_term/N2END[7] Tile_X5Y0_NE_term/N4END[0] Tile_X5Y0_NE_term/N4END[10]
+ Tile_X5Y0_NE_term/N4END[11] Tile_X5Y0_NE_term/N4END[12] Tile_X5Y0_NE_term/N4END[13]
+ Tile_X5Y0_NE_term/N4END[14] Tile_X5Y0_NE_term/N4END[15] Tile_X5Y0_NE_term/N4END[1]
+ Tile_X5Y0_NE_term/N4END[2] Tile_X5Y0_NE_term/N4END[3] Tile_X5Y0_NE_term/N4END[4]
+ Tile_X5Y0_NE_term/N4END[5] Tile_X5Y0_NE_term/N4END[6] Tile_X5Y0_NE_term/N4END[7]
+ Tile_X5Y0_NE_term/N4END[8] Tile_X5Y0_NE_term/N4END[9] Tile_X5Y0_NE_term/S1BEG[0]
+ Tile_X5Y0_NE_term/S1BEG[1] Tile_X5Y0_NE_term/S1BEG[2] Tile_X5Y0_NE_term/S1BEG[3]
+ Tile_X5Y0_NE_term/S2BEGb[0] Tile_X5Y0_NE_term/S2BEGb[1] Tile_X5Y0_NE_term/S2BEGb[2]
+ Tile_X5Y0_NE_term/S2BEGb[3] Tile_X5Y0_NE_term/S2BEGb[4] Tile_X5Y0_NE_term/S2BEGb[5]
+ Tile_X5Y0_NE_term/S2BEGb[6] Tile_X5Y0_NE_term/S2BEGb[7] Tile_X5Y0_NE_term/S2BEG[0]
+ Tile_X5Y0_NE_term/S2BEG[1] Tile_X5Y0_NE_term/S2BEG[2] Tile_X5Y0_NE_term/S2BEG[3]
+ Tile_X5Y0_NE_term/S2BEG[4] Tile_X5Y0_NE_term/S2BEG[5] Tile_X5Y0_NE_term/S2BEG[6]
+ Tile_X5Y0_NE_term/S2BEG[7] Tile_X5Y0_NE_term/S4BEG[0] Tile_X5Y0_NE_term/S4BEG[10]
+ Tile_X5Y0_NE_term/S4BEG[11] Tile_X5Y0_NE_term/S4BEG[12] Tile_X5Y0_NE_term/S4BEG[13]
+ Tile_X5Y0_NE_term/S4BEG[14] Tile_X5Y0_NE_term/S4BEG[15] Tile_X5Y0_NE_term/S4BEG[1]
+ Tile_X5Y0_NE_term/S4BEG[2] Tile_X5Y0_NE_term/S4BEG[3] Tile_X5Y0_NE_term/S4BEG[4]
+ Tile_X5Y0_NE_term/S4BEG[5] Tile_X5Y0_NE_term/S4BEG[6] Tile_X5Y0_NE_term/S4BEG[7]
+ Tile_X5Y0_NE_term/S4BEG[8] Tile_X5Y0_NE_term/S4BEG[9] Tile_X5Y0_NE_term/UserCLK
+ Tile_X4Y1_LUT4AB/W1END[0] Tile_X4Y1_LUT4AB/W1END[1] Tile_X4Y1_LUT4AB/W1END[2] Tile_X4Y1_LUT4AB/W1END[3]
+ Tile_X4Y1_LUT4AB/W2MID[0] Tile_X4Y1_LUT4AB/W2MID[1] Tile_X4Y1_LUT4AB/W2MID[2] Tile_X4Y1_LUT4AB/W2MID[3]
+ Tile_X4Y1_LUT4AB/W2MID[4] Tile_X4Y1_LUT4AB/W2MID[5] Tile_X4Y1_LUT4AB/W2MID[6] Tile_X4Y1_LUT4AB/W2MID[7]
+ Tile_X4Y1_LUT4AB/W2END[0] Tile_X4Y1_LUT4AB/W2END[1] Tile_X4Y1_LUT4AB/W2END[2] Tile_X4Y1_LUT4AB/W2END[3]
+ Tile_X4Y1_LUT4AB/W2END[4] Tile_X4Y1_LUT4AB/W2END[5] Tile_X4Y1_LUT4AB/W2END[6] Tile_X4Y1_LUT4AB/W2END[7]
+ Tile_X4Y1_LUT4AB/W6END[0] Tile_X4Y1_LUT4AB/W6END[10] Tile_X4Y1_LUT4AB/W6END[11]
+ Tile_X4Y1_LUT4AB/W6END[1] Tile_X4Y1_LUT4AB/W6END[2] Tile_X4Y1_LUT4AB/W6END[3] Tile_X4Y1_LUT4AB/W6END[4]
+ Tile_X4Y1_LUT4AB/W6END[5] Tile_X4Y1_LUT4AB/W6END[6] Tile_X4Y1_LUT4AB/W6END[7] Tile_X4Y1_LUT4AB/W6END[8]
+ Tile_X4Y1_LUT4AB/W6END[9] Tile_X4Y1_LUT4AB/WW4END[0] Tile_X4Y1_LUT4AB/WW4END[10]
+ Tile_X4Y1_LUT4AB/WW4END[11] Tile_X4Y1_LUT4AB/WW4END[12] Tile_X4Y1_LUT4AB/WW4END[13]
+ Tile_X4Y1_LUT4AB/WW4END[14] Tile_X4Y1_LUT4AB/WW4END[15] Tile_X4Y1_LUT4AB/WW4END[1]
+ Tile_X4Y1_LUT4AB/WW4END[2] Tile_X4Y1_LUT4AB/WW4END[3] Tile_X4Y1_LUT4AB/WW4END[4]
+ Tile_X4Y1_LUT4AB/WW4END[5] Tile_X4Y1_LUT4AB/WW4END[6] Tile_X4Y1_LUT4AB/WW4END[7]
+ Tile_X4Y1_LUT4AB/WW4END[8] Tile_X4Y1_LUT4AB/WW4END[9] Tile_X4Y2_LUT4AB/E1BEG[0]
+ Tile_X4Y2_LUT4AB/E1BEG[1] Tile_X4Y2_LUT4AB/E1BEG[2] Tile_X4Y2_LUT4AB/E1BEG[3] Tile_X4Y2_LUT4AB/E2BEGb[0]
+ Tile_X4Y2_LUT4AB/E2BEGb[1] Tile_X4Y2_LUT4AB/E2BEGb[2] Tile_X4Y2_LUT4AB/E2BEGb[3]
+ Tile_X4Y2_LUT4AB/E2BEGb[4] Tile_X4Y2_LUT4AB/E2BEGb[5] Tile_X4Y2_LUT4AB/E2BEGb[6]
+ Tile_X4Y2_LUT4AB/E2BEGb[7] Tile_X4Y2_LUT4AB/E2BEG[0] Tile_X4Y2_LUT4AB/E2BEG[1] Tile_X4Y2_LUT4AB/E2BEG[2]
+ Tile_X4Y2_LUT4AB/E2BEG[3] Tile_X4Y2_LUT4AB/E2BEG[4] Tile_X4Y2_LUT4AB/E2BEG[5] Tile_X4Y2_LUT4AB/E2BEG[6]
+ Tile_X4Y2_LUT4AB/E2BEG[7] Tile_X4Y2_LUT4AB/E6BEG[0] Tile_X4Y2_LUT4AB/E6BEG[10] Tile_X4Y2_LUT4AB/E6BEG[11]
+ Tile_X4Y2_LUT4AB/E6BEG[1] Tile_X4Y2_LUT4AB/E6BEG[2] Tile_X4Y2_LUT4AB/E6BEG[3] Tile_X4Y2_LUT4AB/E6BEG[4]
+ Tile_X4Y2_LUT4AB/E6BEG[5] Tile_X4Y2_LUT4AB/E6BEG[6] Tile_X4Y2_LUT4AB/E6BEG[7] Tile_X4Y2_LUT4AB/E6BEG[8]
+ Tile_X4Y2_LUT4AB/E6BEG[9] Tile_X4Y2_LUT4AB/EE4BEG[0] Tile_X4Y2_LUT4AB/EE4BEG[10]
+ Tile_X4Y2_LUT4AB/EE4BEG[11] Tile_X4Y2_LUT4AB/EE4BEG[12] Tile_X4Y2_LUT4AB/EE4BEG[13]
+ Tile_X4Y2_LUT4AB/EE4BEG[14] Tile_X4Y2_LUT4AB/EE4BEG[15] Tile_X4Y2_LUT4AB/EE4BEG[1]
+ Tile_X4Y2_LUT4AB/EE4BEG[2] Tile_X4Y2_LUT4AB/EE4BEG[3] Tile_X4Y2_LUT4AB/EE4BEG[4]
+ Tile_X4Y2_LUT4AB/EE4BEG[5] Tile_X4Y2_LUT4AB/EE4BEG[6] Tile_X4Y2_LUT4AB/EE4BEG[7]
+ Tile_X4Y2_LUT4AB/EE4BEG[8] Tile_X4Y2_LUT4AB/EE4BEG[9] Tile_X4Y2_LUT4AB/FrameData_O[0]
+ Tile_X4Y2_LUT4AB/FrameData_O[10] Tile_X4Y2_LUT4AB/FrameData_O[11] Tile_X4Y2_LUT4AB/FrameData_O[12]
+ Tile_X4Y2_LUT4AB/FrameData_O[13] Tile_X4Y2_LUT4AB/FrameData_O[14] Tile_X4Y2_LUT4AB/FrameData_O[15]
+ Tile_X4Y2_LUT4AB/FrameData_O[16] Tile_X4Y2_LUT4AB/FrameData_O[17] Tile_X4Y2_LUT4AB/FrameData_O[18]
+ Tile_X4Y2_LUT4AB/FrameData_O[19] Tile_X4Y2_LUT4AB/FrameData_O[1] Tile_X4Y2_LUT4AB/FrameData_O[20]
+ Tile_X4Y2_LUT4AB/FrameData_O[21] Tile_X4Y2_LUT4AB/FrameData_O[22] Tile_X4Y2_LUT4AB/FrameData_O[23]
+ Tile_X4Y2_LUT4AB/FrameData_O[24] Tile_X4Y2_LUT4AB/FrameData_O[25] Tile_X4Y2_LUT4AB/FrameData_O[26]
+ Tile_X4Y2_LUT4AB/FrameData_O[27] Tile_X4Y2_LUT4AB/FrameData_O[28] Tile_X4Y2_LUT4AB/FrameData_O[29]
+ Tile_X4Y2_LUT4AB/FrameData_O[2] Tile_X4Y2_LUT4AB/FrameData_O[30] Tile_X4Y2_LUT4AB/FrameData_O[31]
+ Tile_X4Y2_LUT4AB/FrameData_O[3] Tile_X4Y2_LUT4AB/FrameData_O[4] Tile_X4Y2_LUT4AB/FrameData_O[5]
+ Tile_X4Y2_LUT4AB/FrameData_O[6] Tile_X4Y2_LUT4AB/FrameData_O[7] Tile_X4Y2_LUT4AB/FrameData_O[8]
+ Tile_X4Y2_LUT4AB/FrameData_O[9] Tile_X5Y1_IHP_SRAM/Tile_X0Y1_FrameData_O[0] Tile_X5Y1_IHP_SRAM/Tile_X0Y1_FrameData_O[10]
+ Tile_X5Y1_IHP_SRAM/Tile_X0Y1_FrameData_O[11] Tile_X5Y1_IHP_SRAM/Tile_X0Y1_FrameData_O[12]
+ Tile_X5Y1_IHP_SRAM/Tile_X0Y1_FrameData_O[13] Tile_X5Y1_IHP_SRAM/Tile_X0Y1_FrameData_O[14]
+ Tile_X5Y1_IHP_SRAM/Tile_X0Y1_FrameData_O[15] Tile_X5Y1_IHP_SRAM/Tile_X0Y1_FrameData_O[16]
+ Tile_X5Y1_IHP_SRAM/Tile_X0Y1_FrameData_O[17] Tile_X5Y1_IHP_SRAM/Tile_X0Y1_FrameData_O[18]
+ Tile_X5Y1_IHP_SRAM/Tile_X0Y1_FrameData_O[19] Tile_X5Y1_IHP_SRAM/Tile_X0Y1_FrameData_O[1]
+ Tile_X5Y1_IHP_SRAM/Tile_X0Y1_FrameData_O[20] Tile_X5Y1_IHP_SRAM/Tile_X0Y1_FrameData_O[21]
+ Tile_X5Y1_IHP_SRAM/Tile_X0Y1_FrameData_O[22] Tile_X5Y1_IHP_SRAM/Tile_X0Y1_FrameData_O[23]
+ Tile_X5Y1_IHP_SRAM/Tile_X0Y1_FrameData_O[24] Tile_X5Y1_IHP_SRAM/Tile_X0Y1_FrameData_O[25]
+ Tile_X5Y1_IHP_SRAM/Tile_X0Y1_FrameData_O[26] Tile_X5Y1_IHP_SRAM/Tile_X0Y1_FrameData_O[27]
+ Tile_X5Y1_IHP_SRAM/Tile_X0Y1_FrameData_O[28] Tile_X5Y1_IHP_SRAM/Tile_X0Y1_FrameData_O[29]
+ Tile_X5Y1_IHP_SRAM/Tile_X0Y1_FrameData_O[2] Tile_X5Y1_IHP_SRAM/Tile_X0Y1_FrameData_O[30]
+ Tile_X5Y1_IHP_SRAM/Tile_X0Y1_FrameData_O[31] Tile_X5Y1_IHP_SRAM/Tile_X0Y1_FrameData_O[3]
+ Tile_X5Y1_IHP_SRAM/Tile_X0Y1_FrameData_O[4] Tile_X5Y1_IHP_SRAM/Tile_X0Y1_FrameData_O[5]
+ Tile_X5Y1_IHP_SRAM/Tile_X0Y1_FrameData_O[6] Tile_X5Y1_IHP_SRAM/Tile_X0Y1_FrameData_O[7]
+ Tile_X5Y1_IHP_SRAM/Tile_X0Y1_FrameData_O[8] Tile_X5Y1_IHP_SRAM/Tile_X0Y1_FrameData_O[9]
+ Tile_X5Y3_E_TT_IF/FrameStrobe_O[0] Tile_X5Y3_E_TT_IF/FrameStrobe_O[10] Tile_X5Y3_E_TT_IF/FrameStrobe_O[11]
+ Tile_X5Y3_E_TT_IF/FrameStrobe_O[12] Tile_X5Y3_E_TT_IF/FrameStrobe_O[13] Tile_X5Y3_E_TT_IF/FrameStrobe_O[14]
+ Tile_X5Y3_E_TT_IF/FrameStrobe_O[15] Tile_X5Y3_E_TT_IF/FrameStrobe_O[16] Tile_X5Y3_E_TT_IF/FrameStrobe_O[17]
+ Tile_X5Y3_E_TT_IF/FrameStrobe_O[18] Tile_X5Y3_E_TT_IF/FrameStrobe_O[19] Tile_X5Y3_E_TT_IF/FrameStrobe_O[1]
+ Tile_X5Y3_E_TT_IF/FrameStrobe_O[2] Tile_X5Y3_E_TT_IF/FrameStrobe_O[3] Tile_X5Y3_E_TT_IF/FrameStrobe_O[4]
+ Tile_X5Y3_E_TT_IF/FrameStrobe_O[5] Tile_X5Y3_E_TT_IF/FrameStrobe_O[6] Tile_X5Y3_E_TT_IF/FrameStrobe_O[7]
+ Tile_X5Y3_E_TT_IF/FrameStrobe_O[8] Tile_X5Y3_E_TT_IF/FrameStrobe_O[9] Tile_X5Y3_E_TT_IF/N1BEG[0]
+ Tile_X5Y3_E_TT_IF/N1BEG[1] Tile_X5Y3_E_TT_IF/N1BEG[2] Tile_X5Y3_E_TT_IF/N1BEG[3]
+ Tile_X5Y3_E_TT_IF/N2BEGb[0] Tile_X5Y3_E_TT_IF/N2BEGb[1] Tile_X5Y3_E_TT_IF/N2BEGb[2]
+ Tile_X5Y3_E_TT_IF/N2BEGb[3] Tile_X5Y3_E_TT_IF/N2BEGb[4] Tile_X5Y3_E_TT_IF/N2BEGb[5]
+ Tile_X5Y3_E_TT_IF/N2BEGb[6] Tile_X5Y3_E_TT_IF/N2BEGb[7] Tile_X5Y3_E_TT_IF/N2BEG[0]
+ Tile_X5Y3_E_TT_IF/N2BEG[1] Tile_X5Y3_E_TT_IF/N2BEG[2] Tile_X5Y3_E_TT_IF/N2BEG[3]
+ Tile_X5Y3_E_TT_IF/N2BEG[4] Tile_X5Y3_E_TT_IF/N2BEG[5] Tile_X5Y3_E_TT_IF/N2BEG[6]
+ Tile_X5Y3_E_TT_IF/N2BEG[7] Tile_X5Y3_E_TT_IF/N4BEG[0] Tile_X5Y3_E_TT_IF/N4BEG[10]
+ Tile_X5Y3_E_TT_IF/N4BEG[11] Tile_X5Y3_E_TT_IF/N4BEG[12] Tile_X5Y3_E_TT_IF/N4BEG[13]
+ Tile_X5Y3_E_TT_IF/N4BEG[14] Tile_X5Y3_E_TT_IF/N4BEG[15] Tile_X5Y3_E_TT_IF/N4BEG[1]
+ Tile_X5Y3_E_TT_IF/N4BEG[2] Tile_X5Y3_E_TT_IF/N4BEG[3] Tile_X5Y3_E_TT_IF/N4BEG[4]
+ Tile_X5Y3_E_TT_IF/N4BEG[5] Tile_X5Y3_E_TT_IF/N4BEG[6] Tile_X5Y3_E_TT_IF/N4BEG[7]
+ Tile_X5Y3_E_TT_IF/N4BEG[8] Tile_X5Y3_E_TT_IF/N4BEG[9] Tile_X5Y3_E_TT_IF/S1END[0]
+ Tile_X5Y3_E_TT_IF/S1END[1] Tile_X5Y3_E_TT_IF/S1END[2] Tile_X5Y3_E_TT_IF/S1END[3]
+ Tile_X5Y3_E_TT_IF/S2MID[0] Tile_X5Y3_E_TT_IF/S2MID[1] Tile_X5Y3_E_TT_IF/S2MID[2]
+ Tile_X5Y3_E_TT_IF/S2MID[3] Tile_X5Y3_E_TT_IF/S2MID[4] Tile_X5Y3_E_TT_IF/S2MID[5]
+ Tile_X5Y3_E_TT_IF/S2MID[6] Tile_X5Y3_E_TT_IF/S2MID[7] Tile_X5Y3_E_TT_IF/S2END[0]
+ Tile_X5Y3_E_TT_IF/S2END[1] Tile_X5Y3_E_TT_IF/S2END[2] Tile_X5Y3_E_TT_IF/S2END[3]
+ Tile_X5Y3_E_TT_IF/S2END[4] Tile_X5Y3_E_TT_IF/S2END[5] Tile_X5Y3_E_TT_IF/S2END[6]
+ Tile_X5Y3_E_TT_IF/S2END[7] Tile_X5Y3_E_TT_IF/S4END[0] Tile_X5Y3_E_TT_IF/S4END[10]
+ Tile_X5Y3_E_TT_IF/S4END[11] Tile_X5Y3_E_TT_IF/S4END[12] Tile_X5Y3_E_TT_IF/S4END[13]
+ Tile_X5Y3_E_TT_IF/S4END[14] Tile_X5Y3_E_TT_IF/S4END[15] Tile_X5Y3_E_TT_IF/S4END[1]
+ Tile_X5Y3_E_TT_IF/S4END[2] Tile_X5Y3_E_TT_IF/S4END[3] Tile_X5Y3_E_TT_IF/S4END[4]
+ Tile_X5Y3_E_TT_IF/S4END[5] Tile_X5Y3_E_TT_IF/S4END[6] Tile_X5Y3_E_TT_IF/S4END[7]
+ Tile_X5Y3_E_TT_IF/S4END[8] Tile_X5Y3_E_TT_IF/S4END[9] Tile_X5Y3_E_TT_IF/UserCLKo
+ Tile_X4Y2_LUT4AB/W1END[0] Tile_X4Y2_LUT4AB/W1END[1] Tile_X4Y2_LUT4AB/W1END[2] Tile_X4Y2_LUT4AB/W1END[3]
+ Tile_X4Y2_LUT4AB/W2MID[0] Tile_X4Y2_LUT4AB/W2MID[1] Tile_X4Y2_LUT4AB/W2MID[2] Tile_X4Y2_LUT4AB/W2MID[3]
+ Tile_X4Y2_LUT4AB/W2MID[4] Tile_X4Y2_LUT4AB/W2MID[5] Tile_X4Y2_LUT4AB/W2MID[6] Tile_X4Y2_LUT4AB/W2MID[7]
+ Tile_X4Y2_LUT4AB/W2END[0] Tile_X4Y2_LUT4AB/W2END[1] Tile_X4Y2_LUT4AB/W2END[2] Tile_X4Y2_LUT4AB/W2END[3]
+ Tile_X4Y2_LUT4AB/W2END[4] Tile_X4Y2_LUT4AB/W2END[5] Tile_X4Y2_LUT4AB/W2END[6] Tile_X4Y2_LUT4AB/W2END[7]
+ Tile_X4Y2_LUT4AB/W6END[0] Tile_X4Y2_LUT4AB/W6END[10] Tile_X4Y2_LUT4AB/W6END[11]
+ Tile_X4Y2_LUT4AB/W6END[1] Tile_X4Y2_LUT4AB/W6END[2] Tile_X4Y2_LUT4AB/W6END[3] Tile_X4Y2_LUT4AB/W6END[4]
+ Tile_X4Y2_LUT4AB/W6END[5] Tile_X4Y2_LUT4AB/W6END[6] Tile_X4Y2_LUT4AB/W6END[7] Tile_X4Y2_LUT4AB/W6END[8]
+ Tile_X4Y2_LUT4AB/W6END[9] Tile_X4Y2_LUT4AB/WW4END[0] Tile_X4Y2_LUT4AB/WW4END[10]
+ Tile_X4Y2_LUT4AB/WW4END[11] Tile_X4Y2_LUT4AB/WW4END[12] Tile_X4Y2_LUT4AB/WW4END[13]
+ Tile_X4Y2_LUT4AB/WW4END[14] Tile_X4Y2_LUT4AB/WW4END[15] Tile_X4Y2_LUT4AB/WW4END[1]
+ Tile_X4Y2_LUT4AB/WW4END[2] Tile_X4Y2_LUT4AB/WW4END[3] Tile_X4Y2_LUT4AB/WW4END[4]
+ Tile_X4Y2_LUT4AB/WW4END[5] Tile_X4Y2_LUT4AB/WW4END[6] Tile_X4Y2_LUT4AB/WW4END[7]
+ Tile_X4Y2_LUT4AB/WW4END[8] Tile_X4Y2_LUT4AB/WW4END[9] VGND VPWR Tile_X5Y2_WEN_SRAM
+ IHP_SRAM
XTile_X0Y1_W_TT_IF Tile_X0Y1_CLK_TT_PROJECT Tile_X1Y1_LUT4AB/E1END[0] Tile_X1Y1_LUT4AB/E1END[1]
+ Tile_X1Y1_LUT4AB/E1END[2] Tile_X1Y1_LUT4AB/E1END[3] Tile_X1Y1_LUT4AB/E2MID[0] Tile_X1Y1_LUT4AB/E2MID[1]
+ Tile_X1Y1_LUT4AB/E2MID[2] Tile_X1Y1_LUT4AB/E2MID[3] Tile_X1Y1_LUT4AB/E2MID[4] Tile_X1Y1_LUT4AB/E2MID[5]
+ Tile_X1Y1_LUT4AB/E2MID[6] Tile_X1Y1_LUT4AB/E2MID[7] Tile_X1Y1_LUT4AB/E2END[0] Tile_X1Y1_LUT4AB/E2END[1]
+ Tile_X1Y1_LUT4AB/E2END[2] Tile_X1Y1_LUT4AB/E2END[3] Tile_X1Y1_LUT4AB/E2END[4] Tile_X1Y1_LUT4AB/E2END[5]
+ Tile_X1Y1_LUT4AB/E2END[6] Tile_X1Y1_LUT4AB/E2END[7] Tile_X1Y1_LUT4AB/E6END[0] Tile_X1Y1_LUT4AB/E6END[10]
+ Tile_X1Y1_LUT4AB/E6END[11] Tile_X1Y1_LUT4AB/E6END[1] Tile_X1Y1_LUT4AB/E6END[2] Tile_X1Y1_LUT4AB/E6END[3]
+ Tile_X1Y1_LUT4AB/E6END[4] Tile_X1Y1_LUT4AB/E6END[5] Tile_X1Y1_LUT4AB/E6END[6] Tile_X1Y1_LUT4AB/E6END[7]
+ Tile_X1Y1_LUT4AB/E6END[8] Tile_X1Y1_LUT4AB/E6END[9] Tile_X1Y1_LUT4AB/EE4END[0] Tile_X1Y1_LUT4AB/EE4END[10]
+ Tile_X1Y1_LUT4AB/EE4END[11] Tile_X1Y1_LUT4AB/EE4END[12] Tile_X1Y1_LUT4AB/EE4END[13]
+ Tile_X1Y1_LUT4AB/EE4END[14] Tile_X1Y1_LUT4AB/EE4END[15] Tile_X1Y1_LUT4AB/EE4END[1]
+ Tile_X1Y1_LUT4AB/EE4END[2] Tile_X1Y1_LUT4AB/EE4END[3] Tile_X1Y1_LUT4AB/EE4END[4]
+ Tile_X1Y1_LUT4AB/EE4END[5] Tile_X1Y1_LUT4AB/EE4END[6] Tile_X1Y1_LUT4AB/EE4END[7]
+ Tile_X1Y1_LUT4AB/EE4END[8] Tile_X1Y1_LUT4AB/EE4END[9] Tile_X0Y1_ENA_TT_PROJECT FrameData[32]
+ FrameData[42] FrameData[43] FrameData[44] FrameData[45] FrameData[46] FrameData[47]
+ FrameData[48] FrameData[49] FrameData[50] FrameData[51] FrameData[33] FrameData[52]
+ FrameData[53] FrameData[54] FrameData[55] FrameData[56] FrameData[57] FrameData[58]
+ FrameData[59] FrameData[60] FrameData[61] FrameData[34] FrameData[62] FrameData[63]
+ FrameData[35] FrameData[36] FrameData[37] FrameData[38] FrameData[39] FrameData[40]
+ FrameData[41] Tile_X1Y1_LUT4AB/FrameData[0] Tile_X1Y1_LUT4AB/FrameData[10] Tile_X1Y1_LUT4AB/FrameData[11]
+ Tile_X1Y1_LUT4AB/FrameData[12] Tile_X1Y1_LUT4AB/FrameData[13] Tile_X1Y1_LUT4AB/FrameData[14]
+ Tile_X1Y1_LUT4AB/FrameData[15] Tile_X1Y1_LUT4AB/FrameData[16] Tile_X1Y1_LUT4AB/FrameData[17]
+ Tile_X1Y1_LUT4AB/FrameData[18] Tile_X1Y1_LUT4AB/FrameData[19] Tile_X1Y1_LUT4AB/FrameData[1]
+ Tile_X1Y1_LUT4AB/FrameData[20] Tile_X1Y1_LUT4AB/FrameData[21] Tile_X1Y1_LUT4AB/FrameData[22]
+ Tile_X1Y1_LUT4AB/FrameData[23] Tile_X1Y1_LUT4AB/FrameData[24] Tile_X1Y1_LUT4AB/FrameData[25]
+ Tile_X1Y1_LUT4AB/FrameData[26] Tile_X1Y1_LUT4AB/FrameData[27] Tile_X1Y1_LUT4AB/FrameData[28]
+ Tile_X1Y1_LUT4AB/FrameData[29] Tile_X1Y1_LUT4AB/FrameData[2] Tile_X1Y1_LUT4AB/FrameData[30]
+ Tile_X1Y1_LUT4AB/FrameData[31] Tile_X1Y1_LUT4AB/FrameData[3] Tile_X1Y1_LUT4AB/FrameData[4]
+ Tile_X1Y1_LUT4AB/FrameData[5] Tile_X1Y1_LUT4AB/FrameData[6] Tile_X1Y1_LUT4AB/FrameData[7]
+ Tile_X1Y1_LUT4AB/FrameData[8] Tile_X1Y1_LUT4AB/FrameData[9] Tile_X0Y1_W_TT_IF/FrameStrobe[0]
+ Tile_X0Y1_W_TT_IF/FrameStrobe[10] Tile_X0Y1_W_TT_IF/FrameStrobe[11] Tile_X0Y1_W_TT_IF/FrameStrobe[12]
+ Tile_X0Y1_W_TT_IF/FrameStrobe[13] Tile_X0Y1_W_TT_IF/FrameStrobe[14] Tile_X0Y1_W_TT_IF/FrameStrobe[15]
+ Tile_X0Y1_W_TT_IF/FrameStrobe[16] Tile_X0Y1_W_TT_IF/FrameStrobe[17] Tile_X0Y1_W_TT_IF/FrameStrobe[18]
+ Tile_X0Y1_W_TT_IF/FrameStrobe[19] Tile_X0Y1_W_TT_IF/FrameStrobe[1] Tile_X0Y1_W_TT_IF/FrameStrobe[2]
+ Tile_X0Y1_W_TT_IF/FrameStrobe[3] Tile_X0Y1_W_TT_IF/FrameStrobe[4] Tile_X0Y1_W_TT_IF/FrameStrobe[5]
+ Tile_X0Y1_W_TT_IF/FrameStrobe[6] Tile_X0Y1_W_TT_IF/FrameStrobe[7] Tile_X0Y1_W_TT_IF/FrameStrobe[8]
+ Tile_X0Y1_W_TT_IF/FrameStrobe[9] Tile_X0Y0_NW_term/FrameStrobe[0] Tile_X0Y0_NW_term/FrameStrobe[10]
+ Tile_X0Y0_NW_term/FrameStrobe[11] Tile_X0Y0_NW_term/FrameStrobe[12] Tile_X0Y0_NW_term/FrameStrobe[13]
+ Tile_X0Y0_NW_term/FrameStrobe[14] Tile_X0Y0_NW_term/FrameStrobe[15] Tile_X0Y0_NW_term/FrameStrobe[16]
+ Tile_X0Y0_NW_term/FrameStrobe[17] Tile_X0Y0_NW_term/FrameStrobe[18] Tile_X0Y0_NW_term/FrameStrobe[19]
+ Tile_X0Y0_NW_term/FrameStrobe[1] Tile_X0Y0_NW_term/FrameStrobe[2] Tile_X0Y0_NW_term/FrameStrobe[3]
+ Tile_X0Y0_NW_term/FrameStrobe[4] Tile_X0Y0_NW_term/FrameStrobe[5] Tile_X0Y0_NW_term/FrameStrobe[6]
+ Tile_X0Y0_NW_term/FrameStrobe[7] Tile_X0Y0_NW_term/FrameStrobe[8] Tile_X0Y0_NW_term/FrameStrobe[9]
+ Tile_X0Y1_W_TT_IF/N1BEG[0] Tile_X0Y1_W_TT_IF/N1BEG[1] Tile_X0Y1_W_TT_IF/N1BEG[2]
+ Tile_X0Y1_W_TT_IF/N1BEG[3] Tile_X0Y2_W_TT_IF/N1BEG[0] Tile_X0Y2_W_TT_IF/N1BEG[1]
+ Tile_X0Y2_W_TT_IF/N1BEG[2] Tile_X0Y2_W_TT_IF/N1BEG[3] Tile_X0Y1_W_TT_IF/N2BEG[0]
+ Tile_X0Y1_W_TT_IF/N2BEG[1] Tile_X0Y1_W_TT_IF/N2BEG[2] Tile_X0Y1_W_TT_IF/N2BEG[3]
+ Tile_X0Y1_W_TT_IF/N2BEG[4] Tile_X0Y1_W_TT_IF/N2BEG[5] Tile_X0Y1_W_TT_IF/N2BEG[6]
+ Tile_X0Y1_W_TT_IF/N2BEG[7] Tile_X0Y0_NW_term/N2END[0] Tile_X0Y0_NW_term/N2END[1]
+ Tile_X0Y0_NW_term/N2END[2] Tile_X0Y0_NW_term/N2END[3] Tile_X0Y0_NW_term/N2END[4]
+ Tile_X0Y0_NW_term/N2END[5] Tile_X0Y0_NW_term/N2END[6] Tile_X0Y0_NW_term/N2END[7]
+ Tile_X0Y1_W_TT_IF/N2END[0] Tile_X0Y1_W_TT_IF/N2END[1] Tile_X0Y1_W_TT_IF/N2END[2]
+ Tile_X0Y1_W_TT_IF/N2END[3] Tile_X0Y1_W_TT_IF/N2END[4] Tile_X0Y1_W_TT_IF/N2END[5]
+ Tile_X0Y1_W_TT_IF/N2END[6] Tile_X0Y1_W_TT_IF/N2END[7] Tile_X0Y2_W_TT_IF/N2BEG[0]
+ Tile_X0Y2_W_TT_IF/N2BEG[1] Tile_X0Y2_W_TT_IF/N2BEG[2] Tile_X0Y2_W_TT_IF/N2BEG[3]
+ Tile_X0Y2_W_TT_IF/N2BEG[4] Tile_X0Y2_W_TT_IF/N2BEG[5] Tile_X0Y2_W_TT_IF/N2BEG[6]
+ Tile_X0Y2_W_TT_IF/N2BEG[7] Tile_X0Y1_W_TT_IF/N4BEG[0] Tile_X0Y1_W_TT_IF/N4BEG[10]
+ Tile_X0Y1_W_TT_IF/N4BEG[11] Tile_X0Y1_W_TT_IF/N4BEG[12] Tile_X0Y1_W_TT_IF/N4BEG[13]
+ Tile_X0Y1_W_TT_IF/N4BEG[14] Tile_X0Y1_W_TT_IF/N4BEG[15] Tile_X0Y1_W_TT_IF/N4BEG[1]
+ Tile_X0Y1_W_TT_IF/N4BEG[2] Tile_X0Y1_W_TT_IF/N4BEG[3] Tile_X0Y1_W_TT_IF/N4BEG[4]
+ Tile_X0Y1_W_TT_IF/N4BEG[5] Tile_X0Y1_W_TT_IF/N4BEG[6] Tile_X0Y1_W_TT_IF/N4BEG[7]
+ Tile_X0Y1_W_TT_IF/N4BEG[8] Tile_X0Y1_W_TT_IF/N4BEG[9] Tile_X0Y2_W_TT_IF/N4BEG[0]
+ Tile_X0Y2_W_TT_IF/N4BEG[10] Tile_X0Y2_W_TT_IF/N4BEG[11] Tile_X0Y2_W_TT_IF/N4BEG[12]
+ Tile_X0Y2_W_TT_IF/N4BEG[13] Tile_X0Y2_W_TT_IF/N4BEG[14] Tile_X0Y2_W_TT_IF/N4BEG[15]
+ Tile_X0Y2_W_TT_IF/N4BEG[1] Tile_X0Y2_W_TT_IF/N4BEG[2] Tile_X0Y2_W_TT_IF/N4BEG[3]
+ Tile_X0Y2_W_TT_IF/N4BEG[4] Tile_X0Y2_W_TT_IF/N4BEG[5] Tile_X0Y2_W_TT_IF/N4BEG[6]
+ Tile_X0Y2_W_TT_IF/N4BEG[7] Tile_X0Y2_W_TT_IF/N4BEG[8] Tile_X0Y2_W_TT_IF/N4BEG[9]
+ Tile_X0Y1_RST_N_TT_PROJECT Tile_X0Y2_W_TT_IF/S1END[0] Tile_X0Y2_W_TT_IF/S1END[1]
+ Tile_X0Y2_W_TT_IF/S1END[2] Tile_X0Y2_W_TT_IF/S1END[3] Tile_X0Y1_W_TT_IF/S1END[0]
+ Tile_X0Y1_W_TT_IF/S1END[1] Tile_X0Y1_W_TT_IF/S1END[2] Tile_X0Y1_W_TT_IF/S1END[3]
+ Tile_X0Y2_W_TT_IF/S2MID[0] Tile_X0Y2_W_TT_IF/S2MID[1] Tile_X0Y2_W_TT_IF/S2MID[2]
+ Tile_X0Y2_W_TT_IF/S2MID[3] Tile_X0Y2_W_TT_IF/S2MID[4] Tile_X0Y2_W_TT_IF/S2MID[5]
+ Tile_X0Y2_W_TT_IF/S2MID[6] Tile_X0Y2_W_TT_IF/S2MID[7] Tile_X0Y2_W_TT_IF/S2END[0]
+ Tile_X0Y2_W_TT_IF/S2END[1] Tile_X0Y2_W_TT_IF/S2END[2] Tile_X0Y2_W_TT_IF/S2END[3]
+ Tile_X0Y2_W_TT_IF/S2END[4] Tile_X0Y2_W_TT_IF/S2END[5] Tile_X0Y2_W_TT_IF/S2END[6]
+ Tile_X0Y2_W_TT_IF/S2END[7] Tile_X0Y1_W_TT_IF/S2END[0] Tile_X0Y1_W_TT_IF/S2END[1]
+ Tile_X0Y1_W_TT_IF/S2END[2] Tile_X0Y1_W_TT_IF/S2END[3] Tile_X0Y1_W_TT_IF/S2END[4]
+ Tile_X0Y1_W_TT_IF/S2END[5] Tile_X0Y1_W_TT_IF/S2END[6] Tile_X0Y1_W_TT_IF/S2END[7]
+ Tile_X0Y1_W_TT_IF/S2MID[0] Tile_X0Y1_W_TT_IF/S2MID[1] Tile_X0Y1_W_TT_IF/S2MID[2]
+ Tile_X0Y1_W_TT_IF/S2MID[3] Tile_X0Y1_W_TT_IF/S2MID[4] Tile_X0Y1_W_TT_IF/S2MID[5]
+ Tile_X0Y1_W_TT_IF/S2MID[6] Tile_X0Y1_W_TT_IF/S2MID[7] Tile_X0Y2_W_TT_IF/S4END[0]
+ Tile_X0Y2_W_TT_IF/S4END[10] Tile_X0Y2_W_TT_IF/S4END[11] Tile_X0Y2_W_TT_IF/S4END[12]
+ Tile_X0Y2_W_TT_IF/S4END[13] Tile_X0Y2_W_TT_IF/S4END[14] Tile_X0Y2_W_TT_IF/S4END[15]
+ Tile_X0Y2_W_TT_IF/S4END[1] Tile_X0Y2_W_TT_IF/S4END[2] Tile_X0Y2_W_TT_IF/S4END[3]
+ Tile_X0Y2_W_TT_IF/S4END[4] Tile_X0Y2_W_TT_IF/S4END[5] Tile_X0Y2_W_TT_IF/S4END[6]
+ Tile_X0Y2_W_TT_IF/S4END[7] Tile_X0Y2_W_TT_IF/S4END[8] Tile_X0Y2_W_TT_IF/S4END[9]
+ Tile_X0Y1_W_TT_IF/S4END[0] Tile_X0Y1_W_TT_IF/S4END[10] Tile_X0Y1_W_TT_IF/S4END[11]
+ Tile_X0Y1_W_TT_IF/S4END[12] Tile_X0Y1_W_TT_IF/S4END[13] Tile_X0Y1_W_TT_IF/S4END[14]
+ Tile_X0Y1_W_TT_IF/S4END[15] Tile_X0Y1_W_TT_IF/S4END[1] Tile_X0Y1_W_TT_IF/S4END[2]
+ Tile_X0Y1_W_TT_IF/S4END[3] Tile_X0Y1_W_TT_IF/S4END[4] Tile_X0Y1_W_TT_IF/S4END[5]
+ Tile_X0Y1_W_TT_IF/S4END[6] Tile_X0Y1_W_TT_IF/S4END[7] Tile_X0Y1_W_TT_IF/S4END[8]
+ Tile_X0Y1_W_TT_IF/S4END[9] Tile_X0Y1_UIO_IN_TT_PROJECT0 Tile_X0Y1_UIO_IN_TT_PROJECT1
+ Tile_X0Y1_UIO_IN_TT_PROJECT2 Tile_X0Y1_UIO_IN_TT_PROJECT3 Tile_X0Y1_UIO_IN_TT_PROJECT4
+ Tile_X0Y1_UIO_IN_TT_PROJECT5 Tile_X0Y1_UIO_IN_TT_PROJECT6 Tile_X0Y1_UIO_IN_TT_PROJECT7
+ Tile_X0Y1_UIO_OE_TT_PROJECT0 Tile_X0Y1_UIO_OE_TT_PROJECT1 Tile_X0Y1_UIO_OE_TT_PROJECT2
+ Tile_X0Y1_UIO_OE_TT_PROJECT3 Tile_X0Y1_UIO_OE_TT_PROJECT4 Tile_X0Y1_UIO_OE_TT_PROJECT5
+ Tile_X0Y1_UIO_OE_TT_PROJECT6 Tile_X0Y1_UIO_OE_TT_PROJECT7 Tile_X0Y1_UIO_OUT_TT_PROJECT0
+ Tile_X0Y1_UIO_OUT_TT_PROJECT1 Tile_X0Y1_UIO_OUT_TT_PROJECT2 Tile_X0Y1_UIO_OUT_TT_PROJECT3
+ Tile_X0Y1_UIO_OUT_TT_PROJECT4 Tile_X0Y1_UIO_OUT_TT_PROJECT5 Tile_X0Y1_UIO_OUT_TT_PROJECT6
+ Tile_X0Y1_UIO_OUT_TT_PROJECT7 Tile_X0Y1_UI_IN_TT_PROJECT0 Tile_X0Y1_UI_IN_TT_PROJECT1
+ Tile_X0Y1_UI_IN_TT_PROJECT2 Tile_X0Y1_UI_IN_TT_PROJECT3 Tile_X0Y1_UI_IN_TT_PROJECT4
+ Tile_X0Y1_UI_IN_TT_PROJECT5 Tile_X0Y1_UI_IN_TT_PROJECT6 Tile_X0Y1_UI_IN_TT_PROJECT7
+ Tile_X0Y1_UO_OUT_TT_PROJECT0 Tile_X0Y1_UO_OUT_TT_PROJECT1 Tile_X0Y1_UO_OUT_TT_PROJECT2
+ Tile_X0Y1_UO_OUT_TT_PROJECT3 Tile_X0Y1_UO_OUT_TT_PROJECT4 Tile_X0Y1_UO_OUT_TT_PROJECT5
+ Tile_X0Y1_UO_OUT_TT_PROJECT6 Tile_X0Y1_UO_OUT_TT_PROJECT7 Tile_X0Y1_W_TT_IF/UserCLK
+ Tile_X0Y0_NW_term/UserCLK VGND VPWR Tile_X1Y1_LUT4AB/W1BEG[0] Tile_X1Y1_LUT4AB/W1BEG[1]
+ Tile_X1Y1_LUT4AB/W1BEG[2] Tile_X1Y1_LUT4AB/W1BEG[3] Tile_X1Y1_LUT4AB/W2BEGb[0] Tile_X1Y1_LUT4AB/W2BEGb[1]
+ Tile_X1Y1_LUT4AB/W2BEGb[2] Tile_X1Y1_LUT4AB/W2BEGb[3] Tile_X1Y1_LUT4AB/W2BEGb[4]
+ Tile_X1Y1_LUT4AB/W2BEGb[5] Tile_X1Y1_LUT4AB/W2BEGb[6] Tile_X1Y1_LUT4AB/W2BEGb[7]
+ Tile_X1Y1_LUT4AB/W2BEG[0] Tile_X1Y1_LUT4AB/W2BEG[1] Tile_X1Y1_LUT4AB/W2BEG[2] Tile_X1Y1_LUT4AB/W2BEG[3]
+ Tile_X1Y1_LUT4AB/W2BEG[4] Tile_X1Y1_LUT4AB/W2BEG[5] Tile_X1Y1_LUT4AB/W2BEG[6] Tile_X1Y1_LUT4AB/W2BEG[7]
+ Tile_X1Y1_LUT4AB/W6BEG[0] Tile_X1Y1_LUT4AB/W6BEG[10] Tile_X1Y1_LUT4AB/W6BEG[11]
+ Tile_X1Y1_LUT4AB/W6BEG[1] Tile_X1Y1_LUT4AB/W6BEG[2] Tile_X1Y1_LUT4AB/W6BEG[3] Tile_X1Y1_LUT4AB/W6BEG[4]
+ Tile_X1Y1_LUT4AB/W6BEG[5] Tile_X1Y1_LUT4AB/W6BEG[6] Tile_X1Y1_LUT4AB/W6BEG[7] Tile_X1Y1_LUT4AB/W6BEG[8]
+ Tile_X1Y1_LUT4AB/W6BEG[9] Tile_X1Y1_LUT4AB/WW4BEG[0] Tile_X1Y1_LUT4AB/WW4BEG[10]
+ Tile_X1Y1_LUT4AB/WW4BEG[11] Tile_X1Y1_LUT4AB/WW4BEG[12] Tile_X1Y1_LUT4AB/WW4BEG[13]
+ Tile_X1Y1_LUT4AB/WW4BEG[14] Tile_X1Y1_LUT4AB/WW4BEG[15] Tile_X1Y1_LUT4AB/WW4BEG[1]
+ Tile_X1Y1_LUT4AB/WW4BEG[2] Tile_X1Y1_LUT4AB/WW4BEG[3] Tile_X1Y1_LUT4AB/WW4BEG[4]
+ Tile_X1Y1_LUT4AB/WW4BEG[5] Tile_X1Y1_LUT4AB/WW4BEG[6] Tile_X1Y1_LUT4AB/WW4BEG[7]
+ Tile_X1Y1_LUT4AB/WW4BEG[8] Tile_X1Y1_LUT4AB/WW4BEG[9] W_TT_IF
XTile_X2Y3_LUT4AB Tile_X2Y4_LUT4AB/Co Tile_X2Y3_LUT4AB/Co Tile_X3Y3_LUT4AB/E1END[0]
+ Tile_X3Y3_LUT4AB/E1END[1] Tile_X3Y3_LUT4AB/E1END[2] Tile_X3Y3_LUT4AB/E1END[3] Tile_X2Y3_LUT4AB/E1END[0]
+ Tile_X2Y3_LUT4AB/E1END[1] Tile_X2Y3_LUT4AB/E1END[2] Tile_X2Y3_LUT4AB/E1END[3] Tile_X3Y3_LUT4AB/E2MID[0]
+ Tile_X3Y3_LUT4AB/E2MID[1] Tile_X3Y3_LUT4AB/E2MID[2] Tile_X3Y3_LUT4AB/E2MID[3] Tile_X3Y3_LUT4AB/E2MID[4]
+ Tile_X3Y3_LUT4AB/E2MID[5] Tile_X3Y3_LUT4AB/E2MID[6] Tile_X3Y3_LUT4AB/E2MID[7] Tile_X3Y3_LUT4AB/E2END[0]
+ Tile_X3Y3_LUT4AB/E2END[1] Tile_X3Y3_LUT4AB/E2END[2] Tile_X3Y3_LUT4AB/E2END[3] Tile_X3Y3_LUT4AB/E2END[4]
+ Tile_X3Y3_LUT4AB/E2END[5] Tile_X3Y3_LUT4AB/E2END[6] Tile_X3Y3_LUT4AB/E2END[7] Tile_X2Y3_LUT4AB/E2END[0]
+ Tile_X2Y3_LUT4AB/E2END[1] Tile_X2Y3_LUT4AB/E2END[2] Tile_X2Y3_LUT4AB/E2END[3] Tile_X2Y3_LUT4AB/E2END[4]
+ Tile_X2Y3_LUT4AB/E2END[5] Tile_X2Y3_LUT4AB/E2END[6] Tile_X2Y3_LUT4AB/E2END[7] Tile_X2Y3_LUT4AB/E2MID[0]
+ Tile_X2Y3_LUT4AB/E2MID[1] Tile_X2Y3_LUT4AB/E2MID[2] Tile_X2Y3_LUT4AB/E2MID[3] Tile_X2Y3_LUT4AB/E2MID[4]
+ Tile_X2Y3_LUT4AB/E2MID[5] Tile_X2Y3_LUT4AB/E2MID[6] Tile_X2Y3_LUT4AB/E2MID[7] Tile_X3Y3_LUT4AB/E6END[0]
+ Tile_X3Y3_LUT4AB/E6END[10] Tile_X3Y3_LUT4AB/E6END[11] Tile_X3Y3_LUT4AB/E6END[1]
+ Tile_X3Y3_LUT4AB/E6END[2] Tile_X3Y3_LUT4AB/E6END[3] Tile_X3Y3_LUT4AB/E6END[4] Tile_X3Y3_LUT4AB/E6END[5]
+ Tile_X3Y3_LUT4AB/E6END[6] Tile_X3Y3_LUT4AB/E6END[7] Tile_X3Y3_LUT4AB/E6END[8] Tile_X3Y3_LUT4AB/E6END[9]
+ Tile_X2Y3_LUT4AB/E6END[0] Tile_X2Y3_LUT4AB/E6END[10] Tile_X2Y3_LUT4AB/E6END[11]
+ Tile_X2Y3_LUT4AB/E6END[1] Tile_X2Y3_LUT4AB/E6END[2] Tile_X2Y3_LUT4AB/E6END[3] Tile_X2Y3_LUT4AB/E6END[4]
+ Tile_X2Y3_LUT4AB/E6END[5] Tile_X2Y3_LUT4AB/E6END[6] Tile_X2Y3_LUT4AB/E6END[7] Tile_X2Y3_LUT4AB/E6END[8]
+ Tile_X2Y3_LUT4AB/E6END[9] Tile_X3Y3_LUT4AB/EE4END[0] Tile_X3Y3_LUT4AB/EE4END[10]
+ Tile_X3Y3_LUT4AB/EE4END[11] Tile_X3Y3_LUT4AB/EE4END[12] Tile_X3Y3_LUT4AB/EE4END[13]
+ Tile_X3Y3_LUT4AB/EE4END[14] Tile_X3Y3_LUT4AB/EE4END[15] Tile_X3Y3_LUT4AB/EE4END[1]
+ Tile_X3Y3_LUT4AB/EE4END[2] Tile_X3Y3_LUT4AB/EE4END[3] Tile_X3Y3_LUT4AB/EE4END[4]
+ Tile_X3Y3_LUT4AB/EE4END[5] Tile_X3Y3_LUT4AB/EE4END[6] Tile_X3Y3_LUT4AB/EE4END[7]
+ Tile_X3Y3_LUT4AB/EE4END[8] Tile_X3Y3_LUT4AB/EE4END[9] Tile_X2Y3_LUT4AB/EE4END[0]
+ Tile_X2Y3_LUT4AB/EE4END[10] Tile_X2Y3_LUT4AB/EE4END[11] Tile_X2Y3_LUT4AB/EE4END[12]
+ Tile_X2Y3_LUT4AB/EE4END[13] Tile_X2Y3_LUT4AB/EE4END[14] Tile_X2Y3_LUT4AB/EE4END[15]
+ Tile_X2Y3_LUT4AB/EE4END[1] Tile_X2Y3_LUT4AB/EE4END[2] Tile_X2Y3_LUT4AB/EE4END[3]
+ Tile_X2Y3_LUT4AB/EE4END[4] Tile_X2Y3_LUT4AB/EE4END[5] Tile_X2Y3_LUT4AB/EE4END[6]
+ Tile_X2Y3_LUT4AB/EE4END[7] Tile_X2Y3_LUT4AB/EE4END[8] Tile_X2Y3_LUT4AB/EE4END[9]
+ Tile_X2Y3_LUT4AB/FrameData[0] Tile_X2Y3_LUT4AB/FrameData[10] Tile_X2Y3_LUT4AB/FrameData[11]
+ Tile_X2Y3_LUT4AB/FrameData[12] Tile_X2Y3_LUT4AB/FrameData[13] Tile_X2Y3_LUT4AB/FrameData[14]
+ Tile_X2Y3_LUT4AB/FrameData[15] Tile_X2Y3_LUT4AB/FrameData[16] Tile_X2Y3_LUT4AB/FrameData[17]
+ Tile_X2Y3_LUT4AB/FrameData[18] Tile_X2Y3_LUT4AB/FrameData[19] Tile_X2Y3_LUT4AB/FrameData[1]
+ Tile_X2Y3_LUT4AB/FrameData[20] Tile_X2Y3_LUT4AB/FrameData[21] Tile_X2Y3_LUT4AB/FrameData[22]
+ Tile_X2Y3_LUT4AB/FrameData[23] Tile_X2Y3_LUT4AB/FrameData[24] Tile_X2Y3_LUT4AB/FrameData[25]
+ Tile_X2Y3_LUT4AB/FrameData[26] Tile_X2Y3_LUT4AB/FrameData[27] Tile_X2Y3_LUT4AB/FrameData[28]
+ Tile_X2Y3_LUT4AB/FrameData[29] Tile_X2Y3_LUT4AB/FrameData[2] Tile_X2Y3_LUT4AB/FrameData[30]
+ Tile_X2Y3_LUT4AB/FrameData[31] Tile_X2Y3_LUT4AB/FrameData[3] Tile_X2Y3_LUT4AB/FrameData[4]
+ Tile_X2Y3_LUT4AB/FrameData[5] Tile_X2Y3_LUT4AB/FrameData[6] Tile_X2Y3_LUT4AB/FrameData[7]
+ Tile_X2Y3_LUT4AB/FrameData[8] Tile_X2Y3_LUT4AB/FrameData[9] Tile_X3Y3_LUT4AB/FrameData[0]
+ Tile_X3Y3_LUT4AB/FrameData[10] Tile_X3Y3_LUT4AB/FrameData[11] Tile_X3Y3_LUT4AB/FrameData[12]
+ Tile_X3Y3_LUT4AB/FrameData[13] Tile_X3Y3_LUT4AB/FrameData[14] Tile_X3Y3_LUT4AB/FrameData[15]
+ Tile_X3Y3_LUT4AB/FrameData[16] Tile_X3Y3_LUT4AB/FrameData[17] Tile_X3Y3_LUT4AB/FrameData[18]
+ Tile_X3Y3_LUT4AB/FrameData[19] Tile_X3Y3_LUT4AB/FrameData[1] Tile_X3Y3_LUT4AB/FrameData[20]
+ Tile_X3Y3_LUT4AB/FrameData[21] Tile_X3Y3_LUT4AB/FrameData[22] Tile_X3Y3_LUT4AB/FrameData[23]
+ Tile_X3Y3_LUT4AB/FrameData[24] Tile_X3Y3_LUT4AB/FrameData[25] Tile_X3Y3_LUT4AB/FrameData[26]
+ Tile_X3Y3_LUT4AB/FrameData[27] Tile_X3Y3_LUT4AB/FrameData[28] Tile_X3Y3_LUT4AB/FrameData[29]
+ Tile_X3Y3_LUT4AB/FrameData[2] Tile_X3Y3_LUT4AB/FrameData[30] Tile_X3Y3_LUT4AB/FrameData[31]
+ Tile_X3Y3_LUT4AB/FrameData[3] Tile_X3Y3_LUT4AB/FrameData[4] Tile_X3Y3_LUT4AB/FrameData[5]
+ Tile_X3Y3_LUT4AB/FrameData[6] Tile_X3Y3_LUT4AB/FrameData[7] Tile_X3Y3_LUT4AB/FrameData[8]
+ Tile_X3Y3_LUT4AB/FrameData[9] Tile_X2Y3_LUT4AB/FrameStrobe[0] Tile_X2Y3_LUT4AB/FrameStrobe[10]
+ Tile_X2Y3_LUT4AB/FrameStrobe[11] Tile_X2Y3_LUT4AB/FrameStrobe[12] Tile_X2Y3_LUT4AB/FrameStrobe[13]
+ Tile_X2Y3_LUT4AB/FrameStrobe[14] Tile_X2Y3_LUT4AB/FrameStrobe[15] Tile_X2Y3_LUT4AB/FrameStrobe[16]
+ Tile_X2Y3_LUT4AB/FrameStrobe[17] Tile_X2Y3_LUT4AB/FrameStrobe[18] Tile_X2Y3_LUT4AB/FrameStrobe[19]
+ Tile_X2Y3_LUT4AB/FrameStrobe[1] Tile_X2Y3_LUT4AB/FrameStrobe[2] Tile_X2Y3_LUT4AB/FrameStrobe[3]
+ Tile_X2Y3_LUT4AB/FrameStrobe[4] Tile_X2Y3_LUT4AB/FrameStrobe[5] Tile_X2Y3_LUT4AB/FrameStrobe[6]
+ Tile_X2Y3_LUT4AB/FrameStrobe[7] Tile_X2Y3_LUT4AB/FrameStrobe[8] Tile_X2Y3_LUT4AB/FrameStrobe[9]
+ Tile_X2Y2_LUT4AB/FrameStrobe[0] Tile_X2Y2_LUT4AB/FrameStrobe[10] Tile_X2Y2_LUT4AB/FrameStrobe[11]
+ Tile_X2Y2_LUT4AB/FrameStrobe[12] Tile_X2Y2_LUT4AB/FrameStrobe[13] Tile_X2Y2_LUT4AB/FrameStrobe[14]
+ Tile_X2Y2_LUT4AB/FrameStrobe[15] Tile_X2Y2_LUT4AB/FrameStrobe[16] Tile_X2Y2_LUT4AB/FrameStrobe[17]
+ Tile_X2Y2_LUT4AB/FrameStrobe[18] Tile_X2Y2_LUT4AB/FrameStrobe[19] Tile_X2Y2_LUT4AB/FrameStrobe[1]
+ Tile_X2Y2_LUT4AB/FrameStrobe[2] Tile_X2Y2_LUT4AB/FrameStrobe[3] Tile_X2Y2_LUT4AB/FrameStrobe[4]
+ Tile_X2Y2_LUT4AB/FrameStrobe[5] Tile_X2Y2_LUT4AB/FrameStrobe[6] Tile_X2Y2_LUT4AB/FrameStrobe[7]
+ Tile_X2Y2_LUT4AB/FrameStrobe[8] Tile_X2Y2_LUT4AB/FrameStrobe[9] Tile_X2Y3_LUT4AB/N1BEG[0]
+ Tile_X2Y3_LUT4AB/N1BEG[1] Tile_X2Y3_LUT4AB/N1BEG[2] Tile_X2Y3_LUT4AB/N1BEG[3] Tile_X2Y4_LUT4AB/N1BEG[0]
+ Tile_X2Y4_LUT4AB/N1BEG[1] Tile_X2Y4_LUT4AB/N1BEG[2] Tile_X2Y4_LUT4AB/N1BEG[3] Tile_X2Y3_LUT4AB/N2BEG[0]
+ Tile_X2Y3_LUT4AB/N2BEG[1] Tile_X2Y3_LUT4AB/N2BEG[2] Tile_X2Y3_LUT4AB/N2BEG[3] Tile_X2Y3_LUT4AB/N2BEG[4]
+ Tile_X2Y3_LUT4AB/N2BEG[5] Tile_X2Y3_LUT4AB/N2BEG[6] Tile_X2Y3_LUT4AB/N2BEG[7] Tile_X2Y2_LUT4AB/N2END[0]
+ Tile_X2Y2_LUT4AB/N2END[1] Tile_X2Y2_LUT4AB/N2END[2] Tile_X2Y2_LUT4AB/N2END[3] Tile_X2Y2_LUT4AB/N2END[4]
+ Tile_X2Y2_LUT4AB/N2END[5] Tile_X2Y2_LUT4AB/N2END[6] Tile_X2Y2_LUT4AB/N2END[7] Tile_X2Y3_LUT4AB/N2END[0]
+ Tile_X2Y3_LUT4AB/N2END[1] Tile_X2Y3_LUT4AB/N2END[2] Tile_X2Y3_LUT4AB/N2END[3] Tile_X2Y3_LUT4AB/N2END[4]
+ Tile_X2Y3_LUT4AB/N2END[5] Tile_X2Y3_LUT4AB/N2END[6] Tile_X2Y3_LUT4AB/N2END[7] Tile_X2Y4_LUT4AB/N2BEG[0]
+ Tile_X2Y4_LUT4AB/N2BEG[1] Tile_X2Y4_LUT4AB/N2BEG[2] Tile_X2Y4_LUT4AB/N2BEG[3] Tile_X2Y4_LUT4AB/N2BEG[4]
+ Tile_X2Y4_LUT4AB/N2BEG[5] Tile_X2Y4_LUT4AB/N2BEG[6] Tile_X2Y4_LUT4AB/N2BEG[7] Tile_X2Y3_LUT4AB/N4BEG[0]
+ Tile_X2Y3_LUT4AB/N4BEG[10] Tile_X2Y3_LUT4AB/N4BEG[11] Tile_X2Y3_LUT4AB/N4BEG[12]
+ Tile_X2Y3_LUT4AB/N4BEG[13] Tile_X2Y3_LUT4AB/N4BEG[14] Tile_X2Y3_LUT4AB/N4BEG[15]
+ Tile_X2Y3_LUT4AB/N4BEG[1] Tile_X2Y3_LUT4AB/N4BEG[2] Tile_X2Y3_LUT4AB/N4BEG[3] Tile_X2Y3_LUT4AB/N4BEG[4]
+ Tile_X2Y3_LUT4AB/N4BEG[5] Tile_X2Y3_LUT4AB/N4BEG[6] Tile_X2Y3_LUT4AB/N4BEG[7] Tile_X2Y3_LUT4AB/N4BEG[8]
+ Tile_X2Y3_LUT4AB/N4BEG[9] Tile_X2Y4_LUT4AB/N4BEG[0] Tile_X2Y4_LUT4AB/N4BEG[10] Tile_X2Y4_LUT4AB/N4BEG[11]
+ Tile_X2Y4_LUT4AB/N4BEG[12] Tile_X2Y4_LUT4AB/N4BEG[13] Tile_X2Y4_LUT4AB/N4BEG[14]
+ Tile_X2Y4_LUT4AB/N4BEG[15] Tile_X2Y4_LUT4AB/N4BEG[1] Tile_X2Y4_LUT4AB/N4BEG[2] Tile_X2Y4_LUT4AB/N4BEG[3]
+ Tile_X2Y4_LUT4AB/N4BEG[4] Tile_X2Y4_LUT4AB/N4BEG[5] Tile_X2Y4_LUT4AB/N4BEG[6] Tile_X2Y4_LUT4AB/N4BEG[7]
+ Tile_X2Y4_LUT4AB/N4BEG[8] Tile_X2Y4_LUT4AB/N4BEG[9] Tile_X2Y3_LUT4AB/NN4BEG[0] Tile_X2Y3_LUT4AB/NN4BEG[10]
+ Tile_X2Y3_LUT4AB/NN4BEG[11] Tile_X2Y3_LUT4AB/NN4BEG[12] Tile_X2Y3_LUT4AB/NN4BEG[13]
+ Tile_X2Y3_LUT4AB/NN4BEG[14] Tile_X2Y3_LUT4AB/NN4BEG[15] Tile_X2Y3_LUT4AB/NN4BEG[1]
+ Tile_X2Y3_LUT4AB/NN4BEG[2] Tile_X2Y3_LUT4AB/NN4BEG[3] Tile_X2Y3_LUT4AB/NN4BEG[4]
+ Tile_X2Y3_LUT4AB/NN4BEG[5] Tile_X2Y3_LUT4AB/NN4BEG[6] Tile_X2Y3_LUT4AB/NN4BEG[7]
+ Tile_X2Y3_LUT4AB/NN4BEG[8] Tile_X2Y3_LUT4AB/NN4BEG[9] Tile_X2Y4_LUT4AB/NN4BEG[0]
+ Tile_X2Y4_LUT4AB/NN4BEG[10] Tile_X2Y4_LUT4AB/NN4BEG[11] Tile_X2Y4_LUT4AB/NN4BEG[12]
+ Tile_X2Y4_LUT4AB/NN4BEG[13] Tile_X2Y4_LUT4AB/NN4BEG[14] Tile_X2Y4_LUT4AB/NN4BEG[15]
+ Tile_X2Y4_LUT4AB/NN4BEG[1] Tile_X2Y4_LUT4AB/NN4BEG[2] Tile_X2Y4_LUT4AB/NN4BEG[3]
+ Tile_X2Y4_LUT4AB/NN4BEG[4] Tile_X2Y4_LUT4AB/NN4BEG[5] Tile_X2Y4_LUT4AB/NN4BEG[6]
+ Tile_X2Y4_LUT4AB/NN4BEG[7] Tile_X2Y4_LUT4AB/NN4BEG[8] Tile_X2Y4_LUT4AB/NN4BEG[9]
+ Tile_X2Y4_LUT4AB/S1END[0] Tile_X2Y4_LUT4AB/S1END[1] Tile_X2Y4_LUT4AB/S1END[2] Tile_X2Y4_LUT4AB/S1END[3]
+ Tile_X2Y3_LUT4AB/S1END[0] Tile_X2Y3_LUT4AB/S1END[1] Tile_X2Y3_LUT4AB/S1END[2] Tile_X2Y3_LUT4AB/S1END[3]
+ Tile_X2Y4_LUT4AB/S2MID[0] Tile_X2Y4_LUT4AB/S2MID[1] Tile_X2Y4_LUT4AB/S2MID[2] Tile_X2Y4_LUT4AB/S2MID[3]
+ Tile_X2Y4_LUT4AB/S2MID[4] Tile_X2Y4_LUT4AB/S2MID[5] Tile_X2Y4_LUT4AB/S2MID[6] Tile_X2Y4_LUT4AB/S2MID[7]
+ Tile_X2Y4_LUT4AB/S2END[0] Tile_X2Y4_LUT4AB/S2END[1] Tile_X2Y4_LUT4AB/S2END[2] Tile_X2Y4_LUT4AB/S2END[3]
+ Tile_X2Y4_LUT4AB/S2END[4] Tile_X2Y4_LUT4AB/S2END[5] Tile_X2Y4_LUT4AB/S2END[6] Tile_X2Y4_LUT4AB/S2END[7]
+ Tile_X2Y3_LUT4AB/S2END[0] Tile_X2Y3_LUT4AB/S2END[1] Tile_X2Y3_LUT4AB/S2END[2] Tile_X2Y3_LUT4AB/S2END[3]
+ Tile_X2Y3_LUT4AB/S2END[4] Tile_X2Y3_LUT4AB/S2END[5] Tile_X2Y3_LUT4AB/S2END[6] Tile_X2Y3_LUT4AB/S2END[7]
+ Tile_X2Y3_LUT4AB/S2MID[0] Tile_X2Y3_LUT4AB/S2MID[1] Tile_X2Y3_LUT4AB/S2MID[2] Tile_X2Y3_LUT4AB/S2MID[3]
+ Tile_X2Y3_LUT4AB/S2MID[4] Tile_X2Y3_LUT4AB/S2MID[5] Tile_X2Y3_LUT4AB/S2MID[6] Tile_X2Y3_LUT4AB/S2MID[7]
+ Tile_X2Y4_LUT4AB/S4END[0] Tile_X2Y4_LUT4AB/S4END[10] Tile_X2Y4_LUT4AB/S4END[11]
+ Tile_X2Y4_LUT4AB/S4END[12] Tile_X2Y4_LUT4AB/S4END[13] Tile_X2Y4_LUT4AB/S4END[14]
+ Tile_X2Y4_LUT4AB/S4END[15] Tile_X2Y4_LUT4AB/S4END[1] Tile_X2Y4_LUT4AB/S4END[2] Tile_X2Y4_LUT4AB/S4END[3]
+ Tile_X2Y4_LUT4AB/S4END[4] Tile_X2Y4_LUT4AB/S4END[5] Tile_X2Y4_LUT4AB/S4END[6] Tile_X2Y4_LUT4AB/S4END[7]
+ Tile_X2Y4_LUT4AB/S4END[8] Tile_X2Y4_LUT4AB/S4END[9] Tile_X2Y3_LUT4AB/S4END[0] Tile_X2Y3_LUT4AB/S4END[10]
+ Tile_X2Y3_LUT4AB/S4END[11] Tile_X2Y3_LUT4AB/S4END[12] Tile_X2Y3_LUT4AB/S4END[13]
+ Tile_X2Y3_LUT4AB/S4END[14] Tile_X2Y3_LUT4AB/S4END[15] Tile_X2Y3_LUT4AB/S4END[1]
+ Tile_X2Y3_LUT4AB/S4END[2] Tile_X2Y3_LUT4AB/S4END[3] Tile_X2Y3_LUT4AB/S4END[4] Tile_X2Y3_LUT4AB/S4END[5]
+ Tile_X2Y3_LUT4AB/S4END[6] Tile_X2Y3_LUT4AB/S4END[7] Tile_X2Y3_LUT4AB/S4END[8] Tile_X2Y3_LUT4AB/S4END[9]
+ Tile_X2Y4_LUT4AB/SS4END[0] Tile_X2Y4_LUT4AB/SS4END[10] Tile_X2Y4_LUT4AB/SS4END[11]
+ Tile_X2Y4_LUT4AB/SS4END[12] Tile_X2Y4_LUT4AB/SS4END[13] Tile_X2Y4_LUT4AB/SS4END[14]
+ Tile_X2Y4_LUT4AB/SS4END[15] Tile_X2Y4_LUT4AB/SS4END[1] Tile_X2Y4_LUT4AB/SS4END[2]
+ Tile_X2Y4_LUT4AB/SS4END[3] Tile_X2Y4_LUT4AB/SS4END[4] Tile_X2Y4_LUT4AB/SS4END[5]
+ Tile_X2Y4_LUT4AB/SS4END[6] Tile_X2Y4_LUT4AB/SS4END[7] Tile_X2Y4_LUT4AB/SS4END[8]
+ Tile_X2Y4_LUT4AB/SS4END[9] Tile_X2Y3_LUT4AB/SS4END[0] Tile_X2Y3_LUT4AB/SS4END[10]
+ Tile_X2Y3_LUT4AB/SS4END[11] Tile_X2Y3_LUT4AB/SS4END[12] Tile_X2Y3_LUT4AB/SS4END[13]
+ Tile_X2Y3_LUT4AB/SS4END[14] Tile_X2Y3_LUT4AB/SS4END[15] Tile_X2Y3_LUT4AB/SS4END[1]
+ Tile_X2Y3_LUT4AB/SS4END[2] Tile_X2Y3_LUT4AB/SS4END[3] Tile_X2Y3_LUT4AB/SS4END[4]
+ Tile_X2Y3_LUT4AB/SS4END[5] Tile_X2Y3_LUT4AB/SS4END[6] Tile_X2Y3_LUT4AB/SS4END[7]
+ Tile_X2Y3_LUT4AB/SS4END[8] Tile_X2Y3_LUT4AB/SS4END[9] Tile_X2Y3_LUT4AB/UserCLK Tile_X2Y2_LUT4AB/UserCLK
+ VGND VPWR Tile_X2Y3_LUT4AB/W1BEG[0] Tile_X2Y3_LUT4AB/W1BEG[1] Tile_X2Y3_LUT4AB/W1BEG[2]
+ Tile_X2Y3_LUT4AB/W1BEG[3] Tile_X3Y3_LUT4AB/W1BEG[0] Tile_X3Y3_LUT4AB/W1BEG[1] Tile_X3Y3_LUT4AB/W1BEG[2]
+ Tile_X3Y3_LUT4AB/W1BEG[3] Tile_X2Y3_LUT4AB/W2BEG[0] Tile_X2Y3_LUT4AB/W2BEG[1] Tile_X2Y3_LUT4AB/W2BEG[2]
+ Tile_X2Y3_LUT4AB/W2BEG[3] Tile_X2Y3_LUT4AB/W2BEG[4] Tile_X2Y3_LUT4AB/W2BEG[5] Tile_X2Y3_LUT4AB/W2BEG[6]
+ Tile_X2Y3_LUT4AB/W2BEG[7] Tile_X1Y3_LUT4AB/W2END[0] Tile_X1Y3_LUT4AB/W2END[1] Tile_X1Y3_LUT4AB/W2END[2]
+ Tile_X1Y3_LUT4AB/W2END[3] Tile_X1Y3_LUT4AB/W2END[4] Tile_X1Y3_LUT4AB/W2END[5] Tile_X1Y3_LUT4AB/W2END[6]
+ Tile_X1Y3_LUT4AB/W2END[7] Tile_X2Y3_LUT4AB/W2END[0] Tile_X2Y3_LUT4AB/W2END[1] Tile_X2Y3_LUT4AB/W2END[2]
+ Tile_X2Y3_LUT4AB/W2END[3] Tile_X2Y3_LUT4AB/W2END[4] Tile_X2Y3_LUT4AB/W2END[5] Tile_X2Y3_LUT4AB/W2END[6]
+ Tile_X2Y3_LUT4AB/W2END[7] Tile_X3Y3_LUT4AB/W2BEG[0] Tile_X3Y3_LUT4AB/W2BEG[1] Tile_X3Y3_LUT4AB/W2BEG[2]
+ Tile_X3Y3_LUT4AB/W2BEG[3] Tile_X3Y3_LUT4AB/W2BEG[4] Tile_X3Y3_LUT4AB/W2BEG[5] Tile_X3Y3_LUT4AB/W2BEG[6]
+ Tile_X3Y3_LUT4AB/W2BEG[7] Tile_X2Y3_LUT4AB/W6BEG[0] Tile_X2Y3_LUT4AB/W6BEG[10] Tile_X2Y3_LUT4AB/W6BEG[11]
+ Tile_X2Y3_LUT4AB/W6BEG[1] Tile_X2Y3_LUT4AB/W6BEG[2] Tile_X2Y3_LUT4AB/W6BEG[3] Tile_X2Y3_LUT4AB/W6BEG[4]
+ Tile_X2Y3_LUT4AB/W6BEG[5] Tile_X2Y3_LUT4AB/W6BEG[6] Tile_X2Y3_LUT4AB/W6BEG[7] Tile_X2Y3_LUT4AB/W6BEG[8]
+ Tile_X2Y3_LUT4AB/W6BEG[9] Tile_X3Y3_LUT4AB/W6BEG[0] Tile_X3Y3_LUT4AB/W6BEG[10] Tile_X3Y3_LUT4AB/W6BEG[11]
+ Tile_X3Y3_LUT4AB/W6BEG[1] Tile_X3Y3_LUT4AB/W6BEG[2] Tile_X3Y3_LUT4AB/W6BEG[3] Tile_X3Y3_LUT4AB/W6BEG[4]
+ Tile_X3Y3_LUT4AB/W6BEG[5] Tile_X3Y3_LUT4AB/W6BEG[6] Tile_X3Y3_LUT4AB/W6BEG[7] Tile_X3Y3_LUT4AB/W6BEG[8]
+ Tile_X3Y3_LUT4AB/W6BEG[9] Tile_X2Y3_LUT4AB/WW4BEG[0] Tile_X2Y3_LUT4AB/WW4BEG[10]
+ Tile_X2Y3_LUT4AB/WW4BEG[11] Tile_X2Y3_LUT4AB/WW4BEG[12] Tile_X2Y3_LUT4AB/WW4BEG[13]
+ Tile_X2Y3_LUT4AB/WW4BEG[14] Tile_X2Y3_LUT4AB/WW4BEG[15] Tile_X2Y3_LUT4AB/WW4BEG[1]
+ Tile_X2Y3_LUT4AB/WW4BEG[2] Tile_X2Y3_LUT4AB/WW4BEG[3] Tile_X2Y3_LUT4AB/WW4BEG[4]
+ Tile_X2Y3_LUT4AB/WW4BEG[5] Tile_X2Y3_LUT4AB/WW4BEG[6] Tile_X2Y3_LUT4AB/WW4BEG[7]
+ Tile_X2Y3_LUT4AB/WW4BEG[8] Tile_X2Y3_LUT4AB/WW4BEG[9] Tile_X3Y3_LUT4AB/WW4BEG[0]
+ Tile_X3Y3_LUT4AB/WW4BEG[10] Tile_X3Y3_LUT4AB/WW4BEG[11] Tile_X3Y3_LUT4AB/WW4BEG[12]
+ Tile_X3Y3_LUT4AB/WW4BEG[13] Tile_X3Y3_LUT4AB/WW4BEG[14] Tile_X3Y3_LUT4AB/WW4BEG[15]
+ Tile_X3Y3_LUT4AB/WW4BEG[1] Tile_X3Y3_LUT4AB/WW4BEG[2] Tile_X3Y3_LUT4AB/WW4BEG[3]
+ Tile_X3Y3_LUT4AB/WW4BEG[4] Tile_X3Y3_LUT4AB/WW4BEG[5] Tile_X3Y3_LUT4AB/WW4BEG[6]
+ Tile_X3Y3_LUT4AB/WW4BEG[7] Tile_X3Y3_LUT4AB/WW4BEG[8] Tile_X3Y3_LUT4AB/WW4BEG[9]
+ LUT4AB
XTile_X0Y5_W_TT_IF Tile_X0Y5_CLK_TT_PROJECT Tile_X1Y5_LUT4AB/E1END[0] Tile_X1Y5_LUT4AB/E1END[1]
+ Tile_X1Y5_LUT4AB/E1END[2] Tile_X1Y5_LUT4AB/E1END[3] Tile_X1Y5_LUT4AB/E2MID[0] Tile_X1Y5_LUT4AB/E2MID[1]
+ Tile_X1Y5_LUT4AB/E2MID[2] Tile_X1Y5_LUT4AB/E2MID[3] Tile_X1Y5_LUT4AB/E2MID[4] Tile_X1Y5_LUT4AB/E2MID[5]
+ Tile_X1Y5_LUT4AB/E2MID[6] Tile_X1Y5_LUT4AB/E2MID[7] Tile_X1Y5_LUT4AB/E2END[0] Tile_X1Y5_LUT4AB/E2END[1]
+ Tile_X1Y5_LUT4AB/E2END[2] Tile_X1Y5_LUT4AB/E2END[3] Tile_X1Y5_LUT4AB/E2END[4] Tile_X1Y5_LUT4AB/E2END[5]
+ Tile_X1Y5_LUT4AB/E2END[6] Tile_X1Y5_LUT4AB/E2END[7] Tile_X1Y5_LUT4AB/E6END[0] Tile_X1Y5_LUT4AB/E6END[10]
+ Tile_X1Y5_LUT4AB/E6END[11] Tile_X1Y5_LUT4AB/E6END[1] Tile_X1Y5_LUT4AB/E6END[2] Tile_X1Y5_LUT4AB/E6END[3]
+ Tile_X1Y5_LUT4AB/E6END[4] Tile_X1Y5_LUT4AB/E6END[5] Tile_X1Y5_LUT4AB/E6END[6] Tile_X1Y5_LUT4AB/E6END[7]
+ Tile_X1Y5_LUT4AB/E6END[8] Tile_X1Y5_LUT4AB/E6END[9] Tile_X1Y5_LUT4AB/EE4END[0] Tile_X1Y5_LUT4AB/EE4END[10]
+ Tile_X1Y5_LUT4AB/EE4END[11] Tile_X1Y5_LUT4AB/EE4END[12] Tile_X1Y5_LUT4AB/EE4END[13]
+ Tile_X1Y5_LUT4AB/EE4END[14] Tile_X1Y5_LUT4AB/EE4END[15] Tile_X1Y5_LUT4AB/EE4END[1]
+ Tile_X1Y5_LUT4AB/EE4END[2] Tile_X1Y5_LUT4AB/EE4END[3] Tile_X1Y5_LUT4AB/EE4END[4]
+ Tile_X1Y5_LUT4AB/EE4END[5] Tile_X1Y5_LUT4AB/EE4END[6] Tile_X1Y5_LUT4AB/EE4END[7]
+ Tile_X1Y5_LUT4AB/EE4END[8] Tile_X1Y5_LUT4AB/EE4END[9] Tile_X0Y5_ENA_TT_PROJECT FrameData[160]
+ FrameData[170] FrameData[171] FrameData[172] FrameData[173] FrameData[174] FrameData[175]
+ FrameData[176] FrameData[177] FrameData[178] FrameData[179] FrameData[161] FrameData[180]
+ FrameData[181] FrameData[182] FrameData[183] FrameData[184] FrameData[185] FrameData[186]
+ FrameData[187] FrameData[188] FrameData[189] FrameData[162] FrameData[190] FrameData[191]
+ FrameData[163] FrameData[164] FrameData[165] FrameData[166] FrameData[167] FrameData[168]
+ FrameData[169] Tile_X1Y5_LUT4AB/FrameData[0] Tile_X1Y5_LUT4AB/FrameData[10] Tile_X1Y5_LUT4AB/FrameData[11]
+ Tile_X1Y5_LUT4AB/FrameData[12] Tile_X1Y5_LUT4AB/FrameData[13] Tile_X1Y5_LUT4AB/FrameData[14]
+ Tile_X1Y5_LUT4AB/FrameData[15] Tile_X1Y5_LUT4AB/FrameData[16] Tile_X1Y5_LUT4AB/FrameData[17]
+ Tile_X1Y5_LUT4AB/FrameData[18] Tile_X1Y5_LUT4AB/FrameData[19] Tile_X1Y5_LUT4AB/FrameData[1]
+ Tile_X1Y5_LUT4AB/FrameData[20] Tile_X1Y5_LUT4AB/FrameData[21] Tile_X1Y5_LUT4AB/FrameData[22]
+ Tile_X1Y5_LUT4AB/FrameData[23] Tile_X1Y5_LUT4AB/FrameData[24] Tile_X1Y5_LUT4AB/FrameData[25]
+ Tile_X1Y5_LUT4AB/FrameData[26] Tile_X1Y5_LUT4AB/FrameData[27] Tile_X1Y5_LUT4AB/FrameData[28]
+ Tile_X1Y5_LUT4AB/FrameData[29] Tile_X1Y5_LUT4AB/FrameData[2] Tile_X1Y5_LUT4AB/FrameData[30]
+ Tile_X1Y5_LUT4AB/FrameData[31] Tile_X1Y5_LUT4AB/FrameData[3] Tile_X1Y5_LUT4AB/FrameData[4]
+ Tile_X1Y5_LUT4AB/FrameData[5] Tile_X1Y5_LUT4AB/FrameData[6] Tile_X1Y5_LUT4AB/FrameData[7]
+ Tile_X1Y5_LUT4AB/FrameData[8] Tile_X1Y5_LUT4AB/FrameData[9] Tile_X0Y5_W_TT_IF/FrameStrobe[0]
+ Tile_X0Y5_W_TT_IF/FrameStrobe[10] Tile_X0Y5_W_TT_IF/FrameStrobe[11] Tile_X0Y5_W_TT_IF/FrameStrobe[12]
+ Tile_X0Y5_W_TT_IF/FrameStrobe[13] Tile_X0Y5_W_TT_IF/FrameStrobe[14] Tile_X0Y5_W_TT_IF/FrameStrobe[15]
+ Tile_X0Y5_W_TT_IF/FrameStrobe[16] Tile_X0Y5_W_TT_IF/FrameStrobe[17] Tile_X0Y5_W_TT_IF/FrameStrobe[18]
+ Tile_X0Y5_W_TT_IF/FrameStrobe[19] Tile_X0Y5_W_TT_IF/FrameStrobe[1] Tile_X0Y5_W_TT_IF/FrameStrobe[2]
+ Tile_X0Y5_W_TT_IF/FrameStrobe[3] Tile_X0Y5_W_TT_IF/FrameStrobe[4] Tile_X0Y5_W_TT_IF/FrameStrobe[5]
+ Tile_X0Y5_W_TT_IF/FrameStrobe[6] Tile_X0Y5_W_TT_IF/FrameStrobe[7] Tile_X0Y5_W_TT_IF/FrameStrobe[8]
+ Tile_X0Y5_W_TT_IF/FrameStrobe[9] Tile_X0Y4_W_TT_IF/FrameStrobe[0] Tile_X0Y4_W_TT_IF/FrameStrobe[10]
+ Tile_X0Y4_W_TT_IF/FrameStrobe[11] Tile_X0Y4_W_TT_IF/FrameStrobe[12] Tile_X0Y4_W_TT_IF/FrameStrobe[13]
+ Tile_X0Y4_W_TT_IF/FrameStrobe[14] Tile_X0Y4_W_TT_IF/FrameStrobe[15] Tile_X0Y4_W_TT_IF/FrameStrobe[16]
+ Tile_X0Y4_W_TT_IF/FrameStrobe[17] Tile_X0Y4_W_TT_IF/FrameStrobe[18] Tile_X0Y4_W_TT_IF/FrameStrobe[19]
+ Tile_X0Y4_W_TT_IF/FrameStrobe[1] Tile_X0Y4_W_TT_IF/FrameStrobe[2] Tile_X0Y4_W_TT_IF/FrameStrobe[3]
+ Tile_X0Y4_W_TT_IF/FrameStrobe[4] Tile_X0Y4_W_TT_IF/FrameStrobe[5] Tile_X0Y4_W_TT_IF/FrameStrobe[6]
+ Tile_X0Y4_W_TT_IF/FrameStrobe[7] Tile_X0Y4_W_TT_IF/FrameStrobe[8] Tile_X0Y4_W_TT_IF/FrameStrobe[9]
+ Tile_X0Y5_W_TT_IF/N1BEG[0] Tile_X0Y5_W_TT_IF/N1BEG[1] Tile_X0Y5_W_TT_IF/N1BEG[2]
+ Tile_X0Y5_W_TT_IF/N1BEG[3] Tile_X0Y6_W_TT_IF/N1BEG[0] Tile_X0Y6_W_TT_IF/N1BEG[1]
+ Tile_X0Y6_W_TT_IF/N1BEG[2] Tile_X0Y6_W_TT_IF/N1BEG[3] Tile_X0Y5_W_TT_IF/N2BEG[0]
+ Tile_X0Y5_W_TT_IF/N2BEG[1] Tile_X0Y5_W_TT_IF/N2BEG[2] Tile_X0Y5_W_TT_IF/N2BEG[3]
+ Tile_X0Y5_W_TT_IF/N2BEG[4] Tile_X0Y5_W_TT_IF/N2BEG[5] Tile_X0Y5_W_TT_IF/N2BEG[6]
+ Tile_X0Y5_W_TT_IF/N2BEG[7] Tile_X0Y4_W_TT_IF/N2END[0] Tile_X0Y4_W_TT_IF/N2END[1]
+ Tile_X0Y4_W_TT_IF/N2END[2] Tile_X0Y4_W_TT_IF/N2END[3] Tile_X0Y4_W_TT_IF/N2END[4]
+ Tile_X0Y4_W_TT_IF/N2END[5] Tile_X0Y4_W_TT_IF/N2END[6] Tile_X0Y4_W_TT_IF/N2END[7]
+ Tile_X0Y5_W_TT_IF/N2END[0] Tile_X0Y5_W_TT_IF/N2END[1] Tile_X0Y5_W_TT_IF/N2END[2]
+ Tile_X0Y5_W_TT_IF/N2END[3] Tile_X0Y5_W_TT_IF/N2END[4] Tile_X0Y5_W_TT_IF/N2END[5]
+ Tile_X0Y5_W_TT_IF/N2END[6] Tile_X0Y5_W_TT_IF/N2END[7] Tile_X0Y6_W_TT_IF/N2BEG[0]
+ Tile_X0Y6_W_TT_IF/N2BEG[1] Tile_X0Y6_W_TT_IF/N2BEG[2] Tile_X0Y6_W_TT_IF/N2BEG[3]
+ Tile_X0Y6_W_TT_IF/N2BEG[4] Tile_X0Y6_W_TT_IF/N2BEG[5] Tile_X0Y6_W_TT_IF/N2BEG[6]
+ Tile_X0Y6_W_TT_IF/N2BEG[7] Tile_X0Y5_W_TT_IF/N4BEG[0] Tile_X0Y5_W_TT_IF/N4BEG[10]
+ Tile_X0Y5_W_TT_IF/N4BEG[11] Tile_X0Y5_W_TT_IF/N4BEG[12] Tile_X0Y5_W_TT_IF/N4BEG[13]
+ Tile_X0Y5_W_TT_IF/N4BEG[14] Tile_X0Y5_W_TT_IF/N4BEG[15] Tile_X0Y5_W_TT_IF/N4BEG[1]
+ Tile_X0Y5_W_TT_IF/N4BEG[2] Tile_X0Y5_W_TT_IF/N4BEG[3] Tile_X0Y5_W_TT_IF/N4BEG[4]
+ Tile_X0Y5_W_TT_IF/N4BEG[5] Tile_X0Y5_W_TT_IF/N4BEG[6] Tile_X0Y5_W_TT_IF/N4BEG[7]
+ Tile_X0Y5_W_TT_IF/N4BEG[8] Tile_X0Y5_W_TT_IF/N4BEG[9] Tile_X0Y6_W_TT_IF/N4BEG[0]
+ Tile_X0Y6_W_TT_IF/N4BEG[10] Tile_X0Y6_W_TT_IF/N4BEG[11] Tile_X0Y6_W_TT_IF/N4BEG[12]
+ Tile_X0Y6_W_TT_IF/N4BEG[13] Tile_X0Y6_W_TT_IF/N4BEG[14] Tile_X0Y6_W_TT_IF/N4BEG[15]
+ Tile_X0Y6_W_TT_IF/N4BEG[1] Tile_X0Y6_W_TT_IF/N4BEG[2] Tile_X0Y6_W_TT_IF/N4BEG[3]
+ Tile_X0Y6_W_TT_IF/N4BEG[4] Tile_X0Y6_W_TT_IF/N4BEG[5] Tile_X0Y6_W_TT_IF/N4BEG[6]
+ Tile_X0Y6_W_TT_IF/N4BEG[7] Tile_X0Y6_W_TT_IF/N4BEG[8] Tile_X0Y6_W_TT_IF/N4BEG[9]
+ Tile_X0Y5_RST_N_TT_PROJECT Tile_X0Y6_W_TT_IF/S1END[0] Tile_X0Y6_W_TT_IF/S1END[1]
+ Tile_X0Y6_W_TT_IF/S1END[2] Tile_X0Y6_W_TT_IF/S1END[3] Tile_X0Y5_W_TT_IF/S1END[0]
+ Tile_X0Y5_W_TT_IF/S1END[1] Tile_X0Y5_W_TT_IF/S1END[2] Tile_X0Y5_W_TT_IF/S1END[3]
+ Tile_X0Y6_W_TT_IF/S2MID[0] Tile_X0Y6_W_TT_IF/S2MID[1] Tile_X0Y6_W_TT_IF/S2MID[2]
+ Tile_X0Y6_W_TT_IF/S2MID[3] Tile_X0Y6_W_TT_IF/S2MID[4] Tile_X0Y6_W_TT_IF/S2MID[5]
+ Tile_X0Y6_W_TT_IF/S2MID[6] Tile_X0Y6_W_TT_IF/S2MID[7] Tile_X0Y6_W_TT_IF/S2END[0]
+ Tile_X0Y6_W_TT_IF/S2END[1] Tile_X0Y6_W_TT_IF/S2END[2] Tile_X0Y6_W_TT_IF/S2END[3]
+ Tile_X0Y6_W_TT_IF/S2END[4] Tile_X0Y6_W_TT_IF/S2END[5] Tile_X0Y6_W_TT_IF/S2END[6]
+ Tile_X0Y6_W_TT_IF/S2END[7] Tile_X0Y5_W_TT_IF/S2END[0] Tile_X0Y5_W_TT_IF/S2END[1]
+ Tile_X0Y5_W_TT_IF/S2END[2] Tile_X0Y5_W_TT_IF/S2END[3] Tile_X0Y5_W_TT_IF/S2END[4]
+ Tile_X0Y5_W_TT_IF/S2END[5] Tile_X0Y5_W_TT_IF/S2END[6] Tile_X0Y5_W_TT_IF/S2END[7]
+ Tile_X0Y5_W_TT_IF/S2MID[0] Tile_X0Y5_W_TT_IF/S2MID[1] Tile_X0Y5_W_TT_IF/S2MID[2]
+ Tile_X0Y5_W_TT_IF/S2MID[3] Tile_X0Y5_W_TT_IF/S2MID[4] Tile_X0Y5_W_TT_IF/S2MID[5]
+ Tile_X0Y5_W_TT_IF/S2MID[6] Tile_X0Y5_W_TT_IF/S2MID[7] Tile_X0Y6_W_TT_IF/S4END[0]
+ Tile_X0Y6_W_TT_IF/S4END[10] Tile_X0Y6_W_TT_IF/S4END[11] Tile_X0Y6_W_TT_IF/S4END[12]
+ Tile_X0Y6_W_TT_IF/S4END[13] Tile_X0Y6_W_TT_IF/S4END[14] Tile_X0Y6_W_TT_IF/S4END[15]
+ Tile_X0Y6_W_TT_IF/S4END[1] Tile_X0Y6_W_TT_IF/S4END[2] Tile_X0Y6_W_TT_IF/S4END[3]
+ Tile_X0Y6_W_TT_IF/S4END[4] Tile_X0Y6_W_TT_IF/S4END[5] Tile_X0Y6_W_TT_IF/S4END[6]
+ Tile_X0Y6_W_TT_IF/S4END[7] Tile_X0Y6_W_TT_IF/S4END[8] Tile_X0Y6_W_TT_IF/S4END[9]
+ Tile_X0Y5_W_TT_IF/S4END[0] Tile_X0Y5_W_TT_IF/S4END[10] Tile_X0Y5_W_TT_IF/S4END[11]
+ Tile_X0Y5_W_TT_IF/S4END[12] Tile_X0Y5_W_TT_IF/S4END[13] Tile_X0Y5_W_TT_IF/S4END[14]
+ Tile_X0Y5_W_TT_IF/S4END[15] Tile_X0Y5_W_TT_IF/S4END[1] Tile_X0Y5_W_TT_IF/S4END[2]
+ Tile_X0Y5_W_TT_IF/S4END[3] Tile_X0Y5_W_TT_IF/S4END[4] Tile_X0Y5_W_TT_IF/S4END[5]
+ Tile_X0Y5_W_TT_IF/S4END[6] Tile_X0Y5_W_TT_IF/S4END[7] Tile_X0Y5_W_TT_IF/S4END[8]
+ Tile_X0Y5_W_TT_IF/S4END[9] Tile_X0Y5_UIO_IN_TT_PROJECT0 Tile_X0Y5_UIO_IN_TT_PROJECT1
+ Tile_X0Y5_UIO_IN_TT_PROJECT2 Tile_X0Y5_UIO_IN_TT_PROJECT3 Tile_X0Y5_UIO_IN_TT_PROJECT4
+ Tile_X0Y5_UIO_IN_TT_PROJECT5 Tile_X0Y5_UIO_IN_TT_PROJECT6 Tile_X0Y5_UIO_IN_TT_PROJECT7
+ Tile_X0Y5_UIO_OE_TT_PROJECT0 Tile_X0Y5_UIO_OE_TT_PROJECT1 Tile_X0Y5_UIO_OE_TT_PROJECT2
+ Tile_X0Y5_UIO_OE_TT_PROJECT3 Tile_X0Y5_UIO_OE_TT_PROJECT4 Tile_X0Y5_UIO_OE_TT_PROJECT5
+ Tile_X0Y5_UIO_OE_TT_PROJECT6 Tile_X0Y5_UIO_OE_TT_PROJECT7 Tile_X0Y5_UIO_OUT_TT_PROJECT0
+ Tile_X0Y5_UIO_OUT_TT_PROJECT1 Tile_X0Y5_UIO_OUT_TT_PROJECT2 Tile_X0Y5_UIO_OUT_TT_PROJECT3
+ Tile_X0Y5_UIO_OUT_TT_PROJECT4 Tile_X0Y5_UIO_OUT_TT_PROJECT5 Tile_X0Y5_UIO_OUT_TT_PROJECT6
+ Tile_X0Y5_UIO_OUT_TT_PROJECT7 Tile_X0Y5_UI_IN_TT_PROJECT0 Tile_X0Y5_UI_IN_TT_PROJECT1
+ Tile_X0Y5_UI_IN_TT_PROJECT2 Tile_X0Y5_UI_IN_TT_PROJECT3 Tile_X0Y5_UI_IN_TT_PROJECT4
+ Tile_X0Y5_UI_IN_TT_PROJECT5 Tile_X0Y5_UI_IN_TT_PROJECT6 Tile_X0Y5_UI_IN_TT_PROJECT7
+ Tile_X0Y5_UO_OUT_TT_PROJECT0 Tile_X0Y5_UO_OUT_TT_PROJECT1 Tile_X0Y5_UO_OUT_TT_PROJECT2
+ Tile_X0Y5_UO_OUT_TT_PROJECT3 Tile_X0Y5_UO_OUT_TT_PROJECT4 Tile_X0Y5_UO_OUT_TT_PROJECT5
+ Tile_X0Y5_UO_OUT_TT_PROJECT6 Tile_X0Y5_UO_OUT_TT_PROJECT7 Tile_X0Y5_W_TT_IF/UserCLK
+ Tile_X0Y4_W_TT_IF/UserCLK VGND VPWR Tile_X1Y5_LUT4AB/W1BEG[0] Tile_X1Y5_LUT4AB/W1BEG[1]
+ Tile_X1Y5_LUT4AB/W1BEG[2] Tile_X1Y5_LUT4AB/W1BEG[3] Tile_X1Y5_LUT4AB/W2BEGb[0] Tile_X1Y5_LUT4AB/W2BEGb[1]
+ Tile_X1Y5_LUT4AB/W2BEGb[2] Tile_X1Y5_LUT4AB/W2BEGb[3] Tile_X1Y5_LUT4AB/W2BEGb[4]
+ Tile_X1Y5_LUT4AB/W2BEGb[5] Tile_X1Y5_LUT4AB/W2BEGb[6] Tile_X1Y5_LUT4AB/W2BEGb[7]
+ Tile_X1Y5_LUT4AB/W2BEG[0] Tile_X1Y5_LUT4AB/W2BEG[1] Tile_X1Y5_LUT4AB/W2BEG[2] Tile_X1Y5_LUT4AB/W2BEG[3]
+ Tile_X1Y5_LUT4AB/W2BEG[4] Tile_X1Y5_LUT4AB/W2BEG[5] Tile_X1Y5_LUT4AB/W2BEG[6] Tile_X1Y5_LUT4AB/W2BEG[7]
+ Tile_X1Y5_LUT4AB/W6BEG[0] Tile_X1Y5_LUT4AB/W6BEG[10] Tile_X1Y5_LUT4AB/W6BEG[11]
+ Tile_X1Y5_LUT4AB/W6BEG[1] Tile_X1Y5_LUT4AB/W6BEG[2] Tile_X1Y5_LUT4AB/W6BEG[3] Tile_X1Y5_LUT4AB/W6BEG[4]
+ Tile_X1Y5_LUT4AB/W6BEG[5] Tile_X1Y5_LUT4AB/W6BEG[6] Tile_X1Y5_LUT4AB/W6BEG[7] Tile_X1Y5_LUT4AB/W6BEG[8]
+ Tile_X1Y5_LUT4AB/W6BEG[9] Tile_X1Y5_LUT4AB/WW4BEG[0] Tile_X1Y5_LUT4AB/WW4BEG[10]
+ Tile_X1Y5_LUT4AB/WW4BEG[11] Tile_X1Y5_LUT4AB/WW4BEG[12] Tile_X1Y5_LUT4AB/WW4BEG[13]
+ Tile_X1Y5_LUT4AB/WW4BEG[14] Tile_X1Y5_LUT4AB/WW4BEG[15] Tile_X1Y5_LUT4AB/WW4BEG[1]
+ Tile_X1Y5_LUT4AB/WW4BEG[2] Tile_X1Y5_LUT4AB/WW4BEG[3] Tile_X1Y5_LUT4AB/WW4BEG[4]
+ Tile_X1Y5_LUT4AB/WW4BEG[5] Tile_X1Y5_LUT4AB/WW4BEG[6] Tile_X1Y5_LUT4AB/WW4BEG[7]
+ Tile_X1Y5_LUT4AB/WW4BEG[8] Tile_X1Y5_LUT4AB/WW4BEG[9] W_TT_IF
XTile_X1Y7_LUT4AB Tile_X1Y8_LUT4AB/Co Tile_X1Y7_LUT4AB/Co Tile_X2Y7_LUT4AB/E1END[0]
+ Tile_X2Y7_LUT4AB/E1END[1] Tile_X2Y7_LUT4AB/E1END[2] Tile_X2Y7_LUT4AB/E1END[3] Tile_X1Y7_LUT4AB/E1END[0]
+ Tile_X1Y7_LUT4AB/E1END[1] Tile_X1Y7_LUT4AB/E1END[2] Tile_X1Y7_LUT4AB/E1END[3] Tile_X2Y7_LUT4AB/E2MID[0]
+ Tile_X2Y7_LUT4AB/E2MID[1] Tile_X2Y7_LUT4AB/E2MID[2] Tile_X2Y7_LUT4AB/E2MID[3] Tile_X2Y7_LUT4AB/E2MID[4]
+ Tile_X2Y7_LUT4AB/E2MID[5] Tile_X2Y7_LUT4AB/E2MID[6] Tile_X2Y7_LUT4AB/E2MID[7] Tile_X2Y7_LUT4AB/E2END[0]
+ Tile_X2Y7_LUT4AB/E2END[1] Tile_X2Y7_LUT4AB/E2END[2] Tile_X2Y7_LUT4AB/E2END[3] Tile_X2Y7_LUT4AB/E2END[4]
+ Tile_X2Y7_LUT4AB/E2END[5] Tile_X2Y7_LUT4AB/E2END[6] Tile_X2Y7_LUT4AB/E2END[7] Tile_X1Y7_LUT4AB/E2END[0]
+ Tile_X1Y7_LUT4AB/E2END[1] Tile_X1Y7_LUT4AB/E2END[2] Tile_X1Y7_LUT4AB/E2END[3] Tile_X1Y7_LUT4AB/E2END[4]
+ Tile_X1Y7_LUT4AB/E2END[5] Tile_X1Y7_LUT4AB/E2END[6] Tile_X1Y7_LUT4AB/E2END[7] Tile_X1Y7_LUT4AB/E2MID[0]
+ Tile_X1Y7_LUT4AB/E2MID[1] Tile_X1Y7_LUT4AB/E2MID[2] Tile_X1Y7_LUT4AB/E2MID[3] Tile_X1Y7_LUT4AB/E2MID[4]
+ Tile_X1Y7_LUT4AB/E2MID[5] Tile_X1Y7_LUT4AB/E2MID[6] Tile_X1Y7_LUT4AB/E2MID[7] Tile_X2Y7_LUT4AB/E6END[0]
+ Tile_X2Y7_LUT4AB/E6END[10] Tile_X2Y7_LUT4AB/E6END[11] Tile_X2Y7_LUT4AB/E6END[1]
+ Tile_X2Y7_LUT4AB/E6END[2] Tile_X2Y7_LUT4AB/E6END[3] Tile_X2Y7_LUT4AB/E6END[4] Tile_X2Y7_LUT4AB/E6END[5]
+ Tile_X2Y7_LUT4AB/E6END[6] Tile_X2Y7_LUT4AB/E6END[7] Tile_X2Y7_LUT4AB/E6END[8] Tile_X2Y7_LUT4AB/E6END[9]
+ Tile_X1Y7_LUT4AB/E6END[0] Tile_X1Y7_LUT4AB/E6END[10] Tile_X1Y7_LUT4AB/E6END[11]
+ Tile_X1Y7_LUT4AB/E6END[1] Tile_X1Y7_LUT4AB/E6END[2] Tile_X1Y7_LUT4AB/E6END[3] Tile_X1Y7_LUT4AB/E6END[4]
+ Tile_X1Y7_LUT4AB/E6END[5] Tile_X1Y7_LUT4AB/E6END[6] Tile_X1Y7_LUT4AB/E6END[7] Tile_X1Y7_LUT4AB/E6END[8]
+ Tile_X1Y7_LUT4AB/E6END[9] Tile_X2Y7_LUT4AB/EE4END[0] Tile_X2Y7_LUT4AB/EE4END[10]
+ Tile_X2Y7_LUT4AB/EE4END[11] Tile_X2Y7_LUT4AB/EE4END[12] Tile_X2Y7_LUT4AB/EE4END[13]
+ Tile_X2Y7_LUT4AB/EE4END[14] Tile_X2Y7_LUT4AB/EE4END[15] Tile_X2Y7_LUT4AB/EE4END[1]
+ Tile_X2Y7_LUT4AB/EE4END[2] Tile_X2Y7_LUT4AB/EE4END[3] Tile_X2Y7_LUT4AB/EE4END[4]
+ Tile_X2Y7_LUT4AB/EE4END[5] Tile_X2Y7_LUT4AB/EE4END[6] Tile_X2Y7_LUT4AB/EE4END[7]
+ Tile_X2Y7_LUT4AB/EE4END[8] Tile_X2Y7_LUT4AB/EE4END[9] Tile_X1Y7_LUT4AB/EE4END[0]
+ Tile_X1Y7_LUT4AB/EE4END[10] Tile_X1Y7_LUT4AB/EE4END[11] Tile_X1Y7_LUT4AB/EE4END[12]
+ Tile_X1Y7_LUT4AB/EE4END[13] Tile_X1Y7_LUT4AB/EE4END[14] Tile_X1Y7_LUT4AB/EE4END[15]
+ Tile_X1Y7_LUT4AB/EE4END[1] Tile_X1Y7_LUT4AB/EE4END[2] Tile_X1Y7_LUT4AB/EE4END[3]
+ Tile_X1Y7_LUT4AB/EE4END[4] Tile_X1Y7_LUT4AB/EE4END[5] Tile_X1Y7_LUT4AB/EE4END[6]
+ Tile_X1Y7_LUT4AB/EE4END[7] Tile_X1Y7_LUT4AB/EE4END[8] Tile_X1Y7_LUT4AB/EE4END[9]
+ Tile_X1Y7_LUT4AB/FrameData[0] Tile_X1Y7_LUT4AB/FrameData[10] Tile_X1Y7_LUT4AB/FrameData[11]
+ Tile_X1Y7_LUT4AB/FrameData[12] Tile_X1Y7_LUT4AB/FrameData[13] Tile_X1Y7_LUT4AB/FrameData[14]
+ Tile_X1Y7_LUT4AB/FrameData[15] Tile_X1Y7_LUT4AB/FrameData[16] Tile_X1Y7_LUT4AB/FrameData[17]
+ Tile_X1Y7_LUT4AB/FrameData[18] Tile_X1Y7_LUT4AB/FrameData[19] Tile_X1Y7_LUT4AB/FrameData[1]
+ Tile_X1Y7_LUT4AB/FrameData[20] Tile_X1Y7_LUT4AB/FrameData[21] Tile_X1Y7_LUT4AB/FrameData[22]
+ Tile_X1Y7_LUT4AB/FrameData[23] Tile_X1Y7_LUT4AB/FrameData[24] Tile_X1Y7_LUT4AB/FrameData[25]
+ Tile_X1Y7_LUT4AB/FrameData[26] Tile_X1Y7_LUT4AB/FrameData[27] Tile_X1Y7_LUT4AB/FrameData[28]
+ Tile_X1Y7_LUT4AB/FrameData[29] Tile_X1Y7_LUT4AB/FrameData[2] Tile_X1Y7_LUT4AB/FrameData[30]
+ Tile_X1Y7_LUT4AB/FrameData[31] Tile_X1Y7_LUT4AB/FrameData[3] Tile_X1Y7_LUT4AB/FrameData[4]
+ Tile_X1Y7_LUT4AB/FrameData[5] Tile_X1Y7_LUT4AB/FrameData[6] Tile_X1Y7_LUT4AB/FrameData[7]
+ Tile_X1Y7_LUT4AB/FrameData[8] Tile_X1Y7_LUT4AB/FrameData[9] Tile_X2Y7_LUT4AB/FrameData[0]
+ Tile_X2Y7_LUT4AB/FrameData[10] Tile_X2Y7_LUT4AB/FrameData[11] Tile_X2Y7_LUT4AB/FrameData[12]
+ Tile_X2Y7_LUT4AB/FrameData[13] Tile_X2Y7_LUT4AB/FrameData[14] Tile_X2Y7_LUT4AB/FrameData[15]
+ Tile_X2Y7_LUT4AB/FrameData[16] Tile_X2Y7_LUT4AB/FrameData[17] Tile_X2Y7_LUT4AB/FrameData[18]
+ Tile_X2Y7_LUT4AB/FrameData[19] Tile_X2Y7_LUT4AB/FrameData[1] Tile_X2Y7_LUT4AB/FrameData[20]
+ Tile_X2Y7_LUT4AB/FrameData[21] Tile_X2Y7_LUT4AB/FrameData[22] Tile_X2Y7_LUT4AB/FrameData[23]
+ Tile_X2Y7_LUT4AB/FrameData[24] Tile_X2Y7_LUT4AB/FrameData[25] Tile_X2Y7_LUT4AB/FrameData[26]
+ Tile_X2Y7_LUT4AB/FrameData[27] Tile_X2Y7_LUT4AB/FrameData[28] Tile_X2Y7_LUT4AB/FrameData[29]
+ Tile_X2Y7_LUT4AB/FrameData[2] Tile_X2Y7_LUT4AB/FrameData[30] Tile_X2Y7_LUT4AB/FrameData[31]
+ Tile_X2Y7_LUT4AB/FrameData[3] Tile_X2Y7_LUT4AB/FrameData[4] Tile_X2Y7_LUT4AB/FrameData[5]
+ Tile_X2Y7_LUT4AB/FrameData[6] Tile_X2Y7_LUT4AB/FrameData[7] Tile_X2Y7_LUT4AB/FrameData[8]
+ Tile_X2Y7_LUT4AB/FrameData[9] Tile_X1Y7_LUT4AB/FrameStrobe[0] Tile_X1Y7_LUT4AB/FrameStrobe[10]
+ Tile_X1Y7_LUT4AB/FrameStrobe[11] Tile_X1Y7_LUT4AB/FrameStrobe[12] Tile_X1Y7_LUT4AB/FrameStrobe[13]
+ Tile_X1Y7_LUT4AB/FrameStrobe[14] Tile_X1Y7_LUT4AB/FrameStrobe[15] Tile_X1Y7_LUT4AB/FrameStrobe[16]
+ Tile_X1Y7_LUT4AB/FrameStrobe[17] Tile_X1Y7_LUT4AB/FrameStrobe[18] Tile_X1Y7_LUT4AB/FrameStrobe[19]
+ Tile_X1Y7_LUT4AB/FrameStrobe[1] Tile_X1Y7_LUT4AB/FrameStrobe[2] Tile_X1Y7_LUT4AB/FrameStrobe[3]
+ Tile_X1Y7_LUT4AB/FrameStrobe[4] Tile_X1Y7_LUT4AB/FrameStrobe[5] Tile_X1Y7_LUT4AB/FrameStrobe[6]
+ Tile_X1Y7_LUT4AB/FrameStrobe[7] Tile_X1Y7_LUT4AB/FrameStrobe[8] Tile_X1Y7_LUT4AB/FrameStrobe[9]
+ Tile_X1Y6_LUT4AB/FrameStrobe[0] Tile_X1Y6_LUT4AB/FrameStrobe[10] Tile_X1Y6_LUT4AB/FrameStrobe[11]
+ Tile_X1Y6_LUT4AB/FrameStrobe[12] Tile_X1Y6_LUT4AB/FrameStrobe[13] Tile_X1Y6_LUT4AB/FrameStrobe[14]
+ Tile_X1Y6_LUT4AB/FrameStrobe[15] Tile_X1Y6_LUT4AB/FrameStrobe[16] Tile_X1Y6_LUT4AB/FrameStrobe[17]
+ Tile_X1Y6_LUT4AB/FrameStrobe[18] Tile_X1Y6_LUT4AB/FrameStrobe[19] Tile_X1Y6_LUT4AB/FrameStrobe[1]
+ Tile_X1Y6_LUT4AB/FrameStrobe[2] Tile_X1Y6_LUT4AB/FrameStrobe[3] Tile_X1Y6_LUT4AB/FrameStrobe[4]
+ Tile_X1Y6_LUT4AB/FrameStrobe[5] Tile_X1Y6_LUT4AB/FrameStrobe[6] Tile_X1Y6_LUT4AB/FrameStrobe[7]
+ Tile_X1Y6_LUT4AB/FrameStrobe[8] Tile_X1Y6_LUT4AB/FrameStrobe[9] Tile_X1Y7_LUT4AB/N1BEG[0]
+ Tile_X1Y7_LUT4AB/N1BEG[1] Tile_X1Y7_LUT4AB/N1BEG[2] Tile_X1Y7_LUT4AB/N1BEG[3] Tile_X1Y8_LUT4AB/N1BEG[0]
+ Tile_X1Y8_LUT4AB/N1BEG[1] Tile_X1Y8_LUT4AB/N1BEG[2] Tile_X1Y8_LUT4AB/N1BEG[3] Tile_X1Y7_LUT4AB/N2BEG[0]
+ Tile_X1Y7_LUT4AB/N2BEG[1] Tile_X1Y7_LUT4AB/N2BEG[2] Tile_X1Y7_LUT4AB/N2BEG[3] Tile_X1Y7_LUT4AB/N2BEG[4]
+ Tile_X1Y7_LUT4AB/N2BEG[5] Tile_X1Y7_LUT4AB/N2BEG[6] Tile_X1Y7_LUT4AB/N2BEG[7] Tile_X1Y6_LUT4AB/N2END[0]
+ Tile_X1Y6_LUT4AB/N2END[1] Tile_X1Y6_LUT4AB/N2END[2] Tile_X1Y6_LUT4AB/N2END[3] Tile_X1Y6_LUT4AB/N2END[4]
+ Tile_X1Y6_LUT4AB/N2END[5] Tile_X1Y6_LUT4AB/N2END[6] Tile_X1Y6_LUT4AB/N2END[7] Tile_X1Y7_LUT4AB/N2END[0]
+ Tile_X1Y7_LUT4AB/N2END[1] Tile_X1Y7_LUT4AB/N2END[2] Tile_X1Y7_LUT4AB/N2END[3] Tile_X1Y7_LUT4AB/N2END[4]
+ Tile_X1Y7_LUT4AB/N2END[5] Tile_X1Y7_LUT4AB/N2END[6] Tile_X1Y7_LUT4AB/N2END[7] Tile_X1Y8_LUT4AB/N2BEG[0]
+ Tile_X1Y8_LUT4AB/N2BEG[1] Tile_X1Y8_LUT4AB/N2BEG[2] Tile_X1Y8_LUT4AB/N2BEG[3] Tile_X1Y8_LUT4AB/N2BEG[4]
+ Tile_X1Y8_LUT4AB/N2BEG[5] Tile_X1Y8_LUT4AB/N2BEG[6] Tile_X1Y8_LUT4AB/N2BEG[7] Tile_X1Y7_LUT4AB/N4BEG[0]
+ Tile_X1Y7_LUT4AB/N4BEG[10] Tile_X1Y7_LUT4AB/N4BEG[11] Tile_X1Y7_LUT4AB/N4BEG[12]
+ Tile_X1Y7_LUT4AB/N4BEG[13] Tile_X1Y7_LUT4AB/N4BEG[14] Tile_X1Y7_LUT4AB/N4BEG[15]
+ Tile_X1Y7_LUT4AB/N4BEG[1] Tile_X1Y7_LUT4AB/N4BEG[2] Tile_X1Y7_LUT4AB/N4BEG[3] Tile_X1Y7_LUT4AB/N4BEG[4]
+ Tile_X1Y7_LUT4AB/N4BEG[5] Tile_X1Y7_LUT4AB/N4BEG[6] Tile_X1Y7_LUT4AB/N4BEG[7] Tile_X1Y7_LUT4AB/N4BEG[8]
+ Tile_X1Y7_LUT4AB/N4BEG[9] Tile_X1Y8_LUT4AB/N4BEG[0] Tile_X1Y8_LUT4AB/N4BEG[10] Tile_X1Y8_LUT4AB/N4BEG[11]
+ Tile_X1Y8_LUT4AB/N4BEG[12] Tile_X1Y8_LUT4AB/N4BEG[13] Tile_X1Y8_LUT4AB/N4BEG[14]
+ Tile_X1Y8_LUT4AB/N4BEG[15] Tile_X1Y8_LUT4AB/N4BEG[1] Tile_X1Y8_LUT4AB/N4BEG[2] Tile_X1Y8_LUT4AB/N4BEG[3]
+ Tile_X1Y8_LUT4AB/N4BEG[4] Tile_X1Y8_LUT4AB/N4BEG[5] Tile_X1Y8_LUT4AB/N4BEG[6] Tile_X1Y8_LUT4AB/N4BEG[7]
+ Tile_X1Y8_LUT4AB/N4BEG[8] Tile_X1Y8_LUT4AB/N4BEG[9] Tile_X1Y7_LUT4AB/NN4BEG[0] Tile_X1Y7_LUT4AB/NN4BEG[10]
+ Tile_X1Y7_LUT4AB/NN4BEG[11] Tile_X1Y7_LUT4AB/NN4BEG[12] Tile_X1Y7_LUT4AB/NN4BEG[13]
+ Tile_X1Y7_LUT4AB/NN4BEG[14] Tile_X1Y7_LUT4AB/NN4BEG[15] Tile_X1Y7_LUT4AB/NN4BEG[1]
+ Tile_X1Y7_LUT4AB/NN4BEG[2] Tile_X1Y7_LUT4AB/NN4BEG[3] Tile_X1Y7_LUT4AB/NN4BEG[4]
+ Tile_X1Y7_LUT4AB/NN4BEG[5] Tile_X1Y7_LUT4AB/NN4BEG[6] Tile_X1Y7_LUT4AB/NN4BEG[7]
+ Tile_X1Y7_LUT4AB/NN4BEG[8] Tile_X1Y7_LUT4AB/NN4BEG[9] Tile_X1Y8_LUT4AB/NN4BEG[0]
+ Tile_X1Y8_LUT4AB/NN4BEG[10] Tile_X1Y8_LUT4AB/NN4BEG[11] Tile_X1Y8_LUT4AB/NN4BEG[12]
+ Tile_X1Y8_LUT4AB/NN4BEG[13] Tile_X1Y8_LUT4AB/NN4BEG[14] Tile_X1Y8_LUT4AB/NN4BEG[15]
+ Tile_X1Y8_LUT4AB/NN4BEG[1] Tile_X1Y8_LUT4AB/NN4BEG[2] Tile_X1Y8_LUT4AB/NN4BEG[3]
+ Tile_X1Y8_LUT4AB/NN4BEG[4] Tile_X1Y8_LUT4AB/NN4BEG[5] Tile_X1Y8_LUT4AB/NN4BEG[6]
+ Tile_X1Y8_LUT4AB/NN4BEG[7] Tile_X1Y8_LUT4AB/NN4BEG[8] Tile_X1Y8_LUT4AB/NN4BEG[9]
+ Tile_X1Y8_LUT4AB/S1END[0] Tile_X1Y8_LUT4AB/S1END[1] Tile_X1Y8_LUT4AB/S1END[2] Tile_X1Y8_LUT4AB/S1END[3]
+ Tile_X1Y7_LUT4AB/S1END[0] Tile_X1Y7_LUT4AB/S1END[1] Tile_X1Y7_LUT4AB/S1END[2] Tile_X1Y7_LUT4AB/S1END[3]
+ Tile_X1Y8_LUT4AB/S2MID[0] Tile_X1Y8_LUT4AB/S2MID[1] Tile_X1Y8_LUT4AB/S2MID[2] Tile_X1Y8_LUT4AB/S2MID[3]
+ Tile_X1Y8_LUT4AB/S2MID[4] Tile_X1Y8_LUT4AB/S2MID[5] Tile_X1Y8_LUT4AB/S2MID[6] Tile_X1Y8_LUT4AB/S2MID[7]
+ Tile_X1Y8_LUT4AB/S2END[0] Tile_X1Y8_LUT4AB/S2END[1] Tile_X1Y8_LUT4AB/S2END[2] Tile_X1Y8_LUT4AB/S2END[3]
+ Tile_X1Y8_LUT4AB/S2END[4] Tile_X1Y8_LUT4AB/S2END[5] Tile_X1Y8_LUT4AB/S2END[6] Tile_X1Y8_LUT4AB/S2END[7]
+ Tile_X1Y7_LUT4AB/S2END[0] Tile_X1Y7_LUT4AB/S2END[1] Tile_X1Y7_LUT4AB/S2END[2] Tile_X1Y7_LUT4AB/S2END[3]
+ Tile_X1Y7_LUT4AB/S2END[4] Tile_X1Y7_LUT4AB/S2END[5] Tile_X1Y7_LUT4AB/S2END[6] Tile_X1Y7_LUT4AB/S2END[7]
+ Tile_X1Y7_LUT4AB/S2MID[0] Tile_X1Y7_LUT4AB/S2MID[1] Tile_X1Y7_LUT4AB/S2MID[2] Tile_X1Y7_LUT4AB/S2MID[3]
+ Tile_X1Y7_LUT4AB/S2MID[4] Tile_X1Y7_LUT4AB/S2MID[5] Tile_X1Y7_LUT4AB/S2MID[6] Tile_X1Y7_LUT4AB/S2MID[7]
+ Tile_X1Y8_LUT4AB/S4END[0] Tile_X1Y8_LUT4AB/S4END[10] Tile_X1Y8_LUT4AB/S4END[11]
+ Tile_X1Y8_LUT4AB/S4END[12] Tile_X1Y8_LUT4AB/S4END[13] Tile_X1Y8_LUT4AB/S4END[14]
+ Tile_X1Y8_LUT4AB/S4END[15] Tile_X1Y8_LUT4AB/S4END[1] Tile_X1Y8_LUT4AB/S4END[2] Tile_X1Y8_LUT4AB/S4END[3]
+ Tile_X1Y8_LUT4AB/S4END[4] Tile_X1Y8_LUT4AB/S4END[5] Tile_X1Y8_LUT4AB/S4END[6] Tile_X1Y8_LUT4AB/S4END[7]
+ Tile_X1Y8_LUT4AB/S4END[8] Tile_X1Y8_LUT4AB/S4END[9] Tile_X1Y7_LUT4AB/S4END[0] Tile_X1Y7_LUT4AB/S4END[10]
+ Tile_X1Y7_LUT4AB/S4END[11] Tile_X1Y7_LUT4AB/S4END[12] Tile_X1Y7_LUT4AB/S4END[13]
+ Tile_X1Y7_LUT4AB/S4END[14] Tile_X1Y7_LUT4AB/S4END[15] Tile_X1Y7_LUT4AB/S4END[1]
+ Tile_X1Y7_LUT4AB/S4END[2] Tile_X1Y7_LUT4AB/S4END[3] Tile_X1Y7_LUT4AB/S4END[4] Tile_X1Y7_LUT4AB/S4END[5]
+ Tile_X1Y7_LUT4AB/S4END[6] Tile_X1Y7_LUT4AB/S4END[7] Tile_X1Y7_LUT4AB/S4END[8] Tile_X1Y7_LUT4AB/S4END[9]
+ Tile_X1Y8_LUT4AB/SS4END[0] Tile_X1Y8_LUT4AB/SS4END[10] Tile_X1Y8_LUT4AB/SS4END[11]
+ Tile_X1Y8_LUT4AB/SS4END[12] Tile_X1Y8_LUT4AB/SS4END[13] Tile_X1Y8_LUT4AB/SS4END[14]
+ Tile_X1Y8_LUT4AB/SS4END[15] Tile_X1Y8_LUT4AB/SS4END[1] Tile_X1Y8_LUT4AB/SS4END[2]
+ Tile_X1Y8_LUT4AB/SS4END[3] Tile_X1Y8_LUT4AB/SS4END[4] Tile_X1Y8_LUT4AB/SS4END[5]
+ Tile_X1Y8_LUT4AB/SS4END[6] Tile_X1Y8_LUT4AB/SS4END[7] Tile_X1Y8_LUT4AB/SS4END[8]
+ Tile_X1Y8_LUT4AB/SS4END[9] Tile_X1Y7_LUT4AB/SS4END[0] Tile_X1Y7_LUT4AB/SS4END[10]
+ Tile_X1Y7_LUT4AB/SS4END[11] Tile_X1Y7_LUT4AB/SS4END[12] Tile_X1Y7_LUT4AB/SS4END[13]
+ Tile_X1Y7_LUT4AB/SS4END[14] Tile_X1Y7_LUT4AB/SS4END[15] Tile_X1Y7_LUT4AB/SS4END[1]
+ Tile_X1Y7_LUT4AB/SS4END[2] Tile_X1Y7_LUT4AB/SS4END[3] Tile_X1Y7_LUT4AB/SS4END[4]
+ Tile_X1Y7_LUT4AB/SS4END[5] Tile_X1Y7_LUT4AB/SS4END[6] Tile_X1Y7_LUT4AB/SS4END[7]
+ Tile_X1Y7_LUT4AB/SS4END[8] Tile_X1Y7_LUT4AB/SS4END[9] Tile_X1Y7_LUT4AB/UserCLK Tile_X1Y6_LUT4AB/UserCLK
+ VGND VPWR Tile_X1Y7_LUT4AB/W1BEG[0] Tile_X1Y7_LUT4AB/W1BEG[1] Tile_X1Y7_LUT4AB/W1BEG[2]
+ Tile_X1Y7_LUT4AB/W1BEG[3] Tile_X2Y7_LUT4AB/W1BEG[0] Tile_X2Y7_LUT4AB/W1BEG[1] Tile_X2Y7_LUT4AB/W1BEG[2]
+ Tile_X2Y7_LUT4AB/W1BEG[3] Tile_X1Y7_LUT4AB/W2BEG[0] Tile_X1Y7_LUT4AB/W2BEG[1] Tile_X1Y7_LUT4AB/W2BEG[2]
+ Tile_X1Y7_LUT4AB/W2BEG[3] Tile_X1Y7_LUT4AB/W2BEG[4] Tile_X1Y7_LUT4AB/W2BEG[5] Tile_X1Y7_LUT4AB/W2BEG[6]
+ Tile_X1Y7_LUT4AB/W2BEG[7] Tile_X1Y7_LUT4AB/W2BEGb[0] Tile_X1Y7_LUT4AB/W2BEGb[1]
+ Tile_X1Y7_LUT4AB/W2BEGb[2] Tile_X1Y7_LUT4AB/W2BEGb[3] Tile_X1Y7_LUT4AB/W2BEGb[4]
+ Tile_X1Y7_LUT4AB/W2BEGb[5] Tile_X1Y7_LUT4AB/W2BEGb[6] Tile_X1Y7_LUT4AB/W2BEGb[7]
+ Tile_X1Y7_LUT4AB/W2END[0] Tile_X1Y7_LUT4AB/W2END[1] Tile_X1Y7_LUT4AB/W2END[2] Tile_X1Y7_LUT4AB/W2END[3]
+ Tile_X1Y7_LUT4AB/W2END[4] Tile_X1Y7_LUT4AB/W2END[5] Tile_X1Y7_LUT4AB/W2END[6] Tile_X1Y7_LUT4AB/W2END[7]
+ Tile_X2Y7_LUT4AB/W2BEG[0] Tile_X2Y7_LUT4AB/W2BEG[1] Tile_X2Y7_LUT4AB/W2BEG[2] Tile_X2Y7_LUT4AB/W2BEG[3]
+ Tile_X2Y7_LUT4AB/W2BEG[4] Tile_X2Y7_LUT4AB/W2BEG[5] Tile_X2Y7_LUT4AB/W2BEG[6] Tile_X2Y7_LUT4AB/W2BEG[7]
+ Tile_X1Y7_LUT4AB/W6BEG[0] Tile_X1Y7_LUT4AB/W6BEG[10] Tile_X1Y7_LUT4AB/W6BEG[11]
+ Tile_X1Y7_LUT4AB/W6BEG[1] Tile_X1Y7_LUT4AB/W6BEG[2] Tile_X1Y7_LUT4AB/W6BEG[3] Tile_X1Y7_LUT4AB/W6BEG[4]
+ Tile_X1Y7_LUT4AB/W6BEG[5] Tile_X1Y7_LUT4AB/W6BEG[6] Tile_X1Y7_LUT4AB/W6BEG[7] Tile_X1Y7_LUT4AB/W6BEG[8]
+ Tile_X1Y7_LUT4AB/W6BEG[9] Tile_X2Y7_LUT4AB/W6BEG[0] Tile_X2Y7_LUT4AB/W6BEG[10] Tile_X2Y7_LUT4AB/W6BEG[11]
+ Tile_X2Y7_LUT4AB/W6BEG[1] Tile_X2Y7_LUT4AB/W6BEG[2] Tile_X2Y7_LUT4AB/W6BEG[3] Tile_X2Y7_LUT4AB/W6BEG[4]
+ Tile_X2Y7_LUT4AB/W6BEG[5] Tile_X2Y7_LUT4AB/W6BEG[6] Tile_X2Y7_LUT4AB/W6BEG[7] Tile_X2Y7_LUT4AB/W6BEG[8]
+ Tile_X2Y7_LUT4AB/W6BEG[9] Tile_X1Y7_LUT4AB/WW4BEG[0] Tile_X1Y7_LUT4AB/WW4BEG[10]
+ Tile_X1Y7_LUT4AB/WW4BEG[11] Tile_X1Y7_LUT4AB/WW4BEG[12] Tile_X1Y7_LUT4AB/WW4BEG[13]
+ Tile_X1Y7_LUT4AB/WW4BEG[14] Tile_X1Y7_LUT4AB/WW4BEG[15] Tile_X1Y7_LUT4AB/WW4BEG[1]
+ Tile_X1Y7_LUT4AB/WW4BEG[2] Tile_X1Y7_LUT4AB/WW4BEG[3] Tile_X1Y7_LUT4AB/WW4BEG[4]
+ Tile_X1Y7_LUT4AB/WW4BEG[5] Tile_X1Y7_LUT4AB/WW4BEG[6] Tile_X1Y7_LUT4AB/WW4BEG[7]
+ Tile_X1Y7_LUT4AB/WW4BEG[8] Tile_X1Y7_LUT4AB/WW4BEG[9] Tile_X2Y7_LUT4AB/WW4BEG[0]
+ Tile_X2Y7_LUT4AB/WW4BEG[10] Tile_X2Y7_LUT4AB/WW4BEG[11] Tile_X2Y7_LUT4AB/WW4BEG[12]
+ Tile_X2Y7_LUT4AB/WW4BEG[13] Tile_X2Y7_LUT4AB/WW4BEG[14] Tile_X2Y7_LUT4AB/WW4BEG[15]
+ Tile_X2Y7_LUT4AB/WW4BEG[1] Tile_X2Y7_LUT4AB/WW4BEG[2] Tile_X2Y7_LUT4AB/WW4BEG[3]
+ Tile_X2Y7_LUT4AB/WW4BEG[4] Tile_X2Y7_LUT4AB/WW4BEG[5] Tile_X2Y7_LUT4AB/WW4BEG[6]
+ Tile_X2Y7_LUT4AB/WW4BEG[7] Tile_X2Y7_LUT4AB/WW4BEG[8] Tile_X2Y7_LUT4AB/WW4BEG[9]
+ LUT4AB
XTile_X4Y1_LUT4AB Tile_X4Y2_LUT4AB/Co Tile_X4Y0_N_IO4/Ci Tile_X4Y1_LUT4AB/E1BEG[0]
+ Tile_X4Y1_LUT4AB/E1BEG[1] Tile_X4Y1_LUT4AB/E1BEG[2] Tile_X4Y1_LUT4AB/E1BEG[3] Tile_X4Y1_LUT4AB/E1END[0]
+ Tile_X4Y1_LUT4AB/E1END[1] Tile_X4Y1_LUT4AB/E1END[2] Tile_X4Y1_LUT4AB/E1END[3] Tile_X4Y1_LUT4AB/E2BEG[0]
+ Tile_X4Y1_LUT4AB/E2BEG[1] Tile_X4Y1_LUT4AB/E2BEG[2] Tile_X4Y1_LUT4AB/E2BEG[3] Tile_X4Y1_LUT4AB/E2BEG[4]
+ Tile_X4Y1_LUT4AB/E2BEG[5] Tile_X4Y1_LUT4AB/E2BEG[6] Tile_X4Y1_LUT4AB/E2BEG[7] Tile_X4Y1_LUT4AB/E2BEGb[0]
+ Tile_X4Y1_LUT4AB/E2BEGb[1] Tile_X4Y1_LUT4AB/E2BEGb[2] Tile_X4Y1_LUT4AB/E2BEGb[3]
+ Tile_X4Y1_LUT4AB/E2BEGb[4] Tile_X4Y1_LUT4AB/E2BEGb[5] Tile_X4Y1_LUT4AB/E2BEGb[6]
+ Tile_X4Y1_LUT4AB/E2BEGb[7] Tile_X4Y1_LUT4AB/E2END[0] Tile_X4Y1_LUT4AB/E2END[1] Tile_X4Y1_LUT4AB/E2END[2]
+ Tile_X4Y1_LUT4AB/E2END[3] Tile_X4Y1_LUT4AB/E2END[4] Tile_X4Y1_LUT4AB/E2END[5] Tile_X4Y1_LUT4AB/E2END[6]
+ Tile_X4Y1_LUT4AB/E2END[7] Tile_X4Y1_LUT4AB/E2MID[0] Tile_X4Y1_LUT4AB/E2MID[1] Tile_X4Y1_LUT4AB/E2MID[2]
+ Tile_X4Y1_LUT4AB/E2MID[3] Tile_X4Y1_LUT4AB/E2MID[4] Tile_X4Y1_LUT4AB/E2MID[5] Tile_X4Y1_LUT4AB/E2MID[6]
+ Tile_X4Y1_LUT4AB/E2MID[7] Tile_X4Y1_LUT4AB/E6BEG[0] Tile_X4Y1_LUT4AB/E6BEG[10] Tile_X4Y1_LUT4AB/E6BEG[11]
+ Tile_X4Y1_LUT4AB/E6BEG[1] Tile_X4Y1_LUT4AB/E6BEG[2] Tile_X4Y1_LUT4AB/E6BEG[3] Tile_X4Y1_LUT4AB/E6BEG[4]
+ Tile_X4Y1_LUT4AB/E6BEG[5] Tile_X4Y1_LUT4AB/E6BEG[6] Tile_X4Y1_LUT4AB/E6BEG[7] Tile_X4Y1_LUT4AB/E6BEG[8]
+ Tile_X4Y1_LUT4AB/E6BEG[9] Tile_X4Y1_LUT4AB/E6END[0] Tile_X4Y1_LUT4AB/E6END[10] Tile_X4Y1_LUT4AB/E6END[11]
+ Tile_X4Y1_LUT4AB/E6END[1] Tile_X4Y1_LUT4AB/E6END[2] Tile_X4Y1_LUT4AB/E6END[3] Tile_X4Y1_LUT4AB/E6END[4]
+ Tile_X4Y1_LUT4AB/E6END[5] Tile_X4Y1_LUT4AB/E6END[6] Tile_X4Y1_LUT4AB/E6END[7] Tile_X4Y1_LUT4AB/E6END[8]
+ Tile_X4Y1_LUT4AB/E6END[9] Tile_X4Y1_LUT4AB/EE4BEG[0] Tile_X4Y1_LUT4AB/EE4BEG[10]
+ Tile_X4Y1_LUT4AB/EE4BEG[11] Tile_X4Y1_LUT4AB/EE4BEG[12] Tile_X4Y1_LUT4AB/EE4BEG[13]
+ Tile_X4Y1_LUT4AB/EE4BEG[14] Tile_X4Y1_LUT4AB/EE4BEG[15] Tile_X4Y1_LUT4AB/EE4BEG[1]
+ Tile_X4Y1_LUT4AB/EE4BEG[2] Tile_X4Y1_LUT4AB/EE4BEG[3] Tile_X4Y1_LUT4AB/EE4BEG[4]
+ Tile_X4Y1_LUT4AB/EE4BEG[5] Tile_X4Y1_LUT4AB/EE4BEG[6] Tile_X4Y1_LUT4AB/EE4BEG[7]
+ Tile_X4Y1_LUT4AB/EE4BEG[8] Tile_X4Y1_LUT4AB/EE4BEG[9] Tile_X4Y1_LUT4AB/EE4END[0]
+ Tile_X4Y1_LUT4AB/EE4END[10] Tile_X4Y1_LUT4AB/EE4END[11] Tile_X4Y1_LUT4AB/EE4END[12]
+ Tile_X4Y1_LUT4AB/EE4END[13] Tile_X4Y1_LUT4AB/EE4END[14] Tile_X4Y1_LUT4AB/EE4END[15]
+ Tile_X4Y1_LUT4AB/EE4END[1] Tile_X4Y1_LUT4AB/EE4END[2] Tile_X4Y1_LUT4AB/EE4END[3]
+ Tile_X4Y1_LUT4AB/EE4END[4] Tile_X4Y1_LUT4AB/EE4END[5] Tile_X4Y1_LUT4AB/EE4END[6]
+ Tile_X4Y1_LUT4AB/EE4END[7] Tile_X4Y1_LUT4AB/EE4END[8] Tile_X4Y1_LUT4AB/EE4END[9]
+ Tile_X4Y1_LUT4AB/FrameData[0] Tile_X4Y1_LUT4AB/FrameData[10] Tile_X4Y1_LUT4AB/FrameData[11]
+ Tile_X4Y1_LUT4AB/FrameData[12] Tile_X4Y1_LUT4AB/FrameData[13] Tile_X4Y1_LUT4AB/FrameData[14]
+ Tile_X4Y1_LUT4AB/FrameData[15] Tile_X4Y1_LUT4AB/FrameData[16] Tile_X4Y1_LUT4AB/FrameData[17]
+ Tile_X4Y1_LUT4AB/FrameData[18] Tile_X4Y1_LUT4AB/FrameData[19] Tile_X4Y1_LUT4AB/FrameData[1]
+ Tile_X4Y1_LUT4AB/FrameData[20] Tile_X4Y1_LUT4AB/FrameData[21] Tile_X4Y1_LUT4AB/FrameData[22]
+ Tile_X4Y1_LUT4AB/FrameData[23] Tile_X4Y1_LUT4AB/FrameData[24] Tile_X4Y1_LUT4AB/FrameData[25]
+ Tile_X4Y1_LUT4AB/FrameData[26] Tile_X4Y1_LUT4AB/FrameData[27] Tile_X4Y1_LUT4AB/FrameData[28]
+ Tile_X4Y1_LUT4AB/FrameData[29] Tile_X4Y1_LUT4AB/FrameData[2] Tile_X4Y1_LUT4AB/FrameData[30]
+ Tile_X4Y1_LUT4AB/FrameData[31] Tile_X4Y1_LUT4AB/FrameData[3] Tile_X4Y1_LUT4AB/FrameData[4]
+ Tile_X4Y1_LUT4AB/FrameData[5] Tile_X4Y1_LUT4AB/FrameData[6] Tile_X4Y1_LUT4AB/FrameData[7]
+ Tile_X4Y1_LUT4AB/FrameData[8] Tile_X4Y1_LUT4AB/FrameData[9] Tile_X4Y1_LUT4AB/FrameData_O[0]
+ Tile_X4Y1_LUT4AB/FrameData_O[10] Tile_X4Y1_LUT4AB/FrameData_O[11] Tile_X4Y1_LUT4AB/FrameData_O[12]
+ Tile_X4Y1_LUT4AB/FrameData_O[13] Tile_X4Y1_LUT4AB/FrameData_O[14] Tile_X4Y1_LUT4AB/FrameData_O[15]
+ Tile_X4Y1_LUT4AB/FrameData_O[16] Tile_X4Y1_LUT4AB/FrameData_O[17] Tile_X4Y1_LUT4AB/FrameData_O[18]
+ Tile_X4Y1_LUT4AB/FrameData_O[19] Tile_X4Y1_LUT4AB/FrameData_O[1] Tile_X4Y1_LUT4AB/FrameData_O[20]
+ Tile_X4Y1_LUT4AB/FrameData_O[21] Tile_X4Y1_LUT4AB/FrameData_O[22] Tile_X4Y1_LUT4AB/FrameData_O[23]
+ Tile_X4Y1_LUT4AB/FrameData_O[24] Tile_X4Y1_LUT4AB/FrameData_O[25] Tile_X4Y1_LUT4AB/FrameData_O[26]
+ Tile_X4Y1_LUT4AB/FrameData_O[27] Tile_X4Y1_LUT4AB/FrameData_O[28] Tile_X4Y1_LUT4AB/FrameData_O[29]
+ Tile_X4Y1_LUT4AB/FrameData_O[2] Tile_X4Y1_LUT4AB/FrameData_O[30] Tile_X4Y1_LUT4AB/FrameData_O[31]
+ Tile_X4Y1_LUT4AB/FrameData_O[3] Tile_X4Y1_LUT4AB/FrameData_O[4] Tile_X4Y1_LUT4AB/FrameData_O[5]
+ Tile_X4Y1_LUT4AB/FrameData_O[6] Tile_X4Y1_LUT4AB/FrameData_O[7] Tile_X4Y1_LUT4AB/FrameData_O[8]
+ Tile_X4Y1_LUT4AB/FrameData_O[9] Tile_X4Y1_LUT4AB/FrameStrobe[0] Tile_X4Y1_LUT4AB/FrameStrobe[10]
+ Tile_X4Y1_LUT4AB/FrameStrobe[11] Tile_X4Y1_LUT4AB/FrameStrobe[12] Tile_X4Y1_LUT4AB/FrameStrobe[13]
+ Tile_X4Y1_LUT4AB/FrameStrobe[14] Tile_X4Y1_LUT4AB/FrameStrobe[15] Tile_X4Y1_LUT4AB/FrameStrobe[16]
+ Tile_X4Y1_LUT4AB/FrameStrobe[17] Tile_X4Y1_LUT4AB/FrameStrobe[18] Tile_X4Y1_LUT4AB/FrameStrobe[19]
+ Tile_X4Y1_LUT4AB/FrameStrobe[1] Tile_X4Y1_LUT4AB/FrameStrobe[2] Tile_X4Y1_LUT4AB/FrameStrobe[3]
+ Tile_X4Y1_LUT4AB/FrameStrobe[4] Tile_X4Y1_LUT4AB/FrameStrobe[5] Tile_X4Y1_LUT4AB/FrameStrobe[6]
+ Tile_X4Y1_LUT4AB/FrameStrobe[7] Tile_X4Y1_LUT4AB/FrameStrobe[8] Tile_X4Y1_LUT4AB/FrameStrobe[9]
+ Tile_X4Y0_N_IO4/FrameStrobe[0] Tile_X4Y0_N_IO4/FrameStrobe[10] Tile_X4Y0_N_IO4/FrameStrobe[11]
+ Tile_X4Y0_N_IO4/FrameStrobe[12] Tile_X4Y0_N_IO4/FrameStrobe[13] Tile_X4Y0_N_IO4/FrameStrobe[14]
+ Tile_X4Y0_N_IO4/FrameStrobe[15] Tile_X4Y0_N_IO4/FrameStrobe[16] Tile_X4Y0_N_IO4/FrameStrobe[17]
+ Tile_X4Y0_N_IO4/FrameStrobe[18] Tile_X4Y0_N_IO4/FrameStrobe[19] Tile_X4Y0_N_IO4/FrameStrobe[1]
+ Tile_X4Y0_N_IO4/FrameStrobe[2] Tile_X4Y0_N_IO4/FrameStrobe[3] Tile_X4Y0_N_IO4/FrameStrobe[4]
+ Tile_X4Y0_N_IO4/FrameStrobe[5] Tile_X4Y0_N_IO4/FrameStrobe[6] Tile_X4Y0_N_IO4/FrameStrobe[7]
+ Tile_X4Y0_N_IO4/FrameStrobe[8] Tile_X4Y0_N_IO4/FrameStrobe[9] Tile_X4Y0_N_IO4/N1END[0]
+ Tile_X4Y0_N_IO4/N1END[1] Tile_X4Y0_N_IO4/N1END[2] Tile_X4Y0_N_IO4/N1END[3] Tile_X4Y2_LUT4AB/N1BEG[0]
+ Tile_X4Y2_LUT4AB/N1BEG[1] Tile_X4Y2_LUT4AB/N1BEG[2] Tile_X4Y2_LUT4AB/N1BEG[3] Tile_X4Y0_N_IO4/N2MID[0]
+ Tile_X4Y0_N_IO4/N2MID[1] Tile_X4Y0_N_IO4/N2MID[2] Tile_X4Y0_N_IO4/N2MID[3] Tile_X4Y0_N_IO4/N2MID[4]
+ Tile_X4Y0_N_IO4/N2MID[5] Tile_X4Y0_N_IO4/N2MID[6] Tile_X4Y0_N_IO4/N2MID[7] Tile_X4Y0_N_IO4/N2END[0]
+ Tile_X4Y0_N_IO4/N2END[1] Tile_X4Y0_N_IO4/N2END[2] Tile_X4Y0_N_IO4/N2END[3] Tile_X4Y0_N_IO4/N2END[4]
+ Tile_X4Y0_N_IO4/N2END[5] Tile_X4Y0_N_IO4/N2END[6] Tile_X4Y0_N_IO4/N2END[7] Tile_X4Y1_LUT4AB/N2END[0]
+ Tile_X4Y1_LUT4AB/N2END[1] Tile_X4Y1_LUT4AB/N2END[2] Tile_X4Y1_LUT4AB/N2END[3] Tile_X4Y1_LUT4AB/N2END[4]
+ Tile_X4Y1_LUT4AB/N2END[5] Tile_X4Y1_LUT4AB/N2END[6] Tile_X4Y1_LUT4AB/N2END[7] Tile_X4Y2_LUT4AB/N2BEG[0]
+ Tile_X4Y2_LUT4AB/N2BEG[1] Tile_X4Y2_LUT4AB/N2BEG[2] Tile_X4Y2_LUT4AB/N2BEG[3] Tile_X4Y2_LUT4AB/N2BEG[4]
+ Tile_X4Y2_LUT4AB/N2BEG[5] Tile_X4Y2_LUT4AB/N2BEG[6] Tile_X4Y2_LUT4AB/N2BEG[7] Tile_X4Y0_N_IO4/N4END[0]
+ Tile_X4Y0_N_IO4/N4END[10] Tile_X4Y0_N_IO4/N4END[11] Tile_X4Y0_N_IO4/N4END[12] Tile_X4Y0_N_IO4/N4END[13]
+ Tile_X4Y0_N_IO4/N4END[14] Tile_X4Y0_N_IO4/N4END[15] Tile_X4Y0_N_IO4/N4END[1] Tile_X4Y0_N_IO4/N4END[2]
+ Tile_X4Y0_N_IO4/N4END[3] Tile_X4Y0_N_IO4/N4END[4] Tile_X4Y0_N_IO4/N4END[5] Tile_X4Y0_N_IO4/N4END[6]
+ Tile_X4Y0_N_IO4/N4END[7] Tile_X4Y0_N_IO4/N4END[8] Tile_X4Y0_N_IO4/N4END[9] Tile_X4Y2_LUT4AB/N4BEG[0]
+ Tile_X4Y2_LUT4AB/N4BEG[10] Tile_X4Y2_LUT4AB/N4BEG[11] Tile_X4Y2_LUT4AB/N4BEG[12]
+ Tile_X4Y2_LUT4AB/N4BEG[13] Tile_X4Y2_LUT4AB/N4BEG[14] Tile_X4Y2_LUT4AB/N4BEG[15]
+ Tile_X4Y2_LUT4AB/N4BEG[1] Tile_X4Y2_LUT4AB/N4BEG[2] Tile_X4Y2_LUT4AB/N4BEG[3] Tile_X4Y2_LUT4AB/N4BEG[4]
+ Tile_X4Y2_LUT4AB/N4BEG[5] Tile_X4Y2_LUT4AB/N4BEG[6] Tile_X4Y2_LUT4AB/N4BEG[7] Tile_X4Y2_LUT4AB/N4BEG[8]
+ Tile_X4Y2_LUT4AB/N4BEG[9] Tile_X4Y0_N_IO4/NN4END[0] Tile_X4Y0_N_IO4/NN4END[10] Tile_X4Y0_N_IO4/NN4END[11]
+ Tile_X4Y0_N_IO4/NN4END[12] Tile_X4Y0_N_IO4/NN4END[13] Tile_X4Y0_N_IO4/NN4END[14]
+ Tile_X4Y0_N_IO4/NN4END[15] Tile_X4Y0_N_IO4/NN4END[1] Tile_X4Y0_N_IO4/NN4END[2] Tile_X4Y0_N_IO4/NN4END[3]
+ Tile_X4Y0_N_IO4/NN4END[4] Tile_X4Y0_N_IO4/NN4END[5] Tile_X4Y0_N_IO4/NN4END[6] Tile_X4Y0_N_IO4/NN4END[7]
+ Tile_X4Y0_N_IO4/NN4END[8] Tile_X4Y0_N_IO4/NN4END[9] Tile_X4Y2_LUT4AB/NN4BEG[0] Tile_X4Y2_LUT4AB/NN4BEG[10]
+ Tile_X4Y2_LUT4AB/NN4BEG[11] Tile_X4Y2_LUT4AB/NN4BEG[12] Tile_X4Y2_LUT4AB/NN4BEG[13]
+ Tile_X4Y2_LUT4AB/NN4BEG[14] Tile_X4Y2_LUT4AB/NN4BEG[15] Tile_X4Y2_LUT4AB/NN4BEG[1]
+ Tile_X4Y2_LUT4AB/NN4BEG[2] Tile_X4Y2_LUT4AB/NN4BEG[3] Tile_X4Y2_LUT4AB/NN4BEG[4]
+ Tile_X4Y2_LUT4AB/NN4BEG[5] Tile_X4Y2_LUT4AB/NN4BEG[6] Tile_X4Y2_LUT4AB/NN4BEG[7]
+ Tile_X4Y2_LUT4AB/NN4BEG[8] Tile_X4Y2_LUT4AB/NN4BEG[9] Tile_X4Y2_LUT4AB/S1END[0]
+ Tile_X4Y2_LUT4AB/S1END[1] Tile_X4Y2_LUT4AB/S1END[2] Tile_X4Y2_LUT4AB/S1END[3] Tile_X4Y0_N_IO4/S1BEG[0]
+ Tile_X4Y0_N_IO4/S1BEG[1] Tile_X4Y0_N_IO4/S1BEG[2] Tile_X4Y0_N_IO4/S1BEG[3] Tile_X4Y2_LUT4AB/S2MID[0]
+ Tile_X4Y2_LUT4AB/S2MID[1] Tile_X4Y2_LUT4AB/S2MID[2] Tile_X4Y2_LUT4AB/S2MID[3] Tile_X4Y2_LUT4AB/S2MID[4]
+ Tile_X4Y2_LUT4AB/S2MID[5] Tile_X4Y2_LUT4AB/S2MID[6] Tile_X4Y2_LUT4AB/S2MID[7] Tile_X4Y2_LUT4AB/S2END[0]
+ Tile_X4Y2_LUT4AB/S2END[1] Tile_X4Y2_LUT4AB/S2END[2] Tile_X4Y2_LUT4AB/S2END[3] Tile_X4Y2_LUT4AB/S2END[4]
+ Tile_X4Y2_LUT4AB/S2END[5] Tile_X4Y2_LUT4AB/S2END[6] Tile_X4Y2_LUT4AB/S2END[7] Tile_X4Y1_LUT4AB/S2END[0]
+ Tile_X4Y1_LUT4AB/S2END[1] Tile_X4Y1_LUT4AB/S2END[2] Tile_X4Y1_LUT4AB/S2END[3] Tile_X4Y1_LUT4AB/S2END[4]
+ Tile_X4Y1_LUT4AB/S2END[5] Tile_X4Y1_LUT4AB/S2END[6] Tile_X4Y1_LUT4AB/S2END[7] Tile_X4Y0_N_IO4/S2BEG[0]
+ Tile_X4Y0_N_IO4/S2BEG[1] Tile_X4Y0_N_IO4/S2BEG[2] Tile_X4Y0_N_IO4/S2BEG[3] Tile_X4Y0_N_IO4/S2BEG[4]
+ Tile_X4Y0_N_IO4/S2BEG[5] Tile_X4Y0_N_IO4/S2BEG[6] Tile_X4Y0_N_IO4/S2BEG[7] Tile_X4Y2_LUT4AB/S4END[0]
+ Tile_X4Y2_LUT4AB/S4END[10] Tile_X4Y2_LUT4AB/S4END[11] Tile_X4Y2_LUT4AB/S4END[12]
+ Tile_X4Y2_LUT4AB/S4END[13] Tile_X4Y2_LUT4AB/S4END[14] Tile_X4Y2_LUT4AB/S4END[15]
+ Tile_X4Y2_LUT4AB/S4END[1] Tile_X4Y2_LUT4AB/S4END[2] Tile_X4Y2_LUT4AB/S4END[3] Tile_X4Y2_LUT4AB/S4END[4]
+ Tile_X4Y2_LUT4AB/S4END[5] Tile_X4Y2_LUT4AB/S4END[6] Tile_X4Y2_LUT4AB/S4END[7] Tile_X4Y2_LUT4AB/S4END[8]
+ Tile_X4Y2_LUT4AB/S4END[9] Tile_X4Y0_N_IO4/S4BEG[0] Tile_X4Y0_N_IO4/S4BEG[10] Tile_X4Y0_N_IO4/S4BEG[11]
+ Tile_X4Y0_N_IO4/S4BEG[12] Tile_X4Y0_N_IO4/S4BEG[13] Tile_X4Y0_N_IO4/S4BEG[14] Tile_X4Y0_N_IO4/S4BEG[15]
+ Tile_X4Y0_N_IO4/S4BEG[1] Tile_X4Y0_N_IO4/S4BEG[2] Tile_X4Y0_N_IO4/S4BEG[3] Tile_X4Y0_N_IO4/S4BEG[4]
+ Tile_X4Y0_N_IO4/S4BEG[5] Tile_X4Y0_N_IO4/S4BEG[6] Tile_X4Y0_N_IO4/S4BEG[7] Tile_X4Y0_N_IO4/S4BEG[8]
+ Tile_X4Y0_N_IO4/S4BEG[9] Tile_X4Y2_LUT4AB/SS4END[0] Tile_X4Y2_LUT4AB/SS4END[10]
+ Tile_X4Y2_LUT4AB/SS4END[11] Tile_X4Y2_LUT4AB/SS4END[12] Tile_X4Y2_LUT4AB/SS4END[13]
+ Tile_X4Y2_LUT4AB/SS4END[14] Tile_X4Y2_LUT4AB/SS4END[15] Tile_X4Y2_LUT4AB/SS4END[1]
+ Tile_X4Y2_LUT4AB/SS4END[2] Tile_X4Y2_LUT4AB/SS4END[3] Tile_X4Y2_LUT4AB/SS4END[4]
+ Tile_X4Y2_LUT4AB/SS4END[5] Tile_X4Y2_LUT4AB/SS4END[6] Tile_X4Y2_LUT4AB/SS4END[7]
+ Tile_X4Y2_LUT4AB/SS4END[8] Tile_X4Y2_LUT4AB/SS4END[9] Tile_X4Y0_N_IO4/SS4BEG[0]
+ Tile_X4Y0_N_IO4/SS4BEG[10] Tile_X4Y0_N_IO4/SS4BEG[11] Tile_X4Y0_N_IO4/SS4BEG[12]
+ Tile_X4Y0_N_IO4/SS4BEG[13] Tile_X4Y0_N_IO4/SS4BEG[14] Tile_X4Y0_N_IO4/SS4BEG[15]
+ Tile_X4Y0_N_IO4/SS4BEG[1] Tile_X4Y0_N_IO4/SS4BEG[2] Tile_X4Y0_N_IO4/SS4BEG[3] Tile_X4Y0_N_IO4/SS4BEG[4]
+ Tile_X4Y0_N_IO4/SS4BEG[5] Tile_X4Y0_N_IO4/SS4BEG[6] Tile_X4Y0_N_IO4/SS4BEG[7] Tile_X4Y0_N_IO4/SS4BEG[8]
+ Tile_X4Y0_N_IO4/SS4BEG[9] Tile_X4Y1_LUT4AB/UserCLK Tile_X4Y0_N_IO4/UserCLK VGND
+ VPWR Tile_X4Y1_LUT4AB/W1BEG[0] Tile_X4Y1_LUT4AB/W1BEG[1] Tile_X4Y1_LUT4AB/W1BEG[2]
+ Tile_X4Y1_LUT4AB/W1BEG[3] Tile_X4Y1_LUT4AB/W1END[0] Tile_X4Y1_LUT4AB/W1END[1] Tile_X4Y1_LUT4AB/W1END[2]
+ Tile_X4Y1_LUT4AB/W1END[3] Tile_X4Y1_LUT4AB/W2BEG[0] Tile_X4Y1_LUT4AB/W2BEG[1] Tile_X4Y1_LUT4AB/W2BEG[2]
+ Tile_X4Y1_LUT4AB/W2BEG[3] Tile_X4Y1_LUT4AB/W2BEG[4] Tile_X4Y1_LUT4AB/W2BEG[5] Tile_X4Y1_LUT4AB/W2BEG[6]
+ Tile_X4Y1_LUT4AB/W2BEG[7] Tile_X3Y1_LUT4AB/W2END[0] Tile_X3Y1_LUT4AB/W2END[1] Tile_X3Y1_LUT4AB/W2END[2]
+ Tile_X3Y1_LUT4AB/W2END[3] Tile_X3Y1_LUT4AB/W2END[4] Tile_X3Y1_LUT4AB/W2END[5] Tile_X3Y1_LUT4AB/W2END[6]
+ Tile_X3Y1_LUT4AB/W2END[7] Tile_X4Y1_LUT4AB/W2END[0] Tile_X4Y1_LUT4AB/W2END[1] Tile_X4Y1_LUT4AB/W2END[2]
+ Tile_X4Y1_LUT4AB/W2END[3] Tile_X4Y1_LUT4AB/W2END[4] Tile_X4Y1_LUT4AB/W2END[5] Tile_X4Y1_LUT4AB/W2END[6]
+ Tile_X4Y1_LUT4AB/W2END[7] Tile_X4Y1_LUT4AB/W2MID[0] Tile_X4Y1_LUT4AB/W2MID[1] Tile_X4Y1_LUT4AB/W2MID[2]
+ Tile_X4Y1_LUT4AB/W2MID[3] Tile_X4Y1_LUT4AB/W2MID[4] Tile_X4Y1_LUT4AB/W2MID[5] Tile_X4Y1_LUT4AB/W2MID[6]
+ Tile_X4Y1_LUT4AB/W2MID[7] Tile_X4Y1_LUT4AB/W6BEG[0] Tile_X4Y1_LUT4AB/W6BEG[10] Tile_X4Y1_LUT4AB/W6BEG[11]
+ Tile_X4Y1_LUT4AB/W6BEG[1] Tile_X4Y1_LUT4AB/W6BEG[2] Tile_X4Y1_LUT4AB/W6BEG[3] Tile_X4Y1_LUT4AB/W6BEG[4]
+ Tile_X4Y1_LUT4AB/W6BEG[5] Tile_X4Y1_LUT4AB/W6BEG[6] Tile_X4Y1_LUT4AB/W6BEG[7] Tile_X4Y1_LUT4AB/W6BEG[8]
+ Tile_X4Y1_LUT4AB/W6BEG[9] Tile_X4Y1_LUT4AB/W6END[0] Tile_X4Y1_LUT4AB/W6END[10] Tile_X4Y1_LUT4AB/W6END[11]
+ Tile_X4Y1_LUT4AB/W6END[1] Tile_X4Y1_LUT4AB/W6END[2] Tile_X4Y1_LUT4AB/W6END[3] Tile_X4Y1_LUT4AB/W6END[4]
+ Tile_X4Y1_LUT4AB/W6END[5] Tile_X4Y1_LUT4AB/W6END[6] Tile_X4Y1_LUT4AB/W6END[7] Tile_X4Y1_LUT4AB/W6END[8]
+ Tile_X4Y1_LUT4AB/W6END[9] Tile_X4Y1_LUT4AB/WW4BEG[0] Tile_X4Y1_LUT4AB/WW4BEG[10]
+ Tile_X4Y1_LUT4AB/WW4BEG[11] Tile_X4Y1_LUT4AB/WW4BEG[12] Tile_X4Y1_LUT4AB/WW4BEG[13]
+ Tile_X4Y1_LUT4AB/WW4BEG[14] Tile_X4Y1_LUT4AB/WW4BEG[15] Tile_X4Y1_LUT4AB/WW4BEG[1]
+ Tile_X4Y1_LUT4AB/WW4BEG[2] Tile_X4Y1_LUT4AB/WW4BEG[3] Tile_X4Y1_LUT4AB/WW4BEG[4]
+ Tile_X4Y1_LUT4AB/WW4BEG[5] Tile_X4Y1_LUT4AB/WW4BEG[6] Tile_X4Y1_LUT4AB/WW4BEG[7]
+ Tile_X4Y1_LUT4AB/WW4BEG[8] Tile_X4Y1_LUT4AB/WW4BEG[9] Tile_X4Y1_LUT4AB/WW4END[0]
+ Tile_X4Y1_LUT4AB/WW4END[10] Tile_X4Y1_LUT4AB/WW4END[11] Tile_X4Y1_LUT4AB/WW4END[12]
+ Tile_X4Y1_LUT4AB/WW4END[13] Tile_X4Y1_LUT4AB/WW4END[14] Tile_X4Y1_LUT4AB/WW4END[15]
+ Tile_X4Y1_LUT4AB/WW4END[1] Tile_X4Y1_LUT4AB/WW4END[2] Tile_X4Y1_LUT4AB/WW4END[3]
+ Tile_X4Y1_LUT4AB/WW4END[4] Tile_X4Y1_LUT4AB/WW4END[5] Tile_X4Y1_LUT4AB/WW4END[6]
+ Tile_X4Y1_LUT4AB/WW4END[7] Tile_X4Y1_LUT4AB/WW4END[8] Tile_X4Y1_LUT4AB/WW4END[9]
+ LUT4AB
XTile_X3Y5_LUT4AB Tile_X3Y6_LUT4AB/Co Tile_X3Y5_LUT4AB/Co Tile_X4Y5_LUT4AB/E1END[0]
+ Tile_X4Y5_LUT4AB/E1END[1] Tile_X4Y5_LUT4AB/E1END[2] Tile_X4Y5_LUT4AB/E1END[3] Tile_X3Y5_LUT4AB/E1END[0]
+ Tile_X3Y5_LUT4AB/E1END[1] Tile_X3Y5_LUT4AB/E1END[2] Tile_X3Y5_LUT4AB/E1END[3] Tile_X4Y5_LUT4AB/E2MID[0]
+ Tile_X4Y5_LUT4AB/E2MID[1] Tile_X4Y5_LUT4AB/E2MID[2] Tile_X4Y5_LUT4AB/E2MID[3] Tile_X4Y5_LUT4AB/E2MID[4]
+ Tile_X4Y5_LUT4AB/E2MID[5] Tile_X4Y5_LUT4AB/E2MID[6] Tile_X4Y5_LUT4AB/E2MID[7] Tile_X4Y5_LUT4AB/E2END[0]
+ Tile_X4Y5_LUT4AB/E2END[1] Tile_X4Y5_LUT4AB/E2END[2] Tile_X4Y5_LUT4AB/E2END[3] Tile_X4Y5_LUT4AB/E2END[4]
+ Tile_X4Y5_LUT4AB/E2END[5] Tile_X4Y5_LUT4AB/E2END[6] Tile_X4Y5_LUT4AB/E2END[7] Tile_X3Y5_LUT4AB/E2END[0]
+ Tile_X3Y5_LUT4AB/E2END[1] Tile_X3Y5_LUT4AB/E2END[2] Tile_X3Y5_LUT4AB/E2END[3] Tile_X3Y5_LUT4AB/E2END[4]
+ Tile_X3Y5_LUT4AB/E2END[5] Tile_X3Y5_LUT4AB/E2END[6] Tile_X3Y5_LUT4AB/E2END[7] Tile_X3Y5_LUT4AB/E2MID[0]
+ Tile_X3Y5_LUT4AB/E2MID[1] Tile_X3Y5_LUT4AB/E2MID[2] Tile_X3Y5_LUT4AB/E2MID[3] Tile_X3Y5_LUT4AB/E2MID[4]
+ Tile_X3Y5_LUT4AB/E2MID[5] Tile_X3Y5_LUT4AB/E2MID[6] Tile_X3Y5_LUT4AB/E2MID[7] Tile_X4Y5_LUT4AB/E6END[0]
+ Tile_X4Y5_LUT4AB/E6END[10] Tile_X4Y5_LUT4AB/E6END[11] Tile_X4Y5_LUT4AB/E6END[1]
+ Tile_X4Y5_LUT4AB/E6END[2] Tile_X4Y5_LUT4AB/E6END[3] Tile_X4Y5_LUT4AB/E6END[4] Tile_X4Y5_LUT4AB/E6END[5]
+ Tile_X4Y5_LUT4AB/E6END[6] Tile_X4Y5_LUT4AB/E6END[7] Tile_X4Y5_LUT4AB/E6END[8] Tile_X4Y5_LUT4AB/E6END[9]
+ Tile_X3Y5_LUT4AB/E6END[0] Tile_X3Y5_LUT4AB/E6END[10] Tile_X3Y5_LUT4AB/E6END[11]
+ Tile_X3Y5_LUT4AB/E6END[1] Tile_X3Y5_LUT4AB/E6END[2] Tile_X3Y5_LUT4AB/E6END[3] Tile_X3Y5_LUT4AB/E6END[4]
+ Tile_X3Y5_LUT4AB/E6END[5] Tile_X3Y5_LUT4AB/E6END[6] Tile_X3Y5_LUT4AB/E6END[7] Tile_X3Y5_LUT4AB/E6END[8]
+ Tile_X3Y5_LUT4AB/E6END[9] Tile_X4Y5_LUT4AB/EE4END[0] Tile_X4Y5_LUT4AB/EE4END[10]
+ Tile_X4Y5_LUT4AB/EE4END[11] Tile_X4Y5_LUT4AB/EE4END[12] Tile_X4Y5_LUT4AB/EE4END[13]
+ Tile_X4Y5_LUT4AB/EE4END[14] Tile_X4Y5_LUT4AB/EE4END[15] Tile_X4Y5_LUT4AB/EE4END[1]
+ Tile_X4Y5_LUT4AB/EE4END[2] Tile_X4Y5_LUT4AB/EE4END[3] Tile_X4Y5_LUT4AB/EE4END[4]
+ Tile_X4Y5_LUT4AB/EE4END[5] Tile_X4Y5_LUT4AB/EE4END[6] Tile_X4Y5_LUT4AB/EE4END[7]
+ Tile_X4Y5_LUT4AB/EE4END[8] Tile_X4Y5_LUT4AB/EE4END[9] Tile_X3Y5_LUT4AB/EE4END[0]
+ Tile_X3Y5_LUT4AB/EE4END[10] Tile_X3Y5_LUT4AB/EE4END[11] Tile_X3Y5_LUT4AB/EE4END[12]
+ Tile_X3Y5_LUT4AB/EE4END[13] Tile_X3Y5_LUT4AB/EE4END[14] Tile_X3Y5_LUT4AB/EE4END[15]
+ Tile_X3Y5_LUT4AB/EE4END[1] Tile_X3Y5_LUT4AB/EE4END[2] Tile_X3Y5_LUT4AB/EE4END[3]
+ Tile_X3Y5_LUT4AB/EE4END[4] Tile_X3Y5_LUT4AB/EE4END[5] Tile_X3Y5_LUT4AB/EE4END[6]
+ Tile_X3Y5_LUT4AB/EE4END[7] Tile_X3Y5_LUT4AB/EE4END[8] Tile_X3Y5_LUT4AB/EE4END[9]
+ Tile_X3Y5_LUT4AB/FrameData[0] Tile_X3Y5_LUT4AB/FrameData[10] Tile_X3Y5_LUT4AB/FrameData[11]
+ Tile_X3Y5_LUT4AB/FrameData[12] Tile_X3Y5_LUT4AB/FrameData[13] Tile_X3Y5_LUT4AB/FrameData[14]
+ Tile_X3Y5_LUT4AB/FrameData[15] Tile_X3Y5_LUT4AB/FrameData[16] Tile_X3Y5_LUT4AB/FrameData[17]
+ Tile_X3Y5_LUT4AB/FrameData[18] Tile_X3Y5_LUT4AB/FrameData[19] Tile_X3Y5_LUT4AB/FrameData[1]
+ Tile_X3Y5_LUT4AB/FrameData[20] Tile_X3Y5_LUT4AB/FrameData[21] Tile_X3Y5_LUT4AB/FrameData[22]
+ Tile_X3Y5_LUT4AB/FrameData[23] Tile_X3Y5_LUT4AB/FrameData[24] Tile_X3Y5_LUT4AB/FrameData[25]
+ Tile_X3Y5_LUT4AB/FrameData[26] Tile_X3Y5_LUT4AB/FrameData[27] Tile_X3Y5_LUT4AB/FrameData[28]
+ Tile_X3Y5_LUT4AB/FrameData[29] Tile_X3Y5_LUT4AB/FrameData[2] Tile_X3Y5_LUT4AB/FrameData[30]
+ Tile_X3Y5_LUT4AB/FrameData[31] Tile_X3Y5_LUT4AB/FrameData[3] Tile_X3Y5_LUT4AB/FrameData[4]
+ Tile_X3Y5_LUT4AB/FrameData[5] Tile_X3Y5_LUT4AB/FrameData[6] Tile_X3Y5_LUT4AB/FrameData[7]
+ Tile_X3Y5_LUT4AB/FrameData[8] Tile_X3Y5_LUT4AB/FrameData[9] Tile_X4Y5_LUT4AB/FrameData[0]
+ Tile_X4Y5_LUT4AB/FrameData[10] Tile_X4Y5_LUT4AB/FrameData[11] Tile_X4Y5_LUT4AB/FrameData[12]
+ Tile_X4Y5_LUT4AB/FrameData[13] Tile_X4Y5_LUT4AB/FrameData[14] Tile_X4Y5_LUT4AB/FrameData[15]
+ Tile_X4Y5_LUT4AB/FrameData[16] Tile_X4Y5_LUT4AB/FrameData[17] Tile_X4Y5_LUT4AB/FrameData[18]
+ Tile_X4Y5_LUT4AB/FrameData[19] Tile_X4Y5_LUT4AB/FrameData[1] Tile_X4Y5_LUT4AB/FrameData[20]
+ Tile_X4Y5_LUT4AB/FrameData[21] Tile_X4Y5_LUT4AB/FrameData[22] Tile_X4Y5_LUT4AB/FrameData[23]
+ Tile_X4Y5_LUT4AB/FrameData[24] Tile_X4Y5_LUT4AB/FrameData[25] Tile_X4Y5_LUT4AB/FrameData[26]
+ Tile_X4Y5_LUT4AB/FrameData[27] Tile_X4Y5_LUT4AB/FrameData[28] Tile_X4Y5_LUT4AB/FrameData[29]
+ Tile_X4Y5_LUT4AB/FrameData[2] Tile_X4Y5_LUT4AB/FrameData[30] Tile_X4Y5_LUT4AB/FrameData[31]
+ Tile_X4Y5_LUT4AB/FrameData[3] Tile_X4Y5_LUT4AB/FrameData[4] Tile_X4Y5_LUT4AB/FrameData[5]
+ Tile_X4Y5_LUT4AB/FrameData[6] Tile_X4Y5_LUT4AB/FrameData[7] Tile_X4Y5_LUT4AB/FrameData[8]
+ Tile_X4Y5_LUT4AB/FrameData[9] Tile_X3Y5_LUT4AB/FrameStrobe[0] Tile_X3Y5_LUT4AB/FrameStrobe[10]
+ Tile_X3Y5_LUT4AB/FrameStrobe[11] Tile_X3Y5_LUT4AB/FrameStrobe[12] Tile_X3Y5_LUT4AB/FrameStrobe[13]
+ Tile_X3Y5_LUT4AB/FrameStrobe[14] Tile_X3Y5_LUT4AB/FrameStrobe[15] Tile_X3Y5_LUT4AB/FrameStrobe[16]
+ Tile_X3Y5_LUT4AB/FrameStrobe[17] Tile_X3Y5_LUT4AB/FrameStrobe[18] Tile_X3Y5_LUT4AB/FrameStrobe[19]
+ Tile_X3Y5_LUT4AB/FrameStrobe[1] Tile_X3Y5_LUT4AB/FrameStrobe[2] Tile_X3Y5_LUT4AB/FrameStrobe[3]
+ Tile_X3Y5_LUT4AB/FrameStrobe[4] Tile_X3Y5_LUT4AB/FrameStrobe[5] Tile_X3Y5_LUT4AB/FrameStrobe[6]
+ Tile_X3Y5_LUT4AB/FrameStrobe[7] Tile_X3Y5_LUT4AB/FrameStrobe[8] Tile_X3Y5_LUT4AB/FrameStrobe[9]
+ Tile_X3Y4_LUT4AB/FrameStrobe[0] Tile_X3Y4_LUT4AB/FrameStrobe[10] Tile_X3Y4_LUT4AB/FrameStrobe[11]
+ Tile_X3Y4_LUT4AB/FrameStrobe[12] Tile_X3Y4_LUT4AB/FrameStrobe[13] Tile_X3Y4_LUT4AB/FrameStrobe[14]
+ Tile_X3Y4_LUT4AB/FrameStrobe[15] Tile_X3Y4_LUT4AB/FrameStrobe[16] Tile_X3Y4_LUT4AB/FrameStrobe[17]
+ Tile_X3Y4_LUT4AB/FrameStrobe[18] Tile_X3Y4_LUT4AB/FrameStrobe[19] Tile_X3Y4_LUT4AB/FrameStrobe[1]
+ Tile_X3Y4_LUT4AB/FrameStrobe[2] Tile_X3Y4_LUT4AB/FrameStrobe[3] Tile_X3Y4_LUT4AB/FrameStrobe[4]
+ Tile_X3Y4_LUT4AB/FrameStrobe[5] Tile_X3Y4_LUT4AB/FrameStrobe[6] Tile_X3Y4_LUT4AB/FrameStrobe[7]
+ Tile_X3Y4_LUT4AB/FrameStrobe[8] Tile_X3Y4_LUT4AB/FrameStrobe[9] Tile_X3Y5_LUT4AB/N1BEG[0]
+ Tile_X3Y5_LUT4AB/N1BEG[1] Tile_X3Y5_LUT4AB/N1BEG[2] Tile_X3Y5_LUT4AB/N1BEG[3] Tile_X3Y6_LUT4AB/N1BEG[0]
+ Tile_X3Y6_LUT4AB/N1BEG[1] Tile_X3Y6_LUT4AB/N1BEG[2] Tile_X3Y6_LUT4AB/N1BEG[3] Tile_X3Y5_LUT4AB/N2BEG[0]
+ Tile_X3Y5_LUT4AB/N2BEG[1] Tile_X3Y5_LUT4AB/N2BEG[2] Tile_X3Y5_LUT4AB/N2BEG[3] Tile_X3Y5_LUT4AB/N2BEG[4]
+ Tile_X3Y5_LUT4AB/N2BEG[5] Tile_X3Y5_LUT4AB/N2BEG[6] Tile_X3Y5_LUT4AB/N2BEG[7] Tile_X3Y4_LUT4AB/N2END[0]
+ Tile_X3Y4_LUT4AB/N2END[1] Tile_X3Y4_LUT4AB/N2END[2] Tile_X3Y4_LUT4AB/N2END[3] Tile_X3Y4_LUT4AB/N2END[4]
+ Tile_X3Y4_LUT4AB/N2END[5] Tile_X3Y4_LUT4AB/N2END[6] Tile_X3Y4_LUT4AB/N2END[7] Tile_X3Y5_LUT4AB/N2END[0]
+ Tile_X3Y5_LUT4AB/N2END[1] Tile_X3Y5_LUT4AB/N2END[2] Tile_X3Y5_LUT4AB/N2END[3] Tile_X3Y5_LUT4AB/N2END[4]
+ Tile_X3Y5_LUT4AB/N2END[5] Tile_X3Y5_LUT4AB/N2END[6] Tile_X3Y5_LUT4AB/N2END[7] Tile_X3Y6_LUT4AB/N2BEG[0]
+ Tile_X3Y6_LUT4AB/N2BEG[1] Tile_X3Y6_LUT4AB/N2BEG[2] Tile_X3Y6_LUT4AB/N2BEG[3] Tile_X3Y6_LUT4AB/N2BEG[4]
+ Tile_X3Y6_LUT4AB/N2BEG[5] Tile_X3Y6_LUT4AB/N2BEG[6] Tile_X3Y6_LUT4AB/N2BEG[7] Tile_X3Y5_LUT4AB/N4BEG[0]
+ Tile_X3Y5_LUT4AB/N4BEG[10] Tile_X3Y5_LUT4AB/N4BEG[11] Tile_X3Y5_LUT4AB/N4BEG[12]
+ Tile_X3Y5_LUT4AB/N4BEG[13] Tile_X3Y5_LUT4AB/N4BEG[14] Tile_X3Y5_LUT4AB/N4BEG[15]
+ Tile_X3Y5_LUT4AB/N4BEG[1] Tile_X3Y5_LUT4AB/N4BEG[2] Tile_X3Y5_LUT4AB/N4BEG[3] Tile_X3Y5_LUT4AB/N4BEG[4]
+ Tile_X3Y5_LUT4AB/N4BEG[5] Tile_X3Y5_LUT4AB/N4BEG[6] Tile_X3Y5_LUT4AB/N4BEG[7] Tile_X3Y5_LUT4AB/N4BEG[8]
+ Tile_X3Y5_LUT4AB/N4BEG[9] Tile_X3Y6_LUT4AB/N4BEG[0] Tile_X3Y6_LUT4AB/N4BEG[10] Tile_X3Y6_LUT4AB/N4BEG[11]
+ Tile_X3Y6_LUT4AB/N4BEG[12] Tile_X3Y6_LUT4AB/N4BEG[13] Tile_X3Y6_LUT4AB/N4BEG[14]
+ Tile_X3Y6_LUT4AB/N4BEG[15] Tile_X3Y6_LUT4AB/N4BEG[1] Tile_X3Y6_LUT4AB/N4BEG[2] Tile_X3Y6_LUT4AB/N4BEG[3]
+ Tile_X3Y6_LUT4AB/N4BEG[4] Tile_X3Y6_LUT4AB/N4BEG[5] Tile_X3Y6_LUT4AB/N4BEG[6] Tile_X3Y6_LUT4AB/N4BEG[7]
+ Tile_X3Y6_LUT4AB/N4BEG[8] Tile_X3Y6_LUT4AB/N4BEG[9] Tile_X3Y5_LUT4AB/NN4BEG[0] Tile_X3Y5_LUT4AB/NN4BEG[10]
+ Tile_X3Y5_LUT4AB/NN4BEG[11] Tile_X3Y5_LUT4AB/NN4BEG[12] Tile_X3Y5_LUT4AB/NN4BEG[13]
+ Tile_X3Y5_LUT4AB/NN4BEG[14] Tile_X3Y5_LUT4AB/NN4BEG[15] Tile_X3Y5_LUT4AB/NN4BEG[1]
+ Tile_X3Y5_LUT4AB/NN4BEG[2] Tile_X3Y5_LUT4AB/NN4BEG[3] Tile_X3Y5_LUT4AB/NN4BEG[4]
+ Tile_X3Y5_LUT4AB/NN4BEG[5] Tile_X3Y5_LUT4AB/NN4BEG[6] Tile_X3Y5_LUT4AB/NN4BEG[7]
+ Tile_X3Y5_LUT4AB/NN4BEG[8] Tile_X3Y5_LUT4AB/NN4BEG[9] Tile_X3Y6_LUT4AB/NN4BEG[0]
+ Tile_X3Y6_LUT4AB/NN4BEG[10] Tile_X3Y6_LUT4AB/NN4BEG[11] Tile_X3Y6_LUT4AB/NN4BEG[12]
+ Tile_X3Y6_LUT4AB/NN4BEG[13] Tile_X3Y6_LUT4AB/NN4BEG[14] Tile_X3Y6_LUT4AB/NN4BEG[15]
+ Tile_X3Y6_LUT4AB/NN4BEG[1] Tile_X3Y6_LUT4AB/NN4BEG[2] Tile_X3Y6_LUT4AB/NN4BEG[3]
+ Tile_X3Y6_LUT4AB/NN4BEG[4] Tile_X3Y6_LUT4AB/NN4BEG[5] Tile_X3Y6_LUT4AB/NN4BEG[6]
+ Tile_X3Y6_LUT4AB/NN4BEG[7] Tile_X3Y6_LUT4AB/NN4BEG[8] Tile_X3Y6_LUT4AB/NN4BEG[9]
+ Tile_X3Y6_LUT4AB/S1END[0] Tile_X3Y6_LUT4AB/S1END[1] Tile_X3Y6_LUT4AB/S1END[2] Tile_X3Y6_LUT4AB/S1END[3]
+ Tile_X3Y5_LUT4AB/S1END[0] Tile_X3Y5_LUT4AB/S1END[1] Tile_X3Y5_LUT4AB/S1END[2] Tile_X3Y5_LUT4AB/S1END[3]
+ Tile_X3Y6_LUT4AB/S2MID[0] Tile_X3Y6_LUT4AB/S2MID[1] Tile_X3Y6_LUT4AB/S2MID[2] Tile_X3Y6_LUT4AB/S2MID[3]
+ Tile_X3Y6_LUT4AB/S2MID[4] Tile_X3Y6_LUT4AB/S2MID[5] Tile_X3Y6_LUT4AB/S2MID[6] Tile_X3Y6_LUT4AB/S2MID[7]
+ Tile_X3Y6_LUT4AB/S2END[0] Tile_X3Y6_LUT4AB/S2END[1] Tile_X3Y6_LUT4AB/S2END[2] Tile_X3Y6_LUT4AB/S2END[3]
+ Tile_X3Y6_LUT4AB/S2END[4] Tile_X3Y6_LUT4AB/S2END[5] Tile_X3Y6_LUT4AB/S2END[6] Tile_X3Y6_LUT4AB/S2END[7]
+ Tile_X3Y5_LUT4AB/S2END[0] Tile_X3Y5_LUT4AB/S2END[1] Tile_X3Y5_LUT4AB/S2END[2] Tile_X3Y5_LUT4AB/S2END[3]
+ Tile_X3Y5_LUT4AB/S2END[4] Tile_X3Y5_LUT4AB/S2END[5] Tile_X3Y5_LUT4AB/S2END[6] Tile_X3Y5_LUT4AB/S2END[7]
+ Tile_X3Y5_LUT4AB/S2MID[0] Tile_X3Y5_LUT4AB/S2MID[1] Tile_X3Y5_LUT4AB/S2MID[2] Tile_X3Y5_LUT4AB/S2MID[3]
+ Tile_X3Y5_LUT4AB/S2MID[4] Tile_X3Y5_LUT4AB/S2MID[5] Tile_X3Y5_LUT4AB/S2MID[6] Tile_X3Y5_LUT4AB/S2MID[7]
+ Tile_X3Y6_LUT4AB/S4END[0] Tile_X3Y6_LUT4AB/S4END[10] Tile_X3Y6_LUT4AB/S4END[11]
+ Tile_X3Y6_LUT4AB/S4END[12] Tile_X3Y6_LUT4AB/S4END[13] Tile_X3Y6_LUT4AB/S4END[14]
+ Tile_X3Y6_LUT4AB/S4END[15] Tile_X3Y6_LUT4AB/S4END[1] Tile_X3Y6_LUT4AB/S4END[2] Tile_X3Y6_LUT4AB/S4END[3]
+ Tile_X3Y6_LUT4AB/S4END[4] Tile_X3Y6_LUT4AB/S4END[5] Tile_X3Y6_LUT4AB/S4END[6] Tile_X3Y6_LUT4AB/S4END[7]
+ Tile_X3Y6_LUT4AB/S4END[8] Tile_X3Y6_LUT4AB/S4END[9] Tile_X3Y5_LUT4AB/S4END[0] Tile_X3Y5_LUT4AB/S4END[10]
+ Tile_X3Y5_LUT4AB/S4END[11] Tile_X3Y5_LUT4AB/S4END[12] Tile_X3Y5_LUT4AB/S4END[13]
+ Tile_X3Y5_LUT4AB/S4END[14] Tile_X3Y5_LUT4AB/S4END[15] Tile_X3Y5_LUT4AB/S4END[1]
+ Tile_X3Y5_LUT4AB/S4END[2] Tile_X3Y5_LUT4AB/S4END[3] Tile_X3Y5_LUT4AB/S4END[4] Tile_X3Y5_LUT4AB/S4END[5]
+ Tile_X3Y5_LUT4AB/S4END[6] Tile_X3Y5_LUT4AB/S4END[7] Tile_X3Y5_LUT4AB/S4END[8] Tile_X3Y5_LUT4AB/S4END[9]
+ Tile_X3Y6_LUT4AB/SS4END[0] Tile_X3Y6_LUT4AB/SS4END[10] Tile_X3Y6_LUT4AB/SS4END[11]
+ Tile_X3Y6_LUT4AB/SS4END[12] Tile_X3Y6_LUT4AB/SS4END[13] Tile_X3Y6_LUT4AB/SS4END[14]
+ Tile_X3Y6_LUT4AB/SS4END[15] Tile_X3Y6_LUT4AB/SS4END[1] Tile_X3Y6_LUT4AB/SS4END[2]
+ Tile_X3Y6_LUT4AB/SS4END[3] Tile_X3Y6_LUT4AB/SS4END[4] Tile_X3Y6_LUT4AB/SS4END[5]
+ Tile_X3Y6_LUT4AB/SS4END[6] Tile_X3Y6_LUT4AB/SS4END[7] Tile_X3Y6_LUT4AB/SS4END[8]
+ Tile_X3Y6_LUT4AB/SS4END[9] Tile_X3Y5_LUT4AB/SS4END[0] Tile_X3Y5_LUT4AB/SS4END[10]
+ Tile_X3Y5_LUT4AB/SS4END[11] Tile_X3Y5_LUT4AB/SS4END[12] Tile_X3Y5_LUT4AB/SS4END[13]
+ Tile_X3Y5_LUT4AB/SS4END[14] Tile_X3Y5_LUT4AB/SS4END[15] Tile_X3Y5_LUT4AB/SS4END[1]
+ Tile_X3Y5_LUT4AB/SS4END[2] Tile_X3Y5_LUT4AB/SS4END[3] Tile_X3Y5_LUT4AB/SS4END[4]
+ Tile_X3Y5_LUT4AB/SS4END[5] Tile_X3Y5_LUT4AB/SS4END[6] Tile_X3Y5_LUT4AB/SS4END[7]
+ Tile_X3Y5_LUT4AB/SS4END[8] Tile_X3Y5_LUT4AB/SS4END[9] Tile_X3Y5_LUT4AB/UserCLK Tile_X3Y4_LUT4AB/UserCLK
+ VGND VPWR Tile_X3Y5_LUT4AB/W1BEG[0] Tile_X3Y5_LUT4AB/W1BEG[1] Tile_X3Y5_LUT4AB/W1BEG[2]
+ Tile_X3Y5_LUT4AB/W1BEG[3] Tile_X4Y5_LUT4AB/W1BEG[0] Tile_X4Y5_LUT4AB/W1BEG[1] Tile_X4Y5_LUT4AB/W1BEG[2]
+ Tile_X4Y5_LUT4AB/W1BEG[3] Tile_X3Y5_LUT4AB/W2BEG[0] Tile_X3Y5_LUT4AB/W2BEG[1] Tile_X3Y5_LUT4AB/W2BEG[2]
+ Tile_X3Y5_LUT4AB/W2BEG[3] Tile_X3Y5_LUT4AB/W2BEG[4] Tile_X3Y5_LUT4AB/W2BEG[5] Tile_X3Y5_LUT4AB/W2BEG[6]
+ Tile_X3Y5_LUT4AB/W2BEG[7] Tile_X2Y5_LUT4AB/W2END[0] Tile_X2Y5_LUT4AB/W2END[1] Tile_X2Y5_LUT4AB/W2END[2]
+ Tile_X2Y5_LUT4AB/W2END[3] Tile_X2Y5_LUT4AB/W2END[4] Tile_X2Y5_LUT4AB/W2END[5] Tile_X2Y5_LUT4AB/W2END[6]
+ Tile_X2Y5_LUT4AB/W2END[7] Tile_X3Y5_LUT4AB/W2END[0] Tile_X3Y5_LUT4AB/W2END[1] Tile_X3Y5_LUT4AB/W2END[2]
+ Tile_X3Y5_LUT4AB/W2END[3] Tile_X3Y5_LUT4AB/W2END[4] Tile_X3Y5_LUT4AB/W2END[5] Tile_X3Y5_LUT4AB/W2END[6]
+ Tile_X3Y5_LUT4AB/W2END[7] Tile_X4Y5_LUT4AB/W2BEG[0] Tile_X4Y5_LUT4AB/W2BEG[1] Tile_X4Y5_LUT4AB/W2BEG[2]
+ Tile_X4Y5_LUT4AB/W2BEG[3] Tile_X4Y5_LUT4AB/W2BEG[4] Tile_X4Y5_LUT4AB/W2BEG[5] Tile_X4Y5_LUT4AB/W2BEG[6]
+ Tile_X4Y5_LUT4AB/W2BEG[7] Tile_X3Y5_LUT4AB/W6BEG[0] Tile_X3Y5_LUT4AB/W6BEG[10] Tile_X3Y5_LUT4AB/W6BEG[11]
+ Tile_X3Y5_LUT4AB/W6BEG[1] Tile_X3Y5_LUT4AB/W6BEG[2] Tile_X3Y5_LUT4AB/W6BEG[3] Tile_X3Y5_LUT4AB/W6BEG[4]
+ Tile_X3Y5_LUT4AB/W6BEG[5] Tile_X3Y5_LUT4AB/W6BEG[6] Tile_X3Y5_LUT4AB/W6BEG[7] Tile_X3Y5_LUT4AB/W6BEG[8]
+ Tile_X3Y5_LUT4AB/W6BEG[9] Tile_X4Y5_LUT4AB/W6BEG[0] Tile_X4Y5_LUT4AB/W6BEG[10] Tile_X4Y5_LUT4AB/W6BEG[11]
+ Tile_X4Y5_LUT4AB/W6BEG[1] Tile_X4Y5_LUT4AB/W6BEG[2] Tile_X4Y5_LUT4AB/W6BEG[3] Tile_X4Y5_LUT4AB/W6BEG[4]
+ Tile_X4Y5_LUT4AB/W6BEG[5] Tile_X4Y5_LUT4AB/W6BEG[6] Tile_X4Y5_LUT4AB/W6BEG[7] Tile_X4Y5_LUT4AB/W6BEG[8]
+ Tile_X4Y5_LUT4AB/W6BEG[9] Tile_X3Y5_LUT4AB/WW4BEG[0] Tile_X3Y5_LUT4AB/WW4BEG[10]
+ Tile_X3Y5_LUT4AB/WW4BEG[11] Tile_X3Y5_LUT4AB/WW4BEG[12] Tile_X3Y5_LUT4AB/WW4BEG[13]
+ Tile_X3Y5_LUT4AB/WW4BEG[14] Tile_X3Y5_LUT4AB/WW4BEG[15] Tile_X3Y5_LUT4AB/WW4BEG[1]
+ Tile_X3Y5_LUT4AB/WW4BEG[2] Tile_X3Y5_LUT4AB/WW4BEG[3] Tile_X3Y5_LUT4AB/WW4BEG[4]
+ Tile_X3Y5_LUT4AB/WW4BEG[5] Tile_X3Y5_LUT4AB/WW4BEG[6] Tile_X3Y5_LUT4AB/WW4BEG[7]
+ Tile_X3Y5_LUT4AB/WW4BEG[8] Tile_X3Y5_LUT4AB/WW4BEG[9] Tile_X4Y5_LUT4AB/WW4BEG[0]
+ Tile_X4Y5_LUT4AB/WW4BEG[10] Tile_X4Y5_LUT4AB/WW4BEG[11] Tile_X4Y5_LUT4AB/WW4BEG[12]
+ Tile_X4Y5_LUT4AB/WW4BEG[13] Tile_X4Y5_LUT4AB/WW4BEG[14] Tile_X4Y5_LUT4AB/WW4BEG[15]
+ Tile_X4Y5_LUT4AB/WW4BEG[1] Tile_X4Y5_LUT4AB/WW4BEG[2] Tile_X4Y5_LUT4AB/WW4BEG[3]
+ Tile_X4Y5_LUT4AB/WW4BEG[4] Tile_X4Y5_LUT4AB/WW4BEG[5] Tile_X4Y5_LUT4AB/WW4BEG[6]
+ Tile_X4Y5_LUT4AB/WW4BEG[7] Tile_X4Y5_LUT4AB/WW4BEG[8] Tile_X4Y5_LUT4AB/WW4BEG[9]
+ LUT4AB
XTile_X2Y9_S_IO4 Tile_X2Y9_A_I_top Tile_X2Y9_A_O_top Tile_X2Y9_A_T_top Tile_X2Y9_B_I_top
+ Tile_X2Y9_B_O_top Tile_X2Y9_B_T_top Tile_X2Y9_C_I_top Tile_X2Y9_C_O_top Tile_X2Y9_C_T_top
+ Tile_X2Y9_S_IO4/Co Tile_X2Y9_D_I_top Tile_X2Y9_D_O_top Tile_X2Y9_D_T_top Tile_X2Y9_S_IO4/FrameData[0]
+ Tile_X2Y9_S_IO4/FrameData[10] Tile_X2Y9_S_IO4/FrameData[11] Tile_X2Y9_S_IO4/FrameData[12]
+ Tile_X2Y9_S_IO4/FrameData[13] Tile_X2Y9_S_IO4/FrameData[14] Tile_X2Y9_S_IO4/FrameData[15]
+ Tile_X2Y9_S_IO4/FrameData[16] Tile_X2Y9_S_IO4/FrameData[17] Tile_X2Y9_S_IO4/FrameData[18]
+ Tile_X2Y9_S_IO4/FrameData[19] Tile_X2Y9_S_IO4/FrameData[1] Tile_X2Y9_S_IO4/FrameData[20]
+ Tile_X2Y9_S_IO4/FrameData[21] Tile_X2Y9_S_IO4/FrameData[22] Tile_X2Y9_S_IO4/FrameData[23]
+ Tile_X2Y9_S_IO4/FrameData[24] Tile_X2Y9_S_IO4/FrameData[25] Tile_X2Y9_S_IO4/FrameData[26]
+ Tile_X2Y9_S_IO4/FrameData[27] Tile_X2Y9_S_IO4/FrameData[28] Tile_X2Y9_S_IO4/FrameData[29]
+ Tile_X2Y9_S_IO4/FrameData[2] Tile_X2Y9_S_IO4/FrameData[30] Tile_X2Y9_S_IO4/FrameData[31]
+ Tile_X2Y9_S_IO4/FrameData[3] Tile_X2Y9_S_IO4/FrameData[4] Tile_X2Y9_S_IO4/FrameData[5]
+ Tile_X2Y9_S_IO4/FrameData[6] Tile_X2Y9_S_IO4/FrameData[7] Tile_X2Y9_S_IO4/FrameData[8]
+ Tile_X2Y9_S_IO4/FrameData[9] Tile_X3Y9_S_IO4/FrameData[0] Tile_X3Y9_S_IO4/FrameData[10]
+ Tile_X3Y9_S_IO4/FrameData[11] Tile_X3Y9_S_IO4/FrameData[12] Tile_X3Y9_S_IO4/FrameData[13]
+ Tile_X3Y9_S_IO4/FrameData[14] Tile_X3Y9_S_IO4/FrameData[15] Tile_X3Y9_S_IO4/FrameData[16]
+ Tile_X3Y9_S_IO4/FrameData[17] Tile_X3Y9_S_IO4/FrameData[18] Tile_X3Y9_S_IO4/FrameData[19]
+ Tile_X3Y9_S_IO4/FrameData[1] Tile_X3Y9_S_IO4/FrameData[20] Tile_X3Y9_S_IO4/FrameData[21]
+ Tile_X3Y9_S_IO4/FrameData[22] Tile_X3Y9_S_IO4/FrameData[23] Tile_X3Y9_S_IO4/FrameData[24]
+ Tile_X3Y9_S_IO4/FrameData[25] Tile_X3Y9_S_IO4/FrameData[26] Tile_X3Y9_S_IO4/FrameData[27]
+ Tile_X3Y9_S_IO4/FrameData[28] Tile_X3Y9_S_IO4/FrameData[29] Tile_X3Y9_S_IO4/FrameData[2]
+ Tile_X3Y9_S_IO4/FrameData[30] Tile_X3Y9_S_IO4/FrameData[31] Tile_X3Y9_S_IO4/FrameData[3]
+ Tile_X3Y9_S_IO4/FrameData[4] Tile_X3Y9_S_IO4/FrameData[5] Tile_X3Y9_S_IO4/FrameData[6]
+ Tile_X3Y9_S_IO4/FrameData[7] Tile_X3Y9_S_IO4/FrameData[8] Tile_X3Y9_S_IO4/FrameData[9]
+ FrameStrobe[40] FrameStrobe[50] FrameStrobe[51] FrameStrobe[52] FrameStrobe[53]
+ FrameStrobe[54] FrameStrobe[55] FrameStrobe[56] FrameStrobe[57] FrameStrobe[58]
+ FrameStrobe[59] FrameStrobe[41] FrameStrobe[42] FrameStrobe[43] FrameStrobe[44]
+ FrameStrobe[45] FrameStrobe[46] FrameStrobe[47] FrameStrobe[48] FrameStrobe[49]
+ Tile_X2Y8_LUT4AB/FrameStrobe[0] Tile_X2Y8_LUT4AB/FrameStrobe[10] Tile_X2Y8_LUT4AB/FrameStrobe[11]
+ Tile_X2Y8_LUT4AB/FrameStrobe[12] Tile_X2Y8_LUT4AB/FrameStrobe[13] Tile_X2Y8_LUT4AB/FrameStrobe[14]
+ Tile_X2Y8_LUT4AB/FrameStrobe[15] Tile_X2Y8_LUT4AB/FrameStrobe[16] Tile_X2Y8_LUT4AB/FrameStrobe[17]
+ Tile_X2Y8_LUT4AB/FrameStrobe[18] Tile_X2Y8_LUT4AB/FrameStrobe[19] Tile_X2Y8_LUT4AB/FrameStrobe[1]
+ Tile_X2Y8_LUT4AB/FrameStrobe[2] Tile_X2Y8_LUT4AB/FrameStrobe[3] Tile_X2Y8_LUT4AB/FrameStrobe[4]
+ Tile_X2Y8_LUT4AB/FrameStrobe[5] Tile_X2Y8_LUT4AB/FrameStrobe[6] Tile_X2Y8_LUT4AB/FrameStrobe[7]
+ Tile_X2Y8_LUT4AB/FrameStrobe[8] Tile_X2Y8_LUT4AB/FrameStrobe[9] Tile_X2Y9_S_IO4/N1BEG[0]
+ Tile_X2Y9_S_IO4/N1BEG[1] Tile_X2Y9_S_IO4/N1BEG[2] Tile_X2Y9_S_IO4/N1BEG[3] Tile_X2Y9_S_IO4/N2BEG[0]
+ Tile_X2Y9_S_IO4/N2BEG[1] Tile_X2Y9_S_IO4/N2BEG[2] Tile_X2Y9_S_IO4/N2BEG[3] Tile_X2Y9_S_IO4/N2BEG[4]
+ Tile_X2Y9_S_IO4/N2BEG[5] Tile_X2Y9_S_IO4/N2BEG[6] Tile_X2Y9_S_IO4/N2BEG[7] Tile_X2Y9_S_IO4/N2BEGb[0]
+ Tile_X2Y9_S_IO4/N2BEGb[1] Tile_X2Y9_S_IO4/N2BEGb[2] Tile_X2Y9_S_IO4/N2BEGb[3] Tile_X2Y9_S_IO4/N2BEGb[4]
+ Tile_X2Y9_S_IO4/N2BEGb[5] Tile_X2Y9_S_IO4/N2BEGb[6] Tile_X2Y9_S_IO4/N2BEGb[7] Tile_X2Y9_S_IO4/N4BEG[0]
+ Tile_X2Y9_S_IO4/N4BEG[10] Tile_X2Y9_S_IO4/N4BEG[11] Tile_X2Y9_S_IO4/N4BEG[12] Tile_X2Y9_S_IO4/N4BEG[13]
+ Tile_X2Y9_S_IO4/N4BEG[14] Tile_X2Y9_S_IO4/N4BEG[15] Tile_X2Y9_S_IO4/N4BEG[1] Tile_X2Y9_S_IO4/N4BEG[2]
+ Tile_X2Y9_S_IO4/N4BEG[3] Tile_X2Y9_S_IO4/N4BEG[4] Tile_X2Y9_S_IO4/N4BEG[5] Tile_X2Y9_S_IO4/N4BEG[6]
+ Tile_X2Y9_S_IO4/N4BEG[7] Tile_X2Y9_S_IO4/N4BEG[8] Tile_X2Y9_S_IO4/N4BEG[9] Tile_X2Y9_S_IO4/NN4BEG[0]
+ Tile_X2Y9_S_IO4/NN4BEG[10] Tile_X2Y9_S_IO4/NN4BEG[11] Tile_X2Y9_S_IO4/NN4BEG[12]
+ Tile_X2Y9_S_IO4/NN4BEG[13] Tile_X2Y9_S_IO4/NN4BEG[14] Tile_X2Y9_S_IO4/NN4BEG[15]
+ Tile_X2Y9_S_IO4/NN4BEG[1] Tile_X2Y9_S_IO4/NN4BEG[2] Tile_X2Y9_S_IO4/NN4BEG[3] Tile_X2Y9_S_IO4/NN4BEG[4]
+ Tile_X2Y9_S_IO4/NN4BEG[5] Tile_X2Y9_S_IO4/NN4BEG[6] Tile_X2Y9_S_IO4/NN4BEG[7] Tile_X2Y9_S_IO4/NN4BEG[8]
+ Tile_X2Y9_S_IO4/NN4BEG[9] Tile_X2Y9_S_IO4/S1END[0] Tile_X2Y9_S_IO4/S1END[1] Tile_X2Y9_S_IO4/S1END[2]
+ Tile_X2Y9_S_IO4/S1END[3] Tile_X2Y9_S_IO4/S2END[0] Tile_X2Y9_S_IO4/S2END[1] Tile_X2Y9_S_IO4/S2END[2]
+ Tile_X2Y9_S_IO4/S2END[3] Tile_X2Y9_S_IO4/S2END[4] Tile_X2Y9_S_IO4/S2END[5] Tile_X2Y9_S_IO4/S2END[6]
+ Tile_X2Y9_S_IO4/S2END[7] Tile_X2Y9_S_IO4/S2MID[0] Tile_X2Y9_S_IO4/S2MID[1] Tile_X2Y9_S_IO4/S2MID[2]
+ Tile_X2Y9_S_IO4/S2MID[3] Tile_X2Y9_S_IO4/S2MID[4] Tile_X2Y9_S_IO4/S2MID[5] Tile_X2Y9_S_IO4/S2MID[6]
+ Tile_X2Y9_S_IO4/S2MID[7] Tile_X2Y9_S_IO4/S4END[0] Tile_X2Y9_S_IO4/S4END[10] Tile_X2Y9_S_IO4/S4END[11]
+ Tile_X2Y9_S_IO4/S4END[12] Tile_X2Y9_S_IO4/S4END[13] Tile_X2Y9_S_IO4/S4END[14] Tile_X2Y9_S_IO4/S4END[15]
+ Tile_X2Y9_S_IO4/S4END[1] Tile_X2Y9_S_IO4/S4END[2] Tile_X2Y9_S_IO4/S4END[3] Tile_X2Y9_S_IO4/S4END[4]
+ Tile_X2Y9_S_IO4/S4END[5] Tile_X2Y9_S_IO4/S4END[6] Tile_X2Y9_S_IO4/S4END[7] Tile_X2Y9_S_IO4/S4END[8]
+ Tile_X2Y9_S_IO4/S4END[9] Tile_X2Y9_S_IO4/SS4END[0] Tile_X2Y9_S_IO4/SS4END[10] Tile_X2Y9_S_IO4/SS4END[11]
+ Tile_X2Y9_S_IO4/SS4END[12] Tile_X2Y9_S_IO4/SS4END[13] Tile_X2Y9_S_IO4/SS4END[14]
+ Tile_X2Y9_S_IO4/SS4END[15] Tile_X2Y9_S_IO4/SS4END[1] Tile_X2Y9_S_IO4/SS4END[2] Tile_X2Y9_S_IO4/SS4END[3]
+ Tile_X2Y9_S_IO4/SS4END[4] Tile_X2Y9_S_IO4/SS4END[5] Tile_X2Y9_S_IO4/SS4END[6] Tile_X2Y9_S_IO4/SS4END[7]
+ Tile_X2Y9_S_IO4/SS4END[8] Tile_X2Y9_S_IO4/SS4END[9] UserCLK Tile_X2Y9_S_IO4/UserCLKo
+ VGND VPWR S_IO4
XTile_X5Y9_SE_term Tile_X5Y9_SE_term/FrameData[0] Tile_X5Y9_SE_term/FrameData[10]
+ Tile_X5Y9_SE_term/FrameData[11] Tile_X5Y9_SE_term/FrameData[12] Tile_X5Y9_SE_term/FrameData[13]
+ Tile_X5Y9_SE_term/FrameData[14] Tile_X5Y9_SE_term/FrameData[15] Tile_X5Y9_SE_term/FrameData[16]
+ Tile_X5Y9_SE_term/FrameData[17] Tile_X5Y9_SE_term/FrameData[18] Tile_X5Y9_SE_term/FrameData[19]
+ Tile_X5Y9_SE_term/FrameData[1] Tile_X5Y9_SE_term/FrameData[20] Tile_X5Y9_SE_term/FrameData[21]
+ Tile_X5Y9_SE_term/FrameData[22] Tile_X5Y9_SE_term/FrameData[23] Tile_X5Y9_SE_term/FrameData[24]
+ Tile_X5Y9_SE_term/FrameData[25] Tile_X5Y9_SE_term/FrameData[26] Tile_X5Y9_SE_term/FrameData[27]
+ Tile_X5Y9_SE_term/FrameData[28] Tile_X5Y9_SE_term/FrameData[29] Tile_X5Y9_SE_term/FrameData[2]
+ Tile_X5Y9_SE_term/FrameData[30] Tile_X5Y9_SE_term/FrameData[31] Tile_X5Y9_SE_term/FrameData[3]
+ Tile_X5Y9_SE_term/FrameData[4] Tile_X5Y9_SE_term/FrameData[5] Tile_X5Y9_SE_term/FrameData[6]
+ Tile_X5Y9_SE_term/FrameData[7] Tile_X5Y9_SE_term/FrameData[8] Tile_X5Y9_SE_term/FrameData[9]
+ Tile_X5Y9_SE_term/FrameData_O[0] Tile_X5Y9_SE_term/FrameData_O[10] Tile_X5Y9_SE_term/FrameData_O[11]
+ Tile_X5Y9_SE_term/FrameData_O[12] Tile_X5Y9_SE_term/FrameData_O[13] Tile_X5Y9_SE_term/FrameData_O[14]
+ Tile_X5Y9_SE_term/FrameData_O[15] Tile_X5Y9_SE_term/FrameData_O[16] Tile_X5Y9_SE_term/FrameData_O[17]
+ Tile_X5Y9_SE_term/FrameData_O[18] Tile_X5Y9_SE_term/FrameData_O[19] Tile_X5Y9_SE_term/FrameData_O[1]
+ Tile_X5Y9_SE_term/FrameData_O[20] Tile_X5Y9_SE_term/FrameData_O[21] Tile_X5Y9_SE_term/FrameData_O[22]
+ Tile_X5Y9_SE_term/FrameData_O[23] Tile_X5Y9_SE_term/FrameData_O[24] Tile_X5Y9_SE_term/FrameData_O[25]
+ Tile_X5Y9_SE_term/FrameData_O[26] Tile_X5Y9_SE_term/FrameData_O[27] Tile_X5Y9_SE_term/FrameData_O[28]
+ Tile_X5Y9_SE_term/FrameData_O[29] Tile_X5Y9_SE_term/FrameData_O[2] Tile_X5Y9_SE_term/FrameData_O[30]
+ Tile_X5Y9_SE_term/FrameData_O[31] Tile_X5Y9_SE_term/FrameData_O[3] Tile_X5Y9_SE_term/FrameData_O[4]
+ Tile_X5Y9_SE_term/FrameData_O[5] Tile_X5Y9_SE_term/FrameData_O[6] Tile_X5Y9_SE_term/FrameData_O[7]
+ Tile_X5Y9_SE_term/FrameData_O[8] Tile_X5Y9_SE_term/FrameData_O[9] FrameStrobe[100]
+ FrameStrobe[110] FrameStrobe[111] FrameStrobe[112] FrameStrobe[113] FrameStrobe[114]
+ FrameStrobe[115] FrameStrobe[116] FrameStrobe[117] FrameStrobe[118] FrameStrobe[119]
+ FrameStrobe[101] FrameStrobe[102] FrameStrobe[103] FrameStrobe[104] FrameStrobe[105]
+ FrameStrobe[106] FrameStrobe[107] FrameStrobe[108] FrameStrobe[109] Tile_X5Y8_E_TT_IF/FrameStrobe[0]
+ Tile_X5Y8_E_TT_IF/FrameStrobe[10] Tile_X5Y8_E_TT_IF/FrameStrobe[11] Tile_X5Y8_E_TT_IF/FrameStrobe[12]
+ Tile_X5Y8_E_TT_IF/FrameStrobe[13] Tile_X5Y8_E_TT_IF/FrameStrobe[14] Tile_X5Y8_E_TT_IF/FrameStrobe[15]
+ Tile_X5Y8_E_TT_IF/FrameStrobe[16] Tile_X5Y8_E_TT_IF/FrameStrobe[17] Tile_X5Y8_E_TT_IF/FrameStrobe[18]
+ Tile_X5Y8_E_TT_IF/FrameStrobe[19] Tile_X5Y8_E_TT_IF/FrameStrobe[1] Tile_X5Y8_E_TT_IF/FrameStrobe[2]
+ Tile_X5Y8_E_TT_IF/FrameStrobe[3] Tile_X5Y8_E_TT_IF/FrameStrobe[4] Tile_X5Y8_E_TT_IF/FrameStrobe[5]
+ Tile_X5Y8_E_TT_IF/FrameStrobe[6] Tile_X5Y8_E_TT_IF/FrameStrobe[7] Tile_X5Y8_E_TT_IF/FrameStrobe[8]
+ Tile_X5Y8_E_TT_IF/FrameStrobe[9] Tile_X5Y9_SE_term/N1BEG[0] Tile_X5Y9_SE_term/N1BEG[1]
+ Tile_X5Y9_SE_term/N1BEG[2] Tile_X5Y9_SE_term/N1BEG[3] Tile_X5Y9_SE_term/N2BEG[0]
+ Tile_X5Y9_SE_term/N2BEG[1] Tile_X5Y9_SE_term/N2BEG[2] Tile_X5Y9_SE_term/N2BEG[3]
+ Tile_X5Y9_SE_term/N2BEG[4] Tile_X5Y9_SE_term/N2BEG[5] Tile_X5Y9_SE_term/N2BEG[6]
+ Tile_X5Y9_SE_term/N2BEG[7] Tile_X5Y8_E_TT_IF/N2END[0] Tile_X5Y8_E_TT_IF/N2END[1]
+ Tile_X5Y8_E_TT_IF/N2END[2] Tile_X5Y8_E_TT_IF/N2END[3] Tile_X5Y8_E_TT_IF/N2END[4]
+ Tile_X5Y8_E_TT_IF/N2END[5] Tile_X5Y8_E_TT_IF/N2END[6] Tile_X5Y8_E_TT_IF/N2END[7]
+ Tile_X5Y9_SE_term/N4BEG[0] Tile_X5Y9_SE_term/N4BEG[10] Tile_X5Y9_SE_term/N4BEG[11]
+ Tile_X5Y9_SE_term/N4BEG[12] Tile_X5Y9_SE_term/N4BEG[13] Tile_X5Y9_SE_term/N4BEG[14]
+ Tile_X5Y9_SE_term/N4BEG[15] Tile_X5Y9_SE_term/N4BEG[1] Tile_X5Y9_SE_term/N4BEG[2]
+ Tile_X5Y9_SE_term/N4BEG[3] Tile_X5Y9_SE_term/N4BEG[4] Tile_X5Y9_SE_term/N4BEG[5]
+ Tile_X5Y9_SE_term/N4BEG[6] Tile_X5Y9_SE_term/N4BEG[7] Tile_X5Y9_SE_term/N4BEG[8]
+ Tile_X5Y9_SE_term/N4BEG[9] Tile_X5Y9_SE_term/S1END[0] Tile_X5Y9_SE_term/S1END[1]
+ Tile_X5Y9_SE_term/S1END[2] Tile_X5Y9_SE_term/S1END[3] Tile_X5Y9_SE_term/S2END[0]
+ Tile_X5Y9_SE_term/S2END[1] Tile_X5Y9_SE_term/S2END[2] Tile_X5Y9_SE_term/S2END[3]
+ Tile_X5Y9_SE_term/S2END[4] Tile_X5Y9_SE_term/S2END[5] Tile_X5Y9_SE_term/S2END[6]
+ Tile_X5Y9_SE_term/S2END[7] Tile_X5Y9_SE_term/S2MID[0] Tile_X5Y9_SE_term/S2MID[1]
+ Tile_X5Y9_SE_term/S2MID[2] Tile_X5Y9_SE_term/S2MID[3] Tile_X5Y9_SE_term/S2MID[4]
+ Tile_X5Y9_SE_term/S2MID[5] Tile_X5Y9_SE_term/S2MID[6] Tile_X5Y9_SE_term/S2MID[7]
+ Tile_X5Y9_SE_term/S4END[0] Tile_X5Y9_SE_term/S4END[10] Tile_X5Y9_SE_term/S4END[11]
+ Tile_X5Y9_SE_term/S4END[12] Tile_X5Y9_SE_term/S4END[13] Tile_X5Y9_SE_term/S4END[14]
+ Tile_X5Y9_SE_term/S4END[15] Tile_X5Y9_SE_term/S4END[1] Tile_X5Y9_SE_term/S4END[2]
+ Tile_X5Y9_SE_term/S4END[3] Tile_X5Y9_SE_term/S4END[4] Tile_X5Y9_SE_term/S4END[5]
+ Tile_X5Y9_SE_term/S4END[6] Tile_X5Y9_SE_term/S4END[7] Tile_X5Y9_SE_term/S4END[8]
+ Tile_X5Y9_SE_term/S4END[9] UserCLK Tile_X5Y8_E_TT_IF/UserCLK VGND VPWR SE_term
XTile_X1Y2_LUT4AB Tile_X1Y3_LUT4AB/Co Tile_X1Y2_LUT4AB/Co Tile_X2Y2_LUT4AB/E1END[0]
+ Tile_X2Y2_LUT4AB/E1END[1] Tile_X2Y2_LUT4AB/E1END[2] Tile_X2Y2_LUT4AB/E1END[3] Tile_X1Y2_LUT4AB/E1END[0]
+ Tile_X1Y2_LUT4AB/E1END[1] Tile_X1Y2_LUT4AB/E1END[2] Tile_X1Y2_LUT4AB/E1END[3] Tile_X2Y2_LUT4AB/E2MID[0]
+ Tile_X2Y2_LUT4AB/E2MID[1] Tile_X2Y2_LUT4AB/E2MID[2] Tile_X2Y2_LUT4AB/E2MID[3] Tile_X2Y2_LUT4AB/E2MID[4]
+ Tile_X2Y2_LUT4AB/E2MID[5] Tile_X2Y2_LUT4AB/E2MID[6] Tile_X2Y2_LUT4AB/E2MID[7] Tile_X2Y2_LUT4AB/E2END[0]
+ Tile_X2Y2_LUT4AB/E2END[1] Tile_X2Y2_LUT4AB/E2END[2] Tile_X2Y2_LUT4AB/E2END[3] Tile_X2Y2_LUT4AB/E2END[4]
+ Tile_X2Y2_LUT4AB/E2END[5] Tile_X2Y2_LUT4AB/E2END[6] Tile_X2Y2_LUT4AB/E2END[7] Tile_X1Y2_LUT4AB/E2END[0]
+ Tile_X1Y2_LUT4AB/E2END[1] Tile_X1Y2_LUT4AB/E2END[2] Tile_X1Y2_LUT4AB/E2END[3] Tile_X1Y2_LUT4AB/E2END[4]
+ Tile_X1Y2_LUT4AB/E2END[5] Tile_X1Y2_LUT4AB/E2END[6] Tile_X1Y2_LUT4AB/E2END[7] Tile_X1Y2_LUT4AB/E2MID[0]
+ Tile_X1Y2_LUT4AB/E2MID[1] Tile_X1Y2_LUT4AB/E2MID[2] Tile_X1Y2_LUT4AB/E2MID[3] Tile_X1Y2_LUT4AB/E2MID[4]
+ Tile_X1Y2_LUT4AB/E2MID[5] Tile_X1Y2_LUT4AB/E2MID[6] Tile_X1Y2_LUT4AB/E2MID[7] Tile_X2Y2_LUT4AB/E6END[0]
+ Tile_X2Y2_LUT4AB/E6END[10] Tile_X2Y2_LUT4AB/E6END[11] Tile_X2Y2_LUT4AB/E6END[1]
+ Tile_X2Y2_LUT4AB/E6END[2] Tile_X2Y2_LUT4AB/E6END[3] Tile_X2Y2_LUT4AB/E6END[4] Tile_X2Y2_LUT4AB/E6END[5]
+ Tile_X2Y2_LUT4AB/E6END[6] Tile_X2Y2_LUT4AB/E6END[7] Tile_X2Y2_LUT4AB/E6END[8] Tile_X2Y2_LUT4AB/E6END[9]
+ Tile_X1Y2_LUT4AB/E6END[0] Tile_X1Y2_LUT4AB/E6END[10] Tile_X1Y2_LUT4AB/E6END[11]
+ Tile_X1Y2_LUT4AB/E6END[1] Tile_X1Y2_LUT4AB/E6END[2] Tile_X1Y2_LUT4AB/E6END[3] Tile_X1Y2_LUT4AB/E6END[4]
+ Tile_X1Y2_LUT4AB/E6END[5] Tile_X1Y2_LUT4AB/E6END[6] Tile_X1Y2_LUT4AB/E6END[7] Tile_X1Y2_LUT4AB/E6END[8]
+ Tile_X1Y2_LUT4AB/E6END[9] Tile_X2Y2_LUT4AB/EE4END[0] Tile_X2Y2_LUT4AB/EE4END[10]
+ Tile_X2Y2_LUT4AB/EE4END[11] Tile_X2Y2_LUT4AB/EE4END[12] Tile_X2Y2_LUT4AB/EE4END[13]
+ Tile_X2Y2_LUT4AB/EE4END[14] Tile_X2Y2_LUT4AB/EE4END[15] Tile_X2Y2_LUT4AB/EE4END[1]
+ Tile_X2Y2_LUT4AB/EE4END[2] Tile_X2Y2_LUT4AB/EE4END[3] Tile_X2Y2_LUT4AB/EE4END[4]
+ Tile_X2Y2_LUT4AB/EE4END[5] Tile_X2Y2_LUT4AB/EE4END[6] Tile_X2Y2_LUT4AB/EE4END[7]
+ Tile_X2Y2_LUT4AB/EE4END[8] Tile_X2Y2_LUT4AB/EE4END[9] Tile_X1Y2_LUT4AB/EE4END[0]
+ Tile_X1Y2_LUT4AB/EE4END[10] Tile_X1Y2_LUT4AB/EE4END[11] Tile_X1Y2_LUT4AB/EE4END[12]
+ Tile_X1Y2_LUT4AB/EE4END[13] Tile_X1Y2_LUT4AB/EE4END[14] Tile_X1Y2_LUT4AB/EE4END[15]
+ Tile_X1Y2_LUT4AB/EE4END[1] Tile_X1Y2_LUT4AB/EE4END[2] Tile_X1Y2_LUT4AB/EE4END[3]
+ Tile_X1Y2_LUT4AB/EE4END[4] Tile_X1Y2_LUT4AB/EE4END[5] Tile_X1Y2_LUT4AB/EE4END[6]
+ Tile_X1Y2_LUT4AB/EE4END[7] Tile_X1Y2_LUT4AB/EE4END[8] Tile_X1Y2_LUT4AB/EE4END[9]
+ Tile_X1Y2_LUT4AB/FrameData[0] Tile_X1Y2_LUT4AB/FrameData[10] Tile_X1Y2_LUT4AB/FrameData[11]
+ Tile_X1Y2_LUT4AB/FrameData[12] Tile_X1Y2_LUT4AB/FrameData[13] Tile_X1Y2_LUT4AB/FrameData[14]
+ Tile_X1Y2_LUT4AB/FrameData[15] Tile_X1Y2_LUT4AB/FrameData[16] Tile_X1Y2_LUT4AB/FrameData[17]
+ Tile_X1Y2_LUT4AB/FrameData[18] Tile_X1Y2_LUT4AB/FrameData[19] Tile_X1Y2_LUT4AB/FrameData[1]
+ Tile_X1Y2_LUT4AB/FrameData[20] Tile_X1Y2_LUT4AB/FrameData[21] Tile_X1Y2_LUT4AB/FrameData[22]
+ Tile_X1Y2_LUT4AB/FrameData[23] Tile_X1Y2_LUT4AB/FrameData[24] Tile_X1Y2_LUT4AB/FrameData[25]
+ Tile_X1Y2_LUT4AB/FrameData[26] Tile_X1Y2_LUT4AB/FrameData[27] Tile_X1Y2_LUT4AB/FrameData[28]
+ Tile_X1Y2_LUT4AB/FrameData[29] Tile_X1Y2_LUT4AB/FrameData[2] Tile_X1Y2_LUT4AB/FrameData[30]
+ Tile_X1Y2_LUT4AB/FrameData[31] Tile_X1Y2_LUT4AB/FrameData[3] Tile_X1Y2_LUT4AB/FrameData[4]
+ Tile_X1Y2_LUT4AB/FrameData[5] Tile_X1Y2_LUT4AB/FrameData[6] Tile_X1Y2_LUT4AB/FrameData[7]
+ Tile_X1Y2_LUT4AB/FrameData[8] Tile_X1Y2_LUT4AB/FrameData[9] Tile_X2Y2_LUT4AB/FrameData[0]
+ Tile_X2Y2_LUT4AB/FrameData[10] Tile_X2Y2_LUT4AB/FrameData[11] Tile_X2Y2_LUT4AB/FrameData[12]
+ Tile_X2Y2_LUT4AB/FrameData[13] Tile_X2Y2_LUT4AB/FrameData[14] Tile_X2Y2_LUT4AB/FrameData[15]
+ Tile_X2Y2_LUT4AB/FrameData[16] Tile_X2Y2_LUT4AB/FrameData[17] Tile_X2Y2_LUT4AB/FrameData[18]
+ Tile_X2Y2_LUT4AB/FrameData[19] Tile_X2Y2_LUT4AB/FrameData[1] Tile_X2Y2_LUT4AB/FrameData[20]
+ Tile_X2Y2_LUT4AB/FrameData[21] Tile_X2Y2_LUT4AB/FrameData[22] Tile_X2Y2_LUT4AB/FrameData[23]
+ Tile_X2Y2_LUT4AB/FrameData[24] Tile_X2Y2_LUT4AB/FrameData[25] Tile_X2Y2_LUT4AB/FrameData[26]
+ Tile_X2Y2_LUT4AB/FrameData[27] Tile_X2Y2_LUT4AB/FrameData[28] Tile_X2Y2_LUT4AB/FrameData[29]
+ Tile_X2Y2_LUT4AB/FrameData[2] Tile_X2Y2_LUT4AB/FrameData[30] Tile_X2Y2_LUT4AB/FrameData[31]
+ Tile_X2Y2_LUT4AB/FrameData[3] Tile_X2Y2_LUT4AB/FrameData[4] Tile_X2Y2_LUT4AB/FrameData[5]
+ Tile_X2Y2_LUT4AB/FrameData[6] Tile_X2Y2_LUT4AB/FrameData[7] Tile_X2Y2_LUT4AB/FrameData[8]
+ Tile_X2Y2_LUT4AB/FrameData[9] Tile_X1Y2_LUT4AB/FrameStrobe[0] Tile_X1Y2_LUT4AB/FrameStrobe[10]
+ Tile_X1Y2_LUT4AB/FrameStrobe[11] Tile_X1Y2_LUT4AB/FrameStrobe[12] Tile_X1Y2_LUT4AB/FrameStrobe[13]
+ Tile_X1Y2_LUT4AB/FrameStrobe[14] Tile_X1Y2_LUT4AB/FrameStrobe[15] Tile_X1Y2_LUT4AB/FrameStrobe[16]
+ Tile_X1Y2_LUT4AB/FrameStrobe[17] Tile_X1Y2_LUT4AB/FrameStrobe[18] Tile_X1Y2_LUT4AB/FrameStrobe[19]
+ Tile_X1Y2_LUT4AB/FrameStrobe[1] Tile_X1Y2_LUT4AB/FrameStrobe[2] Tile_X1Y2_LUT4AB/FrameStrobe[3]
+ Tile_X1Y2_LUT4AB/FrameStrobe[4] Tile_X1Y2_LUT4AB/FrameStrobe[5] Tile_X1Y2_LUT4AB/FrameStrobe[6]
+ Tile_X1Y2_LUT4AB/FrameStrobe[7] Tile_X1Y2_LUT4AB/FrameStrobe[8] Tile_X1Y2_LUT4AB/FrameStrobe[9]
+ Tile_X1Y1_LUT4AB/FrameStrobe[0] Tile_X1Y1_LUT4AB/FrameStrobe[10] Tile_X1Y1_LUT4AB/FrameStrobe[11]
+ Tile_X1Y1_LUT4AB/FrameStrobe[12] Tile_X1Y1_LUT4AB/FrameStrobe[13] Tile_X1Y1_LUT4AB/FrameStrobe[14]
+ Tile_X1Y1_LUT4AB/FrameStrobe[15] Tile_X1Y1_LUT4AB/FrameStrobe[16] Tile_X1Y1_LUT4AB/FrameStrobe[17]
+ Tile_X1Y1_LUT4AB/FrameStrobe[18] Tile_X1Y1_LUT4AB/FrameStrobe[19] Tile_X1Y1_LUT4AB/FrameStrobe[1]
+ Tile_X1Y1_LUT4AB/FrameStrobe[2] Tile_X1Y1_LUT4AB/FrameStrobe[3] Tile_X1Y1_LUT4AB/FrameStrobe[4]
+ Tile_X1Y1_LUT4AB/FrameStrobe[5] Tile_X1Y1_LUT4AB/FrameStrobe[6] Tile_X1Y1_LUT4AB/FrameStrobe[7]
+ Tile_X1Y1_LUT4AB/FrameStrobe[8] Tile_X1Y1_LUT4AB/FrameStrobe[9] Tile_X1Y2_LUT4AB/N1BEG[0]
+ Tile_X1Y2_LUT4AB/N1BEG[1] Tile_X1Y2_LUT4AB/N1BEG[2] Tile_X1Y2_LUT4AB/N1BEG[3] Tile_X1Y3_LUT4AB/N1BEG[0]
+ Tile_X1Y3_LUT4AB/N1BEG[1] Tile_X1Y3_LUT4AB/N1BEG[2] Tile_X1Y3_LUT4AB/N1BEG[3] Tile_X1Y2_LUT4AB/N2BEG[0]
+ Tile_X1Y2_LUT4AB/N2BEG[1] Tile_X1Y2_LUT4AB/N2BEG[2] Tile_X1Y2_LUT4AB/N2BEG[3] Tile_X1Y2_LUT4AB/N2BEG[4]
+ Tile_X1Y2_LUT4AB/N2BEG[5] Tile_X1Y2_LUT4AB/N2BEG[6] Tile_X1Y2_LUT4AB/N2BEG[7] Tile_X1Y1_LUT4AB/N2END[0]
+ Tile_X1Y1_LUT4AB/N2END[1] Tile_X1Y1_LUT4AB/N2END[2] Tile_X1Y1_LUT4AB/N2END[3] Tile_X1Y1_LUT4AB/N2END[4]
+ Tile_X1Y1_LUT4AB/N2END[5] Tile_X1Y1_LUT4AB/N2END[6] Tile_X1Y1_LUT4AB/N2END[7] Tile_X1Y2_LUT4AB/N2END[0]
+ Tile_X1Y2_LUT4AB/N2END[1] Tile_X1Y2_LUT4AB/N2END[2] Tile_X1Y2_LUT4AB/N2END[3] Tile_X1Y2_LUT4AB/N2END[4]
+ Tile_X1Y2_LUT4AB/N2END[5] Tile_X1Y2_LUT4AB/N2END[6] Tile_X1Y2_LUT4AB/N2END[7] Tile_X1Y3_LUT4AB/N2BEG[0]
+ Tile_X1Y3_LUT4AB/N2BEG[1] Tile_X1Y3_LUT4AB/N2BEG[2] Tile_X1Y3_LUT4AB/N2BEG[3] Tile_X1Y3_LUT4AB/N2BEG[4]
+ Tile_X1Y3_LUT4AB/N2BEG[5] Tile_X1Y3_LUT4AB/N2BEG[6] Tile_X1Y3_LUT4AB/N2BEG[7] Tile_X1Y2_LUT4AB/N4BEG[0]
+ Tile_X1Y2_LUT4AB/N4BEG[10] Tile_X1Y2_LUT4AB/N4BEG[11] Tile_X1Y2_LUT4AB/N4BEG[12]
+ Tile_X1Y2_LUT4AB/N4BEG[13] Tile_X1Y2_LUT4AB/N4BEG[14] Tile_X1Y2_LUT4AB/N4BEG[15]
+ Tile_X1Y2_LUT4AB/N4BEG[1] Tile_X1Y2_LUT4AB/N4BEG[2] Tile_X1Y2_LUT4AB/N4BEG[3] Tile_X1Y2_LUT4AB/N4BEG[4]
+ Tile_X1Y2_LUT4AB/N4BEG[5] Tile_X1Y2_LUT4AB/N4BEG[6] Tile_X1Y2_LUT4AB/N4BEG[7] Tile_X1Y2_LUT4AB/N4BEG[8]
+ Tile_X1Y2_LUT4AB/N4BEG[9] Tile_X1Y3_LUT4AB/N4BEG[0] Tile_X1Y3_LUT4AB/N4BEG[10] Tile_X1Y3_LUT4AB/N4BEG[11]
+ Tile_X1Y3_LUT4AB/N4BEG[12] Tile_X1Y3_LUT4AB/N4BEG[13] Tile_X1Y3_LUT4AB/N4BEG[14]
+ Tile_X1Y3_LUT4AB/N4BEG[15] Tile_X1Y3_LUT4AB/N4BEG[1] Tile_X1Y3_LUT4AB/N4BEG[2] Tile_X1Y3_LUT4AB/N4BEG[3]
+ Tile_X1Y3_LUT4AB/N4BEG[4] Tile_X1Y3_LUT4AB/N4BEG[5] Tile_X1Y3_LUT4AB/N4BEG[6] Tile_X1Y3_LUT4AB/N4BEG[7]
+ Tile_X1Y3_LUT4AB/N4BEG[8] Tile_X1Y3_LUT4AB/N4BEG[9] Tile_X1Y2_LUT4AB/NN4BEG[0] Tile_X1Y2_LUT4AB/NN4BEG[10]
+ Tile_X1Y2_LUT4AB/NN4BEG[11] Tile_X1Y2_LUT4AB/NN4BEG[12] Tile_X1Y2_LUT4AB/NN4BEG[13]
+ Tile_X1Y2_LUT4AB/NN4BEG[14] Tile_X1Y2_LUT4AB/NN4BEG[15] Tile_X1Y2_LUT4AB/NN4BEG[1]
+ Tile_X1Y2_LUT4AB/NN4BEG[2] Tile_X1Y2_LUT4AB/NN4BEG[3] Tile_X1Y2_LUT4AB/NN4BEG[4]
+ Tile_X1Y2_LUT4AB/NN4BEG[5] Tile_X1Y2_LUT4AB/NN4BEG[6] Tile_X1Y2_LUT4AB/NN4BEG[7]
+ Tile_X1Y2_LUT4AB/NN4BEG[8] Tile_X1Y2_LUT4AB/NN4BEG[9] Tile_X1Y3_LUT4AB/NN4BEG[0]
+ Tile_X1Y3_LUT4AB/NN4BEG[10] Tile_X1Y3_LUT4AB/NN4BEG[11] Tile_X1Y3_LUT4AB/NN4BEG[12]
+ Tile_X1Y3_LUT4AB/NN4BEG[13] Tile_X1Y3_LUT4AB/NN4BEG[14] Tile_X1Y3_LUT4AB/NN4BEG[15]
+ Tile_X1Y3_LUT4AB/NN4BEG[1] Tile_X1Y3_LUT4AB/NN4BEG[2] Tile_X1Y3_LUT4AB/NN4BEG[3]
+ Tile_X1Y3_LUT4AB/NN4BEG[4] Tile_X1Y3_LUT4AB/NN4BEG[5] Tile_X1Y3_LUT4AB/NN4BEG[6]
+ Tile_X1Y3_LUT4AB/NN4BEG[7] Tile_X1Y3_LUT4AB/NN4BEG[8] Tile_X1Y3_LUT4AB/NN4BEG[9]
+ Tile_X1Y3_LUT4AB/S1END[0] Tile_X1Y3_LUT4AB/S1END[1] Tile_X1Y3_LUT4AB/S1END[2] Tile_X1Y3_LUT4AB/S1END[3]
+ Tile_X1Y2_LUT4AB/S1END[0] Tile_X1Y2_LUT4AB/S1END[1] Tile_X1Y2_LUT4AB/S1END[2] Tile_X1Y2_LUT4AB/S1END[3]
+ Tile_X1Y3_LUT4AB/S2MID[0] Tile_X1Y3_LUT4AB/S2MID[1] Tile_X1Y3_LUT4AB/S2MID[2] Tile_X1Y3_LUT4AB/S2MID[3]
+ Tile_X1Y3_LUT4AB/S2MID[4] Tile_X1Y3_LUT4AB/S2MID[5] Tile_X1Y3_LUT4AB/S2MID[6] Tile_X1Y3_LUT4AB/S2MID[7]
+ Tile_X1Y3_LUT4AB/S2END[0] Tile_X1Y3_LUT4AB/S2END[1] Tile_X1Y3_LUT4AB/S2END[2] Tile_X1Y3_LUT4AB/S2END[3]
+ Tile_X1Y3_LUT4AB/S2END[4] Tile_X1Y3_LUT4AB/S2END[5] Tile_X1Y3_LUT4AB/S2END[6] Tile_X1Y3_LUT4AB/S2END[7]
+ Tile_X1Y2_LUT4AB/S2END[0] Tile_X1Y2_LUT4AB/S2END[1] Tile_X1Y2_LUT4AB/S2END[2] Tile_X1Y2_LUT4AB/S2END[3]
+ Tile_X1Y2_LUT4AB/S2END[4] Tile_X1Y2_LUT4AB/S2END[5] Tile_X1Y2_LUT4AB/S2END[6] Tile_X1Y2_LUT4AB/S2END[7]
+ Tile_X1Y2_LUT4AB/S2MID[0] Tile_X1Y2_LUT4AB/S2MID[1] Tile_X1Y2_LUT4AB/S2MID[2] Tile_X1Y2_LUT4AB/S2MID[3]
+ Tile_X1Y2_LUT4AB/S2MID[4] Tile_X1Y2_LUT4AB/S2MID[5] Tile_X1Y2_LUT4AB/S2MID[6] Tile_X1Y2_LUT4AB/S2MID[7]
+ Tile_X1Y3_LUT4AB/S4END[0] Tile_X1Y3_LUT4AB/S4END[10] Tile_X1Y3_LUT4AB/S4END[11]
+ Tile_X1Y3_LUT4AB/S4END[12] Tile_X1Y3_LUT4AB/S4END[13] Tile_X1Y3_LUT4AB/S4END[14]
+ Tile_X1Y3_LUT4AB/S4END[15] Tile_X1Y3_LUT4AB/S4END[1] Tile_X1Y3_LUT4AB/S4END[2] Tile_X1Y3_LUT4AB/S4END[3]
+ Tile_X1Y3_LUT4AB/S4END[4] Tile_X1Y3_LUT4AB/S4END[5] Tile_X1Y3_LUT4AB/S4END[6] Tile_X1Y3_LUT4AB/S4END[7]
+ Tile_X1Y3_LUT4AB/S4END[8] Tile_X1Y3_LUT4AB/S4END[9] Tile_X1Y2_LUT4AB/S4END[0] Tile_X1Y2_LUT4AB/S4END[10]
+ Tile_X1Y2_LUT4AB/S4END[11] Tile_X1Y2_LUT4AB/S4END[12] Tile_X1Y2_LUT4AB/S4END[13]
+ Tile_X1Y2_LUT4AB/S4END[14] Tile_X1Y2_LUT4AB/S4END[15] Tile_X1Y2_LUT4AB/S4END[1]
+ Tile_X1Y2_LUT4AB/S4END[2] Tile_X1Y2_LUT4AB/S4END[3] Tile_X1Y2_LUT4AB/S4END[4] Tile_X1Y2_LUT4AB/S4END[5]
+ Tile_X1Y2_LUT4AB/S4END[6] Tile_X1Y2_LUT4AB/S4END[7] Tile_X1Y2_LUT4AB/S4END[8] Tile_X1Y2_LUT4AB/S4END[9]
+ Tile_X1Y3_LUT4AB/SS4END[0] Tile_X1Y3_LUT4AB/SS4END[10] Tile_X1Y3_LUT4AB/SS4END[11]
+ Tile_X1Y3_LUT4AB/SS4END[12] Tile_X1Y3_LUT4AB/SS4END[13] Tile_X1Y3_LUT4AB/SS4END[14]
+ Tile_X1Y3_LUT4AB/SS4END[15] Tile_X1Y3_LUT4AB/SS4END[1] Tile_X1Y3_LUT4AB/SS4END[2]
+ Tile_X1Y3_LUT4AB/SS4END[3] Tile_X1Y3_LUT4AB/SS4END[4] Tile_X1Y3_LUT4AB/SS4END[5]
+ Tile_X1Y3_LUT4AB/SS4END[6] Tile_X1Y3_LUT4AB/SS4END[7] Tile_X1Y3_LUT4AB/SS4END[8]
+ Tile_X1Y3_LUT4AB/SS4END[9] Tile_X1Y2_LUT4AB/SS4END[0] Tile_X1Y2_LUT4AB/SS4END[10]
+ Tile_X1Y2_LUT4AB/SS4END[11] Tile_X1Y2_LUT4AB/SS4END[12] Tile_X1Y2_LUT4AB/SS4END[13]
+ Tile_X1Y2_LUT4AB/SS4END[14] Tile_X1Y2_LUT4AB/SS4END[15] Tile_X1Y2_LUT4AB/SS4END[1]
+ Tile_X1Y2_LUT4AB/SS4END[2] Tile_X1Y2_LUT4AB/SS4END[3] Tile_X1Y2_LUT4AB/SS4END[4]
+ Tile_X1Y2_LUT4AB/SS4END[5] Tile_X1Y2_LUT4AB/SS4END[6] Tile_X1Y2_LUT4AB/SS4END[7]
+ Tile_X1Y2_LUT4AB/SS4END[8] Tile_X1Y2_LUT4AB/SS4END[9] Tile_X1Y2_LUT4AB/UserCLK Tile_X1Y1_LUT4AB/UserCLK
+ VGND VPWR Tile_X1Y2_LUT4AB/W1BEG[0] Tile_X1Y2_LUT4AB/W1BEG[1] Tile_X1Y2_LUT4AB/W1BEG[2]
+ Tile_X1Y2_LUT4AB/W1BEG[3] Tile_X2Y2_LUT4AB/W1BEG[0] Tile_X2Y2_LUT4AB/W1BEG[1] Tile_X2Y2_LUT4AB/W1BEG[2]
+ Tile_X2Y2_LUT4AB/W1BEG[3] Tile_X1Y2_LUT4AB/W2BEG[0] Tile_X1Y2_LUT4AB/W2BEG[1] Tile_X1Y2_LUT4AB/W2BEG[2]
+ Tile_X1Y2_LUT4AB/W2BEG[3] Tile_X1Y2_LUT4AB/W2BEG[4] Tile_X1Y2_LUT4AB/W2BEG[5] Tile_X1Y2_LUT4AB/W2BEG[6]
+ Tile_X1Y2_LUT4AB/W2BEG[7] Tile_X1Y2_LUT4AB/W2BEGb[0] Tile_X1Y2_LUT4AB/W2BEGb[1]
+ Tile_X1Y2_LUT4AB/W2BEGb[2] Tile_X1Y2_LUT4AB/W2BEGb[3] Tile_X1Y2_LUT4AB/W2BEGb[4]
+ Tile_X1Y2_LUT4AB/W2BEGb[5] Tile_X1Y2_LUT4AB/W2BEGb[6] Tile_X1Y2_LUT4AB/W2BEGb[7]
+ Tile_X1Y2_LUT4AB/W2END[0] Tile_X1Y2_LUT4AB/W2END[1] Tile_X1Y2_LUT4AB/W2END[2] Tile_X1Y2_LUT4AB/W2END[3]
+ Tile_X1Y2_LUT4AB/W2END[4] Tile_X1Y2_LUT4AB/W2END[5] Tile_X1Y2_LUT4AB/W2END[6] Tile_X1Y2_LUT4AB/W2END[7]
+ Tile_X2Y2_LUT4AB/W2BEG[0] Tile_X2Y2_LUT4AB/W2BEG[1] Tile_X2Y2_LUT4AB/W2BEG[2] Tile_X2Y2_LUT4AB/W2BEG[3]
+ Tile_X2Y2_LUT4AB/W2BEG[4] Tile_X2Y2_LUT4AB/W2BEG[5] Tile_X2Y2_LUT4AB/W2BEG[6] Tile_X2Y2_LUT4AB/W2BEG[7]
+ Tile_X1Y2_LUT4AB/W6BEG[0] Tile_X1Y2_LUT4AB/W6BEG[10] Tile_X1Y2_LUT4AB/W6BEG[11]
+ Tile_X1Y2_LUT4AB/W6BEG[1] Tile_X1Y2_LUT4AB/W6BEG[2] Tile_X1Y2_LUT4AB/W6BEG[3] Tile_X1Y2_LUT4AB/W6BEG[4]
+ Tile_X1Y2_LUT4AB/W6BEG[5] Tile_X1Y2_LUT4AB/W6BEG[6] Tile_X1Y2_LUT4AB/W6BEG[7] Tile_X1Y2_LUT4AB/W6BEG[8]
+ Tile_X1Y2_LUT4AB/W6BEG[9] Tile_X2Y2_LUT4AB/W6BEG[0] Tile_X2Y2_LUT4AB/W6BEG[10] Tile_X2Y2_LUT4AB/W6BEG[11]
+ Tile_X2Y2_LUT4AB/W6BEG[1] Tile_X2Y2_LUT4AB/W6BEG[2] Tile_X2Y2_LUT4AB/W6BEG[3] Tile_X2Y2_LUT4AB/W6BEG[4]
+ Tile_X2Y2_LUT4AB/W6BEG[5] Tile_X2Y2_LUT4AB/W6BEG[6] Tile_X2Y2_LUT4AB/W6BEG[7] Tile_X2Y2_LUT4AB/W6BEG[8]
+ Tile_X2Y2_LUT4AB/W6BEG[9] Tile_X1Y2_LUT4AB/WW4BEG[0] Tile_X1Y2_LUT4AB/WW4BEG[10]
+ Tile_X1Y2_LUT4AB/WW4BEG[11] Tile_X1Y2_LUT4AB/WW4BEG[12] Tile_X1Y2_LUT4AB/WW4BEG[13]
+ Tile_X1Y2_LUT4AB/WW4BEG[14] Tile_X1Y2_LUT4AB/WW4BEG[15] Tile_X1Y2_LUT4AB/WW4BEG[1]
+ Tile_X1Y2_LUT4AB/WW4BEG[2] Tile_X1Y2_LUT4AB/WW4BEG[3] Tile_X1Y2_LUT4AB/WW4BEG[4]
+ Tile_X1Y2_LUT4AB/WW4BEG[5] Tile_X1Y2_LUT4AB/WW4BEG[6] Tile_X1Y2_LUT4AB/WW4BEG[7]
+ Tile_X1Y2_LUT4AB/WW4BEG[8] Tile_X1Y2_LUT4AB/WW4BEG[9] Tile_X2Y2_LUT4AB/WW4BEG[0]
+ Tile_X2Y2_LUT4AB/WW4BEG[10] Tile_X2Y2_LUT4AB/WW4BEG[11] Tile_X2Y2_LUT4AB/WW4BEG[12]
+ Tile_X2Y2_LUT4AB/WW4BEG[13] Tile_X2Y2_LUT4AB/WW4BEG[14] Tile_X2Y2_LUT4AB/WW4BEG[15]
+ Tile_X2Y2_LUT4AB/WW4BEG[1] Tile_X2Y2_LUT4AB/WW4BEG[2] Tile_X2Y2_LUT4AB/WW4BEG[3]
+ Tile_X2Y2_LUT4AB/WW4BEG[4] Tile_X2Y2_LUT4AB/WW4BEG[5] Tile_X2Y2_LUT4AB/WW4BEG[6]
+ Tile_X2Y2_LUT4AB/WW4BEG[7] Tile_X2Y2_LUT4AB/WW4BEG[8] Tile_X2Y2_LUT4AB/WW4BEG[9]
+ LUT4AB
XTile_X4Y7_LUT4AB Tile_X4Y8_LUT4AB/Co Tile_X4Y7_LUT4AB/Co Tile_X4Y7_LUT4AB/E1BEG[0]
+ Tile_X4Y7_LUT4AB/E1BEG[1] Tile_X4Y7_LUT4AB/E1BEG[2] Tile_X4Y7_LUT4AB/E1BEG[3] Tile_X4Y7_LUT4AB/E1END[0]
+ Tile_X4Y7_LUT4AB/E1END[1] Tile_X4Y7_LUT4AB/E1END[2] Tile_X4Y7_LUT4AB/E1END[3] Tile_X4Y7_LUT4AB/E2BEG[0]
+ Tile_X4Y7_LUT4AB/E2BEG[1] Tile_X4Y7_LUT4AB/E2BEG[2] Tile_X4Y7_LUT4AB/E2BEG[3] Tile_X4Y7_LUT4AB/E2BEG[4]
+ Tile_X4Y7_LUT4AB/E2BEG[5] Tile_X4Y7_LUT4AB/E2BEG[6] Tile_X4Y7_LUT4AB/E2BEG[7] Tile_X5Y7_E_TT_IF/E2END[0]
+ Tile_X5Y7_E_TT_IF/E2END[1] Tile_X5Y7_E_TT_IF/E2END[2] Tile_X5Y7_E_TT_IF/E2END[3]
+ Tile_X5Y7_E_TT_IF/E2END[4] Tile_X5Y7_E_TT_IF/E2END[5] Tile_X5Y7_E_TT_IF/E2END[6]
+ Tile_X5Y7_E_TT_IF/E2END[7] Tile_X4Y7_LUT4AB/E2END[0] Tile_X4Y7_LUT4AB/E2END[1] Tile_X4Y7_LUT4AB/E2END[2]
+ Tile_X4Y7_LUT4AB/E2END[3] Tile_X4Y7_LUT4AB/E2END[4] Tile_X4Y7_LUT4AB/E2END[5] Tile_X4Y7_LUT4AB/E2END[6]
+ Tile_X4Y7_LUT4AB/E2END[7] Tile_X4Y7_LUT4AB/E2MID[0] Tile_X4Y7_LUT4AB/E2MID[1] Tile_X4Y7_LUT4AB/E2MID[2]
+ Tile_X4Y7_LUT4AB/E2MID[3] Tile_X4Y7_LUT4AB/E2MID[4] Tile_X4Y7_LUT4AB/E2MID[5] Tile_X4Y7_LUT4AB/E2MID[6]
+ Tile_X4Y7_LUT4AB/E2MID[7] Tile_X4Y7_LUT4AB/E6BEG[0] Tile_X4Y7_LUT4AB/E6BEG[10] Tile_X4Y7_LUT4AB/E6BEG[11]
+ Tile_X4Y7_LUT4AB/E6BEG[1] Tile_X4Y7_LUT4AB/E6BEG[2] Tile_X4Y7_LUT4AB/E6BEG[3] Tile_X4Y7_LUT4AB/E6BEG[4]
+ Tile_X4Y7_LUT4AB/E6BEG[5] Tile_X4Y7_LUT4AB/E6BEG[6] Tile_X4Y7_LUT4AB/E6BEG[7] Tile_X4Y7_LUT4AB/E6BEG[8]
+ Tile_X4Y7_LUT4AB/E6BEG[9] Tile_X4Y7_LUT4AB/E6END[0] Tile_X4Y7_LUT4AB/E6END[10] Tile_X4Y7_LUT4AB/E6END[11]
+ Tile_X4Y7_LUT4AB/E6END[1] Tile_X4Y7_LUT4AB/E6END[2] Tile_X4Y7_LUT4AB/E6END[3] Tile_X4Y7_LUT4AB/E6END[4]
+ Tile_X4Y7_LUT4AB/E6END[5] Tile_X4Y7_LUT4AB/E6END[6] Tile_X4Y7_LUT4AB/E6END[7] Tile_X4Y7_LUT4AB/E6END[8]
+ Tile_X4Y7_LUT4AB/E6END[9] Tile_X4Y7_LUT4AB/EE4BEG[0] Tile_X4Y7_LUT4AB/EE4BEG[10]
+ Tile_X4Y7_LUT4AB/EE4BEG[11] Tile_X4Y7_LUT4AB/EE4BEG[12] Tile_X4Y7_LUT4AB/EE4BEG[13]
+ Tile_X4Y7_LUT4AB/EE4BEG[14] Tile_X4Y7_LUT4AB/EE4BEG[15] Tile_X4Y7_LUT4AB/EE4BEG[1]
+ Tile_X4Y7_LUT4AB/EE4BEG[2] Tile_X4Y7_LUT4AB/EE4BEG[3] Tile_X4Y7_LUT4AB/EE4BEG[4]
+ Tile_X4Y7_LUT4AB/EE4BEG[5] Tile_X4Y7_LUT4AB/EE4BEG[6] Tile_X4Y7_LUT4AB/EE4BEG[7]
+ Tile_X4Y7_LUT4AB/EE4BEG[8] Tile_X4Y7_LUT4AB/EE4BEG[9] Tile_X4Y7_LUT4AB/EE4END[0]
+ Tile_X4Y7_LUT4AB/EE4END[10] Tile_X4Y7_LUT4AB/EE4END[11] Tile_X4Y7_LUT4AB/EE4END[12]
+ Tile_X4Y7_LUT4AB/EE4END[13] Tile_X4Y7_LUT4AB/EE4END[14] Tile_X4Y7_LUT4AB/EE4END[15]
+ Tile_X4Y7_LUT4AB/EE4END[1] Tile_X4Y7_LUT4AB/EE4END[2] Tile_X4Y7_LUT4AB/EE4END[3]
+ Tile_X4Y7_LUT4AB/EE4END[4] Tile_X4Y7_LUT4AB/EE4END[5] Tile_X4Y7_LUT4AB/EE4END[6]
+ Tile_X4Y7_LUT4AB/EE4END[7] Tile_X4Y7_LUT4AB/EE4END[8] Tile_X4Y7_LUT4AB/EE4END[9]
+ Tile_X4Y7_LUT4AB/FrameData[0] Tile_X4Y7_LUT4AB/FrameData[10] Tile_X4Y7_LUT4AB/FrameData[11]
+ Tile_X4Y7_LUT4AB/FrameData[12] Tile_X4Y7_LUT4AB/FrameData[13] Tile_X4Y7_LUT4AB/FrameData[14]
+ Tile_X4Y7_LUT4AB/FrameData[15] Tile_X4Y7_LUT4AB/FrameData[16] Tile_X4Y7_LUT4AB/FrameData[17]
+ Tile_X4Y7_LUT4AB/FrameData[18] Tile_X4Y7_LUT4AB/FrameData[19] Tile_X4Y7_LUT4AB/FrameData[1]
+ Tile_X4Y7_LUT4AB/FrameData[20] Tile_X4Y7_LUT4AB/FrameData[21] Tile_X4Y7_LUT4AB/FrameData[22]
+ Tile_X4Y7_LUT4AB/FrameData[23] Tile_X4Y7_LUT4AB/FrameData[24] Tile_X4Y7_LUT4AB/FrameData[25]
+ Tile_X4Y7_LUT4AB/FrameData[26] Tile_X4Y7_LUT4AB/FrameData[27] Tile_X4Y7_LUT4AB/FrameData[28]
+ Tile_X4Y7_LUT4AB/FrameData[29] Tile_X4Y7_LUT4AB/FrameData[2] Tile_X4Y7_LUT4AB/FrameData[30]
+ Tile_X4Y7_LUT4AB/FrameData[31] Tile_X4Y7_LUT4AB/FrameData[3] Tile_X4Y7_LUT4AB/FrameData[4]
+ Tile_X4Y7_LUT4AB/FrameData[5] Tile_X4Y7_LUT4AB/FrameData[6] Tile_X4Y7_LUT4AB/FrameData[7]
+ Tile_X4Y7_LUT4AB/FrameData[8] Tile_X4Y7_LUT4AB/FrameData[9] Tile_X5Y7_E_TT_IF/FrameData[0]
+ Tile_X5Y7_E_TT_IF/FrameData[10] Tile_X5Y7_E_TT_IF/FrameData[11] Tile_X5Y7_E_TT_IF/FrameData[12]
+ Tile_X5Y7_E_TT_IF/FrameData[13] Tile_X5Y7_E_TT_IF/FrameData[14] Tile_X5Y7_E_TT_IF/FrameData[15]
+ Tile_X5Y7_E_TT_IF/FrameData[16] Tile_X5Y7_E_TT_IF/FrameData[17] Tile_X5Y7_E_TT_IF/FrameData[18]
+ Tile_X5Y7_E_TT_IF/FrameData[19] Tile_X5Y7_E_TT_IF/FrameData[1] Tile_X5Y7_E_TT_IF/FrameData[20]
+ Tile_X5Y7_E_TT_IF/FrameData[21] Tile_X5Y7_E_TT_IF/FrameData[22] Tile_X5Y7_E_TT_IF/FrameData[23]
+ Tile_X5Y7_E_TT_IF/FrameData[24] Tile_X5Y7_E_TT_IF/FrameData[25] Tile_X5Y7_E_TT_IF/FrameData[26]
+ Tile_X5Y7_E_TT_IF/FrameData[27] Tile_X5Y7_E_TT_IF/FrameData[28] Tile_X5Y7_E_TT_IF/FrameData[29]
+ Tile_X5Y7_E_TT_IF/FrameData[2] Tile_X5Y7_E_TT_IF/FrameData[30] Tile_X5Y7_E_TT_IF/FrameData[31]
+ Tile_X5Y7_E_TT_IF/FrameData[3] Tile_X5Y7_E_TT_IF/FrameData[4] Tile_X5Y7_E_TT_IF/FrameData[5]
+ Tile_X5Y7_E_TT_IF/FrameData[6] Tile_X5Y7_E_TT_IF/FrameData[7] Tile_X5Y7_E_TT_IF/FrameData[8]
+ Tile_X5Y7_E_TT_IF/FrameData[9] Tile_X4Y7_LUT4AB/FrameStrobe[0] Tile_X4Y7_LUT4AB/FrameStrobe[10]
+ Tile_X4Y7_LUT4AB/FrameStrobe[11] Tile_X4Y7_LUT4AB/FrameStrobe[12] Tile_X4Y7_LUT4AB/FrameStrobe[13]
+ Tile_X4Y7_LUT4AB/FrameStrobe[14] Tile_X4Y7_LUT4AB/FrameStrobe[15] Tile_X4Y7_LUT4AB/FrameStrobe[16]
+ Tile_X4Y7_LUT4AB/FrameStrobe[17] Tile_X4Y7_LUT4AB/FrameStrobe[18] Tile_X4Y7_LUT4AB/FrameStrobe[19]
+ Tile_X4Y7_LUT4AB/FrameStrobe[1] Tile_X4Y7_LUT4AB/FrameStrobe[2] Tile_X4Y7_LUT4AB/FrameStrobe[3]
+ Tile_X4Y7_LUT4AB/FrameStrobe[4] Tile_X4Y7_LUT4AB/FrameStrobe[5] Tile_X4Y7_LUT4AB/FrameStrobe[6]
+ Tile_X4Y7_LUT4AB/FrameStrobe[7] Tile_X4Y7_LUT4AB/FrameStrobe[8] Tile_X4Y7_LUT4AB/FrameStrobe[9]
+ Tile_X4Y6_LUT4AB/FrameStrobe[0] Tile_X4Y6_LUT4AB/FrameStrobe[10] Tile_X4Y6_LUT4AB/FrameStrobe[11]
+ Tile_X4Y6_LUT4AB/FrameStrobe[12] Tile_X4Y6_LUT4AB/FrameStrobe[13] Tile_X4Y6_LUT4AB/FrameStrobe[14]
+ Tile_X4Y6_LUT4AB/FrameStrobe[15] Tile_X4Y6_LUT4AB/FrameStrobe[16] Tile_X4Y6_LUT4AB/FrameStrobe[17]
+ Tile_X4Y6_LUT4AB/FrameStrobe[18] Tile_X4Y6_LUT4AB/FrameStrobe[19] Tile_X4Y6_LUT4AB/FrameStrobe[1]
+ Tile_X4Y6_LUT4AB/FrameStrobe[2] Tile_X4Y6_LUT4AB/FrameStrobe[3] Tile_X4Y6_LUT4AB/FrameStrobe[4]
+ Tile_X4Y6_LUT4AB/FrameStrobe[5] Tile_X4Y6_LUT4AB/FrameStrobe[6] Tile_X4Y6_LUT4AB/FrameStrobe[7]
+ Tile_X4Y6_LUT4AB/FrameStrobe[8] Tile_X4Y6_LUT4AB/FrameStrobe[9] Tile_X4Y7_LUT4AB/N1BEG[0]
+ Tile_X4Y7_LUT4AB/N1BEG[1] Tile_X4Y7_LUT4AB/N1BEG[2] Tile_X4Y7_LUT4AB/N1BEG[3] Tile_X4Y8_LUT4AB/N1BEG[0]
+ Tile_X4Y8_LUT4AB/N1BEG[1] Tile_X4Y8_LUT4AB/N1BEG[2] Tile_X4Y8_LUT4AB/N1BEG[3] Tile_X4Y7_LUT4AB/N2BEG[0]
+ Tile_X4Y7_LUT4AB/N2BEG[1] Tile_X4Y7_LUT4AB/N2BEG[2] Tile_X4Y7_LUT4AB/N2BEG[3] Tile_X4Y7_LUT4AB/N2BEG[4]
+ Tile_X4Y7_LUT4AB/N2BEG[5] Tile_X4Y7_LUT4AB/N2BEG[6] Tile_X4Y7_LUT4AB/N2BEG[7] Tile_X4Y6_LUT4AB/N2END[0]
+ Tile_X4Y6_LUT4AB/N2END[1] Tile_X4Y6_LUT4AB/N2END[2] Tile_X4Y6_LUT4AB/N2END[3] Tile_X4Y6_LUT4AB/N2END[4]
+ Tile_X4Y6_LUT4AB/N2END[5] Tile_X4Y6_LUT4AB/N2END[6] Tile_X4Y6_LUT4AB/N2END[7] Tile_X4Y7_LUT4AB/N2END[0]
+ Tile_X4Y7_LUT4AB/N2END[1] Tile_X4Y7_LUT4AB/N2END[2] Tile_X4Y7_LUT4AB/N2END[3] Tile_X4Y7_LUT4AB/N2END[4]
+ Tile_X4Y7_LUT4AB/N2END[5] Tile_X4Y7_LUT4AB/N2END[6] Tile_X4Y7_LUT4AB/N2END[7] Tile_X4Y8_LUT4AB/N2BEG[0]
+ Tile_X4Y8_LUT4AB/N2BEG[1] Tile_X4Y8_LUT4AB/N2BEG[2] Tile_X4Y8_LUT4AB/N2BEG[3] Tile_X4Y8_LUT4AB/N2BEG[4]
+ Tile_X4Y8_LUT4AB/N2BEG[5] Tile_X4Y8_LUT4AB/N2BEG[6] Tile_X4Y8_LUT4AB/N2BEG[7] Tile_X4Y7_LUT4AB/N4BEG[0]
+ Tile_X4Y7_LUT4AB/N4BEG[10] Tile_X4Y7_LUT4AB/N4BEG[11] Tile_X4Y7_LUT4AB/N4BEG[12]
+ Tile_X4Y7_LUT4AB/N4BEG[13] Tile_X4Y7_LUT4AB/N4BEG[14] Tile_X4Y7_LUT4AB/N4BEG[15]
+ Tile_X4Y7_LUT4AB/N4BEG[1] Tile_X4Y7_LUT4AB/N4BEG[2] Tile_X4Y7_LUT4AB/N4BEG[3] Tile_X4Y7_LUT4AB/N4BEG[4]
+ Tile_X4Y7_LUT4AB/N4BEG[5] Tile_X4Y7_LUT4AB/N4BEG[6] Tile_X4Y7_LUT4AB/N4BEG[7] Tile_X4Y7_LUT4AB/N4BEG[8]
+ Tile_X4Y7_LUT4AB/N4BEG[9] Tile_X4Y8_LUT4AB/N4BEG[0] Tile_X4Y8_LUT4AB/N4BEG[10] Tile_X4Y8_LUT4AB/N4BEG[11]
+ Tile_X4Y8_LUT4AB/N4BEG[12] Tile_X4Y8_LUT4AB/N4BEG[13] Tile_X4Y8_LUT4AB/N4BEG[14]
+ Tile_X4Y8_LUT4AB/N4BEG[15] Tile_X4Y8_LUT4AB/N4BEG[1] Tile_X4Y8_LUT4AB/N4BEG[2] Tile_X4Y8_LUT4AB/N4BEG[3]
+ Tile_X4Y8_LUT4AB/N4BEG[4] Tile_X4Y8_LUT4AB/N4BEG[5] Tile_X4Y8_LUT4AB/N4BEG[6] Tile_X4Y8_LUT4AB/N4BEG[7]
+ Tile_X4Y8_LUT4AB/N4BEG[8] Tile_X4Y8_LUT4AB/N4BEG[9] Tile_X4Y7_LUT4AB/NN4BEG[0] Tile_X4Y7_LUT4AB/NN4BEG[10]
+ Tile_X4Y7_LUT4AB/NN4BEG[11] Tile_X4Y7_LUT4AB/NN4BEG[12] Tile_X4Y7_LUT4AB/NN4BEG[13]
+ Tile_X4Y7_LUT4AB/NN4BEG[14] Tile_X4Y7_LUT4AB/NN4BEG[15] Tile_X4Y7_LUT4AB/NN4BEG[1]
+ Tile_X4Y7_LUT4AB/NN4BEG[2] Tile_X4Y7_LUT4AB/NN4BEG[3] Tile_X4Y7_LUT4AB/NN4BEG[4]
+ Tile_X4Y7_LUT4AB/NN4BEG[5] Tile_X4Y7_LUT4AB/NN4BEG[6] Tile_X4Y7_LUT4AB/NN4BEG[7]
+ Tile_X4Y7_LUT4AB/NN4BEG[8] Tile_X4Y7_LUT4AB/NN4BEG[9] Tile_X4Y8_LUT4AB/NN4BEG[0]
+ Tile_X4Y8_LUT4AB/NN4BEG[10] Tile_X4Y8_LUT4AB/NN4BEG[11] Tile_X4Y8_LUT4AB/NN4BEG[12]
+ Tile_X4Y8_LUT4AB/NN4BEG[13] Tile_X4Y8_LUT4AB/NN4BEG[14] Tile_X4Y8_LUT4AB/NN4BEG[15]
+ Tile_X4Y8_LUT4AB/NN4BEG[1] Tile_X4Y8_LUT4AB/NN4BEG[2] Tile_X4Y8_LUT4AB/NN4BEG[3]
+ Tile_X4Y8_LUT4AB/NN4BEG[4] Tile_X4Y8_LUT4AB/NN4BEG[5] Tile_X4Y8_LUT4AB/NN4BEG[6]
+ Tile_X4Y8_LUT4AB/NN4BEG[7] Tile_X4Y8_LUT4AB/NN4BEG[8] Tile_X4Y8_LUT4AB/NN4BEG[9]
+ Tile_X4Y8_LUT4AB/S1END[0] Tile_X4Y8_LUT4AB/S1END[1] Tile_X4Y8_LUT4AB/S1END[2] Tile_X4Y8_LUT4AB/S1END[3]
+ Tile_X4Y7_LUT4AB/S1END[0] Tile_X4Y7_LUT4AB/S1END[1] Tile_X4Y7_LUT4AB/S1END[2] Tile_X4Y7_LUT4AB/S1END[3]
+ Tile_X4Y8_LUT4AB/S2MID[0] Tile_X4Y8_LUT4AB/S2MID[1] Tile_X4Y8_LUT4AB/S2MID[2] Tile_X4Y8_LUT4AB/S2MID[3]
+ Tile_X4Y8_LUT4AB/S2MID[4] Tile_X4Y8_LUT4AB/S2MID[5] Tile_X4Y8_LUT4AB/S2MID[6] Tile_X4Y8_LUT4AB/S2MID[7]
+ Tile_X4Y8_LUT4AB/S2END[0] Tile_X4Y8_LUT4AB/S2END[1] Tile_X4Y8_LUT4AB/S2END[2] Tile_X4Y8_LUT4AB/S2END[3]
+ Tile_X4Y8_LUT4AB/S2END[4] Tile_X4Y8_LUT4AB/S2END[5] Tile_X4Y8_LUT4AB/S2END[6] Tile_X4Y8_LUT4AB/S2END[7]
+ Tile_X4Y7_LUT4AB/S2END[0] Tile_X4Y7_LUT4AB/S2END[1] Tile_X4Y7_LUT4AB/S2END[2] Tile_X4Y7_LUT4AB/S2END[3]
+ Tile_X4Y7_LUT4AB/S2END[4] Tile_X4Y7_LUT4AB/S2END[5] Tile_X4Y7_LUT4AB/S2END[6] Tile_X4Y7_LUT4AB/S2END[7]
+ Tile_X4Y7_LUT4AB/S2MID[0] Tile_X4Y7_LUT4AB/S2MID[1] Tile_X4Y7_LUT4AB/S2MID[2] Tile_X4Y7_LUT4AB/S2MID[3]
+ Tile_X4Y7_LUT4AB/S2MID[4] Tile_X4Y7_LUT4AB/S2MID[5] Tile_X4Y7_LUT4AB/S2MID[6] Tile_X4Y7_LUT4AB/S2MID[7]
+ Tile_X4Y8_LUT4AB/S4END[0] Tile_X4Y8_LUT4AB/S4END[10] Tile_X4Y8_LUT4AB/S4END[11]
+ Tile_X4Y8_LUT4AB/S4END[12] Tile_X4Y8_LUT4AB/S4END[13] Tile_X4Y8_LUT4AB/S4END[14]
+ Tile_X4Y8_LUT4AB/S4END[15] Tile_X4Y8_LUT4AB/S4END[1] Tile_X4Y8_LUT4AB/S4END[2] Tile_X4Y8_LUT4AB/S4END[3]
+ Tile_X4Y8_LUT4AB/S4END[4] Tile_X4Y8_LUT4AB/S4END[5] Tile_X4Y8_LUT4AB/S4END[6] Tile_X4Y8_LUT4AB/S4END[7]
+ Tile_X4Y8_LUT4AB/S4END[8] Tile_X4Y8_LUT4AB/S4END[9] Tile_X4Y7_LUT4AB/S4END[0] Tile_X4Y7_LUT4AB/S4END[10]
+ Tile_X4Y7_LUT4AB/S4END[11] Tile_X4Y7_LUT4AB/S4END[12] Tile_X4Y7_LUT4AB/S4END[13]
+ Tile_X4Y7_LUT4AB/S4END[14] Tile_X4Y7_LUT4AB/S4END[15] Tile_X4Y7_LUT4AB/S4END[1]
+ Tile_X4Y7_LUT4AB/S4END[2] Tile_X4Y7_LUT4AB/S4END[3] Tile_X4Y7_LUT4AB/S4END[4] Tile_X4Y7_LUT4AB/S4END[5]
+ Tile_X4Y7_LUT4AB/S4END[6] Tile_X4Y7_LUT4AB/S4END[7] Tile_X4Y7_LUT4AB/S4END[8] Tile_X4Y7_LUT4AB/S4END[9]
+ Tile_X4Y8_LUT4AB/SS4END[0] Tile_X4Y8_LUT4AB/SS4END[10] Tile_X4Y8_LUT4AB/SS4END[11]
+ Tile_X4Y8_LUT4AB/SS4END[12] Tile_X4Y8_LUT4AB/SS4END[13] Tile_X4Y8_LUT4AB/SS4END[14]
+ Tile_X4Y8_LUT4AB/SS4END[15] Tile_X4Y8_LUT4AB/SS4END[1] Tile_X4Y8_LUT4AB/SS4END[2]
+ Tile_X4Y8_LUT4AB/SS4END[3] Tile_X4Y8_LUT4AB/SS4END[4] Tile_X4Y8_LUT4AB/SS4END[5]
+ Tile_X4Y8_LUT4AB/SS4END[6] Tile_X4Y8_LUT4AB/SS4END[7] Tile_X4Y8_LUT4AB/SS4END[8]
+ Tile_X4Y8_LUT4AB/SS4END[9] Tile_X4Y7_LUT4AB/SS4END[0] Tile_X4Y7_LUT4AB/SS4END[10]
+ Tile_X4Y7_LUT4AB/SS4END[11] Tile_X4Y7_LUT4AB/SS4END[12] Tile_X4Y7_LUT4AB/SS4END[13]
+ Tile_X4Y7_LUT4AB/SS4END[14] Tile_X4Y7_LUT4AB/SS4END[15] Tile_X4Y7_LUT4AB/SS4END[1]
+ Tile_X4Y7_LUT4AB/SS4END[2] Tile_X4Y7_LUT4AB/SS4END[3] Tile_X4Y7_LUT4AB/SS4END[4]
+ Tile_X4Y7_LUT4AB/SS4END[5] Tile_X4Y7_LUT4AB/SS4END[6] Tile_X4Y7_LUT4AB/SS4END[7]
+ Tile_X4Y7_LUT4AB/SS4END[8] Tile_X4Y7_LUT4AB/SS4END[9] Tile_X4Y7_LUT4AB/UserCLK Tile_X4Y6_LUT4AB/UserCLK
+ VGND VPWR Tile_X4Y7_LUT4AB/W1BEG[0] Tile_X4Y7_LUT4AB/W1BEG[1] Tile_X4Y7_LUT4AB/W1BEG[2]
+ Tile_X4Y7_LUT4AB/W1BEG[3] Tile_X4Y7_LUT4AB/W1END[0] Tile_X4Y7_LUT4AB/W1END[1] Tile_X4Y7_LUT4AB/W1END[2]
+ Tile_X4Y7_LUT4AB/W1END[3] Tile_X4Y7_LUT4AB/W2BEG[0] Tile_X4Y7_LUT4AB/W2BEG[1] Tile_X4Y7_LUT4AB/W2BEG[2]
+ Tile_X4Y7_LUT4AB/W2BEG[3] Tile_X4Y7_LUT4AB/W2BEG[4] Tile_X4Y7_LUT4AB/W2BEG[5] Tile_X4Y7_LUT4AB/W2BEG[6]
+ Tile_X4Y7_LUT4AB/W2BEG[7] Tile_X3Y7_LUT4AB/W2END[0] Tile_X3Y7_LUT4AB/W2END[1] Tile_X3Y7_LUT4AB/W2END[2]
+ Tile_X3Y7_LUT4AB/W2END[3] Tile_X3Y7_LUT4AB/W2END[4] Tile_X3Y7_LUT4AB/W2END[5] Tile_X3Y7_LUT4AB/W2END[6]
+ Tile_X3Y7_LUT4AB/W2END[7] Tile_X4Y7_LUT4AB/W2END[0] Tile_X4Y7_LUT4AB/W2END[1] Tile_X4Y7_LUT4AB/W2END[2]
+ Tile_X4Y7_LUT4AB/W2END[3] Tile_X4Y7_LUT4AB/W2END[4] Tile_X4Y7_LUT4AB/W2END[5] Tile_X4Y7_LUT4AB/W2END[6]
+ Tile_X4Y7_LUT4AB/W2END[7] Tile_X4Y7_LUT4AB/W2MID[0] Tile_X4Y7_LUT4AB/W2MID[1] Tile_X4Y7_LUT4AB/W2MID[2]
+ Tile_X4Y7_LUT4AB/W2MID[3] Tile_X4Y7_LUT4AB/W2MID[4] Tile_X4Y7_LUT4AB/W2MID[5] Tile_X4Y7_LUT4AB/W2MID[6]
+ Tile_X4Y7_LUT4AB/W2MID[7] Tile_X4Y7_LUT4AB/W6BEG[0] Tile_X4Y7_LUT4AB/W6BEG[10] Tile_X4Y7_LUT4AB/W6BEG[11]
+ Tile_X4Y7_LUT4AB/W6BEG[1] Tile_X4Y7_LUT4AB/W6BEG[2] Tile_X4Y7_LUT4AB/W6BEG[3] Tile_X4Y7_LUT4AB/W6BEG[4]
+ Tile_X4Y7_LUT4AB/W6BEG[5] Tile_X4Y7_LUT4AB/W6BEG[6] Tile_X4Y7_LUT4AB/W6BEG[7] Tile_X4Y7_LUT4AB/W6BEG[8]
+ Tile_X4Y7_LUT4AB/W6BEG[9] Tile_X4Y7_LUT4AB/W6END[0] Tile_X4Y7_LUT4AB/W6END[10] Tile_X4Y7_LUT4AB/W6END[11]
+ Tile_X4Y7_LUT4AB/W6END[1] Tile_X4Y7_LUT4AB/W6END[2] Tile_X4Y7_LUT4AB/W6END[3] Tile_X4Y7_LUT4AB/W6END[4]
+ Tile_X4Y7_LUT4AB/W6END[5] Tile_X4Y7_LUT4AB/W6END[6] Tile_X4Y7_LUT4AB/W6END[7] Tile_X4Y7_LUT4AB/W6END[8]
+ Tile_X4Y7_LUT4AB/W6END[9] Tile_X4Y7_LUT4AB/WW4BEG[0] Tile_X4Y7_LUT4AB/WW4BEG[10]
+ Tile_X4Y7_LUT4AB/WW4BEG[11] Tile_X4Y7_LUT4AB/WW4BEG[12] Tile_X4Y7_LUT4AB/WW4BEG[13]
+ Tile_X4Y7_LUT4AB/WW4BEG[14] Tile_X4Y7_LUT4AB/WW4BEG[15] Tile_X4Y7_LUT4AB/WW4BEG[1]
+ Tile_X4Y7_LUT4AB/WW4BEG[2] Tile_X4Y7_LUT4AB/WW4BEG[3] Tile_X4Y7_LUT4AB/WW4BEG[4]
+ Tile_X4Y7_LUT4AB/WW4BEG[5] Tile_X4Y7_LUT4AB/WW4BEG[6] Tile_X4Y7_LUT4AB/WW4BEG[7]
+ Tile_X4Y7_LUT4AB/WW4BEG[8] Tile_X4Y7_LUT4AB/WW4BEG[9] Tile_X4Y7_LUT4AB/WW4END[0]
+ Tile_X4Y7_LUT4AB/WW4END[10] Tile_X4Y7_LUT4AB/WW4END[11] Tile_X4Y7_LUT4AB/WW4END[12]
+ Tile_X4Y7_LUT4AB/WW4END[13] Tile_X4Y7_LUT4AB/WW4END[14] Tile_X4Y7_LUT4AB/WW4END[15]
+ Tile_X4Y7_LUT4AB/WW4END[1] Tile_X4Y7_LUT4AB/WW4END[2] Tile_X4Y7_LUT4AB/WW4END[3]
+ Tile_X4Y7_LUT4AB/WW4END[4] Tile_X4Y7_LUT4AB/WW4END[5] Tile_X4Y7_LUT4AB/WW4END[6]
+ Tile_X4Y7_LUT4AB/WW4END[7] Tile_X4Y7_LUT4AB/WW4END[8] Tile_X4Y7_LUT4AB/WW4END[9]
+ LUT4AB
XTile_X5Y6_E_TT_IF Tile_X5Y6_CLK_TT_PROJECT Tile_X4Y6_LUT4AB/E1BEG[0] Tile_X4Y6_LUT4AB/E1BEG[1]
+ Tile_X4Y6_LUT4AB/E1BEG[2] Tile_X4Y6_LUT4AB/E1BEG[3] Tile_X5Y6_E_TT_IF/E2END[0] Tile_X5Y6_E_TT_IF/E2END[1]
+ Tile_X5Y6_E_TT_IF/E2END[2] Tile_X5Y6_E_TT_IF/E2END[3] Tile_X5Y6_E_TT_IF/E2END[4]
+ Tile_X5Y6_E_TT_IF/E2END[5] Tile_X5Y6_E_TT_IF/E2END[6] Tile_X5Y6_E_TT_IF/E2END[7]
+ Tile_X4Y6_LUT4AB/E2BEG[0] Tile_X4Y6_LUT4AB/E2BEG[1] Tile_X4Y6_LUT4AB/E2BEG[2] Tile_X4Y6_LUT4AB/E2BEG[3]
+ Tile_X4Y6_LUT4AB/E2BEG[4] Tile_X4Y6_LUT4AB/E2BEG[5] Tile_X4Y6_LUT4AB/E2BEG[6] Tile_X4Y6_LUT4AB/E2BEG[7]
+ Tile_X4Y6_LUT4AB/E6BEG[0] Tile_X4Y6_LUT4AB/E6BEG[10] Tile_X4Y6_LUT4AB/E6BEG[11]
+ Tile_X4Y6_LUT4AB/E6BEG[1] Tile_X4Y6_LUT4AB/E6BEG[2] Tile_X4Y6_LUT4AB/E6BEG[3] Tile_X4Y6_LUT4AB/E6BEG[4]
+ Tile_X4Y6_LUT4AB/E6BEG[5] Tile_X4Y6_LUT4AB/E6BEG[6] Tile_X4Y6_LUT4AB/E6BEG[7] Tile_X4Y6_LUT4AB/E6BEG[8]
+ Tile_X4Y6_LUT4AB/E6BEG[9] Tile_X4Y6_LUT4AB/EE4BEG[0] Tile_X4Y6_LUT4AB/EE4BEG[10]
+ Tile_X4Y6_LUT4AB/EE4BEG[11] Tile_X4Y6_LUT4AB/EE4BEG[12] Tile_X4Y6_LUT4AB/EE4BEG[13]
+ Tile_X4Y6_LUT4AB/EE4BEG[14] Tile_X4Y6_LUT4AB/EE4BEG[15] Tile_X4Y6_LUT4AB/EE4BEG[1]
+ Tile_X4Y6_LUT4AB/EE4BEG[2] Tile_X4Y6_LUT4AB/EE4BEG[3] Tile_X4Y6_LUT4AB/EE4BEG[4]
+ Tile_X4Y6_LUT4AB/EE4BEG[5] Tile_X4Y6_LUT4AB/EE4BEG[6] Tile_X4Y6_LUT4AB/EE4BEG[7]
+ Tile_X4Y6_LUT4AB/EE4BEG[8] Tile_X4Y6_LUT4AB/EE4BEG[9] Tile_X5Y6_ENA_TT_PROJECT Tile_X5Y6_E_TT_IF/FrameData[0]
+ Tile_X5Y6_E_TT_IF/FrameData[10] Tile_X5Y6_E_TT_IF/FrameData[11] Tile_X5Y6_E_TT_IF/FrameData[12]
+ Tile_X5Y6_E_TT_IF/FrameData[13] Tile_X5Y6_E_TT_IF/FrameData[14] Tile_X5Y6_E_TT_IF/FrameData[15]
+ Tile_X5Y6_E_TT_IF/FrameData[16] Tile_X5Y6_E_TT_IF/FrameData[17] Tile_X5Y6_E_TT_IF/FrameData[18]
+ Tile_X5Y6_E_TT_IF/FrameData[19] Tile_X5Y6_E_TT_IF/FrameData[1] Tile_X5Y6_E_TT_IF/FrameData[20]
+ Tile_X5Y6_E_TT_IF/FrameData[21] Tile_X5Y6_E_TT_IF/FrameData[22] Tile_X5Y6_E_TT_IF/FrameData[23]
+ Tile_X5Y6_E_TT_IF/FrameData[24] Tile_X5Y6_E_TT_IF/FrameData[25] Tile_X5Y6_E_TT_IF/FrameData[26]
+ Tile_X5Y6_E_TT_IF/FrameData[27] Tile_X5Y6_E_TT_IF/FrameData[28] Tile_X5Y6_E_TT_IF/FrameData[29]
+ Tile_X5Y6_E_TT_IF/FrameData[2] Tile_X5Y6_E_TT_IF/FrameData[30] Tile_X5Y6_E_TT_IF/FrameData[31]
+ Tile_X5Y6_E_TT_IF/FrameData[3] Tile_X5Y6_E_TT_IF/FrameData[4] Tile_X5Y6_E_TT_IF/FrameData[5]
+ Tile_X5Y6_E_TT_IF/FrameData[6] Tile_X5Y6_E_TT_IF/FrameData[7] Tile_X5Y6_E_TT_IF/FrameData[8]
+ Tile_X5Y6_E_TT_IF/FrameData[9] Tile_X5Y6_E_TT_IF/FrameData_O[0] Tile_X5Y6_E_TT_IF/FrameData_O[10]
+ Tile_X5Y6_E_TT_IF/FrameData_O[11] Tile_X5Y6_E_TT_IF/FrameData_O[12] Tile_X5Y6_E_TT_IF/FrameData_O[13]
+ Tile_X5Y6_E_TT_IF/FrameData_O[14] Tile_X5Y6_E_TT_IF/FrameData_O[15] Tile_X5Y6_E_TT_IF/FrameData_O[16]
+ Tile_X5Y6_E_TT_IF/FrameData_O[17] Tile_X5Y6_E_TT_IF/FrameData_O[18] Tile_X5Y6_E_TT_IF/FrameData_O[19]
+ Tile_X5Y6_E_TT_IF/FrameData_O[1] Tile_X5Y6_E_TT_IF/FrameData_O[20] Tile_X5Y6_E_TT_IF/FrameData_O[21]
+ Tile_X5Y6_E_TT_IF/FrameData_O[22] Tile_X5Y6_E_TT_IF/FrameData_O[23] Tile_X5Y6_E_TT_IF/FrameData_O[24]
+ Tile_X5Y6_E_TT_IF/FrameData_O[25] Tile_X5Y6_E_TT_IF/FrameData_O[26] Tile_X5Y6_E_TT_IF/FrameData_O[27]
+ Tile_X5Y6_E_TT_IF/FrameData_O[28] Tile_X5Y6_E_TT_IF/FrameData_O[29] Tile_X5Y6_E_TT_IF/FrameData_O[2]
+ Tile_X5Y6_E_TT_IF/FrameData_O[30] Tile_X5Y6_E_TT_IF/FrameData_O[31] Tile_X5Y6_E_TT_IF/FrameData_O[3]
+ Tile_X5Y6_E_TT_IF/FrameData_O[4] Tile_X5Y6_E_TT_IF/FrameData_O[5] Tile_X5Y6_E_TT_IF/FrameData_O[6]
+ Tile_X5Y6_E_TT_IF/FrameData_O[7] Tile_X5Y6_E_TT_IF/FrameData_O[8] Tile_X5Y6_E_TT_IF/FrameData_O[9]
+ Tile_X5Y6_E_TT_IF/FrameStrobe[0] Tile_X5Y6_E_TT_IF/FrameStrobe[10] Tile_X5Y6_E_TT_IF/FrameStrobe[11]
+ Tile_X5Y6_E_TT_IF/FrameStrobe[12] Tile_X5Y6_E_TT_IF/FrameStrobe[13] Tile_X5Y6_E_TT_IF/FrameStrobe[14]
+ Tile_X5Y6_E_TT_IF/FrameStrobe[15] Tile_X5Y6_E_TT_IF/FrameStrobe[16] Tile_X5Y6_E_TT_IF/FrameStrobe[17]
+ Tile_X5Y6_E_TT_IF/FrameStrobe[18] Tile_X5Y6_E_TT_IF/FrameStrobe[19] Tile_X5Y6_E_TT_IF/FrameStrobe[1]
+ Tile_X5Y6_E_TT_IF/FrameStrobe[2] Tile_X5Y6_E_TT_IF/FrameStrobe[3] Tile_X5Y6_E_TT_IF/FrameStrobe[4]
+ Tile_X5Y6_E_TT_IF/FrameStrobe[5] Tile_X5Y6_E_TT_IF/FrameStrobe[6] Tile_X5Y6_E_TT_IF/FrameStrobe[7]
+ Tile_X5Y6_E_TT_IF/FrameStrobe[8] Tile_X5Y6_E_TT_IF/FrameStrobe[9] Tile_X5Y5_E_TT_IF/FrameStrobe[0]
+ Tile_X5Y5_E_TT_IF/FrameStrobe[10] Tile_X5Y5_E_TT_IF/FrameStrobe[11] Tile_X5Y5_E_TT_IF/FrameStrobe[12]
+ Tile_X5Y5_E_TT_IF/FrameStrobe[13] Tile_X5Y5_E_TT_IF/FrameStrobe[14] Tile_X5Y5_E_TT_IF/FrameStrobe[15]
+ Tile_X5Y5_E_TT_IF/FrameStrobe[16] Tile_X5Y5_E_TT_IF/FrameStrobe[17] Tile_X5Y5_E_TT_IF/FrameStrobe[18]
+ Tile_X5Y5_E_TT_IF/FrameStrobe[19] Tile_X5Y5_E_TT_IF/FrameStrobe[1] Tile_X5Y5_E_TT_IF/FrameStrobe[2]
+ Tile_X5Y5_E_TT_IF/FrameStrobe[3] Tile_X5Y5_E_TT_IF/FrameStrobe[4] Tile_X5Y5_E_TT_IF/FrameStrobe[5]
+ Tile_X5Y5_E_TT_IF/FrameStrobe[6] Tile_X5Y5_E_TT_IF/FrameStrobe[7] Tile_X5Y5_E_TT_IF/FrameStrobe[8]
+ Tile_X5Y5_E_TT_IF/FrameStrobe[9] Tile_X5Y6_E_TT_IF/N1BEG[0] Tile_X5Y6_E_TT_IF/N1BEG[1]
+ Tile_X5Y6_E_TT_IF/N1BEG[2] Tile_X5Y6_E_TT_IF/N1BEG[3] Tile_X5Y7_E_TT_IF/N1BEG[0]
+ Tile_X5Y7_E_TT_IF/N1BEG[1] Tile_X5Y7_E_TT_IF/N1BEG[2] Tile_X5Y7_E_TT_IF/N1BEG[3]
+ Tile_X5Y6_E_TT_IF/N2BEG[0] Tile_X5Y6_E_TT_IF/N2BEG[1] Tile_X5Y6_E_TT_IF/N2BEG[2]
+ Tile_X5Y6_E_TT_IF/N2BEG[3] Tile_X5Y6_E_TT_IF/N2BEG[4] Tile_X5Y6_E_TT_IF/N2BEG[5]
+ Tile_X5Y6_E_TT_IF/N2BEG[6] Tile_X5Y6_E_TT_IF/N2BEG[7] Tile_X5Y5_E_TT_IF/N2END[0]
+ Tile_X5Y5_E_TT_IF/N2END[1] Tile_X5Y5_E_TT_IF/N2END[2] Tile_X5Y5_E_TT_IF/N2END[3]
+ Tile_X5Y5_E_TT_IF/N2END[4] Tile_X5Y5_E_TT_IF/N2END[5] Tile_X5Y5_E_TT_IF/N2END[6]
+ Tile_X5Y5_E_TT_IF/N2END[7] Tile_X5Y6_E_TT_IF/N2END[0] Tile_X5Y6_E_TT_IF/N2END[1]
+ Tile_X5Y6_E_TT_IF/N2END[2] Tile_X5Y6_E_TT_IF/N2END[3] Tile_X5Y6_E_TT_IF/N2END[4]
+ Tile_X5Y6_E_TT_IF/N2END[5] Tile_X5Y6_E_TT_IF/N2END[6] Tile_X5Y6_E_TT_IF/N2END[7]
+ Tile_X5Y7_E_TT_IF/N2BEG[0] Tile_X5Y7_E_TT_IF/N2BEG[1] Tile_X5Y7_E_TT_IF/N2BEG[2]
+ Tile_X5Y7_E_TT_IF/N2BEG[3] Tile_X5Y7_E_TT_IF/N2BEG[4] Tile_X5Y7_E_TT_IF/N2BEG[5]
+ Tile_X5Y7_E_TT_IF/N2BEG[6] Tile_X5Y7_E_TT_IF/N2BEG[7] Tile_X5Y6_E_TT_IF/N4BEG[0]
+ Tile_X5Y6_E_TT_IF/N4BEG[10] Tile_X5Y6_E_TT_IF/N4BEG[11] Tile_X5Y6_E_TT_IF/N4BEG[12]
+ Tile_X5Y6_E_TT_IF/N4BEG[13] Tile_X5Y6_E_TT_IF/N4BEG[14] Tile_X5Y6_E_TT_IF/N4BEG[15]
+ Tile_X5Y6_E_TT_IF/N4BEG[1] Tile_X5Y6_E_TT_IF/N4BEG[2] Tile_X5Y6_E_TT_IF/N4BEG[3]
+ Tile_X5Y6_E_TT_IF/N4BEG[4] Tile_X5Y6_E_TT_IF/N4BEG[5] Tile_X5Y6_E_TT_IF/N4BEG[6]
+ Tile_X5Y6_E_TT_IF/N4BEG[7] Tile_X5Y6_E_TT_IF/N4BEG[8] Tile_X5Y6_E_TT_IF/N4BEG[9]
+ Tile_X5Y7_E_TT_IF/N4BEG[0] Tile_X5Y7_E_TT_IF/N4BEG[10] Tile_X5Y7_E_TT_IF/N4BEG[11]
+ Tile_X5Y7_E_TT_IF/N4BEG[12] Tile_X5Y7_E_TT_IF/N4BEG[13] Tile_X5Y7_E_TT_IF/N4BEG[14]
+ Tile_X5Y7_E_TT_IF/N4BEG[15] Tile_X5Y7_E_TT_IF/N4BEG[1] Tile_X5Y7_E_TT_IF/N4BEG[2]
+ Tile_X5Y7_E_TT_IF/N4BEG[3] Tile_X5Y7_E_TT_IF/N4BEG[4] Tile_X5Y7_E_TT_IF/N4BEG[5]
+ Tile_X5Y7_E_TT_IF/N4BEG[6] Tile_X5Y7_E_TT_IF/N4BEG[7] Tile_X5Y7_E_TT_IF/N4BEG[8]
+ Tile_X5Y7_E_TT_IF/N4BEG[9] Tile_X5Y6_RST_N_TT_PROJECT Tile_X5Y7_E_TT_IF/S1END[0]
+ Tile_X5Y7_E_TT_IF/S1END[1] Tile_X5Y7_E_TT_IF/S1END[2] Tile_X5Y7_E_TT_IF/S1END[3]
+ Tile_X5Y6_E_TT_IF/S1END[0] Tile_X5Y6_E_TT_IF/S1END[1] Tile_X5Y6_E_TT_IF/S1END[2]
+ Tile_X5Y6_E_TT_IF/S1END[3] Tile_X5Y7_E_TT_IF/S2MID[0] Tile_X5Y7_E_TT_IF/S2MID[1]
+ Tile_X5Y7_E_TT_IF/S2MID[2] Tile_X5Y7_E_TT_IF/S2MID[3] Tile_X5Y7_E_TT_IF/S2MID[4]
+ Tile_X5Y7_E_TT_IF/S2MID[5] Tile_X5Y7_E_TT_IF/S2MID[6] Tile_X5Y7_E_TT_IF/S2MID[7]
+ Tile_X5Y7_E_TT_IF/S2END[0] Tile_X5Y7_E_TT_IF/S2END[1] Tile_X5Y7_E_TT_IF/S2END[2]
+ Tile_X5Y7_E_TT_IF/S2END[3] Tile_X5Y7_E_TT_IF/S2END[4] Tile_X5Y7_E_TT_IF/S2END[5]
+ Tile_X5Y7_E_TT_IF/S2END[6] Tile_X5Y7_E_TT_IF/S2END[7] Tile_X5Y6_E_TT_IF/S2END[0]
+ Tile_X5Y6_E_TT_IF/S2END[1] Tile_X5Y6_E_TT_IF/S2END[2] Tile_X5Y6_E_TT_IF/S2END[3]
+ Tile_X5Y6_E_TT_IF/S2END[4] Tile_X5Y6_E_TT_IF/S2END[5] Tile_X5Y6_E_TT_IF/S2END[6]
+ Tile_X5Y6_E_TT_IF/S2END[7] Tile_X5Y6_E_TT_IF/S2MID[0] Tile_X5Y6_E_TT_IF/S2MID[1]
+ Tile_X5Y6_E_TT_IF/S2MID[2] Tile_X5Y6_E_TT_IF/S2MID[3] Tile_X5Y6_E_TT_IF/S2MID[4]
+ Tile_X5Y6_E_TT_IF/S2MID[5] Tile_X5Y6_E_TT_IF/S2MID[6] Tile_X5Y6_E_TT_IF/S2MID[7]
+ Tile_X5Y7_E_TT_IF/S4END[0] Tile_X5Y7_E_TT_IF/S4END[10] Tile_X5Y7_E_TT_IF/S4END[11]
+ Tile_X5Y7_E_TT_IF/S4END[12] Tile_X5Y7_E_TT_IF/S4END[13] Tile_X5Y7_E_TT_IF/S4END[14]
+ Tile_X5Y7_E_TT_IF/S4END[15] Tile_X5Y7_E_TT_IF/S4END[1] Tile_X5Y7_E_TT_IF/S4END[2]
+ Tile_X5Y7_E_TT_IF/S4END[3] Tile_X5Y7_E_TT_IF/S4END[4] Tile_X5Y7_E_TT_IF/S4END[5]
+ Tile_X5Y7_E_TT_IF/S4END[6] Tile_X5Y7_E_TT_IF/S4END[7] Tile_X5Y7_E_TT_IF/S4END[8]
+ Tile_X5Y7_E_TT_IF/S4END[9] Tile_X5Y6_E_TT_IF/S4END[0] Tile_X5Y6_E_TT_IF/S4END[10]
+ Tile_X5Y6_E_TT_IF/S4END[11] Tile_X5Y6_E_TT_IF/S4END[12] Tile_X5Y6_E_TT_IF/S4END[13]
+ Tile_X5Y6_E_TT_IF/S4END[14] Tile_X5Y6_E_TT_IF/S4END[15] Tile_X5Y6_E_TT_IF/S4END[1]
+ Tile_X5Y6_E_TT_IF/S4END[2] Tile_X5Y6_E_TT_IF/S4END[3] Tile_X5Y6_E_TT_IF/S4END[4]
+ Tile_X5Y6_E_TT_IF/S4END[5] Tile_X5Y6_E_TT_IF/S4END[6] Tile_X5Y6_E_TT_IF/S4END[7]
+ Tile_X5Y6_E_TT_IF/S4END[8] Tile_X5Y6_E_TT_IF/S4END[9] Tile_X5Y6_UIO_IN_TT_PROJECT0
+ Tile_X5Y6_UIO_IN_TT_PROJECT1 Tile_X5Y6_UIO_IN_TT_PROJECT2 Tile_X5Y6_UIO_IN_TT_PROJECT3
+ Tile_X5Y6_UIO_IN_TT_PROJECT4 Tile_X5Y6_UIO_IN_TT_PROJECT5 Tile_X5Y6_UIO_IN_TT_PROJECT6
+ Tile_X5Y6_UIO_IN_TT_PROJECT7 Tile_X5Y6_UIO_OE_TT_PROJECT0 Tile_X5Y6_UIO_OE_TT_PROJECT1
+ Tile_X5Y6_UIO_OE_TT_PROJECT2 Tile_X5Y6_UIO_OE_TT_PROJECT3 Tile_X5Y6_UIO_OE_TT_PROJECT4
+ Tile_X5Y6_UIO_OE_TT_PROJECT5 Tile_X5Y6_UIO_OE_TT_PROJECT6 Tile_X5Y6_UIO_OE_TT_PROJECT7
+ Tile_X5Y6_UIO_OUT_TT_PROJECT0 Tile_X5Y6_UIO_OUT_TT_PROJECT1 Tile_X5Y6_UIO_OUT_TT_PROJECT2
+ Tile_X5Y6_UIO_OUT_TT_PROJECT3 Tile_X5Y6_UIO_OUT_TT_PROJECT4 Tile_X5Y6_UIO_OUT_TT_PROJECT5
+ Tile_X5Y6_UIO_OUT_TT_PROJECT6 Tile_X5Y6_UIO_OUT_TT_PROJECT7 Tile_X5Y6_UI_IN_TT_PROJECT0
+ Tile_X5Y6_UI_IN_TT_PROJECT1 Tile_X5Y6_UI_IN_TT_PROJECT2 Tile_X5Y6_UI_IN_TT_PROJECT3
+ Tile_X5Y6_UI_IN_TT_PROJECT4 Tile_X5Y6_UI_IN_TT_PROJECT5 Tile_X5Y6_UI_IN_TT_PROJECT6
+ Tile_X5Y6_UI_IN_TT_PROJECT7 Tile_X5Y6_UO_OUT_TT_PROJECT0 Tile_X5Y6_UO_OUT_TT_PROJECT1
+ Tile_X5Y6_UO_OUT_TT_PROJECT2 Tile_X5Y6_UO_OUT_TT_PROJECT3 Tile_X5Y6_UO_OUT_TT_PROJECT4
+ Tile_X5Y6_UO_OUT_TT_PROJECT5 Tile_X5Y6_UO_OUT_TT_PROJECT6 Tile_X5Y6_UO_OUT_TT_PROJECT7
+ Tile_X5Y6_E_TT_IF/UserCLK Tile_X5Y5_E_TT_IF/UserCLK VGND VPWR Tile_X4Y6_LUT4AB/W1END[0]
+ Tile_X4Y6_LUT4AB/W1END[1] Tile_X4Y6_LUT4AB/W1END[2] Tile_X4Y6_LUT4AB/W1END[3] Tile_X4Y6_LUT4AB/W2MID[0]
+ Tile_X4Y6_LUT4AB/W2MID[1] Tile_X4Y6_LUT4AB/W2MID[2] Tile_X4Y6_LUT4AB/W2MID[3] Tile_X4Y6_LUT4AB/W2MID[4]
+ Tile_X4Y6_LUT4AB/W2MID[5] Tile_X4Y6_LUT4AB/W2MID[6] Tile_X4Y6_LUT4AB/W2MID[7] Tile_X4Y6_LUT4AB/W2END[0]
+ Tile_X4Y6_LUT4AB/W2END[1] Tile_X4Y6_LUT4AB/W2END[2] Tile_X4Y6_LUT4AB/W2END[3] Tile_X4Y6_LUT4AB/W2END[4]
+ Tile_X4Y6_LUT4AB/W2END[5] Tile_X4Y6_LUT4AB/W2END[6] Tile_X4Y6_LUT4AB/W2END[7] Tile_X4Y6_LUT4AB/W6END[0]
+ Tile_X4Y6_LUT4AB/W6END[10] Tile_X4Y6_LUT4AB/W6END[11] Tile_X4Y6_LUT4AB/W6END[1]
+ Tile_X4Y6_LUT4AB/W6END[2] Tile_X4Y6_LUT4AB/W6END[3] Tile_X4Y6_LUT4AB/W6END[4] Tile_X4Y6_LUT4AB/W6END[5]
+ Tile_X4Y6_LUT4AB/W6END[6] Tile_X4Y6_LUT4AB/W6END[7] Tile_X4Y6_LUT4AB/W6END[8] Tile_X4Y6_LUT4AB/W6END[9]
+ Tile_X4Y6_LUT4AB/WW4END[0] Tile_X4Y6_LUT4AB/WW4END[10] Tile_X4Y6_LUT4AB/WW4END[11]
+ Tile_X4Y6_LUT4AB/WW4END[12] Tile_X4Y6_LUT4AB/WW4END[13] Tile_X4Y6_LUT4AB/WW4END[14]
+ Tile_X4Y6_LUT4AB/WW4END[15] Tile_X4Y6_LUT4AB/WW4END[1] Tile_X4Y6_LUT4AB/WW4END[2]
+ Tile_X4Y6_LUT4AB/WW4END[3] Tile_X4Y6_LUT4AB/WW4END[4] Tile_X4Y6_LUT4AB/WW4END[5]
+ Tile_X4Y6_LUT4AB/WW4END[6] Tile_X4Y6_LUT4AB/WW4END[7] Tile_X4Y6_LUT4AB/WW4END[8]
+ Tile_X4Y6_LUT4AB/WW4END[9] E_TT_IF
XTile_X1Y0_N_IO4 Tile_X1Y0_A_I_top Tile_X1Y0_A_O_top Tile_X1Y0_A_T_top Tile_X1Y0_B_I_top
+ Tile_X1Y0_B_O_top Tile_X1Y0_B_T_top Tile_X1Y0_C_I_top Tile_X1Y0_C_O_top Tile_X1Y0_C_T_top
+ Tile_X1Y0_N_IO4/Ci Tile_X1Y0_D_I_top Tile_X1Y0_D_O_top Tile_X1Y0_D_T_top Tile_X1Y0_N_IO4/FrameData[0]
+ Tile_X1Y0_N_IO4/FrameData[10] Tile_X1Y0_N_IO4/FrameData[11] Tile_X1Y0_N_IO4/FrameData[12]
+ Tile_X1Y0_N_IO4/FrameData[13] Tile_X1Y0_N_IO4/FrameData[14] Tile_X1Y0_N_IO4/FrameData[15]
+ Tile_X1Y0_N_IO4/FrameData[16] Tile_X1Y0_N_IO4/FrameData[17] Tile_X1Y0_N_IO4/FrameData[18]
+ Tile_X1Y0_N_IO4/FrameData[19] Tile_X1Y0_N_IO4/FrameData[1] Tile_X1Y0_N_IO4/FrameData[20]
+ Tile_X1Y0_N_IO4/FrameData[21] Tile_X1Y0_N_IO4/FrameData[22] Tile_X1Y0_N_IO4/FrameData[23]
+ Tile_X1Y0_N_IO4/FrameData[24] Tile_X1Y0_N_IO4/FrameData[25] Tile_X1Y0_N_IO4/FrameData[26]
+ Tile_X1Y0_N_IO4/FrameData[27] Tile_X1Y0_N_IO4/FrameData[28] Tile_X1Y0_N_IO4/FrameData[29]
+ Tile_X1Y0_N_IO4/FrameData[2] Tile_X1Y0_N_IO4/FrameData[30] Tile_X1Y0_N_IO4/FrameData[31]
+ Tile_X1Y0_N_IO4/FrameData[3] Tile_X1Y0_N_IO4/FrameData[4] Tile_X1Y0_N_IO4/FrameData[5]
+ Tile_X1Y0_N_IO4/FrameData[6] Tile_X1Y0_N_IO4/FrameData[7] Tile_X1Y0_N_IO4/FrameData[8]
+ Tile_X1Y0_N_IO4/FrameData[9] Tile_X2Y0_N_IO4/FrameData[0] Tile_X2Y0_N_IO4/FrameData[10]
+ Tile_X2Y0_N_IO4/FrameData[11] Tile_X2Y0_N_IO4/FrameData[12] Tile_X2Y0_N_IO4/FrameData[13]
+ Tile_X2Y0_N_IO4/FrameData[14] Tile_X2Y0_N_IO4/FrameData[15] Tile_X2Y0_N_IO4/FrameData[16]
+ Tile_X2Y0_N_IO4/FrameData[17] Tile_X2Y0_N_IO4/FrameData[18] Tile_X2Y0_N_IO4/FrameData[19]
+ Tile_X2Y0_N_IO4/FrameData[1] Tile_X2Y0_N_IO4/FrameData[20] Tile_X2Y0_N_IO4/FrameData[21]
+ Tile_X2Y0_N_IO4/FrameData[22] Tile_X2Y0_N_IO4/FrameData[23] Tile_X2Y0_N_IO4/FrameData[24]
+ Tile_X2Y0_N_IO4/FrameData[25] Tile_X2Y0_N_IO4/FrameData[26] Tile_X2Y0_N_IO4/FrameData[27]
+ Tile_X2Y0_N_IO4/FrameData[28] Tile_X2Y0_N_IO4/FrameData[29] Tile_X2Y0_N_IO4/FrameData[2]
+ Tile_X2Y0_N_IO4/FrameData[30] Tile_X2Y0_N_IO4/FrameData[31] Tile_X2Y0_N_IO4/FrameData[3]
+ Tile_X2Y0_N_IO4/FrameData[4] Tile_X2Y0_N_IO4/FrameData[5] Tile_X2Y0_N_IO4/FrameData[6]
+ Tile_X2Y0_N_IO4/FrameData[7] Tile_X2Y0_N_IO4/FrameData[8] Tile_X2Y0_N_IO4/FrameData[9]
+ Tile_X1Y0_N_IO4/FrameStrobe[0] Tile_X1Y0_N_IO4/FrameStrobe[10] Tile_X1Y0_N_IO4/FrameStrobe[11]
+ Tile_X1Y0_N_IO4/FrameStrobe[12] Tile_X1Y0_N_IO4/FrameStrobe[13] Tile_X1Y0_N_IO4/FrameStrobe[14]
+ Tile_X1Y0_N_IO4/FrameStrobe[15] Tile_X1Y0_N_IO4/FrameStrobe[16] Tile_X1Y0_N_IO4/FrameStrobe[17]
+ Tile_X1Y0_N_IO4/FrameStrobe[18] Tile_X1Y0_N_IO4/FrameStrobe[19] Tile_X1Y0_N_IO4/FrameStrobe[1]
+ Tile_X1Y0_N_IO4/FrameStrobe[2] Tile_X1Y0_N_IO4/FrameStrobe[3] Tile_X1Y0_N_IO4/FrameStrobe[4]
+ Tile_X1Y0_N_IO4/FrameStrobe[5] Tile_X1Y0_N_IO4/FrameStrobe[6] Tile_X1Y0_N_IO4/FrameStrobe[7]
+ Tile_X1Y0_N_IO4/FrameStrobe[8] Tile_X1Y0_N_IO4/FrameStrobe[9] Tile_X1Y0_N_IO4/FrameStrobe_O[0]
+ Tile_X1Y0_N_IO4/FrameStrobe_O[10] Tile_X1Y0_N_IO4/FrameStrobe_O[11] Tile_X1Y0_N_IO4/FrameStrobe_O[12]
+ Tile_X1Y0_N_IO4/FrameStrobe_O[13] Tile_X1Y0_N_IO4/FrameStrobe_O[14] Tile_X1Y0_N_IO4/FrameStrobe_O[15]
+ Tile_X1Y0_N_IO4/FrameStrobe_O[16] Tile_X1Y0_N_IO4/FrameStrobe_O[17] Tile_X1Y0_N_IO4/FrameStrobe_O[18]
+ Tile_X1Y0_N_IO4/FrameStrobe_O[19] Tile_X1Y0_N_IO4/FrameStrobe_O[1] Tile_X1Y0_N_IO4/FrameStrobe_O[2]
+ Tile_X1Y0_N_IO4/FrameStrobe_O[3] Tile_X1Y0_N_IO4/FrameStrobe_O[4] Tile_X1Y0_N_IO4/FrameStrobe_O[5]
+ Tile_X1Y0_N_IO4/FrameStrobe_O[6] Tile_X1Y0_N_IO4/FrameStrobe_O[7] Tile_X1Y0_N_IO4/FrameStrobe_O[8]
+ Tile_X1Y0_N_IO4/FrameStrobe_O[9] Tile_X1Y0_N_IO4/N1END[0] Tile_X1Y0_N_IO4/N1END[1]
+ Tile_X1Y0_N_IO4/N1END[2] Tile_X1Y0_N_IO4/N1END[3] Tile_X1Y0_N_IO4/N2END[0] Tile_X1Y0_N_IO4/N2END[1]
+ Tile_X1Y0_N_IO4/N2END[2] Tile_X1Y0_N_IO4/N2END[3] Tile_X1Y0_N_IO4/N2END[4] Tile_X1Y0_N_IO4/N2END[5]
+ Tile_X1Y0_N_IO4/N2END[6] Tile_X1Y0_N_IO4/N2END[7] Tile_X1Y0_N_IO4/N2MID[0] Tile_X1Y0_N_IO4/N2MID[1]
+ Tile_X1Y0_N_IO4/N2MID[2] Tile_X1Y0_N_IO4/N2MID[3] Tile_X1Y0_N_IO4/N2MID[4] Tile_X1Y0_N_IO4/N2MID[5]
+ Tile_X1Y0_N_IO4/N2MID[6] Tile_X1Y0_N_IO4/N2MID[7] Tile_X1Y0_N_IO4/N4END[0] Tile_X1Y0_N_IO4/N4END[10]
+ Tile_X1Y0_N_IO4/N4END[11] Tile_X1Y0_N_IO4/N4END[12] Tile_X1Y0_N_IO4/N4END[13] Tile_X1Y0_N_IO4/N4END[14]
+ Tile_X1Y0_N_IO4/N4END[15] Tile_X1Y0_N_IO4/N4END[1] Tile_X1Y0_N_IO4/N4END[2] Tile_X1Y0_N_IO4/N4END[3]
+ Tile_X1Y0_N_IO4/N4END[4] Tile_X1Y0_N_IO4/N4END[5] Tile_X1Y0_N_IO4/N4END[6] Tile_X1Y0_N_IO4/N4END[7]
+ Tile_X1Y0_N_IO4/N4END[8] Tile_X1Y0_N_IO4/N4END[9] Tile_X1Y0_N_IO4/NN4END[0] Tile_X1Y0_N_IO4/NN4END[10]
+ Tile_X1Y0_N_IO4/NN4END[11] Tile_X1Y0_N_IO4/NN4END[12] Tile_X1Y0_N_IO4/NN4END[13]
+ Tile_X1Y0_N_IO4/NN4END[14] Tile_X1Y0_N_IO4/NN4END[15] Tile_X1Y0_N_IO4/NN4END[1]
+ Tile_X1Y0_N_IO4/NN4END[2] Tile_X1Y0_N_IO4/NN4END[3] Tile_X1Y0_N_IO4/NN4END[4] Tile_X1Y0_N_IO4/NN4END[5]
+ Tile_X1Y0_N_IO4/NN4END[6] Tile_X1Y0_N_IO4/NN4END[7] Tile_X1Y0_N_IO4/NN4END[8] Tile_X1Y0_N_IO4/NN4END[9]
+ Tile_X1Y0_N_IO4/S1BEG[0] Tile_X1Y0_N_IO4/S1BEG[1] Tile_X1Y0_N_IO4/S1BEG[2] Tile_X1Y0_N_IO4/S1BEG[3]
+ Tile_X1Y0_N_IO4/S2BEG[0] Tile_X1Y0_N_IO4/S2BEG[1] Tile_X1Y0_N_IO4/S2BEG[2] Tile_X1Y0_N_IO4/S2BEG[3]
+ Tile_X1Y0_N_IO4/S2BEG[4] Tile_X1Y0_N_IO4/S2BEG[5] Tile_X1Y0_N_IO4/S2BEG[6] Tile_X1Y0_N_IO4/S2BEG[7]
+ Tile_X1Y1_LUT4AB/S2END[0] Tile_X1Y1_LUT4AB/S2END[1] Tile_X1Y1_LUT4AB/S2END[2] Tile_X1Y1_LUT4AB/S2END[3]
+ Tile_X1Y1_LUT4AB/S2END[4] Tile_X1Y1_LUT4AB/S2END[5] Tile_X1Y1_LUT4AB/S2END[6] Tile_X1Y1_LUT4AB/S2END[7]
+ Tile_X1Y0_N_IO4/S4BEG[0] Tile_X1Y0_N_IO4/S4BEG[10] Tile_X1Y0_N_IO4/S4BEG[11] Tile_X1Y0_N_IO4/S4BEG[12]
+ Tile_X1Y0_N_IO4/S4BEG[13] Tile_X1Y0_N_IO4/S4BEG[14] Tile_X1Y0_N_IO4/S4BEG[15] Tile_X1Y0_N_IO4/S4BEG[1]
+ Tile_X1Y0_N_IO4/S4BEG[2] Tile_X1Y0_N_IO4/S4BEG[3] Tile_X1Y0_N_IO4/S4BEG[4] Tile_X1Y0_N_IO4/S4BEG[5]
+ Tile_X1Y0_N_IO4/S4BEG[6] Tile_X1Y0_N_IO4/S4BEG[7] Tile_X1Y0_N_IO4/S4BEG[8] Tile_X1Y0_N_IO4/S4BEG[9]
+ Tile_X1Y0_N_IO4/SS4BEG[0] Tile_X1Y0_N_IO4/SS4BEG[10] Tile_X1Y0_N_IO4/SS4BEG[11]
+ Tile_X1Y0_N_IO4/SS4BEG[12] Tile_X1Y0_N_IO4/SS4BEG[13] Tile_X1Y0_N_IO4/SS4BEG[14]
+ Tile_X1Y0_N_IO4/SS4BEG[15] Tile_X1Y0_N_IO4/SS4BEG[1] Tile_X1Y0_N_IO4/SS4BEG[2] Tile_X1Y0_N_IO4/SS4BEG[3]
+ Tile_X1Y0_N_IO4/SS4BEG[4] Tile_X1Y0_N_IO4/SS4BEG[5] Tile_X1Y0_N_IO4/SS4BEG[6] Tile_X1Y0_N_IO4/SS4BEG[7]
+ Tile_X1Y0_N_IO4/SS4BEG[8] Tile_X1Y0_N_IO4/SS4BEG[9] Tile_X1Y0_N_IO4/UserCLK Tile_X1Y0_N_IO4/UserCLKo
+ VGND VPWR N_IO4
XTile_X2Y4_LUT4AB Tile_X2Y5_LUT4AB/Co Tile_X2Y4_LUT4AB/Co Tile_X3Y4_LUT4AB/E1END[0]
+ Tile_X3Y4_LUT4AB/E1END[1] Tile_X3Y4_LUT4AB/E1END[2] Tile_X3Y4_LUT4AB/E1END[3] Tile_X2Y4_LUT4AB/E1END[0]
+ Tile_X2Y4_LUT4AB/E1END[1] Tile_X2Y4_LUT4AB/E1END[2] Tile_X2Y4_LUT4AB/E1END[3] Tile_X3Y4_LUT4AB/E2MID[0]
+ Tile_X3Y4_LUT4AB/E2MID[1] Tile_X3Y4_LUT4AB/E2MID[2] Tile_X3Y4_LUT4AB/E2MID[3] Tile_X3Y4_LUT4AB/E2MID[4]
+ Tile_X3Y4_LUT4AB/E2MID[5] Tile_X3Y4_LUT4AB/E2MID[6] Tile_X3Y4_LUT4AB/E2MID[7] Tile_X3Y4_LUT4AB/E2END[0]
+ Tile_X3Y4_LUT4AB/E2END[1] Tile_X3Y4_LUT4AB/E2END[2] Tile_X3Y4_LUT4AB/E2END[3] Tile_X3Y4_LUT4AB/E2END[4]
+ Tile_X3Y4_LUT4AB/E2END[5] Tile_X3Y4_LUT4AB/E2END[6] Tile_X3Y4_LUT4AB/E2END[7] Tile_X2Y4_LUT4AB/E2END[0]
+ Tile_X2Y4_LUT4AB/E2END[1] Tile_X2Y4_LUT4AB/E2END[2] Tile_X2Y4_LUT4AB/E2END[3] Tile_X2Y4_LUT4AB/E2END[4]
+ Tile_X2Y4_LUT4AB/E2END[5] Tile_X2Y4_LUT4AB/E2END[6] Tile_X2Y4_LUT4AB/E2END[7] Tile_X2Y4_LUT4AB/E2MID[0]
+ Tile_X2Y4_LUT4AB/E2MID[1] Tile_X2Y4_LUT4AB/E2MID[2] Tile_X2Y4_LUT4AB/E2MID[3] Tile_X2Y4_LUT4AB/E2MID[4]
+ Tile_X2Y4_LUT4AB/E2MID[5] Tile_X2Y4_LUT4AB/E2MID[6] Tile_X2Y4_LUT4AB/E2MID[7] Tile_X3Y4_LUT4AB/E6END[0]
+ Tile_X3Y4_LUT4AB/E6END[10] Tile_X3Y4_LUT4AB/E6END[11] Tile_X3Y4_LUT4AB/E6END[1]
+ Tile_X3Y4_LUT4AB/E6END[2] Tile_X3Y4_LUT4AB/E6END[3] Tile_X3Y4_LUT4AB/E6END[4] Tile_X3Y4_LUT4AB/E6END[5]
+ Tile_X3Y4_LUT4AB/E6END[6] Tile_X3Y4_LUT4AB/E6END[7] Tile_X3Y4_LUT4AB/E6END[8] Tile_X3Y4_LUT4AB/E6END[9]
+ Tile_X2Y4_LUT4AB/E6END[0] Tile_X2Y4_LUT4AB/E6END[10] Tile_X2Y4_LUT4AB/E6END[11]
+ Tile_X2Y4_LUT4AB/E6END[1] Tile_X2Y4_LUT4AB/E6END[2] Tile_X2Y4_LUT4AB/E6END[3] Tile_X2Y4_LUT4AB/E6END[4]
+ Tile_X2Y4_LUT4AB/E6END[5] Tile_X2Y4_LUT4AB/E6END[6] Tile_X2Y4_LUT4AB/E6END[7] Tile_X2Y4_LUT4AB/E6END[8]
+ Tile_X2Y4_LUT4AB/E6END[9] Tile_X3Y4_LUT4AB/EE4END[0] Tile_X3Y4_LUT4AB/EE4END[10]
+ Tile_X3Y4_LUT4AB/EE4END[11] Tile_X3Y4_LUT4AB/EE4END[12] Tile_X3Y4_LUT4AB/EE4END[13]
+ Tile_X3Y4_LUT4AB/EE4END[14] Tile_X3Y4_LUT4AB/EE4END[15] Tile_X3Y4_LUT4AB/EE4END[1]
+ Tile_X3Y4_LUT4AB/EE4END[2] Tile_X3Y4_LUT4AB/EE4END[3] Tile_X3Y4_LUT4AB/EE4END[4]
+ Tile_X3Y4_LUT4AB/EE4END[5] Tile_X3Y4_LUT4AB/EE4END[6] Tile_X3Y4_LUT4AB/EE4END[7]
+ Tile_X3Y4_LUT4AB/EE4END[8] Tile_X3Y4_LUT4AB/EE4END[9] Tile_X2Y4_LUT4AB/EE4END[0]
+ Tile_X2Y4_LUT4AB/EE4END[10] Tile_X2Y4_LUT4AB/EE4END[11] Tile_X2Y4_LUT4AB/EE4END[12]
+ Tile_X2Y4_LUT4AB/EE4END[13] Tile_X2Y4_LUT4AB/EE4END[14] Tile_X2Y4_LUT4AB/EE4END[15]
+ Tile_X2Y4_LUT4AB/EE4END[1] Tile_X2Y4_LUT4AB/EE4END[2] Tile_X2Y4_LUT4AB/EE4END[3]
+ Tile_X2Y4_LUT4AB/EE4END[4] Tile_X2Y4_LUT4AB/EE4END[5] Tile_X2Y4_LUT4AB/EE4END[6]
+ Tile_X2Y4_LUT4AB/EE4END[7] Tile_X2Y4_LUT4AB/EE4END[8] Tile_X2Y4_LUT4AB/EE4END[9]
+ Tile_X2Y4_LUT4AB/FrameData[0] Tile_X2Y4_LUT4AB/FrameData[10] Tile_X2Y4_LUT4AB/FrameData[11]
+ Tile_X2Y4_LUT4AB/FrameData[12] Tile_X2Y4_LUT4AB/FrameData[13] Tile_X2Y4_LUT4AB/FrameData[14]
+ Tile_X2Y4_LUT4AB/FrameData[15] Tile_X2Y4_LUT4AB/FrameData[16] Tile_X2Y4_LUT4AB/FrameData[17]
+ Tile_X2Y4_LUT4AB/FrameData[18] Tile_X2Y4_LUT4AB/FrameData[19] Tile_X2Y4_LUT4AB/FrameData[1]
+ Tile_X2Y4_LUT4AB/FrameData[20] Tile_X2Y4_LUT4AB/FrameData[21] Tile_X2Y4_LUT4AB/FrameData[22]
+ Tile_X2Y4_LUT4AB/FrameData[23] Tile_X2Y4_LUT4AB/FrameData[24] Tile_X2Y4_LUT4AB/FrameData[25]
+ Tile_X2Y4_LUT4AB/FrameData[26] Tile_X2Y4_LUT4AB/FrameData[27] Tile_X2Y4_LUT4AB/FrameData[28]
+ Tile_X2Y4_LUT4AB/FrameData[29] Tile_X2Y4_LUT4AB/FrameData[2] Tile_X2Y4_LUT4AB/FrameData[30]
+ Tile_X2Y4_LUT4AB/FrameData[31] Tile_X2Y4_LUT4AB/FrameData[3] Tile_X2Y4_LUT4AB/FrameData[4]
+ Tile_X2Y4_LUT4AB/FrameData[5] Tile_X2Y4_LUT4AB/FrameData[6] Tile_X2Y4_LUT4AB/FrameData[7]
+ Tile_X2Y4_LUT4AB/FrameData[8] Tile_X2Y4_LUT4AB/FrameData[9] Tile_X3Y4_LUT4AB/FrameData[0]
+ Tile_X3Y4_LUT4AB/FrameData[10] Tile_X3Y4_LUT4AB/FrameData[11] Tile_X3Y4_LUT4AB/FrameData[12]
+ Tile_X3Y4_LUT4AB/FrameData[13] Tile_X3Y4_LUT4AB/FrameData[14] Tile_X3Y4_LUT4AB/FrameData[15]
+ Tile_X3Y4_LUT4AB/FrameData[16] Tile_X3Y4_LUT4AB/FrameData[17] Tile_X3Y4_LUT4AB/FrameData[18]
+ Tile_X3Y4_LUT4AB/FrameData[19] Tile_X3Y4_LUT4AB/FrameData[1] Tile_X3Y4_LUT4AB/FrameData[20]
+ Tile_X3Y4_LUT4AB/FrameData[21] Tile_X3Y4_LUT4AB/FrameData[22] Tile_X3Y4_LUT4AB/FrameData[23]
+ Tile_X3Y4_LUT4AB/FrameData[24] Tile_X3Y4_LUT4AB/FrameData[25] Tile_X3Y4_LUT4AB/FrameData[26]
+ Tile_X3Y4_LUT4AB/FrameData[27] Tile_X3Y4_LUT4AB/FrameData[28] Tile_X3Y4_LUT4AB/FrameData[29]
+ Tile_X3Y4_LUT4AB/FrameData[2] Tile_X3Y4_LUT4AB/FrameData[30] Tile_X3Y4_LUT4AB/FrameData[31]
+ Tile_X3Y4_LUT4AB/FrameData[3] Tile_X3Y4_LUT4AB/FrameData[4] Tile_X3Y4_LUT4AB/FrameData[5]
+ Tile_X3Y4_LUT4AB/FrameData[6] Tile_X3Y4_LUT4AB/FrameData[7] Tile_X3Y4_LUT4AB/FrameData[8]
+ Tile_X3Y4_LUT4AB/FrameData[9] Tile_X2Y4_LUT4AB/FrameStrobe[0] Tile_X2Y4_LUT4AB/FrameStrobe[10]
+ Tile_X2Y4_LUT4AB/FrameStrobe[11] Tile_X2Y4_LUT4AB/FrameStrobe[12] Tile_X2Y4_LUT4AB/FrameStrobe[13]
+ Tile_X2Y4_LUT4AB/FrameStrobe[14] Tile_X2Y4_LUT4AB/FrameStrobe[15] Tile_X2Y4_LUT4AB/FrameStrobe[16]
+ Tile_X2Y4_LUT4AB/FrameStrobe[17] Tile_X2Y4_LUT4AB/FrameStrobe[18] Tile_X2Y4_LUT4AB/FrameStrobe[19]
+ Tile_X2Y4_LUT4AB/FrameStrobe[1] Tile_X2Y4_LUT4AB/FrameStrobe[2] Tile_X2Y4_LUT4AB/FrameStrobe[3]
+ Tile_X2Y4_LUT4AB/FrameStrobe[4] Tile_X2Y4_LUT4AB/FrameStrobe[5] Tile_X2Y4_LUT4AB/FrameStrobe[6]
+ Tile_X2Y4_LUT4AB/FrameStrobe[7] Tile_X2Y4_LUT4AB/FrameStrobe[8] Tile_X2Y4_LUT4AB/FrameStrobe[9]
+ Tile_X2Y3_LUT4AB/FrameStrobe[0] Tile_X2Y3_LUT4AB/FrameStrobe[10] Tile_X2Y3_LUT4AB/FrameStrobe[11]
+ Tile_X2Y3_LUT4AB/FrameStrobe[12] Tile_X2Y3_LUT4AB/FrameStrobe[13] Tile_X2Y3_LUT4AB/FrameStrobe[14]
+ Tile_X2Y3_LUT4AB/FrameStrobe[15] Tile_X2Y3_LUT4AB/FrameStrobe[16] Tile_X2Y3_LUT4AB/FrameStrobe[17]
+ Tile_X2Y3_LUT4AB/FrameStrobe[18] Tile_X2Y3_LUT4AB/FrameStrobe[19] Tile_X2Y3_LUT4AB/FrameStrobe[1]
+ Tile_X2Y3_LUT4AB/FrameStrobe[2] Tile_X2Y3_LUT4AB/FrameStrobe[3] Tile_X2Y3_LUT4AB/FrameStrobe[4]
+ Tile_X2Y3_LUT4AB/FrameStrobe[5] Tile_X2Y3_LUT4AB/FrameStrobe[6] Tile_X2Y3_LUT4AB/FrameStrobe[7]
+ Tile_X2Y3_LUT4AB/FrameStrobe[8] Tile_X2Y3_LUT4AB/FrameStrobe[9] Tile_X2Y4_LUT4AB/N1BEG[0]
+ Tile_X2Y4_LUT4AB/N1BEG[1] Tile_X2Y4_LUT4AB/N1BEG[2] Tile_X2Y4_LUT4AB/N1BEG[3] Tile_X2Y5_LUT4AB/N1BEG[0]
+ Tile_X2Y5_LUT4AB/N1BEG[1] Tile_X2Y5_LUT4AB/N1BEG[2] Tile_X2Y5_LUT4AB/N1BEG[3] Tile_X2Y4_LUT4AB/N2BEG[0]
+ Tile_X2Y4_LUT4AB/N2BEG[1] Tile_X2Y4_LUT4AB/N2BEG[2] Tile_X2Y4_LUT4AB/N2BEG[3] Tile_X2Y4_LUT4AB/N2BEG[4]
+ Tile_X2Y4_LUT4AB/N2BEG[5] Tile_X2Y4_LUT4AB/N2BEG[6] Tile_X2Y4_LUT4AB/N2BEG[7] Tile_X2Y3_LUT4AB/N2END[0]
+ Tile_X2Y3_LUT4AB/N2END[1] Tile_X2Y3_LUT4AB/N2END[2] Tile_X2Y3_LUT4AB/N2END[3] Tile_X2Y3_LUT4AB/N2END[4]
+ Tile_X2Y3_LUT4AB/N2END[5] Tile_X2Y3_LUT4AB/N2END[6] Tile_X2Y3_LUT4AB/N2END[7] Tile_X2Y4_LUT4AB/N2END[0]
+ Tile_X2Y4_LUT4AB/N2END[1] Tile_X2Y4_LUT4AB/N2END[2] Tile_X2Y4_LUT4AB/N2END[3] Tile_X2Y4_LUT4AB/N2END[4]
+ Tile_X2Y4_LUT4AB/N2END[5] Tile_X2Y4_LUT4AB/N2END[6] Tile_X2Y4_LUT4AB/N2END[7] Tile_X2Y5_LUT4AB/N2BEG[0]
+ Tile_X2Y5_LUT4AB/N2BEG[1] Tile_X2Y5_LUT4AB/N2BEG[2] Tile_X2Y5_LUT4AB/N2BEG[3] Tile_X2Y5_LUT4AB/N2BEG[4]
+ Tile_X2Y5_LUT4AB/N2BEG[5] Tile_X2Y5_LUT4AB/N2BEG[6] Tile_X2Y5_LUT4AB/N2BEG[7] Tile_X2Y4_LUT4AB/N4BEG[0]
+ Tile_X2Y4_LUT4AB/N4BEG[10] Tile_X2Y4_LUT4AB/N4BEG[11] Tile_X2Y4_LUT4AB/N4BEG[12]
+ Tile_X2Y4_LUT4AB/N4BEG[13] Tile_X2Y4_LUT4AB/N4BEG[14] Tile_X2Y4_LUT4AB/N4BEG[15]
+ Tile_X2Y4_LUT4AB/N4BEG[1] Tile_X2Y4_LUT4AB/N4BEG[2] Tile_X2Y4_LUT4AB/N4BEG[3] Tile_X2Y4_LUT4AB/N4BEG[4]
+ Tile_X2Y4_LUT4AB/N4BEG[5] Tile_X2Y4_LUT4AB/N4BEG[6] Tile_X2Y4_LUT4AB/N4BEG[7] Tile_X2Y4_LUT4AB/N4BEG[8]
+ Tile_X2Y4_LUT4AB/N4BEG[9] Tile_X2Y5_LUT4AB/N4BEG[0] Tile_X2Y5_LUT4AB/N4BEG[10] Tile_X2Y5_LUT4AB/N4BEG[11]
+ Tile_X2Y5_LUT4AB/N4BEG[12] Tile_X2Y5_LUT4AB/N4BEG[13] Tile_X2Y5_LUT4AB/N4BEG[14]
+ Tile_X2Y5_LUT4AB/N4BEG[15] Tile_X2Y5_LUT4AB/N4BEG[1] Tile_X2Y5_LUT4AB/N4BEG[2] Tile_X2Y5_LUT4AB/N4BEG[3]
+ Tile_X2Y5_LUT4AB/N4BEG[4] Tile_X2Y5_LUT4AB/N4BEG[5] Tile_X2Y5_LUT4AB/N4BEG[6] Tile_X2Y5_LUT4AB/N4BEG[7]
+ Tile_X2Y5_LUT4AB/N4BEG[8] Tile_X2Y5_LUT4AB/N4BEG[9] Tile_X2Y4_LUT4AB/NN4BEG[0] Tile_X2Y4_LUT4AB/NN4BEG[10]
+ Tile_X2Y4_LUT4AB/NN4BEG[11] Tile_X2Y4_LUT4AB/NN4BEG[12] Tile_X2Y4_LUT4AB/NN4BEG[13]
+ Tile_X2Y4_LUT4AB/NN4BEG[14] Tile_X2Y4_LUT4AB/NN4BEG[15] Tile_X2Y4_LUT4AB/NN4BEG[1]
+ Tile_X2Y4_LUT4AB/NN4BEG[2] Tile_X2Y4_LUT4AB/NN4BEG[3] Tile_X2Y4_LUT4AB/NN4BEG[4]
+ Tile_X2Y4_LUT4AB/NN4BEG[5] Tile_X2Y4_LUT4AB/NN4BEG[6] Tile_X2Y4_LUT4AB/NN4BEG[7]
+ Tile_X2Y4_LUT4AB/NN4BEG[8] Tile_X2Y4_LUT4AB/NN4BEG[9] Tile_X2Y5_LUT4AB/NN4BEG[0]
+ Tile_X2Y5_LUT4AB/NN4BEG[10] Tile_X2Y5_LUT4AB/NN4BEG[11] Tile_X2Y5_LUT4AB/NN4BEG[12]
+ Tile_X2Y5_LUT4AB/NN4BEG[13] Tile_X2Y5_LUT4AB/NN4BEG[14] Tile_X2Y5_LUT4AB/NN4BEG[15]
+ Tile_X2Y5_LUT4AB/NN4BEG[1] Tile_X2Y5_LUT4AB/NN4BEG[2] Tile_X2Y5_LUT4AB/NN4BEG[3]
+ Tile_X2Y5_LUT4AB/NN4BEG[4] Tile_X2Y5_LUT4AB/NN4BEG[5] Tile_X2Y5_LUT4AB/NN4BEG[6]
+ Tile_X2Y5_LUT4AB/NN4BEG[7] Tile_X2Y5_LUT4AB/NN4BEG[8] Tile_X2Y5_LUT4AB/NN4BEG[9]
+ Tile_X2Y5_LUT4AB/S1END[0] Tile_X2Y5_LUT4AB/S1END[1] Tile_X2Y5_LUT4AB/S1END[2] Tile_X2Y5_LUT4AB/S1END[3]
+ Tile_X2Y4_LUT4AB/S1END[0] Tile_X2Y4_LUT4AB/S1END[1] Tile_X2Y4_LUT4AB/S1END[2] Tile_X2Y4_LUT4AB/S1END[3]
+ Tile_X2Y5_LUT4AB/S2MID[0] Tile_X2Y5_LUT4AB/S2MID[1] Tile_X2Y5_LUT4AB/S2MID[2] Tile_X2Y5_LUT4AB/S2MID[3]
+ Tile_X2Y5_LUT4AB/S2MID[4] Tile_X2Y5_LUT4AB/S2MID[5] Tile_X2Y5_LUT4AB/S2MID[6] Tile_X2Y5_LUT4AB/S2MID[7]
+ Tile_X2Y5_LUT4AB/S2END[0] Tile_X2Y5_LUT4AB/S2END[1] Tile_X2Y5_LUT4AB/S2END[2] Tile_X2Y5_LUT4AB/S2END[3]
+ Tile_X2Y5_LUT4AB/S2END[4] Tile_X2Y5_LUT4AB/S2END[5] Tile_X2Y5_LUT4AB/S2END[6] Tile_X2Y5_LUT4AB/S2END[7]
+ Tile_X2Y4_LUT4AB/S2END[0] Tile_X2Y4_LUT4AB/S2END[1] Tile_X2Y4_LUT4AB/S2END[2] Tile_X2Y4_LUT4AB/S2END[3]
+ Tile_X2Y4_LUT4AB/S2END[4] Tile_X2Y4_LUT4AB/S2END[5] Tile_X2Y4_LUT4AB/S2END[6] Tile_X2Y4_LUT4AB/S2END[7]
+ Tile_X2Y4_LUT4AB/S2MID[0] Tile_X2Y4_LUT4AB/S2MID[1] Tile_X2Y4_LUT4AB/S2MID[2] Tile_X2Y4_LUT4AB/S2MID[3]
+ Tile_X2Y4_LUT4AB/S2MID[4] Tile_X2Y4_LUT4AB/S2MID[5] Tile_X2Y4_LUT4AB/S2MID[6] Tile_X2Y4_LUT4AB/S2MID[7]
+ Tile_X2Y5_LUT4AB/S4END[0] Tile_X2Y5_LUT4AB/S4END[10] Tile_X2Y5_LUT4AB/S4END[11]
+ Tile_X2Y5_LUT4AB/S4END[12] Tile_X2Y5_LUT4AB/S4END[13] Tile_X2Y5_LUT4AB/S4END[14]
+ Tile_X2Y5_LUT4AB/S4END[15] Tile_X2Y5_LUT4AB/S4END[1] Tile_X2Y5_LUT4AB/S4END[2] Tile_X2Y5_LUT4AB/S4END[3]
+ Tile_X2Y5_LUT4AB/S4END[4] Tile_X2Y5_LUT4AB/S4END[5] Tile_X2Y5_LUT4AB/S4END[6] Tile_X2Y5_LUT4AB/S4END[7]
+ Tile_X2Y5_LUT4AB/S4END[8] Tile_X2Y5_LUT4AB/S4END[9] Tile_X2Y4_LUT4AB/S4END[0] Tile_X2Y4_LUT4AB/S4END[10]
+ Tile_X2Y4_LUT4AB/S4END[11] Tile_X2Y4_LUT4AB/S4END[12] Tile_X2Y4_LUT4AB/S4END[13]
+ Tile_X2Y4_LUT4AB/S4END[14] Tile_X2Y4_LUT4AB/S4END[15] Tile_X2Y4_LUT4AB/S4END[1]
+ Tile_X2Y4_LUT4AB/S4END[2] Tile_X2Y4_LUT4AB/S4END[3] Tile_X2Y4_LUT4AB/S4END[4] Tile_X2Y4_LUT4AB/S4END[5]
+ Tile_X2Y4_LUT4AB/S4END[6] Tile_X2Y4_LUT4AB/S4END[7] Tile_X2Y4_LUT4AB/S4END[8] Tile_X2Y4_LUT4AB/S4END[9]
+ Tile_X2Y5_LUT4AB/SS4END[0] Tile_X2Y5_LUT4AB/SS4END[10] Tile_X2Y5_LUT4AB/SS4END[11]
+ Tile_X2Y5_LUT4AB/SS4END[12] Tile_X2Y5_LUT4AB/SS4END[13] Tile_X2Y5_LUT4AB/SS4END[14]
+ Tile_X2Y5_LUT4AB/SS4END[15] Tile_X2Y5_LUT4AB/SS4END[1] Tile_X2Y5_LUT4AB/SS4END[2]
+ Tile_X2Y5_LUT4AB/SS4END[3] Tile_X2Y5_LUT4AB/SS4END[4] Tile_X2Y5_LUT4AB/SS4END[5]
+ Tile_X2Y5_LUT4AB/SS4END[6] Tile_X2Y5_LUT4AB/SS4END[7] Tile_X2Y5_LUT4AB/SS4END[8]
+ Tile_X2Y5_LUT4AB/SS4END[9] Tile_X2Y4_LUT4AB/SS4END[0] Tile_X2Y4_LUT4AB/SS4END[10]
+ Tile_X2Y4_LUT4AB/SS4END[11] Tile_X2Y4_LUT4AB/SS4END[12] Tile_X2Y4_LUT4AB/SS4END[13]
+ Tile_X2Y4_LUT4AB/SS4END[14] Tile_X2Y4_LUT4AB/SS4END[15] Tile_X2Y4_LUT4AB/SS4END[1]
+ Tile_X2Y4_LUT4AB/SS4END[2] Tile_X2Y4_LUT4AB/SS4END[3] Tile_X2Y4_LUT4AB/SS4END[4]
+ Tile_X2Y4_LUT4AB/SS4END[5] Tile_X2Y4_LUT4AB/SS4END[6] Tile_X2Y4_LUT4AB/SS4END[7]
+ Tile_X2Y4_LUT4AB/SS4END[8] Tile_X2Y4_LUT4AB/SS4END[9] Tile_X2Y4_LUT4AB/UserCLK Tile_X2Y3_LUT4AB/UserCLK
+ VGND VPWR Tile_X2Y4_LUT4AB/W1BEG[0] Tile_X2Y4_LUT4AB/W1BEG[1] Tile_X2Y4_LUT4AB/W1BEG[2]
+ Tile_X2Y4_LUT4AB/W1BEG[3] Tile_X3Y4_LUT4AB/W1BEG[0] Tile_X3Y4_LUT4AB/W1BEG[1] Tile_X3Y4_LUT4AB/W1BEG[2]
+ Tile_X3Y4_LUT4AB/W1BEG[3] Tile_X2Y4_LUT4AB/W2BEG[0] Tile_X2Y4_LUT4AB/W2BEG[1] Tile_X2Y4_LUT4AB/W2BEG[2]
+ Tile_X2Y4_LUT4AB/W2BEG[3] Tile_X2Y4_LUT4AB/W2BEG[4] Tile_X2Y4_LUT4AB/W2BEG[5] Tile_X2Y4_LUT4AB/W2BEG[6]
+ Tile_X2Y4_LUT4AB/W2BEG[7] Tile_X1Y4_LUT4AB/W2END[0] Tile_X1Y4_LUT4AB/W2END[1] Tile_X1Y4_LUT4AB/W2END[2]
+ Tile_X1Y4_LUT4AB/W2END[3] Tile_X1Y4_LUT4AB/W2END[4] Tile_X1Y4_LUT4AB/W2END[5] Tile_X1Y4_LUT4AB/W2END[6]
+ Tile_X1Y4_LUT4AB/W2END[7] Tile_X2Y4_LUT4AB/W2END[0] Tile_X2Y4_LUT4AB/W2END[1] Tile_X2Y4_LUT4AB/W2END[2]
+ Tile_X2Y4_LUT4AB/W2END[3] Tile_X2Y4_LUT4AB/W2END[4] Tile_X2Y4_LUT4AB/W2END[5] Tile_X2Y4_LUT4AB/W2END[6]
+ Tile_X2Y4_LUT4AB/W2END[7] Tile_X3Y4_LUT4AB/W2BEG[0] Tile_X3Y4_LUT4AB/W2BEG[1] Tile_X3Y4_LUT4AB/W2BEG[2]
+ Tile_X3Y4_LUT4AB/W2BEG[3] Tile_X3Y4_LUT4AB/W2BEG[4] Tile_X3Y4_LUT4AB/W2BEG[5] Tile_X3Y4_LUT4AB/W2BEG[6]
+ Tile_X3Y4_LUT4AB/W2BEG[7] Tile_X2Y4_LUT4AB/W6BEG[0] Tile_X2Y4_LUT4AB/W6BEG[10] Tile_X2Y4_LUT4AB/W6BEG[11]
+ Tile_X2Y4_LUT4AB/W6BEG[1] Tile_X2Y4_LUT4AB/W6BEG[2] Tile_X2Y4_LUT4AB/W6BEG[3] Tile_X2Y4_LUT4AB/W6BEG[4]
+ Tile_X2Y4_LUT4AB/W6BEG[5] Tile_X2Y4_LUT4AB/W6BEG[6] Tile_X2Y4_LUT4AB/W6BEG[7] Tile_X2Y4_LUT4AB/W6BEG[8]
+ Tile_X2Y4_LUT4AB/W6BEG[9] Tile_X3Y4_LUT4AB/W6BEG[0] Tile_X3Y4_LUT4AB/W6BEG[10] Tile_X3Y4_LUT4AB/W6BEG[11]
+ Tile_X3Y4_LUT4AB/W6BEG[1] Tile_X3Y4_LUT4AB/W6BEG[2] Tile_X3Y4_LUT4AB/W6BEG[3] Tile_X3Y4_LUT4AB/W6BEG[4]
+ Tile_X3Y4_LUT4AB/W6BEG[5] Tile_X3Y4_LUT4AB/W6BEG[6] Tile_X3Y4_LUT4AB/W6BEG[7] Tile_X3Y4_LUT4AB/W6BEG[8]
+ Tile_X3Y4_LUT4AB/W6BEG[9] Tile_X2Y4_LUT4AB/WW4BEG[0] Tile_X2Y4_LUT4AB/WW4BEG[10]
+ Tile_X2Y4_LUT4AB/WW4BEG[11] Tile_X2Y4_LUT4AB/WW4BEG[12] Tile_X2Y4_LUT4AB/WW4BEG[13]
+ Tile_X2Y4_LUT4AB/WW4BEG[14] Tile_X2Y4_LUT4AB/WW4BEG[15] Tile_X2Y4_LUT4AB/WW4BEG[1]
+ Tile_X2Y4_LUT4AB/WW4BEG[2] Tile_X2Y4_LUT4AB/WW4BEG[3] Tile_X2Y4_LUT4AB/WW4BEG[4]
+ Tile_X2Y4_LUT4AB/WW4BEG[5] Tile_X2Y4_LUT4AB/WW4BEG[6] Tile_X2Y4_LUT4AB/WW4BEG[7]
+ Tile_X2Y4_LUT4AB/WW4BEG[8] Tile_X2Y4_LUT4AB/WW4BEG[9] Tile_X3Y4_LUT4AB/WW4BEG[0]
+ Tile_X3Y4_LUT4AB/WW4BEG[10] Tile_X3Y4_LUT4AB/WW4BEG[11] Tile_X3Y4_LUT4AB/WW4BEG[12]
+ Tile_X3Y4_LUT4AB/WW4BEG[13] Tile_X3Y4_LUT4AB/WW4BEG[14] Tile_X3Y4_LUT4AB/WW4BEG[15]
+ Tile_X3Y4_LUT4AB/WW4BEG[1] Tile_X3Y4_LUT4AB/WW4BEG[2] Tile_X3Y4_LUT4AB/WW4BEG[3]
+ Tile_X3Y4_LUT4AB/WW4BEG[4] Tile_X3Y4_LUT4AB/WW4BEG[5] Tile_X3Y4_LUT4AB/WW4BEG[6]
+ Tile_X3Y4_LUT4AB/WW4BEG[7] Tile_X3Y4_LUT4AB/WW4BEG[8] Tile_X3Y4_LUT4AB/WW4BEG[9]
+ LUT4AB
XTile_X1Y8_LUT4AB Tile_X1Y9_S_IO4/Co Tile_X1Y8_LUT4AB/Co Tile_X2Y8_LUT4AB/E1END[0]
+ Tile_X2Y8_LUT4AB/E1END[1] Tile_X2Y8_LUT4AB/E1END[2] Tile_X2Y8_LUT4AB/E1END[3] Tile_X1Y8_LUT4AB/E1END[0]
+ Tile_X1Y8_LUT4AB/E1END[1] Tile_X1Y8_LUT4AB/E1END[2] Tile_X1Y8_LUT4AB/E1END[3] Tile_X2Y8_LUT4AB/E2MID[0]
+ Tile_X2Y8_LUT4AB/E2MID[1] Tile_X2Y8_LUT4AB/E2MID[2] Tile_X2Y8_LUT4AB/E2MID[3] Tile_X2Y8_LUT4AB/E2MID[4]
+ Tile_X2Y8_LUT4AB/E2MID[5] Tile_X2Y8_LUT4AB/E2MID[6] Tile_X2Y8_LUT4AB/E2MID[7] Tile_X2Y8_LUT4AB/E2END[0]
+ Tile_X2Y8_LUT4AB/E2END[1] Tile_X2Y8_LUT4AB/E2END[2] Tile_X2Y8_LUT4AB/E2END[3] Tile_X2Y8_LUT4AB/E2END[4]
+ Tile_X2Y8_LUT4AB/E2END[5] Tile_X2Y8_LUT4AB/E2END[6] Tile_X2Y8_LUT4AB/E2END[7] Tile_X1Y8_LUT4AB/E2END[0]
+ Tile_X1Y8_LUT4AB/E2END[1] Tile_X1Y8_LUT4AB/E2END[2] Tile_X1Y8_LUT4AB/E2END[3] Tile_X1Y8_LUT4AB/E2END[4]
+ Tile_X1Y8_LUT4AB/E2END[5] Tile_X1Y8_LUT4AB/E2END[6] Tile_X1Y8_LUT4AB/E2END[7] Tile_X1Y8_LUT4AB/E2MID[0]
+ Tile_X1Y8_LUT4AB/E2MID[1] Tile_X1Y8_LUT4AB/E2MID[2] Tile_X1Y8_LUT4AB/E2MID[3] Tile_X1Y8_LUT4AB/E2MID[4]
+ Tile_X1Y8_LUT4AB/E2MID[5] Tile_X1Y8_LUT4AB/E2MID[6] Tile_X1Y8_LUT4AB/E2MID[7] Tile_X2Y8_LUT4AB/E6END[0]
+ Tile_X2Y8_LUT4AB/E6END[10] Tile_X2Y8_LUT4AB/E6END[11] Tile_X2Y8_LUT4AB/E6END[1]
+ Tile_X2Y8_LUT4AB/E6END[2] Tile_X2Y8_LUT4AB/E6END[3] Tile_X2Y8_LUT4AB/E6END[4] Tile_X2Y8_LUT4AB/E6END[5]
+ Tile_X2Y8_LUT4AB/E6END[6] Tile_X2Y8_LUT4AB/E6END[7] Tile_X2Y8_LUT4AB/E6END[8] Tile_X2Y8_LUT4AB/E6END[9]
+ Tile_X1Y8_LUT4AB/E6END[0] Tile_X1Y8_LUT4AB/E6END[10] Tile_X1Y8_LUT4AB/E6END[11]
+ Tile_X1Y8_LUT4AB/E6END[1] Tile_X1Y8_LUT4AB/E6END[2] Tile_X1Y8_LUT4AB/E6END[3] Tile_X1Y8_LUT4AB/E6END[4]
+ Tile_X1Y8_LUT4AB/E6END[5] Tile_X1Y8_LUT4AB/E6END[6] Tile_X1Y8_LUT4AB/E6END[7] Tile_X1Y8_LUT4AB/E6END[8]
+ Tile_X1Y8_LUT4AB/E6END[9] Tile_X2Y8_LUT4AB/EE4END[0] Tile_X2Y8_LUT4AB/EE4END[10]
+ Tile_X2Y8_LUT4AB/EE4END[11] Tile_X2Y8_LUT4AB/EE4END[12] Tile_X2Y8_LUT4AB/EE4END[13]
+ Tile_X2Y8_LUT4AB/EE4END[14] Tile_X2Y8_LUT4AB/EE4END[15] Tile_X2Y8_LUT4AB/EE4END[1]
+ Tile_X2Y8_LUT4AB/EE4END[2] Tile_X2Y8_LUT4AB/EE4END[3] Tile_X2Y8_LUT4AB/EE4END[4]
+ Tile_X2Y8_LUT4AB/EE4END[5] Tile_X2Y8_LUT4AB/EE4END[6] Tile_X2Y8_LUT4AB/EE4END[7]
+ Tile_X2Y8_LUT4AB/EE4END[8] Tile_X2Y8_LUT4AB/EE4END[9] Tile_X1Y8_LUT4AB/EE4END[0]
+ Tile_X1Y8_LUT4AB/EE4END[10] Tile_X1Y8_LUT4AB/EE4END[11] Tile_X1Y8_LUT4AB/EE4END[12]
+ Tile_X1Y8_LUT4AB/EE4END[13] Tile_X1Y8_LUT4AB/EE4END[14] Tile_X1Y8_LUT4AB/EE4END[15]
+ Tile_X1Y8_LUT4AB/EE4END[1] Tile_X1Y8_LUT4AB/EE4END[2] Tile_X1Y8_LUT4AB/EE4END[3]
+ Tile_X1Y8_LUT4AB/EE4END[4] Tile_X1Y8_LUT4AB/EE4END[5] Tile_X1Y8_LUT4AB/EE4END[6]
+ Tile_X1Y8_LUT4AB/EE4END[7] Tile_X1Y8_LUT4AB/EE4END[8] Tile_X1Y8_LUT4AB/EE4END[9]
+ Tile_X1Y8_LUT4AB/FrameData[0] Tile_X1Y8_LUT4AB/FrameData[10] Tile_X1Y8_LUT4AB/FrameData[11]
+ Tile_X1Y8_LUT4AB/FrameData[12] Tile_X1Y8_LUT4AB/FrameData[13] Tile_X1Y8_LUT4AB/FrameData[14]
+ Tile_X1Y8_LUT4AB/FrameData[15] Tile_X1Y8_LUT4AB/FrameData[16] Tile_X1Y8_LUT4AB/FrameData[17]
+ Tile_X1Y8_LUT4AB/FrameData[18] Tile_X1Y8_LUT4AB/FrameData[19] Tile_X1Y8_LUT4AB/FrameData[1]
+ Tile_X1Y8_LUT4AB/FrameData[20] Tile_X1Y8_LUT4AB/FrameData[21] Tile_X1Y8_LUT4AB/FrameData[22]
+ Tile_X1Y8_LUT4AB/FrameData[23] Tile_X1Y8_LUT4AB/FrameData[24] Tile_X1Y8_LUT4AB/FrameData[25]
+ Tile_X1Y8_LUT4AB/FrameData[26] Tile_X1Y8_LUT4AB/FrameData[27] Tile_X1Y8_LUT4AB/FrameData[28]
+ Tile_X1Y8_LUT4AB/FrameData[29] Tile_X1Y8_LUT4AB/FrameData[2] Tile_X1Y8_LUT4AB/FrameData[30]
+ Tile_X1Y8_LUT4AB/FrameData[31] Tile_X1Y8_LUT4AB/FrameData[3] Tile_X1Y8_LUT4AB/FrameData[4]
+ Tile_X1Y8_LUT4AB/FrameData[5] Tile_X1Y8_LUT4AB/FrameData[6] Tile_X1Y8_LUT4AB/FrameData[7]
+ Tile_X1Y8_LUT4AB/FrameData[8] Tile_X1Y8_LUT4AB/FrameData[9] Tile_X2Y8_LUT4AB/FrameData[0]
+ Tile_X2Y8_LUT4AB/FrameData[10] Tile_X2Y8_LUT4AB/FrameData[11] Tile_X2Y8_LUT4AB/FrameData[12]
+ Tile_X2Y8_LUT4AB/FrameData[13] Tile_X2Y8_LUT4AB/FrameData[14] Tile_X2Y8_LUT4AB/FrameData[15]
+ Tile_X2Y8_LUT4AB/FrameData[16] Tile_X2Y8_LUT4AB/FrameData[17] Tile_X2Y8_LUT4AB/FrameData[18]
+ Tile_X2Y8_LUT4AB/FrameData[19] Tile_X2Y8_LUT4AB/FrameData[1] Tile_X2Y8_LUT4AB/FrameData[20]
+ Tile_X2Y8_LUT4AB/FrameData[21] Tile_X2Y8_LUT4AB/FrameData[22] Tile_X2Y8_LUT4AB/FrameData[23]
+ Tile_X2Y8_LUT4AB/FrameData[24] Tile_X2Y8_LUT4AB/FrameData[25] Tile_X2Y8_LUT4AB/FrameData[26]
+ Tile_X2Y8_LUT4AB/FrameData[27] Tile_X2Y8_LUT4AB/FrameData[28] Tile_X2Y8_LUT4AB/FrameData[29]
+ Tile_X2Y8_LUT4AB/FrameData[2] Tile_X2Y8_LUT4AB/FrameData[30] Tile_X2Y8_LUT4AB/FrameData[31]
+ Tile_X2Y8_LUT4AB/FrameData[3] Tile_X2Y8_LUT4AB/FrameData[4] Tile_X2Y8_LUT4AB/FrameData[5]
+ Tile_X2Y8_LUT4AB/FrameData[6] Tile_X2Y8_LUT4AB/FrameData[7] Tile_X2Y8_LUT4AB/FrameData[8]
+ Tile_X2Y8_LUT4AB/FrameData[9] Tile_X1Y8_LUT4AB/FrameStrobe[0] Tile_X1Y8_LUT4AB/FrameStrobe[10]
+ Tile_X1Y8_LUT4AB/FrameStrobe[11] Tile_X1Y8_LUT4AB/FrameStrobe[12] Tile_X1Y8_LUT4AB/FrameStrobe[13]
+ Tile_X1Y8_LUT4AB/FrameStrobe[14] Tile_X1Y8_LUT4AB/FrameStrobe[15] Tile_X1Y8_LUT4AB/FrameStrobe[16]
+ Tile_X1Y8_LUT4AB/FrameStrobe[17] Tile_X1Y8_LUT4AB/FrameStrobe[18] Tile_X1Y8_LUT4AB/FrameStrobe[19]
+ Tile_X1Y8_LUT4AB/FrameStrobe[1] Tile_X1Y8_LUT4AB/FrameStrobe[2] Tile_X1Y8_LUT4AB/FrameStrobe[3]
+ Tile_X1Y8_LUT4AB/FrameStrobe[4] Tile_X1Y8_LUT4AB/FrameStrobe[5] Tile_X1Y8_LUT4AB/FrameStrobe[6]
+ Tile_X1Y8_LUT4AB/FrameStrobe[7] Tile_X1Y8_LUT4AB/FrameStrobe[8] Tile_X1Y8_LUT4AB/FrameStrobe[9]
+ Tile_X1Y7_LUT4AB/FrameStrobe[0] Tile_X1Y7_LUT4AB/FrameStrobe[10] Tile_X1Y7_LUT4AB/FrameStrobe[11]
+ Tile_X1Y7_LUT4AB/FrameStrobe[12] Tile_X1Y7_LUT4AB/FrameStrobe[13] Tile_X1Y7_LUT4AB/FrameStrobe[14]
+ Tile_X1Y7_LUT4AB/FrameStrobe[15] Tile_X1Y7_LUT4AB/FrameStrobe[16] Tile_X1Y7_LUT4AB/FrameStrobe[17]
+ Tile_X1Y7_LUT4AB/FrameStrobe[18] Tile_X1Y7_LUT4AB/FrameStrobe[19] Tile_X1Y7_LUT4AB/FrameStrobe[1]
+ Tile_X1Y7_LUT4AB/FrameStrobe[2] Tile_X1Y7_LUT4AB/FrameStrobe[3] Tile_X1Y7_LUT4AB/FrameStrobe[4]
+ Tile_X1Y7_LUT4AB/FrameStrobe[5] Tile_X1Y7_LUT4AB/FrameStrobe[6] Tile_X1Y7_LUT4AB/FrameStrobe[7]
+ Tile_X1Y7_LUT4AB/FrameStrobe[8] Tile_X1Y7_LUT4AB/FrameStrobe[9] Tile_X1Y8_LUT4AB/N1BEG[0]
+ Tile_X1Y8_LUT4AB/N1BEG[1] Tile_X1Y8_LUT4AB/N1BEG[2] Tile_X1Y8_LUT4AB/N1BEG[3] Tile_X1Y9_S_IO4/N1BEG[0]
+ Tile_X1Y9_S_IO4/N1BEG[1] Tile_X1Y9_S_IO4/N1BEG[2] Tile_X1Y9_S_IO4/N1BEG[3] Tile_X1Y8_LUT4AB/N2BEG[0]
+ Tile_X1Y8_LUT4AB/N2BEG[1] Tile_X1Y8_LUT4AB/N2BEG[2] Tile_X1Y8_LUT4AB/N2BEG[3] Tile_X1Y8_LUT4AB/N2BEG[4]
+ Tile_X1Y8_LUT4AB/N2BEG[5] Tile_X1Y8_LUT4AB/N2BEG[6] Tile_X1Y8_LUT4AB/N2BEG[7] Tile_X1Y7_LUT4AB/N2END[0]
+ Tile_X1Y7_LUT4AB/N2END[1] Tile_X1Y7_LUT4AB/N2END[2] Tile_X1Y7_LUT4AB/N2END[3] Tile_X1Y7_LUT4AB/N2END[4]
+ Tile_X1Y7_LUT4AB/N2END[5] Tile_X1Y7_LUT4AB/N2END[6] Tile_X1Y7_LUT4AB/N2END[7] Tile_X1Y9_S_IO4/N2BEGb[0]
+ Tile_X1Y9_S_IO4/N2BEGb[1] Tile_X1Y9_S_IO4/N2BEGb[2] Tile_X1Y9_S_IO4/N2BEGb[3] Tile_X1Y9_S_IO4/N2BEGb[4]
+ Tile_X1Y9_S_IO4/N2BEGb[5] Tile_X1Y9_S_IO4/N2BEGb[6] Tile_X1Y9_S_IO4/N2BEGb[7] Tile_X1Y9_S_IO4/N2BEG[0]
+ Tile_X1Y9_S_IO4/N2BEG[1] Tile_X1Y9_S_IO4/N2BEG[2] Tile_X1Y9_S_IO4/N2BEG[3] Tile_X1Y9_S_IO4/N2BEG[4]
+ Tile_X1Y9_S_IO4/N2BEG[5] Tile_X1Y9_S_IO4/N2BEG[6] Tile_X1Y9_S_IO4/N2BEG[7] Tile_X1Y8_LUT4AB/N4BEG[0]
+ Tile_X1Y8_LUT4AB/N4BEG[10] Tile_X1Y8_LUT4AB/N4BEG[11] Tile_X1Y8_LUT4AB/N4BEG[12]
+ Tile_X1Y8_LUT4AB/N4BEG[13] Tile_X1Y8_LUT4AB/N4BEG[14] Tile_X1Y8_LUT4AB/N4BEG[15]
+ Tile_X1Y8_LUT4AB/N4BEG[1] Tile_X1Y8_LUT4AB/N4BEG[2] Tile_X1Y8_LUT4AB/N4BEG[3] Tile_X1Y8_LUT4AB/N4BEG[4]
+ Tile_X1Y8_LUT4AB/N4BEG[5] Tile_X1Y8_LUT4AB/N4BEG[6] Tile_X1Y8_LUT4AB/N4BEG[7] Tile_X1Y8_LUT4AB/N4BEG[8]
+ Tile_X1Y8_LUT4AB/N4BEG[9] Tile_X1Y9_S_IO4/N4BEG[0] Tile_X1Y9_S_IO4/N4BEG[10] Tile_X1Y9_S_IO4/N4BEG[11]
+ Tile_X1Y9_S_IO4/N4BEG[12] Tile_X1Y9_S_IO4/N4BEG[13] Tile_X1Y9_S_IO4/N4BEG[14] Tile_X1Y9_S_IO4/N4BEG[15]
+ Tile_X1Y9_S_IO4/N4BEG[1] Tile_X1Y9_S_IO4/N4BEG[2] Tile_X1Y9_S_IO4/N4BEG[3] Tile_X1Y9_S_IO4/N4BEG[4]
+ Tile_X1Y9_S_IO4/N4BEG[5] Tile_X1Y9_S_IO4/N4BEG[6] Tile_X1Y9_S_IO4/N4BEG[7] Tile_X1Y9_S_IO4/N4BEG[8]
+ Tile_X1Y9_S_IO4/N4BEG[9] Tile_X1Y8_LUT4AB/NN4BEG[0] Tile_X1Y8_LUT4AB/NN4BEG[10]
+ Tile_X1Y8_LUT4AB/NN4BEG[11] Tile_X1Y8_LUT4AB/NN4BEG[12] Tile_X1Y8_LUT4AB/NN4BEG[13]
+ Tile_X1Y8_LUT4AB/NN4BEG[14] Tile_X1Y8_LUT4AB/NN4BEG[15] Tile_X1Y8_LUT4AB/NN4BEG[1]
+ Tile_X1Y8_LUT4AB/NN4BEG[2] Tile_X1Y8_LUT4AB/NN4BEG[3] Tile_X1Y8_LUT4AB/NN4BEG[4]
+ Tile_X1Y8_LUT4AB/NN4BEG[5] Tile_X1Y8_LUT4AB/NN4BEG[6] Tile_X1Y8_LUT4AB/NN4BEG[7]
+ Tile_X1Y8_LUT4AB/NN4BEG[8] Tile_X1Y8_LUT4AB/NN4BEG[9] Tile_X1Y9_S_IO4/NN4BEG[0]
+ Tile_X1Y9_S_IO4/NN4BEG[10] Tile_X1Y9_S_IO4/NN4BEG[11] Tile_X1Y9_S_IO4/NN4BEG[12]
+ Tile_X1Y9_S_IO4/NN4BEG[13] Tile_X1Y9_S_IO4/NN4BEG[14] Tile_X1Y9_S_IO4/NN4BEG[15]
+ Tile_X1Y9_S_IO4/NN4BEG[1] Tile_X1Y9_S_IO4/NN4BEG[2] Tile_X1Y9_S_IO4/NN4BEG[3] Tile_X1Y9_S_IO4/NN4BEG[4]
+ Tile_X1Y9_S_IO4/NN4BEG[5] Tile_X1Y9_S_IO4/NN4BEG[6] Tile_X1Y9_S_IO4/NN4BEG[7] Tile_X1Y9_S_IO4/NN4BEG[8]
+ Tile_X1Y9_S_IO4/NN4BEG[9] Tile_X1Y9_S_IO4/S1END[0] Tile_X1Y9_S_IO4/S1END[1] Tile_X1Y9_S_IO4/S1END[2]
+ Tile_X1Y9_S_IO4/S1END[3] Tile_X1Y8_LUT4AB/S1END[0] Tile_X1Y8_LUT4AB/S1END[1] Tile_X1Y8_LUT4AB/S1END[2]
+ Tile_X1Y8_LUT4AB/S1END[3] Tile_X1Y9_S_IO4/S2MID[0] Tile_X1Y9_S_IO4/S2MID[1] Tile_X1Y9_S_IO4/S2MID[2]
+ Tile_X1Y9_S_IO4/S2MID[3] Tile_X1Y9_S_IO4/S2MID[4] Tile_X1Y9_S_IO4/S2MID[5] Tile_X1Y9_S_IO4/S2MID[6]
+ Tile_X1Y9_S_IO4/S2MID[7] Tile_X1Y9_S_IO4/S2END[0] Tile_X1Y9_S_IO4/S2END[1] Tile_X1Y9_S_IO4/S2END[2]
+ Tile_X1Y9_S_IO4/S2END[3] Tile_X1Y9_S_IO4/S2END[4] Tile_X1Y9_S_IO4/S2END[5] Tile_X1Y9_S_IO4/S2END[6]
+ Tile_X1Y9_S_IO4/S2END[7] Tile_X1Y8_LUT4AB/S2END[0] Tile_X1Y8_LUT4AB/S2END[1] Tile_X1Y8_LUT4AB/S2END[2]
+ Tile_X1Y8_LUT4AB/S2END[3] Tile_X1Y8_LUT4AB/S2END[4] Tile_X1Y8_LUT4AB/S2END[5] Tile_X1Y8_LUT4AB/S2END[6]
+ Tile_X1Y8_LUT4AB/S2END[7] Tile_X1Y8_LUT4AB/S2MID[0] Tile_X1Y8_LUT4AB/S2MID[1] Tile_X1Y8_LUT4AB/S2MID[2]
+ Tile_X1Y8_LUT4AB/S2MID[3] Tile_X1Y8_LUT4AB/S2MID[4] Tile_X1Y8_LUT4AB/S2MID[5] Tile_X1Y8_LUT4AB/S2MID[6]
+ Tile_X1Y8_LUT4AB/S2MID[7] Tile_X1Y9_S_IO4/S4END[0] Tile_X1Y9_S_IO4/S4END[10] Tile_X1Y9_S_IO4/S4END[11]
+ Tile_X1Y9_S_IO4/S4END[12] Tile_X1Y9_S_IO4/S4END[13] Tile_X1Y9_S_IO4/S4END[14] Tile_X1Y9_S_IO4/S4END[15]
+ Tile_X1Y9_S_IO4/S4END[1] Tile_X1Y9_S_IO4/S4END[2] Tile_X1Y9_S_IO4/S4END[3] Tile_X1Y9_S_IO4/S4END[4]
+ Tile_X1Y9_S_IO4/S4END[5] Tile_X1Y9_S_IO4/S4END[6] Tile_X1Y9_S_IO4/S4END[7] Tile_X1Y9_S_IO4/S4END[8]
+ Tile_X1Y9_S_IO4/S4END[9] Tile_X1Y8_LUT4AB/S4END[0] Tile_X1Y8_LUT4AB/S4END[10] Tile_X1Y8_LUT4AB/S4END[11]
+ Tile_X1Y8_LUT4AB/S4END[12] Tile_X1Y8_LUT4AB/S4END[13] Tile_X1Y8_LUT4AB/S4END[14]
+ Tile_X1Y8_LUT4AB/S4END[15] Tile_X1Y8_LUT4AB/S4END[1] Tile_X1Y8_LUT4AB/S4END[2] Tile_X1Y8_LUT4AB/S4END[3]
+ Tile_X1Y8_LUT4AB/S4END[4] Tile_X1Y8_LUT4AB/S4END[5] Tile_X1Y8_LUT4AB/S4END[6] Tile_X1Y8_LUT4AB/S4END[7]
+ Tile_X1Y8_LUT4AB/S4END[8] Tile_X1Y8_LUT4AB/S4END[9] Tile_X1Y9_S_IO4/SS4END[0] Tile_X1Y9_S_IO4/SS4END[10]
+ Tile_X1Y9_S_IO4/SS4END[11] Tile_X1Y9_S_IO4/SS4END[12] Tile_X1Y9_S_IO4/SS4END[13]
+ Tile_X1Y9_S_IO4/SS4END[14] Tile_X1Y9_S_IO4/SS4END[15] Tile_X1Y9_S_IO4/SS4END[1]
+ Tile_X1Y9_S_IO4/SS4END[2] Tile_X1Y9_S_IO4/SS4END[3] Tile_X1Y9_S_IO4/SS4END[4] Tile_X1Y9_S_IO4/SS4END[5]
+ Tile_X1Y9_S_IO4/SS4END[6] Tile_X1Y9_S_IO4/SS4END[7] Tile_X1Y9_S_IO4/SS4END[8] Tile_X1Y9_S_IO4/SS4END[9]
+ Tile_X1Y8_LUT4AB/SS4END[0] Tile_X1Y8_LUT4AB/SS4END[10] Tile_X1Y8_LUT4AB/SS4END[11]
+ Tile_X1Y8_LUT4AB/SS4END[12] Tile_X1Y8_LUT4AB/SS4END[13] Tile_X1Y8_LUT4AB/SS4END[14]
+ Tile_X1Y8_LUT4AB/SS4END[15] Tile_X1Y8_LUT4AB/SS4END[1] Tile_X1Y8_LUT4AB/SS4END[2]
+ Tile_X1Y8_LUT4AB/SS4END[3] Tile_X1Y8_LUT4AB/SS4END[4] Tile_X1Y8_LUT4AB/SS4END[5]
+ Tile_X1Y8_LUT4AB/SS4END[6] Tile_X1Y8_LUT4AB/SS4END[7] Tile_X1Y8_LUT4AB/SS4END[8]
+ Tile_X1Y8_LUT4AB/SS4END[9] Tile_X1Y9_S_IO4/UserCLKo Tile_X1Y7_LUT4AB/UserCLK VGND
+ VPWR Tile_X1Y8_LUT4AB/W1BEG[0] Tile_X1Y8_LUT4AB/W1BEG[1] Tile_X1Y8_LUT4AB/W1BEG[2]
+ Tile_X1Y8_LUT4AB/W1BEG[3] Tile_X2Y8_LUT4AB/W1BEG[0] Tile_X2Y8_LUT4AB/W1BEG[1] Tile_X2Y8_LUT4AB/W1BEG[2]
+ Tile_X2Y8_LUT4AB/W1BEG[3] Tile_X1Y8_LUT4AB/W2BEG[0] Tile_X1Y8_LUT4AB/W2BEG[1] Tile_X1Y8_LUT4AB/W2BEG[2]
+ Tile_X1Y8_LUT4AB/W2BEG[3] Tile_X1Y8_LUT4AB/W2BEG[4] Tile_X1Y8_LUT4AB/W2BEG[5] Tile_X1Y8_LUT4AB/W2BEG[6]
+ Tile_X1Y8_LUT4AB/W2BEG[7] Tile_X1Y8_LUT4AB/W2BEGb[0] Tile_X1Y8_LUT4AB/W2BEGb[1]
+ Tile_X1Y8_LUT4AB/W2BEGb[2] Tile_X1Y8_LUT4AB/W2BEGb[3] Tile_X1Y8_LUT4AB/W2BEGb[4]
+ Tile_X1Y8_LUT4AB/W2BEGb[5] Tile_X1Y8_LUT4AB/W2BEGb[6] Tile_X1Y8_LUT4AB/W2BEGb[7]
+ Tile_X1Y8_LUT4AB/W2END[0] Tile_X1Y8_LUT4AB/W2END[1] Tile_X1Y8_LUT4AB/W2END[2] Tile_X1Y8_LUT4AB/W2END[3]
+ Tile_X1Y8_LUT4AB/W2END[4] Tile_X1Y8_LUT4AB/W2END[5] Tile_X1Y8_LUT4AB/W2END[6] Tile_X1Y8_LUT4AB/W2END[7]
+ Tile_X2Y8_LUT4AB/W2BEG[0] Tile_X2Y8_LUT4AB/W2BEG[1] Tile_X2Y8_LUT4AB/W2BEG[2] Tile_X2Y8_LUT4AB/W2BEG[3]
+ Tile_X2Y8_LUT4AB/W2BEG[4] Tile_X2Y8_LUT4AB/W2BEG[5] Tile_X2Y8_LUT4AB/W2BEG[6] Tile_X2Y8_LUT4AB/W2BEG[7]
+ Tile_X1Y8_LUT4AB/W6BEG[0] Tile_X1Y8_LUT4AB/W6BEG[10] Tile_X1Y8_LUT4AB/W6BEG[11]
+ Tile_X1Y8_LUT4AB/W6BEG[1] Tile_X1Y8_LUT4AB/W6BEG[2] Tile_X1Y8_LUT4AB/W6BEG[3] Tile_X1Y8_LUT4AB/W6BEG[4]
+ Tile_X1Y8_LUT4AB/W6BEG[5] Tile_X1Y8_LUT4AB/W6BEG[6] Tile_X1Y8_LUT4AB/W6BEG[7] Tile_X1Y8_LUT4AB/W6BEG[8]
+ Tile_X1Y8_LUT4AB/W6BEG[9] Tile_X2Y8_LUT4AB/W6BEG[0] Tile_X2Y8_LUT4AB/W6BEG[10] Tile_X2Y8_LUT4AB/W6BEG[11]
+ Tile_X2Y8_LUT4AB/W6BEG[1] Tile_X2Y8_LUT4AB/W6BEG[2] Tile_X2Y8_LUT4AB/W6BEG[3] Tile_X2Y8_LUT4AB/W6BEG[4]
+ Tile_X2Y8_LUT4AB/W6BEG[5] Tile_X2Y8_LUT4AB/W6BEG[6] Tile_X2Y8_LUT4AB/W6BEG[7] Tile_X2Y8_LUT4AB/W6BEG[8]
+ Tile_X2Y8_LUT4AB/W6BEG[9] Tile_X1Y8_LUT4AB/WW4BEG[0] Tile_X1Y8_LUT4AB/WW4BEG[10]
+ Tile_X1Y8_LUT4AB/WW4BEG[11] Tile_X1Y8_LUT4AB/WW4BEG[12] Tile_X1Y8_LUT4AB/WW4BEG[13]
+ Tile_X1Y8_LUT4AB/WW4BEG[14] Tile_X1Y8_LUT4AB/WW4BEG[15] Tile_X1Y8_LUT4AB/WW4BEG[1]
+ Tile_X1Y8_LUT4AB/WW4BEG[2] Tile_X1Y8_LUT4AB/WW4BEG[3] Tile_X1Y8_LUT4AB/WW4BEG[4]
+ Tile_X1Y8_LUT4AB/WW4BEG[5] Tile_X1Y8_LUT4AB/WW4BEG[6] Tile_X1Y8_LUT4AB/WW4BEG[7]
+ Tile_X1Y8_LUT4AB/WW4BEG[8] Tile_X1Y8_LUT4AB/WW4BEG[9] Tile_X2Y8_LUT4AB/WW4BEG[0]
+ Tile_X2Y8_LUT4AB/WW4BEG[10] Tile_X2Y8_LUT4AB/WW4BEG[11] Tile_X2Y8_LUT4AB/WW4BEG[12]
+ Tile_X2Y8_LUT4AB/WW4BEG[13] Tile_X2Y8_LUT4AB/WW4BEG[14] Tile_X2Y8_LUT4AB/WW4BEG[15]
+ Tile_X2Y8_LUT4AB/WW4BEG[1] Tile_X2Y8_LUT4AB/WW4BEG[2] Tile_X2Y8_LUT4AB/WW4BEG[3]
+ Tile_X2Y8_LUT4AB/WW4BEG[4] Tile_X2Y8_LUT4AB/WW4BEG[5] Tile_X2Y8_LUT4AB/WW4BEG[6]
+ Tile_X2Y8_LUT4AB/WW4BEG[7] Tile_X2Y8_LUT4AB/WW4BEG[8] Tile_X2Y8_LUT4AB/WW4BEG[9]
+ LUT4AB
XTile_X0Y0_NW_term FrameData[0] FrameData[10] FrameData[11] FrameData[12] FrameData[13]
+ FrameData[14] FrameData[15] FrameData[16] FrameData[17] FrameData[18] FrameData[19]
+ FrameData[1] FrameData[20] FrameData[21] FrameData[22] FrameData[23] FrameData[24]
+ FrameData[25] FrameData[26] FrameData[27] FrameData[28] FrameData[29] FrameData[2]
+ FrameData[30] FrameData[31] FrameData[3] FrameData[4] FrameData[5] FrameData[6]
+ FrameData[7] FrameData[8] FrameData[9] Tile_X1Y0_N_IO4/FrameData[0] Tile_X1Y0_N_IO4/FrameData[10]
+ Tile_X1Y0_N_IO4/FrameData[11] Tile_X1Y0_N_IO4/FrameData[12] Tile_X1Y0_N_IO4/FrameData[13]
+ Tile_X1Y0_N_IO4/FrameData[14] Tile_X1Y0_N_IO4/FrameData[15] Tile_X1Y0_N_IO4/FrameData[16]
+ Tile_X1Y0_N_IO4/FrameData[17] Tile_X1Y0_N_IO4/FrameData[18] Tile_X1Y0_N_IO4/FrameData[19]
+ Tile_X1Y0_N_IO4/FrameData[1] Tile_X1Y0_N_IO4/FrameData[20] Tile_X1Y0_N_IO4/FrameData[21]
+ Tile_X1Y0_N_IO4/FrameData[22] Tile_X1Y0_N_IO4/FrameData[23] Tile_X1Y0_N_IO4/FrameData[24]
+ Tile_X1Y0_N_IO4/FrameData[25] Tile_X1Y0_N_IO4/FrameData[26] Tile_X1Y0_N_IO4/FrameData[27]
+ Tile_X1Y0_N_IO4/FrameData[28] Tile_X1Y0_N_IO4/FrameData[29] Tile_X1Y0_N_IO4/FrameData[2]
+ Tile_X1Y0_N_IO4/FrameData[30] Tile_X1Y0_N_IO4/FrameData[31] Tile_X1Y0_N_IO4/FrameData[3]
+ Tile_X1Y0_N_IO4/FrameData[4] Tile_X1Y0_N_IO4/FrameData[5] Tile_X1Y0_N_IO4/FrameData[6]
+ Tile_X1Y0_N_IO4/FrameData[7] Tile_X1Y0_N_IO4/FrameData[8] Tile_X1Y0_N_IO4/FrameData[9]
+ Tile_X0Y0_NW_term/FrameStrobe[0] Tile_X0Y0_NW_term/FrameStrobe[10] Tile_X0Y0_NW_term/FrameStrobe[11]
+ Tile_X0Y0_NW_term/FrameStrobe[12] Tile_X0Y0_NW_term/FrameStrobe[13] Tile_X0Y0_NW_term/FrameStrobe[14]
+ Tile_X0Y0_NW_term/FrameStrobe[15] Tile_X0Y0_NW_term/FrameStrobe[16] Tile_X0Y0_NW_term/FrameStrobe[17]
+ Tile_X0Y0_NW_term/FrameStrobe[18] Tile_X0Y0_NW_term/FrameStrobe[19] Tile_X0Y0_NW_term/FrameStrobe[1]
+ Tile_X0Y0_NW_term/FrameStrobe[2] Tile_X0Y0_NW_term/FrameStrobe[3] Tile_X0Y0_NW_term/FrameStrobe[4]
+ Tile_X0Y0_NW_term/FrameStrobe[5] Tile_X0Y0_NW_term/FrameStrobe[6] Tile_X0Y0_NW_term/FrameStrobe[7]
+ Tile_X0Y0_NW_term/FrameStrobe[8] Tile_X0Y0_NW_term/FrameStrobe[9] Tile_X0Y0_NW_term/FrameStrobe_O[0]
+ Tile_X0Y0_NW_term/FrameStrobe_O[10] Tile_X0Y0_NW_term/FrameStrobe_O[11] Tile_X0Y0_NW_term/FrameStrobe_O[12]
+ Tile_X0Y0_NW_term/FrameStrobe_O[13] Tile_X0Y0_NW_term/FrameStrobe_O[14] Tile_X0Y0_NW_term/FrameStrobe_O[15]
+ Tile_X0Y0_NW_term/FrameStrobe_O[16] Tile_X0Y0_NW_term/FrameStrobe_O[17] Tile_X0Y0_NW_term/FrameStrobe_O[18]
+ Tile_X0Y0_NW_term/FrameStrobe_O[19] Tile_X0Y0_NW_term/FrameStrobe_O[1] Tile_X0Y0_NW_term/FrameStrobe_O[2]
+ Tile_X0Y0_NW_term/FrameStrobe_O[3] Tile_X0Y0_NW_term/FrameStrobe_O[4] Tile_X0Y0_NW_term/FrameStrobe_O[5]
+ Tile_X0Y0_NW_term/FrameStrobe_O[6] Tile_X0Y0_NW_term/FrameStrobe_O[7] Tile_X0Y0_NW_term/FrameStrobe_O[8]
+ Tile_X0Y0_NW_term/FrameStrobe_O[9] Tile_X0Y1_W_TT_IF/N1BEG[0] Tile_X0Y1_W_TT_IF/N1BEG[1]
+ Tile_X0Y1_W_TT_IF/N1BEG[2] Tile_X0Y1_W_TT_IF/N1BEG[3] Tile_X0Y0_NW_term/N2END[0]
+ Tile_X0Y0_NW_term/N2END[1] Tile_X0Y0_NW_term/N2END[2] Tile_X0Y0_NW_term/N2END[3]
+ Tile_X0Y0_NW_term/N2END[4] Tile_X0Y0_NW_term/N2END[5] Tile_X0Y0_NW_term/N2END[6]
+ Tile_X0Y0_NW_term/N2END[7] Tile_X0Y1_W_TT_IF/N2BEG[0] Tile_X0Y1_W_TT_IF/N2BEG[1]
+ Tile_X0Y1_W_TT_IF/N2BEG[2] Tile_X0Y1_W_TT_IF/N2BEG[3] Tile_X0Y1_W_TT_IF/N2BEG[4]
+ Tile_X0Y1_W_TT_IF/N2BEG[5] Tile_X0Y1_W_TT_IF/N2BEG[6] Tile_X0Y1_W_TT_IF/N2BEG[7]
+ Tile_X0Y1_W_TT_IF/N4BEG[0] Tile_X0Y1_W_TT_IF/N4BEG[10] Tile_X0Y1_W_TT_IF/N4BEG[11]
+ Tile_X0Y1_W_TT_IF/N4BEG[12] Tile_X0Y1_W_TT_IF/N4BEG[13] Tile_X0Y1_W_TT_IF/N4BEG[14]
+ Tile_X0Y1_W_TT_IF/N4BEG[15] Tile_X0Y1_W_TT_IF/N4BEG[1] Tile_X0Y1_W_TT_IF/N4BEG[2]
+ Tile_X0Y1_W_TT_IF/N4BEG[3] Tile_X0Y1_W_TT_IF/N4BEG[4] Tile_X0Y1_W_TT_IF/N4BEG[5]
+ Tile_X0Y1_W_TT_IF/N4BEG[6] Tile_X0Y1_W_TT_IF/N4BEG[7] Tile_X0Y1_W_TT_IF/N4BEG[8]
+ Tile_X0Y1_W_TT_IF/N4BEG[9] Tile_X0Y1_W_TT_IF/S1END[0] Tile_X0Y1_W_TT_IF/S1END[1]
+ Tile_X0Y1_W_TT_IF/S1END[2] Tile_X0Y1_W_TT_IF/S1END[3] Tile_X0Y1_W_TT_IF/S2MID[0]
+ Tile_X0Y1_W_TT_IF/S2MID[1] Tile_X0Y1_W_TT_IF/S2MID[2] Tile_X0Y1_W_TT_IF/S2MID[3]
+ Tile_X0Y1_W_TT_IF/S2MID[4] Tile_X0Y1_W_TT_IF/S2MID[5] Tile_X0Y1_W_TT_IF/S2MID[6]
+ Tile_X0Y1_W_TT_IF/S2MID[7] Tile_X0Y1_W_TT_IF/S2END[0] Tile_X0Y1_W_TT_IF/S2END[1]
+ Tile_X0Y1_W_TT_IF/S2END[2] Tile_X0Y1_W_TT_IF/S2END[3] Tile_X0Y1_W_TT_IF/S2END[4]
+ Tile_X0Y1_W_TT_IF/S2END[5] Tile_X0Y1_W_TT_IF/S2END[6] Tile_X0Y1_W_TT_IF/S2END[7]
+ Tile_X0Y1_W_TT_IF/S4END[0] Tile_X0Y1_W_TT_IF/S4END[10] Tile_X0Y1_W_TT_IF/S4END[11]
+ Tile_X0Y1_W_TT_IF/S4END[12] Tile_X0Y1_W_TT_IF/S4END[13] Tile_X0Y1_W_TT_IF/S4END[14]
+ Tile_X0Y1_W_TT_IF/S4END[15] Tile_X0Y1_W_TT_IF/S4END[1] Tile_X0Y1_W_TT_IF/S4END[2]
+ Tile_X0Y1_W_TT_IF/S4END[3] Tile_X0Y1_W_TT_IF/S4END[4] Tile_X0Y1_W_TT_IF/S4END[5]
+ Tile_X0Y1_W_TT_IF/S4END[6] Tile_X0Y1_W_TT_IF/S4END[7] Tile_X0Y1_W_TT_IF/S4END[8]
+ Tile_X0Y1_W_TT_IF/S4END[9] Tile_X0Y0_NW_term/UserCLK Tile_X0Y0_NW_term/UserCLKo
+ VGND VPWR NW_term
XTile_X4Y2_LUT4AB Tile_X4Y3_LUT4AB/Co Tile_X4Y2_LUT4AB/Co Tile_X4Y2_LUT4AB/E1BEG[0]
+ Tile_X4Y2_LUT4AB/E1BEG[1] Tile_X4Y2_LUT4AB/E1BEG[2] Tile_X4Y2_LUT4AB/E1BEG[3] Tile_X4Y2_LUT4AB/E1END[0]
+ Tile_X4Y2_LUT4AB/E1END[1] Tile_X4Y2_LUT4AB/E1END[2] Tile_X4Y2_LUT4AB/E1END[3] Tile_X4Y2_LUT4AB/E2BEG[0]
+ Tile_X4Y2_LUT4AB/E2BEG[1] Tile_X4Y2_LUT4AB/E2BEG[2] Tile_X4Y2_LUT4AB/E2BEG[3] Tile_X4Y2_LUT4AB/E2BEG[4]
+ Tile_X4Y2_LUT4AB/E2BEG[5] Tile_X4Y2_LUT4AB/E2BEG[6] Tile_X4Y2_LUT4AB/E2BEG[7] Tile_X4Y2_LUT4AB/E2BEGb[0]
+ Tile_X4Y2_LUT4AB/E2BEGb[1] Tile_X4Y2_LUT4AB/E2BEGb[2] Tile_X4Y2_LUT4AB/E2BEGb[3]
+ Tile_X4Y2_LUT4AB/E2BEGb[4] Tile_X4Y2_LUT4AB/E2BEGb[5] Tile_X4Y2_LUT4AB/E2BEGb[6]
+ Tile_X4Y2_LUT4AB/E2BEGb[7] Tile_X4Y2_LUT4AB/E2END[0] Tile_X4Y2_LUT4AB/E2END[1] Tile_X4Y2_LUT4AB/E2END[2]
+ Tile_X4Y2_LUT4AB/E2END[3] Tile_X4Y2_LUT4AB/E2END[4] Tile_X4Y2_LUT4AB/E2END[5] Tile_X4Y2_LUT4AB/E2END[6]
+ Tile_X4Y2_LUT4AB/E2END[7] Tile_X4Y2_LUT4AB/E2MID[0] Tile_X4Y2_LUT4AB/E2MID[1] Tile_X4Y2_LUT4AB/E2MID[2]
+ Tile_X4Y2_LUT4AB/E2MID[3] Tile_X4Y2_LUT4AB/E2MID[4] Tile_X4Y2_LUT4AB/E2MID[5] Tile_X4Y2_LUT4AB/E2MID[6]
+ Tile_X4Y2_LUT4AB/E2MID[7] Tile_X4Y2_LUT4AB/E6BEG[0] Tile_X4Y2_LUT4AB/E6BEG[10] Tile_X4Y2_LUT4AB/E6BEG[11]
+ Tile_X4Y2_LUT4AB/E6BEG[1] Tile_X4Y2_LUT4AB/E6BEG[2] Tile_X4Y2_LUT4AB/E6BEG[3] Tile_X4Y2_LUT4AB/E6BEG[4]
+ Tile_X4Y2_LUT4AB/E6BEG[5] Tile_X4Y2_LUT4AB/E6BEG[6] Tile_X4Y2_LUT4AB/E6BEG[7] Tile_X4Y2_LUT4AB/E6BEG[8]
+ Tile_X4Y2_LUT4AB/E6BEG[9] Tile_X4Y2_LUT4AB/E6END[0] Tile_X4Y2_LUT4AB/E6END[10] Tile_X4Y2_LUT4AB/E6END[11]
+ Tile_X4Y2_LUT4AB/E6END[1] Tile_X4Y2_LUT4AB/E6END[2] Tile_X4Y2_LUT4AB/E6END[3] Tile_X4Y2_LUT4AB/E6END[4]
+ Tile_X4Y2_LUT4AB/E6END[5] Tile_X4Y2_LUT4AB/E6END[6] Tile_X4Y2_LUT4AB/E6END[7] Tile_X4Y2_LUT4AB/E6END[8]
+ Tile_X4Y2_LUT4AB/E6END[9] Tile_X4Y2_LUT4AB/EE4BEG[0] Tile_X4Y2_LUT4AB/EE4BEG[10]
+ Tile_X4Y2_LUT4AB/EE4BEG[11] Tile_X4Y2_LUT4AB/EE4BEG[12] Tile_X4Y2_LUT4AB/EE4BEG[13]
+ Tile_X4Y2_LUT4AB/EE4BEG[14] Tile_X4Y2_LUT4AB/EE4BEG[15] Tile_X4Y2_LUT4AB/EE4BEG[1]
+ Tile_X4Y2_LUT4AB/EE4BEG[2] Tile_X4Y2_LUT4AB/EE4BEG[3] Tile_X4Y2_LUT4AB/EE4BEG[4]
+ Tile_X4Y2_LUT4AB/EE4BEG[5] Tile_X4Y2_LUT4AB/EE4BEG[6] Tile_X4Y2_LUT4AB/EE4BEG[7]
+ Tile_X4Y2_LUT4AB/EE4BEG[8] Tile_X4Y2_LUT4AB/EE4BEG[9] Tile_X4Y2_LUT4AB/EE4END[0]
+ Tile_X4Y2_LUT4AB/EE4END[10] Tile_X4Y2_LUT4AB/EE4END[11] Tile_X4Y2_LUT4AB/EE4END[12]
+ Tile_X4Y2_LUT4AB/EE4END[13] Tile_X4Y2_LUT4AB/EE4END[14] Tile_X4Y2_LUT4AB/EE4END[15]
+ Tile_X4Y2_LUT4AB/EE4END[1] Tile_X4Y2_LUT4AB/EE4END[2] Tile_X4Y2_LUT4AB/EE4END[3]
+ Tile_X4Y2_LUT4AB/EE4END[4] Tile_X4Y2_LUT4AB/EE4END[5] Tile_X4Y2_LUT4AB/EE4END[6]
+ Tile_X4Y2_LUT4AB/EE4END[7] Tile_X4Y2_LUT4AB/EE4END[8] Tile_X4Y2_LUT4AB/EE4END[9]
+ Tile_X4Y2_LUT4AB/FrameData[0] Tile_X4Y2_LUT4AB/FrameData[10] Tile_X4Y2_LUT4AB/FrameData[11]
+ Tile_X4Y2_LUT4AB/FrameData[12] Tile_X4Y2_LUT4AB/FrameData[13] Tile_X4Y2_LUT4AB/FrameData[14]
+ Tile_X4Y2_LUT4AB/FrameData[15] Tile_X4Y2_LUT4AB/FrameData[16] Tile_X4Y2_LUT4AB/FrameData[17]
+ Tile_X4Y2_LUT4AB/FrameData[18] Tile_X4Y2_LUT4AB/FrameData[19] Tile_X4Y2_LUT4AB/FrameData[1]
+ Tile_X4Y2_LUT4AB/FrameData[20] Tile_X4Y2_LUT4AB/FrameData[21] Tile_X4Y2_LUT4AB/FrameData[22]
+ Tile_X4Y2_LUT4AB/FrameData[23] Tile_X4Y2_LUT4AB/FrameData[24] Tile_X4Y2_LUT4AB/FrameData[25]
+ Tile_X4Y2_LUT4AB/FrameData[26] Tile_X4Y2_LUT4AB/FrameData[27] Tile_X4Y2_LUT4AB/FrameData[28]
+ Tile_X4Y2_LUT4AB/FrameData[29] Tile_X4Y2_LUT4AB/FrameData[2] Tile_X4Y2_LUT4AB/FrameData[30]
+ Tile_X4Y2_LUT4AB/FrameData[31] Tile_X4Y2_LUT4AB/FrameData[3] Tile_X4Y2_LUT4AB/FrameData[4]
+ Tile_X4Y2_LUT4AB/FrameData[5] Tile_X4Y2_LUT4AB/FrameData[6] Tile_X4Y2_LUT4AB/FrameData[7]
+ Tile_X4Y2_LUT4AB/FrameData[8] Tile_X4Y2_LUT4AB/FrameData[9] Tile_X4Y2_LUT4AB/FrameData_O[0]
+ Tile_X4Y2_LUT4AB/FrameData_O[10] Tile_X4Y2_LUT4AB/FrameData_O[11] Tile_X4Y2_LUT4AB/FrameData_O[12]
+ Tile_X4Y2_LUT4AB/FrameData_O[13] Tile_X4Y2_LUT4AB/FrameData_O[14] Tile_X4Y2_LUT4AB/FrameData_O[15]
+ Tile_X4Y2_LUT4AB/FrameData_O[16] Tile_X4Y2_LUT4AB/FrameData_O[17] Tile_X4Y2_LUT4AB/FrameData_O[18]
+ Tile_X4Y2_LUT4AB/FrameData_O[19] Tile_X4Y2_LUT4AB/FrameData_O[1] Tile_X4Y2_LUT4AB/FrameData_O[20]
+ Tile_X4Y2_LUT4AB/FrameData_O[21] Tile_X4Y2_LUT4AB/FrameData_O[22] Tile_X4Y2_LUT4AB/FrameData_O[23]
+ Tile_X4Y2_LUT4AB/FrameData_O[24] Tile_X4Y2_LUT4AB/FrameData_O[25] Tile_X4Y2_LUT4AB/FrameData_O[26]
+ Tile_X4Y2_LUT4AB/FrameData_O[27] Tile_X4Y2_LUT4AB/FrameData_O[28] Tile_X4Y2_LUT4AB/FrameData_O[29]
+ Tile_X4Y2_LUT4AB/FrameData_O[2] Tile_X4Y2_LUT4AB/FrameData_O[30] Tile_X4Y2_LUT4AB/FrameData_O[31]
+ Tile_X4Y2_LUT4AB/FrameData_O[3] Tile_X4Y2_LUT4AB/FrameData_O[4] Tile_X4Y2_LUT4AB/FrameData_O[5]
+ Tile_X4Y2_LUT4AB/FrameData_O[6] Tile_X4Y2_LUT4AB/FrameData_O[7] Tile_X4Y2_LUT4AB/FrameData_O[8]
+ Tile_X4Y2_LUT4AB/FrameData_O[9] Tile_X4Y2_LUT4AB/FrameStrobe[0] Tile_X4Y2_LUT4AB/FrameStrobe[10]
+ Tile_X4Y2_LUT4AB/FrameStrobe[11] Tile_X4Y2_LUT4AB/FrameStrobe[12] Tile_X4Y2_LUT4AB/FrameStrobe[13]
+ Tile_X4Y2_LUT4AB/FrameStrobe[14] Tile_X4Y2_LUT4AB/FrameStrobe[15] Tile_X4Y2_LUT4AB/FrameStrobe[16]
+ Tile_X4Y2_LUT4AB/FrameStrobe[17] Tile_X4Y2_LUT4AB/FrameStrobe[18] Tile_X4Y2_LUT4AB/FrameStrobe[19]
+ Tile_X4Y2_LUT4AB/FrameStrobe[1] Tile_X4Y2_LUT4AB/FrameStrobe[2] Tile_X4Y2_LUT4AB/FrameStrobe[3]
+ Tile_X4Y2_LUT4AB/FrameStrobe[4] Tile_X4Y2_LUT4AB/FrameStrobe[5] Tile_X4Y2_LUT4AB/FrameStrobe[6]
+ Tile_X4Y2_LUT4AB/FrameStrobe[7] Tile_X4Y2_LUT4AB/FrameStrobe[8] Tile_X4Y2_LUT4AB/FrameStrobe[9]
+ Tile_X4Y1_LUT4AB/FrameStrobe[0] Tile_X4Y1_LUT4AB/FrameStrobe[10] Tile_X4Y1_LUT4AB/FrameStrobe[11]
+ Tile_X4Y1_LUT4AB/FrameStrobe[12] Tile_X4Y1_LUT4AB/FrameStrobe[13] Tile_X4Y1_LUT4AB/FrameStrobe[14]
+ Tile_X4Y1_LUT4AB/FrameStrobe[15] Tile_X4Y1_LUT4AB/FrameStrobe[16] Tile_X4Y1_LUT4AB/FrameStrobe[17]
+ Tile_X4Y1_LUT4AB/FrameStrobe[18] Tile_X4Y1_LUT4AB/FrameStrobe[19] Tile_X4Y1_LUT4AB/FrameStrobe[1]
+ Tile_X4Y1_LUT4AB/FrameStrobe[2] Tile_X4Y1_LUT4AB/FrameStrobe[3] Tile_X4Y1_LUT4AB/FrameStrobe[4]
+ Tile_X4Y1_LUT4AB/FrameStrobe[5] Tile_X4Y1_LUT4AB/FrameStrobe[6] Tile_X4Y1_LUT4AB/FrameStrobe[7]
+ Tile_X4Y1_LUT4AB/FrameStrobe[8] Tile_X4Y1_LUT4AB/FrameStrobe[9] Tile_X4Y2_LUT4AB/N1BEG[0]
+ Tile_X4Y2_LUT4AB/N1BEG[1] Tile_X4Y2_LUT4AB/N1BEG[2] Tile_X4Y2_LUT4AB/N1BEG[3] Tile_X4Y3_LUT4AB/N1BEG[0]
+ Tile_X4Y3_LUT4AB/N1BEG[1] Tile_X4Y3_LUT4AB/N1BEG[2] Tile_X4Y3_LUT4AB/N1BEG[3] Tile_X4Y2_LUT4AB/N2BEG[0]
+ Tile_X4Y2_LUT4AB/N2BEG[1] Tile_X4Y2_LUT4AB/N2BEG[2] Tile_X4Y2_LUT4AB/N2BEG[3] Tile_X4Y2_LUT4AB/N2BEG[4]
+ Tile_X4Y2_LUT4AB/N2BEG[5] Tile_X4Y2_LUT4AB/N2BEG[6] Tile_X4Y2_LUT4AB/N2BEG[7] Tile_X4Y1_LUT4AB/N2END[0]
+ Tile_X4Y1_LUT4AB/N2END[1] Tile_X4Y1_LUT4AB/N2END[2] Tile_X4Y1_LUT4AB/N2END[3] Tile_X4Y1_LUT4AB/N2END[4]
+ Tile_X4Y1_LUT4AB/N2END[5] Tile_X4Y1_LUT4AB/N2END[6] Tile_X4Y1_LUT4AB/N2END[7] Tile_X4Y2_LUT4AB/N2END[0]
+ Tile_X4Y2_LUT4AB/N2END[1] Tile_X4Y2_LUT4AB/N2END[2] Tile_X4Y2_LUT4AB/N2END[3] Tile_X4Y2_LUT4AB/N2END[4]
+ Tile_X4Y2_LUT4AB/N2END[5] Tile_X4Y2_LUT4AB/N2END[6] Tile_X4Y2_LUT4AB/N2END[7] Tile_X4Y3_LUT4AB/N2BEG[0]
+ Tile_X4Y3_LUT4AB/N2BEG[1] Tile_X4Y3_LUT4AB/N2BEG[2] Tile_X4Y3_LUT4AB/N2BEG[3] Tile_X4Y3_LUT4AB/N2BEG[4]
+ Tile_X4Y3_LUT4AB/N2BEG[5] Tile_X4Y3_LUT4AB/N2BEG[6] Tile_X4Y3_LUT4AB/N2BEG[7] Tile_X4Y2_LUT4AB/N4BEG[0]
+ Tile_X4Y2_LUT4AB/N4BEG[10] Tile_X4Y2_LUT4AB/N4BEG[11] Tile_X4Y2_LUT4AB/N4BEG[12]
+ Tile_X4Y2_LUT4AB/N4BEG[13] Tile_X4Y2_LUT4AB/N4BEG[14] Tile_X4Y2_LUT4AB/N4BEG[15]
+ Tile_X4Y2_LUT4AB/N4BEG[1] Tile_X4Y2_LUT4AB/N4BEG[2] Tile_X4Y2_LUT4AB/N4BEG[3] Tile_X4Y2_LUT4AB/N4BEG[4]
+ Tile_X4Y2_LUT4AB/N4BEG[5] Tile_X4Y2_LUT4AB/N4BEG[6] Tile_X4Y2_LUT4AB/N4BEG[7] Tile_X4Y2_LUT4AB/N4BEG[8]
+ Tile_X4Y2_LUT4AB/N4BEG[9] Tile_X4Y3_LUT4AB/N4BEG[0] Tile_X4Y3_LUT4AB/N4BEG[10] Tile_X4Y3_LUT4AB/N4BEG[11]
+ Tile_X4Y3_LUT4AB/N4BEG[12] Tile_X4Y3_LUT4AB/N4BEG[13] Tile_X4Y3_LUT4AB/N4BEG[14]
+ Tile_X4Y3_LUT4AB/N4BEG[15] Tile_X4Y3_LUT4AB/N4BEG[1] Tile_X4Y3_LUT4AB/N4BEG[2] Tile_X4Y3_LUT4AB/N4BEG[3]
+ Tile_X4Y3_LUT4AB/N4BEG[4] Tile_X4Y3_LUT4AB/N4BEG[5] Tile_X4Y3_LUT4AB/N4BEG[6] Tile_X4Y3_LUT4AB/N4BEG[7]
+ Tile_X4Y3_LUT4AB/N4BEG[8] Tile_X4Y3_LUT4AB/N4BEG[9] Tile_X4Y2_LUT4AB/NN4BEG[0] Tile_X4Y2_LUT4AB/NN4BEG[10]
+ Tile_X4Y2_LUT4AB/NN4BEG[11] Tile_X4Y2_LUT4AB/NN4BEG[12] Tile_X4Y2_LUT4AB/NN4BEG[13]
+ Tile_X4Y2_LUT4AB/NN4BEG[14] Tile_X4Y2_LUT4AB/NN4BEG[15] Tile_X4Y2_LUT4AB/NN4BEG[1]
+ Tile_X4Y2_LUT4AB/NN4BEG[2] Tile_X4Y2_LUT4AB/NN4BEG[3] Tile_X4Y2_LUT4AB/NN4BEG[4]
+ Tile_X4Y2_LUT4AB/NN4BEG[5] Tile_X4Y2_LUT4AB/NN4BEG[6] Tile_X4Y2_LUT4AB/NN4BEG[7]
+ Tile_X4Y2_LUT4AB/NN4BEG[8] Tile_X4Y2_LUT4AB/NN4BEG[9] Tile_X4Y3_LUT4AB/NN4BEG[0]
+ Tile_X4Y3_LUT4AB/NN4BEG[10] Tile_X4Y3_LUT4AB/NN4BEG[11] Tile_X4Y3_LUT4AB/NN4BEG[12]
+ Tile_X4Y3_LUT4AB/NN4BEG[13] Tile_X4Y3_LUT4AB/NN4BEG[14] Tile_X4Y3_LUT4AB/NN4BEG[15]
+ Tile_X4Y3_LUT4AB/NN4BEG[1] Tile_X4Y3_LUT4AB/NN4BEG[2] Tile_X4Y3_LUT4AB/NN4BEG[3]
+ Tile_X4Y3_LUT4AB/NN4BEG[4] Tile_X4Y3_LUT4AB/NN4BEG[5] Tile_X4Y3_LUT4AB/NN4BEG[6]
+ Tile_X4Y3_LUT4AB/NN4BEG[7] Tile_X4Y3_LUT4AB/NN4BEG[8] Tile_X4Y3_LUT4AB/NN4BEG[9]
+ Tile_X4Y3_LUT4AB/S1END[0] Tile_X4Y3_LUT4AB/S1END[1] Tile_X4Y3_LUT4AB/S1END[2] Tile_X4Y3_LUT4AB/S1END[3]
+ Tile_X4Y2_LUT4AB/S1END[0] Tile_X4Y2_LUT4AB/S1END[1] Tile_X4Y2_LUT4AB/S1END[2] Tile_X4Y2_LUT4AB/S1END[3]
+ Tile_X4Y3_LUT4AB/S2MID[0] Tile_X4Y3_LUT4AB/S2MID[1] Tile_X4Y3_LUT4AB/S2MID[2] Tile_X4Y3_LUT4AB/S2MID[3]
+ Tile_X4Y3_LUT4AB/S2MID[4] Tile_X4Y3_LUT4AB/S2MID[5] Tile_X4Y3_LUT4AB/S2MID[6] Tile_X4Y3_LUT4AB/S2MID[7]
+ Tile_X4Y3_LUT4AB/S2END[0] Tile_X4Y3_LUT4AB/S2END[1] Tile_X4Y3_LUT4AB/S2END[2] Tile_X4Y3_LUT4AB/S2END[3]
+ Tile_X4Y3_LUT4AB/S2END[4] Tile_X4Y3_LUT4AB/S2END[5] Tile_X4Y3_LUT4AB/S2END[6] Tile_X4Y3_LUT4AB/S2END[7]
+ Tile_X4Y2_LUT4AB/S2END[0] Tile_X4Y2_LUT4AB/S2END[1] Tile_X4Y2_LUT4AB/S2END[2] Tile_X4Y2_LUT4AB/S2END[3]
+ Tile_X4Y2_LUT4AB/S2END[4] Tile_X4Y2_LUT4AB/S2END[5] Tile_X4Y2_LUT4AB/S2END[6] Tile_X4Y2_LUT4AB/S2END[7]
+ Tile_X4Y2_LUT4AB/S2MID[0] Tile_X4Y2_LUT4AB/S2MID[1] Tile_X4Y2_LUT4AB/S2MID[2] Tile_X4Y2_LUT4AB/S2MID[3]
+ Tile_X4Y2_LUT4AB/S2MID[4] Tile_X4Y2_LUT4AB/S2MID[5] Tile_X4Y2_LUT4AB/S2MID[6] Tile_X4Y2_LUT4AB/S2MID[7]
+ Tile_X4Y3_LUT4AB/S4END[0] Tile_X4Y3_LUT4AB/S4END[10] Tile_X4Y3_LUT4AB/S4END[11]
+ Tile_X4Y3_LUT4AB/S4END[12] Tile_X4Y3_LUT4AB/S4END[13] Tile_X4Y3_LUT4AB/S4END[14]
+ Tile_X4Y3_LUT4AB/S4END[15] Tile_X4Y3_LUT4AB/S4END[1] Tile_X4Y3_LUT4AB/S4END[2] Tile_X4Y3_LUT4AB/S4END[3]
+ Tile_X4Y3_LUT4AB/S4END[4] Tile_X4Y3_LUT4AB/S4END[5] Tile_X4Y3_LUT4AB/S4END[6] Tile_X4Y3_LUT4AB/S4END[7]
+ Tile_X4Y3_LUT4AB/S4END[8] Tile_X4Y3_LUT4AB/S4END[9] Tile_X4Y2_LUT4AB/S4END[0] Tile_X4Y2_LUT4AB/S4END[10]
+ Tile_X4Y2_LUT4AB/S4END[11] Tile_X4Y2_LUT4AB/S4END[12] Tile_X4Y2_LUT4AB/S4END[13]
+ Tile_X4Y2_LUT4AB/S4END[14] Tile_X4Y2_LUT4AB/S4END[15] Tile_X4Y2_LUT4AB/S4END[1]
+ Tile_X4Y2_LUT4AB/S4END[2] Tile_X4Y2_LUT4AB/S4END[3] Tile_X4Y2_LUT4AB/S4END[4] Tile_X4Y2_LUT4AB/S4END[5]
+ Tile_X4Y2_LUT4AB/S4END[6] Tile_X4Y2_LUT4AB/S4END[7] Tile_X4Y2_LUT4AB/S4END[8] Tile_X4Y2_LUT4AB/S4END[9]
+ Tile_X4Y3_LUT4AB/SS4END[0] Tile_X4Y3_LUT4AB/SS4END[10] Tile_X4Y3_LUT4AB/SS4END[11]
+ Tile_X4Y3_LUT4AB/SS4END[12] Tile_X4Y3_LUT4AB/SS4END[13] Tile_X4Y3_LUT4AB/SS4END[14]
+ Tile_X4Y3_LUT4AB/SS4END[15] Tile_X4Y3_LUT4AB/SS4END[1] Tile_X4Y3_LUT4AB/SS4END[2]
+ Tile_X4Y3_LUT4AB/SS4END[3] Tile_X4Y3_LUT4AB/SS4END[4] Tile_X4Y3_LUT4AB/SS4END[5]
+ Tile_X4Y3_LUT4AB/SS4END[6] Tile_X4Y3_LUT4AB/SS4END[7] Tile_X4Y3_LUT4AB/SS4END[8]
+ Tile_X4Y3_LUT4AB/SS4END[9] Tile_X4Y2_LUT4AB/SS4END[0] Tile_X4Y2_LUT4AB/SS4END[10]
+ Tile_X4Y2_LUT4AB/SS4END[11] Tile_X4Y2_LUT4AB/SS4END[12] Tile_X4Y2_LUT4AB/SS4END[13]
+ Tile_X4Y2_LUT4AB/SS4END[14] Tile_X4Y2_LUT4AB/SS4END[15] Tile_X4Y2_LUT4AB/SS4END[1]
+ Tile_X4Y2_LUT4AB/SS4END[2] Tile_X4Y2_LUT4AB/SS4END[3] Tile_X4Y2_LUT4AB/SS4END[4]
+ Tile_X4Y2_LUT4AB/SS4END[5] Tile_X4Y2_LUT4AB/SS4END[6] Tile_X4Y2_LUT4AB/SS4END[7]
+ Tile_X4Y2_LUT4AB/SS4END[8] Tile_X4Y2_LUT4AB/SS4END[9] Tile_X4Y2_LUT4AB/UserCLK Tile_X4Y1_LUT4AB/UserCLK
+ VGND VPWR Tile_X4Y2_LUT4AB/W1BEG[0] Tile_X4Y2_LUT4AB/W1BEG[1] Tile_X4Y2_LUT4AB/W1BEG[2]
+ Tile_X4Y2_LUT4AB/W1BEG[3] Tile_X4Y2_LUT4AB/W1END[0] Tile_X4Y2_LUT4AB/W1END[1] Tile_X4Y2_LUT4AB/W1END[2]
+ Tile_X4Y2_LUT4AB/W1END[3] Tile_X4Y2_LUT4AB/W2BEG[0] Tile_X4Y2_LUT4AB/W2BEG[1] Tile_X4Y2_LUT4AB/W2BEG[2]
+ Tile_X4Y2_LUT4AB/W2BEG[3] Tile_X4Y2_LUT4AB/W2BEG[4] Tile_X4Y2_LUT4AB/W2BEG[5] Tile_X4Y2_LUT4AB/W2BEG[6]
+ Tile_X4Y2_LUT4AB/W2BEG[7] Tile_X3Y2_LUT4AB/W2END[0] Tile_X3Y2_LUT4AB/W2END[1] Tile_X3Y2_LUT4AB/W2END[2]
+ Tile_X3Y2_LUT4AB/W2END[3] Tile_X3Y2_LUT4AB/W2END[4] Tile_X3Y2_LUT4AB/W2END[5] Tile_X3Y2_LUT4AB/W2END[6]
+ Tile_X3Y2_LUT4AB/W2END[7] Tile_X4Y2_LUT4AB/W2END[0] Tile_X4Y2_LUT4AB/W2END[1] Tile_X4Y2_LUT4AB/W2END[2]
+ Tile_X4Y2_LUT4AB/W2END[3] Tile_X4Y2_LUT4AB/W2END[4] Tile_X4Y2_LUT4AB/W2END[5] Tile_X4Y2_LUT4AB/W2END[6]
+ Tile_X4Y2_LUT4AB/W2END[7] Tile_X4Y2_LUT4AB/W2MID[0] Tile_X4Y2_LUT4AB/W2MID[1] Tile_X4Y2_LUT4AB/W2MID[2]
+ Tile_X4Y2_LUT4AB/W2MID[3] Tile_X4Y2_LUT4AB/W2MID[4] Tile_X4Y2_LUT4AB/W2MID[5] Tile_X4Y2_LUT4AB/W2MID[6]
+ Tile_X4Y2_LUT4AB/W2MID[7] Tile_X4Y2_LUT4AB/W6BEG[0] Tile_X4Y2_LUT4AB/W6BEG[10] Tile_X4Y2_LUT4AB/W6BEG[11]
+ Tile_X4Y2_LUT4AB/W6BEG[1] Tile_X4Y2_LUT4AB/W6BEG[2] Tile_X4Y2_LUT4AB/W6BEG[3] Tile_X4Y2_LUT4AB/W6BEG[4]
+ Tile_X4Y2_LUT4AB/W6BEG[5] Tile_X4Y2_LUT4AB/W6BEG[6] Tile_X4Y2_LUT4AB/W6BEG[7] Tile_X4Y2_LUT4AB/W6BEG[8]
+ Tile_X4Y2_LUT4AB/W6BEG[9] Tile_X4Y2_LUT4AB/W6END[0] Tile_X4Y2_LUT4AB/W6END[10] Tile_X4Y2_LUT4AB/W6END[11]
+ Tile_X4Y2_LUT4AB/W6END[1] Tile_X4Y2_LUT4AB/W6END[2] Tile_X4Y2_LUT4AB/W6END[3] Tile_X4Y2_LUT4AB/W6END[4]
+ Tile_X4Y2_LUT4AB/W6END[5] Tile_X4Y2_LUT4AB/W6END[6] Tile_X4Y2_LUT4AB/W6END[7] Tile_X4Y2_LUT4AB/W6END[8]
+ Tile_X4Y2_LUT4AB/W6END[9] Tile_X4Y2_LUT4AB/WW4BEG[0] Tile_X4Y2_LUT4AB/WW4BEG[10]
+ Tile_X4Y2_LUT4AB/WW4BEG[11] Tile_X4Y2_LUT4AB/WW4BEG[12] Tile_X4Y2_LUT4AB/WW4BEG[13]
+ Tile_X4Y2_LUT4AB/WW4BEG[14] Tile_X4Y2_LUT4AB/WW4BEG[15] Tile_X4Y2_LUT4AB/WW4BEG[1]
+ Tile_X4Y2_LUT4AB/WW4BEG[2] Tile_X4Y2_LUT4AB/WW4BEG[3] Tile_X4Y2_LUT4AB/WW4BEG[4]
+ Tile_X4Y2_LUT4AB/WW4BEG[5] Tile_X4Y2_LUT4AB/WW4BEG[6] Tile_X4Y2_LUT4AB/WW4BEG[7]
+ Tile_X4Y2_LUT4AB/WW4BEG[8] Tile_X4Y2_LUT4AB/WW4BEG[9] Tile_X4Y2_LUT4AB/WW4END[0]
+ Tile_X4Y2_LUT4AB/WW4END[10] Tile_X4Y2_LUT4AB/WW4END[11] Tile_X4Y2_LUT4AB/WW4END[12]
+ Tile_X4Y2_LUT4AB/WW4END[13] Tile_X4Y2_LUT4AB/WW4END[14] Tile_X4Y2_LUT4AB/WW4END[15]
+ Tile_X4Y2_LUT4AB/WW4END[1] Tile_X4Y2_LUT4AB/WW4END[2] Tile_X4Y2_LUT4AB/WW4END[3]
+ Tile_X4Y2_LUT4AB/WW4END[4] Tile_X4Y2_LUT4AB/WW4END[5] Tile_X4Y2_LUT4AB/WW4END[6]
+ Tile_X4Y2_LUT4AB/WW4END[7] Tile_X4Y2_LUT4AB/WW4END[8] Tile_X4Y2_LUT4AB/WW4END[9]
+ LUT4AB
XTile_X0Y8_W_TT_IF Tile_X0Y8_CLK_TT_PROJECT Tile_X1Y8_LUT4AB/E1END[0] Tile_X1Y8_LUT4AB/E1END[1]
+ Tile_X1Y8_LUT4AB/E1END[2] Tile_X1Y8_LUT4AB/E1END[3] Tile_X1Y8_LUT4AB/E2MID[0] Tile_X1Y8_LUT4AB/E2MID[1]
+ Tile_X1Y8_LUT4AB/E2MID[2] Tile_X1Y8_LUT4AB/E2MID[3] Tile_X1Y8_LUT4AB/E2MID[4] Tile_X1Y8_LUT4AB/E2MID[5]
+ Tile_X1Y8_LUT4AB/E2MID[6] Tile_X1Y8_LUT4AB/E2MID[7] Tile_X1Y8_LUT4AB/E2END[0] Tile_X1Y8_LUT4AB/E2END[1]
+ Tile_X1Y8_LUT4AB/E2END[2] Tile_X1Y8_LUT4AB/E2END[3] Tile_X1Y8_LUT4AB/E2END[4] Tile_X1Y8_LUT4AB/E2END[5]
+ Tile_X1Y8_LUT4AB/E2END[6] Tile_X1Y8_LUT4AB/E2END[7] Tile_X1Y8_LUT4AB/E6END[0] Tile_X1Y8_LUT4AB/E6END[10]
+ Tile_X1Y8_LUT4AB/E6END[11] Tile_X1Y8_LUT4AB/E6END[1] Tile_X1Y8_LUT4AB/E6END[2] Tile_X1Y8_LUT4AB/E6END[3]
+ Tile_X1Y8_LUT4AB/E6END[4] Tile_X1Y8_LUT4AB/E6END[5] Tile_X1Y8_LUT4AB/E6END[6] Tile_X1Y8_LUT4AB/E6END[7]
+ Tile_X1Y8_LUT4AB/E6END[8] Tile_X1Y8_LUT4AB/E6END[9] Tile_X1Y8_LUT4AB/EE4END[0] Tile_X1Y8_LUT4AB/EE4END[10]
+ Tile_X1Y8_LUT4AB/EE4END[11] Tile_X1Y8_LUT4AB/EE4END[12] Tile_X1Y8_LUT4AB/EE4END[13]
+ Tile_X1Y8_LUT4AB/EE4END[14] Tile_X1Y8_LUT4AB/EE4END[15] Tile_X1Y8_LUT4AB/EE4END[1]
+ Tile_X1Y8_LUT4AB/EE4END[2] Tile_X1Y8_LUT4AB/EE4END[3] Tile_X1Y8_LUT4AB/EE4END[4]
+ Tile_X1Y8_LUT4AB/EE4END[5] Tile_X1Y8_LUT4AB/EE4END[6] Tile_X1Y8_LUT4AB/EE4END[7]
+ Tile_X1Y8_LUT4AB/EE4END[8] Tile_X1Y8_LUT4AB/EE4END[9] Tile_X0Y8_ENA_TT_PROJECT FrameData[256]
+ FrameData[266] FrameData[267] FrameData[268] FrameData[269] FrameData[270] FrameData[271]
+ FrameData[272] FrameData[273] FrameData[274] FrameData[275] FrameData[257] FrameData[276]
+ FrameData[277] FrameData[278] FrameData[279] FrameData[280] FrameData[281] FrameData[282]
+ FrameData[283] FrameData[284] FrameData[285] FrameData[258] FrameData[286] FrameData[287]
+ FrameData[259] FrameData[260] FrameData[261] FrameData[262] FrameData[263] FrameData[264]
+ FrameData[265] Tile_X1Y8_LUT4AB/FrameData[0] Tile_X1Y8_LUT4AB/FrameData[10] Tile_X1Y8_LUT4AB/FrameData[11]
+ Tile_X1Y8_LUT4AB/FrameData[12] Tile_X1Y8_LUT4AB/FrameData[13] Tile_X1Y8_LUT4AB/FrameData[14]
+ Tile_X1Y8_LUT4AB/FrameData[15] Tile_X1Y8_LUT4AB/FrameData[16] Tile_X1Y8_LUT4AB/FrameData[17]
+ Tile_X1Y8_LUT4AB/FrameData[18] Tile_X1Y8_LUT4AB/FrameData[19] Tile_X1Y8_LUT4AB/FrameData[1]
+ Tile_X1Y8_LUT4AB/FrameData[20] Tile_X1Y8_LUT4AB/FrameData[21] Tile_X1Y8_LUT4AB/FrameData[22]
+ Tile_X1Y8_LUT4AB/FrameData[23] Tile_X1Y8_LUT4AB/FrameData[24] Tile_X1Y8_LUT4AB/FrameData[25]
+ Tile_X1Y8_LUT4AB/FrameData[26] Tile_X1Y8_LUT4AB/FrameData[27] Tile_X1Y8_LUT4AB/FrameData[28]
+ Tile_X1Y8_LUT4AB/FrameData[29] Tile_X1Y8_LUT4AB/FrameData[2] Tile_X1Y8_LUT4AB/FrameData[30]
+ Tile_X1Y8_LUT4AB/FrameData[31] Tile_X1Y8_LUT4AB/FrameData[3] Tile_X1Y8_LUT4AB/FrameData[4]
+ Tile_X1Y8_LUT4AB/FrameData[5] Tile_X1Y8_LUT4AB/FrameData[6] Tile_X1Y8_LUT4AB/FrameData[7]
+ Tile_X1Y8_LUT4AB/FrameData[8] Tile_X1Y8_LUT4AB/FrameData[9] Tile_X0Y8_W_TT_IF/FrameStrobe[0]
+ Tile_X0Y8_W_TT_IF/FrameStrobe[10] Tile_X0Y8_W_TT_IF/FrameStrobe[11] Tile_X0Y8_W_TT_IF/FrameStrobe[12]
+ Tile_X0Y8_W_TT_IF/FrameStrobe[13] Tile_X0Y8_W_TT_IF/FrameStrobe[14] Tile_X0Y8_W_TT_IF/FrameStrobe[15]
+ Tile_X0Y8_W_TT_IF/FrameStrobe[16] Tile_X0Y8_W_TT_IF/FrameStrobe[17] Tile_X0Y8_W_TT_IF/FrameStrobe[18]
+ Tile_X0Y8_W_TT_IF/FrameStrobe[19] Tile_X0Y8_W_TT_IF/FrameStrobe[1] Tile_X0Y8_W_TT_IF/FrameStrobe[2]
+ Tile_X0Y8_W_TT_IF/FrameStrobe[3] Tile_X0Y8_W_TT_IF/FrameStrobe[4] Tile_X0Y8_W_TT_IF/FrameStrobe[5]
+ Tile_X0Y8_W_TT_IF/FrameStrobe[6] Tile_X0Y8_W_TT_IF/FrameStrobe[7] Tile_X0Y8_W_TT_IF/FrameStrobe[8]
+ Tile_X0Y8_W_TT_IF/FrameStrobe[9] Tile_X0Y7_W_TT_IF/FrameStrobe[0] Tile_X0Y7_W_TT_IF/FrameStrobe[10]
+ Tile_X0Y7_W_TT_IF/FrameStrobe[11] Tile_X0Y7_W_TT_IF/FrameStrobe[12] Tile_X0Y7_W_TT_IF/FrameStrobe[13]
+ Tile_X0Y7_W_TT_IF/FrameStrobe[14] Tile_X0Y7_W_TT_IF/FrameStrobe[15] Tile_X0Y7_W_TT_IF/FrameStrobe[16]
+ Tile_X0Y7_W_TT_IF/FrameStrobe[17] Tile_X0Y7_W_TT_IF/FrameStrobe[18] Tile_X0Y7_W_TT_IF/FrameStrobe[19]
+ Tile_X0Y7_W_TT_IF/FrameStrobe[1] Tile_X0Y7_W_TT_IF/FrameStrobe[2] Tile_X0Y7_W_TT_IF/FrameStrobe[3]
+ Tile_X0Y7_W_TT_IF/FrameStrobe[4] Tile_X0Y7_W_TT_IF/FrameStrobe[5] Tile_X0Y7_W_TT_IF/FrameStrobe[6]
+ Tile_X0Y7_W_TT_IF/FrameStrobe[7] Tile_X0Y7_W_TT_IF/FrameStrobe[8] Tile_X0Y7_W_TT_IF/FrameStrobe[9]
+ Tile_X0Y8_W_TT_IF/N1BEG[0] Tile_X0Y8_W_TT_IF/N1BEG[1] Tile_X0Y8_W_TT_IF/N1BEG[2]
+ Tile_X0Y8_W_TT_IF/N1BEG[3] Tile_X0Y9_SW_term/N1BEG[0] Tile_X0Y9_SW_term/N1BEG[1]
+ Tile_X0Y9_SW_term/N1BEG[2] Tile_X0Y9_SW_term/N1BEG[3] Tile_X0Y8_W_TT_IF/N2BEG[0]
+ Tile_X0Y8_W_TT_IF/N2BEG[1] Tile_X0Y8_W_TT_IF/N2BEG[2] Tile_X0Y8_W_TT_IF/N2BEG[3]
+ Tile_X0Y8_W_TT_IF/N2BEG[4] Tile_X0Y8_W_TT_IF/N2BEG[5] Tile_X0Y8_W_TT_IF/N2BEG[6]
+ Tile_X0Y8_W_TT_IF/N2BEG[7] Tile_X0Y7_W_TT_IF/N2END[0] Tile_X0Y7_W_TT_IF/N2END[1]
+ Tile_X0Y7_W_TT_IF/N2END[2] Tile_X0Y7_W_TT_IF/N2END[3] Tile_X0Y7_W_TT_IF/N2END[4]
+ Tile_X0Y7_W_TT_IF/N2END[5] Tile_X0Y7_W_TT_IF/N2END[6] Tile_X0Y7_W_TT_IF/N2END[7]
+ Tile_X0Y8_W_TT_IF/N2END[0] Tile_X0Y8_W_TT_IF/N2END[1] Tile_X0Y8_W_TT_IF/N2END[2]
+ Tile_X0Y8_W_TT_IF/N2END[3] Tile_X0Y8_W_TT_IF/N2END[4] Tile_X0Y8_W_TT_IF/N2END[5]
+ Tile_X0Y8_W_TT_IF/N2END[6] Tile_X0Y8_W_TT_IF/N2END[7] Tile_X0Y9_SW_term/N2BEG[0]
+ Tile_X0Y9_SW_term/N2BEG[1] Tile_X0Y9_SW_term/N2BEG[2] Tile_X0Y9_SW_term/N2BEG[3]
+ Tile_X0Y9_SW_term/N2BEG[4] Tile_X0Y9_SW_term/N2BEG[5] Tile_X0Y9_SW_term/N2BEG[6]
+ Tile_X0Y9_SW_term/N2BEG[7] Tile_X0Y8_W_TT_IF/N4BEG[0] Tile_X0Y8_W_TT_IF/N4BEG[10]
+ Tile_X0Y8_W_TT_IF/N4BEG[11] Tile_X0Y8_W_TT_IF/N4BEG[12] Tile_X0Y8_W_TT_IF/N4BEG[13]
+ Tile_X0Y8_W_TT_IF/N4BEG[14] Tile_X0Y8_W_TT_IF/N4BEG[15] Tile_X0Y8_W_TT_IF/N4BEG[1]
+ Tile_X0Y8_W_TT_IF/N4BEG[2] Tile_X0Y8_W_TT_IF/N4BEG[3] Tile_X0Y8_W_TT_IF/N4BEG[4]
+ Tile_X0Y8_W_TT_IF/N4BEG[5] Tile_X0Y8_W_TT_IF/N4BEG[6] Tile_X0Y8_W_TT_IF/N4BEG[7]
+ Tile_X0Y8_W_TT_IF/N4BEG[8] Tile_X0Y8_W_TT_IF/N4BEG[9] Tile_X0Y9_SW_term/N4BEG[0]
+ Tile_X0Y9_SW_term/N4BEG[10] Tile_X0Y9_SW_term/N4BEG[11] Tile_X0Y9_SW_term/N4BEG[12]
+ Tile_X0Y9_SW_term/N4BEG[13] Tile_X0Y9_SW_term/N4BEG[14] Tile_X0Y9_SW_term/N4BEG[15]
+ Tile_X0Y9_SW_term/N4BEG[1] Tile_X0Y9_SW_term/N4BEG[2] Tile_X0Y9_SW_term/N4BEG[3]
+ Tile_X0Y9_SW_term/N4BEG[4] Tile_X0Y9_SW_term/N4BEG[5] Tile_X0Y9_SW_term/N4BEG[6]
+ Tile_X0Y9_SW_term/N4BEG[7] Tile_X0Y9_SW_term/N4BEG[8] Tile_X0Y9_SW_term/N4BEG[9]
+ Tile_X0Y8_RST_N_TT_PROJECT Tile_X0Y9_SW_term/S1END[0] Tile_X0Y9_SW_term/S1END[1]
+ Tile_X0Y9_SW_term/S1END[2] Tile_X0Y9_SW_term/S1END[3] Tile_X0Y8_W_TT_IF/S1END[0]
+ Tile_X0Y8_W_TT_IF/S1END[1] Tile_X0Y8_W_TT_IF/S1END[2] Tile_X0Y8_W_TT_IF/S1END[3]
+ Tile_X0Y9_SW_term/S2MID[0] Tile_X0Y9_SW_term/S2MID[1] Tile_X0Y9_SW_term/S2MID[2]
+ Tile_X0Y9_SW_term/S2MID[3] Tile_X0Y9_SW_term/S2MID[4] Tile_X0Y9_SW_term/S2MID[5]
+ Tile_X0Y9_SW_term/S2MID[6] Tile_X0Y9_SW_term/S2MID[7] Tile_X0Y9_SW_term/S2END[0]
+ Tile_X0Y9_SW_term/S2END[1] Tile_X0Y9_SW_term/S2END[2] Tile_X0Y9_SW_term/S2END[3]
+ Tile_X0Y9_SW_term/S2END[4] Tile_X0Y9_SW_term/S2END[5] Tile_X0Y9_SW_term/S2END[6]
+ Tile_X0Y9_SW_term/S2END[7] Tile_X0Y8_W_TT_IF/S2END[0] Tile_X0Y8_W_TT_IF/S2END[1]
+ Tile_X0Y8_W_TT_IF/S2END[2] Tile_X0Y8_W_TT_IF/S2END[3] Tile_X0Y8_W_TT_IF/S2END[4]
+ Tile_X0Y8_W_TT_IF/S2END[5] Tile_X0Y8_W_TT_IF/S2END[6] Tile_X0Y8_W_TT_IF/S2END[7]
+ Tile_X0Y8_W_TT_IF/S2MID[0] Tile_X0Y8_W_TT_IF/S2MID[1] Tile_X0Y8_W_TT_IF/S2MID[2]
+ Tile_X0Y8_W_TT_IF/S2MID[3] Tile_X0Y8_W_TT_IF/S2MID[4] Tile_X0Y8_W_TT_IF/S2MID[5]
+ Tile_X0Y8_W_TT_IF/S2MID[6] Tile_X0Y8_W_TT_IF/S2MID[7] Tile_X0Y9_SW_term/S4END[0]
+ Tile_X0Y9_SW_term/S4END[10] Tile_X0Y9_SW_term/S4END[11] Tile_X0Y9_SW_term/S4END[12]
+ Tile_X0Y9_SW_term/S4END[13] Tile_X0Y9_SW_term/S4END[14] Tile_X0Y9_SW_term/S4END[15]
+ Tile_X0Y9_SW_term/S4END[1] Tile_X0Y9_SW_term/S4END[2] Tile_X0Y9_SW_term/S4END[3]
+ Tile_X0Y9_SW_term/S4END[4] Tile_X0Y9_SW_term/S4END[5] Tile_X0Y9_SW_term/S4END[6]
+ Tile_X0Y9_SW_term/S4END[7] Tile_X0Y9_SW_term/S4END[8] Tile_X0Y9_SW_term/S4END[9]
+ Tile_X0Y8_W_TT_IF/S4END[0] Tile_X0Y8_W_TT_IF/S4END[10] Tile_X0Y8_W_TT_IF/S4END[11]
+ Tile_X0Y8_W_TT_IF/S4END[12] Tile_X0Y8_W_TT_IF/S4END[13] Tile_X0Y8_W_TT_IF/S4END[14]
+ Tile_X0Y8_W_TT_IF/S4END[15] Tile_X0Y8_W_TT_IF/S4END[1] Tile_X0Y8_W_TT_IF/S4END[2]
+ Tile_X0Y8_W_TT_IF/S4END[3] Tile_X0Y8_W_TT_IF/S4END[4] Tile_X0Y8_W_TT_IF/S4END[5]
+ Tile_X0Y8_W_TT_IF/S4END[6] Tile_X0Y8_W_TT_IF/S4END[7] Tile_X0Y8_W_TT_IF/S4END[8]
+ Tile_X0Y8_W_TT_IF/S4END[9] Tile_X0Y8_UIO_IN_TT_PROJECT0 Tile_X0Y8_UIO_IN_TT_PROJECT1
+ Tile_X0Y8_UIO_IN_TT_PROJECT2 Tile_X0Y8_UIO_IN_TT_PROJECT3 Tile_X0Y8_UIO_IN_TT_PROJECT4
+ Tile_X0Y8_UIO_IN_TT_PROJECT5 Tile_X0Y8_UIO_IN_TT_PROJECT6 Tile_X0Y8_UIO_IN_TT_PROJECT7
+ Tile_X0Y8_UIO_OE_TT_PROJECT0 Tile_X0Y8_UIO_OE_TT_PROJECT1 Tile_X0Y8_UIO_OE_TT_PROJECT2
+ Tile_X0Y8_UIO_OE_TT_PROJECT3 Tile_X0Y8_UIO_OE_TT_PROJECT4 Tile_X0Y8_UIO_OE_TT_PROJECT5
+ Tile_X0Y8_UIO_OE_TT_PROJECT6 Tile_X0Y8_UIO_OE_TT_PROJECT7 Tile_X0Y8_UIO_OUT_TT_PROJECT0
+ Tile_X0Y8_UIO_OUT_TT_PROJECT1 Tile_X0Y8_UIO_OUT_TT_PROJECT2 Tile_X0Y8_UIO_OUT_TT_PROJECT3
+ Tile_X0Y8_UIO_OUT_TT_PROJECT4 Tile_X0Y8_UIO_OUT_TT_PROJECT5 Tile_X0Y8_UIO_OUT_TT_PROJECT6
+ Tile_X0Y8_UIO_OUT_TT_PROJECT7 Tile_X0Y8_UI_IN_TT_PROJECT0 Tile_X0Y8_UI_IN_TT_PROJECT1
+ Tile_X0Y8_UI_IN_TT_PROJECT2 Tile_X0Y8_UI_IN_TT_PROJECT3 Tile_X0Y8_UI_IN_TT_PROJECT4
+ Tile_X0Y8_UI_IN_TT_PROJECT5 Tile_X0Y8_UI_IN_TT_PROJECT6 Tile_X0Y8_UI_IN_TT_PROJECT7
+ Tile_X0Y8_UO_OUT_TT_PROJECT0 Tile_X0Y8_UO_OUT_TT_PROJECT1 Tile_X0Y8_UO_OUT_TT_PROJECT2
+ Tile_X0Y8_UO_OUT_TT_PROJECT3 Tile_X0Y8_UO_OUT_TT_PROJECT4 Tile_X0Y8_UO_OUT_TT_PROJECT5
+ Tile_X0Y8_UO_OUT_TT_PROJECT6 Tile_X0Y8_UO_OUT_TT_PROJECT7 Tile_X0Y8_W_TT_IF/UserCLK
+ Tile_X0Y7_W_TT_IF/UserCLK VGND VPWR Tile_X1Y8_LUT4AB/W1BEG[0] Tile_X1Y8_LUT4AB/W1BEG[1]
+ Tile_X1Y8_LUT4AB/W1BEG[2] Tile_X1Y8_LUT4AB/W1BEG[3] Tile_X1Y8_LUT4AB/W2BEGb[0] Tile_X1Y8_LUT4AB/W2BEGb[1]
+ Tile_X1Y8_LUT4AB/W2BEGb[2] Tile_X1Y8_LUT4AB/W2BEGb[3] Tile_X1Y8_LUT4AB/W2BEGb[4]
+ Tile_X1Y8_LUT4AB/W2BEGb[5] Tile_X1Y8_LUT4AB/W2BEGb[6] Tile_X1Y8_LUT4AB/W2BEGb[7]
+ Tile_X1Y8_LUT4AB/W2BEG[0] Tile_X1Y8_LUT4AB/W2BEG[1] Tile_X1Y8_LUT4AB/W2BEG[2] Tile_X1Y8_LUT4AB/W2BEG[3]
+ Tile_X1Y8_LUT4AB/W2BEG[4] Tile_X1Y8_LUT4AB/W2BEG[5] Tile_X1Y8_LUT4AB/W2BEG[6] Tile_X1Y8_LUT4AB/W2BEG[7]
+ Tile_X1Y8_LUT4AB/W6BEG[0] Tile_X1Y8_LUT4AB/W6BEG[10] Tile_X1Y8_LUT4AB/W6BEG[11]
+ Tile_X1Y8_LUT4AB/W6BEG[1] Tile_X1Y8_LUT4AB/W6BEG[2] Tile_X1Y8_LUT4AB/W6BEG[3] Tile_X1Y8_LUT4AB/W6BEG[4]
+ Tile_X1Y8_LUT4AB/W6BEG[5] Tile_X1Y8_LUT4AB/W6BEG[6] Tile_X1Y8_LUT4AB/W6BEG[7] Tile_X1Y8_LUT4AB/W6BEG[8]
+ Tile_X1Y8_LUT4AB/W6BEG[9] Tile_X1Y8_LUT4AB/WW4BEG[0] Tile_X1Y8_LUT4AB/WW4BEG[10]
+ Tile_X1Y8_LUT4AB/WW4BEG[11] Tile_X1Y8_LUT4AB/WW4BEG[12] Tile_X1Y8_LUT4AB/WW4BEG[13]
+ Tile_X1Y8_LUT4AB/WW4BEG[14] Tile_X1Y8_LUT4AB/WW4BEG[15] Tile_X1Y8_LUT4AB/WW4BEG[1]
+ Tile_X1Y8_LUT4AB/WW4BEG[2] Tile_X1Y8_LUT4AB/WW4BEG[3] Tile_X1Y8_LUT4AB/WW4BEG[4]
+ Tile_X1Y8_LUT4AB/WW4BEG[5] Tile_X1Y8_LUT4AB/WW4BEG[6] Tile_X1Y8_LUT4AB/WW4BEG[7]
+ Tile_X1Y8_LUT4AB/WW4BEG[8] Tile_X1Y8_LUT4AB/WW4BEG[9] W_TT_IF
XTile_X0Y4_W_TT_IF Tile_X0Y4_CLK_TT_PROJECT Tile_X1Y4_LUT4AB/E1END[0] Tile_X1Y4_LUT4AB/E1END[1]
+ Tile_X1Y4_LUT4AB/E1END[2] Tile_X1Y4_LUT4AB/E1END[3] Tile_X1Y4_LUT4AB/E2MID[0] Tile_X1Y4_LUT4AB/E2MID[1]
+ Tile_X1Y4_LUT4AB/E2MID[2] Tile_X1Y4_LUT4AB/E2MID[3] Tile_X1Y4_LUT4AB/E2MID[4] Tile_X1Y4_LUT4AB/E2MID[5]
+ Tile_X1Y4_LUT4AB/E2MID[6] Tile_X1Y4_LUT4AB/E2MID[7] Tile_X1Y4_LUT4AB/E2END[0] Tile_X1Y4_LUT4AB/E2END[1]
+ Tile_X1Y4_LUT4AB/E2END[2] Tile_X1Y4_LUT4AB/E2END[3] Tile_X1Y4_LUT4AB/E2END[4] Tile_X1Y4_LUT4AB/E2END[5]
+ Tile_X1Y4_LUT4AB/E2END[6] Tile_X1Y4_LUT4AB/E2END[7] Tile_X1Y4_LUT4AB/E6END[0] Tile_X1Y4_LUT4AB/E6END[10]
+ Tile_X1Y4_LUT4AB/E6END[11] Tile_X1Y4_LUT4AB/E6END[1] Tile_X1Y4_LUT4AB/E6END[2] Tile_X1Y4_LUT4AB/E6END[3]
+ Tile_X1Y4_LUT4AB/E6END[4] Tile_X1Y4_LUT4AB/E6END[5] Tile_X1Y4_LUT4AB/E6END[6] Tile_X1Y4_LUT4AB/E6END[7]
+ Tile_X1Y4_LUT4AB/E6END[8] Tile_X1Y4_LUT4AB/E6END[9] Tile_X1Y4_LUT4AB/EE4END[0] Tile_X1Y4_LUT4AB/EE4END[10]
+ Tile_X1Y4_LUT4AB/EE4END[11] Tile_X1Y4_LUT4AB/EE4END[12] Tile_X1Y4_LUT4AB/EE4END[13]
+ Tile_X1Y4_LUT4AB/EE4END[14] Tile_X1Y4_LUT4AB/EE4END[15] Tile_X1Y4_LUT4AB/EE4END[1]
+ Tile_X1Y4_LUT4AB/EE4END[2] Tile_X1Y4_LUT4AB/EE4END[3] Tile_X1Y4_LUT4AB/EE4END[4]
+ Tile_X1Y4_LUT4AB/EE4END[5] Tile_X1Y4_LUT4AB/EE4END[6] Tile_X1Y4_LUT4AB/EE4END[7]
+ Tile_X1Y4_LUT4AB/EE4END[8] Tile_X1Y4_LUT4AB/EE4END[9] Tile_X0Y4_ENA_TT_PROJECT FrameData[128]
+ FrameData[138] FrameData[139] FrameData[140] FrameData[141] FrameData[142] FrameData[143]
+ FrameData[144] FrameData[145] FrameData[146] FrameData[147] FrameData[129] FrameData[148]
+ FrameData[149] FrameData[150] FrameData[151] FrameData[152] FrameData[153] FrameData[154]
+ FrameData[155] FrameData[156] FrameData[157] FrameData[130] FrameData[158] FrameData[159]
+ FrameData[131] FrameData[132] FrameData[133] FrameData[134] FrameData[135] FrameData[136]
+ FrameData[137] Tile_X1Y4_LUT4AB/FrameData[0] Tile_X1Y4_LUT4AB/FrameData[10] Tile_X1Y4_LUT4AB/FrameData[11]
+ Tile_X1Y4_LUT4AB/FrameData[12] Tile_X1Y4_LUT4AB/FrameData[13] Tile_X1Y4_LUT4AB/FrameData[14]
+ Tile_X1Y4_LUT4AB/FrameData[15] Tile_X1Y4_LUT4AB/FrameData[16] Tile_X1Y4_LUT4AB/FrameData[17]
+ Tile_X1Y4_LUT4AB/FrameData[18] Tile_X1Y4_LUT4AB/FrameData[19] Tile_X1Y4_LUT4AB/FrameData[1]
+ Tile_X1Y4_LUT4AB/FrameData[20] Tile_X1Y4_LUT4AB/FrameData[21] Tile_X1Y4_LUT4AB/FrameData[22]
+ Tile_X1Y4_LUT4AB/FrameData[23] Tile_X1Y4_LUT4AB/FrameData[24] Tile_X1Y4_LUT4AB/FrameData[25]
+ Tile_X1Y4_LUT4AB/FrameData[26] Tile_X1Y4_LUT4AB/FrameData[27] Tile_X1Y4_LUT4AB/FrameData[28]
+ Tile_X1Y4_LUT4AB/FrameData[29] Tile_X1Y4_LUT4AB/FrameData[2] Tile_X1Y4_LUT4AB/FrameData[30]
+ Tile_X1Y4_LUT4AB/FrameData[31] Tile_X1Y4_LUT4AB/FrameData[3] Tile_X1Y4_LUT4AB/FrameData[4]
+ Tile_X1Y4_LUT4AB/FrameData[5] Tile_X1Y4_LUT4AB/FrameData[6] Tile_X1Y4_LUT4AB/FrameData[7]
+ Tile_X1Y4_LUT4AB/FrameData[8] Tile_X1Y4_LUT4AB/FrameData[9] Tile_X0Y4_W_TT_IF/FrameStrobe[0]
+ Tile_X0Y4_W_TT_IF/FrameStrobe[10] Tile_X0Y4_W_TT_IF/FrameStrobe[11] Tile_X0Y4_W_TT_IF/FrameStrobe[12]
+ Tile_X0Y4_W_TT_IF/FrameStrobe[13] Tile_X0Y4_W_TT_IF/FrameStrobe[14] Tile_X0Y4_W_TT_IF/FrameStrobe[15]
+ Tile_X0Y4_W_TT_IF/FrameStrobe[16] Tile_X0Y4_W_TT_IF/FrameStrobe[17] Tile_X0Y4_W_TT_IF/FrameStrobe[18]
+ Tile_X0Y4_W_TT_IF/FrameStrobe[19] Tile_X0Y4_W_TT_IF/FrameStrobe[1] Tile_X0Y4_W_TT_IF/FrameStrobe[2]
+ Tile_X0Y4_W_TT_IF/FrameStrobe[3] Tile_X0Y4_W_TT_IF/FrameStrobe[4] Tile_X0Y4_W_TT_IF/FrameStrobe[5]
+ Tile_X0Y4_W_TT_IF/FrameStrobe[6] Tile_X0Y4_W_TT_IF/FrameStrobe[7] Tile_X0Y4_W_TT_IF/FrameStrobe[8]
+ Tile_X0Y4_W_TT_IF/FrameStrobe[9] Tile_X0Y3_W_TT_IF/FrameStrobe[0] Tile_X0Y3_W_TT_IF/FrameStrobe[10]
+ Tile_X0Y3_W_TT_IF/FrameStrobe[11] Tile_X0Y3_W_TT_IF/FrameStrobe[12] Tile_X0Y3_W_TT_IF/FrameStrobe[13]
+ Tile_X0Y3_W_TT_IF/FrameStrobe[14] Tile_X0Y3_W_TT_IF/FrameStrobe[15] Tile_X0Y3_W_TT_IF/FrameStrobe[16]
+ Tile_X0Y3_W_TT_IF/FrameStrobe[17] Tile_X0Y3_W_TT_IF/FrameStrobe[18] Tile_X0Y3_W_TT_IF/FrameStrobe[19]
+ Tile_X0Y3_W_TT_IF/FrameStrobe[1] Tile_X0Y3_W_TT_IF/FrameStrobe[2] Tile_X0Y3_W_TT_IF/FrameStrobe[3]
+ Tile_X0Y3_W_TT_IF/FrameStrobe[4] Tile_X0Y3_W_TT_IF/FrameStrobe[5] Tile_X0Y3_W_TT_IF/FrameStrobe[6]
+ Tile_X0Y3_W_TT_IF/FrameStrobe[7] Tile_X0Y3_W_TT_IF/FrameStrobe[8] Tile_X0Y3_W_TT_IF/FrameStrobe[9]
+ Tile_X0Y4_W_TT_IF/N1BEG[0] Tile_X0Y4_W_TT_IF/N1BEG[1] Tile_X0Y4_W_TT_IF/N1BEG[2]
+ Tile_X0Y4_W_TT_IF/N1BEG[3] Tile_X0Y5_W_TT_IF/N1BEG[0] Tile_X0Y5_W_TT_IF/N1BEG[1]
+ Tile_X0Y5_W_TT_IF/N1BEG[2] Tile_X0Y5_W_TT_IF/N1BEG[3] Tile_X0Y4_W_TT_IF/N2BEG[0]
+ Tile_X0Y4_W_TT_IF/N2BEG[1] Tile_X0Y4_W_TT_IF/N2BEG[2] Tile_X0Y4_W_TT_IF/N2BEG[3]
+ Tile_X0Y4_W_TT_IF/N2BEG[4] Tile_X0Y4_W_TT_IF/N2BEG[5] Tile_X0Y4_W_TT_IF/N2BEG[6]
+ Tile_X0Y4_W_TT_IF/N2BEG[7] Tile_X0Y3_W_TT_IF/N2END[0] Tile_X0Y3_W_TT_IF/N2END[1]
+ Tile_X0Y3_W_TT_IF/N2END[2] Tile_X0Y3_W_TT_IF/N2END[3] Tile_X0Y3_W_TT_IF/N2END[4]
+ Tile_X0Y3_W_TT_IF/N2END[5] Tile_X0Y3_W_TT_IF/N2END[6] Tile_X0Y3_W_TT_IF/N2END[7]
+ Tile_X0Y4_W_TT_IF/N2END[0] Tile_X0Y4_W_TT_IF/N2END[1] Tile_X0Y4_W_TT_IF/N2END[2]
+ Tile_X0Y4_W_TT_IF/N2END[3] Tile_X0Y4_W_TT_IF/N2END[4] Tile_X0Y4_W_TT_IF/N2END[5]
+ Tile_X0Y4_W_TT_IF/N2END[6] Tile_X0Y4_W_TT_IF/N2END[7] Tile_X0Y5_W_TT_IF/N2BEG[0]
+ Tile_X0Y5_W_TT_IF/N2BEG[1] Tile_X0Y5_W_TT_IF/N2BEG[2] Tile_X0Y5_W_TT_IF/N2BEG[3]
+ Tile_X0Y5_W_TT_IF/N2BEG[4] Tile_X0Y5_W_TT_IF/N2BEG[5] Tile_X0Y5_W_TT_IF/N2BEG[6]
+ Tile_X0Y5_W_TT_IF/N2BEG[7] Tile_X0Y4_W_TT_IF/N4BEG[0] Tile_X0Y4_W_TT_IF/N4BEG[10]
+ Tile_X0Y4_W_TT_IF/N4BEG[11] Tile_X0Y4_W_TT_IF/N4BEG[12] Tile_X0Y4_W_TT_IF/N4BEG[13]
+ Tile_X0Y4_W_TT_IF/N4BEG[14] Tile_X0Y4_W_TT_IF/N4BEG[15] Tile_X0Y4_W_TT_IF/N4BEG[1]
+ Tile_X0Y4_W_TT_IF/N4BEG[2] Tile_X0Y4_W_TT_IF/N4BEG[3] Tile_X0Y4_W_TT_IF/N4BEG[4]
+ Tile_X0Y4_W_TT_IF/N4BEG[5] Tile_X0Y4_W_TT_IF/N4BEG[6] Tile_X0Y4_W_TT_IF/N4BEG[7]
+ Tile_X0Y4_W_TT_IF/N4BEG[8] Tile_X0Y4_W_TT_IF/N4BEG[9] Tile_X0Y5_W_TT_IF/N4BEG[0]
+ Tile_X0Y5_W_TT_IF/N4BEG[10] Tile_X0Y5_W_TT_IF/N4BEG[11] Tile_X0Y5_W_TT_IF/N4BEG[12]
+ Tile_X0Y5_W_TT_IF/N4BEG[13] Tile_X0Y5_W_TT_IF/N4BEG[14] Tile_X0Y5_W_TT_IF/N4BEG[15]
+ Tile_X0Y5_W_TT_IF/N4BEG[1] Tile_X0Y5_W_TT_IF/N4BEG[2] Tile_X0Y5_W_TT_IF/N4BEG[3]
+ Tile_X0Y5_W_TT_IF/N4BEG[4] Tile_X0Y5_W_TT_IF/N4BEG[5] Tile_X0Y5_W_TT_IF/N4BEG[6]
+ Tile_X0Y5_W_TT_IF/N4BEG[7] Tile_X0Y5_W_TT_IF/N4BEG[8] Tile_X0Y5_W_TT_IF/N4BEG[9]
+ Tile_X0Y4_RST_N_TT_PROJECT Tile_X0Y5_W_TT_IF/S1END[0] Tile_X0Y5_W_TT_IF/S1END[1]
+ Tile_X0Y5_W_TT_IF/S1END[2] Tile_X0Y5_W_TT_IF/S1END[3] Tile_X0Y4_W_TT_IF/S1END[0]
+ Tile_X0Y4_W_TT_IF/S1END[1] Tile_X0Y4_W_TT_IF/S1END[2] Tile_X0Y4_W_TT_IF/S1END[3]
+ Tile_X0Y5_W_TT_IF/S2MID[0] Tile_X0Y5_W_TT_IF/S2MID[1] Tile_X0Y5_W_TT_IF/S2MID[2]
+ Tile_X0Y5_W_TT_IF/S2MID[3] Tile_X0Y5_W_TT_IF/S2MID[4] Tile_X0Y5_W_TT_IF/S2MID[5]
+ Tile_X0Y5_W_TT_IF/S2MID[6] Tile_X0Y5_W_TT_IF/S2MID[7] Tile_X0Y5_W_TT_IF/S2END[0]
+ Tile_X0Y5_W_TT_IF/S2END[1] Tile_X0Y5_W_TT_IF/S2END[2] Tile_X0Y5_W_TT_IF/S2END[3]
+ Tile_X0Y5_W_TT_IF/S2END[4] Tile_X0Y5_W_TT_IF/S2END[5] Tile_X0Y5_W_TT_IF/S2END[6]
+ Tile_X0Y5_W_TT_IF/S2END[7] Tile_X0Y4_W_TT_IF/S2END[0] Tile_X0Y4_W_TT_IF/S2END[1]
+ Tile_X0Y4_W_TT_IF/S2END[2] Tile_X0Y4_W_TT_IF/S2END[3] Tile_X0Y4_W_TT_IF/S2END[4]
+ Tile_X0Y4_W_TT_IF/S2END[5] Tile_X0Y4_W_TT_IF/S2END[6] Tile_X0Y4_W_TT_IF/S2END[7]
+ Tile_X0Y4_W_TT_IF/S2MID[0] Tile_X0Y4_W_TT_IF/S2MID[1] Tile_X0Y4_W_TT_IF/S2MID[2]
+ Tile_X0Y4_W_TT_IF/S2MID[3] Tile_X0Y4_W_TT_IF/S2MID[4] Tile_X0Y4_W_TT_IF/S2MID[5]
+ Tile_X0Y4_W_TT_IF/S2MID[6] Tile_X0Y4_W_TT_IF/S2MID[7] Tile_X0Y5_W_TT_IF/S4END[0]
+ Tile_X0Y5_W_TT_IF/S4END[10] Tile_X0Y5_W_TT_IF/S4END[11] Tile_X0Y5_W_TT_IF/S4END[12]
+ Tile_X0Y5_W_TT_IF/S4END[13] Tile_X0Y5_W_TT_IF/S4END[14] Tile_X0Y5_W_TT_IF/S4END[15]
+ Tile_X0Y5_W_TT_IF/S4END[1] Tile_X0Y5_W_TT_IF/S4END[2] Tile_X0Y5_W_TT_IF/S4END[3]
+ Tile_X0Y5_W_TT_IF/S4END[4] Tile_X0Y5_W_TT_IF/S4END[5] Tile_X0Y5_W_TT_IF/S4END[6]
+ Tile_X0Y5_W_TT_IF/S4END[7] Tile_X0Y5_W_TT_IF/S4END[8] Tile_X0Y5_W_TT_IF/S4END[9]
+ Tile_X0Y4_W_TT_IF/S4END[0] Tile_X0Y4_W_TT_IF/S4END[10] Tile_X0Y4_W_TT_IF/S4END[11]
+ Tile_X0Y4_W_TT_IF/S4END[12] Tile_X0Y4_W_TT_IF/S4END[13] Tile_X0Y4_W_TT_IF/S4END[14]
+ Tile_X0Y4_W_TT_IF/S4END[15] Tile_X0Y4_W_TT_IF/S4END[1] Tile_X0Y4_W_TT_IF/S4END[2]
+ Tile_X0Y4_W_TT_IF/S4END[3] Tile_X0Y4_W_TT_IF/S4END[4] Tile_X0Y4_W_TT_IF/S4END[5]
+ Tile_X0Y4_W_TT_IF/S4END[6] Tile_X0Y4_W_TT_IF/S4END[7] Tile_X0Y4_W_TT_IF/S4END[8]
+ Tile_X0Y4_W_TT_IF/S4END[9] Tile_X0Y4_UIO_IN_TT_PROJECT0 Tile_X0Y4_UIO_IN_TT_PROJECT1
+ Tile_X0Y4_UIO_IN_TT_PROJECT2 Tile_X0Y4_UIO_IN_TT_PROJECT3 Tile_X0Y4_UIO_IN_TT_PROJECT4
+ Tile_X0Y4_UIO_IN_TT_PROJECT5 Tile_X0Y4_UIO_IN_TT_PROJECT6 Tile_X0Y4_UIO_IN_TT_PROJECT7
+ Tile_X0Y4_UIO_OE_TT_PROJECT0 Tile_X0Y4_UIO_OE_TT_PROJECT1 Tile_X0Y4_UIO_OE_TT_PROJECT2
+ Tile_X0Y4_UIO_OE_TT_PROJECT3 Tile_X0Y4_UIO_OE_TT_PROJECT4 Tile_X0Y4_UIO_OE_TT_PROJECT5
+ Tile_X0Y4_UIO_OE_TT_PROJECT6 Tile_X0Y4_UIO_OE_TT_PROJECT7 Tile_X0Y4_UIO_OUT_TT_PROJECT0
+ Tile_X0Y4_UIO_OUT_TT_PROJECT1 Tile_X0Y4_UIO_OUT_TT_PROJECT2 Tile_X0Y4_UIO_OUT_TT_PROJECT3
+ Tile_X0Y4_UIO_OUT_TT_PROJECT4 Tile_X0Y4_UIO_OUT_TT_PROJECT5 Tile_X0Y4_UIO_OUT_TT_PROJECT6
+ Tile_X0Y4_UIO_OUT_TT_PROJECT7 Tile_X0Y4_UI_IN_TT_PROJECT0 Tile_X0Y4_UI_IN_TT_PROJECT1
+ Tile_X0Y4_UI_IN_TT_PROJECT2 Tile_X0Y4_UI_IN_TT_PROJECT3 Tile_X0Y4_UI_IN_TT_PROJECT4
+ Tile_X0Y4_UI_IN_TT_PROJECT5 Tile_X0Y4_UI_IN_TT_PROJECT6 Tile_X0Y4_UI_IN_TT_PROJECT7
+ Tile_X0Y4_UO_OUT_TT_PROJECT0 Tile_X0Y4_UO_OUT_TT_PROJECT1 Tile_X0Y4_UO_OUT_TT_PROJECT2
+ Tile_X0Y4_UO_OUT_TT_PROJECT3 Tile_X0Y4_UO_OUT_TT_PROJECT4 Tile_X0Y4_UO_OUT_TT_PROJECT5
+ Tile_X0Y4_UO_OUT_TT_PROJECT6 Tile_X0Y4_UO_OUT_TT_PROJECT7 Tile_X0Y4_W_TT_IF/UserCLK
+ Tile_X0Y3_W_TT_IF/UserCLK VGND VPWR Tile_X1Y4_LUT4AB/W1BEG[0] Tile_X1Y4_LUT4AB/W1BEG[1]
+ Tile_X1Y4_LUT4AB/W1BEG[2] Tile_X1Y4_LUT4AB/W1BEG[3] Tile_X1Y4_LUT4AB/W2BEGb[0] Tile_X1Y4_LUT4AB/W2BEGb[1]
+ Tile_X1Y4_LUT4AB/W2BEGb[2] Tile_X1Y4_LUT4AB/W2BEGb[3] Tile_X1Y4_LUT4AB/W2BEGb[4]
+ Tile_X1Y4_LUT4AB/W2BEGb[5] Tile_X1Y4_LUT4AB/W2BEGb[6] Tile_X1Y4_LUT4AB/W2BEGb[7]
+ Tile_X1Y4_LUT4AB/W2BEG[0] Tile_X1Y4_LUT4AB/W2BEG[1] Tile_X1Y4_LUT4AB/W2BEG[2] Tile_X1Y4_LUT4AB/W2BEG[3]
+ Tile_X1Y4_LUT4AB/W2BEG[4] Tile_X1Y4_LUT4AB/W2BEG[5] Tile_X1Y4_LUT4AB/W2BEG[6] Tile_X1Y4_LUT4AB/W2BEG[7]
+ Tile_X1Y4_LUT4AB/W6BEG[0] Tile_X1Y4_LUT4AB/W6BEG[10] Tile_X1Y4_LUT4AB/W6BEG[11]
+ Tile_X1Y4_LUT4AB/W6BEG[1] Tile_X1Y4_LUT4AB/W6BEG[2] Tile_X1Y4_LUT4AB/W6BEG[3] Tile_X1Y4_LUT4AB/W6BEG[4]
+ Tile_X1Y4_LUT4AB/W6BEG[5] Tile_X1Y4_LUT4AB/W6BEG[6] Tile_X1Y4_LUT4AB/W6BEG[7] Tile_X1Y4_LUT4AB/W6BEG[8]
+ Tile_X1Y4_LUT4AB/W6BEG[9] Tile_X1Y4_LUT4AB/WW4BEG[0] Tile_X1Y4_LUT4AB/WW4BEG[10]
+ Tile_X1Y4_LUT4AB/WW4BEG[11] Tile_X1Y4_LUT4AB/WW4BEG[12] Tile_X1Y4_LUT4AB/WW4BEG[13]
+ Tile_X1Y4_LUT4AB/WW4BEG[14] Tile_X1Y4_LUT4AB/WW4BEG[15] Tile_X1Y4_LUT4AB/WW4BEG[1]
+ Tile_X1Y4_LUT4AB/WW4BEG[2] Tile_X1Y4_LUT4AB/WW4BEG[3] Tile_X1Y4_LUT4AB/WW4BEG[4]
+ Tile_X1Y4_LUT4AB/WW4BEG[5] Tile_X1Y4_LUT4AB/WW4BEG[6] Tile_X1Y4_LUT4AB/WW4BEG[7]
+ Tile_X1Y4_LUT4AB/WW4BEG[8] Tile_X1Y4_LUT4AB/WW4BEG[9] W_TT_IF
XTile_X3Y6_LUT4AB Tile_X3Y7_LUT4AB/Co Tile_X3Y6_LUT4AB/Co Tile_X4Y6_LUT4AB/E1END[0]
+ Tile_X4Y6_LUT4AB/E1END[1] Tile_X4Y6_LUT4AB/E1END[2] Tile_X4Y6_LUT4AB/E1END[3] Tile_X3Y6_LUT4AB/E1END[0]
+ Tile_X3Y6_LUT4AB/E1END[1] Tile_X3Y6_LUT4AB/E1END[2] Tile_X3Y6_LUT4AB/E1END[3] Tile_X4Y6_LUT4AB/E2MID[0]
+ Tile_X4Y6_LUT4AB/E2MID[1] Tile_X4Y6_LUT4AB/E2MID[2] Tile_X4Y6_LUT4AB/E2MID[3] Tile_X4Y6_LUT4AB/E2MID[4]
+ Tile_X4Y6_LUT4AB/E2MID[5] Tile_X4Y6_LUT4AB/E2MID[6] Tile_X4Y6_LUT4AB/E2MID[7] Tile_X4Y6_LUT4AB/E2END[0]
+ Tile_X4Y6_LUT4AB/E2END[1] Tile_X4Y6_LUT4AB/E2END[2] Tile_X4Y6_LUT4AB/E2END[3] Tile_X4Y6_LUT4AB/E2END[4]
+ Tile_X4Y6_LUT4AB/E2END[5] Tile_X4Y6_LUT4AB/E2END[6] Tile_X4Y6_LUT4AB/E2END[7] Tile_X3Y6_LUT4AB/E2END[0]
+ Tile_X3Y6_LUT4AB/E2END[1] Tile_X3Y6_LUT4AB/E2END[2] Tile_X3Y6_LUT4AB/E2END[3] Tile_X3Y6_LUT4AB/E2END[4]
+ Tile_X3Y6_LUT4AB/E2END[5] Tile_X3Y6_LUT4AB/E2END[6] Tile_X3Y6_LUT4AB/E2END[7] Tile_X3Y6_LUT4AB/E2MID[0]
+ Tile_X3Y6_LUT4AB/E2MID[1] Tile_X3Y6_LUT4AB/E2MID[2] Tile_X3Y6_LUT4AB/E2MID[3] Tile_X3Y6_LUT4AB/E2MID[4]
+ Tile_X3Y6_LUT4AB/E2MID[5] Tile_X3Y6_LUT4AB/E2MID[6] Tile_X3Y6_LUT4AB/E2MID[7] Tile_X4Y6_LUT4AB/E6END[0]
+ Tile_X4Y6_LUT4AB/E6END[10] Tile_X4Y6_LUT4AB/E6END[11] Tile_X4Y6_LUT4AB/E6END[1]
+ Tile_X4Y6_LUT4AB/E6END[2] Tile_X4Y6_LUT4AB/E6END[3] Tile_X4Y6_LUT4AB/E6END[4] Tile_X4Y6_LUT4AB/E6END[5]
+ Tile_X4Y6_LUT4AB/E6END[6] Tile_X4Y6_LUT4AB/E6END[7] Tile_X4Y6_LUT4AB/E6END[8] Tile_X4Y6_LUT4AB/E6END[9]
+ Tile_X3Y6_LUT4AB/E6END[0] Tile_X3Y6_LUT4AB/E6END[10] Tile_X3Y6_LUT4AB/E6END[11]
+ Tile_X3Y6_LUT4AB/E6END[1] Tile_X3Y6_LUT4AB/E6END[2] Tile_X3Y6_LUT4AB/E6END[3] Tile_X3Y6_LUT4AB/E6END[4]
+ Tile_X3Y6_LUT4AB/E6END[5] Tile_X3Y6_LUT4AB/E6END[6] Tile_X3Y6_LUT4AB/E6END[7] Tile_X3Y6_LUT4AB/E6END[8]
+ Tile_X3Y6_LUT4AB/E6END[9] Tile_X4Y6_LUT4AB/EE4END[0] Tile_X4Y6_LUT4AB/EE4END[10]
+ Tile_X4Y6_LUT4AB/EE4END[11] Tile_X4Y6_LUT4AB/EE4END[12] Tile_X4Y6_LUT4AB/EE4END[13]
+ Tile_X4Y6_LUT4AB/EE4END[14] Tile_X4Y6_LUT4AB/EE4END[15] Tile_X4Y6_LUT4AB/EE4END[1]
+ Tile_X4Y6_LUT4AB/EE4END[2] Tile_X4Y6_LUT4AB/EE4END[3] Tile_X4Y6_LUT4AB/EE4END[4]
+ Tile_X4Y6_LUT4AB/EE4END[5] Tile_X4Y6_LUT4AB/EE4END[6] Tile_X4Y6_LUT4AB/EE4END[7]
+ Tile_X4Y6_LUT4AB/EE4END[8] Tile_X4Y6_LUT4AB/EE4END[9] Tile_X3Y6_LUT4AB/EE4END[0]
+ Tile_X3Y6_LUT4AB/EE4END[10] Tile_X3Y6_LUT4AB/EE4END[11] Tile_X3Y6_LUT4AB/EE4END[12]
+ Tile_X3Y6_LUT4AB/EE4END[13] Tile_X3Y6_LUT4AB/EE4END[14] Tile_X3Y6_LUT4AB/EE4END[15]
+ Tile_X3Y6_LUT4AB/EE4END[1] Tile_X3Y6_LUT4AB/EE4END[2] Tile_X3Y6_LUT4AB/EE4END[3]
+ Tile_X3Y6_LUT4AB/EE4END[4] Tile_X3Y6_LUT4AB/EE4END[5] Tile_X3Y6_LUT4AB/EE4END[6]
+ Tile_X3Y6_LUT4AB/EE4END[7] Tile_X3Y6_LUT4AB/EE4END[8] Tile_X3Y6_LUT4AB/EE4END[9]
+ Tile_X3Y6_LUT4AB/FrameData[0] Tile_X3Y6_LUT4AB/FrameData[10] Tile_X3Y6_LUT4AB/FrameData[11]
+ Tile_X3Y6_LUT4AB/FrameData[12] Tile_X3Y6_LUT4AB/FrameData[13] Tile_X3Y6_LUT4AB/FrameData[14]
+ Tile_X3Y6_LUT4AB/FrameData[15] Tile_X3Y6_LUT4AB/FrameData[16] Tile_X3Y6_LUT4AB/FrameData[17]
+ Tile_X3Y6_LUT4AB/FrameData[18] Tile_X3Y6_LUT4AB/FrameData[19] Tile_X3Y6_LUT4AB/FrameData[1]
+ Tile_X3Y6_LUT4AB/FrameData[20] Tile_X3Y6_LUT4AB/FrameData[21] Tile_X3Y6_LUT4AB/FrameData[22]
+ Tile_X3Y6_LUT4AB/FrameData[23] Tile_X3Y6_LUT4AB/FrameData[24] Tile_X3Y6_LUT4AB/FrameData[25]
+ Tile_X3Y6_LUT4AB/FrameData[26] Tile_X3Y6_LUT4AB/FrameData[27] Tile_X3Y6_LUT4AB/FrameData[28]
+ Tile_X3Y6_LUT4AB/FrameData[29] Tile_X3Y6_LUT4AB/FrameData[2] Tile_X3Y6_LUT4AB/FrameData[30]
+ Tile_X3Y6_LUT4AB/FrameData[31] Tile_X3Y6_LUT4AB/FrameData[3] Tile_X3Y6_LUT4AB/FrameData[4]
+ Tile_X3Y6_LUT4AB/FrameData[5] Tile_X3Y6_LUT4AB/FrameData[6] Tile_X3Y6_LUT4AB/FrameData[7]
+ Tile_X3Y6_LUT4AB/FrameData[8] Tile_X3Y6_LUT4AB/FrameData[9] Tile_X4Y6_LUT4AB/FrameData[0]
+ Tile_X4Y6_LUT4AB/FrameData[10] Tile_X4Y6_LUT4AB/FrameData[11] Tile_X4Y6_LUT4AB/FrameData[12]
+ Tile_X4Y6_LUT4AB/FrameData[13] Tile_X4Y6_LUT4AB/FrameData[14] Tile_X4Y6_LUT4AB/FrameData[15]
+ Tile_X4Y6_LUT4AB/FrameData[16] Tile_X4Y6_LUT4AB/FrameData[17] Tile_X4Y6_LUT4AB/FrameData[18]
+ Tile_X4Y6_LUT4AB/FrameData[19] Tile_X4Y6_LUT4AB/FrameData[1] Tile_X4Y6_LUT4AB/FrameData[20]
+ Tile_X4Y6_LUT4AB/FrameData[21] Tile_X4Y6_LUT4AB/FrameData[22] Tile_X4Y6_LUT4AB/FrameData[23]
+ Tile_X4Y6_LUT4AB/FrameData[24] Tile_X4Y6_LUT4AB/FrameData[25] Tile_X4Y6_LUT4AB/FrameData[26]
+ Tile_X4Y6_LUT4AB/FrameData[27] Tile_X4Y6_LUT4AB/FrameData[28] Tile_X4Y6_LUT4AB/FrameData[29]
+ Tile_X4Y6_LUT4AB/FrameData[2] Tile_X4Y6_LUT4AB/FrameData[30] Tile_X4Y6_LUT4AB/FrameData[31]
+ Tile_X4Y6_LUT4AB/FrameData[3] Tile_X4Y6_LUT4AB/FrameData[4] Tile_X4Y6_LUT4AB/FrameData[5]
+ Tile_X4Y6_LUT4AB/FrameData[6] Tile_X4Y6_LUT4AB/FrameData[7] Tile_X4Y6_LUT4AB/FrameData[8]
+ Tile_X4Y6_LUT4AB/FrameData[9] Tile_X3Y6_LUT4AB/FrameStrobe[0] Tile_X3Y6_LUT4AB/FrameStrobe[10]
+ Tile_X3Y6_LUT4AB/FrameStrobe[11] Tile_X3Y6_LUT4AB/FrameStrobe[12] Tile_X3Y6_LUT4AB/FrameStrobe[13]
+ Tile_X3Y6_LUT4AB/FrameStrobe[14] Tile_X3Y6_LUT4AB/FrameStrobe[15] Tile_X3Y6_LUT4AB/FrameStrobe[16]
+ Tile_X3Y6_LUT4AB/FrameStrobe[17] Tile_X3Y6_LUT4AB/FrameStrobe[18] Tile_X3Y6_LUT4AB/FrameStrobe[19]
+ Tile_X3Y6_LUT4AB/FrameStrobe[1] Tile_X3Y6_LUT4AB/FrameStrobe[2] Tile_X3Y6_LUT4AB/FrameStrobe[3]
+ Tile_X3Y6_LUT4AB/FrameStrobe[4] Tile_X3Y6_LUT4AB/FrameStrobe[5] Tile_X3Y6_LUT4AB/FrameStrobe[6]
+ Tile_X3Y6_LUT4AB/FrameStrobe[7] Tile_X3Y6_LUT4AB/FrameStrobe[8] Tile_X3Y6_LUT4AB/FrameStrobe[9]
+ Tile_X3Y5_LUT4AB/FrameStrobe[0] Tile_X3Y5_LUT4AB/FrameStrobe[10] Tile_X3Y5_LUT4AB/FrameStrobe[11]
+ Tile_X3Y5_LUT4AB/FrameStrobe[12] Tile_X3Y5_LUT4AB/FrameStrobe[13] Tile_X3Y5_LUT4AB/FrameStrobe[14]
+ Tile_X3Y5_LUT4AB/FrameStrobe[15] Tile_X3Y5_LUT4AB/FrameStrobe[16] Tile_X3Y5_LUT4AB/FrameStrobe[17]
+ Tile_X3Y5_LUT4AB/FrameStrobe[18] Tile_X3Y5_LUT4AB/FrameStrobe[19] Tile_X3Y5_LUT4AB/FrameStrobe[1]
+ Tile_X3Y5_LUT4AB/FrameStrobe[2] Tile_X3Y5_LUT4AB/FrameStrobe[3] Tile_X3Y5_LUT4AB/FrameStrobe[4]
+ Tile_X3Y5_LUT4AB/FrameStrobe[5] Tile_X3Y5_LUT4AB/FrameStrobe[6] Tile_X3Y5_LUT4AB/FrameStrobe[7]
+ Tile_X3Y5_LUT4AB/FrameStrobe[8] Tile_X3Y5_LUT4AB/FrameStrobe[9] Tile_X3Y6_LUT4AB/N1BEG[0]
+ Tile_X3Y6_LUT4AB/N1BEG[1] Tile_X3Y6_LUT4AB/N1BEG[2] Tile_X3Y6_LUT4AB/N1BEG[3] Tile_X3Y7_LUT4AB/N1BEG[0]
+ Tile_X3Y7_LUT4AB/N1BEG[1] Tile_X3Y7_LUT4AB/N1BEG[2] Tile_X3Y7_LUT4AB/N1BEG[3] Tile_X3Y6_LUT4AB/N2BEG[0]
+ Tile_X3Y6_LUT4AB/N2BEG[1] Tile_X3Y6_LUT4AB/N2BEG[2] Tile_X3Y6_LUT4AB/N2BEG[3] Tile_X3Y6_LUT4AB/N2BEG[4]
+ Tile_X3Y6_LUT4AB/N2BEG[5] Tile_X3Y6_LUT4AB/N2BEG[6] Tile_X3Y6_LUT4AB/N2BEG[7] Tile_X3Y5_LUT4AB/N2END[0]
+ Tile_X3Y5_LUT4AB/N2END[1] Tile_X3Y5_LUT4AB/N2END[2] Tile_X3Y5_LUT4AB/N2END[3] Tile_X3Y5_LUT4AB/N2END[4]
+ Tile_X3Y5_LUT4AB/N2END[5] Tile_X3Y5_LUT4AB/N2END[6] Tile_X3Y5_LUT4AB/N2END[7] Tile_X3Y6_LUT4AB/N2END[0]
+ Tile_X3Y6_LUT4AB/N2END[1] Tile_X3Y6_LUT4AB/N2END[2] Tile_X3Y6_LUT4AB/N2END[3] Tile_X3Y6_LUT4AB/N2END[4]
+ Tile_X3Y6_LUT4AB/N2END[5] Tile_X3Y6_LUT4AB/N2END[6] Tile_X3Y6_LUT4AB/N2END[7] Tile_X3Y7_LUT4AB/N2BEG[0]
+ Tile_X3Y7_LUT4AB/N2BEG[1] Tile_X3Y7_LUT4AB/N2BEG[2] Tile_X3Y7_LUT4AB/N2BEG[3] Tile_X3Y7_LUT4AB/N2BEG[4]
+ Tile_X3Y7_LUT4AB/N2BEG[5] Tile_X3Y7_LUT4AB/N2BEG[6] Tile_X3Y7_LUT4AB/N2BEG[7] Tile_X3Y6_LUT4AB/N4BEG[0]
+ Tile_X3Y6_LUT4AB/N4BEG[10] Tile_X3Y6_LUT4AB/N4BEG[11] Tile_X3Y6_LUT4AB/N4BEG[12]
+ Tile_X3Y6_LUT4AB/N4BEG[13] Tile_X3Y6_LUT4AB/N4BEG[14] Tile_X3Y6_LUT4AB/N4BEG[15]
+ Tile_X3Y6_LUT4AB/N4BEG[1] Tile_X3Y6_LUT4AB/N4BEG[2] Tile_X3Y6_LUT4AB/N4BEG[3] Tile_X3Y6_LUT4AB/N4BEG[4]
+ Tile_X3Y6_LUT4AB/N4BEG[5] Tile_X3Y6_LUT4AB/N4BEG[6] Tile_X3Y6_LUT4AB/N4BEG[7] Tile_X3Y6_LUT4AB/N4BEG[8]
+ Tile_X3Y6_LUT4AB/N4BEG[9] Tile_X3Y7_LUT4AB/N4BEG[0] Tile_X3Y7_LUT4AB/N4BEG[10] Tile_X3Y7_LUT4AB/N4BEG[11]
+ Tile_X3Y7_LUT4AB/N4BEG[12] Tile_X3Y7_LUT4AB/N4BEG[13] Tile_X3Y7_LUT4AB/N4BEG[14]
+ Tile_X3Y7_LUT4AB/N4BEG[15] Tile_X3Y7_LUT4AB/N4BEG[1] Tile_X3Y7_LUT4AB/N4BEG[2] Tile_X3Y7_LUT4AB/N4BEG[3]
+ Tile_X3Y7_LUT4AB/N4BEG[4] Tile_X3Y7_LUT4AB/N4BEG[5] Tile_X3Y7_LUT4AB/N4BEG[6] Tile_X3Y7_LUT4AB/N4BEG[7]
+ Tile_X3Y7_LUT4AB/N4BEG[8] Tile_X3Y7_LUT4AB/N4BEG[9] Tile_X3Y6_LUT4AB/NN4BEG[0] Tile_X3Y6_LUT4AB/NN4BEG[10]
+ Tile_X3Y6_LUT4AB/NN4BEG[11] Tile_X3Y6_LUT4AB/NN4BEG[12] Tile_X3Y6_LUT4AB/NN4BEG[13]
+ Tile_X3Y6_LUT4AB/NN4BEG[14] Tile_X3Y6_LUT4AB/NN4BEG[15] Tile_X3Y6_LUT4AB/NN4BEG[1]
+ Tile_X3Y6_LUT4AB/NN4BEG[2] Tile_X3Y6_LUT4AB/NN4BEG[3] Tile_X3Y6_LUT4AB/NN4BEG[4]
+ Tile_X3Y6_LUT4AB/NN4BEG[5] Tile_X3Y6_LUT4AB/NN4BEG[6] Tile_X3Y6_LUT4AB/NN4BEG[7]
+ Tile_X3Y6_LUT4AB/NN4BEG[8] Tile_X3Y6_LUT4AB/NN4BEG[9] Tile_X3Y7_LUT4AB/NN4BEG[0]
+ Tile_X3Y7_LUT4AB/NN4BEG[10] Tile_X3Y7_LUT4AB/NN4BEG[11] Tile_X3Y7_LUT4AB/NN4BEG[12]
+ Tile_X3Y7_LUT4AB/NN4BEG[13] Tile_X3Y7_LUT4AB/NN4BEG[14] Tile_X3Y7_LUT4AB/NN4BEG[15]
+ Tile_X3Y7_LUT4AB/NN4BEG[1] Tile_X3Y7_LUT4AB/NN4BEG[2] Tile_X3Y7_LUT4AB/NN4BEG[3]
+ Tile_X3Y7_LUT4AB/NN4BEG[4] Tile_X3Y7_LUT4AB/NN4BEG[5] Tile_X3Y7_LUT4AB/NN4BEG[6]
+ Tile_X3Y7_LUT4AB/NN4BEG[7] Tile_X3Y7_LUT4AB/NN4BEG[8] Tile_X3Y7_LUT4AB/NN4BEG[9]
+ Tile_X3Y7_LUT4AB/S1END[0] Tile_X3Y7_LUT4AB/S1END[1] Tile_X3Y7_LUT4AB/S1END[2] Tile_X3Y7_LUT4AB/S1END[3]
+ Tile_X3Y6_LUT4AB/S1END[0] Tile_X3Y6_LUT4AB/S1END[1] Tile_X3Y6_LUT4AB/S1END[2] Tile_X3Y6_LUT4AB/S1END[3]
+ Tile_X3Y7_LUT4AB/S2MID[0] Tile_X3Y7_LUT4AB/S2MID[1] Tile_X3Y7_LUT4AB/S2MID[2] Tile_X3Y7_LUT4AB/S2MID[3]
+ Tile_X3Y7_LUT4AB/S2MID[4] Tile_X3Y7_LUT4AB/S2MID[5] Tile_X3Y7_LUT4AB/S2MID[6] Tile_X3Y7_LUT4AB/S2MID[7]
+ Tile_X3Y7_LUT4AB/S2END[0] Tile_X3Y7_LUT4AB/S2END[1] Tile_X3Y7_LUT4AB/S2END[2] Tile_X3Y7_LUT4AB/S2END[3]
+ Tile_X3Y7_LUT4AB/S2END[4] Tile_X3Y7_LUT4AB/S2END[5] Tile_X3Y7_LUT4AB/S2END[6] Tile_X3Y7_LUT4AB/S2END[7]
+ Tile_X3Y6_LUT4AB/S2END[0] Tile_X3Y6_LUT4AB/S2END[1] Tile_X3Y6_LUT4AB/S2END[2] Tile_X3Y6_LUT4AB/S2END[3]
+ Tile_X3Y6_LUT4AB/S2END[4] Tile_X3Y6_LUT4AB/S2END[5] Tile_X3Y6_LUT4AB/S2END[6] Tile_X3Y6_LUT4AB/S2END[7]
+ Tile_X3Y6_LUT4AB/S2MID[0] Tile_X3Y6_LUT4AB/S2MID[1] Tile_X3Y6_LUT4AB/S2MID[2] Tile_X3Y6_LUT4AB/S2MID[3]
+ Tile_X3Y6_LUT4AB/S2MID[4] Tile_X3Y6_LUT4AB/S2MID[5] Tile_X3Y6_LUT4AB/S2MID[6] Tile_X3Y6_LUT4AB/S2MID[7]
+ Tile_X3Y7_LUT4AB/S4END[0] Tile_X3Y7_LUT4AB/S4END[10] Tile_X3Y7_LUT4AB/S4END[11]
+ Tile_X3Y7_LUT4AB/S4END[12] Tile_X3Y7_LUT4AB/S4END[13] Tile_X3Y7_LUT4AB/S4END[14]
+ Tile_X3Y7_LUT4AB/S4END[15] Tile_X3Y7_LUT4AB/S4END[1] Tile_X3Y7_LUT4AB/S4END[2] Tile_X3Y7_LUT4AB/S4END[3]
+ Tile_X3Y7_LUT4AB/S4END[4] Tile_X3Y7_LUT4AB/S4END[5] Tile_X3Y7_LUT4AB/S4END[6] Tile_X3Y7_LUT4AB/S4END[7]
+ Tile_X3Y7_LUT4AB/S4END[8] Tile_X3Y7_LUT4AB/S4END[9] Tile_X3Y6_LUT4AB/S4END[0] Tile_X3Y6_LUT4AB/S4END[10]
+ Tile_X3Y6_LUT4AB/S4END[11] Tile_X3Y6_LUT4AB/S4END[12] Tile_X3Y6_LUT4AB/S4END[13]
+ Tile_X3Y6_LUT4AB/S4END[14] Tile_X3Y6_LUT4AB/S4END[15] Tile_X3Y6_LUT4AB/S4END[1]
+ Tile_X3Y6_LUT4AB/S4END[2] Tile_X3Y6_LUT4AB/S4END[3] Tile_X3Y6_LUT4AB/S4END[4] Tile_X3Y6_LUT4AB/S4END[5]
+ Tile_X3Y6_LUT4AB/S4END[6] Tile_X3Y6_LUT4AB/S4END[7] Tile_X3Y6_LUT4AB/S4END[8] Tile_X3Y6_LUT4AB/S4END[9]
+ Tile_X3Y7_LUT4AB/SS4END[0] Tile_X3Y7_LUT4AB/SS4END[10] Tile_X3Y7_LUT4AB/SS4END[11]
+ Tile_X3Y7_LUT4AB/SS4END[12] Tile_X3Y7_LUT4AB/SS4END[13] Tile_X3Y7_LUT4AB/SS4END[14]
+ Tile_X3Y7_LUT4AB/SS4END[15] Tile_X3Y7_LUT4AB/SS4END[1] Tile_X3Y7_LUT4AB/SS4END[2]
+ Tile_X3Y7_LUT4AB/SS4END[3] Tile_X3Y7_LUT4AB/SS4END[4] Tile_X3Y7_LUT4AB/SS4END[5]
+ Tile_X3Y7_LUT4AB/SS4END[6] Tile_X3Y7_LUT4AB/SS4END[7] Tile_X3Y7_LUT4AB/SS4END[8]
+ Tile_X3Y7_LUT4AB/SS4END[9] Tile_X3Y6_LUT4AB/SS4END[0] Tile_X3Y6_LUT4AB/SS4END[10]
+ Tile_X3Y6_LUT4AB/SS4END[11] Tile_X3Y6_LUT4AB/SS4END[12] Tile_X3Y6_LUT4AB/SS4END[13]
+ Tile_X3Y6_LUT4AB/SS4END[14] Tile_X3Y6_LUT4AB/SS4END[15] Tile_X3Y6_LUT4AB/SS4END[1]
+ Tile_X3Y6_LUT4AB/SS4END[2] Tile_X3Y6_LUT4AB/SS4END[3] Tile_X3Y6_LUT4AB/SS4END[4]
+ Tile_X3Y6_LUT4AB/SS4END[5] Tile_X3Y6_LUT4AB/SS4END[6] Tile_X3Y6_LUT4AB/SS4END[7]
+ Tile_X3Y6_LUT4AB/SS4END[8] Tile_X3Y6_LUT4AB/SS4END[9] Tile_X3Y6_LUT4AB/UserCLK Tile_X3Y5_LUT4AB/UserCLK
+ VGND VPWR Tile_X3Y6_LUT4AB/W1BEG[0] Tile_X3Y6_LUT4AB/W1BEG[1] Tile_X3Y6_LUT4AB/W1BEG[2]
+ Tile_X3Y6_LUT4AB/W1BEG[3] Tile_X4Y6_LUT4AB/W1BEG[0] Tile_X4Y6_LUT4AB/W1BEG[1] Tile_X4Y6_LUT4AB/W1BEG[2]
+ Tile_X4Y6_LUT4AB/W1BEG[3] Tile_X3Y6_LUT4AB/W2BEG[0] Tile_X3Y6_LUT4AB/W2BEG[1] Tile_X3Y6_LUT4AB/W2BEG[2]
+ Tile_X3Y6_LUT4AB/W2BEG[3] Tile_X3Y6_LUT4AB/W2BEG[4] Tile_X3Y6_LUT4AB/W2BEG[5] Tile_X3Y6_LUT4AB/W2BEG[6]
+ Tile_X3Y6_LUT4AB/W2BEG[7] Tile_X2Y6_LUT4AB/W2END[0] Tile_X2Y6_LUT4AB/W2END[1] Tile_X2Y6_LUT4AB/W2END[2]
+ Tile_X2Y6_LUT4AB/W2END[3] Tile_X2Y6_LUT4AB/W2END[4] Tile_X2Y6_LUT4AB/W2END[5] Tile_X2Y6_LUT4AB/W2END[6]
+ Tile_X2Y6_LUT4AB/W2END[7] Tile_X3Y6_LUT4AB/W2END[0] Tile_X3Y6_LUT4AB/W2END[1] Tile_X3Y6_LUT4AB/W2END[2]
+ Tile_X3Y6_LUT4AB/W2END[3] Tile_X3Y6_LUT4AB/W2END[4] Tile_X3Y6_LUT4AB/W2END[5] Tile_X3Y6_LUT4AB/W2END[6]
+ Tile_X3Y6_LUT4AB/W2END[7] Tile_X4Y6_LUT4AB/W2BEG[0] Tile_X4Y6_LUT4AB/W2BEG[1] Tile_X4Y6_LUT4AB/W2BEG[2]
+ Tile_X4Y6_LUT4AB/W2BEG[3] Tile_X4Y6_LUT4AB/W2BEG[4] Tile_X4Y6_LUT4AB/W2BEG[5] Tile_X4Y6_LUT4AB/W2BEG[6]
+ Tile_X4Y6_LUT4AB/W2BEG[7] Tile_X3Y6_LUT4AB/W6BEG[0] Tile_X3Y6_LUT4AB/W6BEG[10] Tile_X3Y6_LUT4AB/W6BEG[11]
+ Tile_X3Y6_LUT4AB/W6BEG[1] Tile_X3Y6_LUT4AB/W6BEG[2] Tile_X3Y6_LUT4AB/W6BEG[3] Tile_X3Y6_LUT4AB/W6BEG[4]
+ Tile_X3Y6_LUT4AB/W6BEG[5] Tile_X3Y6_LUT4AB/W6BEG[6] Tile_X3Y6_LUT4AB/W6BEG[7] Tile_X3Y6_LUT4AB/W6BEG[8]
+ Tile_X3Y6_LUT4AB/W6BEG[9] Tile_X4Y6_LUT4AB/W6BEG[0] Tile_X4Y6_LUT4AB/W6BEG[10] Tile_X4Y6_LUT4AB/W6BEG[11]
+ Tile_X4Y6_LUT4AB/W6BEG[1] Tile_X4Y6_LUT4AB/W6BEG[2] Tile_X4Y6_LUT4AB/W6BEG[3] Tile_X4Y6_LUT4AB/W6BEG[4]
+ Tile_X4Y6_LUT4AB/W6BEG[5] Tile_X4Y6_LUT4AB/W6BEG[6] Tile_X4Y6_LUT4AB/W6BEG[7] Tile_X4Y6_LUT4AB/W6BEG[8]
+ Tile_X4Y6_LUT4AB/W6BEG[9] Tile_X3Y6_LUT4AB/WW4BEG[0] Tile_X3Y6_LUT4AB/WW4BEG[10]
+ Tile_X3Y6_LUT4AB/WW4BEG[11] Tile_X3Y6_LUT4AB/WW4BEG[12] Tile_X3Y6_LUT4AB/WW4BEG[13]
+ Tile_X3Y6_LUT4AB/WW4BEG[14] Tile_X3Y6_LUT4AB/WW4BEG[15] Tile_X3Y6_LUT4AB/WW4BEG[1]
+ Tile_X3Y6_LUT4AB/WW4BEG[2] Tile_X3Y6_LUT4AB/WW4BEG[3] Tile_X3Y6_LUT4AB/WW4BEG[4]
+ Tile_X3Y6_LUT4AB/WW4BEG[5] Tile_X3Y6_LUT4AB/WW4BEG[6] Tile_X3Y6_LUT4AB/WW4BEG[7]
+ Tile_X3Y6_LUT4AB/WW4BEG[8] Tile_X3Y6_LUT4AB/WW4BEG[9] Tile_X4Y6_LUT4AB/WW4BEG[0]
+ Tile_X4Y6_LUT4AB/WW4BEG[10] Tile_X4Y6_LUT4AB/WW4BEG[11] Tile_X4Y6_LUT4AB/WW4BEG[12]
+ Tile_X4Y6_LUT4AB/WW4BEG[13] Tile_X4Y6_LUT4AB/WW4BEG[14] Tile_X4Y6_LUT4AB/WW4BEG[15]
+ Tile_X4Y6_LUT4AB/WW4BEG[1] Tile_X4Y6_LUT4AB/WW4BEG[2] Tile_X4Y6_LUT4AB/WW4BEG[3]
+ Tile_X4Y6_LUT4AB/WW4BEG[4] Tile_X4Y6_LUT4AB/WW4BEG[5] Tile_X4Y6_LUT4AB/WW4BEG[6]
+ Tile_X4Y6_LUT4AB/WW4BEG[7] Tile_X4Y6_LUT4AB/WW4BEG[8] Tile_X4Y6_LUT4AB/WW4BEG[9]
+ LUT4AB
XTile_X1Y3_LUT4AB Tile_X1Y4_LUT4AB/Co Tile_X1Y3_LUT4AB/Co Tile_X2Y3_LUT4AB/E1END[0]
+ Tile_X2Y3_LUT4AB/E1END[1] Tile_X2Y3_LUT4AB/E1END[2] Tile_X2Y3_LUT4AB/E1END[3] Tile_X1Y3_LUT4AB/E1END[0]
+ Tile_X1Y3_LUT4AB/E1END[1] Tile_X1Y3_LUT4AB/E1END[2] Tile_X1Y3_LUT4AB/E1END[3] Tile_X2Y3_LUT4AB/E2MID[0]
+ Tile_X2Y3_LUT4AB/E2MID[1] Tile_X2Y3_LUT4AB/E2MID[2] Tile_X2Y3_LUT4AB/E2MID[3] Tile_X2Y3_LUT4AB/E2MID[4]
+ Tile_X2Y3_LUT4AB/E2MID[5] Tile_X2Y3_LUT4AB/E2MID[6] Tile_X2Y3_LUT4AB/E2MID[7] Tile_X2Y3_LUT4AB/E2END[0]
+ Tile_X2Y3_LUT4AB/E2END[1] Tile_X2Y3_LUT4AB/E2END[2] Tile_X2Y3_LUT4AB/E2END[3] Tile_X2Y3_LUT4AB/E2END[4]
+ Tile_X2Y3_LUT4AB/E2END[5] Tile_X2Y3_LUT4AB/E2END[6] Tile_X2Y3_LUT4AB/E2END[7] Tile_X1Y3_LUT4AB/E2END[0]
+ Tile_X1Y3_LUT4AB/E2END[1] Tile_X1Y3_LUT4AB/E2END[2] Tile_X1Y3_LUT4AB/E2END[3] Tile_X1Y3_LUT4AB/E2END[4]
+ Tile_X1Y3_LUT4AB/E2END[5] Tile_X1Y3_LUT4AB/E2END[6] Tile_X1Y3_LUT4AB/E2END[7] Tile_X1Y3_LUT4AB/E2MID[0]
+ Tile_X1Y3_LUT4AB/E2MID[1] Tile_X1Y3_LUT4AB/E2MID[2] Tile_X1Y3_LUT4AB/E2MID[3] Tile_X1Y3_LUT4AB/E2MID[4]
+ Tile_X1Y3_LUT4AB/E2MID[5] Tile_X1Y3_LUT4AB/E2MID[6] Tile_X1Y3_LUT4AB/E2MID[7] Tile_X2Y3_LUT4AB/E6END[0]
+ Tile_X2Y3_LUT4AB/E6END[10] Tile_X2Y3_LUT4AB/E6END[11] Tile_X2Y3_LUT4AB/E6END[1]
+ Tile_X2Y3_LUT4AB/E6END[2] Tile_X2Y3_LUT4AB/E6END[3] Tile_X2Y3_LUT4AB/E6END[4] Tile_X2Y3_LUT4AB/E6END[5]
+ Tile_X2Y3_LUT4AB/E6END[6] Tile_X2Y3_LUT4AB/E6END[7] Tile_X2Y3_LUT4AB/E6END[8] Tile_X2Y3_LUT4AB/E6END[9]
+ Tile_X1Y3_LUT4AB/E6END[0] Tile_X1Y3_LUT4AB/E6END[10] Tile_X1Y3_LUT4AB/E6END[11]
+ Tile_X1Y3_LUT4AB/E6END[1] Tile_X1Y3_LUT4AB/E6END[2] Tile_X1Y3_LUT4AB/E6END[3] Tile_X1Y3_LUT4AB/E6END[4]
+ Tile_X1Y3_LUT4AB/E6END[5] Tile_X1Y3_LUT4AB/E6END[6] Tile_X1Y3_LUT4AB/E6END[7] Tile_X1Y3_LUT4AB/E6END[8]
+ Tile_X1Y3_LUT4AB/E6END[9] Tile_X2Y3_LUT4AB/EE4END[0] Tile_X2Y3_LUT4AB/EE4END[10]
+ Tile_X2Y3_LUT4AB/EE4END[11] Tile_X2Y3_LUT4AB/EE4END[12] Tile_X2Y3_LUT4AB/EE4END[13]
+ Tile_X2Y3_LUT4AB/EE4END[14] Tile_X2Y3_LUT4AB/EE4END[15] Tile_X2Y3_LUT4AB/EE4END[1]
+ Tile_X2Y3_LUT4AB/EE4END[2] Tile_X2Y3_LUT4AB/EE4END[3] Tile_X2Y3_LUT4AB/EE4END[4]
+ Tile_X2Y3_LUT4AB/EE4END[5] Tile_X2Y3_LUT4AB/EE4END[6] Tile_X2Y3_LUT4AB/EE4END[7]
+ Tile_X2Y3_LUT4AB/EE4END[8] Tile_X2Y3_LUT4AB/EE4END[9] Tile_X1Y3_LUT4AB/EE4END[0]
+ Tile_X1Y3_LUT4AB/EE4END[10] Tile_X1Y3_LUT4AB/EE4END[11] Tile_X1Y3_LUT4AB/EE4END[12]
+ Tile_X1Y3_LUT4AB/EE4END[13] Tile_X1Y3_LUT4AB/EE4END[14] Tile_X1Y3_LUT4AB/EE4END[15]
+ Tile_X1Y3_LUT4AB/EE4END[1] Tile_X1Y3_LUT4AB/EE4END[2] Tile_X1Y3_LUT4AB/EE4END[3]
+ Tile_X1Y3_LUT4AB/EE4END[4] Tile_X1Y3_LUT4AB/EE4END[5] Tile_X1Y3_LUT4AB/EE4END[6]
+ Tile_X1Y3_LUT4AB/EE4END[7] Tile_X1Y3_LUT4AB/EE4END[8] Tile_X1Y3_LUT4AB/EE4END[9]
+ Tile_X1Y3_LUT4AB/FrameData[0] Tile_X1Y3_LUT4AB/FrameData[10] Tile_X1Y3_LUT4AB/FrameData[11]
+ Tile_X1Y3_LUT4AB/FrameData[12] Tile_X1Y3_LUT4AB/FrameData[13] Tile_X1Y3_LUT4AB/FrameData[14]
+ Tile_X1Y3_LUT4AB/FrameData[15] Tile_X1Y3_LUT4AB/FrameData[16] Tile_X1Y3_LUT4AB/FrameData[17]
+ Tile_X1Y3_LUT4AB/FrameData[18] Tile_X1Y3_LUT4AB/FrameData[19] Tile_X1Y3_LUT4AB/FrameData[1]
+ Tile_X1Y3_LUT4AB/FrameData[20] Tile_X1Y3_LUT4AB/FrameData[21] Tile_X1Y3_LUT4AB/FrameData[22]
+ Tile_X1Y3_LUT4AB/FrameData[23] Tile_X1Y3_LUT4AB/FrameData[24] Tile_X1Y3_LUT4AB/FrameData[25]
+ Tile_X1Y3_LUT4AB/FrameData[26] Tile_X1Y3_LUT4AB/FrameData[27] Tile_X1Y3_LUT4AB/FrameData[28]
+ Tile_X1Y3_LUT4AB/FrameData[29] Tile_X1Y3_LUT4AB/FrameData[2] Tile_X1Y3_LUT4AB/FrameData[30]
+ Tile_X1Y3_LUT4AB/FrameData[31] Tile_X1Y3_LUT4AB/FrameData[3] Tile_X1Y3_LUT4AB/FrameData[4]
+ Tile_X1Y3_LUT4AB/FrameData[5] Tile_X1Y3_LUT4AB/FrameData[6] Tile_X1Y3_LUT4AB/FrameData[7]
+ Tile_X1Y3_LUT4AB/FrameData[8] Tile_X1Y3_LUT4AB/FrameData[9] Tile_X2Y3_LUT4AB/FrameData[0]
+ Tile_X2Y3_LUT4AB/FrameData[10] Tile_X2Y3_LUT4AB/FrameData[11] Tile_X2Y3_LUT4AB/FrameData[12]
+ Tile_X2Y3_LUT4AB/FrameData[13] Tile_X2Y3_LUT4AB/FrameData[14] Tile_X2Y3_LUT4AB/FrameData[15]
+ Tile_X2Y3_LUT4AB/FrameData[16] Tile_X2Y3_LUT4AB/FrameData[17] Tile_X2Y3_LUT4AB/FrameData[18]
+ Tile_X2Y3_LUT4AB/FrameData[19] Tile_X2Y3_LUT4AB/FrameData[1] Tile_X2Y3_LUT4AB/FrameData[20]
+ Tile_X2Y3_LUT4AB/FrameData[21] Tile_X2Y3_LUT4AB/FrameData[22] Tile_X2Y3_LUT4AB/FrameData[23]
+ Tile_X2Y3_LUT4AB/FrameData[24] Tile_X2Y3_LUT4AB/FrameData[25] Tile_X2Y3_LUT4AB/FrameData[26]
+ Tile_X2Y3_LUT4AB/FrameData[27] Tile_X2Y3_LUT4AB/FrameData[28] Tile_X2Y3_LUT4AB/FrameData[29]
+ Tile_X2Y3_LUT4AB/FrameData[2] Tile_X2Y3_LUT4AB/FrameData[30] Tile_X2Y3_LUT4AB/FrameData[31]
+ Tile_X2Y3_LUT4AB/FrameData[3] Tile_X2Y3_LUT4AB/FrameData[4] Tile_X2Y3_LUT4AB/FrameData[5]
+ Tile_X2Y3_LUT4AB/FrameData[6] Tile_X2Y3_LUT4AB/FrameData[7] Tile_X2Y3_LUT4AB/FrameData[8]
+ Tile_X2Y3_LUT4AB/FrameData[9] Tile_X1Y3_LUT4AB/FrameStrobe[0] Tile_X1Y3_LUT4AB/FrameStrobe[10]
+ Tile_X1Y3_LUT4AB/FrameStrobe[11] Tile_X1Y3_LUT4AB/FrameStrobe[12] Tile_X1Y3_LUT4AB/FrameStrobe[13]
+ Tile_X1Y3_LUT4AB/FrameStrobe[14] Tile_X1Y3_LUT4AB/FrameStrobe[15] Tile_X1Y3_LUT4AB/FrameStrobe[16]
+ Tile_X1Y3_LUT4AB/FrameStrobe[17] Tile_X1Y3_LUT4AB/FrameStrobe[18] Tile_X1Y3_LUT4AB/FrameStrobe[19]
+ Tile_X1Y3_LUT4AB/FrameStrobe[1] Tile_X1Y3_LUT4AB/FrameStrobe[2] Tile_X1Y3_LUT4AB/FrameStrobe[3]
+ Tile_X1Y3_LUT4AB/FrameStrobe[4] Tile_X1Y3_LUT4AB/FrameStrobe[5] Tile_X1Y3_LUT4AB/FrameStrobe[6]
+ Tile_X1Y3_LUT4AB/FrameStrobe[7] Tile_X1Y3_LUT4AB/FrameStrobe[8] Tile_X1Y3_LUT4AB/FrameStrobe[9]
+ Tile_X1Y2_LUT4AB/FrameStrobe[0] Tile_X1Y2_LUT4AB/FrameStrobe[10] Tile_X1Y2_LUT4AB/FrameStrobe[11]
+ Tile_X1Y2_LUT4AB/FrameStrobe[12] Tile_X1Y2_LUT4AB/FrameStrobe[13] Tile_X1Y2_LUT4AB/FrameStrobe[14]
+ Tile_X1Y2_LUT4AB/FrameStrobe[15] Tile_X1Y2_LUT4AB/FrameStrobe[16] Tile_X1Y2_LUT4AB/FrameStrobe[17]
+ Tile_X1Y2_LUT4AB/FrameStrobe[18] Tile_X1Y2_LUT4AB/FrameStrobe[19] Tile_X1Y2_LUT4AB/FrameStrobe[1]
+ Tile_X1Y2_LUT4AB/FrameStrobe[2] Tile_X1Y2_LUT4AB/FrameStrobe[3] Tile_X1Y2_LUT4AB/FrameStrobe[4]
+ Tile_X1Y2_LUT4AB/FrameStrobe[5] Tile_X1Y2_LUT4AB/FrameStrobe[6] Tile_X1Y2_LUT4AB/FrameStrobe[7]
+ Tile_X1Y2_LUT4AB/FrameStrobe[8] Tile_X1Y2_LUT4AB/FrameStrobe[9] Tile_X1Y3_LUT4AB/N1BEG[0]
+ Tile_X1Y3_LUT4AB/N1BEG[1] Tile_X1Y3_LUT4AB/N1BEG[2] Tile_X1Y3_LUT4AB/N1BEG[3] Tile_X1Y4_LUT4AB/N1BEG[0]
+ Tile_X1Y4_LUT4AB/N1BEG[1] Tile_X1Y4_LUT4AB/N1BEG[2] Tile_X1Y4_LUT4AB/N1BEG[3] Tile_X1Y3_LUT4AB/N2BEG[0]
+ Tile_X1Y3_LUT4AB/N2BEG[1] Tile_X1Y3_LUT4AB/N2BEG[2] Tile_X1Y3_LUT4AB/N2BEG[3] Tile_X1Y3_LUT4AB/N2BEG[4]
+ Tile_X1Y3_LUT4AB/N2BEG[5] Tile_X1Y3_LUT4AB/N2BEG[6] Tile_X1Y3_LUT4AB/N2BEG[7] Tile_X1Y2_LUT4AB/N2END[0]
+ Tile_X1Y2_LUT4AB/N2END[1] Tile_X1Y2_LUT4AB/N2END[2] Tile_X1Y2_LUT4AB/N2END[3] Tile_X1Y2_LUT4AB/N2END[4]
+ Tile_X1Y2_LUT4AB/N2END[5] Tile_X1Y2_LUT4AB/N2END[6] Tile_X1Y2_LUT4AB/N2END[7] Tile_X1Y3_LUT4AB/N2END[0]
+ Tile_X1Y3_LUT4AB/N2END[1] Tile_X1Y3_LUT4AB/N2END[2] Tile_X1Y3_LUT4AB/N2END[3] Tile_X1Y3_LUT4AB/N2END[4]
+ Tile_X1Y3_LUT4AB/N2END[5] Tile_X1Y3_LUT4AB/N2END[6] Tile_X1Y3_LUT4AB/N2END[7] Tile_X1Y4_LUT4AB/N2BEG[0]
+ Tile_X1Y4_LUT4AB/N2BEG[1] Tile_X1Y4_LUT4AB/N2BEG[2] Tile_X1Y4_LUT4AB/N2BEG[3] Tile_X1Y4_LUT4AB/N2BEG[4]
+ Tile_X1Y4_LUT4AB/N2BEG[5] Tile_X1Y4_LUT4AB/N2BEG[6] Tile_X1Y4_LUT4AB/N2BEG[7] Tile_X1Y3_LUT4AB/N4BEG[0]
+ Tile_X1Y3_LUT4AB/N4BEG[10] Tile_X1Y3_LUT4AB/N4BEG[11] Tile_X1Y3_LUT4AB/N4BEG[12]
+ Tile_X1Y3_LUT4AB/N4BEG[13] Tile_X1Y3_LUT4AB/N4BEG[14] Tile_X1Y3_LUT4AB/N4BEG[15]
+ Tile_X1Y3_LUT4AB/N4BEG[1] Tile_X1Y3_LUT4AB/N4BEG[2] Tile_X1Y3_LUT4AB/N4BEG[3] Tile_X1Y3_LUT4AB/N4BEG[4]
+ Tile_X1Y3_LUT4AB/N4BEG[5] Tile_X1Y3_LUT4AB/N4BEG[6] Tile_X1Y3_LUT4AB/N4BEG[7] Tile_X1Y3_LUT4AB/N4BEG[8]
+ Tile_X1Y3_LUT4AB/N4BEG[9] Tile_X1Y4_LUT4AB/N4BEG[0] Tile_X1Y4_LUT4AB/N4BEG[10] Tile_X1Y4_LUT4AB/N4BEG[11]
+ Tile_X1Y4_LUT4AB/N4BEG[12] Tile_X1Y4_LUT4AB/N4BEG[13] Tile_X1Y4_LUT4AB/N4BEG[14]
+ Tile_X1Y4_LUT4AB/N4BEG[15] Tile_X1Y4_LUT4AB/N4BEG[1] Tile_X1Y4_LUT4AB/N4BEG[2] Tile_X1Y4_LUT4AB/N4BEG[3]
+ Tile_X1Y4_LUT4AB/N4BEG[4] Tile_X1Y4_LUT4AB/N4BEG[5] Tile_X1Y4_LUT4AB/N4BEG[6] Tile_X1Y4_LUT4AB/N4BEG[7]
+ Tile_X1Y4_LUT4AB/N4BEG[8] Tile_X1Y4_LUT4AB/N4BEG[9] Tile_X1Y3_LUT4AB/NN4BEG[0] Tile_X1Y3_LUT4AB/NN4BEG[10]
+ Tile_X1Y3_LUT4AB/NN4BEG[11] Tile_X1Y3_LUT4AB/NN4BEG[12] Tile_X1Y3_LUT4AB/NN4BEG[13]
+ Tile_X1Y3_LUT4AB/NN4BEG[14] Tile_X1Y3_LUT4AB/NN4BEG[15] Tile_X1Y3_LUT4AB/NN4BEG[1]
+ Tile_X1Y3_LUT4AB/NN4BEG[2] Tile_X1Y3_LUT4AB/NN4BEG[3] Tile_X1Y3_LUT4AB/NN4BEG[4]
+ Tile_X1Y3_LUT4AB/NN4BEG[5] Tile_X1Y3_LUT4AB/NN4BEG[6] Tile_X1Y3_LUT4AB/NN4BEG[7]
+ Tile_X1Y3_LUT4AB/NN4BEG[8] Tile_X1Y3_LUT4AB/NN4BEG[9] Tile_X1Y4_LUT4AB/NN4BEG[0]
+ Tile_X1Y4_LUT4AB/NN4BEG[10] Tile_X1Y4_LUT4AB/NN4BEG[11] Tile_X1Y4_LUT4AB/NN4BEG[12]
+ Tile_X1Y4_LUT4AB/NN4BEG[13] Tile_X1Y4_LUT4AB/NN4BEG[14] Tile_X1Y4_LUT4AB/NN4BEG[15]
+ Tile_X1Y4_LUT4AB/NN4BEG[1] Tile_X1Y4_LUT4AB/NN4BEG[2] Tile_X1Y4_LUT4AB/NN4BEG[3]
+ Tile_X1Y4_LUT4AB/NN4BEG[4] Tile_X1Y4_LUT4AB/NN4BEG[5] Tile_X1Y4_LUT4AB/NN4BEG[6]
+ Tile_X1Y4_LUT4AB/NN4BEG[7] Tile_X1Y4_LUT4AB/NN4BEG[8] Tile_X1Y4_LUT4AB/NN4BEG[9]
+ Tile_X1Y4_LUT4AB/S1END[0] Tile_X1Y4_LUT4AB/S1END[1] Tile_X1Y4_LUT4AB/S1END[2] Tile_X1Y4_LUT4AB/S1END[3]
+ Tile_X1Y3_LUT4AB/S1END[0] Tile_X1Y3_LUT4AB/S1END[1] Tile_X1Y3_LUT4AB/S1END[2] Tile_X1Y3_LUT4AB/S1END[3]
+ Tile_X1Y4_LUT4AB/S2MID[0] Tile_X1Y4_LUT4AB/S2MID[1] Tile_X1Y4_LUT4AB/S2MID[2] Tile_X1Y4_LUT4AB/S2MID[3]
+ Tile_X1Y4_LUT4AB/S2MID[4] Tile_X1Y4_LUT4AB/S2MID[5] Tile_X1Y4_LUT4AB/S2MID[6] Tile_X1Y4_LUT4AB/S2MID[7]
+ Tile_X1Y4_LUT4AB/S2END[0] Tile_X1Y4_LUT4AB/S2END[1] Tile_X1Y4_LUT4AB/S2END[2] Tile_X1Y4_LUT4AB/S2END[3]
+ Tile_X1Y4_LUT4AB/S2END[4] Tile_X1Y4_LUT4AB/S2END[5] Tile_X1Y4_LUT4AB/S2END[6] Tile_X1Y4_LUT4AB/S2END[7]
+ Tile_X1Y3_LUT4AB/S2END[0] Tile_X1Y3_LUT4AB/S2END[1] Tile_X1Y3_LUT4AB/S2END[2] Tile_X1Y3_LUT4AB/S2END[3]
+ Tile_X1Y3_LUT4AB/S2END[4] Tile_X1Y3_LUT4AB/S2END[5] Tile_X1Y3_LUT4AB/S2END[6] Tile_X1Y3_LUT4AB/S2END[7]
+ Tile_X1Y3_LUT4AB/S2MID[0] Tile_X1Y3_LUT4AB/S2MID[1] Tile_X1Y3_LUT4AB/S2MID[2] Tile_X1Y3_LUT4AB/S2MID[3]
+ Tile_X1Y3_LUT4AB/S2MID[4] Tile_X1Y3_LUT4AB/S2MID[5] Tile_X1Y3_LUT4AB/S2MID[6] Tile_X1Y3_LUT4AB/S2MID[7]
+ Tile_X1Y4_LUT4AB/S4END[0] Tile_X1Y4_LUT4AB/S4END[10] Tile_X1Y4_LUT4AB/S4END[11]
+ Tile_X1Y4_LUT4AB/S4END[12] Tile_X1Y4_LUT4AB/S4END[13] Tile_X1Y4_LUT4AB/S4END[14]
+ Tile_X1Y4_LUT4AB/S4END[15] Tile_X1Y4_LUT4AB/S4END[1] Tile_X1Y4_LUT4AB/S4END[2] Tile_X1Y4_LUT4AB/S4END[3]
+ Tile_X1Y4_LUT4AB/S4END[4] Tile_X1Y4_LUT4AB/S4END[5] Tile_X1Y4_LUT4AB/S4END[6] Tile_X1Y4_LUT4AB/S4END[7]
+ Tile_X1Y4_LUT4AB/S4END[8] Tile_X1Y4_LUT4AB/S4END[9] Tile_X1Y3_LUT4AB/S4END[0] Tile_X1Y3_LUT4AB/S4END[10]
+ Tile_X1Y3_LUT4AB/S4END[11] Tile_X1Y3_LUT4AB/S4END[12] Tile_X1Y3_LUT4AB/S4END[13]
+ Tile_X1Y3_LUT4AB/S4END[14] Tile_X1Y3_LUT4AB/S4END[15] Tile_X1Y3_LUT4AB/S4END[1]
+ Tile_X1Y3_LUT4AB/S4END[2] Tile_X1Y3_LUT4AB/S4END[3] Tile_X1Y3_LUT4AB/S4END[4] Tile_X1Y3_LUT4AB/S4END[5]
+ Tile_X1Y3_LUT4AB/S4END[6] Tile_X1Y3_LUT4AB/S4END[7] Tile_X1Y3_LUT4AB/S4END[8] Tile_X1Y3_LUT4AB/S4END[9]
+ Tile_X1Y4_LUT4AB/SS4END[0] Tile_X1Y4_LUT4AB/SS4END[10] Tile_X1Y4_LUT4AB/SS4END[11]
+ Tile_X1Y4_LUT4AB/SS4END[12] Tile_X1Y4_LUT4AB/SS4END[13] Tile_X1Y4_LUT4AB/SS4END[14]
+ Tile_X1Y4_LUT4AB/SS4END[15] Tile_X1Y4_LUT4AB/SS4END[1] Tile_X1Y4_LUT4AB/SS4END[2]
+ Tile_X1Y4_LUT4AB/SS4END[3] Tile_X1Y4_LUT4AB/SS4END[4] Tile_X1Y4_LUT4AB/SS4END[5]
+ Tile_X1Y4_LUT4AB/SS4END[6] Tile_X1Y4_LUT4AB/SS4END[7] Tile_X1Y4_LUT4AB/SS4END[8]
+ Tile_X1Y4_LUT4AB/SS4END[9] Tile_X1Y3_LUT4AB/SS4END[0] Tile_X1Y3_LUT4AB/SS4END[10]
+ Tile_X1Y3_LUT4AB/SS4END[11] Tile_X1Y3_LUT4AB/SS4END[12] Tile_X1Y3_LUT4AB/SS4END[13]
+ Tile_X1Y3_LUT4AB/SS4END[14] Tile_X1Y3_LUT4AB/SS4END[15] Tile_X1Y3_LUT4AB/SS4END[1]
+ Tile_X1Y3_LUT4AB/SS4END[2] Tile_X1Y3_LUT4AB/SS4END[3] Tile_X1Y3_LUT4AB/SS4END[4]
+ Tile_X1Y3_LUT4AB/SS4END[5] Tile_X1Y3_LUT4AB/SS4END[6] Tile_X1Y3_LUT4AB/SS4END[7]
+ Tile_X1Y3_LUT4AB/SS4END[8] Tile_X1Y3_LUT4AB/SS4END[9] Tile_X1Y3_LUT4AB/UserCLK Tile_X1Y2_LUT4AB/UserCLK
+ VGND VPWR Tile_X1Y3_LUT4AB/W1BEG[0] Tile_X1Y3_LUT4AB/W1BEG[1] Tile_X1Y3_LUT4AB/W1BEG[2]
+ Tile_X1Y3_LUT4AB/W1BEG[3] Tile_X2Y3_LUT4AB/W1BEG[0] Tile_X2Y3_LUT4AB/W1BEG[1] Tile_X2Y3_LUT4AB/W1BEG[2]
+ Tile_X2Y3_LUT4AB/W1BEG[3] Tile_X1Y3_LUT4AB/W2BEG[0] Tile_X1Y3_LUT4AB/W2BEG[1] Tile_X1Y3_LUT4AB/W2BEG[2]
+ Tile_X1Y3_LUT4AB/W2BEG[3] Tile_X1Y3_LUT4AB/W2BEG[4] Tile_X1Y3_LUT4AB/W2BEG[5] Tile_X1Y3_LUT4AB/W2BEG[6]
+ Tile_X1Y3_LUT4AB/W2BEG[7] Tile_X1Y3_LUT4AB/W2BEGb[0] Tile_X1Y3_LUT4AB/W2BEGb[1]
+ Tile_X1Y3_LUT4AB/W2BEGb[2] Tile_X1Y3_LUT4AB/W2BEGb[3] Tile_X1Y3_LUT4AB/W2BEGb[4]
+ Tile_X1Y3_LUT4AB/W2BEGb[5] Tile_X1Y3_LUT4AB/W2BEGb[6] Tile_X1Y3_LUT4AB/W2BEGb[7]
+ Tile_X1Y3_LUT4AB/W2END[0] Tile_X1Y3_LUT4AB/W2END[1] Tile_X1Y3_LUT4AB/W2END[2] Tile_X1Y3_LUT4AB/W2END[3]
+ Tile_X1Y3_LUT4AB/W2END[4] Tile_X1Y3_LUT4AB/W2END[5] Tile_X1Y3_LUT4AB/W2END[6] Tile_X1Y3_LUT4AB/W2END[7]
+ Tile_X2Y3_LUT4AB/W2BEG[0] Tile_X2Y3_LUT4AB/W2BEG[1] Tile_X2Y3_LUT4AB/W2BEG[2] Tile_X2Y3_LUT4AB/W2BEG[3]
+ Tile_X2Y3_LUT4AB/W2BEG[4] Tile_X2Y3_LUT4AB/W2BEG[5] Tile_X2Y3_LUT4AB/W2BEG[6] Tile_X2Y3_LUT4AB/W2BEG[7]
+ Tile_X1Y3_LUT4AB/W6BEG[0] Tile_X1Y3_LUT4AB/W6BEG[10] Tile_X1Y3_LUT4AB/W6BEG[11]
+ Tile_X1Y3_LUT4AB/W6BEG[1] Tile_X1Y3_LUT4AB/W6BEG[2] Tile_X1Y3_LUT4AB/W6BEG[3] Tile_X1Y3_LUT4AB/W6BEG[4]
+ Tile_X1Y3_LUT4AB/W6BEG[5] Tile_X1Y3_LUT4AB/W6BEG[6] Tile_X1Y3_LUT4AB/W6BEG[7] Tile_X1Y3_LUT4AB/W6BEG[8]
+ Tile_X1Y3_LUT4AB/W6BEG[9] Tile_X2Y3_LUT4AB/W6BEG[0] Tile_X2Y3_LUT4AB/W6BEG[10] Tile_X2Y3_LUT4AB/W6BEG[11]
+ Tile_X2Y3_LUT4AB/W6BEG[1] Tile_X2Y3_LUT4AB/W6BEG[2] Tile_X2Y3_LUT4AB/W6BEG[3] Tile_X2Y3_LUT4AB/W6BEG[4]
+ Tile_X2Y3_LUT4AB/W6BEG[5] Tile_X2Y3_LUT4AB/W6BEG[6] Tile_X2Y3_LUT4AB/W6BEG[7] Tile_X2Y3_LUT4AB/W6BEG[8]
+ Tile_X2Y3_LUT4AB/W6BEG[9] Tile_X1Y3_LUT4AB/WW4BEG[0] Tile_X1Y3_LUT4AB/WW4BEG[10]
+ Tile_X1Y3_LUT4AB/WW4BEG[11] Tile_X1Y3_LUT4AB/WW4BEG[12] Tile_X1Y3_LUT4AB/WW4BEG[13]
+ Tile_X1Y3_LUT4AB/WW4BEG[14] Tile_X1Y3_LUT4AB/WW4BEG[15] Tile_X1Y3_LUT4AB/WW4BEG[1]
+ Tile_X1Y3_LUT4AB/WW4BEG[2] Tile_X1Y3_LUT4AB/WW4BEG[3] Tile_X1Y3_LUT4AB/WW4BEG[4]
+ Tile_X1Y3_LUT4AB/WW4BEG[5] Tile_X1Y3_LUT4AB/WW4BEG[6] Tile_X1Y3_LUT4AB/WW4BEG[7]
+ Tile_X1Y3_LUT4AB/WW4BEG[8] Tile_X1Y3_LUT4AB/WW4BEG[9] Tile_X2Y3_LUT4AB/WW4BEG[0]
+ Tile_X2Y3_LUT4AB/WW4BEG[10] Tile_X2Y3_LUT4AB/WW4BEG[11] Tile_X2Y3_LUT4AB/WW4BEG[12]
+ Tile_X2Y3_LUT4AB/WW4BEG[13] Tile_X2Y3_LUT4AB/WW4BEG[14] Tile_X2Y3_LUT4AB/WW4BEG[15]
+ Tile_X2Y3_LUT4AB/WW4BEG[1] Tile_X2Y3_LUT4AB/WW4BEG[2] Tile_X2Y3_LUT4AB/WW4BEG[3]
+ Tile_X2Y3_LUT4AB/WW4BEG[4] Tile_X2Y3_LUT4AB/WW4BEG[5] Tile_X2Y3_LUT4AB/WW4BEG[6]
+ Tile_X2Y3_LUT4AB/WW4BEG[7] Tile_X2Y3_LUT4AB/WW4BEG[8] Tile_X2Y3_LUT4AB/WW4BEG[9]
+ LUT4AB
XTile_X4Y8_LUT4AB Tile_X4Y9_S_IO4/Co Tile_X4Y8_LUT4AB/Co Tile_X4Y8_LUT4AB/E1BEG[0]
+ Tile_X4Y8_LUT4AB/E1BEG[1] Tile_X4Y8_LUT4AB/E1BEG[2] Tile_X4Y8_LUT4AB/E1BEG[3] Tile_X4Y8_LUT4AB/E1END[0]
+ Tile_X4Y8_LUT4AB/E1END[1] Tile_X4Y8_LUT4AB/E1END[2] Tile_X4Y8_LUT4AB/E1END[3] Tile_X4Y8_LUT4AB/E2BEG[0]
+ Tile_X4Y8_LUT4AB/E2BEG[1] Tile_X4Y8_LUT4AB/E2BEG[2] Tile_X4Y8_LUT4AB/E2BEG[3] Tile_X4Y8_LUT4AB/E2BEG[4]
+ Tile_X4Y8_LUT4AB/E2BEG[5] Tile_X4Y8_LUT4AB/E2BEG[6] Tile_X4Y8_LUT4AB/E2BEG[7] Tile_X5Y8_E_TT_IF/E2END[0]
+ Tile_X5Y8_E_TT_IF/E2END[1] Tile_X5Y8_E_TT_IF/E2END[2] Tile_X5Y8_E_TT_IF/E2END[3]
+ Tile_X5Y8_E_TT_IF/E2END[4] Tile_X5Y8_E_TT_IF/E2END[5] Tile_X5Y8_E_TT_IF/E2END[6]
+ Tile_X5Y8_E_TT_IF/E2END[7] Tile_X4Y8_LUT4AB/E2END[0] Tile_X4Y8_LUT4AB/E2END[1] Tile_X4Y8_LUT4AB/E2END[2]
+ Tile_X4Y8_LUT4AB/E2END[3] Tile_X4Y8_LUT4AB/E2END[4] Tile_X4Y8_LUT4AB/E2END[5] Tile_X4Y8_LUT4AB/E2END[6]
+ Tile_X4Y8_LUT4AB/E2END[7] Tile_X4Y8_LUT4AB/E2MID[0] Tile_X4Y8_LUT4AB/E2MID[1] Tile_X4Y8_LUT4AB/E2MID[2]
+ Tile_X4Y8_LUT4AB/E2MID[3] Tile_X4Y8_LUT4AB/E2MID[4] Tile_X4Y8_LUT4AB/E2MID[5] Tile_X4Y8_LUT4AB/E2MID[6]
+ Tile_X4Y8_LUT4AB/E2MID[7] Tile_X4Y8_LUT4AB/E6BEG[0] Tile_X4Y8_LUT4AB/E6BEG[10] Tile_X4Y8_LUT4AB/E6BEG[11]
+ Tile_X4Y8_LUT4AB/E6BEG[1] Tile_X4Y8_LUT4AB/E6BEG[2] Tile_X4Y8_LUT4AB/E6BEG[3] Tile_X4Y8_LUT4AB/E6BEG[4]
+ Tile_X4Y8_LUT4AB/E6BEG[5] Tile_X4Y8_LUT4AB/E6BEG[6] Tile_X4Y8_LUT4AB/E6BEG[7] Tile_X4Y8_LUT4AB/E6BEG[8]
+ Tile_X4Y8_LUT4AB/E6BEG[9] Tile_X4Y8_LUT4AB/E6END[0] Tile_X4Y8_LUT4AB/E6END[10] Tile_X4Y8_LUT4AB/E6END[11]
+ Tile_X4Y8_LUT4AB/E6END[1] Tile_X4Y8_LUT4AB/E6END[2] Tile_X4Y8_LUT4AB/E6END[3] Tile_X4Y8_LUT4AB/E6END[4]
+ Tile_X4Y8_LUT4AB/E6END[5] Tile_X4Y8_LUT4AB/E6END[6] Tile_X4Y8_LUT4AB/E6END[7] Tile_X4Y8_LUT4AB/E6END[8]
+ Tile_X4Y8_LUT4AB/E6END[9] Tile_X4Y8_LUT4AB/EE4BEG[0] Tile_X4Y8_LUT4AB/EE4BEG[10]
+ Tile_X4Y8_LUT4AB/EE4BEG[11] Tile_X4Y8_LUT4AB/EE4BEG[12] Tile_X4Y8_LUT4AB/EE4BEG[13]
+ Tile_X4Y8_LUT4AB/EE4BEG[14] Tile_X4Y8_LUT4AB/EE4BEG[15] Tile_X4Y8_LUT4AB/EE4BEG[1]
+ Tile_X4Y8_LUT4AB/EE4BEG[2] Tile_X4Y8_LUT4AB/EE4BEG[3] Tile_X4Y8_LUT4AB/EE4BEG[4]
+ Tile_X4Y8_LUT4AB/EE4BEG[5] Tile_X4Y8_LUT4AB/EE4BEG[6] Tile_X4Y8_LUT4AB/EE4BEG[7]
+ Tile_X4Y8_LUT4AB/EE4BEG[8] Tile_X4Y8_LUT4AB/EE4BEG[9] Tile_X4Y8_LUT4AB/EE4END[0]
+ Tile_X4Y8_LUT4AB/EE4END[10] Tile_X4Y8_LUT4AB/EE4END[11] Tile_X4Y8_LUT4AB/EE4END[12]
+ Tile_X4Y8_LUT4AB/EE4END[13] Tile_X4Y8_LUT4AB/EE4END[14] Tile_X4Y8_LUT4AB/EE4END[15]
+ Tile_X4Y8_LUT4AB/EE4END[1] Tile_X4Y8_LUT4AB/EE4END[2] Tile_X4Y8_LUT4AB/EE4END[3]
+ Tile_X4Y8_LUT4AB/EE4END[4] Tile_X4Y8_LUT4AB/EE4END[5] Tile_X4Y8_LUT4AB/EE4END[6]
+ Tile_X4Y8_LUT4AB/EE4END[7] Tile_X4Y8_LUT4AB/EE4END[8] Tile_X4Y8_LUT4AB/EE4END[9]
+ Tile_X4Y8_LUT4AB/FrameData[0] Tile_X4Y8_LUT4AB/FrameData[10] Tile_X4Y8_LUT4AB/FrameData[11]
+ Tile_X4Y8_LUT4AB/FrameData[12] Tile_X4Y8_LUT4AB/FrameData[13] Tile_X4Y8_LUT4AB/FrameData[14]
+ Tile_X4Y8_LUT4AB/FrameData[15] Tile_X4Y8_LUT4AB/FrameData[16] Tile_X4Y8_LUT4AB/FrameData[17]
+ Tile_X4Y8_LUT4AB/FrameData[18] Tile_X4Y8_LUT4AB/FrameData[19] Tile_X4Y8_LUT4AB/FrameData[1]
+ Tile_X4Y8_LUT4AB/FrameData[20] Tile_X4Y8_LUT4AB/FrameData[21] Tile_X4Y8_LUT4AB/FrameData[22]
+ Tile_X4Y8_LUT4AB/FrameData[23] Tile_X4Y8_LUT4AB/FrameData[24] Tile_X4Y8_LUT4AB/FrameData[25]
+ Tile_X4Y8_LUT4AB/FrameData[26] Tile_X4Y8_LUT4AB/FrameData[27] Tile_X4Y8_LUT4AB/FrameData[28]
+ Tile_X4Y8_LUT4AB/FrameData[29] Tile_X4Y8_LUT4AB/FrameData[2] Tile_X4Y8_LUT4AB/FrameData[30]
+ Tile_X4Y8_LUT4AB/FrameData[31] Tile_X4Y8_LUT4AB/FrameData[3] Tile_X4Y8_LUT4AB/FrameData[4]
+ Tile_X4Y8_LUT4AB/FrameData[5] Tile_X4Y8_LUT4AB/FrameData[6] Tile_X4Y8_LUT4AB/FrameData[7]
+ Tile_X4Y8_LUT4AB/FrameData[8] Tile_X4Y8_LUT4AB/FrameData[9] Tile_X5Y8_E_TT_IF/FrameData[0]
+ Tile_X5Y8_E_TT_IF/FrameData[10] Tile_X5Y8_E_TT_IF/FrameData[11] Tile_X5Y8_E_TT_IF/FrameData[12]
+ Tile_X5Y8_E_TT_IF/FrameData[13] Tile_X5Y8_E_TT_IF/FrameData[14] Tile_X5Y8_E_TT_IF/FrameData[15]
+ Tile_X5Y8_E_TT_IF/FrameData[16] Tile_X5Y8_E_TT_IF/FrameData[17] Tile_X5Y8_E_TT_IF/FrameData[18]
+ Tile_X5Y8_E_TT_IF/FrameData[19] Tile_X5Y8_E_TT_IF/FrameData[1] Tile_X5Y8_E_TT_IF/FrameData[20]
+ Tile_X5Y8_E_TT_IF/FrameData[21] Tile_X5Y8_E_TT_IF/FrameData[22] Tile_X5Y8_E_TT_IF/FrameData[23]
+ Tile_X5Y8_E_TT_IF/FrameData[24] Tile_X5Y8_E_TT_IF/FrameData[25] Tile_X5Y8_E_TT_IF/FrameData[26]
+ Tile_X5Y8_E_TT_IF/FrameData[27] Tile_X5Y8_E_TT_IF/FrameData[28] Tile_X5Y8_E_TT_IF/FrameData[29]
+ Tile_X5Y8_E_TT_IF/FrameData[2] Tile_X5Y8_E_TT_IF/FrameData[30] Tile_X5Y8_E_TT_IF/FrameData[31]
+ Tile_X5Y8_E_TT_IF/FrameData[3] Tile_X5Y8_E_TT_IF/FrameData[4] Tile_X5Y8_E_TT_IF/FrameData[5]
+ Tile_X5Y8_E_TT_IF/FrameData[6] Tile_X5Y8_E_TT_IF/FrameData[7] Tile_X5Y8_E_TT_IF/FrameData[8]
+ Tile_X5Y8_E_TT_IF/FrameData[9] Tile_X4Y8_LUT4AB/FrameStrobe[0] Tile_X4Y8_LUT4AB/FrameStrobe[10]
+ Tile_X4Y8_LUT4AB/FrameStrobe[11] Tile_X4Y8_LUT4AB/FrameStrobe[12] Tile_X4Y8_LUT4AB/FrameStrobe[13]
+ Tile_X4Y8_LUT4AB/FrameStrobe[14] Tile_X4Y8_LUT4AB/FrameStrobe[15] Tile_X4Y8_LUT4AB/FrameStrobe[16]
+ Tile_X4Y8_LUT4AB/FrameStrobe[17] Tile_X4Y8_LUT4AB/FrameStrobe[18] Tile_X4Y8_LUT4AB/FrameStrobe[19]
+ Tile_X4Y8_LUT4AB/FrameStrobe[1] Tile_X4Y8_LUT4AB/FrameStrobe[2] Tile_X4Y8_LUT4AB/FrameStrobe[3]
+ Tile_X4Y8_LUT4AB/FrameStrobe[4] Tile_X4Y8_LUT4AB/FrameStrobe[5] Tile_X4Y8_LUT4AB/FrameStrobe[6]
+ Tile_X4Y8_LUT4AB/FrameStrobe[7] Tile_X4Y8_LUT4AB/FrameStrobe[8] Tile_X4Y8_LUT4AB/FrameStrobe[9]
+ Tile_X4Y7_LUT4AB/FrameStrobe[0] Tile_X4Y7_LUT4AB/FrameStrobe[10] Tile_X4Y7_LUT4AB/FrameStrobe[11]
+ Tile_X4Y7_LUT4AB/FrameStrobe[12] Tile_X4Y7_LUT4AB/FrameStrobe[13] Tile_X4Y7_LUT4AB/FrameStrobe[14]
+ Tile_X4Y7_LUT4AB/FrameStrobe[15] Tile_X4Y7_LUT4AB/FrameStrobe[16] Tile_X4Y7_LUT4AB/FrameStrobe[17]
+ Tile_X4Y7_LUT4AB/FrameStrobe[18] Tile_X4Y7_LUT4AB/FrameStrobe[19] Tile_X4Y7_LUT4AB/FrameStrobe[1]
+ Tile_X4Y7_LUT4AB/FrameStrobe[2] Tile_X4Y7_LUT4AB/FrameStrobe[3] Tile_X4Y7_LUT4AB/FrameStrobe[4]
+ Tile_X4Y7_LUT4AB/FrameStrobe[5] Tile_X4Y7_LUT4AB/FrameStrobe[6] Tile_X4Y7_LUT4AB/FrameStrobe[7]
+ Tile_X4Y7_LUT4AB/FrameStrobe[8] Tile_X4Y7_LUT4AB/FrameStrobe[9] Tile_X4Y8_LUT4AB/N1BEG[0]
+ Tile_X4Y8_LUT4AB/N1BEG[1] Tile_X4Y8_LUT4AB/N1BEG[2] Tile_X4Y8_LUT4AB/N1BEG[3] Tile_X4Y9_S_IO4/N1BEG[0]
+ Tile_X4Y9_S_IO4/N1BEG[1] Tile_X4Y9_S_IO4/N1BEG[2] Tile_X4Y9_S_IO4/N1BEG[3] Tile_X4Y8_LUT4AB/N2BEG[0]
+ Tile_X4Y8_LUT4AB/N2BEG[1] Tile_X4Y8_LUT4AB/N2BEG[2] Tile_X4Y8_LUT4AB/N2BEG[3] Tile_X4Y8_LUT4AB/N2BEG[4]
+ Tile_X4Y8_LUT4AB/N2BEG[5] Tile_X4Y8_LUT4AB/N2BEG[6] Tile_X4Y8_LUT4AB/N2BEG[7] Tile_X4Y7_LUT4AB/N2END[0]
+ Tile_X4Y7_LUT4AB/N2END[1] Tile_X4Y7_LUT4AB/N2END[2] Tile_X4Y7_LUT4AB/N2END[3] Tile_X4Y7_LUT4AB/N2END[4]
+ Tile_X4Y7_LUT4AB/N2END[5] Tile_X4Y7_LUT4AB/N2END[6] Tile_X4Y7_LUT4AB/N2END[7] Tile_X4Y9_S_IO4/N2BEGb[0]
+ Tile_X4Y9_S_IO4/N2BEGb[1] Tile_X4Y9_S_IO4/N2BEGb[2] Tile_X4Y9_S_IO4/N2BEGb[3] Tile_X4Y9_S_IO4/N2BEGb[4]
+ Tile_X4Y9_S_IO4/N2BEGb[5] Tile_X4Y9_S_IO4/N2BEGb[6] Tile_X4Y9_S_IO4/N2BEGb[7] Tile_X4Y9_S_IO4/N2BEG[0]
+ Tile_X4Y9_S_IO4/N2BEG[1] Tile_X4Y9_S_IO4/N2BEG[2] Tile_X4Y9_S_IO4/N2BEG[3] Tile_X4Y9_S_IO4/N2BEG[4]
+ Tile_X4Y9_S_IO4/N2BEG[5] Tile_X4Y9_S_IO4/N2BEG[6] Tile_X4Y9_S_IO4/N2BEG[7] Tile_X4Y8_LUT4AB/N4BEG[0]
+ Tile_X4Y8_LUT4AB/N4BEG[10] Tile_X4Y8_LUT4AB/N4BEG[11] Tile_X4Y8_LUT4AB/N4BEG[12]
+ Tile_X4Y8_LUT4AB/N4BEG[13] Tile_X4Y8_LUT4AB/N4BEG[14] Tile_X4Y8_LUT4AB/N4BEG[15]
+ Tile_X4Y8_LUT4AB/N4BEG[1] Tile_X4Y8_LUT4AB/N4BEG[2] Tile_X4Y8_LUT4AB/N4BEG[3] Tile_X4Y8_LUT4AB/N4BEG[4]
+ Tile_X4Y8_LUT4AB/N4BEG[5] Tile_X4Y8_LUT4AB/N4BEG[6] Tile_X4Y8_LUT4AB/N4BEG[7] Tile_X4Y8_LUT4AB/N4BEG[8]
+ Tile_X4Y8_LUT4AB/N4BEG[9] Tile_X4Y9_S_IO4/N4BEG[0] Tile_X4Y9_S_IO4/N4BEG[10] Tile_X4Y9_S_IO4/N4BEG[11]
+ Tile_X4Y9_S_IO4/N4BEG[12] Tile_X4Y9_S_IO4/N4BEG[13] Tile_X4Y9_S_IO4/N4BEG[14] Tile_X4Y9_S_IO4/N4BEG[15]
+ Tile_X4Y9_S_IO4/N4BEG[1] Tile_X4Y9_S_IO4/N4BEG[2] Tile_X4Y9_S_IO4/N4BEG[3] Tile_X4Y9_S_IO4/N4BEG[4]
+ Tile_X4Y9_S_IO4/N4BEG[5] Tile_X4Y9_S_IO4/N4BEG[6] Tile_X4Y9_S_IO4/N4BEG[7] Tile_X4Y9_S_IO4/N4BEG[8]
+ Tile_X4Y9_S_IO4/N4BEG[9] Tile_X4Y8_LUT4AB/NN4BEG[0] Tile_X4Y8_LUT4AB/NN4BEG[10]
+ Tile_X4Y8_LUT4AB/NN4BEG[11] Tile_X4Y8_LUT4AB/NN4BEG[12] Tile_X4Y8_LUT4AB/NN4BEG[13]
+ Tile_X4Y8_LUT4AB/NN4BEG[14] Tile_X4Y8_LUT4AB/NN4BEG[15] Tile_X4Y8_LUT4AB/NN4BEG[1]
+ Tile_X4Y8_LUT4AB/NN4BEG[2] Tile_X4Y8_LUT4AB/NN4BEG[3] Tile_X4Y8_LUT4AB/NN4BEG[4]
+ Tile_X4Y8_LUT4AB/NN4BEG[5] Tile_X4Y8_LUT4AB/NN4BEG[6] Tile_X4Y8_LUT4AB/NN4BEG[7]
+ Tile_X4Y8_LUT4AB/NN4BEG[8] Tile_X4Y8_LUT4AB/NN4BEG[9] Tile_X4Y9_S_IO4/NN4BEG[0]
+ Tile_X4Y9_S_IO4/NN4BEG[10] Tile_X4Y9_S_IO4/NN4BEG[11] Tile_X4Y9_S_IO4/NN4BEG[12]
+ Tile_X4Y9_S_IO4/NN4BEG[13] Tile_X4Y9_S_IO4/NN4BEG[14] Tile_X4Y9_S_IO4/NN4BEG[15]
+ Tile_X4Y9_S_IO4/NN4BEG[1] Tile_X4Y9_S_IO4/NN4BEG[2] Tile_X4Y9_S_IO4/NN4BEG[3] Tile_X4Y9_S_IO4/NN4BEG[4]
+ Tile_X4Y9_S_IO4/NN4BEG[5] Tile_X4Y9_S_IO4/NN4BEG[6] Tile_X4Y9_S_IO4/NN4BEG[7] Tile_X4Y9_S_IO4/NN4BEG[8]
+ Tile_X4Y9_S_IO4/NN4BEG[9] Tile_X4Y9_S_IO4/S1END[0] Tile_X4Y9_S_IO4/S1END[1] Tile_X4Y9_S_IO4/S1END[2]
+ Tile_X4Y9_S_IO4/S1END[3] Tile_X4Y8_LUT4AB/S1END[0] Tile_X4Y8_LUT4AB/S1END[1] Tile_X4Y8_LUT4AB/S1END[2]
+ Tile_X4Y8_LUT4AB/S1END[3] Tile_X4Y9_S_IO4/S2MID[0] Tile_X4Y9_S_IO4/S2MID[1] Tile_X4Y9_S_IO4/S2MID[2]
+ Tile_X4Y9_S_IO4/S2MID[3] Tile_X4Y9_S_IO4/S2MID[4] Tile_X4Y9_S_IO4/S2MID[5] Tile_X4Y9_S_IO4/S2MID[6]
+ Tile_X4Y9_S_IO4/S2MID[7] Tile_X4Y9_S_IO4/S2END[0] Tile_X4Y9_S_IO4/S2END[1] Tile_X4Y9_S_IO4/S2END[2]
+ Tile_X4Y9_S_IO4/S2END[3] Tile_X4Y9_S_IO4/S2END[4] Tile_X4Y9_S_IO4/S2END[5] Tile_X4Y9_S_IO4/S2END[6]
+ Tile_X4Y9_S_IO4/S2END[7] Tile_X4Y8_LUT4AB/S2END[0] Tile_X4Y8_LUT4AB/S2END[1] Tile_X4Y8_LUT4AB/S2END[2]
+ Tile_X4Y8_LUT4AB/S2END[3] Tile_X4Y8_LUT4AB/S2END[4] Tile_X4Y8_LUT4AB/S2END[5] Tile_X4Y8_LUT4AB/S2END[6]
+ Tile_X4Y8_LUT4AB/S2END[7] Tile_X4Y8_LUT4AB/S2MID[0] Tile_X4Y8_LUT4AB/S2MID[1] Tile_X4Y8_LUT4AB/S2MID[2]
+ Tile_X4Y8_LUT4AB/S2MID[3] Tile_X4Y8_LUT4AB/S2MID[4] Tile_X4Y8_LUT4AB/S2MID[5] Tile_X4Y8_LUT4AB/S2MID[6]
+ Tile_X4Y8_LUT4AB/S2MID[7] Tile_X4Y9_S_IO4/S4END[0] Tile_X4Y9_S_IO4/S4END[10] Tile_X4Y9_S_IO4/S4END[11]
+ Tile_X4Y9_S_IO4/S4END[12] Tile_X4Y9_S_IO4/S4END[13] Tile_X4Y9_S_IO4/S4END[14] Tile_X4Y9_S_IO4/S4END[15]
+ Tile_X4Y9_S_IO4/S4END[1] Tile_X4Y9_S_IO4/S4END[2] Tile_X4Y9_S_IO4/S4END[3] Tile_X4Y9_S_IO4/S4END[4]
+ Tile_X4Y9_S_IO4/S4END[5] Tile_X4Y9_S_IO4/S4END[6] Tile_X4Y9_S_IO4/S4END[7] Tile_X4Y9_S_IO4/S4END[8]
+ Tile_X4Y9_S_IO4/S4END[9] Tile_X4Y8_LUT4AB/S4END[0] Tile_X4Y8_LUT4AB/S4END[10] Tile_X4Y8_LUT4AB/S4END[11]
+ Tile_X4Y8_LUT4AB/S4END[12] Tile_X4Y8_LUT4AB/S4END[13] Tile_X4Y8_LUT4AB/S4END[14]
+ Tile_X4Y8_LUT4AB/S4END[15] Tile_X4Y8_LUT4AB/S4END[1] Tile_X4Y8_LUT4AB/S4END[2] Tile_X4Y8_LUT4AB/S4END[3]
+ Tile_X4Y8_LUT4AB/S4END[4] Tile_X4Y8_LUT4AB/S4END[5] Tile_X4Y8_LUT4AB/S4END[6] Tile_X4Y8_LUT4AB/S4END[7]
+ Tile_X4Y8_LUT4AB/S4END[8] Tile_X4Y8_LUT4AB/S4END[9] Tile_X4Y9_S_IO4/SS4END[0] Tile_X4Y9_S_IO4/SS4END[10]
+ Tile_X4Y9_S_IO4/SS4END[11] Tile_X4Y9_S_IO4/SS4END[12] Tile_X4Y9_S_IO4/SS4END[13]
+ Tile_X4Y9_S_IO4/SS4END[14] Tile_X4Y9_S_IO4/SS4END[15] Tile_X4Y9_S_IO4/SS4END[1]
+ Tile_X4Y9_S_IO4/SS4END[2] Tile_X4Y9_S_IO4/SS4END[3] Tile_X4Y9_S_IO4/SS4END[4] Tile_X4Y9_S_IO4/SS4END[5]
+ Tile_X4Y9_S_IO4/SS4END[6] Tile_X4Y9_S_IO4/SS4END[7] Tile_X4Y9_S_IO4/SS4END[8] Tile_X4Y9_S_IO4/SS4END[9]
+ Tile_X4Y8_LUT4AB/SS4END[0] Tile_X4Y8_LUT4AB/SS4END[10] Tile_X4Y8_LUT4AB/SS4END[11]
+ Tile_X4Y8_LUT4AB/SS4END[12] Tile_X4Y8_LUT4AB/SS4END[13] Tile_X4Y8_LUT4AB/SS4END[14]
+ Tile_X4Y8_LUT4AB/SS4END[15] Tile_X4Y8_LUT4AB/SS4END[1] Tile_X4Y8_LUT4AB/SS4END[2]
+ Tile_X4Y8_LUT4AB/SS4END[3] Tile_X4Y8_LUT4AB/SS4END[4] Tile_X4Y8_LUT4AB/SS4END[5]
+ Tile_X4Y8_LUT4AB/SS4END[6] Tile_X4Y8_LUT4AB/SS4END[7] Tile_X4Y8_LUT4AB/SS4END[8]
+ Tile_X4Y8_LUT4AB/SS4END[9] Tile_X4Y9_S_IO4/UserCLKo Tile_X4Y7_LUT4AB/UserCLK VGND
+ VPWR Tile_X4Y8_LUT4AB/W1BEG[0] Tile_X4Y8_LUT4AB/W1BEG[1] Tile_X4Y8_LUT4AB/W1BEG[2]
+ Tile_X4Y8_LUT4AB/W1BEG[3] Tile_X4Y8_LUT4AB/W1END[0] Tile_X4Y8_LUT4AB/W1END[1] Tile_X4Y8_LUT4AB/W1END[2]
+ Tile_X4Y8_LUT4AB/W1END[3] Tile_X4Y8_LUT4AB/W2BEG[0] Tile_X4Y8_LUT4AB/W2BEG[1] Tile_X4Y8_LUT4AB/W2BEG[2]
+ Tile_X4Y8_LUT4AB/W2BEG[3] Tile_X4Y8_LUT4AB/W2BEG[4] Tile_X4Y8_LUT4AB/W2BEG[5] Tile_X4Y8_LUT4AB/W2BEG[6]
+ Tile_X4Y8_LUT4AB/W2BEG[7] Tile_X3Y8_LUT4AB/W2END[0] Tile_X3Y8_LUT4AB/W2END[1] Tile_X3Y8_LUT4AB/W2END[2]
+ Tile_X3Y8_LUT4AB/W2END[3] Tile_X3Y8_LUT4AB/W2END[4] Tile_X3Y8_LUT4AB/W2END[5] Tile_X3Y8_LUT4AB/W2END[6]
+ Tile_X3Y8_LUT4AB/W2END[7] Tile_X4Y8_LUT4AB/W2END[0] Tile_X4Y8_LUT4AB/W2END[1] Tile_X4Y8_LUT4AB/W2END[2]
+ Tile_X4Y8_LUT4AB/W2END[3] Tile_X4Y8_LUT4AB/W2END[4] Tile_X4Y8_LUT4AB/W2END[5] Tile_X4Y8_LUT4AB/W2END[6]
+ Tile_X4Y8_LUT4AB/W2END[7] Tile_X4Y8_LUT4AB/W2MID[0] Tile_X4Y8_LUT4AB/W2MID[1] Tile_X4Y8_LUT4AB/W2MID[2]
+ Tile_X4Y8_LUT4AB/W2MID[3] Tile_X4Y8_LUT4AB/W2MID[4] Tile_X4Y8_LUT4AB/W2MID[5] Tile_X4Y8_LUT4AB/W2MID[6]
+ Tile_X4Y8_LUT4AB/W2MID[7] Tile_X4Y8_LUT4AB/W6BEG[0] Tile_X4Y8_LUT4AB/W6BEG[10] Tile_X4Y8_LUT4AB/W6BEG[11]
+ Tile_X4Y8_LUT4AB/W6BEG[1] Tile_X4Y8_LUT4AB/W6BEG[2] Tile_X4Y8_LUT4AB/W6BEG[3] Tile_X4Y8_LUT4AB/W6BEG[4]
+ Tile_X4Y8_LUT4AB/W6BEG[5] Tile_X4Y8_LUT4AB/W6BEG[6] Tile_X4Y8_LUT4AB/W6BEG[7] Tile_X4Y8_LUT4AB/W6BEG[8]
+ Tile_X4Y8_LUT4AB/W6BEG[9] Tile_X4Y8_LUT4AB/W6END[0] Tile_X4Y8_LUT4AB/W6END[10] Tile_X4Y8_LUT4AB/W6END[11]
+ Tile_X4Y8_LUT4AB/W6END[1] Tile_X4Y8_LUT4AB/W6END[2] Tile_X4Y8_LUT4AB/W6END[3] Tile_X4Y8_LUT4AB/W6END[4]
+ Tile_X4Y8_LUT4AB/W6END[5] Tile_X4Y8_LUT4AB/W6END[6] Tile_X4Y8_LUT4AB/W6END[7] Tile_X4Y8_LUT4AB/W6END[8]
+ Tile_X4Y8_LUT4AB/W6END[9] Tile_X4Y8_LUT4AB/WW4BEG[0] Tile_X4Y8_LUT4AB/WW4BEG[10]
+ Tile_X4Y8_LUT4AB/WW4BEG[11] Tile_X4Y8_LUT4AB/WW4BEG[12] Tile_X4Y8_LUT4AB/WW4BEG[13]
+ Tile_X4Y8_LUT4AB/WW4BEG[14] Tile_X4Y8_LUT4AB/WW4BEG[15] Tile_X4Y8_LUT4AB/WW4BEG[1]
+ Tile_X4Y8_LUT4AB/WW4BEG[2] Tile_X4Y8_LUT4AB/WW4BEG[3] Tile_X4Y8_LUT4AB/WW4BEG[4]
+ Tile_X4Y8_LUT4AB/WW4BEG[5] Tile_X4Y8_LUT4AB/WW4BEG[6] Tile_X4Y8_LUT4AB/WW4BEG[7]
+ Tile_X4Y8_LUT4AB/WW4BEG[8] Tile_X4Y8_LUT4AB/WW4BEG[9] Tile_X4Y8_LUT4AB/WW4END[0]
+ Tile_X4Y8_LUT4AB/WW4END[10] Tile_X4Y8_LUT4AB/WW4END[11] Tile_X4Y8_LUT4AB/WW4END[12]
+ Tile_X4Y8_LUT4AB/WW4END[13] Tile_X4Y8_LUT4AB/WW4END[14] Tile_X4Y8_LUT4AB/WW4END[15]
+ Tile_X4Y8_LUT4AB/WW4END[1] Tile_X4Y8_LUT4AB/WW4END[2] Tile_X4Y8_LUT4AB/WW4END[3]
+ Tile_X4Y8_LUT4AB/WW4END[4] Tile_X4Y8_LUT4AB/WW4END[5] Tile_X4Y8_LUT4AB/WW4END[6]
+ Tile_X4Y8_LUT4AB/WW4END[7] Tile_X4Y8_LUT4AB/WW4END[8] Tile_X4Y8_LUT4AB/WW4END[9]
+ LUT4AB
XTile_X1Y9_S_IO4 Tile_X1Y9_A_I_top Tile_X1Y9_A_O_top Tile_X1Y9_A_T_top Tile_X1Y9_B_I_top
+ Tile_X1Y9_B_O_top Tile_X1Y9_B_T_top Tile_X1Y9_C_I_top Tile_X1Y9_C_O_top Tile_X1Y9_C_T_top
+ Tile_X1Y9_S_IO4/Co Tile_X1Y9_D_I_top Tile_X1Y9_D_O_top Tile_X1Y9_D_T_top Tile_X1Y9_S_IO4/FrameData[0]
+ Tile_X1Y9_S_IO4/FrameData[10] Tile_X1Y9_S_IO4/FrameData[11] Tile_X1Y9_S_IO4/FrameData[12]
+ Tile_X1Y9_S_IO4/FrameData[13] Tile_X1Y9_S_IO4/FrameData[14] Tile_X1Y9_S_IO4/FrameData[15]
+ Tile_X1Y9_S_IO4/FrameData[16] Tile_X1Y9_S_IO4/FrameData[17] Tile_X1Y9_S_IO4/FrameData[18]
+ Tile_X1Y9_S_IO4/FrameData[19] Tile_X1Y9_S_IO4/FrameData[1] Tile_X1Y9_S_IO4/FrameData[20]
+ Tile_X1Y9_S_IO4/FrameData[21] Tile_X1Y9_S_IO4/FrameData[22] Tile_X1Y9_S_IO4/FrameData[23]
+ Tile_X1Y9_S_IO4/FrameData[24] Tile_X1Y9_S_IO4/FrameData[25] Tile_X1Y9_S_IO4/FrameData[26]
+ Tile_X1Y9_S_IO4/FrameData[27] Tile_X1Y9_S_IO4/FrameData[28] Tile_X1Y9_S_IO4/FrameData[29]
+ Tile_X1Y9_S_IO4/FrameData[2] Tile_X1Y9_S_IO4/FrameData[30] Tile_X1Y9_S_IO4/FrameData[31]
+ Tile_X1Y9_S_IO4/FrameData[3] Tile_X1Y9_S_IO4/FrameData[4] Tile_X1Y9_S_IO4/FrameData[5]
+ Tile_X1Y9_S_IO4/FrameData[6] Tile_X1Y9_S_IO4/FrameData[7] Tile_X1Y9_S_IO4/FrameData[8]
+ Tile_X1Y9_S_IO4/FrameData[9] Tile_X2Y9_S_IO4/FrameData[0] Tile_X2Y9_S_IO4/FrameData[10]
+ Tile_X2Y9_S_IO4/FrameData[11] Tile_X2Y9_S_IO4/FrameData[12] Tile_X2Y9_S_IO4/FrameData[13]
+ Tile_X2Y9_S_IO4/FrameData[14] Tile_X2Y9_S_IO4/FrameData[15] Tile_X2Y9_S_IO4/FrameData[16]
+ Tile_X2Y9_S_IO4/FrameData[17] Tile_X2Y9_S_IO4/FrameData[18] Tile_X2Y9_S_IO4/FrameData[19]
+ Tile_X2Y9_S_IO4/FrameData[1] Tile_X2Y9_S_IO4/FrameData[20] Tile_X2Y9_S_IO4/FrameData[21]
+ Tile_X2Y9_S_IO4/FrameData[22] Tile_X2Y9_S_IO4/FrameData[23] Tile_X2Y9_S_IO4/FrameData[24]
+ Tile_X2Y9_S_IO4/FrameData[25] Tile_X2Y9_S_IO4/FrameData[26] Tile_X2Y9_S_IO4/FrameData[27]
+ Tile_X2Y9_S_IO4/FrameData[28] Tile_X2Y9_S_IO4/FrameData[29] Tile_X2Y9_S_IO4/FrameData[2]
+ Tile_X2Y9_S_IO4/FrameData[30] Tile_X2Y9_S_IO4/FrameData[31] Tile_X2Y9_S_IO4/FrameData[3]
+ Tile_X2Y9_S_IO4/FrameData[4] Tile_X2Y9_S_IO4/FrameData[5] Tile_X2Y9_S_IO4/FrameData[6]
+ Tile_X2Y9_S_IO4/FrameData[7] Tile_X2Y9_S_IO4/FrameData[8] Tile_X2Y9_S_IO4/FrameData[9]
+ FrameStrobe[20] FrameStrobe[30] FrameStrobe[31] FrameStrobe[32] FrameStrobe[33]
+ FrameStrobe[34] FrameStrobe[35] FrameStrobe[36] FrameStrobe[37] FrameStrobe[38]
+ FrameStrobe[39] FrameStrobe[21] FrameStrobe[22] FrameStrobe[23] FrameStrobe[24]
+ FrameStrobe[25] FrameStrobe[26] FrameStrobe[27] FrameStrobe[28] FrameStrobe[29]
+ Tile_X1Y8_LUT4AB/FrameStrobe[0] Tile_X1Y8_LUT4AB/FrameStrobe[10] Tile_X1Y8_LUT4AB/FrameStrobe[11]
+ Tile_X1Y8_LUT4AB/FrameStrobe[12] Tile_X1Y8_LUT4AB/FrameStrobe[13] Tile_X1Y8_LUT4AB/FrameStrobe[14]
+ Tile_X1Y8_LUT4AB/FrameStrobe[15] Tile_X1Y8_LUT4AB/FrameStrobe[16] Tile_X1Y8_LUT4AB/FrameStrobe[17]
+ Tile_X1Y8_LUT4AB/FrameStrobe[18] Tile_X1Y8_LUT4AB/FrameStrobe[19] Tile_X1Y8_LUT4AB/FrameStrobe[1]
+ Tile_X1Y8_LUT4AB/FrameStrobe[2] Tile_X1Y8_LUT4AB/FrameStrobe[3] Tile_X1Y8_LUT4AB/FrameStrobe[4]
+ Tile_X1Y8_LUT4AB/FrameStrobe[5] Tile_X1Y8_LUT4AB/FrameStrobe[6] Tile_X1Y8_LUT4AB/FrameStrobe[7]
+ Tile_X1Y8_LUT4AB/FrameStrobe[8] Tile_X1Y8_LUT4AB/FrameStrobe[9] Tile_X1Y9_S_IO4/N1BEG[0]
+ Tile_X1Y9_S_IO4/N1BEG[1] Tile_X1Y9_S_IO4/N1BEG[2] Tile_X1Y9_S_IO4/N1BEG[3] Tile_X1Y9_S_IO4/N2BEG[0]
+ Tile_X1Y9_S_IO4/N2BEG[1] Tile_X1Y9_S_IO4/N2BEG[2] Tile_X1Y9_S_IO4/N2BEG[3] Tile_X1Y9_S_IO4/N2BEG[4]
+ Tile_X1Y9_S_IO4/N2BEG[5] Tile_X1Y9_S_IO4/N2BEG[6] Tile_X1Y9_S_IO4/N2BEG[7] Tile_X1Y9_S_IO4/N2BEGb[0]
+ Tile_X1Y9_S_IO4/N2BEGb[1] Tile_X1Y9_S_IO4/N2BEGb[2] Tile_X1Y9_S_IO4/N2BEGb[3] Tile_X1Y9_S_IO4/N2BEGb[4]
+ Tile_X1Y9_S_IO4/N2BEGb[5] Tile_X1Y9_S_IO4/N2BEGb[6] Tile_X1Y9_S_IO4/N2BEGb[7] Tile_X1Y9_S_IO4/N4BEG[0]
+ Tile_X1Y9_S_IO4/N4BEG[10] Tile_X1Y9_S_IO4/N4BEG[11] Tile_X1Y9_S_IO4/N4BEG[12] Tile_X1Y9_S_IO4/N4BEG[13]
+ Tile_X1Y9_S_IO4/N4BEG[14] Tile_X1Y9_S_IO4/N4BEG[15] Tile_X1Y9_S_IO4/N4BEG[1] Tile_X1Y9_S_IO4/N4BEG[2]
+ Tile_X1Y9_S_IO4/N4BEG[3] Tile_X1Y9_S_IO4/N4BEG[4] Tile_X1Y9_S_IO4/N4BEG[5] Tile_X1Y9_S_IO4/N4BEG[6]
+ Tile_X1Y9_S_IO4/N4BEG[7] Tile_X1Y9_S_IO4/N4BEG[8] Tile_X1Y9_S_IO4/N4BEG[9] Tile_X1Y9_S_IO4/NN4BEG[0]
+ Tile_X1Y9_S_IO4/NN4BEG[10] Tile_X1Y9_S_IO4/NN4BEG[11] Tile_X1Y9_S_IO4/NN4BEG[12]
+ Tile_X1Y9_S_IO4/NN4BEG[13] Tile_X1Y9_S_IO4/NN4BEG[14] Tile_X1Y9_S_IO4/NN4BEG[15]
+ Tile_X1Y9_S_IO4/NN4BEG[1] Tile_X1Y9_S_IO4/NN4BEG[2] Tile_X1Y9_S_IO4/NN4BEG[3] Tile_X1Y9_S_IO4/NN4BEG[4]
+ Tile_X1Y9_S_IO4/NN4BEG[5] Tile_X1Y9_S_IO4/NN4BEG[6] Tile_X1Y9_S_IO4/NN4BEG[7] Tile_X1Y9_S_IO4/NN4BEG[8]
+ Tile_X1Y9_S_IO4/NN4BEG[9] Tile_X1Y9_S_IO4/S1END[0] Tile_X1Y9_S_IO4/S1END[1] Tile_X1Y9_S_IO4/S1END[2]
+ Tile_X1Y9_S_IO4/S1END[3] Tile_X1Y9_S_IO4/S2END[0] Tile_X1Y9_S_IO4/S2END[1] Tile_X1Y9_S_IO4/S2END[2]
+ Tile_X1Y9_S_IO4/S2END[3] Tile_X1Y9_S_IO4/S2END[4] Tile_X1Y9_S_IO4/S2END[5] Tile_X1Y9_S_IO4/S2END[6]
+ Tile_X1Y9_S_IO4/S2END[7] Tile_X1Y9_S_IO4/S2MID[0] Tile_X1Y9_S_IO4/S2MID[1] Tile_X1Y9_S_IO4/S2MID[2]
+ Tile_X1Y9_S_IO4/S2MID[3] Tile_X1Y9_S_IO4/S2MID[4] Tile_X1Y9_S_IO4/S2MID[5] Tile_X1Y9_S_IO4/S2MID[6]
+ Tile_X1Y9_S_IO4/S2MID[7] Tile_X1Y9_S_IO4/S4END[0] Tile_X1Y9_S_IO4/S4END[10] Tile_X1Y9_S_IO4/S4END[11]
+ Tile_X1Y9_S_IO4/S4END[12] Tile_X1Y9_S_IO4/S4END[13] Tile_X1Y9_S_IO4/S4END[14] Tile_X1Y9_S_IO4/S4END[15]
+ Tile_X1Y9_S_IO4/S4END[1] Tile_X1Y9_S_IO4/S4END[2] Tile_X1Y9_S_IO4/S4END[3] Tile_X1Y9_S_IO4/S4END[4]
+ Tile_X1Y9_S_IO4/S4END[5] Tile_X1Y9_S_IO4/S4END[6] Tile_X1Y9_S_IO4/S4END[7] Tile_X1Y9_S_IO4/S4END[8]
+ Tile_X1Y9_S_IO4/S4END[9] Tile_X1Y9_S_IO4/SS4END[0] Tile_X1Y9_S_IO4/SS4END[10] Tile_X1Y9_S_IO4/SS4END[11]
+ Tile_X1Y9_S_IO4/SS4END[12] Tile_X1Y9_S_IO4/SS4END[13] Tile_X1Y9_S_IO4/SS4END[14]
+ Tile_X1Y9_S_IO4/SS4END[15] Tile_X1Y9_S_IO4/SS4END[1] Tile_X1Y9_S_IO4/SS4END[2] Tile_X1Y9_S_IO4/SS4END[3]
+ Tile_X1Y9_S_IO4/SS4END[4] Tile_X1Y9_S_IO4/SS4END[5] Tile_X1Y9_S_IO4/SS4END[6] Tile_X1Y9_S_IO4/SS4END[7]
+ Tile_X1Y9_S_IO4/SS4END[8] Tile_X1Y9_S_IO4/SS4END[9] UserCLK Tile_X1Y9_S_IO4/UserCLKo
+ VGND VPWR S_IO4
XTile_X3Y1_LUT4AB Tile_X3Y2_LUT4AB/Co Tile_X3Y0_N_IO4/Ci Tile_X4Y1_LUT4AB/E1END[0]
+ Tile_X4Y1_LUT4AB/E1END[1] Tile_X4Y1_LUT4AB/E1END[2] Tile_X4Y1_LUT4AB/E1END[3] Tile_X3Y1_LUT4AB/E1END[0]
+ Tile_X3Y1_LUT4AB/E1END[1] Tile_X3Y1_LUT4AB/E1END[2] Tile_X3Y1_LUT4AB/E1END[3] Tile_X4Y1_LUT4AB/E2MID[0]
+ Tile_X4Y1_LUT4AB/E2MID[1] Tile_X4Y1_LUT4AB/E2MID[2] Tile_X4Y1_LUT4AB/E2MID[3] Tile_X4Y1_LUT4AB/E2MID[4]
+ Tile_X4Y1_LUT4AB/E2MID[5] Tile_X4Y1_LUT4AB/E2MID[6] Tile_X4Y1_LUT4AB/E2MID[7] Tile_X4Y1_LUT4AB/E2END[0]
+ Tile_X4Y1_LUT4AB/E2END[1] Tile_X4Y1_LUT4AB/E2END[2] Tile_X4Y1_LUT4AB/E2END[3] Tile_X4Y1_LUT4AB/E2END[4]
+ Tile_X4Y1_LUT4AB/E2END[5] Tile_X4Y1_LUT4AB/E2END[6] Tile_X4Y1_LUT4AB/E2END[7] Tile_X3Y1_LUT4AB/E2END[0]
+ Tile_X3Y1_LUT4AB/E2END[1] Tile_X3Y1_LUT4AB/E2END[2] Tile_X3Y1_LUT4AB/E2END[3] Tile_X3Y1_LUT4AB/E2END[4]
+ Tile_X3Y1_LUT4AB/E2END[5] Tile_X3Y1_LUT4AB/E2END[6] Tile_X3Y1_LUT4AB/E2END[7] Tile_X3Y1_LUT4AB/E2MID[0]
+ Tile_X3Y1_LUT4AB/E2MID[1] Tile_X3Y1_LUT4AB/E2MID[2] Tile_X3Y1_LUT4AB/E2MID[3] Tile_X3Y1_LUT4AB/E2MID[4]
+ Tile_X3Y1_LUT4AB/E2MID[5] Tile_X3Y1_LUT4AB/E2MID[6] Tile_X3Y1_LUT4AB/E2MID[7] Tile_X4Y1_LUT4AB/E6END[0]
+ Tile_X4Y1_LUT4AB/E6END[10] Tile_X4Y1_LUT4AB/E6END[11] Tile_X4Y1_LUT4AB/E6END[1]
+ Tile_X4Y1_LUT4AB/E6END[2] Tile_X4Y1_LUT4AB/E6END[3] Tile_X4Y1_LUT4AB/E6END[4] Tile_X4Y1_LUT4AB/E6END[5]
+ Tile_X4Y1_LUT4AB/E6END[6] Tile_X4Y1_LUT4AB/E6END[7] Tile_X4Y1_LUT4AB/E6END[8] Tile_X4Y1_LUT4AB/E6END[9]
+ Tile_X3Y1_LUT4AB/E6END[0] Tile_X3Y1_LUT4AB/E6END[10] Tile_X3Y1_LUT4AB/E6END[11]
+ Tile_X3Y1_LUT4AB/E6END[1] Tile_X3Y1_LUT4AB/E6END[2] Tile_X3Y1_LUT4AB/E6END[3] Tile_X3Y1_LUT4AB/E6END[4]
+ Tile_X3Y1_LUT4AB/E6END[5] Tile_X3Y1_LUT4AB/E6END[6] Tile_X3Y1_LUT4AB/E6END[7] Tile_X3Y1_LUT4AB/E6END[8]
+ Tile_X3Y1_LUT4AB/E6END[9] Tile_X4Y1_LUT4AB/EE4END[0] Tile_X4Y1_LUT4AB/EE4END[10]
+ Tile_X4Y1_LUT4AB/EE4END[11] Tile_X4Y1_LUT4AB/EE4END[12] Tile_X4Y1_LUT4AB/EE4END[13]
+ Tile_X4Y1_LUT4AB/EE4END[14] Tile_X4Y1_LUT4AB/EE4END[15] Tile_X4Y1_LUT4AB/EE4END[1]
+ Tile_X4Y1_LUT4AB/EE4END[2] Tile_X4Y1_LUT4AB/EE4END[3] Tile_X4Y1_LUT4AB/EE4END[4]
+ Tile_X4Y1_LUT4AB/EE4END[5] Tile_X4Y1_LUT4AB/EE4END[6] Tile_X4Y1_LUT4AB/EE4END[7]
+ Tile_X4Y1_LUT4AB/EE4END[8] Tile_X4Y1_LUT4AB/EE4END[9] Tile_X3Y1_LUT4AB/EE4END[0]
+ Tile_X3Y1_LUT4AB/EE4END[10] Tile_X3Y1_LUT4AB/EE4END[11] Tile_X3Y1_LUT4AB/EE4END[12]
+ Tile_X3Y1_LUT4AB/EE4END[13] Tile_X3Y1_LUT4AB/EE4END[14] Tile_X3Y1_LUT4AB/EE4END[15]
+ Tile_X3Y1_LUT4AB/EE4END[1] Tile_X3Y1_LUT4AB/EE4END[2] Tile_X3Y1_LUT4AB/EE4END[3]
+ Tile_X3Y1_LUT4AB/EE4END[4] Tile_X3Y1_LUT4AB/EE4END[5] Tile_X3Y1_LUT4AB/EE4END[6]
+ Tile_X3Y1_LUT4AB/EE4END[7] Tile_X3Y1_LUT4AB/EE4END[8] Tile_X3Y1_LUT4AB/EE4END[9]
+ Tile_X3Y1_LUT4AB/FrameData[0] Tile_X3Y1_LUT4AB/FrameData[10] Tile_X3Y1_LUT4AB/FrameData[11]
+ Tile_X3Y1_LUT4AB/FrameData[12] Tile_X3Y1_LUT4AB/FrameData[13] Tile_X3Y1_LUT4AB/FrameData[14]
+ Tile_X3Y1_LUT4AB/FrameData[15] Tile_X3Y1_LUT4AB/FrameData[16] Tile_X3Y1_LUT4AB/FrameData[17]
+ Tile_X3Y1_LUT4AB/FrameData[18] Tile_X3Y1_LUT4AB/FrameData[19] Tile_X3Y1_LUT4AB/FrameData[1]
+ Tile_X3Y1_LUT4AB/FrameData[20] Tile_X3Y1_LUT4AB/FrameData[21] Tile_X3Y1_LUT4AB/FrameData[22]
+ Tile_X3Y1_LUT4AB/FrameData[23] Tile_X3Y1_LUT4AB/FrameData[24] Tile_X3Y1_LUT4AB/FrameData[25]
+ Tile_X3Y1_LUT4AB/FrameData[26] Tile_X3Y1_LUT4AB/FrameData[27] Tile_X3Y1_LUT4AB/FrameData[28]
+ Tile_X3Y1_LUT4AB/FrameData[29] Tile_X3Y1_LUT4AB/FrameData[2] Tile_X3Y1_LUT4AB/FrameData[30]
+ Tile_X3Y1_LUT4AB/FrameData[31] Tile_X3Y1_LUT4AB/FrameData[3] Tile_X3Y1_LUT4AB/FrameData[4]
+ Tile_X3Y1_LUT4AB/FrameData[5] Tile_X3Y1_LUT4AB/FrameData[6] Tile_X3Y1_LUT4AB/FrameData[7]
+ Tile_X3Y1_LUT4AB/FrameData[8] Tile_X3Y1_LUT4AB/FrameData[9] Tile_X4Y1_LUT4AB/FrameData[0]
+ Tile_X4Y1_LUT4AB/FrameData[10] Tile_X4Y1_LUT4AB/FrameData[11] Tile_X4Y1_LUT4AB/FrameData[12]
+ Tile_X4Y1_LUT4AB/FrameData[13] Tile_X4Y1_LUT4AB/FrameData[14] Tile_X4Y1_LUT4AB/FrameData[15]
+ Tile_X4Y1_LUT4AB/FrameData[16] Tile_X4Y1_LUT4AB/FrameData[17] Tile_X4Y1_LUT4AB/FrameData[18]
+ Tile_X4Y1_LUT4AB/FrameData[19] Tile_X4Y1_LUT4AB/FrameData[1] Tile_X4Y1_LUT4AB/FrameData[20]
+ Tile_X4Y1_LUT4AB/FrameData[21] Tile_X4Y1_LUT4AB/FrameData[22] Tile_X4Y1_LUT4AB/FrameData[23]
+ Tile_X4Y1_LUT4AB/FrameData[24] Tile_X4Y1_LUT4AB/FrameData[25] Tile_X4Y1_LUT4AB/FrameData[26]
+ Tile_X4Y1_LUT4AB/FrameData[27] Tile_X4Y1_LUT4AB/FrameData[28] Tile_X4Y1_LUT4AB/FrameData[29]
+ Tile_X4Y1_LUT4AB/FrameData[2] Tile_X4Y1_LUT4AB/FrameData[30] Tile_X4Y1_LUT4AB/FrameData[31]
+ Tile_X4Y1_LUT4AB/FrameData[3] Tile_X4Y1_LUT4AB/FrameData[4] Tile_X4Y1_LUT4AB/FrameData[5]
+ Tile_X4Y1_LUT4AB/FrameData[6] Tile_X4Y1_LUT4AB/FrameData[7] Tile_X4Y1_LUT4AB/FrameData[8]
+ Tile_X4Y1_LUT4AB/FrameData[9] Tile_X3Y1_LUT4AB/FrameStrobe[0] Tile_X3Y1_LUT4AB/FrameStrobe[10]
+ Tile_X3Y1_LUT4AB/FrameStrobe[11] Tile_X3Y1_LUT4AB/FrameStrobe[12] Tile_X3Y1_LUT4AB/FrameStrobe[13]
+ Tile_X3Y1_LUT4AB/FrameStrobe[14] Tile_X3Y1_LUT4AB/FrameStrobe[15] Tile_X3Y1_LUT4AB/FrameStrobe[16]
+ Tile_X3Y1_LUT4AB/FrameStrobe[17] Tile_X3Y1_LUT4AB/FrameStrobe[18] Tile_X3Y1_LUT4AB/FrameStrobe[19]
+ Tile_X3Y1_LUT4AB/FrameStrobe[1] Tile_X3Y1_LUT4AB/FrameStrobe[2] Tile_X3Y1_LUT4AB/FrameStrobe[3]
+ Tile_X3Y1_LUT4AB/FrameStrobe[4] Tile_X3Y1_LUT4AB/FrameStrobe[5] Tile_X3Y1_LUT4AB/FrameStrobe[6]
+ Tile_X3Y1_LUT4AB/FrameStrobe[7] Tile_X3Y1_LUT4AB/FrameStrobe[8] Tile_X3Y1_LUT4AB/FrameStrobe[9]
+ Tile_X3Y0_N_IO4/FrameStrobe[0] Tile_X3Y0_N_IO4/FrameStrobe[10] Tile_X3Y0_N_IO4/FrameStrobe[11]
+ Tile_X3Y0_N_IO4/FrameStrobe[12] Tile_X3Y0_N_IO4/FrameStrobe[13] Tile_X3Y0_N_IO4/FrameStrobe[14]
+ Tile_X3Y0_N_IO4/FrameStrobe[15] Tile_X3Y0_N_IO4/FrameStrobe[16] Tile_X3Y0_N_IO4/FrameStrobe[17]
+ Tile_X3Y0_N_IO4/FrameStrobe[18] Tile_X3Y0_N_IO4/FrameStrobe[19] Tile_X3Y0_N_IO4/FrameStrobe[1]
+ Tile_X3Y0_N_IO4/FrameStrobe[2] Tile_X3Y0_N_IO4/FrameStrobe[3] Tile_X3Y0_N_IO4/FrameStrobe[4]
+ Tile_X3Y0_N_IO4/FrameStrobe[5] Tile_X3Y0_N_IO4/FrameStrobe[6] Tile_X3Y0_N_IO4/FrameStrobe[7]
+ Tile_X3Y0_N_IO4/FrameStrobe[8] Tile_X3Y0_N_IO4/FrameStrobe[9] Tile_X3Y0_N_IO4/N1END[0]
+ Tile_X3Y0_N_IO4/N1END[1] Tile_X3Y0_N_IO4/N1END[2] Tile_X3Y0_N_IO4/N1END[3] Tile_X3Y2_LUT4AB/N1BEG[0]
+ Tile_X3Y2_LUT4AB/N1BEG[1] Tile_X3Y2_LUT4AB/N1BEG[2] Tile_X3Y2_LUT4AB/N1BEG[3] Tile_X3Y0_N_IO4/N2MID[0]
+ Tile_X3Y0_N_IO4/N2MID[1] Tile_X3Y0_N_IO4/N2MID[2] Tile_X3Y0_N_IO4/N2MID[3] Tile_X3Y0_N_IO4/N2MID[4]
+ Tile_X3Y0_N_IO4/N2MID[5] Tile_X3Y0_N_IO4/N2MID[6] Tile_X3Y0_N_IO4/N2MID[7] Tile_X3Y0_N_IO4/N2END[0]
+ Tile_X3Y0_N_IO4/N2END[1] Tile_X3Y0_N_IO4/N2END[2] Tile_X3Y0_N_IO4/N2END[3] Tile_X3Y0_N_IO4/N2END[4]
+ Tile_X3Y0_N_IO4/N2END[5] Tile_X3Y0_N_IO4/N2END[6] Tile_X3Y0_N_IO4/N2END[7] Tile_X3Y1_LUT4AB/N2END[0]
+ Tile_X3Y1_LUT4AB/N2END[1] Tile_X3Y1_LUT4AB/N2END[2] Tile_X3Y1_LUT4AB/N2END[3] Tile_X3Y1_LUT4AB/N2END[4]
+ Tile_X3Y1_LUT4AB/N2END[5] Tile_X3Y1_LUT4AB/N2END[6] Tile_X3Y1_LUT4AB/N2END[7] Tile_X3Y2_LUT4AB/N2BEG[0]
+ Tile_X3Y2_LUT4AB/N2BEG[1] Tile_X3Y2_LUT4AB/N2BEG[2] Tile_X3Y2_LUT4AB/N2BEG[3] Tile_X3Y2_LUT4AB/N2BEG[4]
+ Tile_X3Y2_LUT4AB/N2BEG[5] Tile_X3Y2_LUT4AB/N2BEG[6] Tile_X3Y2_LUT4AB/N2BEG[7] Tile_X3Y0_N_IO4/N4END[0]
+ Tile_X3Y0_N_IO4/N4END[10] Tile_X3Y0_N_IO4/N4END[11] Tile_X3Y0_N_IO4/N4END[12] Tile_X3Y0_N_IO4/N4END[13]
+ Tile_X3Y0_N_IO4/N4END[14] Tile_X3Y0_N_IO4/N4END[15] Tile_X3Y0_N_IO4/N4END[1] Tile_X3Y0_N_IO4/N4END[2]
+ Tile_X3Y0_N_IO4/N4END[3] Tile_X3Y0_N_IO4/N4END[4] Tile_X3Y0_N_IO4/N4END[5] Tile_X3Y0_N_IO4/N4END[6]
+ Tile_X3Y0_N_IO4/N4END[7] Tile_X3Y0_N_IO4/N4END[8] Tile_X3Y0_N_IO4/N4END[9] Tile_X3Y2_LUT4AB/N4BEG[0]
+ Tile_X3Y2_LUT4AB/N4BEG[10] Tile_X3Y2_LUT4AB/N4BEG[11] Tile_X3Y2_LUT4AB/N4BEG[12]
+ Tile_X3Y2_LUT4AB/N4BEG[13] Tile_X3Y2_LUT4AB/N4BEG[14] Tile_X3Y2_LUT4AB/N4BEG[15]
+ Tile_X3Y2_LUT4AB/N4BEG[1] Tile_X3Y2_LUT4AB/N4BEG[2] Tile_X3Y2_LUT4AB/N4BEG[3] Tile_X3Y2_LUT4AB/N4BEG[4]
+ Tile_X3Y2_LUT4AB/N4BEG[5] Tile_X3Y2_LUT4AB/N4BEG[6] Tile_X3Y2_LUT4AB/N4BEG[7] Tile_X3Y2_LUT4AB/N4BEG[8]
+ Tile_X3Y2_LUT4AB/N4BEG[9] Tile_X3Y0_N_IO4/NN4END[0] Tile_X3Y0_N_IO4/NN4END[10] Tile_X3Y0_N_IO4/NN4END[11]
+ Tile_X3Y0_N_IO4/NN4END[12] Tile_X3Y0_N_IO4/NN4END[13] Tile_X3Y0_N_IO4/NN4END[14]
+ Tile_X3Y0_N_IO4/NN4END[15] Tile_X3Y0_N_IO4/NN4END[1] Tile_X3Y0_N_IO4/NN4END[2] Tile_X3Y0_N_IO4/NN4END[3]
+ Tile_X3Y0_N_IO4/NN4END[4] Tile_X3Y0_N_IO4/NN4END[5] Tile_X3Y0_N_IO4/NN4END[6] Tile_X3Y0_N_IO4/NN4END[7]
+ Tile_X3Y0_N_IO4/NN4END[8] Tile_X3Y0_N_IO4/NN4END[9] Tile_X3Y2_LUT4AB/NN4BEG[0] Tile_X3Y2_LUT4AB/NN4BEG[10]
+ Tile_X3Y2_LUT4AB/NN4BEG[11] Tile_X3Y2_LUT4AB/NN4BEG[12] Tile_X3Y2_LUT4AB/NN4BEG[13]
+ Tile_X3Y2_LUT4AB/NN4BEG[14] Tile_X3Y2_LUT4AB/NN4BEG[15] Tile_X3Y2_LUT4AB/NN4BEG[1]
+ Tile_X3Y2_LUT4AB/NN4BEG[2] Tile_X3Y2_LUT4AB/NN4BEG[3] Tile_X3Y2_LUT4AB/NN4BEG[4]
+ Tile_X3Y2_LUT4AB/NN4BEG[5] Tile_X3Y2_LUT4AB/NN4BEG[6] Tile_X3Y2_LUT4AB/NN4BEG[7]
+ Tile_X3Y2_LUT4AB/NN4BEG[8] Tile_X3Y2_LUT4AB/NN4BEG[9] Tile_X3Y2_LUT4AB/S1END[0]
+ Tile_X3Y2_LUT4AB/S1END[1] Tile_X3Y2_LUT4AB/S1END[2] Tile_X3Y2_LUT4AB/S1END[3] Tile_X3Y0_N_IO4/S1BEG[0]
+ Tile_X3Y0_N_IO4/S1BEG[1] Tile_X3Y0_N_IO4/S1BEG[2] Tile_X3Y0_N_IO4/S1BEG[3] Tile_X3Y2_LUT4AB/S2MID[0]
+ Tile_X3Y2_LUT4AB/S2MID[1] Tile_X3Y2_LUT4AB/S2MID[2] Tile_X3Y2_LUT4AB/S2MID[3] Tile_X3Y2_LUT4AB/S2MID[4]
+ Tile_X3Y2_LUT4AB/S2MID[5] Tile_X3Y2_LUT4AB/S2MID[6] Tile_X3Y2_LUT4AB/S2MID[7] Tile_X3Y2_LUT4AB/S2END[0]
+ Tile_X3Y2_LUT4AB/S2END[1] Tile_X3Y2_LUT4AB/S2END[2] Tile_X3Y2_LUT4AB/S2END[3] Tile_X3Y2_LUT4AB/S2END[4]
+ Tile_X3Y2_LUT4AB/S2END[5] Tile_X3Y2_LUT4AB/S2END[6] Tile_X3Y2_LUT4AB/S2END[7] Tile_X3Y1_LUT4AB/S2END[0]
+ Tile_X3Y1_LUT4AB/S2END[1] Tile_X3Y1_LUT4AB/S2END[2] Tile_X3Y1_LUT4AB/S2END[3] Tile_X3Y1_LUT4AB/S2END[4]
+ Tile_X3Y1_LUT4AB/S2END[5] Tile_X3Y1_LUT4AB/S2END[6] Tile_X3Y1_LUT4AB/S2END[7] Tile_X3Y0_N_IO4/S2BEG[0]
+ Tile_X3Y0_N_IO4/S2BEG[1] Tile_X3Y0_N_IO4/S2BEG[2] Tile_X3Y0_N_IO4/S2BEG[3] Tile_X3Y0_N_IO4/S2BEG[4]
+ Tile_X3Y0_N_IO4/S2BEG[5] Tile_X3Y0_N_IO4/S2BEG[6] Tile_X3Y0_N_IO4/S2BEG[7] Tile_X3Y2_LUT4AB/S4END[0]
+ Tile_X3Y2_LUT4AB/S4END[10] Tile_X3Y2_LUT4AB/S4END[11] Tile_X3Y2_LUT4AB/S4END[12]
+ Tile_X3Y2_LUT4AB/S4END[13] Tile_X3Y2_LUT4AB/S4END[14] Tile_X3Y2_LUT4AB/S4END[15]
+ Tile_X3Y2_LUT4AB/S4END[1] Tile_X3Y2_LUT4AB/S4END[2] Tile_X3Y2_LUT4AB/S4END[3] Tile_X3Y2_LUT4AB/S4END[4]
+ Tile_X3Y2_LUT4AB/S4END[5] Tile_X3Y2_LUT4AB/S4END[6] Tile_X3Y2_LUT4AB/S4END[7] Tile_X3Y2_LUT4AB/S4END[8]
+ Tile_X3Y2_LUT4AB/S4END[9] Tile_X3Y0_N_IO4/S4BEG[0] Tile_X3Y0_N_IO4/S4BEG[10] Tile_X3Y0_N_IO4/S4BEG[11]
+ Tile_X3Y0_N_IO4/S4BEG[12] Tile_X3Y0_N_IO4/S4BEG[13] Tile_X3Y0_N_IO4/S4BEG[14] Tile_X3Y0_N_IO4/S4BEG[15]
+ Tile_X3Y0_N_IO4/S4BEG[1] Tile_X3Y0_N_IO4/S4BEG[2] Tile_X3Y0_N_IO4/S4BEG[3] Tile_X3Y0_N_IO4/S4BEG[4]
+ Tile_X3Y0_N_IO4/S4BEG[5] Tile_X3Y0_N_IO4/S4BEG[6] Tile_X3Y0_N_IO4/S4BEG[7] Tile_X3Y0_N_IO4/S4BEG[8]
+ Tile_X3Y0_N_IO4/S4BEG[9] Tile_X3Y2_LUT4AB/SS4END[0] Tile_X3Y2_LUT4AB/SS4END[10]
+ Tile_X3Y2_LUT4AB/SS4END[11] Tile_X3Y2_LUT4AB/SS4END[12] Tile_X3Y2_LUT4AB/SS4END[13]
+ Tile_X3Y2_LUT4AB/SS4END[14] Tile_X3Y2_LUT4AB/SS4END[15] Tile_X3Y2_LUT4AB/SS4END[1]
+ Tile_X3Y2_LUT4AB/SS4END[2] Tile_X3Y2_LUT4AB/SS4END[3] Tile_X3Y2_LUT4AB/SS4END[4]
+ Tile_X3Y2_LUT4AB/SS4END[5] Tile_X3Y2_LUT4AB/SS4END[6] Tile_X3Y2_LUT4AB/SS4END[7]
+ Tile_X3Y2_LUT4AB/SS4END[8] Tile_X3Y2_LUT4AB/SS4END[9] Tile_X3Y0_N_IO4/SS4BEG[0]
+ Tile_X3Y0_N_IO4/SS4BEG[10] Tile_X3Y0_N_IO4/SS4BEG[11] Tile_X3Y0_N_IO4/SS4BEG[12]
+ Tile_X3Y0_N_IO4/SS4BEG[13] Tile_X3Y0_N_IO4/SS4BEG[14] Tile_X3Y0_N_IO4/SS4BEG[15]
+ Tile_X3Y0_N_IO4/SS4BEG[1] Tile_X3Y0_N_IO4/SS4BEG[2] Tile_X3Y0_N_IO4/SS4BEG[3] Tile_X3Y0_N_IO4/SS4BEG[4]
+ Tile_X3Y0_N_IO4/SS4BEG[5] Tile_X3Y0_N_IO4/SS4BEG[6] Tile_X3Y0_N_IO4/SS4BEG[7] Tile_X3Y0_N_IO4/SS4BEG[8]
+ Tile_X3Y0_N_IO4/SS4BEG[9] Tile_X3Y1_LUT4AB/UserCLK Tile_X3Y0_N_IO4/UserCLK VGND
+ VPWR Tile_X3Y1_LUT4AB/W1BEG[0] Tile_X3Y1_LUT4AB/W1BEG[1] Tile_X3Y1_LUT4AB/W1BEG[2]
+ Tile_X3Y1_LUT4AB/W1BEG[3] Tile_X4Y1_LUT4AB/W1BEG[0] Tile_X4Y1_LUT4AB/W1BEG[1] Tile_X4Y1_LUT4AB/W1BEG[2]
+ Tile_X4Y1_LUT4AB/W1BEG[3] Tile_X3Y1_LUT4AB/W2BEG[0] Tile_X3Y1_LUT4AB/W2BEG[1] Tile_X3Y1_LUT4AB/W2BEG[2]
+ Tile_X3Y1_LUT4AB/W2BEG[3] Tile_X3Y1_LUT4AB/W2BEG[4] Tile_X3Y1_LUT4AB/W2BEG[5] Tile_X3Y1_LUT4AB/W2BEG[6]
+ Tile_X3Y1_LUT4AB/W2BEG[7] Tile_X2Y1_LUT4AB/W2END[0] Tile_X2Y1_LUT4AB/W2END[1] Tile_X2Y1_LUT4AB/W2END[2]
+ Tile_X2Y1_LUT4AB/W2END[3] Tile_X2Y1_LUT4AB/W2END[4] Tile_X2Y1_LUT4AB/W2END[5] Tile_X2Y1_LUT4AB/W2END[6]
+ Tile_X2Y1_LUT4AB/W2END[7] Tile_X3Y1_LUT4AB/W2END[0] Tile_X3Y1_LUT4AB/W2END[1] Tile_X3Y1_LUT4AB/W2END[2]
+ Tile_X3Y1_LUT4AB/W2END[3] Tile_X3Y1_LUT4AB/W2END[4] Tile_X3Y1_LUT4AB/W2END[5] Tile_X3Y1_LUT4AB/W2END[6]
+ Tile_X3Y1_LUT4AB/W2END[7] Tile_X4Y1_LUT4AB/W2BEG[0] Tile_X4Y1_LUT4AB/W2BEG[1] Tile_X4Y1_LUT4AB/W2BEG[2]
+ Tile_X4Y1_LUT4AB/W2BEG[3] Tile_X4Y1_LUT4AB/W2BEG[4] Tile_X4Y1_LUT4AB/W2BEG[5] Tile_X4Y1_LUT4AB/W2BEG[6]
+ Tile_X4Y1_LUT4AB/W2BEG[7] Tile_X3Y1_LUT4AB/W6BEG[0] Tile_X3Y1_LUT4AB/W6BEG[10] Tile_X3Y1_LUT4AB/W6BEG[11]
+ Tile_X3Y1_LUT4AB/W6BEG[1] Tile_X3Y1_LUT4AB/W6BEG[2] Tile_X3Y1_LUT4AB/W6BEG[3] Tile_X3Y1_LUT4AB/W6BEG[4]
+ Tile_X3Y1_LUT4AB/W6BEG[5] Tile_X3Y1_LUT4AB/W6BEG[6] Tile_X3Y1_LUT4AB/W6BEG[7] Tile_X3Y1_LUT4AB/W6BEG[8]
+ Tile_X3Y1_LUT4AB/W6BEG[9] Tile_X4Y1_LUT4AB/W6BEG[0] Tile_X4Y1_LUT4AB/W6BEG[10] Tile_X4Y1_LUT4AB/W6BEG[11]
+ Tile_X4Y1_LUT4AB/W6BEG[1] Tile_X4Y1_LUT4AB/W6BEG[2] Tile_X4Y1_LUT4AB/W6BEG[3] Tile_X4Y1_LUT4AB/W6BEG[4]
+ Tile_X4Y1_LUT4AB/W6BEG[5] Tile_X4Y1_LUT4AB/W6BEG[6] Tile_X4Y1_LUT4AB/W6BEG[7] Tile_X4Y1_LUT4AB/W6BEG[8]
+ Tile_X4Y1_LUT4AB/W6BEG[9] Tile_X3Y1_LUT4AB/WW4BEG[0] Tile_X3Y1_LUT4AB/WW4BEG[10]
+ Tile_X3Y1_LUT4AB/WW4BEG[11] Tile_X3Y1_LUT4AB/WW4BEG[12] Tile_X3Y1_LUT4AB/WW4BEG[13]
+ Tile_X3Y1_LUT4AB/WW4BEG[14] Tile_X3Y1_LUT4AB/WW4BEG[15] Tile_X3Y1_LUT4AB/WW4BEG[1]
+ Tile_X3Y1_LUT4AB/WW4BEG[2] Tile_X3Y1_LUT4AB/WW4BEG[3] Tile_X3Y1_LUT4AB/WW4BEG[4]
+ Tile_X3Y1_LUT4AB/WW4BEG[5] Tile_X3Y1_LUT4AB/WW4BEG[6] Tile_X3Y1_LUT4AB/WW4BEG[7]
+ Tile_X3Y1_LUT4AB/WW4BEG[8] Tile_X3Y1_LUT4AB/WW4BEG[9] Tile_X4Y1_LUT4AB/WW4BEG[0]
+ Tile_X4Y1_LUT4AB/WW4BEG[10] Tile_X4Y1_LUT4AB/WW4BEG[11] Tile_X4Y1_LUT4AB/WW4BEG[12]
+ Tile_X4Y1_LUT4AB/WW4BEG[13] Tile_X4Y1_LUT4AB/WW4BEG[14] Tile_X4Y1_LUT4AB/WW4BEG[15]
+ Tile_X4Y1_LUT4AB/WW4BEG[1] Tile_X4Y1_LUT4AB/WW4BEG[2] Tile_X4Y1_LUT4AB/WW4BEG[3]
+ Tile_X4Y1_LUT4AB/WW4BEG[4] Tile_X4Y1_LUT4AB/WW4BEG[5] Tile_X4Y1_LUT4AB/WW4BEG[6]
+ Tile_X4Y1_LUT4AB/WW4BEG[7] Tile_X4Y1_LUT4AB/WW4BEG[8] Tile_X4Y1_LUT4AB/WW4BEG[9]
+ LUT4AB
XTile_X2Y5_LUT4AB Tile_X2Y6_LUT4AB/Co Tile_X2Y5_LUT4AB/Co Tile_X3Y5_LUT4AB/E1END[0]
+ Tile_X3Y5_LUT4AB/E1END[1] Tile_X3Y5_LUT4AB/E1END[2] Tile_X3Y5_LUT4AB/E1END[3] Tile_X2Y5_LUT4AB/E1END[0]
+ Tile_X2Y5_LUT4AB/E1END[1] Tile_X2Y5_LUT4AB/E1END[2] Tile_X2Y5_LUT4AB/E1END[3] Tile_X3Y5_LUT4AB/E2MID[0]
+ Tile_X3Y5_LUT4AB/E2MID[1] Tile_X3Y5_LUT4AB/E2MID[2] Tile_X3Y5_LUT4AB/E2MID[3] Tile_X3Y5_LUT4AB/E2MID[4]
+ Tile_X3Y5_LUT4AB/E2MID[5] Tile_X3Y5_LUT4AB/E2MID[6] Tile_X3Y5_LUT4AB/E2MID[7] Tile_X3Y5_LUT4AB/E2END[0]
+ Tile_X3Y5_LUT4AB/E2END[1] Tile_X3Y5_LUT4AB/E2END[2] Tile_X3Y5_LUT4AB/E2END[3] Tile_X3Y5_LUT4AB/E2END[4]
+ Tile_X3Y5_LUT4AB/E2END[5] Tile_X3Y5_LUT4AB/E2END[6] Tile_X3Y5_LUT4AB/E2END[7] Tile_X2Y5_LUT4AB/E2END[0]
+ Tile_X2Y5_LUT4AB/E2END[1] Tile_X2Y5_LUT4AB/E2END[2] Tile_X2Y5_LUT4AB/E2END[3] Tile_X2Y5_LUT4AB/E2END[4]
+ Tile_X2Y5_LUT4AB/E2END[5] Tile_X2Y5_LUT4AB/E2END[6] Tile_X2Y5_LUT4AB/E2END[7] Tile_X2Y5_LUT4AB/E2MID[0]
+ Tile_X2Y5_LUT4AB/E2MID[1] Tile_X2Y5_LUT4AB/E2MID[2] Tile_X2Y5_LUT4AB/E2MID[3] Tile_X2Y5_LUT4AB/E2MID[4]
+ Tile_X2Y5_LUT4AB/E2MID[5] Tile_X2Y5_LUT4AB/E2MID[6] Tile_X2Y5_LUT4AB/E2MID[7] Tile_X3Y5_LUT4AB/E6END[0]
+ Tile_X3Y5_LUT4AB/E6END[10] Tile_X3Y5_LUT4AB/E6END[11] Tile_X3Y5_LUT4AB/E6END[1]
+ Tile_X3Y5_LUT4AB/E6END[2] Tile_X3Y5_LUT4AB/E6END[3] Tile_X3Y5_LUT4AB/E6END[4] Tile_X3Y5_LUT4AB/E6END[5]
+ Tile_X3Y5_LUT4AB/E6END[6] Tile_X3Y5_LUT4AB/E6END[7] Tile_X3Y5_LUT4AB/E6END[8] Tile_X3Y5_LUT4AB/E6END[9]
+ Tile_X2Y5_LUT4AB/E6END[0] Tile_X2Y5_LUT4AB/E6END[10] Tile_X2Y5_LUT4AB/E6END[11]
+ Tile_X2Y5_LUT4AB/E6END[1] Tile_X2Y5_LUT4AB/E6END[2] Tile_X2Y5_LUT4AB/E6END[3] Tile_X2Y5_LUT4AB/E6END[4]
+ Tile_X2Y5_LUT4AB/E6END[5] Tile_X2Y5_LUT4AB/E6END[6] Tile_X2Y5_LUT4AB/E6END[7] Tile_X2Y5_LUT4AB/E6END[8]
+ Tile_X2Y5_LUT4AB/E6END[9] Tile_X3Y5_LUT4AB/EE4END[0] Tile_X3Y5_LUT4AB/EE4END[10]
+ Tile_X3Y5_LUT4AB/EE4END[11] Tile_X3Y5_LUT4AB/EE4END[12] Tile_X3Y5_LUT4AB/EE4END[13]
+ Tile_X3Y5_LUT4AB/EE4END[14] Tile_X3Y5_LUT4AB/EE4END[15] Tile_X3Y5_LUT4AB/EE4END[1]
+ Tile_X3Y5_LUT4AB/EE4END[2] Tile_X3Y5_LUT4AB/EE4END[3] Tile_X3Y5_LUT4AB/EE4END[4]
+ Tile_X3Y5_LUT4AB/EE4END[5] Tile_X3Y5_LUT4AB/EE4END[6] Tile_X3Y5_LUT4AB/EE4END[7]
+ Tile_X3Y5_LUT4AB/EE4END[8] Tile_X3Y5_LUT4AB/EE4END[9] Tile_X2Y5_LUT4AB/EE4END[0]
+ Tile_X2Y5_LUT4AB/EE4END[10] Tile_X2Y5_LUT4AB/EE4END[11] Tile_X2Y5_LUT4AB/EE4END[12]
+ Tile_X2Y5_LUT4AB/EE4END[13] Tile_X2Y5_LUT4AB/EE4END[14] Tile_X2Y5_LUT4AB/EE4END[15]
+ Tile_X2Y5_LUT4AB/EE4END[1] Tile_X2Y5_LUT4AB/EE4END[2] Tile_X2Y5_LUT4AB/EE4END[3]
+ Tile_X2Y5_LUT4AB/EE4END[4] Tile_X2Y5_LUT4AB/EE4END[5] Tile_X2Y5_LUT4AB/EE4END[6]
+ Tile_X2Y5_LUT4AB/EE4END[7] Tile_X2Y5_LUT4AB/EE4END[8] Tile_X2Y5_LUT4AB/EE4END[9]
+ Tile_X2Y5_LUT4AB/FrameData[0] Tile_X2Y5_LUT4AB/FrameData[10] Tile_X2Y5_LUT4AB/FrameData[11]
+ Tile_X2Y5_LUT4AB/FrameData[12] Tile_X2Y5_LUT4AB/FrameData[13] Tile_X2Y5_LUT4AB/FrameData[14]
+ Tile_X2Y5_LUT4AB/FrameData[15] Tile_X2Y5_LUT4AB/FrameData[16] Tile_X2Y5_LUT4AB/FrameData[17]
+ Tile_X2Y5_LUT4AB/FrameData[18] Tile_X2Y5_LUT4AB/FrameData[19] Tile_X2Y5_LUT4AB/FrameData[1]
+ Tile_X2Y5_LUT4AB/FrameData[20] Tile_X2Y5_LUT4AB/FrameData[21] Tile_X2Y5_LUT4AB/FrameData[22]
+ Tile_X2Y5_LUT4AB/FrameData[23] Tile_X2Y5_LUT4AB/FrameData[24] Tile_X2Y5_LUT4AB/FrameData[25]
+ Tile_X2Y5_LUT4AB/FrameData[26] Tile_X2Y5_LUT4AB/FrameData[27] Tile_X2Y5_LUT4AB/FrameData[28]
+ Tile_X2Y5_LUT4AB/FrameData[29] Tile_X2Y5_LUT4AB/FrameData[2] Tile_X2Y5_LUT4AB/FrameData[30]
+ Tile_X2Y5_LUT4AB/FrameData[31] Tile_X2Y5_LUT4AB/FrameData[3] Tile_X2Y5_LUT4AB/FrameData[4]
+ Tile_X2Y5_LUT4AB/FrameData[5] Tile_X2Y5_LUT4AB/FrameData[6] Tile_X2Y5_LUT4AB/FrameData[7]
+ Tile_X2Y5_LUT4AB/FrameData[8] Tile_X2Y5_LUT4AB/FrameData[9] Tile_X3Y5_LUT4AB/FrameData[0]
+ Tile_X3Y5_LUT4AB/FrameData[10] Tile_X3Y5_LUT4AB/FrameData[11] Tile_X3Y5_LUT4AB/FrameData[12]
+ Tile_X3Y5_LUT4AB/FrameData[13] Tile_X3Y5_LUT4AB/FrameData[14] Tile_X3Y5_LUT4AB/FrameData[15]
+ Tile_X3Y5_LUT4AB/FrameData[16] Tile_X3Y5_LUT4AB/FrameData[17] Tile_X3Y5_LUT4AB/FrameData[18]
+ Tile_X3Y5_LUT4AB/FrameData[19] Tile_X3Y5_LUT4AB/FrameData[1] Tile_X3Y5_LUT4AB/FrameData[20]
+ Tile_X3Y5_LUT4AB/FrameData[21] Tile_X3Y5_LUT4AB/FrameData[22] Tile_X3Y5_LUT4AB/FrameData[23]
+ Tile_X3Y5_LUT4AB/FrameData[24] Tile_X3Y5_LUT4AB/FrameData[25] Tile_X3Y5_LUT4AB/FrameData[26]
+ Tile_X3Y5_LUT4AB/FrameData[27] Tile_X3Y5_LUT4AB/FrameData[28] Tile_X3Y5_LUT4AB/FrameData[29]
+ Tile_X3Y5_LUT4AB/FrameData[2] Tile_X3Y5_LUT4AB/FrameData[30] Tile_X3Y5_LUT4AB/FrameData[31]
+ Tile_X3Y5_LUT4AB/FrameData[3] Tile_X3Y5_LUT4AB/FrameData[4] Tile_X3Y5_LUT4AB/FrameData[5]
+ Tile_X3Y5_LUT4AB/FrameData[6] Tile_X3Y5_LUT4AB/FrameData[7] Tile_X3Y5_LUT4AB/FrameData[8]
+ Tile_X3Y5_LUT4AB/FrameData[9] Tile_X2Y5_LUT4AB/FrameStrobe[0] Tile_X2Y5_LUT4AB/FrameStrobe[10]
+ Tile_X2Y5_LUT4AB/FrameStrobe[11] Tile_X2Y5_LUT4AB/FrameStrobe[12] Tile_X2Y5_LUT4AB/FrameStrobe[13]
+ Tile_X2Y5_LUT4AB/FrameStrobe[14] Tile_X2Y5_LUT4AB/FrameStrobe[15] Tile_X2Y5_LUT4AB/FrameStrobe[16]
+ Tile_X2Y5_LUT4AB/FrameStrobe[17] Tile_X2Y5_LUT4AB/FrameStrobe[18] Tile_X2Y5_LUT4AB/FrameStrobe[19]
+ Tile_X2Y5_LUT4AB/FrameStrobe[1] Tile_X2Y5_LUT4AB/FrameStrobe[2] Tile_X2Y5_LUT4AB/FrameStrobe[3]
+ Tile_X2Y5_LUT4AB/FrameStrobe[4] Tile_X2Y5_LUT4AB/FrameStrobe[5] Tile_X2Y5_LUT4AB/FrameStrobe[6]
+ Tile_X2Y5_LUT4AB/FrameStrobe[7] Tile_X2Y5_LUT4AB/FrameStrobe[8] Tile_X2Y5_LUT4AB/FrameStrobe[9]
+ Tile_X2Y4_LUT4AB/FrameStrobe[0] Tile_X2Y4_LUT4AB/FrameStrobe[10] Tile_X2Y4_LUT4AB/FrameStrobe[11]
+ Tile_X2Y4_LUT4AB/FrameStrobe[12] Tile_X2Y4_LUT4AB/FrameStrobe[13] Tile_X2Y4_LUT4AB/FrameStrobe[14]
+ Tile_X2Y4_LUT4AB/FrameStrobe[15] Tile_X2Y4_LUT4AB/FrameStrobe[16] Tile_X2Y4_LUT4AB/FrameStrobe[17]
+ Tile_X2Y4_LUT4AB/FrameStrobe[18] Tile_X2Y4_LUT4AB/FrameStrobe[19] Tile_X2Y4_LUT4AB/FrameStrobe[1]
+ Tile_X2Y4_LUT4AB/FrameStrobe[2] Tile_X2Y4_LUT4AB/FrameStrobe[3] Tile_X2Y4_LUT4AB/FrameStrobe[4]
+ Tile_X2Y4_LUT4AB/FrameStrobe[5] Tile_X2Y4_LUT4AB/FrameStrobe[6] Tile_X2Y4_LUT4AB/FrameStrobe[7]
+ Tile_X2Y4_LUT4AB/FrameStrobe[8] Tile_X2Y4_LUT4AB/FrameStrobe[9] Tile_X2Y5_LUT4AB/N1BEG[0]
+ Tile_X2Y5_LUT4AB/N1BEG[1] Tile_X2Y5_LUT4AB/N1BEG[2] Tile_X2Y5_LUT4AB/N1BEG[3] Tile_X2Y6_LUT4AB/N1BEG[0]
+ Tile_X2Y6_LUT4AB/N1BEG[1] Tile_X2Y6_LUT4AB/N1BEG[2] Tile_X2Y6_LUT4AB/N1BEG[3] Tile_X2Y5_LUT4AB/N2BEG[0]
+ Tile_X2Y5_LUT4AB/N2BEG[1] Tile_X2Y5_LUT4AB/N2BEG[2] Tile_X2Y5_LUT4AB/N2BEG[3] Tile_X2Y5_LUT4AB/N2BEG[4]
+ Tile_X2Y5_LUT4AB/N2BEG[5] Tile_X2Y5_LUT4AB/N2BEG[6] Tile_X2Y5_LUT4AB/N2BEG[7] Tile_X2Y4_LUT4AB/N2END[0]
+ Tile_X2Y4_LUT4AB/N2END[1] Tile_X2Y4_LUT4AB/N2END[2] Tile_X2Y4_LUT4AB/N2END[3] Tile_X2Y4_LUT4AB/N2END[4]
+ Tile_X2Y4_LUT4AB/N2END[5] Tile_X2Y4_LUT4AB/N2END[6] Tile_X2Y4_LUT4AB/N2END[7] Tile_X2Y5_LUT4AB/N2END[0]
+ Tile_X2Y5_LUT4AB/N2END[1] Tile_X2Y5_LUT4AB/N2END[2] Tile_X2Y5_LUT4AB/N2END[3] Tile_X2Y5_LUT4AB/N2END[4]
+ Tile_X2Y5_LUT4AB/N2END[5] Tile_X2Y5_LUT4AB/N2END[6] Tile_X2Y5_LUT4AB/N2END[7] Tile_X2Y6_LUT4AB/N2BEG[0]
+ Tile_X2Y6_LUT4AB/N2BEG[1] Tile_X2Y6_LUT4AB/N2BEG[2] Tile_X2Y6_LUT4AB/N2BEG[3] Tile_X2Y6_LUT4AB/N2BEG[4]
+ Tile_X2Y6_LUT4AB/N2BEG[5] Tile_X2Y6_LUT4AB/N2BEG[6] Tile_X2Y6_LUT4AB/N2BEG[7] Tile_X2Y5_LUT4AB/N4BEG[0]
+ Tile_X2Y5_LUT4AB/N4BEG[10] Tile_X2Y5_LUT4AB/N4BEG[11] Tile_X2Y5_LUT4AB/N4BEG[12]
+ Tile_X2Y5_LUT4AB/N4BEG[13] Tile_X2Y5_LUT4AB/N4BEG[14] Tile_X2Y5_LUT4AB/N4BEG[15]
+ Tile_X2Y5_LUT4AB/N4BEG[1] Tile_X2Y5_LUT4AB/N4BEG[2] Tile_X2Y5_LUT4AB/N4BEG[3] Tile_X2Y5_LUT4AB/N4BEG[4]
+ Tile_X2Y5_LUT4AB/N4BEG[5] Tile_X2Y5_LUT4AB/N4BEG[6] Tile_X2Y5_LUT4AB/N4BEG[7] Tile_X2Y5_LUT4AB/N4BEG[8]
+ Tile_X2Y5_LUT4AB/N4BEG[9] Tile_X2Y6_LUT4AB/N4BEG[0] Tile_X2Y6_LUT4AB/N4BEG[10] Tile_X2Y6_LUT4AB/N4BEG[11]
+ Tile_X2Y6_LUT4AB/N4BEG[12] Tile_X2Y6_LUT4AB/N4BEG[13] Tile_X2Y6_LUT4AB/N4BEG[14]
+ Tile_X2Y6_LUT4AB/N4BEG[15] Tile_X2Y6_LUT4AB/N4BEG[1] Tile_X2Y6_LUT4AB/N4BEG[2] Tile_X2Y6_LUT4AB/N4BEG[3]
+ Tile_X2Y6_LUT4AB/N4BEG[4] Tile_X2Y6_LUT4AB/N4BEG[5] Tile_X2Y6_LUT4AB/N4BEG[6] Tile_X2Y6_LUT4AB/N4BEG[7]
+ Tile_X2Y6_LUT4AB/N4BEG[8] Tile_X2Y6_LUT4AB/N4BEG[9] Tile_X2Y5_LUT4AB/NN4BEG[0] Tile_X2Y5_LUT4AB/NN4BEG[10]
+ Tile_X2Y5_LUT4AB/NN4BEG[11] Tile_X2Y5_LUT4AB/NN4BEG[12] Tile_X2Y5_LUT4AB/NN4BEG[13]
+ Tile_X2Y5_LUT4AB/NN4BEG[14] Tile_X2Y5_LUT4AB/NN4BEG[15] Tile_X2Y5_LUT4AB/NN4BEG[1]
+ Tile_X2Y5_LUT4AB/NN4BEG[2] Tile_X2Y5_LUT4AB/NN4BEG[3] Tile_X2Y5_LUT4AB/NN4BEG[4]
+ Tile_X2Y5_LUT4AB/NN4BEG[5] Tile_X2Y5_LUT4AB/NN4BEG[6] Tile_X2Y5_LUT4AB/NN4BEG[7]
+ Tile_X2Y5_LUT4AB/NN4BEG[8] Tile_X2Y5_LUT4AB/NN4BEG[9] Tile_X2Y6_LUT4AB/NN4BEG[0]
+ Tile_X2Y6_LUT4AB/NN4BEG[10] Tile_X2Y6_LUT4AB/NN4BEG[11] Tile_X2Y6_LUT4AB/NN4BEG[12]
+ Tile_X2Y6_LUT4AB/NN4BEG[13] Tile_X2Y6_LUT4AB/NN4BEG[14] Tile_X2Y6_LUT4AB/NN4BEG[15]
+ Tile_X2Y6_LUT4AB/NN4BEG[1] Tile_X2Y6_LUT4AB/NN4BEG[2] Tile_X2Y6_LUT4AB/NN4BEG[3]
+ Tile_X2Y6_LUT4AB/NN4BEG[4] Tile_X2Y6_LUT4AB/NN4BEG[5] Tile_X2Y6_LUT4AB/NN4BEG[6]
+ Tile_X2Y6_LUT4AB/NN4BEG[7] Tile_X2Y6_LUT4AB/NN4BEG[8] Tile_X2Y6_LUT4AB/NN4BEG[9]
+ Tile_X2Y6_LUT4AB/S1END[0] Tile_X2Y6_LUT4AB/S1END[1] Tile_X2Y6_LUT4AB/S1END[2] Tile_X2Y6_LUT4AB/S1END[3]
+ Tile_X2Y5_LUT4AB/S1END[0] Tile_X2Y5_LUT4AB/S1END[1] Tile_X2Y5_LUT4AB/S1END[2] Tile_X2Y5_LUT4AB/S1END[3]
+ Tile_X2Y6_LUT4AB/S2MID[0] Tile_X2Y6_LUT4AB/S2MID[1] Tile_X2Y6_LUT4AB/S2MID[2] Tile_X2Y6_LUT4AB/S2MID[3]
+ Tile_X2Y6_LUT4AB/S2MID[4] Tile_X2Y6_LUT4AB/S2MID[5] Tile_X2Y6_LUT4AB/S2MID[6] Tile_X2Y6_LUT4AB/S2MID[7]
+ Tile_X2Y6_LUT4AB/S2END[0] Tile_X2Y6_LUT4AB/S2END[1] Tile_X2Y6_LUT4AB/S2END[2] Tile_X2Y6_LUT4AB/S2END[3]
+ Tile_X2Y6_LUT4AB/S2END[4] Tile_X2Y6_LUT4AB/S2END[5] Tile_X2Y6_LUT4AB/S2END[6] Tile_X2Y6_LUT4AB/S2END[7]
+ Tile_X2Y5_LUT4AB/S2END[0] Tile_X2Y5_LUT4AB/S2END[1] Tile_X2Y5_LUT4AB/S2END[2] Tile_X2Y5_LUT4AB/S2END[3]
+ Tile_X2Y5_LUT4AB/S2END[4] Tile_X2Y5_LUT4AB/S2END[5] Tile_X2Y5_LUT4AB/S2END[6] Tile_X2Y5_LUT4AB/S2END[7]
+ Tile_X2Y5_LUT4AB/S2MID[0] Tile_X2Y5_LUT4AB/S2MID[1] Tile_X2Y5_LUT4AB/S2MID[2] Tile_X2Y5_LUT4AB/S2MID[3]
+ Tile_X2Y5_LUT4AB/S2MID[4] Tile_X2Y5_LUT4AB/S2MID[5] Tile_X2Y5_LUT4AB/S2MID[6] Tile_X2Y5_LUT4AB/S2MID[7]
+ Tile_X2Y6_LUT4AB/S4END[0] Tile_X2Y6_LUT4AB/S4END[10] Tile_X2Y6_LUT4AB/S4END[11]
+ Tile_X2Y6_LUT4AB/S4END[12] Tile_X2Y6_LUT4AB/S4END[13] Tile_X2Y6_LUT4AB/S4END[14]
+ Tile_X2Y6_LUT4AB/S4END[15] Tile_X2Y6_LUT4AB/S4END[1] Tile_X2Y6_LUT4AB/S4END[2] Tile_X2Y6_LUT4AB/S4END[3]
+ Tile_X2Y6_LUT4AB/S4END[4] Tile_X2Y6_LUT4AB/S4END[5] Tile_X2Y6_LUT4AB/S4END[6] Tile_X2Y6_LUT4AB/S4END[7]
+ Tile_X2Y6_LUT4AB/S4END[8] Tile_X2Y6_LUT4AB/S4END[9] Tile_X2Y5_LUT4AB/S4END[0] Tile_X2Y5_LUT4AB/S4END[10]
+ Tile_X2Y5_LUT4AB/S4END[11] Tile_X2Y5_LUT4AB/S4END[12] Tile_X2Y5_LUT4AB/S4END[13]
+ Tile_X2Y5_LUT4AB/S4END[14] Tile_X2Y5_LUT4AB/S4END[15] Tile_X2Y5_LUT4AB/S4END[1]
+ Tile_X2Y5_LUT4AB/S4END[2] Tile_X2Y5_LUT4AB/S4END[3] Tile_X2Y5_LUT4AB/S4END[4] Tile_X2Y5_LUT4AB/S4END[5]
+ Tile_X2Y5_LUT4AB/S4END[6] Tile_X2Y5_LUT4AB/S4END[7] Tile_X2Y5_LUT4AB/S4END[8] Tile_X2Y5_LUT4AB/S4END[9]
+ Tile_X2Y6_LUT4AB/SS4END[0] Tile_X2Y6_LUT4AB/SS4END[10] Tile_X2Y6_LUT4AB/SS4END[11]
+ Tile_X2Y6_LUT4AB/SS4END[12] Tile_X2Y6_LUT4AB/SS4END[13] Tile_X2Y6_LUT4AB/SS4END[14]
+ Tile_X2Y6_LUT4AB/SS4END[15] Tile_X2Y6_LUT4AB/SS4END[1] Tile_X2Y6_LUT4AB/SS4END[2]
+ Tile_X2Y6_LUT4AB/SS4END[3] Tile_X2Y6_LUT4AB/SS4END[4] Tile_X2Y6_LUT4AB/SS4END[5]
+ Tile_X2Y6_LUT4AB/SS4END[6] Tile_X2Y6_LUT4AB/SS4END[7] Tile_X2Y6_LUT4AB/SS4END[8]
+ Tile_X2Y6_LUT4AB/SS4END[9] Tile_X2Y5_LUT4AB/SS4END[0] Tile_X2Y5_LUT4AB/SS4END[10]
+ Tile_X2Y5_LUT4AB/SS4END[11] Tile_X2Y5_LUT4AB/SS4END[12] Tile_X2Y5_LUT4AB/SS4END[13]
+ Tile_X2Y5_LUT4AB/SS4END[14] Tile_X2Y5_LUT4AB/SS4END[15] Tile_X2Y5_LUT4AB/SS4END[1]
+ Tile_X2Y5_LUT4AB/SS4END[2] Tile_X2Y5_LUT4AB/SS4END[3] Tile_X2Y5_LUT4AB/SS4END[4]
+ Tile_X2Y5_LUT4AB/SS4END[5] Tile_X2Y5_LUT4AB/SS4END[6] Tile_X2Y5_LUT4AB/SS4END[7]
+ Tile_X2Y5_LUT4AB/SS4END[8] Tile_X2Y5_LUT4AB/SS4END[9] Tile_X2Y5_LUT4AB/UserCLK Tile_X2Y4_LUT4AB/UserCLK
+ VGND VPWR Tile_X2Y5_LUT4AB/W1BEG[0] Tile_X2Y5_LUT4AB/W1BEG[1] Tile_X2Y5_LUT4AB/W1BEG[2]
+ Tile_X2Y5_LUT4AB/W1BEG[3] Tile_X3Y5_LUT4AB/W1BEG[0] Tile_X3Y5_LUT4AB/W1BEG[1] Tile_X3Y5_LUT4AB/W1BEG[2]
+ Tile_X3Y5_LUT4AB/W1BEG[3] Tile_X2Y5_LUT4AB/W2BEG[0] Tile_X2Y5_LUT4AB/W2BEG[1] Tile_X2Y5_LUT4AB/W2BEG[2]
+ Tile_X2Y5_LUT4AB/W2BEG[3] Tile_X2Y5_LUT4AB/W2BEG[4] Tile_X2Y5_LUT4AB/W2BEG[5] Tile_X2Y5_LUT4AB/W2BEG[6]
+ Tile_X2Y5_LUT4AB/W2BEG[7] Tile_X1Y5_LUT4AB/W2END[0] Tile_X1Y5_LUT4AB/W2END[1] Tile_X1Y5_LUT4AB/W2END[2]
+ Tile_X1Y5_LUT4AB/W2END[3] Tile_X1Y5_LUT4AB/W2END[4] Tile_X1Y5_LUT4AB/W2END[5] Tile_X1Y5_LUT4AB/W2END[6]
+ Tile_X1Y5_LUT4AB/W2END[7] Tile_X2Y5_LUT4AB/W2END[0] Tile_X2Y5_LUT4AB/W2END[1] Tile_X2Y5_LUT4AB/W2END[2]
+ Tile_X2Y5_LUT4AB/W2END[3] Tile_X2Y5_LUT4AB/W2END[4] Tile_X2Y5_LUT4AB/W2END[5] Tile_X2Y5_LUT4AB/W2END[6]
+ Tile_X2Y5_LUT4AB/W2END[7] Tile_X3Y5_LUT4AB/W2BEG[0] Tile_X3Y5_LUT4AB/W2BEG[1] Tile_X3Y5_LUT4AB/W2BEG[2]
+ Tile_X3Y5_LUT4AB/W2BEG[3] Tile_X3Y5_LUT4AB/W2BEG[4] Tile_X3Y5_LUT4AB/W2BEG[5] Tile_X3Y5_LUT4AB/W2BEG[6]
+ Tile_X3Y5_LUT4AB/W2BEG[7] Tile_X2Y5_LUT4AB/W6BEG[0] Tile_X2Y5_LUT4AB/W6BEG[10] Tile_X2Y5_LUT4AB/W6BEG[11]
+ Tile_X2Y5_LUT4AB/W6BEG[1] Tile_X2Y5_LUT4AB/W6BEG[2] Tile_X2Y5_LUT4AB/W6BEG[3] Tile_X2Y5_LUT4AB/W6BEG[4]
+ Tile_X2Y5_LUT4AB/W6BEG[5] Tile_X2Y5_LUT4AB/W6BEG[6] Tile_X2Y5_LUT4AB/W6BEG[7] Tile_X2Y5_LUT4AB/W6BEG[8]
+ Tile_X2Y5_LUT4AB/W6BEG[9] Tile_X3Y5_LUT4AB/W6BEG[0] Tile_X3Y5_LUT4AB/W6BEG[10] Tile_X3Y5_LUT4AB/W6BEG[11]
+ Tile_X3Y5_LUT4AB/W6BEG[1] Tile_X3Y5_LUT4AB/W6BEG[2] Tile_X3Y5_LUT4AB/W6BEG[3] Tile_X3Y5_LUT4AB/W6BEG[4]
+ Tile_X3Y5_LUT4AB/W6BEG[5] Tile_X3Y5_LUT4AB/W6BEG[6] Tile_X3Y5_LUT4AB/W6BEG[7] Tile_X3Y5_LUT4AB/W6BEG[8]
+ Tile_X3Y5_LUT4AB/W6BEG[9] Tile_X2Y5_LUT4AB/WW4BEG[0] Tile_X2Y5_LUT4AB/WW4BEG[10]
+ Tile_X2Y5_LUT4AB/WW4BEG[11] Tile_X2Y5_LUT4AB/WW4BEG[12] Tile_X2Y5_LUT4AB/WW4BEG[13]
+ Tile_X2Y5_LUT4AB/WW4BEG[14] Tile_X2Y5_LUT4AB/WW4BEG[15] Tile_X2Y5_LUT4AB/WW4BEG[1]
+ Tile_X2Y5_LUT4AB/WW4BEG[2] Tile_X2Y5_LUT4AB/WW4BEG[3] Tile_X2Y5_LUT4AB/WW4BEG[4]
+ Tile_X2Y5_LUT4AB/WW4BEG[5] Tile_X2Y5_LUT4AB/WW4BEG[6] Tile_X2Y5_LUT4AB/WW4BEG[7]
+ Tile_X2Y5_LUT4AB/WW4BEG[8] Tile_X2Y5_LUT4AB/WW4BEG[9] Tile_X3Y5_LUT4AB/WW4BEG[0]
+ Tile_X3Y5_LUT4AB/WW4BEG[10] Tile_X3Y5_LUT4AB/WW4BEG[11] Tile_X3Y5_LUT4AB/WW4BEG[12]
+ Tile_X3Y5_LUT4AB/WW4BEG[13] Tile_X3Y5_LUT4AB/WW4BEG[14] Tile_X3Y5_LUT4AB/WW4BEG[15]
+ Tile_X3Y5_LUT4AB/WW4BEG[1] Tile_X3Y5_LUT4AB/WW4BEG[2] Tile_X3Y5_LUT4AB/WW4BEG[3]
+ Tile_X3Y5_LUT4AB/WW4BEG[4] Tile_X3Y5_LUT4AB/WW4BEG[5] Tile_X3Y5_LUT4AB/WW4BEG[6]
+ Tile_X3Y5_LUT4AB/WW4BEG[7] Tile_X3Y5_LUT4AB/WW4BEG[8] Tile_X3Y5_LUT4AB/WW4BEG[9]
+ LUT4AB
XTile_X4Y0_N_IO4 Tile_X4Y0_A_I_top Tile_X4Y0_A_O_top Tile_X4Y0_A_T_top Tile_X4Y0_B_I_top
+ Tile_X4Y0_B_O_top Tile_X4Y0_B_T_top Tile_X4Y0_C_I_top Tile_X4Y0_C_O_top Tile_X4Y0_C_T_top
+ Tile_X4Y0_N_IO4/Ci Tile_X4Y0_D_I_top Tile_X4Y0_D_O_top Tile_X4Y0_D_T_top Tile_X4Y0_N_IO4/FrameData[0]
+ Tile_X4Y0_N_IO4/FrameData[10] Tile_X4Y0_N_IO4/FrameData[11] Tile_X4Y0_N_IO4/FrameData[12]
+ Tile_X4Y0_N_IO4/FrameData[13] Tile_X4Y0_N_IO4/FrameData[14] Tile_X4Y0_N_IO4/FrameData[15]
+ Tile_X4Y0_N_IO4/FrameData[16] Tile_X4Y0_N_IO4/FrameData[17] Tile_X4Y0_N_IO4/FrameData[18]
+ Tile_X4Y0_N_IO4/FrameData[19] Tile_X4Y0_N_IO4/FrameData[1] Tile_X4Y0_N_IO4/FrameData[20]
+ Tile_X4Y0_N_IO4/FrameData[21] Tile_X4Y0_N_IO4/FrameData[22] Tile_X4Y0_N_IO4/FrameData[23]
+ Tile_X4Y0_N_IO4/FrameData[24] Tile_X4Y0_N_IO4/FrameData[25] Tile_X4Y0_N_IO4/FrameData[26]
+ Tile_X4Y0_N_IO4/FrameData[27] Tile_X4Y0_N_IO4/FrameData[28] Tile_X4Y0_N_IO4/FrameData[29]
+ Tile_X4Y0_N_IO4/FrameData[2] Tile_X4Y0_N_IO4/FrameData[30] Tile_X4Y0_N_IO4/FrameData[31]
+ Tile_X4Y0_N_IO4/FrameData[3] Tile_X4Y0_N_IO4/FrameData[4] Tile_X4Y0_N_IO4/FrameData[5]
+ Tile_X4Y0_N_IO4/FrameData[6] Tile_X4Y0_N_IO4/FrameData[7] Tile_X4Y0_N_IO4/FrameData[8]
+ Tile_X4Y0_N_IO4/FrameData[9] Tile_X5Y0_NE_term/FrameData[0] Tile_X5Y0_NE_term/FrameData[10]
+ Tile_X5Y0_NE_term/FrameData[11] Tile_X5Y0_NE_term/FrameData[12] Tile_X5Y0_NE_term/FrameData[13]
+ Tile_X5Y0_NE_term/FrameData[14] Tile_X5Y0_NE_term/FrameData[15] Tile_X5Y0_NE_term/FrameData[16]
+ Tile_X5Y0_NE_term/FrameData[17] Tile_X5Y0_NE_term/FrameData[18] Tile_X5Y0_NE_term/FrameData[19]
+ Tile_X5Y0_NE_term/FrameData[1] Tile_X5Y0_NE_term/FrameData[20] Tile_X5Y0_NE_term/FrameData[21]
+ Tile_X5Y0_NE_term/FrameData[22] Tile_X5Y0_NE_term/FrameData[23] Tile_X5Y0_NE_term/FrameData[24]
+ Tile_X5Y0_NE_term/FrameData[25] Tile_X5Y0_NE_term/FrameData[26] Tile_X5Y0_NE_term/FrameData[27]
+ Tile_X5Y0_NE_term/FrameData[28] Tile_X5Y0_NE_term/FrameData[29] Tile_X5Y0_NE_term/FrameData[2]
+ Tile_X5Y0_NE_term/FrameData[30] Tile_X5Y0_NE_term/FrameData[31] Tile_X5Y0_NE_term/FrameData[3]
+ Tile_X5Y0_NE_term/FrameData[4] Tile_X5Y0_NE_term/FrameData[5] Tile_X5Y0_NE_term/FrameData[6]
+ Tile_X5Y0_NE_term/FrameData[7] Tile_X5Y0_NE_term/FrameData[8] Tile_X5Y0_NE_term/FrameData[9]
+ Tile_X4Y0_N_IO4/FrameStrobe[0] Tile_X4Y0_N_IO4/FrameStrobe[10] Tile_X4Y0_N_IO4/FrameStrobe[11]
+ Tile_X4Y0_N_IO4/FrameStrobe[12] Tile_X4Y0_N_IO4/FrameStrobe[13] Tile_X4Y0_N_IO4/FrameStrobe[14]
+ Tile_X4Y0_N_IO4/FrameStrobe[15] Tile_X4Y0_N_IO4/FrameStrobe[16] Tile_X4Y0_N_IO4/FrameStrobe[17]
+ Tile_X4Y0_N_IO4/FrameStrobe[18] Tile_X4Y0_N_IO4/FrameStrobe[19] Tile_X4Y0_N_IO4/FrameStrobe[1]
+ Tile_X4Y0_N_IO4/FrameStrobe[2] Tile_X4Y0_N_IO4/FrameStrobe[3] Tile_X4Y0_N_IO4/FrameStrobe[4]
+ Tile_X4Y0_N_IO4/FrameStrobe[5] Tile_X4Y0_N_IO4/FrameStrobe[6] Tile_X4Y0_N_IO4/FrameStrobe[7]
+ Tile_X4Y0_N_IO4/FrameStrobe[8] Tile_X4Y0_N_IO4/FrameStrobe[9] Tile_X4Y0_N_IO4/FrameStrobe_O[0]
+ Tile_X4Y0_N_IO4/FrameStrobe_O[10] Tile_X4Y0_N_IO4/FrameStrobe_O[11] Tile_X4Y0_N_IO4/FrameStrobe_O[12]
+ Tile_X4Y0_N_IO4/FrameStrobe_O[13] Tile_X4Y0_N_IO4/FrameStrobe_O[14] Tile_X4Y0_N_IO4/FrameStrobe_O[15]
+ Tile_X4Y0_N_IO4/FrameStrobe_O[16] Tile_X4Y0_N_IO4/FrameStrobe_O[17] Tile_X4Y0_N_IO4/FrameStrobe_O[18]
+ Tile_X4Y0_N_IO4/FrameStrobe_O[19] Tile_X4Y0_N_IO4/FrameStrobe_O[1] Tile_X4Y0_N_IO4/FrameStrobe_O[2]
+ Tile_X4Y0_N_IO4/FrameStrobe_O[3] Tile_X4Y0_N_IO4/FrameStrobe_O[4] Tile_X4Y0_N_IO4/FrameStrobe_O[5]
+ Tile_X4Y0_N_IO4/FrameStrobe_O[6] Tile_X4Y0_N_IO4/FrameStrobe_O[7] Tile_X4Y0_N_IO4/FrameStrobe_O[8]
+ Tile_X4Y0_N_IO4/FrameStrobe_O[9] Tile_X4Y0_N_IO4/N1END[0] Tile_X4Y0_N_IO4/N1END[1]
+ Tile_X4Y0_N_IO4/N1END[2] Tile_X4Y0_N_IO4/N1END[3] Tile_X4Y0_N_IO4/N2END[0] Tile_X4Y0_N_IO4/N2END[1]
+ Tile_X4Y0_N_IO4/N2END[2] Tile_X4Y0_N_IO4/N2END[3] Tile_X4Y0_N_IO4/N2END[4] Tile_X4Y0_N_IO4/N2END[5]
+ Tile_X4Y0_N_IO4/N2END[6] Tile_X4Y0_N_IO4/N2END[7] Tile_X4Y0_N_IO4/N2MID[0] Tile_X4Y0_N_IO4/N2MID[1]
+ Tile_X4Y0_N_IO4/N2MID[2] Tile_X4Y0_N_IO4/N2MID[3] Tile_X4Y0_N_IO4/N2MID[4] Tile_X4Y0_N_IO4/N2MID[5]
+ Tile_X4Y0_N_IO4/N2MID[6] Tile_X4Y0_N_IO4/N2MID[7] Tile_X4Y0_N_IO4/N4END[0] Tile_X4Y0_N_IO4/N4END[10]
+ Tile_X4Y0_N_IO4/N4END[11] Tile_X4Y0_N_IO4/N4END[12] Tile_X4Y0_N_IO4/N4END[13] Tile_X4Y0_N_IO4/N4END[14]
+ Tile_X4Y0_N_IO4/N4END[15] Tile_X4Y0_N_IO4/N4END[1] Tile_X4Y0_N_IO4/N4END[2] Tile_X4Y0_N_IO4/N4END[3]
+ Tile_X4Y0_N_IO4/N4END[4] Tile_X4Y0_N_IO4/N4END[5] Tile_X4Y0_N_IO4/N4END[6] Tile_X4Y0_N_IO4/N4END[7]
+ Tile_X4Y0_N_IO4/N4END[8] Tile_X4Y0_N_IO4/N4END[9] Tile_X4Y0_N_IO4/NN4END[0] Tile_X4Y0_N_IO4/NN4END[10]
+ Tile_X4Y0_N_IO4/NN4END[11] Tile_X4Y0_N_IO4/NN4END[12] Tile_X4Y0_N_IO4/NN4END[13]
+ Tile_X4Y0_N_IO4/NN4END[14] Tile_X4Y0_N_IO4/NN4END[15] Tile_X4Y0_N_IO4/NN4END[1]
+ Tile_X4Y0_N_IO4/NN4END[2] Tile_X4Y0_N_IO4/NN4END[3] Tile_X4Y0_N_IO4/NN4END[4] Tile_X4Y0_N_IO4/NN4END[5]
+ Tile_X4Y0_N_IO4/NN4END[6] Tile_X4Y0_N_IO4/NN4END[7] Tile_X4Y0_N_IO4/NN4END[8] Tile_X4Y0_N_IO4/NN4END[9]
+ Tile_X4Y0_N_IO4/S1BEG[0] Tile_X4Y0_N_IO4/S1BEG[1] Tile_X4Y0_N_IO4/S1BEG[2] Tile_X4Y0_N_IO4/S1BEG[3]
+ Tile_X4Y0_N_IO4/S2BEG[0] Tile_X4Y0_N_IO4/S2BEG[1] Tile_X4Y0_N_IO4/S2BEG[2] Tile_X4Y0_N_IO4/S2BEG[3]
+ Tile_X4Y0_N_IO4/S2BEG[4] Tile_X4Y0_N_IO4/S2BEG[5] Tile_X4Y0_N_IO4/S2BEG[6] Tile_X4Y0_N_IO4/S2BEG[7]
+ Tile_X4Y1_LUT4AB/S2END[0] Tile_X4Y1_LUT4AB/S2END[1] Tile_X4Y1_LUT4AB/S2END[2] Tile_X4Y1_LUT4AB/S2END[3]
+ Tile_X4Y1_LUT4AB/S2END[4] Tile_X4Y1_LUT4AB/S2END[5] Tile_X4Y1_LUT4AB/S2END[6] Tile_X4Y1_LUT4AB/S2END[7]
+ Tile_X4Y0_N_IO4/S4BEG[0] Tile_X4Y0_N_IO4/S4BEG[10] Tile_X4Y0_N_IO4/S4BEG[11] Tile_X4Y0_N_IO4/S4BEG[12]
+ Tile_X4Y0_N_IO4/S4BEG[13] Tile_X4Y0_N_IO4/S4BEG[14] Tile_X4Y0_N_IO4/S4BEG[15] Tile_X4Y0_N_IO4/S4BEG[1]
+ Tile_X4Y0_N_IO4/S4BEG[2] Tile_X4Y0_N_IO4/S4BEG[3] Tile_X4Y0_N_IO4/S4BEG[4] Tile_X4Y0_N_IO4/S4BEG[5]
+ Tile_X4Y0_N_IO4/S4BEG[6] Tile_X4Y0_N_IO4/S4BEG[7] Tile_X4Y0_N_IO4/S4BEG[8] Tile_X4Y0_N_IO4/S4BEG[9]
+ Tile_X4Y0_N_IO4/SS4BEG[0] Tile_X4Y0_N_IO4/SS4BEG[10] Tile_X4Y0_N_IO4/SS4BEG[11]
+ Tile_X4Y0_N_IO4/SS4BEG[12] Tile_X4Y0_N_IO4/SS4BEG[13] Tile_X4Y0_N_IO4/SS4BEG[14]
+ Tile_X4Y0_N_IO4/SS4BEG[15] Tile_X4Y0_N_IO4/SS4BEG[1] Tile_X4Y0_N_IO4/SS4BEG[2] Tile_X4Y0_N_IO4/SS4BEG[3]
+ Tile_X4Y0_N_IO4/SS4BEG[4] Tile_X4Y0_N_IO4/SS4BEG[5] Tile_X4Y0_N_IO4/SS4BEG[6] Tile_X4Y0_N_IO4/SS4BEG[7]
+ Tile_X4Y0_N_IO4/SS4BEG[8] Tile_X4Y0_N_IO4/SS4BEG[9] Tile_X4Y0_N_IO4/UserCLK Tile_X4Y0_N_IO4/UserCLKo
+ VGND VPWR N_IO4
XTile_X4Y3_LUT4AB Tile_X4Y4_LUT4AB/Co Tile_X4Y3_LUT4AB/Co Tile_X4Y3_LUT4AB/E1BEG[0]
+ Tile_X4Y3_LUT4AB/E1BEG[1] Tile_X4Y3_LUT4AB/E1BEG[2] Tile_X4Y3_LUT4AB/E1BEG[3] Tile_X4Y3_LUT4AB/E1END[0]
+ Tile_X4Y3_LUT4AB/E1END[1] Tile_X4Y3_LUT4AB/E1END[2] Tile_X4Y3_LUT4AB/E1END[3] Tile_X4Y3_LUT4AB/E2BEG[0]
+ Tile_X4Y3_LUT4AB/E2BEG[1] Tile_X4Y3_LUT4AB/E2BEG[2] Tile_X4Y3_LUT4AB/E2BEG[3] Tile_X4Y3_LUT4AB/E2BEG[4]
+ Tile_X4Y3_LUT4AB/E2BEG[5] Tile_X4Y3_LUT4AB/E2BEG[6] Tile_X4Y3_LUT4AB/E2BEG[7] Tile_X5Y3_E_TT_IF/E2END[0]
+ Tile_X5Y3_E_TT_IF/E2END[1] Tile_X5Y3_E_TT_IF/E2END[2] Tile_X5Y3_E_TT_IF/E2END[3]
+ Tile_X5Y3_E_TT_IF/E2END[4] Tile_X5Y3_E_TT_IF/E2END[5] Tile_X5Y3_E_TT_IF/E2END[6]
+ Tile_X5Y3_E_TT_IF/E2END[7] Tile_X4Y3_LUT4AB/E2END[0] Tile_X4Y3_LUT4AB/E2END[1] Tile_X4Y3_LUT4AB/E2END[2]
+ Tile_X4Y3_LUT4AB/E2END[3] Tile_X4Y3_LUT4AB/E2END[4] Tile_X4Y3_LUT4AB/E2END[5] Tile_X4Y3_LUT4AB/E2END[6]
+ Tile_X4Y3_LUT4AB/E2END[7] Tile_X4Y3_LUT4AB/E2MID[0] Tile_X4Y3_LUT4AB/E2MID[1] Tile_X4Y3_LUT4AB/E2MID[2]
+ Tile_X4Y3_LUT4AB/E2MID[3] Tile_X4Y3_LUT4AB/E2MID[4] Tile_X4Y3_LUT4AB/E2MID[5] Tile_X4Y3_LUT4AB/E2MID[6]
+ Tile_X4Y3_LUT4AB/E2MID[7] Tile_X4Y3_LUT4AB/E6BEG[0] Tile_X4Y3_LUT4AB/E6BEG[10] Tile_X4Y3_LUT4AB/E6BEG[11]
+ Tile_X4Y3_LUT4AB/E6BEG[1] Tile_X4Y3_LUT4AB/E6BEG[2] Tile_X4Y3_LUT4AB/E6BEG[3] Tile_X4Y3_LUT4AB/E6BEG[4]
+ Tile_X4Y3_LUT4AB/E6BEG[5] Tile_X4Y3_LUT4AB/E6BEG[6] Tile_X4Y3_LUT4AB/E6BEG[7] Tile_X4Y3_LUT4AB/E6BEG[8]
+ Tile_X4Y3_LUT4AB/E6BEG[9] Tile_X4Y3_LUT4AB/E6END[0] Tile_X4Y3_LUT4AB/E6END[10] Tile_X4Y3_LUT4AB/E6END[11]
+ Tile_X4Y3_LUT4AB/E6END[1] Tile_X4Y3_LUT4AB/E6END[2] Tile_X4Y3_LUT4AB/E6END[3] Tile_X4Y3_LUT4AB/E6END[4]
+ Tile_X4Y3_LUT4AB/E6END[5] Tile_X4Y3_LUT4AB/E6END[6] Tile_X4Y3_LUT4AB/E6END[7] Tile_X4Y3_LUT4AB/E6END[8]
+ Tile_X4Y3_LUT4AB/E6END[9] Tile_X4Y3_LUT4AB/EE4BEG[0] Tile_X4Y3_LUT4AB/EE4BEG[10]
+ Tile_X4Y3_LUT4AB/EE4BEG[11] Tile_X4Y3_LUT4AB/EE4BEG[12] Tile_X4Y3_LUT4AB/EE4BEG[13]
+ Tile_X4Y3_LUT4AB/EE4BEG[14] Tile_X4Y3_LUT4AB/EE4BEG[15] Tile_X4Y3_LUT4AB/EE4BEG[1]
+ Tile_X4Y3_LUT4AB/EE4BEG[2] Tile_X4Y3_LUT4AB/EE4BEG[3] Tile_X4Y3_LUT4AB/EE4BEG[4]
+ Tile_X4Y3_LUT4AB/EE4BEG[5] Tile_X4Y3_LUT4AB/EE4BEG[6] Tile_X4Y3_LUT4AB/EE4BEG[7]
+ Tile_X4Y3_LUT4AB/EE4BEG[8] Tile_X4Y3_LUT4AB/EE4BEG[9] Tile_X4Y3_LUT4AB/EE4END[0]
+ Tile_X4Y3_LUT4AB/EE4END[10] Tile_X4Y3_LUT4AB/EE4END[11] Tile_X4Y3_LUT4AB/EE4END[12]
+ Tile_X4Y3_LUT4AB/EE4END[13] Tile_X4Y3_LUT4AB/EE4END[14] Tile_X4Y3_LUT4AB/EE4END[15]
+ Tile_X4Y3_LUT4AB/EE4END[1] Tile_X4Y3_LUT4AB/EE4END[2] Tile_X4Y3_LUT4AB/EE4END[3]
+ Tile_X4Y3_LUT4AB/EE4END[4] Tile_X4Y3_LUT4AB/EE4END[5] Tile_X4Y3_LUT4AB/EE4END[6]
+ Tile_X4Y3_LUT4AB/EE4END[7] Tile_X4Y3_LUT4AB/EE4END[8] Tile_X4Y3_LUT4AB/EE4END[9]
+ Tile_X4Y3_LUT4AB/FrameData[0] Tile_X4Y3_LUT4AB/FrameData[10] Tile_X4Y3_LUT4AB/FrameData[11]
+ Tile_X4Y3_LUT4AB/FrameData[12] Tile_X4Y3_LUT4AB/FrameData[13] Tile_X4Y3_LUT4AB/FrameData[14]
+ Tile_X4Y3_LUT4AB/FrameData[15] Tile_X4Y3_LUT4AB/FrameData[16] Tile_X4Y3_LUT4AB/FrameData[17]
+ Tile_X4Y3_LUT4AB/FrameData[18] Tile_X4Y3_LUT4AB/FrameData[19] Tile_X4Y3_LUT4AB/FrameData[1]
+ Tile_X4Y3_LUT4AB/FrameData[20] Tile_X4Y3_LUT4AB/FrameData[21] Tile_X4Y3_LUT4AB/FrameData[22]
+ Tile_X4Y3_LUT4AB/FrameData[23] Tile_X4Y3_LUT4AB/FrameData[24] Tile_X4Y3_LUT4AB/FrameData[25]
+ Tile_X4Y3_LUT4AB/FrameData[26] Tile_X4Y3_LUT4AB/FrameData[27] Tile_X4Y3_LUT4AB/FrameData[28]
+ Tile_X4Y3_LUT4AB/FrameData[29] Tile_X4Y3_LUT4AB/FrameData[2] Tile_X4Y3_LUT4AB/FrameData[30]
+ Tile_X4Y3_LUT4AB/FrameData[31] Tile_X4Y3_LUT4AB/FrameData[3] Tile_X4Y3_LUT4AB/FrameData[4]
+ Tile_X4Y3_LUT4AB/FrameData[5] Tile_X4Y3_LUT4AB/FrameData[6] Tile_X4Y3_LUT4AB/FrameData[7]
+ Tile_X4Y3_LUT4AB/FrameData[8] Tile_X4Y3_LUT4AB/FrameData[9] Tile_X5Y3_E_TT_IF/FrameData[0]
+ Tile_X5Y3_E_TT_IF/FrameData[10] Tile_X5Y3_E_TT_IF/FrameData[11] Tile_X5Y3_E_TT_IF/FrameData[12]
+ Tile_X5Y3_E_TT_IF/FrameData[13] Tile_X5Y3_E_TT_IF/FrameData[14] Tile_X5Y3_E_TT_IF/FrameData[15]
+ Tile_X5Y3_E_TT_IF/FrameData[16] Tile_X5Y3_E_TT_IF/FrameData[17] Tile_X5Y3_E_TT_IF/FrameData[18]
+ Tile_X5Y3_E_TT_IF/FrameData[19] Tile_X5Y3_E_TT_IF/FrameData[1] Tile_X5Y3_E_TT_IF/FrameData[20]
+ Tile_X5Y3_E_TT_IF/FrameData[21] Tile_X5Y3_E_TT_IF/FrameData[22] Tile_X5Y3_E_TT_IF/FrameData[23]
+ Tile_X5Y3_E_TT_IF/FrameData[24] Tile_X5Y3_E_TT_IF/FrameData[25] Tile_X5Y3_E_TT_IF/FrameData[26]
+ Tile_X5Y3_E_TT_IF/FrameData[27] Tile_X5Y3_E_TT_IF/FrameData[28] Tile_X5Y3_E_TT_IF/FrameData[29]
+ Tile_X5Y3_E_TT_IF/FrameData[2] Tile_X5Y3_E_TT_IF/FrameData[30] Tile_X5Y3_E_TT_IF/FrameData[31]
+ Tile_X5Y3_E_TT_IF/FrameData[3] Tile_X5Y3_E_TT_IF/FrameData[4] Tile_X5Y3_E_TT_IF/FrameData[5]
+ Tile_X5Y3_E_TT_IF/FrameData[6] Tile_X5Y3_E_TT_IF/FrameData[7] Tile_X5Y3_E_TT_IF/FrameData[8]
+ Tile_X5Y3_E_TT_IF/FrameData[9] Tile_X4Y3_LUT4AB/FrameStrobe[0] Tile_X4Y3_LUT4AB/FrameStrobe[10]
+ Tile_X4Y3_LUT4AB/FrameStrobe[11] Tile_X4Y3_LUT4AB/FrameStrobe[12] Tile_X4Y3_LUT4AB/FrameStrobe[13]
+ Tile_X4Y3_LUT4AB/FrameStrobe[14] Tile_X4Y3_LUT4AB/FrameStrobe[15] Tile_X4Y3_LUT4AB/FrameStrobe[16]
+ Tile_X4Y3_LUT4AB/FrameStrobe[17] Tile_X4Y3_LUT4AB/FrameStrobe[18] Tile_X4Y3_LUT4AB/FrameStrobe[19]
+ Tile_X4Y3_LUT4AB/FrameStrobe[1] Tile_X4Y3_LUT4AB/FrameStrobe[2] Tile_X4Y3_LUT4AB/FrameStrobe[3]
+ Tile_X4Y3_LUT4AB/FrameStrobe[4] Tile_X4Y3_LUT4AB/FrameStrobe[5] Tile_X4Y3_LUT4AB/FrameStrobe[6]
+ Tile_X4Y3_LUT4AB/FrameStrobe[7] Tile_X4Y3_LUT4AB/FrameStrobe[8] Tile_X4Y3_LUT4AB/FrameStrobe[9]
+ Tile_X4Y2_LUT4AB/FrameStrobe[0] Tile_X4Y2_LUT4AB/FrameStrobe[10] Tile_X4Y2_LUT4AB/FrameStrobe[11]
+ Tile_X4Y2_LUT4AB/FrameStrobe[12] Tile_X4Y2_LUT4AB/FrameStrobe[13] Tile_X4Y2_LUT4AB/FrameStrobe[14]
+ Tile_X4Y2_LUT4AB/FrameStrobe[15] Tile_X4Y2_LUT4AB/FrameStrobe[16] Tile_X4Y2_LUT4AB/FrameStrobe[17]
+ Tile_X4Y2_LUT4AB/FrameStrobe[18] Tile_X4Y2_LUT4AB/FrameStrobe[19] Tile_X4Y2_LUT4AB/FrameStrobe[1]
+ Tile_X4Y2_LUT4AB/FrameStrobe[2] Tile_X4Y2_LUT4AB/FrameStrobe[3] Tile_X4Y2_LUT4AB/FrameStrobe[4]
+ Tile_X4Y2_LUT4AB/FrameStrobe[5] Tile_X4Y2_LUT4AB/FrameStrobe[6] Tile_X4Y2_LUT4AB/FrameStrobe[7]
+ Tile_X4Y2_LUT4AB/FrameStrobe[8] Tile_X4Y2_LUT4AB/FrameStrobe[9] Tile_X4Y3_LUT4AB/N1BEG[0]
+ Tile_X4Y3_LUT4AB/N1BEG[1] Tile_X4Y3_LUT4AB/N1BEG[2] Tile_X4Y3_LUT4AB/N1BEG[3] Tile_X4Y4_LUT4AB/N1BEG[0]
+ Tile_X4Y4_LUT4AB/N1BEG[1] Tile_X4Y4_LUT4AB/N1BEG[2] Tile_X4Y4_LUT4AB/N1BEG[3] Tile_X4Y3_LUT4AB/N2BEG[0]
+ Tile_X4Y3_LUT4AB/N2BEG[1] Tile_X4Y3_LUT4AB/N2BEG[2] Tile_X4Y3_LUT4AB/N2BEG[3] Tile_X4Y3_LUT4AB/N2BEG[4]
+ Tile_X4Y3_LUT4AB/N2BEG[5] Tile_X4Y3_LUT4AB/N2BEG[6] Tile_X4Y3_LUT4AB/N2BEG[7] Tile_X4Y2_LUT4AB/N2END[0]
+ Tile_X4Y2_LUT4AB/N2END[1] Tile_X4Y2_LUT4AB/N2END[2] Tile_X4Y2_LUT4AB/N2END[3] Tile_X4Y2_LUT4AB/N2END[4]
+ Tile_X4Y2_LUT4AB/N2END[5] Tile_X4Y2_LUT4AB/N2END[6] Tile_X4Y2_LUT4AB/N2END[7] Tile_X4Y3_LUT4AB/N2END[0]
+ Tile_X4Y3_LUT4AB/N2END[1] Tile_X4Y3_LUT4AB/N2END[2] Tile_X4Y3_LUT4AB/N2END[3] Tile_X4Y3_LUT4AB/N2END[4]
+ Tile_X4Y3_LUT4AB/N2END[5] Tile_X4Y3_LUT4AB/N2END[6] Tile_X4Y3_LUT4AB/N2END[7] Tile_X4Y4_LUT4AB/N2BEG[0]
+ Tile_X4Y4_LUT4AB/N2BEG[1] Tile_X4Y4_LUT4AB/N2BEG[2] Tile_X4Y4_LUT4AB/N2BEG[3] Tile_X4Y4_LUT4AB/N2BEG[4]
+ Tile_X4Y4_LUT4AB/N2BEG[5] Tile_X4Y4_LUT4AB/N2BEG[6] Tile_X4Y4_LUT4AB/N2BEG[7] Tile_X4Y3_LUT4AB/N4BEG[0]
+ Tile_X4Y3_LUT4AB/N4BEG[10] Tile_X4Y3_LUT4AB/N4BEG[11] Tile_X4Y3_LUT4AB/N4BEG[12]
+ Tile_X4Y3_LUT4AB/N4BEG[13] Tile_X4Y3_LUT4AB/N4BEG[14] Tile_X4Y3_LUT4AB/N4BEG[15]
+ Tile_X4Y3_LUT4AB/N4BEG[1] Tile_X4Y3_LUT4AB/N4BEG[2] Tile_X4Y3_LUT4AB/N4BEG[3] Tile_X4Y3_LUT4AB/N4BEG[4]
+ Tile_X4Y3_LUT4AB/N4BEG[5] Tile_X4Y3_LUT4AB/N4BEG[6] Tile_X4Y3_LUT4AB/N4BEG[7] Tile_X4Y3_LUT4AB/N4BEG[8]
+ Tile_X4Y3_LUT4AB/N4BEG[9] Tile_X4Y4_LUT4AB/N4BEG[0] Tile_X4Y4_LUT4AB/N4BEG[10] Tile_X4Y4_LUT4AB/N4BEG[11]
+ Tile_X4Y4_LUT4AB/N4BEG[12] Tile_X4Y4_LUT4AB/N4BEG[13] Tile_X4Y4_LUT4AB/N4BEG[14]
+ Tile_X4Y4_LUT4AB/N4BEG[15] Tile_X4Y4_LUT4AB/N4BEG[1] Tile_X4Y4_LUT4AB/N4BEG[2] Tile_X4Y4_LUT4AB/N4BEG[3]
+ Tile_X4Y4_LUT4AB/N4BEG[4] Tile_X4Y4_LUT4AB/N4BEG[5] Tile_X4Y4_LUT4AB/N4BEG[6] Tile_X4Y4_LUT4AB/N4BEG[7]
+ Tile_X4Y4_LUT4AB/N4BEG[8] Tile_X4Y4_LUT4AB/N4BEG[9] Tile_X4Y3_LUT4AB/NN4BEG[0] Tile_X4Y3_LUT4AB/NN4BEG[10]
+ Tile_X4Y3_LUT4AB/NN4BEG[11] Tile_X4Y3_LUT4AB/NN4BEG[12] Tile_X4Y3_LUT4AB/NN4BEG[13]
+ Tile_X4Y3_LUT4AB/NN4BEG[14] Tile_X4Y3_LUT4AB/NN4BEG[15] Tile_X4Y3_LUT4AB/NN4BEG[1]
+ Tile_X4Y3_LUT4AB/NN4BEG[2] Tile_X4Y3_LUT4AB/NN4BEG[3] Tile_X4Y3_LUT4AB/NN4BEG[4]
+ Tile_X4Y3_LUT4AB/NN4BEG[5] Tile_X4Y3_LUT4AB/NN4BEG[6] Tile_X4Y3_LUT4AB/NN4BEG[7]
+ Tile_X4Y3_LUT4AB/NN4BEG[8] Tile_X4Y3_LUT4AB/NN4BEG[9] Tile_X4Y4_LUT4AB/NN4BEG[0]
+ Tile_X4Y4_LUT4AB/NN4BEG[10] Tile_X4Y4_LUT4AB/NN4BEG[11] Tile_X4Y4_LUT4AB/NN4BEG[12]
+ Tile_X4Y4_LUT4AB/NN4BEG[13] Tile_X4Y4_LUT4AB/NN4BEG[14] Tile_X4Y4_LUT4AB/NN4BEG[15]
+ Tile_X4Y4_LUT4AB/NN4BEG[1] Tile_X4Y4_LUT4AB/NN4BEG[2] Tile_X4Y4_LUT4AB/NN4BEG[3]
+ Tile_X4Y4_LUT4AB/NN4BEG[4] Tile_X4Y4_LUT4AB/NN4BEG[5] Tile_X4Y4_LUT4AB/NN4BEG[6]
+ Tile_X4Y4_LUT4AB/NN4BEG[7] Tile_X4Y4_LUT4AB/NN4BEG[8] Tile_X4Y4_LUT4AB/NN4BEG[9]
+ Tile_X4Y4_LUT4AB/S1END[0] Tile_X4Y4_LUT4AB/S1END[1] Tile_X4Y4_LUT4AB/S1END[2] Tile_X4Y4_LUT4AB/S1END[3]
+ Tile_X4Y3_LUT4AB/S1END[0] Tile_X4Y3_LUT4AB/S1END[1] Tile_X4Y3_LUT4AB/S1END[2] Tile_X4Y3_LUT4AB/S1END[3]
+ Tile_X4Y4_LUT4AB/S2MID[0] Tile_X4Y4_LUT4AB/S2MID[1] Tile_X4Y4_LUT4AB/S2MID[2] Tile_X4Y4_LUT4AB/S2MID[3]
+ Tile_X4Y4_LUT4AB/S2MID[4] Tile_X4Y4_LUT4AB/S2MID[5] Tile_X4Y4_LUT4AB/S2MID[6] Tile_X4Y4_LUT4AB/S2MID[7]
+ Tile_X4Y4_LUT4AB/S2END[0] Tile_X4Y4_LUT4AB/S2END[1] Tile_X4Y4_LUT4AB/S2END[2] Tile_X4Y4_LUT4AB/S2END[3]
+ Tile_X4Y4_LUT4AB/S2END[4] Tile_X4Y4_LUT4AB/S2END[5] Tile_X4Y4_LUT4AB/S2END[6] Tile_X4Y4_LUT4AB/S2END[7]
+ Tile_X4Y3_LUT4AB/S2END[0] Tile_X4Y3_LUT4AB/S2END[1] Tile_X4Y3_LUT4AB/S2END[2] Tile_X4Y3_LUT4AB/S2END[3]
+ Tile_X4Y3_LUT4AB/S2END[4] Tile_X4Y3_LUT4AB/S2END[5] Tile_X4Y3_LUT4AB/S2END[6] Tile_X4Y3_LUT4AB/S2END[7]
+ Tile_X4Y3_LUT4AB/S2MID[0] Tile_X4Y3_LUT4AB/S2MID[1] Tile_X4Y3_LUT4AB/S2MID[2] Tile_X4Y3_LUT4AB/S2MID[3]
+ Tile_X4Y3_LUT4AB/S2MID[4] Tile_X4Y3_LUT4AB/S2MID[5] Tile_X4Y3_LUT4AB/S2MID[6] Tile_X4Y3_LUT4AB/S2MID[7]
+ Tile_X4Y4_LUT4AB/S4END[0] Tile_X4Y4_LUT4AB/S4END[10] Tile_X4Y4_LUT4AB/S4END[11]
+ Tile_X4Y4_LUT4AB/S4END[12] Tile_X4Y4_LUT4AB/S4END[13] Tile_X4Y4_LUT4AB/S4END[14]
+ Tile_X4Y4_LUT4AB/S4END[15] Tile_X4Y4_LUT4AB/S4END[1] Tile_X4Y4_LUT4AB/S4END[2] Tile_X4Y4_LUT4AB/S4END[3]
+ Tile_X4Y4_LUT4AB/S4END[4] Tile_X4Y4_LUT4AB/S4END[5] Tile_X4Y4_LUT4AB/S4END[6] Tile_X4Y4_LUT4AB/S4END[7]
+ Tile_X4Y4_LUT4AB/S4END[8] Tile_X4Y4_LUT4AB/S4END[9] Tile_X4Y3_LUT4AB/S4END[0] Tile_X4Y3_LUT4AB/S4END[10]
+ Tile_X4Y3_LUT4AB/S4END[11] Tile_X4Y3_LUT4AB/S4END[12] Tile_X4Y3_LUT4AB/S4END[13]
+ Tile_X4Y3_LUT4AB/S4END[14] Tile_X4Y3_LUT4AB/S4END[15] Tile_X4Y3_LUT4AB/S4END[1]
+ Tile_X4Y3_LUT4AB/S4END[2] Tile_X4Y3_LUT4AB/S4END[3] Tile_X4Y3_LUT4AB/S4END[4] Tile_X4Y3_LUT4AB/S4END[5]
+ Tile_X4Y3_LUT4AB/S4END[6] Tile_X4Y3_LUT4AB/S4END[7] Tile_X4Y3_LUT4AB/S4END[8] Tile_X4Y3_LUT4AB/S4END[9]
+ Tile_X4Y4_LUT4AB/SS4END[0] Tile_X4Y4_LUT4AB/SS4END[10] Tile_X4Y4_LUT4AB/SS4END[11]
+ Tile_X4Y4_LUT4AB/SS4END[12] Tile_X4Y4_LUT4AB/SS4END[13] Tile_X4Y4_LUT4AB/SS4END[14]
+ Tile_X4Y4_LUT4AB/SS4END[15] Tile_X4Y4_LUT4AB/SS4END[1] Tile_X4Y4_LUT4AB/SS4END[2]
+ Tile_X4Y4_LUT4AB/SS4END[3] Tile_X4Y4_LUT4AB/SS4END[4] Tile_X4Y4_LUT4AB/SS4END[5]
+ Tile_X4Y4_LUT4AB/SS4END[6] Tile_X4Y4_LUT4AB/SS4END[7] Tile_X4Y4_LUT4AB/SS4END[8]
+ Tile_X4Y4_LUT4AB/SS4END[9] Tile_X4Y3_LUT4AB/SS4END[0] Tile_X4Y3_LUT4AB/SS4END[10]
+ Tile_X4Y3_LUT4AB/SS4END[11] Tile_X4Y3_LUT4AB/SS4END[12] Tile_X4Y3_LUT4AB/SS4END[13]
+ Tile_X4Y3_LUT4AB/SS4END[14] Tile_X4Y3_LUT4AB/SS4END[15] Tile_X4Y3_LUT4AB/SS4END[1]
+ Tile_X4Y3_LUT4AB/SS4END[2] Tile_X4Y3_LUT4AB/SS4END[3] Tile_X4Y3_LUT4AB/SS4END[4]
+ Tile_X4Y3_LUT4AB/SS4END[5] Tile_X4Y3_LUT4AB/SS4END[6] Tile_X4Y3_LUT4AB/SS4END[7]
+ Tile_X4Y3_LUT4AB/SS4END[8] Tile_X4Y3_LUT4AB/SS4END[9] Tile_X4Y3_LUT4AB/UserCLK Tile_X4Y2_LUT4AB/UserCLK
+ VGND VPWR Tile_X4Y3_LUT4AB/W1BEG[0] Tile_X4Y3_LUT4AB/W1BEG[1] Tile_X4Y3_LUT4AB/W1BEG[2]
+ Tile_X4Y3_LUT4AB/W1BEG[3] Tile_X4Y3_LUT4AB/W1END[0] Tile_X4Y3_LUT4AB/W1END[1] Tile_X4Y3_LUT4AB/W1END[2]
+ Tile_X4Y3_LUT4AB/W1END[3] Tile_X4Y3_LUT4AB/W2BEG[0] Tile_X4Y3_LUT4AB/W2BEG[1] Tile_X4Y3_LUT4AB/W2BEG[2]
+ Tile_X4Y3_LUT4AB/W2BEG[3] Tile_X4Y3_LUT4AB/W2BEG[4] Tile_X4Y3_LUT4AB/W2BEG[5] Tile_X4Y3_LUT4AB/W2BEG[6]
+ Tile_X4Y3_LUT4AB/W2BEG[7] Tile_X3Y3_LUT4AB/W2END[0] Tile_X3Y3_LUT4AB/W2END[1] Tile_X3Y3_LUT4AB/W2END[2]
+ Tile_X3Y3_LUT4AB/W2END[3] Tile_X3Y3_LUT4AB/W2END[4] Tile_X3Y3_LUT4AB/W2END[5] Tile_X3Y3_LUT4AB/W2END[6]
+ Tile_X3Y3_LUT4AB/W2END[7] Tile_X4Y3_LUT4AB/W2END[0] Tile_X4Y3_LUT4AB/W2END[1] Tile_X4Y3_LUT4AB/W2END[2]
+ Tile_X4Y3_LUT4AB/W2END[3] Tile_X4Y3_LUT4AB/W2END[4] Tile_X4Y3_LUT4AB/W2END[5] Tile_X4Y3_LUT4AB/W2END[6]
+ Tile_X4Y3_LUT4AB/W2END[7] Tile_X4Y3_LUT4AB/W2MID[0] Tile_X4Y3_LUT4AB/W2MID[1] Tile_X4Y3_LUT4AB/W2MID[2]
+ Tile_X4Y3_LUT4AB/W2MID[3] Tile_X4Y3_LUT4AB/W2MID[4] Tile_X4Y3_LUT4AB/W2MID[5] Tile_X4Y3_LUT4AB/W2MID[6]
+ Tile_X4Y3_LUT4AB/W2MID[7] Tile_X4Y3_LUT4AB/W6BEG[0] Tile_X4Y3_LUT4AB/W6BEG[10] Tile_X4Y3_LUT4AB/W6BEG[11]
+ Tile_X4Y3_LUT4AB/W6BEG[1] Tile_X4Y3_LUT4AB/W6BEG[2] Tile_X4Y3_LUT4AB/W6BEG[3] Tile_X4Y3_LUT4AB/W6BEG[4]
+ Tile_X4Y3_LUT4AB/W6BEG[5] Tile_X4Y3_LUT4AB/W6BEG[6] Tile_X4Y3_LUT4AB/W6BEG[7] Tile_X4Y3_LUT4AB/W6BEG[8]
+ Tile_X4Y3_LUT4AB/W6BEG[9] Tile_X4Y3_LUT4AB/W6END[0] Tile_X4Y3_LUT4AB/W6END[10] Tile_X4Y3_LUT4AB/W6END[11]
+ Tile_X4Y3_LUT4AB/W6END[1] Tile_X4Y3_LUT4AB/W6END[2] Tile_X4Y3_LUT4AB/W6END[3] Tile_X4Y3_LUT4AB/W6END[4]
+ Tile_X4Y3_LUT4AB/W6END[5] Tile_X4Y3_LUT4AB/W6END[6] Tile_X4Y3_LUT4AB/W6END[7] Tile_X4Y3_LUT4AB/W6END[8]
+ Tile_X4Y3_LUT4AB/W6END[9] Tile_X4Y3_LUT4AB/WW4BEG[0] Tile_X4Y3_LUT4AB/WW4BEG[10]
+ Tile_X4Y3_LUT4AB/WW4BEG[11] Tile_X4Y3_LUT4AB/WW4BEG[12] Tile_X4Y3_LUT4AB/WW4BEG[13]
+ Tile_X4Y3_LUT4AB/WW4BEG[14] Tile_X4Y3_LUT4AB/WW4BEG[15] Tile_X4Y3_LUT4AB/WW4BEG[1]
+ Tile_X4Y3_LUT4AB/WW4BEG[2] Tile_X4Y3_LUT4AB/WW4BEG[3] Tile_X4Y3_LUT4AB/WW4BEG[4]
+ Tile_X4Y3_LUT4AB/WW4BEG[5] Tile_X4Y3_LUT4AB/WW4BEG[6] Tile_X4Y3_LUT4AB/WW4BEG[7]
+ Tile_X4Y3_LUT4AB/WW4BEG[8] Tile_X4Y3_LUT4AB/WW4BEG[9] Tile_X4Y3_LUT4AB/WW4END[0]
+ Tile_X4Y3_LUT4AB/WW4END[10] Tile_X4Y3_LUT4AB/WW4END[11] Tile_X4Y3_LUT4AB/WW4END[12]
+ Tile_X4Y3_LUT4AB/WW4END[13] Tile_X4Y3_LUT4AB/WW4END[14] Tile_X4Y3_LUT4AB/WW4END[15]
+ Tile_X4Y3_LUT4AB/WW4END[1] Tile_X4Y3_LUT4AB/WW4END[2] Tile_X4Y3_LUT4AB/WW4END[3]
+ Tile_X4Y3_LUT4AB/WW4END[4] Tile_X4Y3_LUT4AB/WW4END[5] Tile_X4Y3_LUT4AB/WW4END[6]
+ Tile_X4Y3_LUT4AB/WW4END[7] Tile_X4Y3_LUT4AB/WW4END[8] Tile_X4Y3_LUT4AB/WW4END[9]
+ LUT4AB
XTile_X5Y5_E_TT_IF Tile_X5Y5_CLK_TT_PROJECT Tile_X4Y5_LUT4AB/E1BEG[0] Tile_X4Y5_LUT4AB/E1BEG[1]
+ Tile_X4Y5_LUT4AB/E1BEG[2] Tile_X4Y5_LUT4AB/E1BEG[3] Tile_X5Y5_E_TT_IF/E2END[0] Tile_X5Y5_E_TT_IF/E2END[1]
+ Tile_X5Y5_E_TT_IF/E2END[2] Tile_X5Y5_E_TT_IF/E2END[3] Tile_X5Y5_E_TT_IF/E2END[4]
+ Tile_X5Y5_E_TT_IF/E2END[5] Tile_X5Y5_E_TT_IF/E2END[6] Tile_X5Y5_E_TT_IF/E2END[7]
+ Tile_X4Y5_LUT4AB/E2BEG[0] Tile_X4Y5_LUT4AB/E2BEG[1] Tile_X4Y5_LUT4AB/E2BEG[2] Tile_X4Y5_LUT4AB/E2BEG[3]
+ Tile_X4Y5_LUT4AB/E2BEG[4] Tile_X4Y5_LUT4AB/E2BEG[5] Tile_X4Y5_LUT4AB/E2BEG[6] Tile_X4Y5_LUT4AB/E2BEG[7]
+ Tile_X4Y5_LUT4AB/E6BEG[0] Tile_X4Y5_LUT4AB/E6BEG[10] Tile_X4Y5_LUT4AB/E6BEG[11]
+ Tile_X4Y5_LUT4AB/E6BEG[1] Tile_X4Y5_LUT4AB/E6BEG[2] Tile_X4Y5_LUT4AB/E6BEG[3] Tile_X4Y5_LUT4AB/E6BEG[4]
+ Tile_X4Y5_LUT4AB/E6BEG[5] Tile_X4Y5_LUT4AB/E6BEG[6] Tile_X4Y5_LUT4AB/E6BEG[7] Tile_X4Y5_LUT4AB/E6BEG[8]
+ Tile_X4Y5_LUT4AB/E6BEG[9] Tile_X4Y5_LUT4AB/EE4BEG[0] Tile_X4Y5_LUT4AB/EE4BEG[10]
+ Tile_X4Y5_LUT4AB/EE4BEG[11] Tile_X4Y5_LUT4AB/EE4BEG[12] Tile_X4Y5_LUT4AB/EE4BEG[13]
+ Tile_X4Y5_LUT4AB/EE4BEG[14] Tile_X4Y5_LUT4AB/EE4BEG[15] Tile_X4Y5_LUT4AB/EE4BEG[1]
+ Tile_X4Y5_LUT4AB/EE4BEG[2] Tile_X4Y5_LUT4AB/EE4BEG[3] Tile_X4Y5_LUT4AB/EE4BEG[4]
+ Tile_X4Y5_LUT4AB/EE4BEG[5] Tile_X4Y5_LUT4AB/EE4BEG[6] Tile_X4Y5_LUT4AB/EE4BEG[7]
+ Tile_X4Y5_LUT4AB/EE4BEG[8] Tile_X4Y5_LUT4AB/EE4BEG[9] Tile_X5Y5_ENA_TT_PROJECT Tile_X5Y5_E_TT_IF/FrameData[0]
+ Tile_X5Y5_E_TT_IF/FrameData[10] Tile_X5Y5_E_TT_IF/FrameData[11] Tile_X5Y5_E_TT_IF/FrameData[12]
+ Tile_X5Y5_E_TT_IF/FrameData[13] Tile_X5Y5_E_TT_IF/FrameData[14] Tile_X5Y5_E_TT_IF/FrameData[15]
+ Tile_X5Y5_E_TT_IF/FrameData[16] Tile_X5Y5_E_TT_IF/FrameData[17] Tile_X5Y5_E_TT_IF/FrameData[18]
+ Tile_X5Y5_E_TT_IF/FrameData[19] Tile_X5Y5_E_TT_IF/FrameData[1] Tile_X5Y5_E_TT_IF/FrameData[20]
+ Tile_X5Y5_E_TT_IF/FrameData[21] Tile_X5Y5_E_TT_IF/FrameData[22] Tile_X5Y5_E_TT_IF/FrameData[23]
+ Tile_X5Y5_E_TT_IF/FrameData[24] Tile_X5Y5_E_TT_IF/FrameData[25] Tile_X5Y5_E_TT_IF/FrameData[26]
+ Tile_X5Y5_E_TT_IF/FrameData[27] Tile_X5Y5_E_TT_IF/FrameData[28] Tile_X5Y5_E_TT_IF/FrameData[29]
+ Tile_X5Y5_E_TT_IF/FrameData[2] Tile_X5Y5_E_TT_IF/FrameData[30] Tile_X5Y5_E_TT_IF/FrameData[31]
+ Tile_X5Y5_E_TT_IF/FrameData[3] Tile_X5Y5_E_TT_IF/FrameData[4] Tile_X5Y5_E_TT_IF/FrameData[5]
+ Tile_X5Y5_E_TT_IF/FrameData[6] Tile_X5Y5_E_TT_IF/FrameData[7] Tile_X5Y5_E_TT_IF/FrameData[8]
+ Tile_X5Y5_E_TT_IF/FrameData[9] Tile_X5Y5_E_TT_IF/FrameData_O[0] Tile_X5Y5_E_TT_IF/FrameData_O[10]
+ Tile_X5Y5_E_TT_IF/FrameData_O[11] Tile_X5Y5_E_TT_IF/FrameData_O[12] Tile_X5Y5_E_TT_IF/FrameData_O[13]
+ Tile_X5Y5_E_TT_IF/FrameData_O[14] Tile_X5Y5_E_TT_IF/FrameData_O[15] Tile_X5Y5_E_TT_IF/FrameData_O[16]
+ Tile_X5Y5_E_TT_IF/FrameData_O[17] Tile_X5Y5_E_TT_IF/FrameData_O[18] Tile_X5Y5_E_TT_IF/FrameData_O[19]
+ Tile_X5Y5_E_TT_IF/FrameData_O[1] Tile_X5Y5_E_TT_IF/FrameData_O[20] Tile_X5Y5_E_TT_IF/FrameData_O[21]
+ Tile_X5Y5_E_TT_IF/FrameData_O[22] Tile_X5Y5_E_TT_IF/FrameData_O[23] Tile_X5Y5_E_TT_IF/FrameData_O[24]
+ Tile_X5Y5_E_TT_IF/FrameData_O[25] Tile_X5Y5_E_TT_IF/FrameData_O[26] Tile_X5Y5_E_TT_IF/FrameData_O[27]
+ Tile_X5Y5_E_TT_IF/FrameData_O[28] Tile_X5Y5_E_TT_IF/FrameData_O[29] Tile_X5Y5_E_TT_IF/FrameData_O[2]
+ Tile_X5Y5_E_TT_IF/FrameData_O[30] Tile_X5Y5_E_TT_IF/FrameData_O[31] Tile_X5Y5_E_TT_IF/FrameData_O[3]
+ Tile_X5Y5_E_TT_IF/FrameData_O[4] Tile_X5Y5_E_TT_IF/FrameData_O[5] Tile_X5Y5_E_TT_IF/FrameData_O[6]
+ Tile_X5Y5_E_TT_IF/FrameData_O[7] Tile_X5Y5_E_TT_IF/FrameData_O[8] Tile_X5Y5_E_TT_IF/FrameData_O[9]
+ Tile_X5Y5_E_TT_IF/FrameStrobe[0] Tile_X5Y5_E_TT_IF/FrameStrobe[10] Tile_X5Y5_E_TT_IF/FrameStrobe[11]
+ Tile_X5Y5_E_TT_IF/FrameStrobe[12] Tile_X5Y5_E_TT_IF/FrameStrobe[13] Tile_X5Y5_E_TT_IF/FrameStrobe[14]
+ Tile_X5Y5_E_TT_IF/FrameStrobe[15] Tile_X5Y5_E_TT_IF/FrameStrobe[16] Tile_X5Y5_E_TT_IF/FrameStrobe[17]
+ Tile_X5Y5_E_TT_IF/FrameStrobe[18] Tile_X5Y5_E_TT_IF/FrameStrobe[19] Tile_X5Y5_E_TT_IF/FrameStrobe[1]
+ Tile_X5Y5_E_TT_IF/FrameStrobe[2] Tile_X5Y5_E_TT_IF/FrameStrobe[3] Tile_X5Y5_E_TT_IF/FrameStrobe[4]
+ Tile_X5Y5_E_TT_IF/FrameStrobe[5] Tile_X5Y5_E_TT_IF/FrameStrobe[6] Tile_X5Y5_E_TT_IF/FrameStrobe[7]
+ Tile_X5Y5_E_TT_IF/FrameStrobe[8] Tile_X5Y5_E_TT_IF/FrameStrobe[9] Tile_X5Y4_E_TT_IF/FrameStrobe[0]
+ Tile_X5Y4_E_TT_IF/FrameStrobe[10] Tile_X5Y4_E_TT_IF/FrameStrobe[11] Tile_X5Y4_E_TT_IF/FrameStrobe[12]
+ Tile_X5Y4_E_TT_IF/FrameStrobe[13] Tile_X5Y4_E_TT_IF/FrameStrobe[14] Tile_X5Y4_E_TT_IF/FrameStrobe[15]
+ Tile_X5Y4_E_TT_IF/FrameStrobe[16] Tile_X5Y4_E_TT_IF/FrameStrobe[17] Tile_X5Y4_E_TT_IF/FrameStrobe[18]
+ Tile_X5Y4_E_TT_IF/FrameStrobe[19] Tile_X5Y4_E_TT_IF/FrameStrobe[1] Tile_X5Y4_E_TT_IF/FrameStrobe[2]
+ Tile_X5Y4_E_TT_IF/FrameStrobe[3] Tile_X5Y4_E_TT_IF/FrameStrobe[4] Tile_X5Y4_E_TT_IF/FrameStrobe[5]
+ Tile_X5Y4_E_TT_IF/FrameStrobe[6] Tile_X5Y4_E_TT_IF/FrameStrobe[7] Tile_X5Y4_E_TT_IF/FrameStrobe[8]
+ Tile_X5Y4_E_TT_IF/FrameStrobe[9] Tile_X5Y5_E_TT_IF/N1BEG[0] Tile_X5Y5_E_TT_IF/N1BEG[1]
+ Tile_X5Y5_E_TT_IF/N1BEG[2] Tile_X5Y5_E_TT_IF/N1BEG[3] Tile_X5Y6_E_TT_IF/N1BEG[0]
+ Tile_X5Y6_E_TT_IF/N1BEG[1] Tile_X5Y6_E_TT_IF/N1BEG[2] Tile_X5Y6_E_TT_IF/N1BEG[3]
+ Tile_X5Y5_E_TT_IF/N2BEG[0] Tile_X5Y5_E_TT_IF/N2BEG[1] Tile_X5Y5_E_TT_IF/N2BEG[2]
+ Tile_X5Y5_E_TT_IF/N2BEG[3] Tile_X5Y5_E_TT_IF/N2BEG[4] Tile_X5Y5_E_TT_IF/N2BEG[5]
+ Tile_X5Y5_E_TT_IF/N2BEG[6] Tile_X5Y5_E_TT_IF/N2BEG[7] Tile_X5Y4_E_TT_IF/N2END[0]
+ Tile_X5Y4_E_TT_IF/N2END[1] Tile_X5Y4_E_TT_IF/N2END[2] Tile_X5Y4_E_TT_IF/N2END[3]
+ Tile_X5Y4_E_TT_IF/N2END[4] Tile_X5Y4_E_TT_IF/N2END[5] Tile_X5Y4_E_TT_IF/N2END[6]
+ Tile_X5Y4_E_TT_IF/N2END[7] Tile_X5Y5_E_TT_IF/N2END[0] Tile_X5Y5_E_TT_IF/N2END[1]
+ Tile_X5Y5_E_TT_IF/N2END[2] Tile_X5Y5_E_TT_IF/N2END[3] Tile_X5Y5_E_TT_IF/N2END[4]
+ Tile_X5Y5_E_TT_IF/N2END[5] Tile_X5Y5_E_TT_IF/N2END[6] Tile_X5Y5_E_TT_IF/N2END[7]
+ Tile_X5Y6_E_TT_IF/N2BEG[0] Tile_X5Y6_E_TT_IF/N2BEG[1] Tile_X5Y6_E_TT_IF/N2BEG[2]
+ Tile_X5Y6_E_TT_IF/N2BEG[3] Tile_X5Y6_E_TT_IF/N2BEG[4] Tile_X5Y6_E_TT_IF/N2BEG[5]
+ Tile_X5Y6_E_TT_IF/N2BEG[6] Tile_X5Y6_E_TT_IF/N2BEG[7] Tile_X5Y5_E_TT_IF/N4BEG[0]
+ Tile_X5Y5_E_TT_IF/N4BEG[10] Tile_X5Y5_E_TT_IF/N4BEG[11] Tile_X5Y5_E_TT_IF/N4BEG[12]
+ Tile_X5Y5_E_TT_IF/N4BEG[13] Tile_X5Y5_E_TT_IF/N4BEG[14] Tile_X5Y5_E_TT_IF/N4BEG[15]
+ Tile_X5Y5_E_TT_IF/N4BEG[1] Tile_X5Y5_E_TT_IF/N4BEG[2] Tile_X5Y5_E_TT_IF/N4BEG[3]
+ Tile_X5Y5_E_TT_IF/N4BEG[4] Tile_X5Y5_E_TT_IF/N4BEG[5] Tile_X5Y5_E_TT_IF/N4BEG[6]
+ Tile_X5Y5_E_TT_IF/N4BEG[7] Tile_X5Y5_E_TT_IF/N4BEG[8] Tile_X5Y5_E_TT_IF/N4BEG[9]
+ Tile_X5Y6_E_TT_IF/N4BEG[0] Tile_X5Y6_E_TT_IF/N4BEG[10] Tile_X5Y6_E_TT_IF/N4BEG[11]
+ Tile_X5Y6_E_TT_IF/N4BEG[12] Tile_X5Y6_E_TT_IF/N4BEG[13] Tile_X5Y6_E_TT_IF/N4BEG[14]
+ Tile_X5Y6_E_TT_IF/N4BEG[15] Tile_X5Y6_E_TT_IF/N4BEG[1] Tile_X5Y6_E_TT_IF/N4BEG[2]
+ Tile_X5Y6_E_TT_IF/N4BEG[3] Tile_X5Y6_E_TT_IF/N4BEG[4] Tile_X5Y6_E_TT_IF/N4BEG[5]
+ Tile_X5Y6_E_TT_IF/N4BEG[6] Tile_X5Y6_E_TT_IF/N4BEG[7] Tile_X5Y6_E_TT_IF/N4BEG[8]
+ Tile_X5Y6_E_TT_IF/N4BEG[9] Tile_X5Y5_RST_N_TT_PROJECT Tile_X5Y6_E_TT_IF/S1END[0]
+ Tile_X5Y6_E_TT_IF/S1END[1] Tile_X5Y6_E_TT_IF/S1END[2] Tile_X5Y6_E_TT_IF/S1END[3]
+ Tile_X5Y5_E_TT_IF/S1END[0] Tile_X5Y5_E_TT_IF/S1END[1] Tile_X5Y5_E_TT_IF/S1END[2]
+ Tile_X5Y5_E_TT_IF/S1END[3] Tile_X5Y6_E_TT_IF/S2MID[0] Tile_X5Y6_E_TT_IF/S2MID[1]
+ Tile_X5Y6_E_TT_IF/S2MID[2] Tile_X5Y6_E_TT_IF/S2MID[3] Tile_X5Y6_E_TT_IF/S2MID[4]
+ Tile_X5Y6_E_TT_IF/S2MID[5] Tile_X5Y6_E_TT_IF/S2MID[6] Tile_X5Y6_E_TT_IF/S2MID[7]
+ Tile_X5Y6_E_TT_IF/S2END[0] Tile_X5Y6_E_TT_IF/S2END[1] Tile_X5Y6_E_TT_IF/S2END[2]
+ Tile_X5Y6_E_TT_IF/S2END[3] Tile_X5Y6_E_TT_IF/S2END[4] Tile_X5Y6_E_TT_IF/S2END[5]
+ Tile_X5Y6_E_TT_IF/S2END[6] Tile_X5Y6_E_TT_IF/S2END[7] Tile_X5Y5_E_TT_IF/S2END[0]
+ Tile_X5Y5_E_TT_IF/S2END[1] Tile_X5Y5_E_TT_IF/S2END[2] Tile_X5Y5_E_TT_IF/S2END[3]
+ Tile_X5Y5_E_TT_IF/S2END[4] Tile_X5Y5_E_TT_IF/S2END[5] Tile_X5Y5_E_TT_IF/S2END[6]
+ Tile_X5Y5_E_TT_IF/S2END[7] Tile_X5Y5_E_TT_IF/S2MID[0] Tile_X5Y5_E_TT_IF/S2MID[1]
+ Tile_X5Y5_E_TT_IF/S2MID[2] Tile_X5Y5_E_TT_IF/S2MID[3] Tile_X5Y5_E_TT_IF/S2MID[4]
+ Tile_X5Y5_E_TT_IF/S2MID[5] Tile_X5Y5_E_TT_IF/S2MID[6] Tile_X5Y5_E_TT_IF/S2MID[7]
+ Tile_X5Y6_E_TT_IF/S4END[0] Tile_X5Y6_E_TT_IF/S4END[10] Tile_X5Y6_E_TT_IF/S4END[11]
+ Tile_X5Y6_E_TT_IF/S4END[12] Tile_X5Y6_E_TT_IF/S4END[13] Tile_X5Y6_E_TT_IF/S4END[14]
+ Tile_X5Y6_E_TT_IF/S4END[15] Tile_X5Y6_E_TT_IF/S4END[1] Tile_X5Y6_E_TT_IF/S4END[2]
+ Tile_X5Y6_E_TT_IF/S4END[3] Tile_X5Y6_E_TT_IF/S4END[4] Tile_X5Y6_E_TT_IF/S4END[5]
+ Tile_X5Y6_E_TT_IF/S4END[6] Tile_X5Y6_E_TT_IF/S4END[7] Tile_X5Y6_E_TT_IF/S4END[8]
+ Tile_X5Y6_E_TT_IF/S4END[9] Tile_X5Y5_E_TT_IF/S4END[0] Tile_X5Y5_E_TT_IF/S4END[10]
+ Tile_X5Y5_E_TT_IF/S4END[11] Tile_X5Y5_E_TT_IF/S4END[12] Tile_X5Y5_E_TT_IF/S4END[13]
+ Tile_X5Y5_E_TT_IF/S4END[14] Tile_X5Y5_E_TT_IF/S4END[15] Tile_X5Y5_E_TT_IF/S4END[1]
+ Tile_X5Y5_E_TT_IF/S4END[2] Tile_X5Y5_E_TT_IF/S4END[3] Tile_X5Y5_E_TT_IF/S4END[4]
+ Tile_X5Y5_E_TT_IF/S4END[5] Tile_X5Y5_E_TT_IF/S4END[6] Tile_X5Y5_E_TT_IF/S4END[7]
+ Tile_X5Y5_E_TT_IF/S4END[8] Tile_X5Y5_E_TT_IF/S4END[9] Tile_X5Y5_UIO_IN_TT_PROJECT0
+ Tile_X5Y5_UIO_IN_TT_PROJECT1 Tile_X5Y5_UIO_IN_TT_PROJECT2 Tile_X5Y5_UIO_IN_TT_PROJECT3
+ Tile_X5Y5_UIO_IN_TT_PROJECT4 Tile_X5Y5_UIO_IN_TT_PROJECT5 Tile_X5Y5_UIO_IN_TT_PROJECT6
+ Tile_X5Y5_UIO_IN_TT_PROJECT7 Tile_X5Y5_UIO_OE_TT_PROJECT0 Tile_X5Y5_UIO_OE_TT_PROJECT1
+ Tile_X5Y5_UIO_OE_TT_PROJECT2 Tile_X5Y5_UIO_OE_TT_PROJECT3 Tile_X5Y5_UIO_OE_TT_PROJECT4
+ Tile_X5Y5_UIO_OE_TT_PROJECT5 Tile_X5Y5_UIO_OE_TT_PROJECT6 Tile_X5Y5_UIO_OE_TT_PROJECT7
+ Tile_X5Y5_UIO_OUT_TT_PROJECT0 Tile_X5Y5_UIO_OUT_TT_PROJECT1 Tile_X5Y5_UIO_OUT_TT_PROJECT2
+ Tile_X5Y5_UIO_OUT_TT_PROJECT3 Tile_X5Y5_UIO_OUT_TT_PROJECT4 Tile_X5Y5_UIO_OUT_TT_PROJECT5
+ Tile_X5Y5_UIO_OUT_TT_PROJECT6 Tile_X5Y5_UIO_OUT_TT_PROJECT7 Tile_X5Y5_UI_IN_TT_PROJECT0
+ Tile_X5Y5_UI_IN_TT_PROJECT1 Tile_X5Y5_UI_IN_TT_PROJECT2 Tile_X5Y5_UI_IN_TT_PROJECT3
+ Tile_X5Y5_UI_IN_TT_PROJECT4 Tile_X5Y5_UI_IN_TT_PROJECT5 Tile_X5Y5_UI_IN_TT_PROJECT6
+ Tile_X5Y5_UI_IN_TT_PROJECT7 Tile_X5Y5_UO_OUT_TT_PROJECT0 Tile_X5Y5_UO_OUT_TT_PROJECT1
+ Tile_X5Y5_UO_OUT_TT_PROJECT2 Tile_X5Y5_UO_OUT_TT_PROJECT3 Tile_X5Y5_UO_OUT_TT_PROJECT4
+ Tile_X5Y5_UO_OUT_TT_PROJECT5 Tile_X5Y5_UO_OUT_TT_PROJECT6 Tile_X5Y5_UO_OUT_TT_PROJECT7
+ Tile_X5Y5_E_TT_IF/UserCLK Tile_X5Y4_E_TT_IF/UserCLK VGND VPWR Tile_X4Y5_LUT4AB/W1END[0]
+ Tile_X4Y5_LUT4AB/W1END[1] Tile_X4Y5_LUT4AB/W1END[2] Tile_X4Y5_LUT4AB/W1END[3] Tile_X4Y5_LUT4AB/W2MID[0]
+ Tile_X4Y5_LUT4AB/W2MID[1] Tile_X4Y5_LUT4AB/W2MID[2] Tile_X4Y5_LUT4AB/W2MID[3] Tile_X4Y5_LUT4AB/W2MID[4]
+ Tile_X4Y5_LUT4AB/W2MID[5] Tile_X4Y5_LUT4AB/W2MID[6] Tile_X4Y5_LUT4AB/W2MID[7] Tile_X4Y5_LUT4AB/W2END[0]
+ Tile_X4Y5_LUT4AB/W2END[1] Tile_X4Y5_LUT4AB/W2END[2] Tile_X4Y5_LUT4AB/W2END[3] Tile_X4Y5_LUT4AB/W2END[4]
+ Tile_X4Y5_LUT4AB/W2END[5] Tile_X4Y5_LUT4AB/W2END[6] Tile_X4Y5_LUT4AB/W2END[7] Tile_X4Y5_LUT4AB/W6END[0]
+ Tile_X4Y5_LUT4AB/W6END[10] Tile_X4Y5_LUT4AB/W6END[11] Tile_X4Y5_LUT4AB/W6END[1]
+ Tile_X4Y5_LUT4AB/W6END[2] Tile_X4Y5_LUT4AB/W6END[3] Tile_X4Y5_LUT4AB/W6END[4] Tile_X4Y5_LUT4AB/W6END[5]
+ Tile_X4Y5_LUT4AB/W6END[6] Tile_X4Y5_LUT4AB/W6END[7] Tile_X4Y5_LUT4AB/W6END[8] Tile_X4Y5_LUT4AB/W6END[9]
+ Tile_X4Y5_LUT4AB/WW4END[0] Tile_X4Y5_LUT4AB/WW4END[10] Tile_X4Y5_LUT4AB/WW4END[11]
+ Tile_X4Y5_LUT4AB/WW4END[12] Tile_X4Y5_LUT4AB/WW4END[13] Tile_X4Y5_LUT4AB/WW4END[14]
+ Tile_X4Y5_LUT4AB/WW4END[15] Tile_X4Y5_LUT4AB/WW4END[1] Tile_X4Y5_LUT4AB/WW4END[2]
+ Tile_X4Y5_LUT4AB/WW4END[3] Tile_X4Y5_LUT4AB/WW4END[4] Tile_X4Y5_LUT4AB/WW4END[5]
+ Tile_X4Y5_LUT4AB/WW4END[6] Tile_X4Y5_LUT4AB/WW4END[7] Tile_X4Y5_LUT4AB/WW4END[8]
+ Tile_X4Y5_LUT4AB/WW4END[9] E_TT_IF
XTile_X3Y7_LUT4AB Tile_X3Y8_LUT4AB/Co Tile_X3Y7_LUT4AB/Co Tile_X4Y7_LUT4AB/E1END[0]
+ Tile_X4Y7_LUT4AB/E1END[1] Tile_X4Y7_LUT4AB/E1END[2] Tile_X4Y7_LUT4AB/E1END[3] Tile_X3Y7_LUT4AB/E1END[0]
+ Tile_X3Y7_LUT4AB/E1END[1] Tile_X3Y7_LUT4AB/E1END[2] Tile_X3Y7_LUT4AB/E1END[3] Tile_X4Y7_LUT4AB/E2MID[0]
+ Tile_X4Y7_LUT4AB/E2MID[1] Tile_X4Y7_LUT4AB/E2MID[2] Tile_X4Y7_LUT4AB/E2MID[3] Tile_X4Y7_LUT4AB/E2MID[4]
+ Tile_X4Y7_LUT4AB/E2MID[5] Tile_X4Y7_LUT4AB/E2MID[6] Tile_X4Y7_LUT4AB/E2MID[7] Tile_X4Y7_LUT4AB/E2END[0]
+ Tile_X4Y7_LUT4AB/E2END[1] Tile_X4Y7_LUT4AB/E2END[2] Tile_X4Y7_LUT4AB/E2END[3] Tile_X4Y7_LUT4AB/E2END[4]
+ Tile_X4Y7_LUT4AB/E2END[5] Tile_X4Y7_LUT4AB/E2END[6] Tile_X4Y7_LUT4AB/E2END[7] Tile_X3Y7_LUT4AB/E2END[0]
+ Tile_X3Y7_LUT4AB/E2END[1] Tile_X3Y7_LUT4AB/E2END[2] Tile_X3Y7_LUT4AB/E2END[3] Tile_X3Y7_LUT4AB/E2END[4]
+ Tile_X3Y7_LUT4AB/E2END[5] Tile_X3Y7_LUT4AB/E2END[6] Tile_X3Y7_LUT4AB/E2END[7] Tile_X3Y7_LUT4AB/E2MID[0]
+ Tile_X3Y7_LUT4AB/E2MID[1] Tile_X3Y7_LUT4AB/E2MID[2] Tile_X3Y7_LUT4AB/E2MID[3] Tile_X3Y7_LUT4AB/E2MID[4]
+ Tile_X3Y7_LUT4AB/E2MID[5] Tile_X3Y7_LUT4AB/E2MID[6] Tile_X3Y7_LUT4AB/E2MID[7] Tile_X4Y7_LUT4AB/E6END[0]
+ Tile_X4Y7_LUT4AB/E6END[10] Tile_X4Y7_LUT4AB/E6END[11] Tile_X4Y7_LUT4AB/E6END[1]
+ Tile_X4Y7_LUT4AB/E6END[2] Tile_X4Y7_LUT4AB/E6END[3] Tile_X4Y7_LUT4AB/E6END[4] Tile_X4Y7_LUT4AB/E6END[5]
+ Tile_X4Y7_LUT4AB/E6END[6] Tile_X4Y7_LUT4AB/E6END[7] Tile_X4Y7_LUT4AB/E6END[8] Tile_X4Y7_LUT4AB/E6END[9]
+ Tile_X3Y7_LUT4AB/E6END[0] Tile_X3Y7_LUT4AB/E6END[10] Tile_X3Y7_LUT4AB/E6END[11]
+ Tile_X3Y7_LUT4AB/E6END[1] Tile_X3Y7_LUT4AB/E6END[2] Tile_X3Y7_LUT4AB/E6END[3] Tile_X3Y7_LUT4AB/E6END[4]
+ Tile_X3Y7_LUT4AB/E6END[5] Tile_X3Y7_LUT4AB/E6END[6] Tile_X3Y7_LUT4AB/E6END[7] Tile_X3Y7_LUT4AB/E6END[8]
+ Tile_X3Y7_LUT4AB/E6END[9] Tile_X4Y7_LUT4AB/EE4END[0] Tile_X4Y7_LUT4AB/EE4END[10]
+ Tile_X4Y7_LUT4AB/EE4END[11] Tile_X4Y7_LUT4AB/EE4END[12] Tile_X4Y7_LUT4AB/EE4END[13]
+ Tile_X4Y7_LUT4AB/EE4END[14] Tile_X4Y7_LUT4AB/EE4END[15] Tile_X4Y7_LUT4AB/EE4END[1]
+ Tile_X4Y7_LUT4AB/EE4END[2] Tile_X4Y7_LUT4AB/EE4END[3] Tile_X4Y7_LUT4AB/EE4END[4]
+ Tile_X4Y7_LUT4AB/EE4END[5] Tile_X4Y7_LUT4AB/EE4END[6] Tile_X4Y7_LUT4AB/EE4END[7]
+ Tile_X4Y7_LUT4AB/EE4END[8] Tile_X4Y7_LUT4AB/EE4END[9] Tile_X3Y7_LUT4AB/EE4END[0]
+ Tile_X3Y7_LUT4AB/EE4END[10] Tile_X3Y7_LUT4AB/EE4END[11] Tile_X3Y7_LUT4AB/EE4END[12]
+ Tile_X3Y7_LUT4AB/EE4END[13] Tile_X3Y7_LUT4AB/EE4END[14] Tile_X3Y7_LUT4AB/EE4END[15]
+ Tile_X3Y7_LUT4AB/EE4END[1] Tile_X3Y7_LUT4AB/EE4END[2] Tile_X3Y7_LUT4AB/EE4END[3]
+ Tile_X3Y7_LUT4AB/EE4END[4] Tile_X3Y7_LUT4AB/EE4END[5] Tile_X3Y7_LUT4AB/EE4END[6]
+ Tile_X3Y7_LUT4AB/EE4END[7] Tile_X3Y7_LUT4AB/EE4END[8] Tile_X3Y7_LUT4AB/EE4END[9]
+ Tile_X3Y7_LUT4AB/FrameData[0] Tile_X3Y7_LUT4AB/FrameData[10] Tile_X3Y7_LUT4AB/FrameData[11]
+ Tile_X3Y7_LUT4AB/FrameData[12] Tile_X3Y7_LUT4AB/FrameData[13] Tile_X3Y7_LUT4AB/FrameData[14]
+ Tile_X3Y7_LUT4AB/FrameData[15] Tile_X3Y7_LUT4AB/FrameData[16] Tile_X3Y7_LUT4AB/FrameData[17]
+ Tile_X3Y7_LUT4AB/FrameData[18] Tile_X3Y7_LUT4AB/FrameData[19] Tile_X3Y7_LUT4AB/FrameData[1]
+ Tile_X3Y7_LUT4AB/FrameData[20] Tile_X3Y7_LUT4AB/FrameData[21] Tile_X3Y7_LUT4AB/FrameData[22]
+ Tile_X3Y7_LUT4AB/FrameData[23] Tile_X3Y7_LUT4AB/FrameData[24] Tile_X3Y7_LUT4AB/FrameData[25]
+ Tile_X3Y7_LUT4AB/FrameData[26] Tile_X3Y7_LUT4AB/FrameData[27] Tile_X3Y7_LUT4AB/FrameData[28]
+ Tile_X3Y7_LUT4AB/FrameData[29] Tile_X3Y7_LUT4AB/FrameData[2] Tile_X3Y7_LUT4AB/FrameData[30]
+ Tile_X3Y7_LUT4AB/FrameData[31] Tile_X3Y7_LUT4AB/FrameData[3] Tile_X3Y7_LUT4AB/FrameData[4]
+ Tile_X3Y7_LUT4AB/FrameData[5] Tile_X3Y7_LUT4AB/FrameData[6] Tile_X3Y7_LUT4AB/FrameData[7]
+ Tile_X3Y7_LUT4AB/FrameData[8] Tile_X3Y7_LUT4AB/FrameData[9] Tile_X4Y7_LUT4AB/FrameData[0]
+ Tile_X4Y7_LUT4AB/FrameData[10] Tile_X4Y7_LUT4AB/FrameData[11] Tile_X4Y7_LUT4AB/FrameData[12]
+ Tile_X4Y7_LUT4AB/FrameData[13] Tile_X4Y7_LUT4AB/FrameData[14] Tile_X4Y7_LUT4AB/FrameData[15]
+ Tile_X4Y7_LUT4AB/FrameData[16] Tile_X4Y7_LUT4AB/FrameData[17] Tile_X4Y7_LUT4AB/FrameData[18]
+ Tile_X4Y7_LUT4AB/FrameData[19] Tile_X4Y7_LUT4AB/FrameData[1] Tile_X4Y7_LUT4AB/FrameData[20]
+ Tile_X4Y7_LUT4AB/FrameData[21] Tile_X4Y7_LUT4AB/FrameData[22] Tile_X4Y7_LUT4AB/FrameData[23]
+ Tile_X4Y7_LUT4AB/FrameData[24] Tile_X4Y7_LUT4AB/FrameData[25] Tile_X4Y7_LUT4AB/FrameData[26]
+ Tile_X4Y7_LUT4AB/FrameData[27] Tile_X4Y7_LUT4AB/FrameData[28] Tile_X4Y7_LUT4AB/FrameData[29]
+ Tile_X4Y7_LUT4AB/FrameData[2] Tile_X4Y7_LUT4AB/FrameData[30] Tile_X4Y7_LUT4AB/FrameData[31]
+ Tile_X4Y7_LUT4AB/FrameData[3] Tile_X4Y7_LUT4AB/FrameData[4] Tile_X4Y7_LUT4AB/FrameData[5]
+ Tile_X4Y7_LUT4AB/FrameData[6] Tile_X4Y7_LUT4AB/FrameData[7] Tile_X4Y7_LUT4AB/FrameData[8]
+ Tile_X4Y7_LUT4AB/FrameData[9] Tile_X3Y7_LUT4AB/FrameStrobe[0] Tile_X3Y7_LUT4AB/FrameStrobe[10]
+ Tile_X3Y7_LUT4AB/FrameStrobe[11] Tile_X3Y7_LUT4AB/FrameStrobe[12] Tile_X3Y7_LUT4AB/FrameStrobe[13]
+ Tile_X3Y7_LUT4AB/FrameStrobe[14] Tile_X3Y7_LUT4AB/FrameStrobe[15] Tile_X3Y7_LUT4AB/FrameStrobe[16]
+ Tile_X3Y7_LUT4AB/FrameStrobe[17] Tile_X3Y7_LUT4AB/FrameStrobe[18] Tile_X3Y7_LUT4AB/FrameStrobe[19]
+ Tile_X3Y7_LUT4AB/FrameStrobe[1] Tile_X3Y7_LUT4AB/FrameStrobe[2] Tile_X3Y7_LUT4AB/FrameStrobe[3]
+ Tile_X3Y7_LUT4AB/FrameStrobe[4] Tile_X3Y7_LUT4AB/FrameStrobe[5] Tile_X3Y7_LUT4AB/FrameStrobe[6]
+ Tile_X3Y7_LUT4AB/FrameStrobe[7] Tile_X3Y7_LUT4AB/FrameStrobe[8] Tile_X3Y7_LUT4AB/FrameStrobe[9]
+ Tile_X3Y6_LUT4AB/FrameStrobe[0] Tile_X3Y6_LUT4AB/FrameStrobe[10] Tile_X3Y6_LUT4AB/FrameStrobe[11]
+ Tile_X3Y6_LUT4AB/FrameStrobe[12] Tile_X3Y6_LUT4AB/FrameStrobe[13] Tile_X3Y6_LUT4AB/FrameStrobe[14]
+ Tile_X3Y6_LUT4AB/FrameStrobe[15] Tile_X3Y6_LUT4AB/FrameStrobe[16] Tile_X3Y6_LUT4AB/FrameStrobe[17]
+ Tile_X3Y6_LUT4AB/FrameStrobe[18] Tile_X3Y6_LUT4AB/FrameStrobe[19] Tile_X3Y6_LUT4AB/FrameStrobe[1]
+ Tile_X3Y6_LUT4AB/FrameStrobe[2] Tile_X3Y6_LUT4AB/FrameStrobe[3] Tile_X3Y6_LUT4AB/FrameStrobe[4]
+ Tile_X3Y6_LUT4AB/FrameStrobe[5] Tile_X3Y6_LUT4AB/FrameStrobe[6] Tile_X3Y6_LUT4AB/FrameStrobe[7]
+ Tile_X3Y6_LUT4AB/FrameStrobe[8] Tile_X3Y6_LUT4AB/FrameStrobe[9] Tile_X3Y7_LUT4AB/N1BEG[0]
+ Tile_X3Y7_LUT4AB/N1BEG[1] Tile_X3Y7_LUT4AB/N1BEG[2] Tile_X3Y7_LUT4AB/N1BEG[3] Tile_X3Y8_LUT4AB/N1BEG[0]
+ Tile_X3Y8_LUT4AB/N1BEG[1] Tile_X3Y8_LUT4AB/N1BEG[2] Tile_X3Y8_LUT4AB/N1BEG[3] Tile_X3Y7_LUT4AB/N2BEG[0]
+ Tile_X3Y7_LUT4AB/N2BEG[1] Tile_X3Y7_LUT4AB/N2BEG[2] Tile_X3Y7_LUT4AB/N2BEG[3] Tile_X3Y7_LUT4AB/N2BEG[4]
+ Tile_X3Y7_LUT4AB/N2BEG[5] Tile_X3Y7_LUT4AB/N2BEG[6] Tile_X3Y7_LUT4AB/N2BEG[7] Tile_X3Y6_LUT4AB/N2END[0]
+ Tile_X3Y6_LUT4AB/N2END[1] Tile_X3Y6_LUT4AB/N2END[2] Tile_X3Y6_LUT4AB/N2END[3] Tile_X3Y6_LUT4AB/N2END[4]
+ Tile_X3Y6_LUT4AB/N2END[5] Tile_X3Y6_LUT4AB/N2END[6] Tile_X3Y6_LUT4AB/N2END[7] Tile_X3Y7_LUT4AB/N2END[0]
+ Tile_X3Y7_LUT4AB/N2END[1] Tile_X3Y7_LUT4AB/N2END[2] Tile_X3Y7_LUT4AB/N2END[3] Tile_X3Y7_LUT4AB/N2END[4]
+ Tile_X3Y7_LUT4AB/N2END[5] Tile_X3Y7_LUT4AB/N2END[6] Tile_X3Y7_LUT4AB/N2END[7] Tile_X3Y8_LUT4AB/N2BEG[0]
+ Tile_X3Y8_LUT4AB/N2BEG[1] Tile_X3Y8_LUT4AB/N2BEG[2] Tile_X3Y8_LUT4AB/N2BEG[3] Tile_X3Y8_LUT4AB/N2BEG[4]
+ Tile_X3Y8_LUT4AB/N2BEG[5] Tile_X3Y8_LUT4AB/N2BEG[6] Tile_X3Y8_LUT4AB/N2BEG[7] Tile_X3Y7_LUT4AB/N4BEG[0]
+ Tile_X3Y7_LUT4AB/N4BEG[10] Tile_X3Y7_LUT4AB/N4BEG[11] Tile_X3Y7_LUT4AB/N4BEG[12]
+ Tile_X3Y7_LUT4AB/N4BEG[13] Tile_X3Y7_LUT4AB/N4BEG[14] Tile_X3Y7_LUT4AB/N4BEG[15]
+ Tile_X3Y7_LUT4AB/N4BEG[1] Tile_X3Y7_LUT4AB/N4BEG[2] Tile_X3Y7_LUT4AB/N4BEG[3] Tile_X3Y7_LUT4AB/N4BEG[4]
+ Tile_X3Y7_LUT4AB/N4BEG[5] Tile_X3Y7_LUT4AB/N4BEG[6] Tile_X3Y7_LUT4AB/N4BEG[7] Tile_X3Y7_LUT4AB/N4BEG[8]
+ Tile_X3Y7_LUT4AB/N4BEG[9] Tile_X3Y8_LUT4AB/N4BEG[0] Tile_X3Y8_LUT4AB/N4BEG[10] Tile_X3Y8_LUT4AB/N4BEG[11]
+ Tile_X3Y8_LUT4AB/N4BEG[12] Tile_X3Y8_LUT4AB/N4BEG[13] Tile_X3Y8_LUT4AB/N4BEG[14]
+ Tile_X3Y8_LUT4AB/N4BEG[15] Tile_X3Y8_LUT4AB/N4BEG[1] Tile_X3Y8_LUT4AB/N4BEG[2] Tile_X3Y8_LUT4AB/N4BEG[3]
+ Tile_X3Y8_LUT4AB/N4BEG[4] Tile_X3Y8_LUT4AB/N4BEG[5] Tile_X3Y8_LUT4AB/N4BEG[6] Tile_X3Y8_LUT4AB/N4BEG[7]
+ Tile_X3Y8_LUT4AB/N4BEG[8] Tile_X3Y8_LUT4AB/N4BEG[9] Tile_X3Y7_LUT4AB/NN4BEG[0] Tile_X3Y7_LUT4AB/NN4BEG[10]
+ Tile_X3Y7_LUT4AB/NN4BEG[11] Tile_X3Y7_LUT4AB/NN4BEG[12] Tile_X3Y7_LUT4AB/NN4BEG[13]
+ Tile_X3Y7_LUT4AB/NN4BEG[14] Tile_X3Y7_LUT4AB/NN4BEG[15] Tile_X3Y7_LUT4AB/NN4BEG[1]
+ Tile_X3Y7_LUT4AB/NN4BEG[2] Tile_X3Y7_LUT4AB/NN4BEG[3] Tile_X3Y7_LUT4AB/NN4BEG[4]
+ Tile_X3Y7_LUT4AB/NN4BEG[5] Tile_X3Y7_LUT4AB/NN4BEG[6] Tile_X3Y7_LUT4AB/NN4BEG[7]
+ Tile_X3Y7_LUT4AB/NN4BEG[8] Tile_X3Y7_LUT4AB/NN4BEG[9] Tile_X3Y8_LUT4AB/NN4BEG[0]
+ Tile_X3Y8_LUT4AB/NN4BEG[10] Tile_X3Y8_LUT4AB/NN4BEG[11] Tile_X3Y8_LUT4AB/NN4BEG[12]
+ Tile_X3Y8_LUT4AB/NN4BEG[13] Tile_X3Y8_LUT4AB/NN4BEG[14] Tile_X3Y8_LUT4AB/NN4BEG[15]
+ Tile_X3Y8_LUT4AB/NN4BEG[1] Tile_X3Y8_LUT4AB/NN4BEG[2] Tile_X3Y8_LUT4AB/NN4BEG[3]
+ Tile_X3Y8_LUT4AB/NN4BEG[4] Tile_X3Y8_LUT4AB/NN4BEG[5] Tile_X3Y8_LUT4AB/NN4BEG[6]
+ Tile_X3Y8_LUT4AB/NN4BEG[7] Tile_X3Y8_LUT4AB/NN4BEG[8] Tile_X3Y8_LUT4AB/NN4BEG[9]
+ Tile_X3Y8_LUT4AB/S1END[0] Tile_X3Y8_LUT4AB/S1END[1] Tile_X3Y8_LUT4AB/S1END[2] Tile_X3Y8_LUT4AB/S1END[3]
+ Tile_X3Y7_LUT4AB/S1END[0] Tile_X3Y7_LUT4AB/S1END[1] Tile_X3Y7_LUT4AB/S1END[2] Tile_X3Y7_LUT4AB/S1END[3]
+ Tile_X3Y8_LUT4AB/S2MID[0] Tile_X3Y8_LUT4AB/S2MID[1] Tile_X3Y8_LUT4AB/S2MID[2] Tile_X3Y8_LUT4AB/S2MID[3]
+ Tile_X3Y8_LUT4AB/S2MID[4] Tile_X3Y8_LUT4AB/S2MID[5] Tile_X3Y8_LUT4AB/S2MID[6] Tile_X3Y8_LUT4AB/S2MID[7]
+ Tile_X3Y8_LUT4AB/S2END[0] Tile_X3Y8_LUT4AB/S2END[1] Tile_X3Y8_LUT4AB/S2END[2] Tile_X3Y8_LUT4AB/S2END[3]
+ Tile_X3Y8_LUT4AB/S2END[4] Tile_X3Y8_LUT4AB/S2END[5] Tile_X3Y8_LUT4AB/S2END[6] Tile_X3Y8_LUT4AB/S2END[7]
+ Tile_X3Y7_LUT4AB/S2END[0] Tile_X3Y7_LUT4AB/S2END[1] Tile_X3Y7_LUT4AB/S2END[2] Tile_X3Y7_LUT4AB/S2END[3]
+ Tile_X3Y7_LUT4AB/S2END[4] Tile_X3Y7_LUT4AB/S2END[5] Tile_X3Y7_LUT4AB/S2END[6] Tile_X3Y7_LUT4AB/S2END[7]
+ Tile_X3Y7_LUT4AB/S2MID[0] Tile_X3Y7_LUT4AB/S2MID[1] Tile_X3Y7_LUT4AB/S2MID[2] Tile_X3Y7_LUT4AB/S2MID[3]
+ Tile_X3Y7_LUT4AB/S2MID[4] Tile_X3Y7_LUT4AB/S2MID[5] Tile_X3Y7_LUT4AB/S2MID[6] Tile_X3Y7_LUT4AB/S2MID[7]
+ Tile_X3Y8_LUT4AB/S4END[0] Tile_X3Y8_LUT4AB/S4END[10] Tile_X3Y8_LUT4AB/S4END[11]
+ Tile_X3Y8_LUT4AB/S4END[12] Tile_X3Y8_LUT4AB/S4END[13] Tile_X3Y8_LUT4AB/S4END[14]
+ Tile_X3Y8_LUT4AB/S4END[15] Tile_X3Y8_LUT4AB/S4END[1] Tile_X3Y8_LUT4AB/S4END[2] Tile_X3Y8_LUT4AB/S4END[3]
+ Tile_X3Y8_LUT4AB/S4END[4] Tile_X3Y8_LUT4AB/S4END[5] Tile_X3Y8_LUT4AB/S4END[6] Tile_X3Y8_LUT4AB/S4END[7]
+ Tile_X3Y8_LUT4AB/S4END[8] Tile_X3Y8_LUT4AB/S4END[9] Tile_X3Y7_LUT4AB/S4END[0] Tile_X3Y7_LUT4AB/S4END[10]
+ Tile_X3Y7_LUT4AB/S4END[11] Tile_X3Y7_LUT4AB/S4END[12] Tile_X3Y7_LUT4AB/S4END[13]
+ Tile_X3Y7_LUT4AB/S4END[14] Tile_X3Y7_LUT4AB/S4END[15] Tile_X3Y7_LUT4AB/S4END[1]
+ Tile_X3Y7_LUT4AB/S4END[2] Tile_X3Y7_LUT4AB/S4END[3] Tile_X3Y7_LUT4AB/S4END[4] Tile_X3Y7_LUT4AB/S4END[5]
+ Tile_X3Y7_LUT4AB/S4END[6] Tile_X3Y7_LUT4AB/S4END[7] Tile_X3Y7_LUT4AB/S4END[8] Tile_X3Y7_LUT4AB/S4END[9]
+ Tile_X3Y8_LUT4AB/SS4END[0] Tile_X3Y8_LUT4AB/SS4END[10] Tile_X3Y8_LUT4AB/SS4END[11]
+ Tile_X3Y8_LUT4AB/SS4END[12] Tile_X3Y8_LUT4AB/SS4END[13] Tile_X3Y8_LUT4AB/SS4END[14]
+ Tile_X3Y8_LUT4AB/SS4END[15] Tile_X3Y8_LUT4AB/SS4END[1] Tile_X3Y8_LUT4AB/SS4END[2]
+ Tile_X3Y8_LUT4AB/SS4END[3] Tile_X3Y8_LUT4AB/SS4END[4] Tile_X3Y8_LUT4AB/SS4END[5]
+ Tile_X3Y8_LUT4AB/SS4END[6] Tile_X3Y8_LUT4AB/SS4END[7] Tile_X3Y8_LUT4AB/SS4END[8]
+ Tile_X3Y8_LUT4AB/SS4END[9] Tile_X3Y7_LUT4AB/SS4END[0] Tile_X3Y7_LUT4AB/SS4END[10]
+ Tile_X3Y7_LUT4AB/SS4END[11] Tile_X3Y7_LUT4AB/SS4END[12] Tile_X3Y7_LUT4AB/SS4END[13]
+ Tile_X3Y7_LUT4AB/SS4END[14] Tile_X3Y7_LUT4AB/SS4END[15] Tile_X3Y7_LUT4AB/SS4END[1]
+ Tile_X3Y7_LUT4AB/SS4END[2] Tile_X3Y7_LUT4AB/SS4END[3] Tile_X3Y7_LUT4AB/SS4END[4]
+ Tile_X3Y7_LUT4AB/SS4END[5] Tile_X3Y7_LUT4AB/SS4END[6] Tile_X3Y7_LUT4AB/SS4END[7]
+ Tile_X3Y7_LUT4AB/SS4END[8] Tile_X3Y7_LUT4AB/SS4END[9] Tile_X3Y7_LUT4AB/UserCLK Tile_X3Y6_LUT4AB/UserCLK
+ VGND VPWR Tile_X3Y7_LUT4AB/W1BEG[0] Tile_X3Y7_LUT4AB/W1BEG[1] Tile_X3Y7_LUT4AB/W1BEG[2]
+ Tile_X3Y7_LUT4AB/W1BEG[3] Tile_X4Y7_LUT4AB/W1BEG[0] Tile_X4Y7_LUT4AB/W1BEG[1] Tile_X4Y7_LUT4AB/W1BEG[2]
+ Tile_X4Y7_LUT4AB/W1BEG[3] Tile_X3Y7_LUT4AB/W2BEG[0] Tile_X3Y7_LUT4AB/W2BEG[1] Tile_X3Y7_LUT4AB/W2BEG[2]
+ Tile_X3Y7_LUT4AB/W2BEG[3] Tile_X3Y7_LUT4AB/W2BEG[4] Tile_X3Y7_LUT4AB/W2BEG[5] Tile_X3Y7_LUT4AB/W2BEG[6]
+ Tile_X3Y7_LUT4AB/W2BEG[7] Tile_X2Y7_LUT4AB/W2END[0] Tile_X2Y7_LUT4AB/W2END[1] Tile_X2Y7_LUT4AB/W2END[2]
+ Tile_X2Y7_LUT4AB/W2END[3] Tile_X2Y7_LUT4AB/W2END[4] Tile_X2Y7_LUT4AB/W2END[5] Tile_X2Y7_LUT4AB/W2END[6]
+ Tile_X2Y7_LUT4AB/W2END[7] Tile_X3Y7_LUT4AB/W2END[0] Tile_X3Y7_LUT4AB/W2END[1] Tile_X3Y7_LUT4AB/W2END[2]
+ Tile_X3Y7_LUT4AB/W2END[3] Tile_X3Y7_LUT4AB/W2END[4] Tile_X3Y7_LUT4AB/W2END[5] Tile_X3Y7_LUT4AB/W2END[6]
+ Tile_X3Y7_LUT4AB/W2END[7] Tile_X4Y7_LUT4AB/W2BEG[0] Tile_X4Y7_LUT4AB/W2BEG[1] Tile_X4Y7_LUT4AB/W2BEG[2]
+ Tile_X4Y7_LUT4AB/W2BEG[3] Tile_X4Y7_LUT4AB/W2BEG[4] Tile_X4Y7_LUT4AB/W2BEG[5] Tile_X4Y7_LUT4AB/W2BEG[6]
+ Tile_X4Y7_LUT4AB/W2BEG[7] Tile_X3Y7_LUT4AB/W6BEG[0] Tile_X3Y7_LUT4AB/W6BEG[10] Tile_X3Y7_LUT4AB/W6BEG[11]
+ Tile_X3Y7_LUT4AB/W6BEG[1] Tile_X3Y7_LUT4AB/W6BEG[2] Tile_X3Y7_LUT4AB/W6BEG[3] Tile_X3Y7_LUT4AB/W6BEG[4]
+ Tile_X3Y7_LUT4AB/W6BEG[5] Tile_X3Y7_LUT4AB/W6BEG[6] Tile_X3Y7_LUT4AB/W6BEG[7] Tile_X3Y7_LUT4AB/W6BEG[8]
+ Tile_X3Y7_LUT4AB/W6BEG[9] Tile_X4Y7_LUT4AB/W6BEG[0] Tile_X4Y7_LUT4AB/W6BEG[10] Tile_X4Y7_LUT4AB/W6BEG[11]
+ Tile_X4Y7_LUT4AB/W6BEG[1] Tile_X4Y7_LUT4AB/W6BEG[2] Tile_X4Y7_LUT4AB/W6BEG[3] Tile_X4Y7_LUT4AB/W6BEG[4]
+ Tile_X4Y7_LUT4AB/W6BEG[5] Tile_X4Y7_LUT4AB/W6BEG[6] Tile_X4Y7_LUT4AB/W6BEG[7] Tile_X4Y7_LUT4AB/W6BEG[8]
+ Tile_X4Y7_LUT4AB/W6BEG[9] Tile_X3Y7_LUT4AB/WW4BEG[0] Tile_X3Y7_LUT4AB/WW4BEG[10]
+ Tile_X3Y7_LUT4AB/WW4BEG[11] Tile_X3Y7_LUT4AB/WW4BEG[12] Tile_X3Y7_LUT4AB/WW4BEG[13]
+ Tile_X3Y7_LUT4AB/WW4BEG[14] Tile_X3Y7_LUT4AB/WW4BEG[15] Tile_X3Y7_LUT4AB/WW4BEG[1]
+ Tile_X3Y7_LUT4AB/WW4BEG[2] Tile_X3Y7_LUT4AB/WW4BEG[3] Tile_X3Y7_LUT4AB/WW4BEG[4]
+ Tile_X3Y7_LUT4AB/WW4BEG[5] Tile_X3Y7_LUT4AB/WW4BEG[6] Tile_X3Y7_LUT4AB/WW4BEG[7]
+ Tile_X3Y7_LUT4AB/WW4BEG[8] Tile_X3Y7_LUT4AB/WW4BEG[9] Tile_X4Y7_LUT4AB/WW4BEG[0]
+ Tile_X4Y7_LUT4AB/WW4BEG[10] Tile_X4Y7_LUT4AB/WW4BEG[11] Tile_X4Y7_LUT4AB/WW4BEG[12]
+ Tile_X4Y7_LUT4AB/WW4BEG[13] Tile_X4Y7_LUT4AB/WW4BEG[14] Tile_X4Y7_LUT4AB/WW4BEG[15]
+ Tile_X4Y7_LUT4AB/WW4BEG[1] Tile_X4Y7_LUT4AB/WW4BEG[2] Tile_X4Y7_LUT4AB/WW4BEG[3]
+ Tile_X4Y7_LUT4AB/WW4BEG[4] Tile_X4Y7_LUT4AB/WW4BEG[5] Tile_X4Y7_LUT4AB/WW4BEG[6]
+ Tile_X4Y7_LUT4AB/WW4BEG[7] Tile_X4Y7_LUT4AB/WW4BEG[8] Tile_X4Y7_LUT4AB/WW4BEG[9]
+ LUT4AB
XTile_X1Y4_LUT4AB Tile_X1Y5_LUT4AB/Co Tile_X1Y4_LUT4AB/Co Tile_X2Y4_LUT4AB/E1END[0]
+ Tile_X2Y4_LUT4AB/E1END[1] Tile_X2Y4_LUT4AB/E1END[2] Tile_X2Y4_LUT4AB/E1END[3] Tile_X1Y4_LUT4AB/E1END[0]
+ Tile_X1Y4_LUT4AB/E1END[1] Tile_X1Y4_LUT4AB/E1END[2] Tile_X1Y4_LUT4AB/E1END[3] Tile_X2Y4_LUT4AB/E2MID[0]
+ Tile_X2Y4_LUT4AB/E2MID[1] Tile_X2Y4_LUT4AB/E2MID[2] Tile_X2Y4_LUT4AB/E2MID[3] Tile_X2Y4_LUT4AB/E2MID[4]
+ Tile_X2Y4_LUT4AB/E2MID[5] Tile_X2Y4_LUT4AB/E2MID[6] Tile_X2Y4_LUT4AB/E2MID[7] Tile_X2Y4_LUT4AB/E2END[0]
+ Tile_X2Y4_LUT4AB/E2END[1] Tile_X2Y4_LUT4AB/E2END[2] Tile_X2Y4_LUT4AB/E2END[3] Tile_X2Y4_LUT4AB/E2END[4]
+ Tile_X2Y4_LUT4AB/E2END[5] Tile_X2Y4_LUT4AB/E2END[6] Tile_X2Y4_LUT4AB/E2END[7] Tile_X1Y4_LUT4AB/E2END[0]
+ Tile_X1Y4_LUT4AB/E2END[1] Tile_X1Y4_LUT4AB/E2END[2] Tile_X1Y4_LUT4AB/E2END[3] Tile_X1Y4_LUT4AB/E2END[4]
+ Tile_X1Y4_LUT4AB/E2END[5] Tile_X1Y4_LUT4AB/E2END[6] Tile_X1Y4_LUT4AB/E2END[7] Tile_X1Y4_LUT4AB/E2MID[0]
+ Tile_X1Y4_LUT4AB/E2MID[1] Tile_X1Y4_LUT4AB/E2MID[2] Tile_X1Y4_LUT4AB/E2MID[3] Tile_X1Y4_LUT4AB/E2MID[4]
+ Tile_X1Y4_LUT4AB/E2MID[5] Tile_X1Y4_LUT4AB/E2MID[6] Tile_X1Y4_LUT4AB/E2MID[7] Tile_X2Y4_LUT4AB/E6END[0]
+ Tile_X2Y4_LUT4AB/E6END[10] Tile_X2Y4_LUT4AB/E6END[11] Tile_X2Y4_LUT4AB/E6END[1]
+ Tile_X2Y4_LUT4AB/E6END[2] Tile_X2Y4_LUT4AB/E6END[3] Tile_X2Y4_LUT4AB/E6END[4] Tile_X2Y4_LUT4AB/E6END[5]
+ Tile_X2Y4_LUT4AB/E6END[6] Tile_X2Y4_LUT4AB/E6END[7] Tile_X2Y4_LUT4AB/E6END[8] Tile_X2Y4_LUT4AB/E6END[9]
+ Tile_X1Y4_LUT4AB/E6END[0] Tile_X1Y4_LUT4AB/E6END[10] Tile_X1Y4_LUT4AB/E6END[11]
+ Tile_X1Y4_LUT4AB/E6END[1] Tile_X1Y4_LUT4AB/E6END[2] Tile_X1Y4_LUT4AB/E6END[3] Tile_X1Y4_LUT4AB/E6END[4]
+ Tile_X1Y4_LUT4AB/E6END[5] Tile_X1Y4_LUT4AB/E6END[6] Tile_X1Y4_LUT4AB/E6END[7] Tile_X1Y4_LUT4AB/E6END[8]
+ Tile_X1Y4_LUT4AB/E6END[9] Tile_X2Y4_LUT4AB/EE4END[0] Tile_X2Y4_LUT4AB/EE4END[10]
+ Tile_X2Y4_LUT4AB/EE4END[11] Tile_X2Y4_LUT4AB/EE4END[12] Tile_X2Y4_LUT4AB/EE4END[13]
+ Tile_X2Y4_LUT4AB/EE4END[14] Tile_X2Y4_LUT4AB/EE4END[15] Tile_X2Y4_LUT4AB/EE4END[1]
+ Tile_X2Y4_LUT4AB/EE4END[2] Tile_X2Y4_LUT4AB/EE4END[3] Tile_X2Y4_LUT4AB/EE4END[4]
+ Tile_X2Y4_LUT4AB/EE4END[5] Tile_X2Y4_LUT4AB/EE4END[6] Tile_X2Y4_LUT4AB/EE4END[7]
+ Tile_X2Y4_LUT4AB/EE4END[8] Tile_X2Y4_LUT4AB/EE4END[9] Tile_X1Y4_LUT4AB/EE4END[0]
+ Tile_X1Y4_LUT4AB/EE4END[10] Tile_X1Y4_LUT4AB/EE4END[11] Tile_X1Y4_LUT4AB/EE4END[12]
+ Tile_X1Y4_LUT4AB/EE4END[13] Tile_X1Y4_LUT4AB/EE4END[14] Tile_X1Y4_LUT4AB/EE4END[15]
+ Tile_X1Y4_LUT4AB/EE4END[1] Tile_X1Y4_LUT4AB/EE4END[2] Tile_X1Y4_LUT4AB/EE4END[3]
+ Tile_X1Y4_LUT4AB/EE4END[4] Tile_X1Y4_LUT4AB/EE4END[5] Tile_X1Y4_LUT4AB/EE4END[6]
+ Tile_X1Y4_LUT4AB/EE4END[7] Tile_X1Y4_LUT4AB/EE4END[8] Tile_X1Y4_LUT4AB/EE4END[9]
+ Tile_X1Y4_LUT4AB/FrameData[0] Tile_X1Y4_LUT4AB/FrameData[10] Tile_X1Y4_LUT4AB/FrameData[11]
+ Tile_X1Y4_LUT4AB/FrameData[12] Tile_X1Y4_LUT4AB/FrameData[13] Tile_X1Y4_LUT4AB/FrameData[14]
+ Tile_X1Y4_LUT4AB/FrameData[15] Tile_X1Y4_LUT4AB/FrameData[16] Tile_X1Y4_LUT4AB/FrameData[17]
+ Tile_X1Y4_LUT4AB/FrameData[18] Tile_X1Y4_LUT4AB/FrameData[19] Tile_X1Y4_LUT4AB/FrameData[1]
+ Tile_X1Y4_LUT4AB/FrameData[20] Tile_X1Y4_LUT4AB/FrameData[21] Tile_X1Y4_LUT4AB/FrameData[22]
+ Tile_X1Y4_LUT4AB/FrameData[23] Tile_X1Y4_LUT4AB/FrameData[24] Tile_X1Y4_LUT4AB/FrameData[25]
+ Tile_X1Y4_LUT4AB/FrameData[26] Tile_X1Y4_LUT4AB/FrameData[27] Tile_X1Y4_LUT4AB/FrameData[28]
+ Tile_X1Y4_LUT4AB/FrameData[29] Tile_X1Y4_LUT4AB/FrameData[2] Tile_X1Y4_LUT4AB/FrameData[30]
+ Tile_X1Y4_LUT4AB/FrameData[31] Tile_X1Y4_LUT4AB/FrameData[3] Tile_X1Y4_LUT4AB/FrameData[4]
+ Tile_X1Y4_LUT4AB/FrameData[5] Tile_X1Y4_LUT4AB/FrameData[6] Tile_X1Y4_LUT4AB/FrameData[7]
+ Tile_X1Y4_LUT4AB/FrameData[8] Tile_X1Y4_LUT4AB/FrameData[9] Tile_X2Y4_LUT4AB/FrameData[0]
+ Tile_X2Y4_LUT4AB/FrameData[10] Tile_X2Y4_LUT4AB/FrameData[11] Tile_X2Y4_LUT4AB/FrameData[12]
+ Tile_X2Y4_LUT4AB/FrameData[13] Tile_X2Y4_LUT4AB/FrameData[14] Tile_X2Y4_LUT4AB/FrameData[15]
+ Tile_X2Y4_LUT4AB/FrameData[16] Tile_X2Y4_LUT4AB/FrameData[17] Tile_X2Y4_LUT4AB/FrameData[18]
+ Tile_X2Y4_LUT4AB/FrameData[19] Tile_X2Y4_LUT4AB/FrameData[1] Tile_X2Y4_LUT4AB/FrameData[20]
+ Tile_X2Y4_LUT4AB/FrameData[21] Tile_X2Y4_LUT4AB/FrameData[22] Tile_X2Y4_LUT4AB/FrameData[23]
+ Tile_X2Y4_LUT4AB/FrameData[24] Tile_X2Y4_LUT4AB/FrameData[25] Tile_X2Y4_LUT4AB/FrameData[26]
+ Tile_X2Y4_LUT4AB/FrameData[27] Tile_X2Y4_LUT4AB/FrameData[28] Tile_X2Y4_LUT4AB/FrameData[29]
+ Tile_X2Y4_LUT4AB/FrameData[2] Tile_X2Y4_LUT4AB/FrameData[30] Tile_X2Y4_LUT4AB/FrameData[31]
+ Tile_X2Y4_LUT4AB/FrameData[3] Tile_X2Y4_LUT4AB/FrameData[4] Tile_X2Y4_LUT4AB/FrameData[5]
+ Tile_X2Y4_LUT4AB/FrameData[6] Tile_X2Y4_LUT4AB/FrameData[7] Tile_X2Y4_LUT4AB/FrameData[8]
+ Tile_X2Y4_LUT4AB/FrameData[9] Tile_X1Y4_LUT4AB/FrameStrobe[0] Tile_X1Y4_LUT4AB/FrameStrobe[10]
+ Tile_X1Y4_LUT4AB/FrameStrobe[11] Tile_X1Y4_LUT4AB/FrameStrobe[12] Tile_X1Y4_LUT4AB/FrameStrobe[13]
+ Tile_X1Y4_LUT4AB/FrameStrobe[14] Tile_X1Y4_LUT4AB/FrameStrobe[15] Tile_X1Y4_LUT4AB/FrameStrobe[16]
+ Tile_X1Y4_LUT4AB/FrameStrobe[17] Tile_X1Y4_LUT4AB/FrameStrobe[18] Tile_X1Y4_LUT4AB/FrameStrobe[19]
+ Tile_X1Y4_LUT4AB/FrameStrobe[1] Tile_X1Y4_LUT4AB/FrameStrobe[2] Tile_X1Y4_LUT4AB/FrameStrobe[3]
+ Tile_X1Y4_LUT4AB/FrameStrobe[4] Tile_X1Y4_LUT4AB/FrameStrobe[5] Tile_X1Y4_LUT4AB/FrameStrobe[6]
+ Tile_X1Y4_LUT4AB/FrameStrobe[7] Tile_X1Y4_LUT4AB/FrameStrobe[8] Tile_X1Y4_LUT4AB/FrameStrobe[9]
+ Tile_X1Y3_LUT4AB/FrameStrobe[0] Tile_X1Y3_LUT4AB/FrameStrobe[10] Tile_X1Y3_LUT4AB/FrameStrobe[11]
+ Tile_X1Y3_LUT4AB/FrameStrobe[12] Tile_X1Y3_LUT4AB/FrameStrobe[13] Tile_X1Y3_LUT4AB/FrameStrobe[14]
+ Tile_X1Y3_LUT4AB/FrameStrobe[15] Tile_X1Y3_LUT4AB/FrameStrobe[16] Tile_X1Y3_LUT4AB/FrameStrobe[17]
+ Tile_X1Y3_LUT4AB/FrameStrobe[18] Tile_X1Y3_LUT4AB/FrameStrobe[19] Tile_X1Y3_LUT4AB/FrameStrobe[1]
+ Tile_X1Y3_LUT4AB/FrameStrobe[2] Tile_X1Y3_LUT4AB/FrameStrobe[3] Tile_X1Y3_LUT4AB/FrameStrobe[4]
+ Tile_X1Y3_LUT4AB/FrameStrobe[5] Tile_X1Y3_LUT4AB/FrameStrobe[6] Tile_X1Y3_LUT4AB/FrameStrobe[7]
+ Tile_X1Y3_LUT4AB/FrameStrobe[8] Tile_X1Y3_LUT4AB/FrameStrobe[9] Tile_X1Y4_LUT4AB/N1BEG[0]
+ Tile_X1Y4_LUT4AB/N1BEG[1] Tile_X1Y4_LUT4AB/N1BEG[2] Tile_X1Y4_LUT4AB/N1BEG[3] Tile_X1Y5_LUT4AB/N1BEG[0]
+ Tile_X1Y5_LUT4AB/N1BEG[1] Tile_X1Y5_LUT4AB/N1BEG[2] Tile_X1Y5_LUT4AB/N1BEG[3] Tile_X1Y4_LUT4AB/N2BEG[0]
+ Tile_X1Y4_LUT4AB/N2BEG[1] Tile_X1Y4_LUT4AB/N2BEG[2] Tile_X1Y4_LUT4AB/N2BEG[3] Tile_X1Y4_LUT4AB/N2BEG[4]
+ Tile_X1Y4_LUT4AB/N2BEG[5] Tile_X1Y4_LUT4AB/N2BEG[6] Tile_X1Y4_LUT4AB/N2BEG[7] Tile_X1Y3_LUT4AB/N2END[0]
+ Tile_X1Y3_LUT4AB/N2END[1] Tile_X1Y3_LUT4AB/N2END[2] Tile_X1Y3_LUT4AB/N2END[3] Tile_X1Y3_LUT4AB/N2END[4]
+ Tile_X1Y3_LUT4AB/N2END[5] Tile_X1Y3_LUT4AB/N2END[6] Tile_X1Y3_LUT4AB/N2END[7] Tile_X1Y4_LUT4AB/N2END[0]
+ Tile_X1Y4_LUT4AB/N2END[1] Tile_X1Y4_LUT4AB/N2END[2] Tile_X1Y4_LUT4AB/N2END[3] Tile_X1Y4_LUT4AB/N2END[4]
+ Tile_X1Y4_LUT4AB/N2END[5] Tile_X1Y4_LUT4AB/N2END[6] Tile_X1Y4_LUT4AB/N2END[7] Tile_X1Y5_LUT4AB/N2BEG[0]
+ Tile_X1Y5_LUT4AB/N2BEG[1] Tile_X1Y5_LUT4AB/N2BEG[2] Tile_X1Y5_LUT4AB/N2BEG[3] Tile_X1Y5_LUT4AB/N2BEG[4]
+ Tile_X1Y5_LUT4AB/N2BEG[5] Tile_X1Y5_LUT4AB/N2BEG[6] Tile_X1Y5_LUT4AB/N2BEG[7] Tile_X1Y4_LUT4AB/N4BEG[0]
+ Tile_X1Y4_LUT4AB/N4BEG[10] Tile_X1Y4_LUT4AB/N4BEG[11] Tile_X1Y4_LUT4AB/N4BEG[12]
+ Tile_X1Y4_LUT4AB/N4BEG[13] Tile_X1Y4_LUT4AB/N4BEG[14] Tile_X1Y4_LUT4AB/N4BEG[15]
+ Tile_X1Y4_LUT4AB/N4BEG[1] Tile_X1Y4_LUT4AB/N4BEG[2] Tile_X1Y4_LUT4AB/N4BEG[3] Tile_X1Y4_LUT4AB/N4BEG[4]
+ Tile_X1Y4_LUT4AB/N4BEG[5] Tile_X1Y4_LUT4AB/N4BEG[6] Tile_X1Y4_LUT4AB/N4BEG[7] Tile_X1Y4_LUT4AB/N4BEG[8]
+ Tile_X1Y4_LUT4AB/N4BEG[9] Tile_X1Y5_LUT4AB/N4BEG[0] Tile_X1Y5_LUT4AB/N4BEG[10] Tile_X1Y5_LUT4AB/N4BEG[11]
+ Tile_X1Y5_LUT4AB/N4BEG[12] Tile_X1Y5_LUT4AB/N4BEG[13] Tile_X1Y5_LUT4AB/N4BEG[14]
+ Tile_X1Y5_LUT4AB/N4BEG[15] Tile_X1Y5_LUT4AB/N4BEG[1] Tile_X1Y5_LUT4AB/N4BEG[2] Tile_X1Y5_LUT4AB/N4BEG[3]
+ Tile_X1Y5_LUT4AB/N4BEG[4] Tile_X1Y5_LUT4AB/N4BEG[5] Tile_X1Y5_LUT4AB/N4BEG[6] Tile_X1Y5_LUT4AB/N4BEG[7]
+ Tile_X1Y5_LUT4AB/N4BEG[8] Tile_X1Y5_LUT4AB/N4BEG[9] Tile_X1Y4_LUT4AB/NN4BEG[0] Tile_X1Y4_LUT4AB/NN4BEG[10]
+ Tile_X1Y4_LUT4AB/NN4BEG[11] Tile_X1Y4_LUT4AB/NN4BEG[12] Tile_X1Y4_LUT4AB/NN4BEG[13]
+ Tile_X1Y4_LUT4AB/NN4BEG[14] Tile_X1Y4_LUT4AB/NN4BEG[15] Tile_X1Y4_LUT4AB/NN4BEG[1]
+ Tile_X1Y4_LUT4AB/NN4BEG[2] Tile_X1Y4_LUT4AB/NN4BEG[3] Tile_X1Y4_LUT4AB/NN4BEG[4]
+ Tile_X1Y4_LUT4AB/NN4BEG[5] Tile_X1Y4_LUT4AB/NN4BEG[6] Tile_X1Y4_LUT4AB/NN4BEG[7]
+ Tile_X1Y4_LUT4AB/NN4BEG[8] Tile_X1Y4_LUT4AB/NN4BEG[9] Tile_X1Y5_LUT4AB/NN4BEG[0]
+ Tile_X1Y5_LUT4AB/NN4BEG[10] Tile_X1Y5_LUT4AB/NN4BEG[11] Tile_X1Y5_LUT4AB/NN4BEG[12]
+ Tile_X1Y5_LUT4AB/NN4BEG[13] Tile_X1Y5_LUT4AB/NN4BEG[14] Tile_X1Y5_LUT4AB/NN4BEG[15]
+ Tile_X1Y5_LUT4AB/NN4BEG[1] Tile_X1Y5_LUT4AB/NN4BEG[2] Tile_X1Y5_LUT4AB/NN4BEG[3]
+ Tile_X1Y5_LUT4AB/NN4BEG[4] Tile_X1Y5_LUT4AB/NN4BEG[5] Tile_X1Y5_LUT4AB/NN4BEG[6]
+ Tile_X1Y5_LUT4AB/NN4BEG[7] Tile_X1Y5_LUT4AB/NN4BEG[8] Tile_X1Y5_LUT4AB/NN4BEG[9]
+ Tile_X1Y5_LUT4AB/S1END[0] Tile_X1Y5_LUT4AB/S1END[1] Tile_X1Y5_LUT4AB/S1END[2] Tile_X1Y5_LUT4AB/S1END[3]
+ Tile_X1Y4_LUT4AB/S1END[0] Tile_X1Y4_LUT4AB/S1END[1] Tile_X1Y4_LUT4AB/S1END[2] Tile_X1Y4_LUT4AB/S1END[3]
+ Tile_X1Y5_LUT4AB/S2MID[0] Tile_X1Y5_LUT4AB/S2MID[1] Tile_X1Y5_LUT4AB/S2MID[2] Tile_X1Y5_LUT4AB/S2MID[3]
+ Tile_X1Y5_LUT4AB/S2MID[4] Tile_X1Y5_LUT4AB/S2MID[5] Tile_X1Y5_LUT4AB/S2MID[6] Tile_X1Y5_LUT4AB/S2MID[7]
+ Tile_X1Y5_LUT4AB/S2END[0] Tile_X1Y5_LUT4AB/S2END[1] Tile_X1Y5_LUT4AB/S2END[2] Tile_X1Y5_LUT4AB/S2END[3]
+ Tile_X1Y5_LUT4AB/S2END[4] Tile_X1Y5_LUT4AB/S2END[5] Tile_X1Y5_LUT4AB/S2END[6] Tile_X1Y5_LUT4AB/S2END[7]
+ Tile_X1Y4_LUT4AB/S2END[0] Tile_X1Y4_LUT4AB/S2END[1] Tile_X1Y4_LUT4AB/S2END[2] Tile_X1Y4_LUT4AB/S2END[3]
+ Tile_X1Y4_LUT4AB/S2END[4] Tile_X1Y4_LUT4AB/S2END[5] Tile_X1Y4_LUT4AB/S2END[6] Tile_X1Y4_LUT4AB/S2END[7]
+ Tile_X1Y4_LUT4AB/S2MID[0] Tile_X1Y4_LUT4AB/S2MID[1] Tile_X1Y4_LUT4AB/S2MID[2] Tile_X1Y4_LUT4AB/S2MID[3]
+ Tile_X1Y4_LUT4AB/S2MID[4] Tile_X1Y4_LUT4AB/S2MID[5] Tile_X1Y4_LUT4AB/S2MID[6] Tile_X1Y4_LUT4AB/S2MID[7]
+ Tile_X1Y5_LUT4AB/S4END[0] Tile_X1Y5_LUT4AB/S4END[10] Tile_X1Y5_LUT4AB/S4END[11]
+ Tile_X1Y5_LUT4AB/S4END[12] Tile_X1Y5_LUT4AB/S4END[13] Tile_X1Y5_LUT4AB/S4END[14]
+ Tile_X1Y5_LUT4AB/S4END[15] Tile_X1Y5_LUT4AB/S4END[1] Tile_X1Y5_LUT4AB/S4END[2] Tile_X1Y5_LUT4AB/S4END[3]
+ Tile_X1Y5_LUT4AB/S4END[4] Tile_X1Y5_LUT4AB/S4END[5] Tile_X1Y5_LUT4AB/S4END[6] Tile_X1Y5_LUT4AB/S4END[7]
+ Tile_X1Y5_LUT4AB/S4END[8] Tile_X1Y5_LUT4AB/S4END[9] Tile_X1Y4_LUT4AB/S4END[0] Tile_X1Y4_LUT4AB/S4END[10]
+ Tile_X1Y4_LUT4AB/S4END[11] Tile_X1Y4_LUT4AB/S4END[12] Tile_X1Y4_LUT4AB/S4END[13]
+ Tile_X1Y4_LUT4AB/S4END[14] Tile_X1Y4_LUT4AB/S4END[15] Tile_X1Y4_LUT4AB/S4END[1]
+ Tile_X1Y4_LUT4AB/S4END[2] Tile_X1Y4_LUT4AB/S4END[3] Tile_X1Y4_LUT4AB/S4END[4] Tile_X1Y4_LUT4AB/S4END[5]
+ Tile_X1Y4_LUT4AB/S4END[6] Tile_X1Y4_LUT4AB/S4END[7] Tile_X1Y4_LUT4AB/S4END[8] Tile_X1Y4_LUT4AB/S4END[9]
+ Tile_X1Y5_LUT4AB/SS4END[0] Tile_X1Y5_LUT4AB/SS4END[10] Tile_X1Y5_LUT4AB/SS4END[11]
+ Tile_X1Y5_LUT4AB/SS4END[12] Tile_X1Y5_LUT4AB/SS4END[13] Tile_X1Y5_LUT4AB/SS4END[14]
+ Tile_X1Y5_LUT4AB/SS4END[15] Tile_X1Y5_LUT4AB/SS4END[1] Tile_X1Y5_LUT4AB/SS4END[2]
+ Tile_X1Y5_LUT4AB/SS4END[3] Tile_X1Y5_LUT4AB/SS4END[4] Tile_X1Y5_LUT4AB/SS4END[5]
+ Tile_X1Y5_LUT4AB/SS4END[6] Tile_X1Y5_LUT4AB/SS4END[7] Tile_X1Y5_LUT4AB/SS4END[8]
+ Tile_X1Y5_LUT4AB/SS4END[9] Tile_X1Y4_LUT4AB/SS4END[0] Tile_X1Y4_LUT4AB/SS4END[10]
+ Tile_X1Y4_LUT4AB/SS4END[11] Tile_X1Y4_LUT4AB/SS4END[12] Tile_X1Y4_LUT4AB/SS4END[13]
+ Tile_X1Y4_LUT4AB/SS4END[14] Tile_X1Y4_LUT4AB/SS4END[15] Tile_X1Y4_LUT4AB/SS4END[1]
+ Tile_X1Y4_LUT4AB/SS4END[2] Tile_X1Y4_LUT4AB/SS4END[3] Tile_X1Y4_LUT4AB/SS4END[4]
+ Tile_X1Y4_LUT4AB/SS4END[5] Tile_X1Y4_LUT4AB/SS4END[6] Tile_X1Y4_LUT4AB/SS4END[7]
+ Tile_X1Y4_LUT4AB/SS4END[8] Tile_X1Y4_LUT4AB/SS4END[9] Tile_X1Y4_LUT4AB/UserCLK Tile_X1Y3_LUT4AB/UserCLK
+ VGND VPWR Tile_X1Y4_LUT4AB/W1BEG[0] Tile_X1Y4_LUT4AB/W1BEG[1] Tile_X1Y4_LUT4AB/W1BEG[2]
+ Tile_X1Y4_LUT4AB/W1BEG[3] Tile_X2Y4_LUT4AB/W1BEG[0] Tile_X2Y4_LUT4AB/W1BEG[1] Tile_X2Y4_LUT4AB/W1BEG[2]
+ Tile_X2Y4_LUT4AB/W1BEG[3] Tile_X1Y4_LUT4AB/W2BEG[0] Tile_X1Y4_LUT4AB/W2BEG[1] Tile_X1Y4_LUT4AB/W2BEG[2]
+ Tile_X1Y4_LUT4AB/W2BEG[3] Tile_X1Y4_LUT4AB/W2BEG[4] Tile_X1Y4_LUT4AB/W2BEG[5] Tile_X1Y4_LUT4AB/W2BEG[6]
+ Tile_X1Y4_LUT4AB/W2BEG[7] Tile_X1Y4_LUT4AB/W2BEGb[0] Tile_X1Y4_LUT4AB/W2BEGb[1]
+ Tile_X1Y4_LUT4AB/W2BEGb[2] Tile_X1Y4_LUT4AB/W2BEGb[3] Tile_X1Y4_LUT4AB/W2BEGb[4]
+ Tile_X1Y4_LUT4AB/W2BEGb[5] Tile_X1Y4_LUT4AB/W2BEGb[6] Tile_X1Y4_LUT4AB/W2BEGb[7]
+ Tile_X1Y4_LUT4AB/W2END[0] Tile_X1Y4_LUT4AB/W2END[1] Tile_X1Y4_LUT4AB/W2END[2] Tile_X1Y4_LUT4AB/W2END[3]
+ Tile_X1Y4_LUT4AB/W2END[4] Tile_X1Y4_LUT4AB/W2END[5] Tile_X1Y4_LUT4AB/W2END[6] Tile_X1Y4_LUT4AB/W2END[7]
+ Tile_X2Y4_LUT4AB/W2BEG[0] Tile_X2Y4_LUT4AB/W2BEG[1] Tile_X2Y4_LUT4AB/W2BEG[2] Tile_X2Y4_LUT4AB/W2BEG[3]
+ Tile_X2Y4_LUT4AB/W2BEG[4] Tile_X2Y4_LUT4AB/W2BEG[5] Tile_X2Y4_LUT4AB/W2BEG[6] Tile_X2Y4_LUT4AB/W2BEG[7]
+ Tile_X1Y4_LUT4AB/W6BEG[0] Tile_X1Y4_LUT4AB/W6BEG[10] Tile_X1Y4_LUT4AB/W6BEG[11]
+ Tile_X1Y4_LUT4AB/W6BEG[1] Tile_X1Y4_LUT4AB/W6BEG[2] Tile_X1Y4_LUT4AB/W6BEG[3] Tile_X1Y4_LUT4AB/W6BEG[4]
+ Tile_X1Y4_LUT4AB/W6BEG[5] Tile_X1Y4_LUT4AB/W6BEG[6] Tile_X1Y4_LUT4AB/W6BEG[7] Tile_X1Y4_LUT4AB/W6BEG[8]
+ Tile_X1Y4_LUT4AB/W6BEG[9] Tile_X2Y4_LUT4AB/W6BEG[0] Tile_X2Y4_LUT4AB/W6BEG[10] Tile_X2Y4_LUT4AB/W6BEG[11]
+ Tile_X2Y4_LUT4AB/W6BEG[1] Tile_X2Y4_LUT4AB/W6BEG[2] Tile_X2Y4_LUT4AB/W6BEG[3] Tile_X2Y4_LUT4AB/W6BEG[4]
+ Tile_X2Y4_LUT4AB/W6BEG[5] Tile_X2Y4_LUT4AB/W6BEG[6] Tile_X2Y4_LUT4AB/W6BEG[7] Tile_X2Y4_LUT4AB/W6BEG[8]
+ Tile_X2Y4_LUT4AB/W6BEG[9] Tile_X1Y4_LUT4AB/WW4BEG[0] Tile_X1Y4_LUT4AB/WW4BEG[10]
+ Tile_X1Y4_LUT4AB/WW4BEG[11] Tile_X1Y4_LUT4AB/WW4BEG[12] Tile_X1Y4_LUT4AB/WW4BEG[13]
+ Tile_X1Y4_LUT4AB/WW4BEG[14] Tile_X1Y4_LUT4AB/WW4BEG[15] Tile_X1Y4_LUT4AB/WW4BEG[1]
+ Tile_X1Y4_LUT4AB/WW4BEG[2] Tile_X1Y4_LUT4AB/WW4BEG[3] Tile_X1Y4_LUT4AB/WW4BEG[4]
+ Tile_X1Y4_LUT4AB/WW4BEG[5] Tile_X1Y4_LUT4AB/WW4BEG[6] Tile_X1Y4_LUT4AB/WW4BEG[7]
+ Tile_X1Y4_LUT4AB/WW4BEG[8] Tile_X1Y4_LUT4AB/WW4BEG[9] Tile_X2Y4_LUT4AB/WW4BEG[0]
+ Tile_X2Y4_LUT4AB/WW4BEG[10] Tile_X2Y4_LUT4AB/WW4BEG[11] Tile_X2Y4_LUT4AB/WW4BEG[12]
+ Tile_X2Y4_LUT4AB/WW4BEG[13] Tile_X2Y4_LUT4AB/WW4BEG[14] Tile_X2Y4_LUT4AB/WW4BEG[15]
+ Tile_X2Y4_LUT4AB/WW4BEG[1] Tile_X2Y4_LUT4AB/WW4BEG[2] Tile_X2Y4_LUT4AB/WW4BEG[3]
+ Tile_X2Y4_LUT4AB/WW4BEG[4] Tile_X2Y4_LUT4AB/WW4BEG[5] Tile_X2Y4_LUT4AB/WW4BEG[6]
+ Tile_X2Y4_LUT4AB/WW4BEG[7] Tile_X2Y4_LUT4AB/WW4BEG[8] Tile_X2Y4_LUT4AB/WW4BEG[9]
+ LUT4AB
XTile_X0Y7_W_TT_IF Tile_X0Y7_CLK_TT_PROJECT Tile_X1Y7_LUT4AB/E1END[0] Tile_X1Y7_LUT4AB/E1END[1]
+ Tile_X1Y7_LUT4AB/E1END[2] Tile_X1Y7_LUT4AB/E1END[3] Tile_X1Y7_LUT4AB/E2MID[0] Tile_X1Y7_LUT4AB/E2MID[1]
+ Tile_X1Y7_LUT4AB/E2MID[2] Tile_X1Y7_LUT4AB/E2MID[3] Tile_X1Y7_LUT4AB/E2MID[4] Tile_X1Y7_LUT4AB/E2MID[5]
+ Tile_X1Y7_LUT4AB/E2MID[6] Tile_X1Y7_LUT4AB/E2MID[7] Tile_X1Y7_LUT4AB/E2END[0] Tile_X1Y7_LUT4AB/E2END[1]
+ Tile_X1Y7_LUT4AB/E2END[2] Tile_X1Y7_LUT4AB/E2END[3] Tile_X1Y7_LUT4AB/E2END[4] Tile_X1Y7_LUT4AB/E2END[5]
+ Tile_X1Y7_LUT4AB/E2END[6] Tile_X1Y7_LUT4AB/E2END[7] Tile_X1Y7_LUT4AB/E6END[0] Tile_X1Y7_LUT4AB/E6END[10]
+ Tile_X1Y7_LUT4AB/E6END[11] Tile_X1Y7_LUT4AB/E6END[1] Tile_X1Y7_LUT4AB/E6END[2] Tile_X1Y7_LUT4AB/E6END[3]
+ Tile_X1Y7_LUT4AB/E6END[4] Tile_X1Y7_LUT4AB/E6END[5] Tile_X1Y7_LUT4AB/E6END[6] Tile_X1Y7_LUT4AB/E6END[7]
+ Tile_X1Y7_LUT4AB/E6END[8] Tile_X1Y7_LUT4AB/E6END[9] Tile_X1Y7_LUT4AB/EE4END[0] Tile_X1Y7_LUT4AB/EE4END[10]
+ Tile_X1Y7_LUT4AB/EE4END[11] Tile_X1Y7_LUT4AB/EE4END[12] Tile_X1Y7_LUT4AB/EE4END[13]
+ Tile_X1Y7_LUT4AB/EE4END[14] Tile_X1Y7_LUT4AB/EE4END[15] Tile_X1Y7_LUT4AB/EE4END[1]
+ Tile_X1Y7_LUT4AB/EE4END[2] Tile_X1Y7_LUT4AB/EE4END[3] Tile_X1Y7_LUT4AB/EE4END[4]
+ Tile_X1Y7_LUT4AB/EE4END[5] Tile_X1Y7_LUT4AB/EE4END[6] Tile_X1Y7_LUT4AB/EE4END[7]
+ Tile_X1Y7_LUT4AB/EE4END[8] Tile_X1Y7_LUT4AB/EE4END[9] Tile_X0Y7_ENA_TT_PROJECT FrameData[224]
+ FrameData[234] FrameData[235] FrameData[236] FrameData[237] FrameData[238] FrameData[239]
+ FrameData[240] FrameData[241] FrameData[242] FrameData[243] FrameData[225] FrameData[244]
+ FrameData[245] FrameData[246] FrameData[247] FrameData[248] FrameData[249] FrameData[250]
+ FrameData[251] FrameData[252] FrameData[253] FrameData[226] FrameData[254] FrameData[255]
+ FrameData[227] FrameData[228] FrameData[229] FrameData[230] FrameData[231] FrameData[232]
+ FrameData[233] Tile_X1Y7_LUT4AB/FrameData[0] Tile_X1Y7_LUT4AB/FrameData[10] Tile_X1Y7_LUT4AB/FrameData[11]
+ Tile_X1Y7_LUT4AB/FrameData[12] Tile_X1Y7_LUT4AB/FrameData[13] Tile_X1Y7_LUT4AB/FrameData[14]
+ Tile_X1Y7_LUT4AB/FrameData[15] Tile_X1Y7_LUT4AB/FrameData[16] Tile_X1Y7_LUT4AB/FrameData[17]
+ Tile_X1Y7_LUT4AB/FrameData[18] Tile_X1Y7_LUT4AB/FrameData[19] Tile_X1Y7_LUT4AB/FrameData[1]
+ Tile_X1Y7_LUT4AB/FrameData[20] Tile_X1Y7_LUT4AB/FrameData[21] Tile_X1Y7_LUT4AB/FrameData[22]
+ Tile_X1Y7_LUT4AB/FrameData[23] Tile_X1Y7_LUT4AB/FrameData[24] Tile_X1Y7_LUT4AB/FrameData[25]
+ Tile_X1Y7_LUT4AB/FrameData[26] Tile_X1Y7_LUT4AB/FrameData[27] Tile_X1Y7_LUT4AB/FrameData[28]
+ Tile_X1Y7_LUT4AB/FrameData[29] Tile_X1Y7_LUT4AB/FrameData[2] Tile_X1Y7_LUT4AB/FrameData[30]
+ Tile_X1Y7_LUT4AB/FrameData[31] Tile_X1Y7_LUT4AB/FrameData[3] Tile_X1Y7_LUT4AB/FrameData[4]
+ Tile_X1Y7_LUT4AB/FrameData[5] Tile_X1Y7_LUT4AB/FrameData[6] Tile_X1Y7_LUT4AB/FrameData[7]
+ Tile_X1Y7_LUT4AB/FrameData[8] Tile_X1Y7_LUT4AB/FrameData[9] Tile_X0Y7_W_TT_IF/FrameStrobe[0]
+ Tile_X0Y7_W_TT_IF/FrameStrobe[10] Tile_X0Y7_W_TT_IF/FrameStrobe[11] Tile_X0Y7_W_TT_IF/FrameStrobe[12]
+ Tile_X0Y7_W_TT_IF/FrameStrobe[13] Tile_X0Y7_W_TT_IF/FrameStrobe[14] Tile_X0Y7_W_TT_IF/FrameStrobe[15]
+ Tile_X0Y7_W_TT_IF/FrameStrobe[16] Tile_X0Y7_W_TT_IF/FrameStrobe[17] Tile_X0Y7_W_TT_IF/FrameStrobe[18]
+ Tile_X0Y7_W_TT_IF/FrameStrobe[19] Tile_X0Y7_W_TT_IF/FrameStrobe[1] Tile_X0Y7_W_TT_IF/FrameStrobe[2]
+ Tile_X0Y7_W_TT_IF/FrameStrobe[3] Tile_X0Y7_W_TT_IF/FrameStrobe[4] Tile_X0Y7_W_TT_IF/FrameStrobe[5]
+ Tile_X0Y7_W_TT_IF/FrameStrobe[6] Tile_X0Y7_W_TT_IF/FrameStrobe[7] Tile_X0Y7_W_TT_IF/FrameStrobe[8]
+ Tile_X0Y7_W_TT_IF/FrameStrobe[9] Tile_X0Y6_W_TT_IF/FrameStrobe[0] Tile_X0Y6_W_TT_IF/FrameStrobe[10]
+ Tile_X0Y6_W_TT_IF/FrameStrobe[11] Tile_X0Y6_W_TT_IF/FrameStrobe[12] Tile_X0Y6_W_TT_IF/FrameStrobe[13]
+ Tile_X0Y6_W_TT_IF/FrameStrobe[14] Tile_X0Y6_W_TT_IF/FrameStrobe[15] Tile_X0Y6_W_TT_IF/FrameStrobe[16]
+ Tile_X0Y6_W_TT_IF/FrameStrobe[17] Tile_X0Y6_W_TT_IF/FrameStrobe[18] Tile_X0Y6_W_TT_IF/FrameStrobe[19]
+ Tile_X0Y6_W_TT_IF/FrameStrobe[1] Tile_X0Y6_W_TT_IF/FrameStrobe[2] Tile_X0Y6_W_TT_IF/FrameStrobe[3]
+ Tile_X0Y6_W_TT_IF/FrameStrobe[4] Tile_X0Y6_W_TT_IF/FrameStrobe[5] Tile_X0Y6_W_TT_IF/FrameStrobe[6]
+ Tile_X0Y6_W_TT_IF/FrameStrobe[7] Tile_X0Y6_W_TT_IF/FrameStrobe[8] Tile_X0Y6_W_TT_IF/FrameStrobe[9]
+ Tile_X0Y7_W_TT_IF/N1BEG[0] Tile_X0Y7_W_TT_IF/N1BEG[1] Tile_X0Y7_W_TT_IF/N1BEG[2]
+ Tile_X0Y7_W_TT_IF/N1BEG[3] Tile_X0Y8_W_TT_IF/N1BEG[0] Tile_X0Y8_W_TT_IF/N1BEG[1]
+ Tile_X0Y8_W_TT_IF/N1BEG[2] Tile_X0Y8_W_TT_IF/N1BEG[3] Tile_X0Y7_W_TT_IF/N2BEG[0]
+ Tile_X0Y7_W_TT_IF/N2BEG[1] Tile_X0Y7_W_TT_IF/N2BEG[2] Tile_X0Y7_W_TT_IF/N2BEG[3]
+ Tile_X0Y7_W_TT_IF/N2BEG[4] Tile_X0Y7_W_TT_IF/N2BEG[5] Tile_X0Y7_W_TT_IF/N2BEG[6]
+ Tile_X0Y7_W_TT_IF/N2BEG[7] Tile_X0Y6_W_TT_IF/N2END[0] Tile_X0Y6_W_TT_IF/N2END[1]
+ Tile_X0Y6_W_TT_IF/N2END[2] Tile_X0Y6_W_TT_IF/N2END[3] Tile_X0Y6_W_TT_IF/N2END[4]
+ Tile_X0Y6_W_TT_IF/N2END[5] Tile_X0Y6_W_TT_IF/N2END[6] Tile_X0Y6_W_TT_IF/N2END[7]
+ Tile_X0Y7_W_TT_IF/N2END[0] Tile_X0Y7_W_TT_IF/N2END[1] Tile_X0Y7_W_TT_IF/N2END[2]
+ Tile_X0Y7_W_TT_IF/N2END[3] Tile_X0Y7_W_TT_IF/N2END[4] Tile_X0Y7_W_TT_IF/N2END[5]
+ Tile_X0Y7_W_TT_IF/N2END[6] Tile_X0Y7_W_TT_IF/N2END[7] Tile_X0Y8_W_TT_IF/N2BEG[0]
+ Tile_X0Y8_W_TT_IF/N2BEG[1] Tile_X0Y8_W_TT_IF/N2BEG[2] Tile_X0Y8_W_TT_IF/N2BEG[3]
+ Tile_X0Y8_W_TT_IF/N2BEG[4] Tile_X0Y8_W_TT_IF/N2BEG[5] Tile_X0Y8_W_TT_IF/N2BEG[6]
+ Tile_X0Y8_W_TT_IF/N2BEG[7] Tile_X0Y7_W_TT_IF/N4BEG[0] Tile_X0Y7_W_TT_IF/N4BEG[10]
+ Tile_X0Y7_W_TT_IF/N4BEG[11] Tile_X0Y7_W_TT_IF/N4BEG[12] Tile_X0Y7_W_TT_IF/N4BEG[13]
+ Tile_X0Y7_W_TT_IF/N4BEG[14] Tile_X0Y7_W_TT_IF/N4BEG[15] Tile_X0Y7_W_TT_IF/N4BEG[1]
+ Tile_X0Y7_W_TT_IF/N4BEG[2] Tile_X0Y7_W_TT_IF/N4BEG[3] Tile_X0Y7_W_TT_IF/N4BEG[4]
+ Tile_X0Y7_W_TT_IF/N4BEG[5] Tile_X0Y7_W_TT_IF/N4BEG[6] Tile_X0Y7_W_TT_IF/N4BEG[7]
+ Tile_X0Y7_W_TT_IF/N4BEG[8] Tile_X0Y7_W_TT_IF/N4BEG[9] Tile_X0Y8_W_TT_IF/N4BEG[0]
+ Tile_X0Y8_W_TT_IF/N4BEG[10] Tile_X0Y8_W_TT_IF/N4BEG[11] Tile_X0Y8_W_TT_IF/N4BEG[12]
+ Tile_X0Y8_W_TT_IF/N4BEG[13] Tile_X0Y8_W_TT_IF/N4BEG[14] Tile_X0Y8_W_TT_IF/N4BEG[15]
+ Tile_X0Y8_W_TT_IF/N4BEG[1] Tile_X0Y8_W_TT_IF/N4BEG[2] Tile_X0Y8_W_TT_IF/N4BEG[3]
+ Tile_X0Y8_W_TT_IF/N4BEG[4] Tile_X0Y8_W_TT_IF/N4BEG[5] Tile_X0Y8_W_TT_IF/N4BEG[6]
+ Tile_X0Y8_W_TT_IF/N4BEG[7] Tile_X0Y8_W_TT_IF/N4BEG[8] Tile_X0Y8_W_TT_IF/N4BEG[9]
+ Tile_X0Y7_RST_N_TT_PROJECT Tile_X0Y8_W_TT_IF/S1END[0] Tile_X0Y8_W_TT_IF/S1END[1]
+ Tile_X0Y8_W_TT_IF/S1END[2] Tile_X0Y8_W_TT_IF/S1END[3] Tile_X0Y7_W_TT_IF/S1END[0]
+ Tile_X0Y7_W_TT_IF/S1END[1] Tile_X0Y7_W_TT_IF/S1END[2] Tile_X0Y7_W_TT_IF/S1END[3]
+ Tile_X0Y8_W_TT_IF/S2MID[0] Tile_X0Y8_W_TT_IF/S2MID[1] Tile_X0Y8_W_TT_IF/S2MID[2]
+ Tile_X0Y8_W_TT_IF/S2MID[3] Tile_X0Y8_W_TT_IF/S2MID[4] Tile_X0Y8_W_TT_IF/S2MID[5]
+ Tile_X0Y8_W_TT_IF/S2MID[6] Tile_X0Y8_W_TT_IF/S2MID[7] Tile_X0Y8_W_TT_IF/S2END[0]
+ Tile_X0Y8_W_TT_IF/S2END[1] Tile_X0Y8_W_TT_IF/S2END[2] Tile_X0Y8_W_TT_IF/S2END[3]
+ Tile_X0Y8_W_TT_IF/S2END[4] Tile_X0Y8_W_TT_IF/S2END[5] Tile_X0Y8_W_TT_IF/S2END[6]
+ Tile_X0Y8_W_TT_IF/S2END[7] Tile_X0Y7_W_TT_IF/S2END[0] Tile_X0Y7_W_TT_IF/S2END[1]
+ Tile_X0Y7_W_TT_IF/S2END[2] Tile_X0Y7_W_TT_IF/S2END[3] Tile_X0Y7_W_TT_IF/S2END[4]
+ Tile_X0Y7_W_TT_IF/S2END[5] Tile_X0Y7_W_TT_IF/S2END[6] Tile_X0Y7_W_TT_IF/S2END[7]
+ Tile_X0Y7_W_TT_IF/S2MID[0] Tile_X0Y7_W_TT_IF/S2MID[1] Tile_X0Y7_W_TT_IF/S2MID[2]
+ Tile_X0Y7_W_TT_IF/S2MID[3] Tile_X0Y7_W_TT_IF/S2MID[4] Tile_X0Y7_W_TT_IF/S2MID[5]
+ Tile_X0Y7_W_TT_IF/S2MID[6] Tile_X0Y7_W_TT_IF/S2MID[7] Tile_X0Y8_W_TT_IF/S4END[0]
+ Tile_X0Y8_W_TT_IF/S4END[10] Tile_X0Y8_W_TT_IF/S4END[11] Tile_X0Y8_W_TT_IF/S4END[12]
+ Tile_X0Y8_W_TT_IF/S4END[13] Tile_X0Y8_W_TT_IF/S4END[14] Tile_X0Y8_W_TT_IF/S4END[15]
+ Tile_X0Y8_W_TT_IF/S4END[1] Tile_X0Y8_W_TT_IF/S4END[2] Tile_X0Y8_W_TT_IF/S4END[3]
+ Tile_X0Y8_W_TT_IF/S4END[4] Tile_X0Y8_W_TT_IF/S4END[5] Tile_X0Y8_W_TT_IF/S4END[6]
+ Tile_X0Y8_W_TT_IF/S4END[7] Tile_X0Y8_W_TT_IF/S4END[8] Tile_X0Y8_W_TT_IF/S4END[9]
+ Tile_X0Y7_W_TT_IF/S4END[0] Tile_X0Y7_W_TT_IF/S4END[10] Tile_X0Y7_W_TT_IF/S4END[11]
+ Tile_X0Y7_W_TT_IF/S4END[12] Tile_X0Y7_W_TT_IF/S4END[13] Tile_X0Y7_W_TT_IF/S4END[14]
+ Tile_X0Y7_W_TT_IF/S4END[15] Tile_X0Y7_W_TT_IF/S4END[1] Tile_X0Y7_W_TT_IF/S4END[2]
+ Tile_X0Y7_W_TT_IF/S4END[3] Tile_X0Y7_W_TT_IF/S4END[4] Tile_X0Y7_W_TT_IF/S4END[5]
+ Tile_X0Y7_W_TT_IF/S4END[6] Tile_X0Y7_W_TT_IF/S4END[7] Tile_X0Y7_W_TT_IF/S4END[8]
+ Tile_X0Y7_W_TT_IF/S4END[9] Tile_X0Y7_UIO_IN_TT_PROJECT0 Tile_X0Y7_UIO_IN_TT_PROJECT1
+ Tile_X0Y7_UIO_IN_TT_PROJECT2 Tile_X0Y7_UIO_IN_TT_PROJECT3 Tile_X0Y7_UIO_IN_TT_PROJECT4
+ Tile_X0Y7_UIO_IN_TT_PROJECT5 Tile_X0Y7_UIO_IN_TT_PROJECT6 Tile_X0Y7_UIO_IN_TT_PROJECT7
+ Tile_X0Y7_UIO_OE_TT_PROJECT0 Tile_X0Y7_UIO_OE_TT_PROJECT1 Tile_X0Y7_UIO_OE_TT_PROJECT2
+ Tile_X0Y7_UIO_OE_TT_PROJECT3 Tile_X0Y7_UIO_OE_TT_PROJECT4 Tile_X0Y7_UIO_OE_TT_PROJECT5
+ Tile_X0Y7_UIO_OE_TT_PROJECT6 Tile_X0Y7_UIO_OE_TT_PROJECT7 Tile_X0Y7_UIO_OUT_TT_PROJECT0
+ Tile_X0Y7_UIO_OUT_TT_PROJECT1 Tile_X0Y7_UIO_OUT_TT_PROJECT2 Tile_X0Y7_UIO_OUT_TT_PROJECT3
+ Tile_X0Y7_UIO_OUT_TT_PROJECT4 Tile_X0Y7_UIO_OUT_TT_PROJECT5 Tile_X0Y7_UIO_OUT_TT_PROJECT6
+ Tile_X0Y7_UIO_OUT_TT_PROJECT7 Tile_X0Y7_UI_IN_TT_PROJECT0 Tile_X0Y7_UI_IN_TT_PROJECT1
+ Tile_X0Y7_UI_IN_TT_PROJECT2 Tile_X0Y7_UI_IN_TT_PROJECT3 Tile_X0Y7_UI_IN_TT_PROJECT4
+ Tile_X0Y7_UI_IN_TT_PROJECT5 Tile_X0Y7_UI_IN_TT_PROJECT6 Tile_X0Y7_UI_IN_TT_PROJECT7
+ Tile_X0Y7_UO_OUT_TT_PROJECT0 Tile_X0Y7_UO_OUT_TT_PROJECT1 Tile_X0Y7_UO_OUT_TT_PROJECT2
+ Tile_X0Y7_UO_OUT_TT_PROJECT3 Tile_X0Y7_UO_OUT_TT_PROJECT4 Tile_X0Y7_UO_OUT_TT_PROJECT5
+ Tile_X0Y7_UO_OUT_TT_PROJECT6 Tile_X0Y7_UO_OUT_TT_PROJECT7 Tile_X0Y7_W_TT_IF/UserCLK
+ Tile_X0Y6_W_TT_IF/UserCLK VGND VPWR Tile_X1Y7_LUT4AB/W1BEG[0] Tile_X1Y7_LUT4AB/W1BEG[1]
+ Tile_X1Y7_LUT4AB/W1BEG[2] Tile_X1Y7_LUT4AB/W1BEG[3] Tile_X1Y7_LUT4AB/W2BEGb[0] Tile_X1Y7_LUT4AB/W2BEGb[1]
+ Tile_X1Y7_LUT4AB/W2BEGb[2] Tile_X1Y7_LUT4AB/W2BEGb[3] Tile_X1Y7_LUT4AB/W2BEGb[4]
+ Tile_X1Y7_LUT4AB/W2BEGb[5] Tile_X1Y7_LUT4AB/W2BEGb[6] Tile_X1Y7_LUT4AB/W2BEGb[7]
+ Tile_X1Y7_LUT4AB/W2BEG[0] Tile_X1Y7_LUT4AB/W2BEG[1] Tile_X1Y7_LUT4AB/W2BEG[2] Tile_X1Y7_LUT4AB/W2BEG[3]
+ Tile_X1Y7_LUT4AB/W2BEG[4] Tile_X1Y7_LUT4AB/W2BEG[5] Tile_X1Y7_LUT4AB/W2BEG[6] Tile_X1Y7_LUT4AB/W2BEG[7]
+ Tile_X1Y7_LUT4AB/W6BEG[0] Tile_X1Y7_LUT4AB/W6BEG[10] Tile_X1Y7_LUT4AB/W6BEG[11]
+ Tile_X1Y7_LUT4AB/W6BEG[1] Tile_X1Y7_LUT4AB/W6BEG[2] Tile_X1Y7_LUT4AB/W6BEG[3] Tile_X1Y7_LUT4AB/W6BEG[4]
+ Tile_X1Y7_LUT4AB/W6BEG[5] Tile_X1Y7_LUT4AB/W6BEG[6] Tile_X1Y7_LUT4AB/W6BEG[7] Tile_X1Y7_LUT4AB/W6BEG[8]
+ Tile_X1Y7_LUT4AB/W6BEG[9] Tile_X1Y7_LUT4AB/WW4BEG[0] Tile_X1Y7_LUT4AB/WW4BEG[10]
+ Tile_X1Y7_LUT4AB/WW4BEG[11] Tile_X1Y7_LUT4AB/WW4BEG[12] Tile_X1Y7_LUT4AB/WW4BEG[13]
+ Tile_X1Y7_LUT4AB/WW4BEG[14] Tile_X1Y7_LUT4AB/WW4BEG[15] Tile_X1Y7_LUT4AB/WW4BEG[1]
+ Tile_X1Y7_LUT4AB/WW4BEG[2] Tile_X1Y7_LUT4AB/WW4BEG[3] Tile_X1Y7_LUT4AB/WW4BEG[4]
+ Tile_X1Y7_LUT4AB/WW4BEG[5] Tile_X1Y7_LUT4AB/WW4BEG[6] Tile_X1Y7_LUT4AB/WW4BEG[7]
+ Tile_X1Y7_LUT4AB/WW4BEG[8] Tile_X1Y7_LUT4AB/WW4BEG[9] W_TT_IF
XTile_X0Y3_W_TT_IF Tile_X0Y3_CLK_TT_PROJECT Tile_X1Y3_LUT4AB/E1END[0] Tile_X1Y3_LUT4AB/E1END[1]
+ Tile_X1Y3_LUT4AB/E1END[2] Tile_X1Y3_LUT4AB/E1END[3] Tile_X1Y3_LUT4AB/E2MID[0] Tile_X1Y3_LUT4AB/E2MID[1]
+ Tile_X1Y3_LUT4AB/E2MID[2] Tile_X1Y3_LUT4AB/E2MID[3] Tile_X1Y3_LUT4AB/E2MID[4] Tile_X1Y3_LUT4AB/E2MID[5]
+ Tile_X1Y3_LUT4AB/E2MID[6] Tile_X1Y3_LUT4AB/E2MID[7] Tile_X1Y3_LUT4AB/E2END[0] Tile_X1Y3_LUT4AB/E2END[1]
+ Tile_X1Y3_LUT4AB/E2END[2] Tile_X1Y3_LUT4AB/E2END[3] Tile_X1Y3_LUT4AB/E2END[4] Tile_X1Y3_LUT4AB/E2END[5]
+ Tile_X1Y3_LUT4AB/E2END[6] Tile_X1Y3_LUT4AB/E2END[7] Tile_X1Y3_LUT4AB/E6END[0] Tile_X1Y3_LUT4AB/E6END[10]
+ Tile_X1Y3_LUT4AB/E6END[11] Tile_X1Y3_LUT4AB/E6END[1] Tile_X1Y3_LUT4AB/E6END[2] Tile_X1Y3_LUT4AB/E6END[3]
+ Tile_X1Y3_LUT4AB/E6END[4] Tile_X1Y3_LUT4AB/E6END[5] Tile_X1Y3_LUT4AB/E6END[6] Tile_X1Y3_LUT4AB/E6END[7]
+ Tile_X1Y3_LUT4AB/E6END[8] Tile_X1Y3_LUT4AB/E6END[9] Tile_X1Y3_LUT4AB/EE4END[0] Tile_X1Y3_LUT4AB/EE4END[10]
+ Tile_X1Y3_LUT4AB/EE4END[11] Tile_X1Y3_LUT4AB/EE4END[12] Tile_X1Y3_LUT4AB/EE4END[13]
+ Tile_X1Y3_LUT4AB/EE4END[14] Tile_X1Y3_LUT4AB/EE4END[15] Tile_X1Y3_LUT4AB/EE4END[1]
+ Tile_X1Y3_LUT4AB/EE4END[2] Tile_X1Y3_LUT4AB/EE4END[3] Tile_X1Y3_LUT4AB/EE4END[4]
+ Tile_X1Y3_LUT4AB/EE4END[5] Tile_X1Y3_LUT4AB/EE4END[6] Tile_X1Y3_LUT4AB/EE4END[7]
+ Tile_X1Y3_LUT4AB/EE4END[8] Tile_X1Y3_LUT4AB/EE4END[9] Tile_X0Y3_ENA_TT_PROJECT FrameData[96]
+ FrameData[106] FrameData[107] FrameData[108] FrameData[109] FrameData[110] FrameData[111]
+ FrameData[112] FrameData[113] FrameData[114] FrameData[115] FrameData[97] FrameData[116]
+ FrameData[117] FrameData[118] FrameData[119] FrameData[120] FrameData[121] FrameData[122]
+ FrameData[123] FrameData[124] FrameData[125] FrameData[98] FrameData[126] FrameData[127]
+ FrameData[99] FrameData[100] FrameData[101] FrameData[102] FrameData[103] FrameData[104]
+ FrameData[105] Tile_X1Y3_LUT4AB/FrameData[0] Tile_X1Y3_LUT4AB/FrameData[10] Tile_X1Y3_LUT4AB/FrameData[11]
+ Tile_X1Y3_LUT4AB/FrameData[12] Tile_X1Y3_LUT4AB/FrameData[13] Tile_X1Y3_LUT4AB/FrameData[14]
+ Tile_X1Y3_LUT4AB/FrameData[15] Tile_X1Y3_LUT4AB/FrameData[16] Tile_X1Y3_LUT4AB/FrameData[17]
+ Tile_X1Y3_LUT4AB/FrameData[18] Tile_X1Y3_LUT4AB/FrameData[19] Tile_X1Y3_LUT4AB/FrameData[1]
+ Tile_X1Y3_LUT4AB/FrameData[20] Tile_X1Y3_LUT4AB/FrameData[21] Tile_X1Y3_LUT4AB/FrameData[22]
+ Tile_X1Y3_LUT4AB/FrameData[23] Tile_X1Y3_LUT4AB/FrameData[24] Tile_X1Y3_LUT4AB/FrameData[25]
+ Tile_X1Y3_LUT4AB/FrameData[26] Tile_X1Y3_LUT4AB/FrameData[27] Tile_X1Y3_LUT4AB/FrameData[28]
+ Tile_X1Y3_LUT4AB/FrameData[29] Tile_X1Y3_LUT4AB/FrameData[2] Tile_X1Y3_LUT4AB/FrameData[30]
+ Tile_X1Y3_LUT4AB/FrameData[31] Tile_X1Y3_LUT4AB/FrameData[3] Tile_X1Y3_LUT4AB/FrameData[4]
+ Tile_X1Y3_LUT4AB/FrameData[5] Tile_X1Y3_LUT4AB/FrameData[6] Tile_X1Y3_LUT4AB/FrameData[7]
+ Tile_X1Y3_LUT4AB/FrameData[8] Tile_X1Y3_LUT4AB/FrameData[9] Tile_X0Y3_W_TT_IF/FrameStrobe[0]
+ Tile_X0Y3_W_TT_IF/FrameStrobe[10] Tile_X0Y3_W_TT_IF/FrameStrobe[11] Tile_X0Y3_W_TT_IF/FrameStrobe[12]
+ Tile_X0Y3_W_TT_IF/FrameStrobe[13] Tile_X0Y3_W_TT_IF/FrameStrobe[14] Tile_X0Y3_W_TT_IF/FrameStrobe[15]
+ Tile_X0Y3_W_TT_IF/FrameStrobe[16] Tile_X0Y3_W_TT_IF/FrameStrobe[17] Tile_X0Y3_W_TT_IF/FrameStrobe[18]
+ Tile_X0Y3_W_TT_IF/FrameStrobe[19] Tile_X0Y3_W_TT_IF/FrameStrobe[1] Tile_X0Y3_W_TT_IF/FrameStrobe[2]
+ Tile_X0Y3_W_TT_IF/FrameStrobe[3] Tile_X0Y3_W_TT_IF/FrameStrobe[4] Tile_X0Y3_W_TT_IF/FrameStrobe[5]
+ Tile_X0Y3_W_TT_IF/FrameStrobe[6] Tile_X0Y3_W_TT_IF/FrameStrobe[7] Tile_X0Y3_W_TT_IF/FrameStrobe[8]
+ Tile_X0Y3_W_TT_IF/FrameStrobe[9] Tile_X0Y2_W_TT_IF/FrameStrobe[0] Tile_X0Y2_W_TT_IF/FrameStrobe[10]
+ Tile_X0Y2_W_TT_IF/FrameStrobe[11] Tile_X0Y2_W_TT_IF/FrameStrobe[12] Tile_X0Y2_W_TT_IF/FrameStrobe[13]
+ Tile_X0Y2_W_TT_IF/FrameStrobe[14] Tile_X0Y2_W_TT_IF/FrameStrobe[15] Tile_X0Y2_W_TT_IF/FrameStrobe[16]
+ Tile_X0Y2_W_TT_IF/FrameStrobe[17] Tile_X0Y2_W_TT_IF/FrameStrobe[18] Tile_X0Y2_W_TT_IF/FrameStrobe[19]
+ Tile_X0Y2_W_TT_IF/FrameStrobe[1] Tile_X0Y2_W_TT_IF/FrameStrobe[2] Tile_X0Y2_W_TT_IF/FrameStrobe[3]
+ Tile_X0Y2_W_TT_IF/FrameStrobe[4] Tile_X0Y2_W_TT_IF/FrameStrobe[5] Tile_X0Y2_W_TT_IF/FrameStrobe[6]
+ Tile_X0Y2_W_TT_IF/FrameStrobe[7] Tile_X0Y2_W_TT_IF/FrameStrobe[8] Tile_X0Y2_W_TT_IF/FrameStrobe[9]
+ Tile_X0Y3_W_TT_IF/N1BEG[0] Tile_X0Y3_W_TT_IF/N1BEG[1] Tile_X0Y3_W_TT_IF/N1BEG[2]
+ Tile_X0Y3_W_TT_IF/N1BEG[3] Tile_X0Y4_W_TT_IF/N1BEG[0] Tile_X0Y4_W_TT_IF/N1BEG[1]
+ Tile_X0Y4_W_TT_IF/N1BEG[2] Tile_X0Y4_W_TT_IF/N1BEG[3] Tile_X0Y3_W_TT_IF/N2BEG[0]
+ Tile_X0Y3_W_TT_IF/N2BEG[1] Tile_X0Y3_W_TT_IF/N2BEG[2] Tile_X0Y3_W_TT_IF/N2BEG[3]
+ Tile_X0Y3_W_TT_IF/N2BEG[4] Tile_X0Y3_W_TT_IF/N2BEG[5] Tile_X0Y3_W_TT_IF/N2BEG[6]
+ Tile_X0Y3_W_TT_IF/N2BEG[7] Tile_X0Y2_W_TT_IF/N2END[0] Tile_X0Y2_W_TT_IF/N2END[1]
+ Tile_X0Y2_W_TT_IF/N2END[2] Tile_X0Y2_W_TT_IF/N2END[3] Tile_X0Y2_W_TT_IF/N2END[4]
+ Tile_X0Y2_W_TT_IF/N2END[5] Tile_X0Y2_W_TT_IF/N2END[6] Tile_X0Y2_W_TT_IF/N2END[7]
+ Tile_X0Y3_W_TT_IF/N2END[0] Tile_X0Y3_W_TT_IF/N2END[1] Tile_X0Y3_W_TT_IF/N2END[2]
+ Tile_X0Y3_W_TT_IF/N2END[3] Tile_X0Y3_W_TT_IF/N2END[4] Tile_X0Y3_W_TT_IF/N2END[5]
+ Tile_X0Y3_W_TT_IF/N2END[6] Tile_X0Y3_W_TT_IF/N2END[7] Tile_X0Y4_W_TT_IF/N2BEG[0]
+ Tile_X0Y4_W_TT_IF/N2BEG[1] Tile_X0Y4_W_TT_IF/N2BEG[2] Tile_X0Y4_W_TT_IF/N2BEG[3]
+ Tile_X0Y4_W_TT_IF/N2BEG[4] Tile_X0Y4_W_TT_IF/N2BEG[5] Tile_X0Y4_W_TT_IF/N2BEG[6]
+ Tile_X0Y4_W_TT_IF/N2BEG[7] Tile_X0Y3_W_TT_IF/N4BEG[0] Tile_X0Y3_W_TT_IF/N4BEG[10]
+ Tile_X0Y3_W_TT_IF/N4BEG[11] Tile_X0Y3_W_TT_IF/N4BEG[12] Tile_X0Y3_W_TT_IF/N4BEG[13]
+ Tile_X0Y3_W_TT_IF/N4BEG[14] Tile_X0Y3_W_TT_IF/N4BEG[15] Tile_X0Y3_W_TT_IF/N4BEG[1]
+ Tile_X0Y3_W_TT_IF/N4BEG[2] Tile_X0Y3_W_TT_IF/N4BEG[3] Tile_X0Y3_W_TT_IF/N4BEG[4]
+ Tile_X0Y3_W_TT_IF/N4BEG[5] Tile_X0Y3_W_TT_IF/N4BEG[6] Tile_X0Y3_W_TT_IF/N4BEG[7]
+ Tile_X0Y3_W_TT_IF/N4BEG[8] Tile_X0Y3_W_TT_IF/N4BEG[9] Tile_X0Y4_W_TT_IF/N4BEG[0]
+ Tile_X0Y4_W_TT_IF/N4BEG[10] Tile_X0Y4_W_TT_IF/N4BEG[11] Tile_X0Y4_W_TT_IF/N4BEG[12]
+ Tile_X0Y4_W_TT_IF/N4BEG[13] Tile_X0Y4_W_TT_IF/N4BEG[14] Tile_X0Y4_W_TT_IF/N4BEG[15]
+ Tile_X0Y4_W_TT_IF/N4BEG[1] Tile_X0Y4_W_TT_IF/N4BEG[2] Tile_X0Y4_W_TT_IF/N4BEG[3]
+ Tile_X0Y4_W_TT_IF/N4BEG[4] Tile_X0Y4_W_TT_IF/N4BEG[5] Tile_X0Y4_W_TT_IF/N4BEG[6]
+ Tile_X0Y4_W_TT_IF/N4BEG[7] Tile_X0Y4_W_TT_IF/N4BEG[8] Tile_X0Y4_W_TT_IF/N4BEG[9]
+ Tile_X0Y3_RST_N_TT_PROJECT Tile_X0Y4_W_TT_IF/S1END[0] Tile_X0Y4_W_TT_IF/S1END[1]
+ Tile_X0Y4_W_TT_IF/S1END[2] Tile_X0Y4_W_TT_IF/S1END[3] Tile_X0Y3_W_TT_IF/S1END[0]
+ Tile_X0Y3_W_TT_IF/S1END[1] Tile_X0Y3_W_TT_IF/S1END[2] Tile_X0Y3_W_TT_IF/S1END[3]
+ Tile_X0Y4_W_TT_IF/S2MID[0] Tile_X0Y4_W_TT_IF/S2MID[1] Tile_X0Y4_W_TT_IF/S2MID[2]
+ Tile_X0Y4_W_TT_IF/S2MID[3] Tile_X0Y4_W_TT_IF/S2MID[4] Tile_X0Y4_W_TT_IF/S2MID[5]
+ Tile_X0Y4_W_TT_IF/S2MID[6] Tile_X0Y4_W_TT_IF/S2MID[7] Tile_X0Y4_W_TT_IF/S2END[0]
+ Tile_X0Y4_W_TT_IF/S2END[1] Tile_X0Y4_W_TT_IF/S2END[2] Tile_X0Y4_W_TT_IF/S2END[3]
+ Tile_X0Y4_W_TT_IF/S2END[4] Tile_X0Y4_W_TT_IF/S2END[5] Tile_X0Y4_W_TT_IF/S2END[6]
+ Tile_X0Y4_W_TT_IF/S2END[7] Tile_X0Y3_W_TT_IF/S2END[0] Tile_X0Y3_W_TT_IF/S2END[1]
+ Tile_X0Y3_W_TT_IF/S2END[2] Tile_X0Y3_W_TT_IF/S2END[3] Tile_X0Y3_W_TT_IF/S2END[4]
+ Tile_X0Y3_W_TT_IF/S2END[5] Tile_X0Y3_W_TT_IF/S2END[6] Tile_X0Y3_W_TT_IF/S2END[7]
+ Tile_X0Y3_W_TT_IF/S2MID[0] Tile_X0Y3_W_TT_IF/S2MID[1] Tile_X0Y3_W_TT_IF/S2MID[2]
+ Tile_X0Y3_W_TT_IF/S2MID[3] Tile_X0Y3_W_TT_IF/S2MID[4] Tile_X0Y3_W_TT_IF/S2MID[5]
+ Tile_X0Y3_W_TT_IF/S2MID[6] Tile_X0Y3_W_TT_IF/S2MID[7] Tile_X0Y4_W_TT_IF/S4END[0]
+ Tile_X0Y4_W_TT_IF/S4END[10] Tile_X0Y4_W_TT_IF/S4END[11] Tile_X0Y4_W_TT_IF/S4END[12]
+ Tile_X0Y4_W_TT_IF/S4END[13] Tile_X0Y4_W_TT_IF/S4END[14] Tile_X0Y4_W_TT_IF/S4END[15]
+ Tile_X0Y4_W_TT_IF/S4END[1] Tile_X0Y4_W_TT_IF/S4END[2] Tile_X0Y4_W_TT_IF/S4END[3]
+ Tile_X0Y4_W_TT_IF/S4END[4] Tile_X0Y4_W_TT_IF/S4END[5] Tile_X0Y4_W_TT_IF/S4END[6]
+ Tile_X0Y4_W_TT_IF/S4END[7] Tile_X0Y4_W_TT_IF/S4END[8] Tile_X0Y4_W_TT_IF/S4END[9]
+ Tile_X0Y3_W_TT_IF/S4END[0] Tile_X0Y3_W_TT_IF/S4END[10] Tile_X0Y3_W_TT_IF/S4END[11]
+ Tile_X0Y3_W_TT_IF/S4END[12] Tile_X0Y3_W_TT_IF/S4END[13] Tile_X0Y3_W_TT_IF/S4END[14]
+ Tile_X0Y3_W_TT_IF/S4END[15] Tile_X0Y3_W_TT_IF/S4END[1] Tile_X0Y3_W_TT_IF/S4END[2]
+ Tile_X0Y3_W_TT_IF/S4END[3] Tile_X0Y3_W_TT_IF/S4END[4] Tile_X0Y3_W_TT_IF/S4END[5]
+ Tile_X0Y3_W_TT_IF/S4END[6] Tile_X0Y3_W_TT_IF/S4END[7] Tile_X0Y3_W_TT_IF/S4END[8]
+ Tile_X0Y3_W_TT_IF/S4END[9] Tile_X0Y3_UIO_IN_TT_PROJECT0 Tile_X0Y3_UIO_IN_TT_PROJECT1
+ Tile_X0Y3_UIO_IN_TT_PROJECT2 Tile_X0Y3_UIO_IN_TT_PROJECT3 Tile_X0Y3_UIO_IN_TT_PROJECT4
+ Tile_X0Y3_UIO_IN_TT_PROJECT5 Tile_X0Y3_UIO_IN_TT_PROJECT6 Tile_X0Y3_UIO_IN_TT_PROJECT7
+ Tile_X0Y3_UIO_OE_TT_PROJECT0 Tile_X0Y3_UIO_OE_TT_PROJECT1 Tile_X0Y3_UIO_OE_TT_PROJECT2
+ Tile_X0Y3_UIO_OE_TT_PROJECT3 Tile_X0Y3_UIO_OE_TT_PROJECT4 Tile_X0Y3_UIO_OE_TT_PROJECT5
+ Tile_X0Y3_UIO_OE_TT_PROJECT6 Tile_X0Y3_UIO_OE_TT_PROJECT7 Tile_X0Y3_UIO_OUT_TT_PROJECT0
+ Tile_X0Y3_UIO_OUT_TT_PROJECT1 Tile_X0Y3_UIO_OUT_TT_PROJECT2 Tile_X0Y3_UIO_OUT_TT_PROJECT3
+ Tile_X0Y3_UIO_OUT_TT_PROJECT4 Tile_X0Y3_UIO_OUT_TT_PROJECT5 Tile_X0Y3_UIO_OUT_TT_PROJECT6
+ Tile_X0Y3_UIO_OUT_TT_PROJECT7 Tile_X0Y3_UI_IN_TT_PROJECT0 Tile_X0Y3_UI_IN_TT_PROJECT1
+ Tile_X0Y3_UI_IN_TT_PROJECT2 Tile_X0Y3_UI_IN_TT_PROJECT3 Tile_X0Y3_UI_IN_TT_PROJECT4
+ Tile_X0Y3_UI_IN_TT_PROJECT5 Tile_X0Y3_UI_IN_TT_PROJECT6 Tile_X0Y3_UI_IN_TT_PROJECT7
+ Tile_X0Y3_UO_OUT_TT_PROJECT0 Tile_X0Y3_UO_OUT_TT_PROJECT1 Tile_X0Y3_UO_OUT_TT_PROJECT2
+ Tile_X0Y3_UO_OUT_TT_PROJECT3 Tile_X0Y3_UO_OUT_TT_PROJECT4 Tile_X0Y3_UO_OUT_TT_PROJECT5
+ Tile_X0Y3_UO_OUT_TT_PROJECT6 Tile_X0Y3_UO_OUT_TT_PROJECT7 Tile_X0Y3_W_TT_IF/UserCLK
+ Tile_X0Y2_W_TT_IF/UserCLK VGND VPWR Tile_X1Y3_LUT4AB/W1BEG[0] Tile_X1Y3_LUT4AB/W1BEG[1]
+ Tile_X1Y3_LUT4AB/W1BEG[2] Tile_X1Y3_LUT4AB/W1BEG[3] Tile_X1Y3_LUT4AB/W2BEGb[0] Tile_X1Y3_LUT4AB/W2BEGb[1]
+ Tile_X1Y3_LUT4AB/W2BEGb[2] Tile_X1Y3_LUT4AB/W2BEGb[3] Tile_X1Y3_LUT4AB/W2BEGb[4]
+ Tile_X1Y3_LUT4AB/W2BEGb[5] Tile_X1Y3_LUT4AB/W2BEGb[6] Tile_X1Y3_LUT4AB/W2BEGb[7]
+ Tile_X1Y3_LUT4AB/W2BEG[0] Tile_X1Y3_LUT4AB/W2BEG[1] Tile_X1Y3_LUT4AB/W2BEG[2] Tile_X1Y3_LUT4AB/W2BEG[3]
+ Tile_X1Y3_LUT4AB/W2BEG[4] Tile_X1Y3_LUT4AB/W2BEG[5] Tile_X1Y3_LUT4AB/W2BEG[6] Tile_X1Y3_LUT4AB/W2BEG[7]
+ Tile_X1Y3_LUT4AB/W6BEG[0] Tile_X1Y3_LUT4AB/W6BEG[10] Tile_X1Y3_LUT4AB/W6BEG[11]
+ Tile_X1Y3_LUT4AB/W6BEG[1] Tile_X1Y3_LUT4AB/W6BEG[2] Tile_X1Y3_LUT4AB/W6BEG[3] Tile_X1Y3_LUT4AB/W6BEG[4]
+ Tile_X1Y3_LUT4AB/W6BEG[5] Tile_X1Y3_LUT4AB/W6BEG[6] Tile_X1Y3_LUT4AB/W6BEG[7] Tile_X1Y3_LUT4AB/W6BEG[8]
+ Tile_X1Y3_LUT4AB/W6BEG[9] Tile_X1Y3_LUT4AB/WW4BEG[0] Tile_X1Y3_LUT4AB/WW4BEG[10]
+ Tile_X1Y3_LUT4AB/WW4BEG[11] Tile_X1Y3_LUT4AB/WW4BEG[12] Tile_X1Y3_LUT4AB/WW4BEG[13]
+ Tile_X1Y3_LUT4AB/WW4BEG[14] Tile_X1Y3_LUT4AB/WW4BEG[15] Tile_X1Y3_LUT4AB/WW4BEG[1]
+ Tile_X1Y3_LUT4AB/WW4BEG[2] Tile_X1Y3_LUT4AB/WW4BEG[3] Tile_X1Y3_LUT4AB/WW4BEG[4]
+ Tile_X1Y3_LUT4AB/WW4BEG[5] Tile_X1Y3_LUT4AB/WW4BEG[6] Tile_X1Y3_LUT4AB/WW4BEG[7]
+ Tile_X1Y3_LUT4AB/WW4BEG[8] Tile_X1Y3_LUT4AB/WW4BEG[9] W_TT_IF
XTile_X3Y2_LUT4AB Tile_X3Y3_LUT4AB/Co Tile_X3Y2_LUT4AB/Co Tile_X4Y2_LUT4AB/E1END[0]
+ Tile_X4Y2_LUT4AB/E1END[1] Tile_X4Y2_LUT4AB/E1END[2] Tile_X4Y2_LUT4AB/E1END[3] Tile_X3Y2_LUT4AB/E1END[0]
+ Tile_X3Y2_LUT4AB/E1END[1] Tile_X3Y2_LUT4AB/E1END[2] Tile_X3Y2_LUT4AB/E1END[3] Tile_X4Y2_LUT4AB/E2MID[0]
+ Tile_X4Y2_LUT4AB/E2MID[1] Tile_X4Y2_LUT4AB/E2MID[2] Tile_X4Y2_LUT4AB/E2MID[3] Tile_X4Y2_LUT4AB/E2MID[4]
+ Tile_X4Y2_LUT4AB/E2MID[5] Tile_X4Y2_LUT4AB/E2MID[6] Tile_X4Y2_LUT4AB/E2MID[7] Tile_X4Y2_LUT4AB/E2END[0]
+ Tile_X4Y2_LUT4AB/E2END[1] Tile_X4Y2_LUT4AB/E2END[2] Tile_X4Y2_LUT4AB/E2END[3] Tile_X4Y2_LUT4AB/E2END[4]
+ Tile_X4Y2_LUT4AB/E2END[5] Tile_X4Y2_LUT4AB/E2END[6] Tile_X4Y2_LUT4AB/E2END[7] Tile_X3Y2_LUT4AB/E2END[0]
+ Tile_X3Y2_LUT4AB/E2END[1] Tile_X3Y2_LUT4AB/E2END[2] Tile_X3Y2_LUT4AB/E2END[3] Tile_X3Y2_LUT4AB/E2END[4]
+ Tile_X3Y2_LUT4AB/E2END[5] Tile_X3Y2_LUT4AB/E2END[6] Tile_X3Y2_LUT4AB/E2END[7] Tile_X3Y2_LUT4AB/E2MID[0]
+ Tile_X3Y2_LUT4AB/E2MID[1] Tile_X3Y2_LUT4AB/E2MID[2] Tile_X3Y2_LUT4AB/E2MID[3] Tile_X3Y2_LUT4AB/E2MID[4]
+ Tile_X3Y2_LUT4AB/E2MID[5] Tile_X3Y2_LUT4AB/E2MID[6] Tile_X3Y2_LUT4AB/E2MID[7] Tile_X4Y2_LUT4AB/E6END[0]
+ Tile_X4Y2_LUT4AB/E6END[10] Tile_X4Y2_LUT4AB/E6END[11] Tile_X4Y2_LUT4AB/E6END[1]
+ Tile_X4Y2_LUT4AB/E6END[2] Tile_X4Y2_LUT4AB/E6END[3] Tile_X4Y2_LUT4AB/E6END[4] Tile_X4Y2_LUT4AB/E6END[5]
+ Tile_X4Y2_LUT4AB/E6END[6] Tile_X4Y2_LUT4AB/E6END[7] Tile_X4Y2_LUT4AB/E6END[8] Tile_X4Y2_LUT4AB/E6END[9]
+ Tile_X3Y2_LUT4AB/E6END[0] Tile_X3Y2_LUT4AB/E6END[10] Tile_X3Y2_LUT4AB/E6END[11]
+ Tile_X3Y2_LUT4AB/E6END[1] Tile_X3Y2_LUT4AB/E6END[2] Tile_X3Y2_LUT4AB/E6END[3] Tile_X3Y2_LUT4AB/E6END[4]
+ Tile_X3Y2_LUT4AB/E6END[5] Tile_X3Y2_LUT4AB/E6END[6] Tile_X3Y2_LUT4AB/E6END[7] Tile_X3Y2_LUT4AB/E6END[8]
+ Tile_X3Y2_LUT4AB/E6END[9] Tile_X4Y2_LUT4AB/EE4END[0] Tile_X4Y2_LUT4AB/EE4END[10]
+ Tile_X4Y2_LUT4AB/EE4END[11] Tile_X4Y2_LUT4AB/EE4END[12] Tile_X4Y2_LUT4AB/EE4END[13]
+ Tile_X4Y2_LUT4AB/EE4END[14] Tile_X4Y2_LUT4AB/EE4END[15] Tile_X4Y2_LUT4AB/EE4END[1]
+ Tile_X4Y2_LUT4AB/EE4END[2] Tile_X4Y2_LUT4AB/EE4END[3] Tile_X4Y2_LUT4AB/EE4END[4]
+ Tile_X4Y2_LUT4AB/EE4END[5] Tile_X4Y2_LUT4AB/EE4END[6] Tile_X4Y2_LUT4AB/EE4END[7]
+ Tile_X4Y2_LUT4AB/EE4END[8] Tile_X4Y2_LUT4AB/EE4END[9] Tile_X3Y2_LUT4AB/EE4END[0]
+ Tile_X3Y2_LUT4AB/EE4END[10] Tile_X3Y2_LUT4AB/EE4END[11] Tile_X3Y2_LUT4AB/EE4END[12]
+ Tile_X3Y2_LUT4AB/EE4END[13] Tile_X3Y2_LUT4AB/EE4END[14] Tile_X3Y2_LUT4AB/EE4END[15]
+ Tile_X3Y2_LUT4AB/EE4END[1] Tile_X3Y2_LUT4AB/EE4END[2] Tile_X3Y2_LUT4AB/EE4END[3]
+ Tile_X3Y2_LUT4AB/EE4END[4] Tile_X3Y2_LUT4AB/EE4END[5] Tile_X3Y2_LUT4AB/EE4END[6]
+ Tile_X3Y2_LUT4AB/EE4END[7] Tile_X3Y2_LUT4AB/EE4END[8] Tile_X3Y2_LUT4AB/EE4END[9]
+ Tile_X3Y2_LUT4AB/FrameData[0] Tile_X3Y2_LUT4AB/FrameData[10] Tile_X3Y2_LUT4AB/FrameData[11]
+ Tile_X3Y2_LUT4AB/FrameData[12] Tile_X3Y2_LUT4AB/FrameData[13] Tile_X3Y2_LUT4AB/FrameData[14]
+ Tile_X3Y2_LUT4AB/FrameData[15] Tile_X3Y2_LUT4AB/FrameData[16] Tile_X3Y2_LUT4AB/FrameData[17]
+ Tile_X3Y2_LUT4AB/FrameData[18] Tile_X3Y2_LUT4AB/FrameData[19] Tile_X3Y2_LUT4AB/FrameData[1]
+ Tile_X3Y2_LUT4AB/FrameData[20] Tile_X3Y2_LUT4AB/FrameData[21] Tile_X3Y2_LUT4AB/FrameData[22]
+ Tile_X3Y2_LUT4AB/FrameData[23] Tile_X3Y2_LUT4AB/FrameData[24] Tile_X3Y2_LUT4AB/FrameData[25]
+ Tile_X3Y2_LUT4AB/FrameData[26] Tile_X3Y2_LUT4AB/FrameData[27] Tile_X3Y2_LUT4AB/FrameData[28]
+ Tile_X3Y2_LUT4AB/FrameData[29] Tile_X3Y2_LUT4AB/FrameData[2] Tile_X3Y2_LUT4AB/FrameData[30]
+ Tile_X3Y2_LUT4AB/FrameData[31] Tile_X3Y2_LUT4AB/FrameData[3] Tile_X3Y2_LUT4AB/FrameData[4]
+ Tile_X3Y2_LUT4AB/FrameData[5] Tile_X3Y2_LUT4AB/FrameData[6] Tile_X3Y2_LUT4AB/FrameData[7]
+ Tile_X3Y2_LUT4AB/FrameData[8] Tile_X3Y2_LUT4AB/FrameData[9] Tile_X4Y2_LUT4AB/FrameData[0]
+ Tile_X4Y2_LUT4AB/FrameData[10] Tile_X4Y2_LUT4AB/FrameData[11] Tile_X4Y2_LUT4AB/FrameData[12]
+ Tile_X4Y2_LUT4AB/FrameData[13] Tile_X4Y2_LUT4AB/FrameData[14] Tile_X4Y2_LUT4AB/FrameData[15]
+ Tile_X4Y2_LUT4AB/FrameData[16] Tile_X4Y2_LUT4AB/FrameData[17] Tile_X4Y2_LUT4AB/FrameData[18]
+ Tile_X4Y2_LUT4AB/FrameData[19] Tile_X4Y2_LUT4AB/FrameData[1] Tile_X4Y2_LUT4AB/FrameData[20]
+ Tile_X4Y2_LUT4AB/FrameData[21] Tile_X4Y2_LUT4AB/FrameData[22] Tile_X4Y2_LUT4AB/FrameData[23]
+ Tile_X4Y2_LUT4AB/FrameData[24] Tile_X4Y2_LUT4AB/FrameData[25] Tile_X4Y2_LUT4AB/FrameData[26]
+ Tile_X4Y2_LUT4AB/FrameData[27] Tile_X4Y2_LUT4AB/FrameData[28] Tile_X4Y2_LUT4AB/FrameData[29]
+ Tile_X4Y2_LUT4AB/FrameData[2] Tile_X4Y2_LUT4AB/FrameData[30] Tile_X4Y2_LUT4AB/FrameData[31]
+ Tile_X4Y2_LUT4AB/FrameData[3] Tile_X4Y2_LUT4AB/FrameData[4] Tile_X4Y2_LUT4AB/FrameData[5]
+ Tile_X4Y2_LUT4AB/FrameData[6] Tile_X4Y2_LUT4AB/FrameData[7] Tile_X4Y2_LUT4AB/FrameData[8]
+ Tile_X4Y2_LUT4AB/FrameData[9] Tile_X3Y2_LUT4AB/FrameStrobe[0] Tile_X3Y2_LUT4AB/FrameStrobe[10]
+ Tile_X3Y2_LUT4AB/FrameStrobe[11] Tile_X3Y2_LUT4AB/FrameStrobe[12] Tile_X3Y2_LUT4AB/FrameStrobe[13]
+ Tile_X3Y2_LUT4AB/FrameStrobe[14] Tile_X3Y2_LUT4AB/FrameStrobe[15] Tile_X3Y2_LUT4AB/FrameStrobe[16]
+ Tile_X3Y2_LUT4AB/FrameStrobe[17] Tile_X3Y2_LUT4AB/FrameStrobe[18] Tile_X3Y2_LUT4AB/FrameStrobe[19]
+ Tile_X3Y2_LUT4AB/FrameStrobe[1] Tile_X3Y2_LUT4AB/FrameStrobe[2] Tile_X3Y2_LUT4AB/FrameStrobe[3]
+ Tile_X3Y2_LUT4AB/FrameStrobe[4] Tile_X3Y2_LUT4AB/FrameStrobe[5] Tile_X3Y2_LUT4AB/FrameStrobe[6]
+ Tile_X3Y2_LUT4AB/FrameStrobe[7] Tile_X3Y2_LUT4AB/FrameStrobe[8] Tile_X3Y2_LUT4AB/FrameStrobe[9]
+ Tile_X3Y1_LUT4AB/FrameStrobe[0] Tile_X3Y1_LUT4AB/FrameStrobe[10] Tile_X3Y1_LUT4AB/FrameStrobe[11]
+ Tile_X3Y1_LUT4AB/FrameStrobe[12] Tile_X3Y1_LUT4AB/FrameStrobe[13] Tile_X3Y1_LUT4AB/FrameStrobe[14]
+ Tile_X3Y1_LUT4AB/FrameStrobe[15] Tile_X3Y1_LUT4AB/FrameStrobe[16] Tile_X3Y1_LUT4AB/FrameStrobe[17]
+ Tile_X3Y1_LUT4AB/FrameStrobe[18] Tile_X3Y1_LUT4AB/FrameStrobe[19] Tile_X3Y1_LUT4AB/FrameStrobe[1]
+ Tile_X3Y1_LUT4AB/FrameStrobe[2] Tile_X3Y1_LUT4AB/FrameStrobe[3] Tile_X3Y1_LUT4AB/FrameStrobe[4]
+ Tile_X3Y1_LUT4AB/FrameStrobe[5] Tile_X3Y1_LUT4AB/FrameStrobe[6] Tile_X3Y1_LUT4AB/FrameStrobe[7]
+ Tile_X3Y1_LUT4AB/FrameStrobe[8] Tile_X3Y1_LUT4AB/FrameStrobe[9] Tile_X3Y2_LUT4AB/N1BEG[0]
+ Tile_X3Y2_LUT4AB/N1BEG[1] Tile_X3Y2_LUT4AB/N1BEG[2] Tile_X3Y2_LUT4AB/N1BEG[3] Tile_X3Y3_LUT4AB/N1BEG[0]
+ Tile_X3Y3_LUT4AB/N1BEG[1] Tile_X3Y3_LUT4AB/N1BEG[2] Tile_X3Y3_LUT4AB/N1BEG[3] Tile_X3Y2_LUT4AB/N2BEG[0]
+ Tile_X3Y2_LUT4AB/N2BEG[1] Tile_X3Y2_LUT4AB/N2BEG[2] Tile_X3Y2_LUT4AB/N2BEG[3] Tile_X3Y2_LUT4AB/N2BEG[4]
+ Tile_X3Y2_LUT4AB/N2BEG[5] Tile_X3Y2_LUT4AB/N2BEG[6] Tile_X3Y2_LUT4AB/N2BEG[7] Tile_X3Y1_LUT4AB/N2END[0]
+ Tile_X3Y1_LUT4AB/N2END[1] Tile_X3Y1_LUT4AB/N2END[2] Tile_X3Y1_LUT4AB/N2END[3] Tile_X3Y1_LUT4AB/N2END[4]
+ Tile_X3Y1_LUT4AB/N2END[5] Tile_X3Y1_LUT4AB/N2END[6] Tile_X3Y1_LUT4AB/N2END[7] Tile_X3Y2_LUT4AB/N2END[0]
+ Tile_X3Y2_LUT4AB/N2END[1] Tile_X3Y2_LUT4AB/N2END[2] Tile_X3Y2_LUT4AB/N2END[3] Tile_X3Y2_LUT4AB/N2END[4]
+ Tile_X3Y2_LUT4AB/N2END[5] Tile_X3Y2_LUT4AB/N2END[6] Tile_X3Y2_LUT4AB/N2END[7] Tile_X3Y3_LUT4AB/N2BEG[0]
+ Tile_X3Y3_LUT4AB/N2BEG[1] Tile_X3Y3_LUT4AB/N2BEG[2] Tile_X3Y3_LUT4AB/N2BEG[3] Tile_X3Y3_LUT4AB/N2BEG[4]
+ Tile_X3Y3_LUT4AB/N2BEG[5] Tile_X3Y3_LUT4AB/N2BEG[6] Tile_X3Y3_LUT4AB/N2BEG[7] Tile_X3Y2_LUT4AB/N4BEG[0]
+ Tile_X3Y2_LUT4AB/N4BEG[10] Tile_X3Y2_LUT4AB/N4BEG[11] Tile_X3Y2_LUT4AB/N4BEG[12]
+ Tile_X3Y2_LUT4AB/N4BEG[13] Tile_X3Y2_LUT4AB/N4BEG[14] Tile_X3Y2_LUT4AB/N4BEG[15]
+ Tile_X3Y2_LUT4AB/N4BEG[1] Tile_X3Y2_LUT4AB/N4BEG[2] Tile_X3Y2_LUT4AB/N4BEG[3] Tile_X3Y2_LUT4AB/N4BEG[4]
+ Tile_X3Y2_LUT4AB/N4BEG[5] Tile_X3Y2_LUT4AB/N4BEG[6] Tile_X3Y2_LUT4AB/N4BEG[7] Tile_X3Y2_LUT4AB/N4BEG[8]
+ Tile_X3Y2_LUT4AB/N4BEG[9] Tile_X3Y3_LUT4AB/N4BEG[0] Tile_X3Y3_LUT4AB/N4BEG[10] Tile_X3Y3_LUT4AB/N4BEG[11]
+ Tile_X3Y3_LUT4AB/N4BEG[12] Tile_X3Y3_LUT4AB/N4BEG[13] Tile_X3Y3_LUT4AB/N4BEG[14]
+ Tile_X3Y3_LUT4AB/N4BEG[15] Tile_X3Y3_LUT4AB/N4BEG[1] Tile_X3Y3_LUT4AB/N4BEG[2] Tile_X3Y3_LUT4AB/N4BEG[3]
+ Tile_X3Y3_LUT4AB/N4BEG[4] Tile_X3Y3_LUT4AB/N4BEG[5] Tile_X3Y3_LUT4AB/N4BEG[6] Tile_X3Y3_LUT4AB/N4BEG[7]
+ Tile_X3Y3_LUT4AB/N4BEG[8] Tile_X3Y3_LUT4AB/N4BEG[9] Tile_X3Y2_LUT4AB/NN4BEG[0] Tile_X3Y2_LUT4AB/NN4BEG[10]
+ Tile_X3Y2_LUT4AB/NN4BEG[11] Tile_X3Y2_LUT4AB/NN4BEG[12] Tile_X3Y2_LUT4AB/NN4BEG[13]
+ Tile_X3Y2_LUT4AB/NN4BEG[14] Tile_X3Y2_LUT4AB/NN4BEG[15] Tile_X3Y2_LUT4AB/NN4BEG[1]
+ Tile_X3Y2_LUT4AB/NN4BEG[2] Tile_X3Y2_LUT4AB/NN4BEG[3] Tile_X3Y2_LUT4AB/NN4BEG[4]
+ Tile_X3Y2_LUT4AB/NN4BEG[5] Tile_X3Y2_LUT4AB/NN4BEG[6] Tile_X3Y2_LUT4AB/NN4BEG[7]
+ Tile_X3Y2_LUT4AB/NN4BEG[8] Tile_X3Y2_LUT4AB/NN4BEG[9] Tile_X3Y3_LUT4AB/NN4BEG[0]
+ Tile_X3Y3_LUT4AB/NN4BEG[10] Tile_X3Y3_LUT4AB/NN4BEG[11] Tile_X3Y3_LUT4AB/NN4BEG[12]
+ Tile_X3Y3_LUT4AB/NN4BEG[13] Tile_X3Y3_LUT4AB/NN4BEG[14] Tile_X3Y3_LUT4AB/NN4BEG[15]
+ Tile_X3Y3_LUT4AB/NN4BEG[1] Tile_X3Y3_LUT4AB/NN4BEG[2] Tile_X3Y3_LUT4AB/NN4BEG[3]
+ Tile_X3Y3_LUT4AB/NN4BEG[4] Tile_X3Y3_LUT4AB/NN4BEG[5] Tile_X3Y3_LUT4AB/NN4BEG[6]
+ Tile_X3Y3_LUT4AB/NN4BEG[7] Tile_X3Y3_LUT4AB/NN4BEG[8] Tile_X3Y3_LUT4AB/NN4BEG[9]
+ Tile_X3Y3_LUT4AB/S1END[0] Tile_X3Y3_LUT4AB/S1END[1] Tile_X3Y3_LUT4AB/S1END[2] Tile_X3Y3_LUT4AB/S1END[3]
+ Tile_X3Y2_LUT4AB/S1END[0] Tile_X3Y2_LUT4AB/S1END[1] Tile_X3Y2_LUT4AB/S1END[2] Tile_X3Y2_LUT4AB/S1END[3]
+ Tile_X3Y3_LUT4AB/S2MID[0] Tile_X3Y3_LUT4AB/S2MID[1] Tile_X3Y3_LUT4AB/S2MID[2] Tile_X3Y3_LUT4AB/S2MID[3]
+ Tile_X3Y3_LUT4AB/S2MID[4] Tile_X3Y3_LUT4AB/S2MID[5] Tile_X3Y3_LUT4AB/S2MID[6] Tile_X3Y3_LUT4AB/S2MID[7]
+ Tile_X3Y3_LUT4AB/S2END[0] Tile_X3Y3_LUT4AB/S2END[1] Tile_X3Y3_LUT4AB/S2END[2] Tile_X3Y3_LUT4AB/S2END[3]
+ Tile_X3Y3_LUT4AB/S2END[4] Tile_X3Y3_LUT4AB/S2END[5] Tile_X3Y3_LUT4AB/S2END[6] Tile_X3Y3_LUT4AB/S2END[7]
+ Tile_X3Y2_LUT4AB/S2END[0] Tile_X3Y2_LUT4AB/S2END[1] Tile_X3Y2_LUT4AB/S2END[2] Tile_X3Y2_LUT4AB/S2END[3]
+ Tile_X3Y2_LUT4AB/S2END[4] Tile_X3Y2_LUT4AB/S2END[5] Tile_X3Y2_LUT4AB/S2END[6] Tile_X3Y2_LUT4AB/S2END[7]
+ Tile_X3Y2_LUT4AB/S2MID[0] Tile_X3Y2_LUT4AB/S2MID[1] Tile_X3Y2_LUT4AB/S2MID[2] Tile_X3Y2_LUT4AB/S2MID[3]
+ Tile_X3Y2_LUT4AB/S2MID[4] Tile_X3Y2_LUT4AB/S2MID[5] Tile_X3Y2_LUT4AB/S2MID[6] Tile_X3Y2_LUT4AB/S2MID[7]
+ Tile_X3Y3_LUT4AB/S4END[0] Tile_X3Y3_LUT4AB/S4END[10] Tile_X3Y3_LUT4AB/S4END[11]
+ Tile_X3Y3_LUT4AB/S4END[12] Tile_X3Y3_LUT4AB/S4END[13] Tile_X3Y3_LUT4AB/S4END[14]
+ Tile_X3Y3_LUT4AB/S4END[15] Tile_X3Y3_LUT4AB/S4END[1] Tile_X3Y3_LUT4AB/S4END[2] Tile_X3Y3_LUT4AB/S4END[3]
+ Tile_X3Y3_LUT4AB/S4END[4] Tile_X3Y3_LUT4AB/S4END[5] Tile_X3Y3_LUT4AB/S4END[6] Tile_X3Y3_LUT4AB/S4END[7]
+ Tile_X3Y3_LUT4AB/S4END[8] Tile_X3Y3_LUT4AB/S4END[9] Tile_X3Y2_LUT4AB/S4END[0] Tile_X3Y2_LUT4AB/S4END[10]
+ Tile_X3Y2_LUT4AB/S4END[11] Tile_X3Y2_LUT4AB/S4END[12] Tile_X3Y2_LUT4AB/S4END[13]
+ Tile_X3Y2_LUT4AB/S4END[14] Tile_X3Y2_LUT4AB/S4END[15] Tile_X3Y2_LUT4AB/S4END[1]
+ Tile_X3Y2_LUT4AB/S4END[2] Tile_X3Y2_LUT4AB/S4END[3] Tile_X3Y2_LUT4AB/S4END[4] Tile_X3Y2_LUT4AB/S4END[5]
+ Tile_X3Y2_LUT4AB/S4END[6] Tile_X3Y2_LUT4AB/S4END[7] Tile_X3Y2_LUT4AB/S4END[8] Tile_X3Y2_LUT4AB/S4END[9]
+ Tile_X3Y3_LUT4AB/SS4END[0] Tile_X3Y3_LUT4AB/SS4END[10] Tile_X3Y3_LUT4AB/SS4END[11]
+ Tile_X3Y3_LUT4AB/SS4END[12] Tile_X3Y3_LUT4AB/SS4END[13] Tile_X3Y3_LUT4AB/SS4END[14]
+ Tile_X3Y3_LUT4AB/SS4END[15] Tile_X3Y3_LUT4AB/SS4END[1] Tile_X3Y3_LUT4AB/SS4END[2]
+ Tile_X3Y3_LUT4AB/SS4END[3] Tile_X3Y3_LUT4AB/SS4END[4] Tile_X3Y3_LUT4AB/SS4END[5]
+ Tile_X3Y3_LUT4AB/SS4END[6] Tile_X3Y3_LUT4AB/SS4END[7] Tile_X3Y3_LUT4AB/SS4END[8]
+ Tile_X3Y3_LUT4AB/SS4END[9] Tile_X3Y2_LUT4AB/SS4END[0] Tile_X3Y2_LUT4AB/SS4END[10]
+ Tile_X3Y2_LUT4AB/SS4END[11] Tile_X3Y2_LUT4AB/SS4END[12] Tile_X3Y2_LUT4AB/SS4END[13]
+ Tile_X3Y2_LUT4AB/SS4END[14] Tile_X3Y2_LUT4AB/SS4END[15] Tile_X3Y2_LUT4AB/SS4END[1]
+ Tile_X3Y2_LUT4AB/SS4END[2] Tile_X3Y2_LUT4AB/SS4END[3] Tile_X3Y2_LUT4AB/SS4END[4]
+ Tile_X3Y2_LUT4AB/SS4END[5] Tile_X3Y2_LUT4AB/SS4END[6] Tile_X3Y2_LUT4AB/SS4END[7]
+ Tile_X3Y2_LUT4AB/SS4END[8] Tile_X3Y2_LUT4AB/SS4END[9] Tile_X3Y2_LUT4AB/UserCLK Tile_X3Y1_LUT4AB/UserCLK
+ VGND VPWR Tile_X3Y2_LUT4AB/W1BEG[0] Tile_X3Y2_LUT4AB/W1BEG[1] Tile_X3Y2_LUT4AB/W1BEG[2]
+ Tile_X3Y2_LUT4AB/W1BEG[3] Tile_X4Y2_LUT4AB/W1BEG[0] Tile_X4Y2_LUT4AB/W1BEG[1] Tile_X4Y2_LUT4AB/W1BEG[2]
+ Tile_X4Y2_LUT4AB/W1BEG[3] Tile_X3Y2_LUT4AB/W2BEG[0] Tile_X3Y2_LUT4AB/W2BEG[1] Tile_X3Y2_LUT4AB/W2BEG[2]
+ Tile_X3Y2_LUT4AB/W2BEG[3] Tile_X3Y2_LUT4AB/W2BEG[4] Tile_X3Y2_LUT4AB/W2BEG[5] Tile_X3Y2_LUT4AB/W2BEG[6]
+ Tile_X3Y2_LUT4AB/W2BEG[7] Tile_X2Y2_LUT4AB/W2END[0] Tile_X2Y2_LUT4AB/W2END[1] Tile_X2Y2_LUT4AB/W2END[2]
+ Tile_X2Y2_LUT4AB/W2END[3] Tile_X2Y2_LUT4AB/W2END[4] Tile_X2Y2_LUT4AB/W2END[5] Tile_X2Y2_LUT4AB/W2END[6]
+ Tile_X2Y2_LUT4AB/W2END[7] Tile_X3Y2_LUT4AB/W2END[0] Tile_X3Y2_LUT4AB/W2END[1] Tile_X3Y2_LUT4AB/W2END[2]
+ Tile_X3Y2_LUT4AB/W2END[3] Tile_X3Y2_LUT4AB/W2END[4] Tile_X3Y2_LUT4AB/W2END[5] Tile_X3Y2_LUT4AB/W2END[6]
+ Tile_X3Y2_LUT4AB/W2END[7] Tile_X4Y2_LUT4AB/W2BEG[0] Tile_X4Y2_LUT4AB/W2BEG[1] Tile_X4Y2_LUT4AB/W2BEG[2]
+ Tile_X4Y2_LUT4AB/W2BEG[3] Tile_X4Y2_LUT4AB/W2BEG[4] Tile_X4Y2_LUT4AB/W2BEG[5] Tile_X4Y2_LUT4AB/W2BEG[6]
+ Tile_X4Y2_LUT4AB/W2BEG[7] Tile_X3Y2_LUT4AB/W6BEG[0] Tile_X3Y2_LUT4AB/W6BEG[10] Tile_X3Y2_LUT4AB/W6BEG[11]
+ Tile_X3Y2_LUT4AB/W6BEG[1] Tile_X3Y2_LUT4AB/W6BEG[2] Tile_X3Y2_LUT4AB/W6BEG[3] Tile_X3Y2_LUT4AB/W6BEG[4]
+ Tile_X3Y2_LUT4AB/W6BEG[5] Tile_X3Y2_LUT4AB/W6BEG[6] Tile_X3Y2_LUT4AB/W6BEG[7] Tile_X3Y2_LUT4AB/W6BEG[8]
+ Tile_X3Y2_LUT4AB/W6BEG[9] Tile_X4Y2_LUT4AB/W6BEG[0] Tile_X4Y2_LUT4AB/W6BEG[10] Tile_X4Y2_LUT4AB/W6BEG[11]
+ Tile_X4Y2_LUT4AB/W6BEG[1] Tile_X4Y2_LUT4AB/W6BEG[2] Tile_X4Y2_LUT4AB/W6BEG[3] Tile_X4Y2_LUT4AB/W6BEG[4]
+ Tile_X4Y2_LUT4AB/W6BEG[5] Tile_X4Y2_LUT4AB/W6BEG[6] Tile_X4Y2_LUT4AB/W6BEG[7] Tile_X4Y2_LUT4AB/W6BEG[8]
+ Tile_X4Y2_LUT4AB/W6BEG[9] Tile_X3Y2_LUT4AB/WW4BEG[0] Tile_X3Y2_LUT4AB/WW4BEG[10]
+ Tile_X3Y2_LUT4AB/WW4BEG[11] Tile_X3Y2_LUT4AB/WW4BEG[12] Tile_X3Y2_LUT4AB/WW4BEG[13]
+ Tile_X3Y2_LUT4AB/WW4BEG[14] Tile_X3Y2_LUT4AB/WW4BEG[15] Tile_X3Y2_LUT4AB/WW4BEG[1]
+ Tile_X3Y2_LUT4AB/WW4BEG[2] Tile_X3Y2_LUT4AB/WW4BEG[3] Tile_X3Y2_LUT4AB/WW4BEG[4]
+ Tile_X3Y2_LUT4AB/WW4BEG[5] Tile_X3Y2_LUT4AB/WW4BEG[6] Tile_X3Y2_LUT4AB/WW4BEG[7]
+ Tile_X3Y2_LUT4AB/WW4BEG[8] Tile_X3Y2_LUT4AB/WW4BEG[9] Tile_X4Y2_LUT4AB/WW4BEG[0]
+ Tile_X4Y2_LUT4AB/WW4BEG[10] Tile_X4Y2_LUT4AB/WW4BEG[11] Tile_X4Y2_LUT4AB/WW4BEG[12]
+ Tile_X4Y2_LUT4AB/WW4BEG[13] Tile_X4Y2_LUT4AB/WW4BEG[14] Tile_X4Y2_LUT4AB/WW4BEG[15]
+ Tile_X4Y2_LUT4AB/WW4BEG[1] Tile_X4Y2_LUT4AB/WW4BEG[2] Tile_X4Y2_LUT4AB/WW4BEG[3]
+ Tile_X4Y2_LUT4AB/WW4BEG[4] Tile_X4Y2_LUT4AB/WW4BEG[5] Tile_X4Y2_LUT4AB/WW4BEG[6]
+ Tile_X4Y2_LUT4AB/WW4BEG[7] Tile_X4Y2_LUT4AB/WW4BEG[8] Tile_X4Y2_LUT4AB/WW4BEG[9]
+ LUT4AB
XTile_X2Y6_LUT4AB Tile_X2Y7_LUT4AB/Co Tile_X2Y6_LUT4AB/Co Tile_X3Y6_LUT4AB/E1END[0]
+ Tile_X3Y6_LUT4AB/E1END[1] Tile_X3Y6_LUT4AB/E1END[2] Tile_X3Y6_LUT4AB/E1END[3] Tile_X2Y6_LUT4AB/E1END[0]
+ Tile_X2Y6_LUT4AB/E1END[1] Tile_X2Y6_LUT4AB/E1END[2] Tile_X2Y6_LUT4AB/E1END[3] Tile_X3Y6_LUT4AB/E2MID[0]
+ Tile_X3Y6_LUT4AB/E2MID[1] Tile_X3Y6_LUT4AB/E2MID[2] Tile_X3Y6_LUT4AB/E2MID[3] Tile_X3Y6_LUT4AB/E2MID[4]
+ Tile_X3Y6_LUT4AB/E2MID[5] Tile_X3Y6_LUT4AB/E2MID[6] Tile_X3Y6_LUT4AB/E2MID[7] Tile_X3Y6_LUT4AB/E2END[0]
+ Tile_X3Y6_LUT4AB/E2END[1] Tile_X3Y6_LUT4AB/E2END[2] Tile_X3Y6_LUT4AB/E2END[3] Tile_X3Y6_LUT4AB/E2END[4]
+ Tile_X3Y6_LUT4AB/E2END[5] Tile_X3Y6_LUT4AB/E2END[6] Tile_X3Y6_LUT4AB/E2END[7] Tile_X2Y6_LUT4AB/E2END[0]
+ Tile_X2Y6_LUT4AB/E2END[1] Tile_X2Y6_LUT4AB/E2END[2] Tile_X2Y6_LUT4AB/E2END[3] Tile_X2Y6_LUT4AB/E2END[4]
+ Tile_X2Y6_LUT4AB/E2END[5] Tile_X2Y6_LUT4AB/E2END[6] Tile_X2Y6_LUT4AB/E2END[7] Tile_X2Y6_LUT4AB/E2MID[0]
+ Tile_X2Y6_LUT4AB/E2MID[1] Tile_X2Y6_LUT4AB/E2MID[2] Tile_X2Y6_LUT4AB/E2MID[3] Tile_X2Y6_LUT4AB/E2MID[4]
+ Tile_X2Y6_LUT4AB/E2MID[5] Tile_X2Y6_LUT4AB/E2MID[6] Tile_X2Y6_LUT4AB/E2MID[7] Tile_X3Y6_LUT4AB/E6END[0]
+ Tile_X3Y6_LUT4AB/E6END[10] Tile_X3Y6_LUT4AB/E6END[11] Tile_X3Y6_LUT4AB/E6END[1]
+ Tile_X3Y6_LUT4AB/E6END[2] Tile_X3Y6_LUT4AB/E6END[3] Tile_X3Y6_LUT4AB/E6END[4] Tile_X3Y6_LUT4AB/E6END[5]
+ Tile_X3Y6_LUT4AB/E6END[6] Tile_X3Y6_LUT4AB/E6END[7] Tile_X3Y6_LUT4AB/E6END[8] Tile_X3Y6_LUT4AB/E6END[9]
+ Tile_X2Y6_LUT4AB/E6END[0] Tile_X2Y6_LUT4AB/E6END[10] Tile_X2Y6_LUT4AB/E6END[11]
+ Tile_X2Y6_LUT4AB/E6END[1] Tile_X2Y6_LUT4AB/E6END[2] Tile_X2Y6_LUT4AB/E6END[3] Tile_X2Y6_LUT4AB/E6END[4]
+ Tile_X2Y6_LUT4AB/E6END[5] Tile_X2Y6_LUT4AB/E6END[6] Tile_X2Y6_LUT4AB/E6END[7] Tile_X2Y6_LUT4AB/E6END[8]
+ Tile_X2Y6_LUT4AB/E6END[9] Tile_X3Y6_LUT4AB/EE4END[0] Tile_X3Y6_LUT4AB/EE4END[10]
+ Tile_X3Y6_LUT4AB/EE4END[11] Tile_X3Y6_LUT4AB/EE4END[12] Tile_X3Y6_LUT4AB/EE4END[13]
+ Tile_X3Y6_LUT4AB/EE4END[14] Tile_X3Y6_LUT4AB/EE4END[15] Tile_X3Y6_LUT4AB/EE4END[1]
+ Tile_X3Y6_LUT4AB/EE4END[2] Tile_X3Y6_LUT4AB/EE4END[3] Tile_X3Y6_LUT4AB/EE4END[4]
+ Tile_X3Y6_LUT4AB/EE4END[5] Tile_X3Y6_LUT4AB/EE4END[6] Tile_X3Y6_LUT4AB/EE4END[7]
+ Tile_X3Y6_LUT4AB/EE4END[8] Tile_X3Y6_LUT4AB/EE4END[9] Tile_X2Y6_LUT4AB/EE4END[0]
+ Tile_X2Y6_LUT4AB/EE4END[10] Tile_X2Y6_LUT4AB/EE4END[11] Tile_X2Y6_LUT4AB/EE4END[12]
+ Tile_X2Y6_LUT4AB/EE4END[13] Tile_X2Y6_LUT4AB/EE4END[14] Tile_X2Y6_LUT4AB/EE4END[15]
+ Tile_X2Y6_LUT4AB/EE4END[1] Tile_X2Y6_LUT4AB/EE4END[2] Tile_X2Y6_LUT4AB/EE4END[3]
+ Tile_X2Y6_LUT4AB/EE4END[4] Tile_X2Y6_LUT4AB/EE4END[5] Tile_X2Y6_LUT4AB/EE4END[6]
+ Tile_X2Y6_LUT4AB/EE4END[7] Tile_X2Y6_LUT4AB/EE4END[8] Tile_X2Y6_LUT4AB/EE4END[9]
+ Tile_X2Y6_LUT4AB/FrameData[0] Tile_X2Y6_LUT4AB/FrameData[10] Tile_X2Y6_LUT4AB/FrameData[11]
+ Tile_X2Y6_LUT4AB/FrameData[12] Tile_X2Y6_LUT4AB/FrameData[13] Tile_X2Y6_LUT4AB/FrameData[14]
+ Tile_X2Y6_LUT4AB/FrameData[15] Tile_X2Y6_LUT4AB/FrameData[16] Tile_X2Y6_LUT4AB/FrameData[17]
+ Tile_X2Y6_LUT4AB/FrameData[18] Tile_X2Y6_LUT4AB/FrameData[19] Tile_X2Y6_LUT4AB/FrameData[1]
+ Tile_X2Y6_LUT4AB/FrameData[20] Tile_X2Y6_LUT4AB/FrameData[21] Tile_X2Y6_LUT4AB/FrameData[22]
+ Tile_X2Y6_LUT4AB/FrameData[23] Tile_X2Y6_LUT4AB/FrameData[24] Tile_X2Y6_LUT4AB/FrameData[25]
+ Tile_X2Y6_LUT4AB/FrameData[26] Tile_X2Y6_LUT4AB/FrameData[27] Tile_X2Y6_LUT4AB/FrameData[28]
+ Tile_X2Y6_LUT4AB/FrameData[29] Tile_X2Y6_LUT4AB/FrameData[2] Tile_X2Y6_LUT4AB/FrameData[30]
+ Tile_X2Y6_LUT4AB/FrameData[31] Tile_X2Y6_LUT4AB/FrameData[3] Tile_X2Y6_LUT4AB/FrameData[4]
+ Tile_X2Y6_LUT4AB/FrameData[5] Tile_X2Y6_LUT4AB/FrameData[6] Tile_X2Y6_LUT4AB/FrameData[7]
+ Tile_X2Y6_LUT4AB/FrameData[8] Tile_X2Y6_LUT4AB/FrameData[9] Tile_X3Y6_LUT4AB/FrameData[0]
+ Tile_X3Y6_LUT4AB/FrameData[10] Tile_X3Y6_LUT4AB/FrameData[11] Tile_X3Y6_LUT4AB/FrameData[12]
+ Tile_X3Y6_LUT4AB/FrameData[13] Tile_X3Y6_LUT4AB/FrameData[14] Tile_X3Y6_LUT4AB/FrameData[15]
+ Tile_X3Y6_LUT4AB/FrameData[16] Tile_X3Y6_LUT4AB/FrameData[17] Tile_X3Y6_LUT4AB/FrameData[18]
+ Tile_X3Y6_LUT4AB/FrameData[19] Tile_X3Y6_LUT4AB/FrameData[1] Tile_X3Y6_LUT4AB/FrameData[20]
+ Tile_X3Y6_LUT4AB/FrameData[21] Tile_X3Y6_LUT4AB/FrameData[22] Tile_X3Y6_LUT4AB/FrameData[23]
+ Tile_X3Y6_LUT4AB/FrameData[24] Tile_X3Y6_LUT4AB/FrameData[25] Tile_X3Y6_LUT4AB/FrameData[26]
+ Tile_X3Y6_LUT4AB/FrameData[27] Tile_X3Y6_LUT4AB/FrameData[28] Tile_X3Y6_LUT4AB/FrameData[29]
+ Tile_X3Y6_LUT4AB/FrameData[2] Tile_X3Y6_LUT4AB/FrameData[30] Tile_X3Y6_LUT4AB/FrameData[31]
+ Tile_X3Y6_LUT4AB/FrameData[3] Tile_X3Y6_LUT4AB/FrameData[4] Tile_X3Y6_LUT4AB/FrameData[5]
+ Tile_X3Y6_LUT4AB/FrameData[6] Tile_X3Y6_LUT4AB/FrameData[7] Tile_X3Y6_LUT4AB/FrameData[8]
+ Tile_X3Y6_LUT4AB/FrameData[9] Tile_X2Y6_LUT4AB/FrameStrobe[0] Tile_X2Y6_LUT4AB/FrameStrobe[10]
+ Tile_X2Y6_LUT4AB/FrameStrobe[11] Tile_X2Y6_LUT4AB/FrameStrobe[12] Tile_X2Y6_LUT4AB/FrameStrobe[13]
+ Tile_X2Y6_LUT4AB/FrameStrobe[14] Tile_X2Y6_LUT4AB/FrameStrobe[15] Tile_X2Y6_LUT4AB/FrameStrobe[16]
+ Tile_X2Y6_LUT4AB/FrameStrobe[17] Tile_X2Y6_LUT4AB/FrameStrobe[18] Tile_X2Y6_LUT4AB/FrameStrobe[19]
+ Tile_X2Y6_LUT4AB/FrameStrobe[1] Tile_X2Y6_LUT4AB/FrameStrobe[2] Tile_X2Y6_LUT4AB/FrameStrobe[3]
+ Tile_X2Y6_LUT4AB/FrameStrobe[4] Tile_X2Y6_LUT4AB/FrameStrobe[5] Tile_X2Y6_LUT4AB/FrameStrobe[6]
+ Tile_X2Y6_LUT4AB/FrameStrobe[7] Tile_X2Y6_LUT4AB/FrameStrobe[8] Tile_X2Y6_LUT4AB/FrameStrobe[9]
+ Tile_X2Y5_LUT4AB/FrameStrobe[0] Tile_X2Y5_LUT4AB/FrameStrobe[10] Tile_X2Y5_LUT4AB/FrameStrobe[11]
+ Tile_X2Y5_LUT4AB/FrameStrobe[12] Tile_X2Y5_LUT4AB/FrameStrobe[13] Tile_X2Y5_LUT4AB/FrameStrobe[14]
+ Tile_X2Y5_LUT4AB/FrameStrobe[15] Tile_X2Y5_LUT4AB/FrameStrobe[16] Tile_X2Y5_LUT4AB/FrameStrobe[17]
+ Tile_X2Y5_LUT4AB/FrameStrobe[18] Tile_X2Y5_LUT4AB/FrameStrobe[19] Tile_X2Y5_LUT4AB/FrameStrobe[1]
+ Tile_X2Y5_LUT4AB/FrameStrobe[2] Tile_X2Y5_LUT4AB/FrameStrobe[3] Tile_X2Y5_LUT4AB/FrameStrobe[4]
+ Tile_X2Y5_LUT4AB/FrameStrobe[5] Tile_X2Y5_LUT4AB/FrameStrobe[6] Tile_X2Y5_LUT4AB/FrameStrobe[7]
+ Tile_X2Y5_LUT4AB/FrameStrobe[8] Tile_X2Y5_LUT4AB/FrameStrobe[9] Tile_X2Y6_LUT4AB/N1BEG[0]
+ Tile_X2Y6_LUT4AB/N1BEG[1] Tile_X2Y6_LUT4AB/N1BEG[2] Tile_X2Y6_LUT4AB/N1BEG[3] Tile_X2Y7_LUT4AB/N1BEG[0]
+ Tile_X2Y7_LUT4AB/N1BEG[1] Tile_X2Y7_LUT4AB/N1BEG[2] Tile_X2Y7_LUT4AB/N1BEG[3] Tile_X2Y6_LUT4AB/N2BEG[0]
+ Tile_X2Y6_LUT4AB/N2BEG[1] Tile_X2Y6_LUT4AB/N2BEG[2] Tile_X2Y6_LUT4AB/N2BEG[3] Tile_X2Y6_LUT4AB/N2BEG[4]
+ Tile_X2Y6_LUT4AB/N2BEG[5] Tile_X2Y6_LUT4AB/N2BEG[6] Tile_X2Y6_LUT4AB/N2BEG[7] Tile_X2Y5_LUT4AB/N2END[0]
+ Tile_X2Y5_LUT4AB/N2END[1] Tile_X2Y5_LUT4AB/N2END[2] Tile_X2Y5_LUT4AB/N2END[3] Tile_X2Y5_LUT4AB/N2END[4]
+ Tile_X2Y5_LUT4AB/N2END[5] Tile_X2Y5_LUT4AB/N2END[6] Tile_X2Y5_LUT4AB/N2END[7] Tile_X2Y6_LUT4AB/N2END[0]
+ Tile_X2Y6_LUT4AB/N2END[1] Tile_X2Y6_LUT4AB/N2END[2] Tile_X2Y6_LUT4AB/N2END[3] Tile_X2Y6_LUT4AB/N2END[4]
+ Tile_X2Y6_LUT4AB/N2END[5] Tile_X2Y6_LUT4AB/N2END[6] Tile_X2Y6_LUT4AB/N2END[7] Tile_X2Y7_LUT4AB/N2BEG[0]
+ Tile_X2Y7_LUT4AB/N2BEG[1] Tile_X2Y7_LUT4AB/N2BEG[2] Tile_X2Y7_LUT4AB/N2BEG[3] Tile_X2Y7_LUT4AB/N2BEG[4]
+ Tile_X2Y7_LUT4AB/N2BEG[5] Tile_X2Y7_LUT4AB/N2BEG[6] Tile_X2Y7_LUT4AB/N2BEG[7] Tile_X2Y6_LUT4AB/N4BEG[0]
+ Tile_X2Y6_LUT4AB/N4BEG[10] Tile_X2Y6_LUT4AB/N4BEG[11] Tile_X2Y6_LUT4AB/N4BEG[12]
+ Tile_X2Y6_LUT4AB/N4BEG[13] Tile_X2Y6_LUT4AB/N4BEG[14] Tile_X2Y6_LUT4AB/N4BEG[15]
+ Tile_X2Y6_LUT4AB/N4BEG[1] Tile_X2Y6_LUT4AB/N4BEG[2] Tile_X2Y6_LUT4AB/N4BEG[3] Tile_X2Y6_LUT4AB/N4BEG[4]
+ Tile_X2Y6_LUT4AB/N4BEG[5] Tile_X2Y6_LUT4AB/N4BEG[6] Tile_X2Y6_LUT4AB/N4BEG[7] Tile_X2Y6_LUT4AB/N4BEG[8]
+ Tile_X2Y6_LUT4AB/N4BEG[9] Tile_X2Y7_LUT4AB/N4BEG[0] Tile_X2Y7_LUT4AB/N4BEG[10] Tile_X2Y7_LUT4AB/N4BEG[11]
+ Tile_X2Y7_LUT4AB/N4BEG[12] Tile_X2Y7_LUT4AB/N4BEG[13] Tile_X2Y7_LUT4AB/N4BEG[14]
+ Tile_X2Y7_LUT4AB/N4BEG[15] Tile_X2Y7_LUT4AB/N4BEG[1] Tile_X2Y7_LUT4AB/N4BEG[2] Tile_X2Y7_LUT4AB/N4BEG[3]
+ Tile_X2Y7_LUT4AB/N4BEG[4] Tile_X2Y7_LUT4AB/N4BEG[5] Tile_X2Y7_LUT4AB/N4BEG[6] Tile_X2Y7_LUT4AB/N4BEG[7]
+ Tile_X2Y7_LUT4AB/N4BEG[8] Tile_X2Y7_LUT4AB/N4BEG[9] Tile_X2Y6_LUT4AB/NN4BEG[0] Tile_X2Y6_LUT4AB/NN4BEG[10]
+ Tile_X2Y6_LUT4AB/NN4BEG[11] Tile_X2Y6_LUT4AB/NN4BEG[12] Tile_X2Y6_LUT4AB/NN4BEG[13]
+ Tile_X2Y6_LUT4AB/NN4BEG[14] Tile_X2Y6_LUT4AB/NN4BEG[15] Tile_X2Y6_LUT4AB/NN4BEG[1]
+ Tile_X2Y6_LUT4AB/NN4BEG[2] Tile_X2Y6_LUT4AB/NN4BEG[3] Tile_X2Y6_LUT4AB/NN4BEG[4]
+ Tile_X2Y6_LUT4AB/NN4BEG[5] Tile_X2Y6_LUT4AB/NN4BEG[6] Tile_X2Y6_LUT4AB/NN4BEG[7]
+ Tile_X2Y6_LUT4AB/NN4BEG[8] Tile_X2Y6_LUT4AB/NN4BEG[9] Tile_X2Y7_LUT4AB/NN4BEG[0]
+ Tile_X2Y7_LUT4AB/NN4BEG[10] Tile_X2Y7_LUT4AB/NN4BEG[11] Tile_X2Y7_LUT4AB/NN4BEG[12]
+ Tile_X2Y7_LUT4AB/NN4BEG[13] Tile_X2Y7_LUT4AB/NN4BEG[14] Tile_X2Y7_LUT4AB/NN4BEG[15]
+ Tile_X2Y7_LUT4AB/NN4BEG[1] Tile_X2Y7_LUT4AB/NN4BEG[2] Tile_X2Y7_LUT4AB/NN4BEG[3]
+ Tile_X2Y7_LUT4AB/NN4BEG[4] Tile_X2Y7_LUT4AB/NN4BEG[5] Tile_X2Y7_LUT4AB/NN4BEG[6]
+ Tile_X2Y7_LUT4AB/NN4BEG[7] Tile_X2Y7_LUT4AB/NN4BEG[8] Tile_X2Y7_LUT4AB/NN4BEG[9]
+ Tile_X2Y7_LUT4AB/S1END[0] Tile_X2Y7_LUT4AB/S1END[1] Tile_X2Y7_LUT4AB/S1END[2] Tile_X2Y7_LUT4AB/S1END[3]
+ Tile_X2Y6_LUT4AB/S1END[0] Tile_X2Y6_LUT4AB/S1END[1] Tile_X2Y6_LUT4AB/S1END[2] Tile_X2Y6_LUT4AB/S1END[3]
+ Tile_X2Y7_LUT4AB/S2MID[0] Tile_X2Y7_LUT4AB/S2MID[1] Tile_X2Y7_LUT4AB/S2MID[2] Tile_X2Y7_LUT4AB/S2MID[3]
+ Tile_X2Y7_LUT4AB/S2MID[4] Tile_X2Y7_LUT4AB/S2MID[5] Tile_X2Y7_LUT4AB/S2MID[6] Tile_X2Y7_LUT4AB/S2MID[7]
+ Tile_X2Y7_LUT4AB/S2END[0] Tile_X2Y7_LUT4AB/S2END[1] Tile_X2Y7_LUT4AB/S2END[2] Tile_X2Y7_LUT4AB/S2END[3]
+ Tile_X2Y7_LUT4AB/S2END[4] Tile_X2Y7_LUT4AB/S2END[5] Tile_X2Y7_LUT4AB/S2END[6] Tile_X2Y7_LUT4AB/S2END[7]
+ Tile_X2Y6_LUT4AB/S2END[0] Tile_X2Y6_LUT4AB/S2END[1] Tile_X2Y6_LUT4AB/S2END[2] Tile_X2Y6_LUT4AB/S2END[3]
+ Tile_X2Y6_LUT4AB/S2END[4] Tile_X2Y6_LUT4AB/S2END[5] Tile_X2Y6_LUT4AB/S2END[6] Tile_X2Y6_LUT4AB/S2END[7]
+ Tile_X2Y6_LUT4AB/S2MID[0] Tile_X2Y6_LUT4AB/S2MID[1] Tile_X2Y6_LUT4AB/S2MID[2] Tile_X2Y6_LUT4AB/S2MID[3]
+ Tile_X2Y6_LUT4AB/S2MID[4] Tile_X2Y6_LUT4AB/S2MID[5] Tile_X2Y6_LUT4AB/S2MID[6] Tile_X2Y6_LUT4AB/S2MID[7]
+ Tile_X2Y7_LUT4AB/S4END[0] Tile_X2Y7_LUT4AB/S4END[10] Tile_X2Y7_LUT4AB/S4END[11]
+ Tile_X2Y7_LUT4AB/S4END[12] Tile_X2Y7_LUT4AB/S4END[13] Tile_X2Y7_LUT4AB/S4END[14]
+ Tile_X2Y7_LUT4AB/S4END[15] Tile_X2Y7_LUT4AB/S4END[1] Tile_X2Y7_LUT4AB/S4END[2] Tile_X2Y7_LUT4AB/S4END[3]
+ Tile_X2Y7_LUT4AB/S4END[4] Tile_X2Y7_LUT4AB/S4END[5] Tile_X2Y7_LUT4AB/S4END[6] Tile_X2Y7_LUT4AB/S4END[7]
+ Tile_X2Y7_LUT4AB/S4END[8] Tile_X2Y7_LUT4AB/S4END[9] Tile_X2Y6_LUT4AB/S4END[0] Tile_X2Y6_LUT4AB/S4END[10]
+ Tile_X2Y6_LUT4AB/S4END[11] Tile_X2Y6_LUT4AB/S4END[12] Tile_X2Y6_LUT4AB/S4END[13]
+ Tile_X2Y6_LUT4AB/S4END[14] Tile_X2Y6_LUT4AB/S4END[15] Tile_X2Y6_LUT4AB/S4END[1]
+ Tile_X2Y6_LUT4AB/S4END[2] Tile_X2Y6_LUT4AB/S4END[3] Tile_X2Y6_LUT4AB/S4END[4] Tile_X2Y6_LUT4AB/S4END[5]
+ Tile_X2Y6_LUT4AB/S4END[6] Tile_X2Y6_LUT4AB/S4END[7] Tile_X2Y6_LUT4AB/S4END[8] Tile_X2Y6_LUT4AB/S4END[9]
+ Tile_X2Y7_LUT4AB/SS4END[0] Tile_X2Y7_LUT4AB/SS4END[10] Tile_X2Y7_LUT4AB/SS4END[11]
+ Tile_X2Y7_LUT4AB/SS4END[12] Tile_X2Y7_LUT4AB/SS4END[13] Tile_X2Y7_LUT4AB/SS4END[14]
+ Tile_X2Y7_LUT4AB/SS4END[15] Tile_X2Y7_LUT4AB/SS4END[1] Tile_X2Y7_LUT4AB/SS4END[2]
+ Tile_X2Y7_LUT4AB/SS4END[3] Tile_X2Y7_LUT4AB/SS4END[4] Tile_X2Y7_LUT4AB/SS4END[5]
+ Tile_X2Y7_LUT4AB/SS4END[6] Tile_X2Y7_LUT4AB/SS4END[7] Tile_X2Y7_LUT4AB/SS4END[8]
+ Tile_X2Y7_LUT4AB/SS4END[9] Tile_X2Y6_LUT4AB/SS4END[0] Tile_X2Y6_LUT4AB/SS4END[10]
+ Tile_X2Y6_LUT4AB/SS4END[11] Tile_X2Y6_LUT4AB/SS4END[12] Tile_X2Y6_LUT4AB/SS4END[13]
+ Tile_X2Y6_LUT4AB/SS4END[14] Tile_X2Y6_LUT4AB/SS4END[15] Tile_X2Y6_LUT4AB/SS4END[1]
+ Tile_X2Y6_LUT4AB/SS4END[2] Tile_X2Y6_LUT4AB/SS4END[3] Tile_X2Y6_LUT4AB/SS4END[4]
+ Tile_X2Y6_LUT4AB/SS4END[5] Tile_X2Y6_LUT4AB/SS4END[6] Tile_X2Y6_LUT4AB/SS4END[7]
+ Tile_X2Y6_LUT4AB/SS4END[8] Tile_X2Y6_LUT4AB/SS4END[9] Tile_X2Y6_LUT4AB/UserCLK Tile_X2Y5_LUT4AB/UserCLK
+ VGND VPWR Tile_X2Y6_LUT4AB/W1BEG[0] Tile_X2Y6_LUT4AB/W1BEG[1] Tile_X2Y6_LUT4AB/W1BEG[2]
+ Tile_X2Y6_LUT4AB/W1BEG[3] Tile_X3Y6_LUT4AB/W1BEG[0] Tile_X3Y6_LUT4AB/W1BEG[1] Tile_X3Y6_LUT4AB/W1BEG[2]
+ Tile_X3Y6_LUT4AB/W1BEG[3] Tile_X2Y6_LUT4AB/W2BEG[0] Tile_X2Y6_LUT4AB/W2BEG[1] Tile_X2Y6_LUT4AB/W2BEG[2]
+ Tile_X2Y6_LUT4AB/W2BEG[3] Tile_X2Y6_LUT4AB/W2BEG[4] Tile_X2Y6_LUT4AB/W2BEG[5] Tile_X2Y6_LUT4AB/W2BEG[6]
+ Tile_X2Y6_LUT4AB/W2BEG[7] Tile_X1Y6_LUT4AB/W2END[0] Tile_X1Y6_LUT4AB/W2END[1] Tile_X1Y6_LUT4AB/W2END[2]
+ Tile_X1Y6_LUT4AB/W2END[3] Tile_X1Y6_LUT4AB/W2END[4] Tile_X1Y6_LUT4AB/W2END[5] Tile_X1Y6_LUT4AB/W2END[6]
+ Tile_X1Y6_LUT4AB/W2END[7] Tile_X2Y6_LUT4AB/W2END[0] Tile_X2Y6_LUT4AB/W2END[1] Tile_X2Y6_LUT4AB/W2END[2]
+ Tile_X2Y6_LUT4AB/W2END[3] Tile_X2Y6_LUT4AB/W2END[4] Tile_X2Y6_LUT4AB/W2END[5] Tile_X2Y6_LUT4AB/W2END[6]
+ Tile_X2Y6_LUT4AB/W2END[7] Tile_X3Y6_LUT4AB/W2BEG[0] Tile_X3Y6_LUT4AB/W2BEG[1] Tile_X3Y6_LUT4AB/W2BEG[2]
+ Tile_X3Y6_LUT4AB/W2BEG[3] Tile_X3Y6_LUT4AB/W2BEG[4] Tile_X3Y6_LUT4AB/W2BEG[5] Tile_X3Y6_LUT4AB/W2BEG[6]
+ Tile_X3Y6_LUT4AB/W2BEG[7] Tile_X2Y6_LUT4AB/W6BEG[0] Tile_X2Y6_LUT4AB/W6BEG[10] Tile_X2Y6_LUT4AB/W6BEG[11]
+ Tile_X2Y6_LUT4AB/W6BEG[1] Tile_X2Y6_LUT4AB/W6BEG[2] Tile_X2Y6_LUT4AB/W6BEG[3] Tile_X2Y6_LUT4AB/W6BEG[4]
+ Tile_X2Y6_LUT4AB/W6BEG[5] Tile_X2Y6_LUT4AB/W6BEG[6] Tile_X2Y6_LUT4AB/W6BEG[7] Tile_X2Y6_LUT4AB/W6BEG[8]
+ Tile_X2Y6_LUT4AB/W6BEG[9] Tile_X3Y6_LUT4AB/W6BEG[0] Tile_X3Y6_LUT4AB/W6BEG[10] Tile_X3Y6_LUT4AB/W6BEG[11]
+ Tile_X3Y6_LUT4AB/W6BEG[1] Tile_X3Y6_LUT4AB/W6BEG[2] Tile_X3Y6_LUT4AB/W6BEG[3] Tile_X3Y6_LUT4AB/W6BEG[4]
+ Tile_X3Y6_LUT4AB/W6BEG[5] Tile_X3Y6_LUT4AB/W6BEG[6] Tile_X3Y6_LUT4AB/W6BEG[7] Tile_X3Y6_LUT4AB/W6BEG[8]
+ Tile_X3Y6_LUT4AB/W6BEG[9] Tile_X2Y6_LUT4AB/WW4BEG[0] Tile_X2Y6_LUT4AB/WW4BEG[10]
+ Tile_X2Y6_LUT4AB/WW4BEG[11] Tile_X2Y6_LUT4AB/WW4BEG[12] Tile_X2Y6_LUT4AB/WW4BEG[13]
+ Tile_X2Y6_LUT4AB/WW4BEG[14] Tile_X2Y6_LUT4AB/WW4BEG[15] Tile_X2Y6_LUT4AB/WW4BEG[1]
+ Tile_X2Y6_LUT4AB/WW4BEG[2] Tile_X2Y6_LUT4AB/WW4BEG[3] Tile_X2Y6_LUT4AB/WW4BEG[4]
+ Tile_X2Y6_LUT4AB/WW4BEG[5] Tile_X2Y6_LUT4AB/WW4BEG[6] Tile_X2Y6_LUT4AB/WW4BEG[7]
+ Tile_X2Y6_LUT4AB/WW4BEG[8] Tile_X2Y6_LUT4AB/WW4BEG[9] Tile_X3Y6_LUT4AB/WW4BEG[0]
+ Tile_X3Y6_LUT4AB/WW4BEG[10] Tile_X3Y6_LUT4AB/WW4BEG[11] Tile_X3Y6_LUT4AB/WW4BEG[12]
+ Tile_X3Y6_LUT4AB/WW4BEG[13] Tile_X3Y6_LUT4AB/WW4BEG[14] Tile_X3Y6_LUT4AB/WW4BEG[15]
+ Tile_X3Y6_LUT4AB/WW4BEG[1] Tile_X3Y6_LUT4AB/WW4BEG[2] Tile_X3Y6_LUT4AB/WW4BEG[3]
+ Tile_X3Y6_LUT4AB/WW4BEG[4] Tile_X3Y6_LUT4AB/WW4BEG[5] Tile_X3Y6_LUT4AB/WW4BEG[6]
+ Tile_X3Y6_LUT4AB/WW4BEG[7] Tile_X3Y6_LUT4AB/WW4BEG[8] Tile_X3Y6_LUT4AB/WW4BEG[9]
+ LUT4AB
XTile_X5Y0_NE_term Tile_X5Y0_NE_term/FrameData[0] Tile_X5Y0_NE_term/FrameData[10]
+ Tile_X5Y0_NE_term/FrameData[11] Tile_X5Y0_NE_term/FrameData[12] Tile_X5Y0_NE_term/FrameData[13]
+ Tile_X5Y0_NE_term/FrameData[14] Tile_X5Y0_NE_term/FrameData[15] Tile_X5Y0_NE_term/FrameData[16]
+ Tile_X5Y0_NE_term/FrameData[17] Tile_X5Y0_NE_term/FrameData[18] Tile_X5Y0_NE_term/FrameData[19]
+ Tile_X5Y0_NE_term/FrameData[1] Tile_X5Y0_NE_term/FrameData[20] Tile_X5Y0_NE_term/FrameData[21]
+ Tile_X5Y0_NE_term/FrameData[22] Tile_X5Y0_NE_term/FrameData[23] Tile_X5Y0_NE_term/FrameData[24]
+ Tile_X5Y0_NE_term/FrameData[25] Tile_X5Y0_NE_term/FrameData[26] Tile_X5Y0_NE_term/FrameData[27]
+ Tile_X5Y0_NE_term/FrameData[28] Tile_X5Y0_NE_term/FrameData[29] Tile_X5Y0_NE_term/FrameData[2]
+ Tile_X5Y0_NE_term/FrameData[30] Tile_X5Y0_NE_term/FrameData[31] Tile_X5Y0_NE_term/FrameData[3]
+ Tile_X5Y0_NE_term/FrameData[4] Tile_X5Y0_NE_term/FrameData[5] Tile_X5Y0_NE_term/FrameData[6]
+ Tile_X5Y0_NE_term/FrameData[7] Tile_X5Y0_NE_term/FrameData[8] Tile_X5Y0_NE_term/FrameData[9]
+ Tile_X5Y0_NE_term/FrameData_O[0] Tile_X5Y0_NE_term/FrameData_O[10] Tile_X5Y0_NE_term/FrameData_O[11]
+ Tile_X5Y0_NE_term/FrameData_O[12] Tile_X5Y0_NE_term/FrameData_O[13] Tile_X5Y0_NE_term/FrameData_O[14]
+ Tile_X5Y0_NE_term/FrameData_O[15] Tile_X5Y0_NE_term/FrameData_O[16] Tile_X5Y0_NE_term/FrameData_O[17]
+ Tile_X5Y0_NE_term/FrameData_O[18] Tile_X5Y0_NE_term/FrameData_O[19] Tile_X5Y0_NE_term/FrameData_O[1]
+ Tile_X5Y0_NE_term/FrameData_O[20] Tile_X5Y0_NE_term/FrameData_O[21] Tile_X5Y0_NE_term/FrameData_O[22]
+ Tile_X5Y0_NE_term/FrameData_O[23] Tile_X5Y0_NE_term/FrameData_O[24] Tile_X5Y0_NE_term/FrameData_O[25]
+ Tile_X5Y0_NE_term/FrameData_O[26] Tile_X5Y0_NE_term/FrameData_O[27] Tile_X5Y0_NE_term/FrameData_O[28]
+ Tile_X5Y0_NE_term/FrameData_O[29] Tile_X5Y0_NE_term/FrameData_O[2] Tile_X5Y0_NE_term/FrameData_O[30]
+ Tile_X5Y0_NE_term/FrameData_O[31] Tile_X5Y0_NE_term/FrameData_O[3] Tile_X5Y0_NE_term/FrameData_O[4]
+ Tile_X5Y0_NE_term/FrameData_O[5] Tile_X5Y0_NE_term/FrameData_O[6] Tile_X5Y0_NE_term/FrameData_O[7]
+ Tile_X5Y0_NE_term/FrameData_O[8] Tile_X5Y0_NE_term/FrameData_O[9] Tile_X5Y0_NE_term/FrameStrobe[0]
+ Tile_X5Y0_NE_term/FrameStrobe[10] Tile_X5Y0_NE_term/FrameStrobe[11] Tile_X5Y0_NE_term/FrameStrobe[12]
+ Tile_X5Y0_NE_term/FrameStrobe[13] Tile_X5Y0_NE_term/FrameStrobe[14] Tile_X5Y0_NE_term/FrameStrobe[15]
+ Tile_X5Y0_NE_term/FrameStrobe[16] Tile_X5Y0_NE_term/FrameStrobe[17] Tile_X5Y0_NE_term/FrameStrobe[18]
+ Tile_X5Y0_NE_term/FrameStrobe[19] Tile_X5Y0_NE_term/FrameStrobe[1] Tile_X5Y0_NE_term/FrameStrobe[2]
+ Tile_X5Y0_NE_term/FrameStrobe[3] Tile_X5Y0_NE_term/FrameStrobe[4] Tile_X5Y0_NE_term/FrameStrobe[5]
+ Tile_X5Y0_NE_term/FrameStrobe[6] Tile_X5Y0_NE_term/FrameStrobe[7] Tile_X5Y0_NE_term/FrameStrobe[8]
+ Tile_X5Y0_NE_term/FrameStrobe[9] Tile_X5Y0_NE_term/FrameStrobe_O[0] Tile_X5Y0_NE_term/FrameStrobe_O[10]
+ Tile_X5Y0_NE_term/FrameStrobe_O[11] Tile_X5Y0_NE_term/FrameStrobe_O[12] Tile_X5Y0_NE_term/FrameStrobe_O[13]
+ Tile_X5Y0_NE_term/FrameStrobe_O[14] Tile_X5Y0_NE_term/FrameStrobe_O[15] Tile_X5Y0_NE_term/FrameStrobe_O[16]
+ Tile_X5Y0_NE_term/FrameStrobe_O[17] Tile_X5Y0_NE_term/FrameStrobe_O[18] Tile_X5Y0_NE_term/FrameStrobe_O[19]
+ Tile_X5Y0_NE_term/FrameStrobe_O[1] Tile_X5Y0_NE_term/FrameStrobe_O[2] Tile_X5Y0_NE_term/FrameStrobe_O[3]
+ Tile_X5Y0_NE_term/FrameStrobe_O[4] Tile_X5Y0_NE_term/FrameStrobe_O[5] Tile_X5Y0_NE_term/FrameStrobe_O[6]
+ Tile_X5Y0_NE_term/FrameStrobe_O[7] Tile_X5Y0_NE_term/FrameStrobe_O[8] Tile_X5Y0_NE_term/FrameStrobe_O[9]
+ Tile_X5Y0_NE_term/N1END[0] Tile_X5Y0_NE_term/N1END[1] Tile_X5Y0_NE_term/N1END[2]
+ Tile_X5Y0_NE_term/N1END[3] Tile_X5Y0_NE_term/N2END[0] Tile_X5Y0_NE_term/N2END[1]
+ Tile_X5Y0_NE_term/N2END[2] Tile_X5Y0_NE_term/N2END[3] Tile_X5Y0_NE_term/N2END[4]
+ Tile_X5Y0_NE_term/N2END[5] Tile_X5Y0_NE_term/N2END[6] Tile_X5Y0_NE_term/N2END[7]
+ Tile_X5Y0_NE_term/N2MID[0] Tile_X5Y0_NE_term/N2MID[1] Tile_X5Y0_NE_term/N2MID[2]
+ Tile_X5Y0_NE_term/N2MID[3] Tile_X5Y0_NE_term/N2MID[4] Tile_X5Y0_NE_term/N2MID[5]
+ Tile_X5Y0_NE_term/N2MID[6] Tile_X5Y0_NE_term/N2MID[7] Tile_X5Y0_NE_term/N4END[0]
+ Tile_X5Y0_NE_term/N4END[10] Tile_X5Y0_NE_term/N4END[11] Tile_X5Y0_NE_term/N4END[12]
+ Tile_X5Y0_NE_term/N4END[13] Tile_X5Y0_NE_term/N4END[14] Tile_X5Y0_NE_term/N4END[15]
+ Tile_X5Y0_NE_term/N4END[1] Tile_X5Y0_NE_term/N4END[2] Tile_X5Y0_NE_term/N4END[3]
+ Tile_X5Y0_NE_term/N4END[4] Tile_X5Y0_NE_term/N4END[5] Tile_X5Y0_NE_term/N4END[6]
+ Tile_X5Y0_NE_term/N4END[7] Tile_X5Y0_NE_term/N4END[8] Tile_X5Y0_NE_term/N4END[9]
+ Tile_X5Y0_NE_term/S1BEG[0] Tile_X5Y0_NE_term/S1BEG[1] Tile_X5Y0_NE_term/S1BEG[2]
+ Tile_X5Y0_NE_term/S1BEG[3] Tile_X5Y0_NE_term/S2BEG[0] Tile_X5Y0_NE_term/S2BEG[1]
+ Tile_X5Y0_NE_term/S2BEG[2] Tile_X5Y0_NE_term/S2BEG[3] Tile_X5Y0_NE_term/S2BEG[4]
+ Tile_X5Y0_NE_term/S2BEG[5] Tile_X5Y0_NE_term/S2BEG[6] Tile_X5Y0_NE_term/S2BEG[7]
+ Tile_X5Y0_NE_term/S2BEGb[0] Tile_X5Y0_NE_term/S2BEGb[1] Tile_X5Y0_NE_term/S2BEGb[2]
+ Tile_X5Y0_NE_term/S2BEGb[3] Tile_X5Y0_NE_term/S2BEGb[4] Tile_X5Y0_NE_term/S2BEGb[5]
+ Tile_X5Y0_NE_term/S2BEGb[6] Tile_X5Y0_NE_term/S2BEGb[7] Tile_X5Y0_NE_term/S4BEG[0]
+ Tile_X5Y0_NE_term/S4BEG[10] Tile_X5Y0_NE_term/S4BEG[11] Tile_X5Y0_NE_term/S4BEG[12]
+ Tile_X5Y0_NE_term/S4BEG[13] Tile_X5Y0_NE_term/S4BEG[14] Tile_X5Y0_NE_term/S4BEG[15]
+ Tile_X5Y0_NE_term/S4BEG[1] Tile_X5Y0_NE_term/S4BEG[2] Tile_X5Y0_NE_term/S4BEG[3]
+ Tile_X5Y0_NE_term/S4BEG[4] Tile_X5Y0_NE_term/S4BEG[5] Tile_X5Y0_NE_term/S4BEG[6]
+ Tile_X5Y0_NE_term/S4BEG[7] Tile_X5Y0_NE_term/S4BEG[8] Tile_X5Y0_NE_term/S4BEG[9]
+ Tile_X5Y0_NE_term/UserCLK Tile_X5Y0_NE_term/UserCLKo VGND VPWR NE_term
XTile_X4Y9_S_IO4 Tile_X4Y9_A_I_top Tile_X4Y9_A_O_top Tile_X4Y9_A_T_top Tile_X4Y9_B_I_top
+ Tile_X4Y9_B_O_top Tile_X4Y9_B_T_top Tile_X4Y9_C_I_top Tile_X4Y9_C_O_top Tile_X4Y9_C_T_top
+ Tile_X4Y9_S_IO4/Co Tile_X4Y9_D_I_top Tile_X4Y9_D_O_top Tile_X4Y9_D_T_top Tile_X4Y9_S_IO4/FrameData[0]
+ Tile_X4Y9_S_IO4/FrameData[10] Tile_X4Y9_S_IO4/FrameData[11] Tile_X4Y9_S_IO4/FrameData[12]
+ Tile_X4Y9_S_IO4/FrameData[13] Tile_X4Y9_S_IO4/FrameData[14] Tile_X4Y9_S_IO4/FrameData[15]
+ Tile_X4Y9_S_IO4/FrameData[16] Tile_X4Y9_S_IO4/FrameData[17] Tile_X4Y9_S_IO4/FrameData[18]
+ Tile_X4Y9_S_IO4/FrameData[19] Tile_X4Y9_S_IO4/FrameData[1] Tile_X4Y9_S_IO4/FrameData[20]
+ Tile_X4Y9_S_IO4/FrameData[21] Tile_X4Y9_S_IO4/FrameData[22] Tile_X4Y9_S_IO4/FrameData[23]
+ Tile_X4Y9_S_IO4/FrameData[24] Tile_X4Y9_S_IO4/FrameData[25] Tile_X4Y9_S_IO4/FrameData[26]
+ Tile_X4Y9_S_IO4/FrameData[27] Tile_X4Y9_S_IO4/FrameData[28] Tile_X4Y9_S_IO4/FrameData[29]
+ Tile_X4Y9_S_IO4/FrameData[2] Tile_X4Y9_S_IO4/FrameData[30] Tile_X4Y9_S_IO4/FrameData[31]
+ Tile_X4Y9_S_IO4/FrameData[3] Tile_X4Y9_S_IO4/FrameData[4] Tile_X4Y9_S_IO4/FrameData[5]
+ Tile_X4Y9_S_IO4/FrameData[6] Tile_X4Y9_S_IO4/FrameData[7] Tile_X4Y9_S_IO4/FrameData[8]
+ Tile_X4Y9_S_IO4/FrameData[9] Tile_X5Y9_SE_term/FrameData[0] Tile_X5Y9_SE_term/FrameData[10]
+ Tile_X5Y9_SE_term/FrameData[11] Tile_X5Y9_SE_term/FrameData[12] Tile_X5Y9_SE_term/FrameData[13]
+ Tile_X5Y9_SE_term/FrameData[14] Tile_X5Y9_SE_term/FrameData[15] Tile_X5Y9_SE_term/FrameData[16]
+ Tile_X5Y9_SE_term/FrameData[17] Tile_X5Y9_SE_term/FrameData[18] Tile_X5Y9_SE_term/FrameData[19]
+ Tile_X5Y9_SE_term/FrameData[1] Tile_X5Y9_SE_term/FrameData[20] Tile_X5Y9_SE_term/FrameData[21]
+ Tile_X5Y9_SE_term/FrameData[22] Tile_X5Y9_SE_term/FrameData[23] Tile_X5Y9_SE_term/FrameData[24]
+ Tile_X5Y9_SE_term/FrameData[25] Tile_X5Y9_SE_term/FrameData[26] Tile_X5Y9_SE_term/FrameData[27]
+ Tile_X5Y9_SE_term/FrameData[28] Tile_X5Y9_SE_term/FrameData[29] Tile_X5Y9_SE_term/FrameData[2]
+ Tile_X5Y9_SE_term/FrameData[30] Tile_X5Y9_SE_term/FrameData[31] Tile_X5Y9_SE_term/FrameData[3]
+ Tile_X5Y9_SE_term/FrameData[4] Tile_X5Y9_SE_term/FrameData[5] Tile_X5Y9_SE_term/FrameData[6]
+ Tile_X5Y9_SE_term/FrameData[7] Tile_X5Y9_SE_term/FrameData[8] Tile_X5Y9_SE_term/FrameData[9]
+ FrameStrobe[80] FrameStrobe[90] FrameStrobe[91] FrameStrobe[92] FrameStrobe[93]
+ FrameStrobe[94] FrameStrobe[95] FrameStrobe[96] FrameStrobe[97] FrameStrobe[98]
+ FrameStrobe[99] FrameStrobe[81] FrameStrobe[82] FrameStrobe[83] FrameStrobe[84]
+ FrameStrobe[85] FrameStrobe[86] FrameStrobe[87] FrameStrobe[88] FrameStrobe[89]
+ Tile_X4Y8_LUT4AB/FrameStrobe[0] Tile_X4Y8_LUT4AB/FrameStrobe[10] Tile_X4Y8_LUT4AB/FrameStrobe[11]
+ Tile_X4Y8_LUT4AB/FrameStrobe[12] Tile_X4Y8_LUT4AB/FrameStrobe[13] Tile_X4Y8_LUT4AB/FrameStrobe[14]
+ Tile_X4Y8_LUT4AB/FrameStrobe[15] Tile_X4Y8_LUT4AB/FrameStrobe[16] Tile_X4Y8_LUT4AB/FrameStrobe[17]
+ Tile_X4Y8_LUT4AB/FrameStrobe[18] Tile_X4Y8_LUT4AB/FrameStrobe[19] Tile_X4Y8_LUT4AB/FrameStrobe[1]
+ Tile_X4Y8_LUT4AB/FrameStrobe[2] Tile_X4Y8_LUT4AB/FrameStrobe[3] Tile_X4Y8_LUT4AB/FrameStrobe[4]
+ Tile_X4Y8_LUT4AB/FrameStrobe[5] Tile_X4Y8_LUT4AB/FrameStrobe[6] Tile_X4Y8_LUT4AB/FrameStrobe[7]
+ Tile_X4Y8_LUT4AB/FrameStrobe[8] Tile_X4Y8_LUT4AB/FrameStrobe[9] Tile_X4Y9_S_IO4/N1BEG[0]
+ Tile_X4Y9_S_IO4/N1BEG[1] Tile_X4Y9_S_IO4/N1BEG[2] Tile_X4Y9_S_IO4/N1BEG[3] Tile_X4Y9_S_IO4/N2BEG[0]
+ Tile_X4Y9_S_IO4/N2BEG[1] Tile_X4Y9_S_IO4/N2BEG[2] Tile_X4Y9_S_IO4/N2BEG[3] Tile_X4Y9_S_IO4/N2BEG[4]
+ Tile_X4Y9_S_IO4/N2BEG[5] Tile_X4Y9_S_IO4/N2BEG[6] Tile_X4Y9_S_IO4/N2BEG[7] Tile_X4Y9_S_IO4/N2BEGb[0]
+ Tile_X4Y9_S_IO4/N2BEGb[1] Tile_X4Y9_S_IO4/N2BEGb[2] Tile_X4Y9_S_IO4/N2BEGb[3] Tile_X4Y9_S_IO4/N2BEGb[4]
+ Tile_X4Y9_S_IO4/N2BEGb[5] Tile_X4Y9_S_IO4/N2BEGb[6] Tile_X4Y9_S_IO4/N2BEGb[7] Tile_X4Y9_S_IO4/N4BEG[0]
+ Tile_X4Y9_S_IO4/N4BEG[10] Tile_X4Y9_S_IO4/N4BEG[11] Tile_X4Y9_S_IO4/N4BEG[12] Tile_X4Y9_S_IO4/N4BEG[13]
+ Tile_X4Y9_S_IO4/N4BEG[14] Tile_X4Y9_S_IO4/N4BEG[15] Tile_X4Y9_S_IO4/N4BEG[1] Tile_X4Y9_S_IO4/N4BEG[2]
+ Tile_X4Y9_S_IO4/N4BEG[3] Tile_X4Y9_S_IO4/N4BEG[4] Tile_X4Y9_S_IO4/N4BEG[5] Tile_X4Y9_S_IO4/N4BEG[6]
+ Tile_X4Y9_S_IO4/N4BEG[7] Tile_X4Y9_S_IO4/N4BEG[8] Tile_X4Y9_S_IO4/N4BEG[9] Tile_X4Y9_S_IO4/NN4BEG[0]
+ Tile_X4Y9_S_IO4/NN4BEG[10] Tile_X4Y9_S_IO4/NN4BEG[11] Tile_X4Y9_S_IO4/NN4BEG[12]
+ Tile_X4Y9_S_IO4/NN4BEG[13] Tile_X4Y9_S_IO4/NN4BEG[14] Tile_X4Y9_S_IO4/NN4BEG[15]
+ Tile_X4Y9_S_IO4/NN4BEG[1] Tile_X4Y9_S_IO4/NN4BEG[2] Tile_X4Y9_S_IO4/NN4BEG[3] Tile_X4Y9_S_IO4/NN4BEG[4]
+ Tile_X4Y9_S_IO4/NN4BEG[5] Tile_X4Y9_S_IO4/NN4BEG[6] Tile_X4Y9_S_IO4/NN4BEG[7] Tile_X4Y9_S_IO4/NN4BEG[8]
+ Tile_X4Y9_S_IO4/NN4BEG[9] Tile_X4Y9_S_IO4/S1END[0] Tile_X4Y9_S_IO4/S1END[1] Tile_X4Y9_S_IO4/S1END[2]
+ Tile_X4Y9_S_IO4/S1END[3] Tile_X4Y9_S_IO4/S2END[0] Tile_X4Y9_S_IO4/S2END[1] Tile_X4Y9_S_IO4/S2END[2]
+ Tile_X4Y9_S_IO4/S2END[3] Tile_X4Y9_S_IO4/S2END[4] Tile_X4Y9_S_IO4/S2END[5] Tile_X4Y9_S_IO4/S2END[6]
+ Tile_X4Y9_S_IO4/S2END[7] Tile_X4Y9_S_IO4/S2MID[0] Tile_X4Y9_S_IO4/S2MID[1] Tile_X4Y9_S_IO4/S2MID[2]
+ Tile_X4Y9_S_IO4/S2MID[3] Tile_X4Y9_S_IO4/S2MID[4] Tile_X4Y9_S_IO4/S2MID[5] Tile_X4Y9_S_IO4/S2MID[6]
+ Tile_X4Y9_S_IO4/S2MID[7] Tile_X4Y9_S_IO4/S4END[0] Tile_X4Y9_S_IO4/S4END[10] Tile_X4Y9_S_IO4/S4END[11]
+ Tile_X4Y9_S_IO4/S4END[12] Tile_X4Y9_S_IO4/S4END[13] Tile_X4Y9_S_IO4/S4END[14] Tile_X4Y9_S_IO4/S4END[15]
+ Tile_X4Y9_S_IO4/S4END[1] Tile_X4Y9_S_IO4/S4END[2] Tile_X4Y9_S_IO4/S4END[3] Tile_X4Y9_S_IO4/S4END[4]
+ Tile_X4Y9_S_IO4/S4END[5] Tile_X4Y9_S_IO4/S4END[6] Tile_X4Y9_S_IO4/S4END[7] Tile_X4Y9_S_IO4/S4END[8]
+ Tile_X4Y9_S_IO4/S4END[9] Tile_X4Y9_S_IO4/SS4END[0] Tile_X4Y9_S_IO4/SS4END[10] Tile_X4Y9_S_IO4/SS4END[11]
+ Tile_X4Y9_S_IO4/SS4END[12] Tile_X4Y9_S_IO4/SS4END[13] Tile_X4Y9_S_IO4/SS4END[14]
+ Tile_X4Y9_S_IO4/SS4END[15] Tile_X4Y9_S_IO4/SS4END[1] Tile_X4Y9_S_IO4/SS4END[2] Tile_X4Y9_S_IO4/SS4END[3]
+ Tile_X4Y9_S_IO4/SS4END[4] Tile_X4Y9_S_IO4/SS4END[5] Tile_X4Y9_S_IO4/SS4END[6] Tile_X4Y9_S_IO4/SS4END[7]
+ Tile_X4Y9_S_IO4/SS4END[8] Tile_X4Y9_S_IO4/SS4END[9] UserCLK Tile_X4Y9_S_IO4/UserCLKo
+ VGND VPWR S_IO4
XTile_X4Y4_LUT4AB Tile_X4Y5_LUT4AB/Co Tile_X4Y4_LUT4AB/Co Tile_X4Y4_LUT4AB/E1BEG[0]
+ Tile_X4Y4_LUT4AB/E1BEG[1] Tile_X4Y4_LUT4AB/E1BEG[2] Tile_X4Y4_LUT4AB/E1BEG[3] Tile_X4Y4_LUT4AB/E1END[0]
+ Tile_X4Y4_LUT4AB/E1END[1] Tile_X4Y4_LUT4AB/E1END[2] Tile_X4Y4_LUT4AB/E1END[3] Tile_X4Y4_LUT4AB/E2BEG[0]
+ Tile_X4Y4_LUT4AB/E2BEG[1] Tile_X4Y4_LUT4AB/E2BEG[2] Tile_X4Y4_LUT4AB/E2BEG[3] Tile_X4Y4_LUT4AB/E2BEG[4]
+ Tile_X4Y4_LUT4AB/E2BEG[5] Tile_X4Y4_LUT4AB/E2BEG[6] Tile_X4Y4_LUT4AB/E2BEG[7] Tile_X5Y4_E_TT_IF/E2END[0]
+ Tile_X5Y4_E_TT_IF/E2END[1] Tile_X5Y4_E_TT_IF/E2END[2] Tile_X5Y4_E_TT_IF/E2END[3]
+ Tile_X5Y4_E_TT_IF/E2END[4] Tile_X5Y4_E_TT_IF/E2END[5] Tile_X5Y4_E_TT_IF/E2END[6]
+ Tile_X5Y4_E_TT_IF/E2END[7] Tile_X4Y4_LUT4AB/E2END[0] Tile_X4Y4_LUT4AB/E2END[1] Tile_X4Y4_LUT4AB/E2END[2]
+ Tile_X4Y4_LUT4AB/E2END[3] Tile_X4Y4_LUT4AB/E2END[4] Tile_X4Y4_LUT4AB/E2END[5] Tile_X4Y4_LUT4AB/E2END[6]
+ Tile_X4Y4_LUT4AB/E2END[7] Tile_X4Y4_LUT4AB/E2MID[0] Tile_X4Y4_LUT4AB/E2MID[1] Tile_X4Y4_LUT4AB/E2MID[2]
+ Tile_X4Y4_LUT4AB/E2MID[3] Tile_X4Y4_LUT4AB/E2MID[4] Tile_X4Y4_LUT4AB/E2MID[5] Tile_X4Y4_LUT4AB/E2MID[6]
+ Tile_X4Y4_LUT4AB/E2MID[7] Tile_X4Y4_LUT4AB/E6BEG[0] Tile_X4Y4_LUT4AB/E6BEG[10] Tile_X4Y4_LUT4AB/E6BEG[11]
+ Tile_X4Y4_LUT4AB/E6BEG[1] Tile_X4Y4_LUT4AB/E6BEG[2] Tile_X4Y4_LUT4AB/E6BEG[3] Tile_X4Y4_LUT4AB/E6BEG[4]
+ Tile_X4Y4_LUT4AB/E6BEG[5] Tile_X4Y4_LUT4AB/E6BEG[6] Tile_X4Y4_LUT4AB/E6BEG[7] Tile_X4Y4_LUT4AB/E6BEG[8]
+ Tile_X4Y4_LUT4AB/E6BEG[9] Tile_X4Y4_LUT4AB/E6END[0] Tile_X4Y4_LUT4AB/E6END[10] Tile_X4Y4_LUT4AB/E6END[11]
+ Tile_X4Y4_LUT4AB/E6END[1] Tile_X4Y4_LUT4AB/E6END[2] Tile_X4Y4_LUT4AB/E6END[3] Tile_X4Y4_LUT4AB/E6END[4]
+ Tile_X4Y4_LUT4AB/E6END[5] Tile_X4Y4_LUT4AB/E6END[6] Tile_X4Y4_LUT4AB/E6END[7] Tile_X4Y4_LUT4AB/E6END[8]
+ Tile_X4Y4_LUT4AB/E6END[9] Tile_X4Y4_LUT4AB/EE4BEG[0] Tile_X4Y4_LUT4AB/EE4BEG[10]
+ Tile_X4Y4_LUT4AB/EE4BEG[11] Tile_X4Y4_LUT4AB/EE4BEG[12] Tile_X4Y4_LUT4AB/EE4BEG[13]
+ Tile_X4Y4_LUT4AB/EE4BEG[14] Tile_X4Y4_LUT4AB/EE4BEG[15] Tile_X4Y4_LUT4AB/EE4BEG[1]
+ Tile_X4Y4_LUT4AB/EE4BEG[2] Tile_X4Y4_LUT4AB/EE4BEG[3] Tile_X4Y4_LUT4AB/EE4BEG[4]
+ Tile_X4Y4_LUT4AB/EE4BEG[5] Tile_X4Y4_LUT4AB/EE4BEG[6] Tile_X4Y4_LUT4AB/EE4BEG[7]
+ Tile_X4Y4_LUT4AB/EE4BEG[8] Tile_X4Y4_LUT4AB/EE4BEG[9] Tile_X4Y4_LUT4AB/EE4END[0]
+ Tile_X4Y4_LUT4AB/EE4END[10] Tile_X4Y4_LUT4AB/EE4END[11] Tile_X4Y4_LUT4AB/EE4END[12]
+ Tile_X4Y4_LUT4AB/EE4END[13] Tile_X4Y4_LUT4AB/EE4END[14] Tile_X4Y4_LUT4AB/EE4END[15]
+ Tile_X4Y4_LUT4AB/EE4END[1] Tile_X4Y4_LUT4AB/EE4END[2] Tile_X4Y4_LUT4AB/EE4END[3]
+ Tile_X4Y4_LUT4AB/EE4END[4] Tile_X4Y4_LUT4AB/EE4END[5] Tile_X4Y4_LUT4AB/EE4END[6]
+ Tile_X4Y4_LUT4AB/EE4END[7] Tile_X4Y4_LUT4AB/EE4END[8] Tile_X4Y4_LUT4AB/EE4END[9]
+ Tile_X4Y4_LUT4AB/FrameData[0] Tile_X4Y4_LUT4AB/FrameData[10] Tile_X4Y4_LUT4AB/FrameData[11]
+ Tile_X4Y4_LUT4AB/FrameData[12] Tile_X4Y4_LUT4AB/FrameData[13] Tile_X4Y4_LUT4AB/FrameData[14]
+ Tile_X4Y4_LUT4AB/FrameData[15] Tile_X4Y4_LUT4AB/FrameData[16] Tile_X4Y4_LUT4AB/FrameData[17]
+ Tile_X4Y4_LUT4AB/FrameData[18] Tile_X4Y4_LUT4AB/FrameData[19] Tile_X4Y4_LUT4AB/FrameData[1]
+ Tile_X4Y4_LUT4AB/FrameData[20] Tile_X4Y4_LUT4AB/FrameData[21] Tile_X4Y4_LUT4AB/FrameData[22]
+ Tile_X4Y4_LUT4AB/FrameData[23] Tile_X4Y4_LUT4AB/FrameData[24] Tile_X4Y4_LUT4AB/FrameData[25]
+ Tile_X4Y4_LUT4AB/FrameData[26] Tile_X4Y4_LUT4AB/FrameData[27] Tile_X4Y4_LUT4AB/FrameData[28]
+ Tile_X4Y4_LUT4AB/FrameData[29] Tile_X4Y4_LUT4AB/FrameData[2] Tile_X4Y4_LUT4AB/FrameData[30]
+ Tile_X4Y4_LUT4AB/FrameData[31] Tile_X4Y4_LUT4AB/FrameData[3] Tile_X4Y4_LUT4AB/FrameData[4]
+ Tile_X4Y4_LUT4AB/FrameData[5] Tile_X4Y4_LUT4AB/FrameData[6] Tile_X4Y4_LUT4AB/FrameData[7]
+ Tile_X4Y4_LUT4AB/FrameData[8] Tile_X4Y4_LUT4AB/FrameData[9] Tile_X5Y4_E_TT_IF/FrameData[0]
+ Tile_X5Y4_E_TT_IF/FrameData[10] Tile_X5Y4_E_TT_IF/FrameData[11] Tile_X5Y4_E_TT_IF/FrameData[12]
+ Tile_X5Y4_E_TT_IF/FrameData[13] Tile_X5Y4_E_TT_IF/FrameData[14] Tile_X5Y4_E_TT_IF/FrameData[15]
+ Tile_X5Y4_E_TT_IF/FrameData[16] Tile_X5Y4_E_TT_IF/FrameData[17] Tile_X5Y4_E_TT_IF/FrameData[18]
+ Tile_X5Y4_E_TT_IF/FrameData[19] Tile_X5Y4_E_TT_IF/FrameData[1] Tile_X5Y4_E_TT_IF/FrameData[20]
+ Tile_X5Y4_E_TT_IF/FrameData[21] Tile_X5Y4_E_TT_IF/FrameData[22] Tile_X5Y4_E_TT_IF/FrameData[23]
+ Tile_X5Y4_E_TT_IF/FrameData[24] Tile_X5Y4_E_TT_IF/FrameData[25] Tile_X5Y4_E_TT_IF/FrameData[26]
+ Tile_X5Y4_E_TT_IF/FrameData[27] Tile_X5Y4_E_TT_IF/FrameData[28] Tile_X5Y4_E_TT_IF/FrameData[29]
+ Tile_X5Y4_E_TT_IF/FrameData[2] Tile_X5Y4_E_TT_IF/FrameData[30] Tile_X5Y4_E_TT_IF/FrameData[31]
+ Tile_X5Y4_E_TT_IF/FrameData[3] Tile_X5Y4_E_TT_IF/FrameData[4] Tile_X5Y4_E_TT_IF/FrameData[5]
+ Tile_X5Y4_E_TT_IF/FrameData[6] Tile_X5Y4_E_TT_IF/FrameData[7] Tile_X5Y4_E_TT_IF/FrameData[8]
+ Tile_X5Y4_E_TT_IF/FrameData[9] Tile_X4Y4_LUT4AB/FrameStrobe[0] Tile_X4Y4_LUT4AB/FrameStrobe[10]
+ Tile_X4Y4_LUT4AB/FrameStrobe[11] Tile_X4Y4_LUT4AB/FrameStrobe[12] Tile_X4Y4_LUT4AB/FrameStrobe[13]
+ Tile_X4Y4_LUT4AB/FrameStrobe[14] Tile_X4Y4_LUT4AB/FrameStrobe[15] Tile_X4Y4_LUT4AB/FrameStrobe[16]
+ Tile_X4Y4_LUT4AB/FrameStrobe[17] Tile_X4Y4_LUT4AB/FrameStrobe[18] Tile_X4Y4_LUT4AB/FrameStrobe[19]
+ Tile_X4Y4_LUT4AB/FrameStrobe[1] Tile_X4Y4_LUT4AB/FrameStrobe[2] Tile_X4Y4_LUT4AB/FrameStrobe[3]
+ Tile_X4Y4_LUT4AB/FrameStrobe[4] Tile_X4Y4_LUT4AB/FrameStrobe[5] Tile_X4Y4_LUT4AB/FrameStrobe[6]
+ Tile_X4Y4_LUT4AB/FrameStrobe[7] Tile_X4Y4_LUT4AB/FrameStrobe[8] Tile_X4Y4_LUT4AB/FrameStrobe[9]
+ Tile_X4Y3_LUT4AB/FrameStrobe[0] Tile_X4Y3_LUT4AB/FrameStrobe[10] Tile_X4Y3_LUT4AB/FrameStrobe[11]
+ Tile_X4Y3_LUT4AB/FrameStrobe[12] Tile_X4Y3_LUT4AB/FrameStrobe[13] Tile_X4Y3_LUT4AB/FrameStrobe[14]
+ Tile_X4Y3_LUT4AB/FrameStrobe[15] Tile_X4Y3_LUT4AB/FrameStrobe[16] Tile_X4Y3_LUT4AB/FrameStrobe[17]
+ Tile_X4Y3_LUT4AB/FrameStrobe[18] Tile_X4Y3_LUT4AB/FrameStrobe[19] Tile_X4Y3_LUT4AB/FrameStrobe[1]
+ Tile_X4Y3_LUT4AB/FrameStrobe[2] Tile_X4Y3_LUT4AB/FrameStrobe[3] Tile_X4Y3_LUT4AB/FrameStrobe[4]
+ Tile_X4Y3_LUT4AB/FrameStrobe[5] Tile_X4Y3_LUT4AB/FrameStrobe[6] Tile_X4Y3_LUT4AB/FrameStrobe[7]
+ Tile_X4Y3_LUT4AB/FrameStrobe[8] Tile_X4Y3_LUT4AB/FrameStrobe[9] Tile_X4Y4_LUT4AB/N1BEG[0]
+ Tile_X4Y4_LUT4AB/N1BEG[1] Tile_X4Y4_LUT4AB/N1BEG[2] Tile_X4Y4_LUT4AB/N1BEG[3] Tile_X4Y5_LUT4AB/N1BEG[0]
+ Tile_X4Y5_LUT4AB/N1BEG[1] Tile_X4Y5_LUT4AB/N1BEG[2] Tile_X4Y5_LUT4AB/N1BEG[3] Tile_X4Y4_LUT4AB/N2BEG[0]
+ Tile_X4Y4_LUT4AB/N2BEG[1] Tile_X4Y4_LUT4AB/N2BEG[2] Tile_X4Y4_LUT4AB/N2BEG[3] Tile_X4Y4_LUT4AB/N2BEG[4]
+ Tile_X4Y4_LUT4AB/N2BEG[5] Tile_X4Y4_LUT4AB/N2BEG[6] Tile_X4Y4_LUT4AB/N2BEG[7] Tile_X4Y3_LUT4AB/N2END[0]
+ Tile_X4Y3_LUT4AB/N2END[1] Tile_X4Y3_LUT4AB/N2END[2] Tile_X4Y3_LUT4AB/N2END[3] Tile_X4Y3_LUT4AB/N2END[4]
+ Tile_X4Y3_LUT4AB/N2END[5] Tile_X4Y3_LUT4AB/N2END[6] Tile_X4Y3_LUT4AB/N2END[7] Tile_X4Y4_LUT4AB/N2END[0]
+ Tile_X4Y4_LUT4AB/N2END[1] Tile_X4Y4_LUT4AB/N2END[2] Tile_X4Y4_LUT4AB/N2END[3] Tile_X4Y4_LUT4AB/N2END[4]
+ Tile_X4Y4_LUT4AB/N2END[5] Tile_X4Y4_LUT4AB/N2END[6] Tile_X4Y4_LUT4AB/N2END[7] Tile_X4Y5_LUT4AB/N2BEG[0]
+ Tile_X4Y5_LUT4AB/N2BEG[1] Tile_X4Y5_LUT4AB/N2BEG[2] Tile_X4Y5_LUT4AB/N2BEG[3] Tile_X4Y5_LUT4AB/N2BEG[4]
+ Tile_X4Y5_LUT4AB/N2BEG[5] Tile_X4Y5_LUT4AB/N2BEG[6] Tile_X4Y5_LUT4AB/N2BEG[7] Tile_X4Y4_LUT4AB/N4BEG[0]
+ Tile_X4Y4_LUT4AB/N4BEG[10] Tile_X4Y4_LUT4AB/N4BEG[11] Tile_X4Y4_LUT4AB/N4BEG[12]
+ Tile_X4Y4_LUT4AB/N4BEG[13] Tile_X4Y4_LUT4AB/N4BEG[14] Tile_X4Y4_LUT4AB/N4BEG[15]
+ Tile_X4Y4_LUT4AB/N4BEG[1] Tile_X4Y4_LUT4AB/N4BEG[2] Tile_X4Y4_LUT4AB/N4BEG[3] Tile_X4Y4_LUT4AB/N4BEG[4]
+ Tile_X4Y4_LUT4AB/N4BEG[5] Tile_X4Y4_LUT4AB/N4BEG[6] Tile_X4Y4_LUT4AB/N4BEG[7] Tile_X4Y4_LUT4AB/N4BEG[8]
+ Tile_X4Y4_LUT4AB/N4BEG[9] Tile_X4Y5_LUT4AB/N4BEG[0] Tile_X4Y5_LUT4AB/N4BEG[10] Tile_X4Y5_LUT4AB/N4BEG[11]
+ Tile_X4Y5_LUT4AB/N4BEG[12] Tile_X4Y5_LUT4AB/N4BEG[13] Tile_X4Y5_LUT4AB/N4BEG[14]
+ Tile_X4Y5_LUT4AB/N4BEG[15] Tile_X4Y5_LUT4AB/N4BEG[1] Tile_X4Y5_LUT4AB/N4BEG[2] Tile_X4Y5_LUT4AB/N4BEG[3]
+ Tile_X4Y5_LUT4AB/N4BEG[4] Tile_X4Y5_LUT4AB/N4BEG[5] Tile_X4Y5_LUT4AB/N4BEG[6] Tile_X4Y5_LUT4AB/N4BEG[7]
+ Tile_X4Y5_LUT4AB/N4BEG[8] Tile_X4Y5_LUT4AB/N4BEG[9] Tile_X4Y4_LUT4AB/NN4BEG[0] Tile_X4Y4_LUT4AB/NN4BEG[10]
+ Tile_X4Y4_LUT4AB/NN4BEG[11] Tile_X4Y4_LUT4AB/NN4BEG[12] Tile_X4Y4_LUT4AB/NN4BEG[13]
+ Tile_X4Y4_LUT4AB/NN4BEG[14] Tile_X4Y4_LUT4AB/NN4BEG[15] Tile_X4Y4_LUT4AB/NN4BEG[1]
+ Tile_X4Y4_LUT4AB/NN4BEG[2] Tile_X4Y4_LUT4AB/NN4BEG[3] Tile_X4Y4_LUT4AB/NN4BEG[4]
+ Tile_X4Y4_LUT4AB/NN4BEG[5] Tile_X4Y4_LUT4AB/NN4BEG[6] Tile_X4Y4_LUT4AB/NN4BEG[7]
+ Tile_X4Y4_LUT4AB/NN4BEG[8] Tile_X4Y4_LUT4AB/NN4BEG[9] Tile_X4Y5_LUT4AB/NN4BEG[0]
+ Tile_X4Y5_LUT4AB/NN4BEG[10] Tile_X4Y5_LUT4AB/NN4BEG[11] Tile_X4Y5_LUT4AB/NN4BEG[12]
+ Tile_X4Y5_LUT4AB/NN4BEG[13] Tile_X4Y5_LUT4AB/NN4BEG[14] Tile_X4Y5_LUT4AB/NN4BEG[15]
+ Tile_X4Y5_LUT4AB/NN4BEG[1] Tile_X4Y5_LUT4AB/NN4BEG[2] Tile_X4Y5_LUT4AB/NN4BEG[3]
+ Tile_X4Y5_LUT4AB/NN4BEG[4] Tile_X4Y5_LUT4AB/NN4BEG[5] Tile_X4Y5_LUT4AB/NN4BEG[6]
+ Tile_X4Y5_LUT4AB/NN4BEG[7] Tile_X4Y5_LUT4AB/NN4BEG[8] Tile_X4Y5_LUT4AB/NN4BEG[9]
+ Tile_X4Y5_LUT4AB/S1END[0] Tile_X4Y5_LUT4AB/S1END[1] Tile_X4Y5_LUT4AB/S1END[2] Tile_X4Y5_LUT4AB/S1END[3]
+ Tile_X4Y4_LUT4AB/S1END[0] Tile_X4Y4_LUT4AB/S1END[1] Tile_X4Y4_LUT4AB/S1END[2] Tile_X4Y4_LUT4AB/S1END[3]
+ Tile_X4Y5_LUT4AB/S2MID[0] Tile_X4Y5_LUT4AB/S2MID[1] Tile_X4Y5_LUT4AB/S2MID[2] Tile_X4Y5_LUT4AB/S2MID[3]
+ Tile_X4Y5_LUT4AB/S2MID[4] Tile_X4Y5_LUT4AB/S2MID[5] Tile_X4Y5_LUT4AB/S2MID[6] Tile_X4Y5_LUT4AB/S2MID[7]
+ Tile_X4Y5_LUT4AB/S2END[0] Tile_X4Y5_LUT4AB/S2END[1] Tile_X4Y5_LUT4AB/S2END[2] Tile_X4Y5_LUT4AB/S2END[3]
+ Tile_X4Y5_LUT4AB/S2END[4] Tile_X4Y5_LUT4AB/S2END[5] Tile_X4Y5_LUT4AB/S2END[6] Tile_X4Y5_LUT4AB/S2END[7]
+ Tile_X4Y4_LUT4AB/S2END[0] Tile_X4Y4_LUT4AB/S2END[1] Tile_X4Y4_LUT4AB/S2END[2] Tile_X4Y4_LUT4AB/S2END[3]
+ Tile_X4Y4_LUT4AB/S2END[4] Tile_X4Y4_LUT4AB/S2END[5] Tile_X4Y4_LUT4AB/S2END[6] Tile_X4Y4_LUT4AB/S2END[7]
+ Tile_X4Y4_LUT4AB/S2MID[0] Tile_X4Y4_LUT4AB/S2MID[1] Tile_X4Y4_LUT4AB/S2MID[2] Tile_X4Y4_LUT4AB/S2MID[3]
+ Tile_X4Y4_LUT4AB/S2MID[4] Tile_X4Y4_LUT4AB/S2MID[5] Tile_X4Y4_LUT4AB/S2MID[6] Tile_X4Y4_LUT4AB/S2MID[7]
+ Tile_X4Y5_LUT4AB/S4END[0] Tile_X4Y5_LUT4AB/S4END[10] Tile_X4Y5_LUT4AB/S4END[11]
+ Tile_X4Y5_LUT4AB/S4END[12] Tile_X4Y5_LUT4AB/S4END[13] Tile_X4Y5_LUT4AB/S4END[14]
+ Tile_X4Y5_LUT4AB/S4END[15] Tile_X4Y5_LUT4AB/S4END[1] Tile_X4Y5_LUT4AB/S4END[2] Tile_X4Y5_LUT4AB/S4END[3]
+ Tile_X4Y5_LUT4AB/S4END[4] Tile_X4Y5_LUT4AB/S4END[5] Tile_X4Y5_LUT4AB/S4END[6] Tile_X4Y5_LUT4AB/S4END[7]
+ Tile_X4Y5_LUT4AB/S4END[8] Tile_X4Y5_LUT4AB/S4END[9] Tile_X4Y4_LUT4AB/S4END[0] Tile_X4Y4_LUT4AB/S4END[10]
+ Tile_X4Y4_LUT4AB/S4END[11] Tile_X4Y4_LUT4AB/S4END[12] Tile_X4Y4_LUT4AB/S4END[13]
+ Tile_X4Y4_LUT4AB/S4END[14] Tile_X4Y4_LUT4AB/S4END[15] Tile_X4Y4_LUT4AB/S4END[1]
+ Tile_X4Y4_LUT4AB/S4END[2] Tile_X4Y4_LUT4AB/S4END[3] Tile_X4Y4_LUT4AB/S4END[4] Tile_X4Y4_LUT4AB/S4END[5]
+ Tile_X4Y4_LUT4AB/S4END[6] Tile_X4Y4_LUT4AB/S4END[7] Tile_X4Y4_LUT4AB/S4END[8] Tile_X4Y4_LUT4AB/S4END[9]
+ Tile_X4Y5_LUT4AB/SS4END[0] Tile_X4Y5_LUT4AB/SS4END[10] Tile_X4Y5_LUT4AB/SS4END[11]
+ Tile_X4Y5_LUT4AB/SS4END[12] Tile_X4Y5_LUT4AB/SS4END[13] Tile_X4Y5_LUT4AB/SS4END[14]
+ Tile_X4Y5_LUT4AB/SS4END[15] Tile_X4Y5_LUT4AB/SS4END[1] Tile_X4Y5_LUT4AB/SS4END[2]
+ Tile_X4Y5_LUT4AB/SS4END[3] Tile_X4Y5_LUT4AB/SS4END[4] Tile_X4Y5_LUT4AB/SS4END[5]
+ Tile_X4Y5_LUT4AB/SS4END[6] Tile_X4Y5_LUT4AB/SS4END[7] Tile_X4Y5_LUT4AB/SS4END[8]
+ Tile_X4Y5_LUT4AB/SS4END[9] Tile_X4Y4_LUT4AB/SS4END[0] Tile_X4Y4_LUT4AB/SS4END[10]
+ Tile_X4Y4_LUT4AB/SS4END[11] Tile_X4Y4_LUT4AB/SS4END[12] Tile_X4Y4_LUT4AB/SS4END[13]
+ Tile_X4Y4_LUT4AB/SS4END[14] Tile_X4Y4_LUT4AB/SS4END[15] Tile_X4Y4_LUT4AB/SS4END[1]
+ Tile_X4Y4_LUT4AB/SS4END[2] Tile_X4Y4_LUT4AB/SS4END[3] Tile_X4Y4_LUT4AB/SS4END[4]
+ Tile_X4Y4_LUT4AB/SS4END[5] Tile_X4Y4_LUT4AB/SS4END[6] Tile_X4Y4_LUT4AB/SS4END[7]
+ Tile_X4Y4_LUT4AB/SS4END[8] Tile_X4Y4_LUT4AB/SS4END[9] Tile_X4Y4_LUT4AB/UserCLK Tile_X4Y3_LUT4AB/UserCLK
+ VGND VPWR Tile_X4Y4_LUT4AB/W1BEG[0] Tile_X4Y4_LUT4AB/W1BEG[1] Tile_X4Y4_LUT4AB/W1BEG[2]
+ Tile_X4Y4_LUT4AB/W1BEG[3] Tile_X4Y4_LUT4AB/W1END[0] Tile_X4Y4_LUT4AB/W1END[1] Tile_X4Y4_LUT4AB/W1END[2]
+ Tile_X4Y4_LUT4AB/W1END[3] Tile_X4Y4_LUT4AB/W2BEG[0] Tile_X4Y4_LUT4AB/W2BEG[1] Tile_X4Y4_LUT4AB/W2BEG[2]
+ Tile_X4Y4_LUT4AB/W2BEG[3] Tile_X4Y4_LUT4AB/W2BEG[4] Tile_X4Y4_LUT4AB/W2BEG[5] Tile_X4Y4_LUT4AB/W2BEG[6]
+ Tile_X4Y4_LUT4AB/W2BEG[7] Tile_X3Y4_LUT4AB/W2END[0] Tile_X3Y4_LUT4AB/W2END[1] Tile_X3Y4_LUT4AB/W2END[2]
+ Tile_X3Y4_LUT4AB/W2END[3] Tile_X3Y4_LUT4AB/W2END[4] Tile_X3Y4_LUT4AB/W2END[5] Tile_X3Y4_LUT4AB/W2END[6]
+ Tile_X3Y4_LUT4AB/W2END[7] Tile_X4Y4_LUT4AB/W2END[0] Tile_X4Y4_LUT4AB/W2END[1] Tile_X4Y4_LUT4AB/W2END[2]
+ Tile_X4Y4_LUT4AB/W2END[3] Tile_X4Y4_LUT4AB/W2END[4] Tile_X4Y4_LUT4AB/W2END[5] Tile_X4Y4_LUT4AB/W2END[6]
+ Tile_X4Y4_LUT4AB/W2END[7] Tile_X4Y4_LUT4AB/W2MID[0] Tile_X4Y4_LUT4AB/W2MID[1] Tile_X4Y4_LUT4AB/W2MID[2]
+ Tile_X4Y4_LUT4AB/W2MID[3] Tile_X4Y4_LUT4AB/W2MID[4] Tile_X4Y4_LUT4AB/W2MID[5] Tile_X4Y4_LUT4AB/W2MID[6]
+ Tile_X4Y4_LUT4AB/W2MID[7] Tile_X4Y4_LUT4AB/W6BEG[0] Tile_X4Y4_LUT4AB/W6BEG[10] Tile_X4Y4_LUT4AB/W6BEG[11]
+ Tile_X4Y4_LUT4AB/W6BEG[1] Tile_X4Y4_LUT4AB/W6BEG[2] Tile_X4Y4_LUT4AB/W6BEG[3] Tile_X4Y4_LUT4AB/W6BEG[4]
+ Tile_X4Y4_LUT4AB/W6BEG[5] Tile_X4Y4_LUT4AB/W6BEG[6] Tile_X4Y4_LUT4AB/W6BEG[7] Tile_X4Y4_LUT4AB/W6BEG[8]
+ Tile_X4Y4_LUT4AB/W6BEG[9] Tile_X4Y4_LUT4AB/W6END[0] Tile_X4Y4_LUT4AB/W6END[10] Tile_X4Y4_LUT4AB/W6END[11]
+ Tile_X4Y4_LUT4AB/W6END[1] Tile_X4Y4_LUT4AB/W6END[2] Tile_X4Y4_LUT4AB/W6END[3] Tile_X4Y4_LUT4AB/W6END[4]
+ Tile_X4Y4_LUT4AB/W6END[5] Tile_X4Y4_LUT4AB/W6END[6] Tile_X4Y4_LUT4AB/W6END[7] Tile_X4Y4_LUT4AB/W6END[8]
+ Tile_X4Y4_LUT4AB/W6END[9] Tile_X4Y4_LUT4AB/WW4BEG[0] Tile_X4Y4_LUT4AB/WW4BEG[10]
+ Tile_X4Y4_LUT4AB/WW4BEG[11] Tile_X4Y4_LUT4AB/WW4BEG[12] Tile_X4Y4_LUT4AB/WW4BEG[13]
+ Tile_X4Y4_LUT4AB/WW4BEG[14] Tile_X4Y4_LUT4AB/WW4BEG[15] Tile_X4Y4_LUT4AB/WW4BEG[1]
+ Tile_X4Y4_LUT4AB/WW4BEG[2] Tile_X4Y4_LUT4AB/WW4BEG[3] Tile_X4Y4_LUT4AB/WW4BEG[4]
+ Tile_X4Y4_LUT4AB/WW4BEG[5] Tile_X4Y4_LUT4AB/WW4BEG[6] Tile_X4Y4_LUT4AB/WW4BEG[7]
+ Tile_X4Y4_LUT4AB/WW4BEG[8] Tile_X4Y4_LUT4AB/WW4BEG[9] Tile_X4Y4_LUT4AB/WW4END[0]
+ Tile_X4Y4_LUT4AB/WW4END[10] Tile_X4Y4_LUT4AB/WW4END[11] Tile_X4Y4_LUT4AB/WW4END[12]
+ Tile_X4Y4_LUT4AB/WW4END[13] Tile_X4Y4_LUT4AB/WW4END[14] Tile_X4Y4_LUT4AB/WW4END[15]
+ Tile_X4Y4_LUT4AB/WW4END[1] Tile_X4Y4_LUT4AB/WW4END[2] Tile_X4Y4_LUT4AB/WW4END[3]
+ Tile_X4Y4_LUT4AB/WW4END[4] Tile_X4Y4_LUT4AB/WW4END[5] Tile_X4Y4_LUT4AB/WW4END[6]
+ Tile_X4Y4_LUT4AB/WW4END[7] Tile_X4Y4_LUT4AB/WW4END[8] Tile_X4Y4_LUT4AB/WW4END[9]
+ LUT4AB
XTile_X3Y8_LUT4AB Tile_X3Y9_S_IO4/Co Tile_X3Y8_LUT4AB/Co Tile_X4Y8_LUT4AB/E1END[0]
+ Tile_X4Y8_LUT4AB/E1END[1] Tile_X4Y8_LUT4AB/E1END[2] Tile_X4Y8_LUT4AB/E1END[3] Tile_X3Y8_LUT4AB/E1END[0]
+ Tile_X3Y8_LUT4AB/E1END[1] Tile_X3Y8_LUT4AB/E1END[2] Tile_X3Y8_LUT4AB/E1END[3] Tile_X4Y8_LUT4AB/E2MID[0]
+ Tile_X4Y8_LUT4AB/E2MID[1] Tile_X4Y8_LUT4AB/E2MID[2] Tile_X4Y8_LUT4AB/E2MID[3] Tile_X4Y8_LUT4AB/E2MID[4]
+ Tile_X4Y8_LUT4AB/E2MID[5] Tile_X4Y8_LUT4AB/E2MID[6] Tile_X4Y8_LUT4AB/E2MID[7] Tile_X4Y8_LUT4AB/E2END[0]
+ Tile_X4Y8_LUT4AB/E2END[1] Tile_X4Y8_LUT4AB/E2END[2] Tile_X4Y8_LUT4AB/E2END[3] Tile_X4Y8_LUT4AB/E2END[4]
+ Tile_X4Y8_LUT4AB/E2END[5] Tile_X4Y8_LUT4AB/E2END[6] Tile_X4Y8_LUT4AB/E2END[7] Tile_X3Y8_LUT4AB/E2END[0]
+ Tile_X3Y8_LUT4AB/E2END[1] Tile_X3Y8_LUT4AB/E2END[2] Tile_X3Y8_LUT4AB/E2END[3] Tile_X3Y8_LUT4AB/E2END[4]
+ Tile_X3Y8_LUT4AB/E2END[5] Tile_X3Y8_LUT4AB/E2END[6] Tile_X3Y8_LUT4AB/E2END[7] Tile_X3Y8_LUT4AB/E2MID[0]
+ Tile_X3Y8_LUT4AB/E2MID[1] Tile_X3Y8_LUT4AB/E2MID[2] Tile_X3Y8_LUT4AB/E2MID[3] Tile_X3Y8_LUT4AB/E2MID[4]
+ Tile_X3Y8_LUT4AB/E2MID[5] Tile_X3Y8_LUT4AB/E2MID[6] Tile_X3Y8_LUT4AB/E2MID[7] Tile_X4Y8_LUT4AB/E6END[0]
+ Tile_X4Y8_LUT4AB/E6END[10] Tile_X4Y8_LUT4AB/E6END[11] Tile_X4Y8_LUT4AB/E6END[1]
+ Tile_X4Y8_LUT4AB/E6END[2] Tile_X4Y8_LUT4AB/E6END[3] Tile_X4Y8_LUT4AB/E6END[4] Tile_X4Y8_LUT4AB/E6END[5]
+ Tile_X4Y8_LUT4AB/E6END[6] Tile_X4Y8_LUT4AB/E6END[7] Tile_X4Y8_LUT4AB/E6END[8] Tile_X4Y8_LUT4AB/E6END[9]
+ Tile_X3Y8_LUT4AB/E6END[0] Tile_X3Y8_LUT4AB/E6END[10] Tile_X3Y8_LUT4AB/E6END[11]
+ Tile_X3Y8_LUT4AB/E6END[1] Tile_X3Y8_LUT4AB/E6END[2] Tile_X3Y8_LUT4AB/E6END[3] Tile_X3Y8_LUT4AB/E6END[4]
+ Tile_X3Y8_LUT4AB/E6END[5] Tile_X3Y8_LUT4AB/E6END[6] Tile_X3Y8_LUT4AB/E6END[7] Tile_X3Y8_LUT4AB/E6END[8]
+ Tile_X3Y8_LUT4AB/E6END[9] Tile_X4Y8_LUT4AB/EE4END[0] Tile_X4Y8_LUT4AB/EE4END[10]
+ Tile_X4Y8_LUT4AB/EE4END[11] Tile_X4Y8_LUT4AB/EE4END[12] Tile_X4Y8_LUT4AB/EE4END[13]
+ Tile_X4Y8_LUT4AB/EE4END[14] Tile_X4Y8_LUT4AB/EE4END[15] Tile_X4Y8_LUT4AB/EE4END[1]
+ Tile_X4Y8_LUT4AB/EE4END[2] Tile_X4Y8_LUT4AB/EE4END[3] Tile_X4Y8_LUT4AB/EE4END[4]
+ Tile_X4Y8_LUT4AB/EE4END[5] Tile_X4Y8_LUT4AB/EE4END[6] Tile_X4Y8_LUT4AB/EE4END[7]
+ Tile_X4Y8_LUT4AB/EE4END[8] Tile_X4Y8_LUT4AB/EE4END[9] Tile_X3Y8_LUT4AB/EE4END[0]
+ Tile_X3Y8_LUT4AB/EE4END[10] Tile_X3Y8_LUT4AB/EE4END[11] Tile_X3Y8_LUT4AB/EE4END[12]
+ Tile_X3Y8_LUT4AB/EE4END[13] Tile_X3Y8_LUT4AB/EE4END[14] Tile_X3Y8_LUT4AB/EE4END[15]
+ Tile_X3Y8_LUT4AB/EE4END[1] Tile_X3Y8_LUT4AB/EE4END[2] Tile_X3Y8_LUT4AB/EE4END[3]
+ Tile_X3Y8_LUT4AB/EE4END[4] Tile_X3Y8_LUT4AB/EE4END[5] Tile_X3Y8_LUT4AB/EE4END[6]
+ Tile_X3Y8_LUT4AB/EE4END[7] Tile_X3Y8_LUT4AB/EE4END[8] Tile_X3Y8_LUT4AB/EE4END[9]
+ Tile_X3Y8_LUT4AB/FrameData[0] Tile_X3Y8_LUT4AB/FrameData[10] Tile_X3Y8_LUT4AB/FrameData[11]
+ Tile_X3Y8_LUT4AB/FrameData[12] Tile_X3Y8_LUT4AB/FrameData[13] Tile_X3Y8_LUT4AB/FrameData[14]
+ Tile_X3Y8_LUT4AB/FrameData[15] Tile_X3Y8_LUT4AB/FrameData[16] Tile_X3Y8_LUT4AB/FrameData[17]
+ Tile_X3Y8_LUT4AB/FrameData[18] Tile_X3Y8_LUT4AB/FrameData[19] Tile_X3Y8_LUT4AB/FrameData[1]
+ Tile_X3Y8_LUT4AB/FrameData[20] Tile_X3Y8_LUT4AB/FrameData[21] Tile_X3Y8_LUT4AB/FrameData[22]
+ Tile_X3Y8_LUT4AB/FrameData[23] Tile_X3Y8_LUT4AB/FrameData[24] Tile_X3Y8_LUT4AB/FrameData[25]
+ Tile_X3Y8_LUT4AB/FrameData[26] Tile_X3Y8_LUT4AB/FrameData[27] Tile_X3Y8_LUT4AB/FrameData[28]
+ Tile_X3Y8_LUT4AB/FrameData[29] Tile_X3Y8_LUT4AB/FrameData[2] Tile_X3Y8_LUT4AB/FrameData[30]
+ Tile_X3Y8_LUT4AB/FrameData[31] Tile_X3Y8_LUT4AB/FrameData[3] Tile_X3Y8_LUT4AB/FrameData[4]
+ Tile_X3Y8_LUT4AB/FrameData[5] Tile_X3Y8_LUT4AB/FrameData[6] Tile_X3Y8_LUT4AB/FrameData[7]
+ Tile_X3Y8_LUT4AB/FrameData[8] Tile_X3Y8_LUT4AB/FrameData[9] Tile_X4Y8_LUT4AB/FrameData[0]
+ Tile_X4Y8_LUT4AB/FrameData[10] Tile_X4Y8_LUT4AB/FrameData[11] Tile_X4Y8_LUT4AB/FrameData[12]
+ Tile_X4Y8_LUT4AB/FrameData[13] Tile_X4Y8_LUT4AB/FrameData[14] Tile_X4Y8_LUT4AB/FrameData[15]
+ Tile_X4Y8_LUT4AB/FrameData[16] Tile_X4Y8_LUT4AB/FrameData[17] Tile_X4Y8_LUT4AB/FrameData[18]
+ Tile_X4Y8_LUT4AB/FrameData[19] Tile_X4Y8_LUT4AB/FrameData[1] Tile_X4Y8_LUT4AB/FrameData[20]
+ Tile_X4Y8_LUT4AB/FrameData[21] Tile_X4Y8_LUT4AB/FrameData[22] Tile_X4Y8_LUT4AB/FrameData[23]
+ Tile_X4Y8_LUT4AB/FrameData[24] Tile_X4Y8_LUT4AB/FrameData[25] Tile_X4Y8_LUT4AB/FrameData[26]
+ Tile_X4Y8_LUT4AB/FrameData[27] Tile_X4Y8_LUT4AB/FrameData[28] Tile_X4Y8_LUT4AB/FrameData[29]
+ Tile_X4Y8_LUT4AB/FrameData[2] Tile_X4Y8_LUT4AB/FrameData[30] Tile_X4Y8_LUT4AB/FrameData[31]
+ Tile_X4Y8_LUT4AB/FrameData[3] Tile_X4Y8_LUT4AB/FrameData[4] Tile_X4Y8_LUT4AB/FrameData[5]
+ Tile_X4Y8_LUT4AB/FrameData[6] Tile_X4Y8_LUT4AB/FrameData[7] Tile_X4Y8_LUT4AB/FrameData[8]
+ Tile_X4Y8_LUT4AB/FrameData[9] Tile_X3Y8_LUT4AB/FrameStrobe[0] Tile_X3Y8_LUT4AB/FrameStrobe[10]
+ Tile_X3Y8_LUT4AB/FrameStrobe[11] Tile_X3Y8_LUT4AB/FrameStrobe[12] Tile_X3Y8_LUT4AB/FrameStrobe[13]
+ Tile_X3Y8_LUT4AB/FrameStrobe[14] Tile_X3Y8_LUT4AB/FrameStrobe[15] Tile_X3Y8_LUT4AB/FrameStrobe[16]
+ Tile_X3Y8_LUT4AB/FrameStrobe[17] Tile_X3Y8_LUT4AB/FrameStrobe[18] Tile_X3Y8_LUT4AB/FrameStrobe[19]
+ Tile_X3Y8_LUT4AB/FrameStrobe[1] Tile_X3Y8_LUT4AB/FrameStrobe[2] Tile_X3Y8_LUT4AB/FrameStrobe[3]
+ Tile_X3Y8_LUT4AB/FrameStrobe[4] Tile_X3Y8_LUT4AB/FrameStrobe[5] Tile_X3Y8_LUT4AB/FrameStrobe[6]
+ Tile_X3Y8_LUT4AB/FrameStrobe[7] Tile_X3Y8_LUT4AB/FrameStrobe[8] Tile_X3Y8_LUT4AB/FrameStrobe[9]
+ Tile_X3Y7_LUT4AB/FrameStrobe[0] Tile_X3Y7_LUT4AB/FrameStrobe[10] Tile_X3Y7_LUT4AB/FrameStrobe[11]
+ Tile_X3Y7_LUT4AB/FrameStrobe[12] Tile_X3Y7_LUT4AB/FrameStrobe[13] Tile_X3Y7_LUT4AB/FrameStrobe[14]
+ Tile_X3Y7_LUT4AB/FrameStrobe[15] Tile_X3Y7_LUT4AB/FrameStrobe[16] Tile_X3Y7_LUT4AB/FrameStrobe[17]
+ Tile_X3Y7_LUT4AB/FrameStrobe[18] Tile_X3Y7_LUT4AB/FrameStrobe[19] Tile_X3Y7_LUT4AB/FrameStrobe[1]
+ Tile_X3Y7_LUT4AB/FrameStrobe[2] Tile_X3Y7_LUT4AB/FrameStrobe[3] Tile_X3Y7_LUT4AB/FrameStrobe[4]
+ Tile_X3Y7_LUT4AB/FrameStrobe[5] Tile_X3Y7_LUT4AB/FrameStrobe[6] Tile_X3Y7_LUT4AB/FrameStrobe[7]
+ Tile_X3Y7_LUT4AB/FrameStrobe[8] Tile_X3Y7_LUT4AB/FrameStrobe[9] Tile_X3Y8_LUT4AB/N1BEG[0]
+ Tile_X3Y8_LUT4AB/N1BEG[1] Tile_X3Y8_LUT4AB/N1BEG[2] Tile_X3Y8_LUT4AB/N1BEG[3] Tile_X3Y9_S_IO4/N1BEG[0]
+ Tile_X3Y9_S_IO4/N1BEG[1] Tile_X3Y9_S_IO4/N1BEG[2] Tile_X3Y9_S_IO4/N1BEG[3] Tile_X3Y8_LUT4AB/N2BEG[0]
+ Tile_X3Y8_LUT4AB/N2BEG[1] Tile_X3Y8_LUT4AB/N2BEG[2] Tile_X3Y8_LUT4AB/N2BEG[3] Tile_X3Y8_LUT4AB/N2BEG[4]
+ Tile_X3Y8_LUT4AB/N2BEG[5] Tile_X3Y8_LUT4AB/N2BEG[6] Tile_X3Y8_LUT4AB/N2BEG[7] Tile_X3Y7_LUT4AB/N2END[0]
+ Tile_X3Y7_LUT4AB/N2END[1] Tile_X3Y7_LUT4AB/N2END[2] Tile_X3Y7_LUT4AB/N2END[3] Tile_X3Y7_LUT4AB/N2END[4]
+ Tile_X3Y7_LUT4AB/N2END[5] Tile_X3Y7_LUT4AB/N2END[6] Tile_X3Y7_LUT4AB/N2END[7] Tile_X3Y9_S_IO4/N2BEGb[0]
+ Tile_X3Y9_S_IO4/N2BEGb[1] Tile_X3Y9_S_IO4/N2BEGb[2] Tile_X3Y9_S_IO4/N2BEGb[3] Tile_X3Y9_S_IO4/N2BEGb[4]
+ Tile_X3Y9_S_IO4/N2BEGb[5] Tile_X3Y9_S_IO4/N2BEGb[6] Tile_X3Y9_S_IO4/N2BEGb[7] Tile_X3Y9_S_IO4/N2BEG[0]
+ Tile_X3Y9_S_IO4/N2BEG[1] Tile_X3Y9_S_IO4/N2BEG[2] Tile_X3Y9_S_IO4/N2BEG[3] Tile_X3Y9_S_IO4/N2BEG[4]
+ Tile_X3Y9_S_IO4/N2BEG[5] Tile_X3Y9_S_IO4/N2BEG[6] Tile_X3Y9_S_IO4/N2BEG[7] Tile_X3Y8_LUT4AB/N4BEG[0]
+ Tile_X3Y8_LUT4AB/N4BEG[10] Tile_X3Y8_LUT4AB/N4BEG[11] Tile_X3Y8_LUT4AB/N4BEG[12]
+ Tile_X3Y8_LUT4AB/N4BEG[13] Tile_X3Y8_LUT4AB/N4BEG[14] Tile_X3Y8_LUT4AB/N4BEG[15]
+ Tile_X3Y8_LUT4AB/N4BEG[1] Tile_X3Y8_LUT4AB/N4BEG[2] Tile_X3Y8_LUT4AB/N4BEG[3] Tile_X3Y8_LUT4AB/N4BEG[4]
+ Tile_X3Y8_LUT4AB/N4BEG[5] Tile_X3Y8_LUT4AB/N4BEG[6] Tile_X3Y8_LUT4AB/N4BEG[7] Tile_X3Y8_LUT4AB/N4BEG[8]
+ Tile_X3Y8_LUT4AB/N4BEG[9] Tile_X3Y9_S_IO4/N4BEG[0] Tile_X3Y9_S_IO4/N4BEG[10] Tile_X3Y9_S_IO4/N4BEG[11]
+ Tile_X3Y9_S_IO4/N4BEG[12] Tile_X3Y9_S_IO4/N4BEG[13] Tile_X3Y9_S_IO4/N4BEG[14] Tile_X3Y9_S_IO4/N4BEG[15]
+ Tile_X3Y9_S_IO4/N4BEG[1] Tile_X3Y9_S_IO4/N4BEG[2] Tile_X3Y9_S_IO4/N4BEG[3] Tile_X3Y9_S_IO4/N4BEG[4]
+ Tile_X3Y9_S_IO4/N4BEG[5] Tile_X3Y9_S_IO4/N4BEG[6] Tile_X3Y9_S_IO4/N4BEG[7] Tile_X3Y9_S_IO4/N4BEG[8]
+ Tile_X3Y9_S_IO4/N4BEG[9] Tile_X3Y8_LUT4AB/NN4BEG[0] Tile_X3Y8_LUT4AB/NN4BEG[10]
+ Tile_X3Y8_LUT4AB/NN4BEG[11] Tile_X3Y8_LUT4AB/NN4BEG[12] Tile_X3Y8_LUT4AB/NN4BEG[13]
+ Tile_X3Y8_LUT4AB/NN4BEG[14] Tile_X3Y8_LUT4AB/NN4BEG[15] Tile_X3Y8_LUT4AB/NN4BEG[1]
+ Tile_X3Y8_LUT4AB/NN4BEG[2] Tile_X3Y8_LUT4AB/NN4BEG[3] Tile_X3Y8_LUT4AB/NN4BEG[4]
+ Tile_X3Y8_LUT4AB/NN4BEG[5] Tile_X3Y8_LUT4AB/NN4BEG[6] Tile_X3Y8_LUT4AB/NN4BEG[7]
+ Tile_X3Y8_LUT4AB/NN4BEG[8] Tile_X3Y8_LUT4AB/NN4BEG[9] Tile_X3Y9_S_IO4/NN4BEG[0]
+ Tile_X3Y9_S_IO4/NN4BEG[10] Tile_X3Y9_S_IO4/NN4BEG[11] Tile_X3Y9_S_IO4/NN4BEG[12]
+ Tile_X3Y9_S_IO4/NN4BEG[13] Tile_X3Y9_S_IO4/NN4BEG[14] Tile_X3Y9_S_IO4/NN4BEG[15]
+ Tile_X3Y9_S_IO4/NN4BEG[1] Tile_X3Y9_S_IO4/NN4BEG[2] Tile_X3Y9_S_IO4/NN4BEG[3] Tile_X3Y9_S_IO4/NN4BEG[4]
+ Tile_X3Y9_S_IO4/NN4BEG[5] Tile_X3Y9_S_IO4/NN4BEG[6] Tile_X3Y9_S_IO4/NN4BEG[7] Tile_X3Y9_S_IO4/NN4BEG[8]
+ Tile_X3Y9_S_IO4/NN4BEG[9] Tile_X3Y9_S_IO4/S1END[0] Tile_X3Y9_S_IO4/S1END[1] Tile_X3Y9_S_IO4/S1END[2]
+ Tile_X3Y9_S_IO4/S1END[3] Tile_X3Y8_LUT4AB/S1END[0] Tile_X3Y8_LUT4AB/S1END[1] Tile_X3Y8_LUT4AB/S1END[2]
+ Tile_X3Y8_LUT4AB/S1END[3] Tile_X3Y9_S_IO4/S2MID[0] Tile_X3Y9_S_IO4/S2MID[1] Tile_X3Y9_S_IO4/S2MID[2]
+ Tile_X3Y9_S_IO4/S2MID[3] Tile_X3Y9_S_IO4/S2MID[4] Tile_X3Y9_S_IO4/S2MID[5] Tile_X3Y9_S_IO4/S2MID[6]
+ Tile_X3Y9_S_IO4/S2MID[7] Tile_X3Y9_S_IO4/S2END[0] Tile_X3Y9_S_IO4/S2END[1] Tile_X3Y9_S_IO4/S2END[2]
+ Tile_X3Y9_S_IO4/S2END[3] Tile_X3Y9_S_IO4/S2END[4] Tile_X3Y9_S_IO4/S2END[5] Tile_X3Y9_S_IO4/S2END[6]
+ Tile_X3Y9_S_IO4/S2END[7] Tile_X3Y8_LUT4AB/S2END[0] Tile_X3Y8_LUT4AB/S2END[1] Tile_X3Y8_LUT4AB/S2END[2]
+ Tile_X3Y8_LUT4AB/S2END[3] Tile_X3Y8_LUT4AB/S2END[4] Tile_X3Y8_LUT4AB/S2END[5] Tile_X3Y8_LUT4AB/S2END[6]
+ Tile_X3Y8_LUT4AB/S2END[7] Tile_X3Y8_LUT4AB/S2MID[0] Tile_X3Y8_LUT4AB/S2MID[1] Tile_X3Y8_LUT4AB/S2MID[2]
+ Tile_X3Y8_LUT4AB/S2MID[3] Tile_X3Y8_LUT4AB/S2MID[4] Tile_X3Y8_LUT4AB/S2MID[5] Tile_X3Y8_LUT4AB/S2MID[6]
+ Tile_X3Y8_LUT4AB/S2MID[7] Tile_X3Y9_S_IO4/S4END[0] Tile_X3Y9_S_IO4/S4END[10] Tile_X3Y9_S_IO4/S4END[11]
+ Tile_X3Y9_S_IO4/S4END[12] Tile_X3Y9_S_IO4/S4END[13] Tile_X3Y9_S_IO4/S4END[14] Tile_X3Y9_S_IO4/S4END[15]
+ Tile_X3Y9_S_IO4/S4END[1] Tile_X3Y9_S_IO4/S4END[2] Tile_X3Y9_S_IO4/S4END[3] Tile_X3Y9_S_IO4/S4END[4]
+ Tile_X3Y9_S_IO4/S4END[5] Tile_X3Y9_S_IO4/S4END[6] Tile_X3Y9_S_IO4/S4END[7] Tile_X3Y9_S_IO4/S4END[8]
+ Tile_X3Y9_S_IO4/S4END[9] Tile_X3Y8_LUT4AB/S4END[0] Tile_X3Y8_LUT4AB/S4END[10] Tile_X3Y8_LUT4AB/S4END[11]
+ Tile_X3Y8_LUT4AB/S4END[12] Tile_X3Y8_LUT4AB/S4END[13] Tile_X3Y8_LUT4AB/S4END[14]
+ Tile_X3Y8_LUT4AB/S4END[15] Tile_X3Y8_LUT4AB/S4END[1] Tile_X3Y8_LUT4AB/S4END[2] Tile_X3Y8_LUT4AB/S4END[3]
+ Tile_X3Y8_LUT4AB/S4END[4] Tile_X3Y8_LUT4AB/S4END[5] Tile_X3Y8_LUT4AB/S4END[6] Tile_X3Y8_LUT4AB/S4END[7]
+ Tile_X3Y8_LUT4AB/S4END[8] Tile_X3Y8_LUT4AB/S4END[9] Tile_X3Y9_S_IO4/SS4END[0] Tile_X3Y9_S_IO4/SS4END[10]
+ Tile_X3Y9_S_IO4/SS4END[11] Tile_X3Y9_S_IO4/SS4END[12] Tile_X3Y9_S_IO4/SS4END[13]
+ Tile_X3Y9_S_IO4/SS4END[14] Tile_X3Y9_S_IO4/SS4END[15] Tile_X3Y9_S_IO4/SS4END[1]
+ Tile_X3Y9_S_IO4/SS4END[2] Tile_X3Y9_S_IO4/SS4END[3] Tile_X3Y9_S_IO4/SS4END[4] Tile_X3Y9_S_IO4/SS4END[5]
+ Tile_X3Y9_S_IO4/SS4END[6] Tile_X3Y9_S_IO4/SS4END[7] Tile_X3Y9_S_IO4/SS4END[8] Tile_X3Y9_S_IO4/SS4END[9]
+ Tile_X3Y8_LUT4AB/SS4END[0] Tile_X3Y8_LUT4AB/SS4END[10] Tile_X3Y8_LUT4AB/SS4END[11]
+ Tile_X3Y8_LUT4AB/SS4END[12] Tile_X3Y8_LUT4AB/SS4END[13] Tile_X3Y8_LUT4AB/SS4END[14]
+ Tile_X3Y8_LUT4AB/SS4END[15] Tile_X3Y8_LUT4AB/SS4END[1] Tile_X3Y8_LUT4AB/SS4END[2]
+ Tile_X3Y8_LUT4AB/SS4END[3] Tile_X3Y8_LUT4AB/SS4END[4] Tile_X3Y8_LUT4AB/SS4END[5]
+ Tile_X3Y8_LUT4AB/SS4END[6] Tile_X3Y8_LUT4AB/SS4END[7] Tile_X3Y8_LUT4AB/SS4END[8]
+ Tile_X3Y8_LUT4AB/SS4END[9] Tile_X3Y9_S_IO4/UserCLKo Tile_X3Y7_LUT4AB/UserCLK VGND
+ VPWR Tile_X3Y8_LUT4AB/W1BEG[0] Tile_X3Y8_LUT4AB/W1BEG[1] Tile_X3Y8_LUT4AB/W1BEG[2]
+ Tile_X3Y8_LUT4AB/W1BEG[3] Tile_X4Y8_LUT4AB/W1BEG[0] Tile_X4Y8_LUT4AB/W1BEG[1] Tile_X4Y8_LUT4AB/W1BEG[2]
+ Tile_X4Y8_LUT4AB/W1BEG[3] Tile_X3Y8_LUT4AB/W2BEG[0] Tile_X3Y8_LUT4AB/W2BEG[1] Tile_X3Y8_LUT4AB/W2BEG[2]
+ Tile_X3Y8_LUT4AB/W2BEG[3] Tile_X3Y8_LUT4AB/W2BEG[4] Tile_X3Y8_LUT4AB/W2BEG[5] Tile_X3Y8_LUT4AB/W2BEG[6]
+ Tile_X3Y8_LUT4AB/W2BEG[7] Tile_X2Y8_LUT4AB/W2END[0] Tile_X2Y8_LUT4AB/W2END[1] Tile_X2Y8_LUT4AB/W2END[2]
+ Tile_X2Y8_LUT4AB/W2END[3] Tile_X2Y8_LUT4AB/W2END[4] Tile_X2Y8_LUT4AB/W2END[5] Tile_X2Y8_LUT4AB/W2END[6]
+ Tile_X2Y8_LUT4AB/W2END[7] Tile_X3Y8_LUT4AB/W2END[0] Tile_X3Y8_LUT4AB/W2END[1] Tile_X3Y8_LUT4AB/W2END[2]
+ Tile_X3Y8_LUT4AB/W2END[3] Tile_X3Y8_LUT4AB/W2END[4] Tile_X3Y8_LUT4AB/W2END[5] Tile_X3Y8_LUT4AB/W2END[6]
+ Tile_X3Y8_LUT4AB/W2END[7] Tile_X4Y8_LUT4AB/W2BEG[0] Tile_X4Y8_LUT4AB/W2BEG[1] Tile_X4Y8_LUT4AB/W2BEG[2]
+ Tile_X4Y8_LUT4AB/W2BEG[3] Tile_X4Y8_LUT4AB/W2BEG[4] Tile_X4Y8_LUT4AB/W2BEG[5] Tile_X4Y8_LUT4AB/W2BEG[6]
+ Tile_X4Y8_LUT4AB/W2BEG[7] Tile_X3Y8_LUT4AB/W6BEG[0] Tile_X3Y8_LUT4AB/W6BEG[10] Tile_X3Y8_LUT4AB/W6BEG[11]
+ Tile_X3Y8_LUT4AB/W6BEG[1] Tile_X3Y8_LUT4AB/W6BEG[2] Tile_X3Y8_LUT4AB/W6BEG[3] Tile_X3Y8_LUT4AB/W6BEG[4]
+ Tile_X3Y8_LUT4AB/W6BEG[5] Tile_X3Y8_LUT4AB/W6BEG[6] Tile_X3Y8_LUT4AB/W6BEG[7] Tile_X3Y8_LUT4AB/W6BEG[8]
+ Tile_X3Y8_LUT4AB/W6BEG[9] Tile_X4Y8_LUT4AB/W6BEG[0] Tile_X4Y8_LUT4AB/W6BEG[10] Tile_X4Y8_LUT4AB/W6BEG[11]
+ Tile_X4Y8_LUT4AB/W6BEG[1] Tile_X4Y8_LUT4AB/W6BEG[2] Tile_X4Y8_LUT4AB/W6BEG[3] Tile_X4Y8_LUT4AB/W6BEG[4]
+ Tile_X4Y8_LUT4AB/W6BEG[5] Tile_X4Y8_LUT4AB/W6BEG[6] Tile_X4Y8_LUT4AB/W6BEG[7] Tile_X4Y8_LUT4AB/W6BEG[8]
+ Tile_X4Y8_LUT4AB/W6BEG[9] Tile_X3Y8_LUT4AB/WW4BEG[0] Tile_X3Y8_LUT4AB/WW4BEG[10]
+ Tile_X3Y8_LUT4AB/WW4BEG[11] Tile_X3Y8_LUT4AB/WW4BEG[12] Tile_X3Y8_LUT4AB/WW4BEG[13]
+ Tile_X3Y8_LUT4AB/WW4BEG[14] Tile_X3Y8_LUT4AB/WW4BEG[15] Tile_X3Y8_LUT4AB/WW4BEG[1]
+ Tile_X3Y8_LUT4AB/WW4BEG[2] Tile_X3Y8_LUT4AB/WW4BEG[3] Tile_X3Y8_LUT4AB/WW4BEG[4]
+ Tile_X3Y8_LUT4AB/WW4BEG[5] Tile_X3Y8_LUT4AB/WW4BEG[6] Tile_X3Y8_LUT4AB/WW4BEG[7]
+ Tile_X3Y8_LUT4AB/WW4BEG[8] Tile_X3Y8_LUT4AB/WW4BEG[9] Tile_X4Y8_LUT4AB/WW4BEG[0]
+ Tile_X4Y8_LUT4AB/WW4BEG[10] Tile_X4Y8_LUT4AB/WW4BEG[11] Tile_X4Y8_LUT4AB/WW4BEG[12]
+ Tile_X4Y8_LUT4AB/WW4BEG[13] Tile_X4Y8_LUT4AB/WW4BEG[14] Tile_X4Y8_LUT4AB/WW4BEG[15]
+ Tile_X4Y8_LUT4AB/WW4BEG[1] Tile_X4Y8_LUT4AB/WW4BEG[2] Tile_X4Y8_LUT4AB/WW4BEG[3]
+ Tile_X4Y8_LUT4AB/WW4BEG[4] Tile_X4Y8_LUT4AB/WW4BEG[5] Tile_X4Y8_LUT4AB/WW4BEG[6]
+ Tile_X4Y8_LUT4AB/WW4BEG[7] Tile_X4Y8_LUT4AB/WW4BEG[8] Tile_X4Y8_LUT4AB/WW4BEG[9]
+ LUT4AB
XTile_X3Y0_N_IO4 Tile_X3Y0_A_I_top Tile_X3Y0_A_O_top Tile_X3Y0_A_T_top Tile_X3Y0_B_I_top
+ Tile_X3Y0_B_O_top Tile_X3Y0_B_T_top Tile_X3Y0_C_I_top Tile_X3Y0_C_O_top Tile_X3Y0_C_T_top
+ Tile_X3Y0_N_IO4/Ci Tile_X3Y0_D_I_top Tile_X3Y0_D_O_top Tile_X3Y0_D_T_top Tile_X3Y0_N_IO4/FrameData[0]
+ Tile_X3Y0_N_IO4/FrameData[10] Tile_X3Y0_N_IO4/FrameData[11] Tile_X3Y0_N_IO4/FrameData[12]
+ Tile_X3Y0_N_IO4/FrameData[13] Tile_X3Y0_N_IO4/FrameData[14] Tile_X3Y0_N_IO4/FrameData[15]
+ Tile_X3Y0_N_IO4/FrameData[16] Tile_X3Y0_N_IO4/FrameData[17] Tile_X3Y0_N_IO4/FrameData[18]
+ Tile_X3Y0_N_IO4/FrameData[19] Tile_X3Y0_N_IO4/FrameData[1] Tile_X3Y0_N_IO4/FrameData[20]
+ Tile_X3Y0_N_IO4/FrameData[21] Tile_X3Y0_N_IO4/FrameData[22] Tile_X3Y0_N_IO4/FrameData[23]
+ Tile_X3Y0_N_IO4/FrameData[24] Tile_X3Y0_N_IO4/FrameData[25] Tile_X3Y0_N_IO4/FrameData[26]
+ Tile_X3Y0_N_IO4/FrameData[27] Tile_X3Y0_N_IO4/FrameData[28] Tile_X3Y0_N_IO4/FrameData[29]
+ Tile_X3Y0_N_IO4/FrameData[2] Tile_X3Y0_N_IO4/FrameData[30] Tile_X3Y0_N_IO4/FrameData[31]
+ Tile_X3Y0_N_IO4/FrameData[3] Tile_X3Y0_N_IO4/FrameData[4] Tile_X3Y0_N_IO4/FrameData[5]
+ Tile_X3Y0_N_IO4/FrameData[6] Tile_X3Y0_N_IO4/FrameData[7] Tile_X3Y0_N_IO4/FrameData[8]
+ Tile_X3Y0_N_IO4/FrameData[9] Tile_X4Y0_N_IO4/FrameData[0] Tile_X4Y0_N_IO4/FrameData[10]
+ Tile_X4Y0_N_IO4/FrameData[11] Tile_X4Y0_N_IO4/FrameData[12] Tile_X4Y0_N_IO4/FrameData[13]
+ Tile_X4Y0_N_IO4/FrameData[14] Tile_X4Y0_N_IO4/FrameData[15] Tile_X4Y0_N_IO4/FrameData[16]
+ Tile_X4Y0_N_IO4/FrameData[17] Tile_X4Y0_N_IO4/FrameData[18] Tile_X4Y0_N_IO4/FrameData[19]
+ Tile_X4Y0_N_IO4/FrameData[1] Tile_X4Y0_N_IO4/FrameData[20] Tile_X4Y0_N_IO4/FrameData[21]
+ Tile_X4Y0_N_IO4/FrameData[22] Tile_X4Y0_N_IO4/FrameData[23] Tile_X4Y0_N_IO4/FrameData[24]
+ Tile_X4Y0_N_IO4/FrameData[25] Tile_X4Y0_N_IO4/FrameData[26] Tile_X4Y0_N_IO4/FrameData[27]
+ Tile_X4Y0_N_IO4/FrameData[28] Tile_X4Y0_N_IO4/FrameData[29] Tile_X4Y0_N_IO4/FrameData[2]
+ Tile_X4Y0_N_IO4/FrameData[30] Tile_X4Y0_N_IO4/FrameData[31] Tile_X4Y0_N_IO4/FrameData[3]
+ Tile_X4Y0_N_IO4/FrameData[4] Tile_X4Y0_N_IO4/FrameData[5] Tile_X4Y0_N_IO4/FrameData[6]
+ Tile_X4Y0_N_IO4/FrameData[7] Tile_X4Y0_N_IO4/FrameData[8] Tile_X4Y0_N_IO4/FrameData[9]
+ Tile_X3Y0_N_IO4/FrameStrobe[0] Tile_X3Y0_N_IO4/FrameStrobe[10] Tile_X3Y0_N_IO4/FrameStrobe[11]
+ Tile_X3Y0_N_IO4/FrameStrobe[12] Tile_X3Y0_N_IO4/FrameStrobe[13] Tile_X3Y0_N_IO4/FrameStrobe[14]
+ Tile_X3Y0_N_IO4/FrameStrobe[15] Tile_X3Y0_N_IO4/FrameStrobe[16] Tile_X3Y0_N_IO4/FrameStrobe[17]
+ Tile_X3Y0_N_IO4/FrameStrobe[18] Tile_X3Y0_N_IO4/FrameStrobe[19] Tile_X3Y0_N_IO4/FrameStrobe[1]
+ Tile_X3Y0_N_IO4/FrameStrobe[2] Tile_X3Y0_N_IO4/FrameStrobe[3] Tile_X3Y0_N_IO4/FrameStrobe[4]
+ Tile_X3Y0_N_IO4/FrameStrobe[5] Tile_X3Y0_N_IO4/FrameStrobe[6] Tile_X3Y0_N_IO4/FrameStrobe[7]
+ Tile_X3Y0_N_IO4/FrameStrobe[8] Tile_X3Y0_N_IO4/FrameStrobe[9] Tile_X3Y0_N_IO4/FrameStrobe_O[0]
+ Tile_X3Y0_N_IO4/FrameStrobe_O[10] Tile_X3Y0_N_IO4/FrameStrobe_O[11] Tile_X3Y0_N_IO4/FrameStrobe_O[12]
+ Tile_X3Y0_N_IO4/FrameStrobe_O[13] Tile_X3Y0_N_IO4/FrameStrobe_O[14] Tile_X3Y0_N_IO4/FrameStrobe_O[15]
+ Tile_X3Y0_N_IO4/FrameStrobe_O[16] Tile_X3Y0_N_IO4/FrameStrobe_O[17] Tile_X3Y0_N_IO4/FrameStrobe_O[18]
+ Tile_X3Y0_N_IO4/FrameStrobe_O[19] Tile_X3Y0_N_IO4/FrameStrobe_O[1] Tile_X3Y0_N_IO4/FrameStrobe_O[2]
+ Tile_X3Y0_N_IO4/FrameStrobe_O[3] Tile_X3Y0_N_IO4/FrameStrobe_O[4] Tile_X3Y0_N_IO4/FrameStrobe_O[5]
+ Tile_X3Y0_N_IO4/FrameStrobe_O[6] Tile_X3Y0_N_IO4/FrameStrobe_O[7] Tile_X3Y0_N_IO4/FrameStrobe_O[8]
+ Tile_X3Y0_N_IO4/FrameStrobe_O[9] Tile_X3Y0_N_IO4/N1END[0] Tile_X3Y0_N_IO4/N1END[1]
+ Tile_X3Y0_N_IO4/N1END[2] Tile_X3Y0_N_IO4/N1END[3] Tile_X3Y0_N_IO4/N2END[0] Tile_X3Y0_N_IO4/N2END[1]
+ Tile_X3Y0_N_IO4/N2END[2] Tile_X3Y0_N_IO4/N2END[3] Tile_X3Y0_N_IO4/N2END[4] Tile_X3Y0_N_IO4/N2END[5]
+ Tile_X3Y0_N_IO4/N2END[6] Tile_X3Y0_N_IO4/N2END[7] Tile_X3Y0_N_IO4/N2MID[0] Tile_X3Y0_N_IO4/N2MID[1]
+ Tile_X3Y0_N_IO4/N2MID[2] Tile_X3Y0_N_IO4/N2MID[3] Tile_X3Y0_N_IO4/N2MID[4] Tile_X3Y0_N_IO4/N2MID[5]
+ Tile_X3Y0_N_IO4/N2MID[6] Tile_X3Y0_N_IO4/N2MID[7] Tile_X3Y0_N_IO4/N4END[0] Tile_X3Y0_N_IO4/N4END[10]
+ Tile_X3Y0_N_IO4/N4END[11] Tile_X3Y0_N_IO4/N4END[12] Tile_X3Y0_N_IO4/N4END[13] Tile_X3Y0_N_IO4/N4END[14]
+ Tile_X3Y0_N_IO4/N4END[15] Tile_X3Y0_N_IO4/N4END[1] Tile_X3Y0_N_IO4/N4END[2] Tile_X3Y0_N_IO4/N4END[3]
+ Tile_X3Y0_N_IO4/N4END[4] Tile_X3Y0_N_IO4/N4END[5] Tile_X3Y0_N_IO4/N4END[6] Tile_X3Y0_N_IO4/N4END[7]
+ Tile_X3Y0_N_IO4/N4END[8] Tile_X3Y0_N_IO4/N4END[9] Tile_X3Y0_N_IO4/NN4END[0] Tile_X3Y0_N_IO4/NN4END[10]
+ Tile_X3Y0_N_IO4/NN4END[11] Tile_X3Y0_N_IO4/NN4END[12] Tile_X3Y0_N_IO4/NN4END[13]
+ Tile_X3Y0_N_IO4/NN4END[14] Tile_X3Y0_N_IO4/NN4END[15] Tile_X3Y0_N_IO4/NN4END[1]
+ Tile_X3Y0_N_IO4/NN4END[2] Tile_X3Y0_N_IO4/NN4END[3] Tile_X3Y0_N_IO4/NN4END[4] Tile_X3Y0_N_IO4/NN4END[5]
+ Tile_X3Y0_N_IO4/NN4END[6] Tile_X3Y0_N_IO4/NN4END[7] Tile_X3Y0_N_IO4/NN4END[8] Tile_X3Y0_N_IO4/NN4END[9]
+ Tile_X3Y0_N_IO4/S1BEG[0] Tile_X3Y0_N_IO4/S1BEG[1] Tile_X3Y0_N_IO4/S1BEG[2] Tile_X3Y0_N_IO4/S1BEG[3]
+ Tile_X3Y0_N_IO4/S2BEG[0] Tile_X3Y0_N_IO4/S2BEG[1] Tile_X3Y0_N_IO4/S2BEG[2] Tile_X3Y0_N_IO4/S2BEG[3]
+ Tile_X3Y0_N_IO4/S2BEG[4] Tile_X3Y0_N_IO4/S2BEG[5] Tile_X3Y0_N_IO4/S2BEG[6] Tile_X3Y0_N_IO4/S2BEG[7]
+ Tile_X3Y1_LUT4AB/S2END[0] Tile_X3Y1_LUT4AB/S2END[1] Tile_X3Y1_LUT4AB/S2END[2] Tile_X3Y1_LUT4AB/S2END[3]
+ Tile_X3Y1_LUT4AB/S2END[4] Tile_X3Y1_LUT4AB/S2END[5] Tile_X3Y1_LUT4AB/S2END[6] Tile_X3Y1_LUT4AB/S2END[7]
+ Tile_X3Y0_N_IO4/S4BEG[0] Tile_X3Y0_N_IO4/S4BEG[10] Tile_X3Y0_N_IO4/S4BEG[11] Tile_X3Y0_N_IO4/S4BEG[12]
+ Tile_X3Y0_N_IO4/S4BEG[13] Tile_X3Y0_N_IO4/S4BEG[14] Tile_X3Y0_N_IO4/S4BEG[15] Tile_X3Y0_N_IO4/S4BEG[1]
+ Tile_X3Y0_N_IO4/S4BEG[2] Tile_X3Y0_N_IO4/S4BEG[3] Tile_X3Y0_N_IO4/S4BEG[4] Tile_X3Y0_N_IO4/S4BEG[5]
+ Tile_X3Y0_N_IO4/S4BEG[6] Tile_X3Y0_N_IO4/S4BEG[7] Tile_X3Y0_N_IO4/S4BEG[8] Tile_X3Y0_N_IO4/S4BEG[9]
+ Tile_X3Y0_N_IO4/SS4BEG[0] Tile_X3Y0_N_IO4/SS4BEG[10] Tile_X3Y0_N_IO4/SS4BEG[11]
+ Tile_X3Y0_N_IO4/SS4BEG[12] Tile_X3Y0_N_IO4/SS4BEG[13] Tile_X3Y0_N_IO4/SS4BEG[14]
+ Tile_X3Y0_N_IO4/SS4BEG[15] Tile_X3Y0_N_IO4/SS4BEG[1] Tile_X3Y0_N_IO4/SS4BEG[2] Tile_X3Y0_N_IO4/SS4BEG[3]
+ Tile_X3Y0_N_IO4/SS4BEG[4] Tile_X3Y0_N_IO4/SS4BEG[5] Tile_X3Y0_N_IO4/SS4BEG[6] Tile_X3Y0_N_IO4/SS4BEG[7]
+ Tile_X3Y0_N_IO4/SS4BEG[8] Tile_X3Y0_N_IO4/SS4BEG[9] Tile_X3Y0_N_IO4/UserCLK Tile_X3Y0_N_IO4/UserCLKo
+ VGND VPWR N_IO4
XTile_X2Y1_LUT4AB Tile_X2Y2_LUT4AB/Co Tile_X2Y0_N_IO4/Ci Tile_X3Y1_LUT4AB/E1END[0]
+ Tile_X3Y1_LUT4AB/E1END[1] Tile_X3Y1_LUT4AB/E1END[2] Tile_X3Y1_LUT4AB/E1END[3] Tile_X2Y1_LUT4AB/E1END[0]
+ Tile_X2Y1_LUT4AB/E1END[1] Tile_X2Y1_LUT4AB/E1END[2] Tile_X2Y1_LUT4AB/E1END[3] Tile_X3Y1_LUT4AB/E2MID[0]
+ Tile_X3Y1_LUT4AB/E2MID[1] Tile_X3Y1_LUT4AB/E2MID[2] Tile_X3Y1_LUT4AB/E2MID[3] Tile_X3Y1_LUT4AB/E2MID[4]
+ Tile_X3Y1_LUT4AB/E2MID[5] Tile_X3Y1_LUT4AB/E2MID[6] Tile_X3Y1_LUT4AB/E2MID[7] Tile_X3Y1_LUT4AB/E2END[0]
+ Tile_X3Y1_LUT4AB/E2END[1] Tile_X3Y1_LUT4AB/E2END[2] Tile_X3Y1_LUT4AB/E2END[3] Tile_X3Y1_LUT4AB/E2END[4]
+ Tile_X3Y1_LUT4AB/E2END[5] Tile_X3Y1_LUT4AB/E2END[6] Tile_X3Y1_LUT4AB/E2END[7] Tile_X2Y1_LUT4AB/E2END[0]
+ Tile_X2Y1_LUT4AB/E2END[1] Tile_X2Y1_LUT4AB/E2END[2] Tile_X2Y1_LUT4AB/E2END[3] Tile_X2Y1_LUT4AB/E2END[4]
+ Tile_X2Y1_LUT4AB/E2END[5] Tile_X2Y1_LUT4AB/E2END[6] Tile_X2Y1_LUT4AB/E2END[7] Tile_X2Y1_LUT4AB/E2MID[0]
+ Tile_X2Y1_LUT4AB/E2MID[1] Tile_X2Y1_LUT4AB/E2MID[2] Tile_X2Y1_LUT4AB/E2MID[3] Tile_X2Y1_LUT4AB/E2MID[4]
+ Tile_X2Y1_LUT4AB/E2MID[5] Tile_X2Y1_LUT4AB/E2MID[6] Tile_X2Y1_LUT4AB/E2MID[7] Tile_X3Y1_LUT4AB/E6END[0]
+ Tile_X3Y1_LUT4AB/E6END[10] Tile_X3Y1_LUT4AB/E6END[11] Tile_X3Y1_LUT4AB/E6END[1]
+ Tile_X3Y1_LUT4AB/E6END[2] Tile_X3Y1_LUT4AB/E6END[3] Tile_X3Y1_LUT4AB/E6END[4] Tile_X3Y1_LUT4AB/E6END[5]
+ Tile_X3Y1_LUT4AB/E6END[6] Tile_X3Y1_LUT4AB/E6END[7] Tile_X3Y1_LUT4AB/E6END[8] Tile_X3Y1_LUT4AB/E6END[9]
+ Tile_X2Y1_LUT4AB/E6END[0] Tile_X2Y1_LUT4AB/E6END[10] Tile_X2Y1_LUT4AB/E6END[11]
+ Tile_X2Y1_LUT4AB/E6END[1] Tile_X2Y1_LUT4AB/E6END[2] Tile_X2Y1_LUT4AB/E6END[3] Tile_X2Y1_LUT4AB/E6END[4]
+ Tile_X2Y1_LUT4AB/E6END[5] Tile_X2Y1_LUT4AB/E6END[6] Tile_X2Y1_LUT4AB/E6END[7] Tile_X2Y1_LUT4AB/E6END[8]
+ Tile_X2Y1_LUT4AB/E6END[9] Tile_X3Y1_LUT4AB/EE4END[0] Tile_X3Y1_LUT4AB/EE4END[10]
+ Tile_X3Y1_LUT4AB/EE4END[11] Tile_X3Y1_LUT4AB/EE4END[12] Tile_X3Y1_LUT4AB/EE4END[13]
+ Tile_X3Y1_LUT4AB/EE4END[14] Tile_X3Y1_LUT4AB/EE4END[15] Tile_X3Y1_LUT4AB/EE4END[1]
+ Tile_X3Y1_LUT4AB/EE4END[2] Tile_X3Y1_LUT4AB/EE4END[3] Tile_X3Y1_LUT4AB/EE4END[4]
+ Tile_X3Y1_LUT4AB/EE4END[5] Tile_X3Y1_LUT4AB/EE4END[6] Tile_X3Y1_LUT4AB/EE4END[7]
+ Tile_X3Y1_LUT4AB/EE4END[8] Tile_X3Y1_LUT4AB/EE4END[9] Tile_X2Y1_LUT4AB/EE4END[0]
+ Tile_X2Y1_LUT4AB/EE4END[10] Tile_X2Y1_LUT4AB/EE4END[11] Tile_X2Y1_LUT4AB/EE4END[12]
+ Tile_X2Y1_LUT4AB/EE4END[13] Tile_X2Y1_LUT4AB/EE4END[14] Tile_X2Y1_LUT4AB/EE4END[15]
+ Tile_X2Y1_LUT4AB/EE4END[1] Tile_X2Y1_LUT4AB/EE4END[2] Tile_X2Y1_LUT4AB/EE4END[3]
+ Tile_X2Y1_LUT4AB/EE4END[4] Tile_X2Y1_LUT4AB/EE4END[5] Tile_X2Y1_LUT4AB/EE4END[6]
+ Tile_X2Y1_LUT4AB/EE4END[7] Tile_X2Y1_LUT4AB/EE4END[8] Tile_X2Y1_LUT4AB/EE4END[9]
+ Tile_X2Y1_LUT4AB/FrameData[0] Tile_X2Y1_LUT4AB/FrameData[10] Tile_X2Y1_LUT4AB/FrameData[11]
+ Tile_X2Y1_LUT4AB/FrameData[12] Tile_X2Y1_LUT4AB/FrameData[13] Tile_X2Y1_LUT4AB/FrameData[14]
+ Tile_X2Y1_LUT4AB/FrameData[15] Tile_X2Y1_LUT4AB/FrameData[16] Tile_X2Y1_LUT4AB/FrameData[17]
+ Tile_X2Y1_LUT4AB/FrameData[18] Tile_X2Y1_LUT4AB/FrameData[19] Tile_X2Y1_LUT4AB/FrameData[1]
+ Tile_X2Y1_LUT4AB/FrameData[20] Tile_X2Y1_LUT4AB/FrameData[21] Tile_X2Y1_LUT4AB/FrameData[22]
+ Tile_X2Y1_LUT4AB/FrameData[23] Tile_X2Y1_LUT4AB/FrameData[24] Tile_X2Y1_LUT4AB/FrameData[25]
+ Tile_X2Y1_LUT4AB/FrameData[26] Tile_X2Y1_LUT4AB/FrameData[27] Tile_X2Y1_LUT4AB/FrameData[28]
+ Tile_X2Y1_LUT4AB/FrameData[29] Tile_X2Y1_LUT4AB/FrameData[2] Tile_X2Y1_LUT4AB/FrameData[30]
+ Tile_X2Y1_LUT4AB/FrameData[31] Tile_X2Y1_LUT4AB/FrameData[3] Tile_X2Y1_LUT4AB/FrameData[4]
+ Tile_X2Y1_LUT4AB/FrameData[5] Tile_X2Y1_LUT4AB/FrameData[6] Tile_X2Y1_LUT4AB/FrameData[7]
+ Tile_X2Y1_LUT4AB/FrameData[8] Tile_X2Y1_LUT4AB/FrameData[9] Tile_X3Y1_LUT4AB/FrameData[0]
+ Tile_X3Y1_LUT4AB/FrameData[10] Tile_X3Y1_LUT4AB/FrameData[11] Tile_X3Y1_LUT4AB/FrameData[12]
+ Tile_X3Y1_LUT4AB/FrameData[13] Tile_X3Y1_LUT4AB/FrameData[14] Tile_X3Y1_LUT4AB/FrameData[15]
+ Tile_X3Y1_LUT4AB/FrameData[16] Tile_X3Y1_LUT4AB/FrameData[17] Tile_X3Y1_LUT4AB/FrameData[18]
+ Tile_X3Y1_LUT4AB/FrameData[19] Tile_X3Y1_LUT4AB/FrameData[1] Tile_X3Y1_LUT4AB/FrameData[20]
+ Tile_X3Y1_LUT4AB/FrameData[21] Tile_X3Y1_LUT4AB/FrameData[22] Tile_X3Y1_LUT4AB/FrameData[23]
+ Tile_X3Y1_LUT4AB/FrameData[24] Tile_X3Y1_LUT4AB/FrameData[25] Tile_X3Y1_LUT4AB/FrameData[26]
+ Tile_X3Y1_LUT4AB/FrameData[27] Tile_X3Y1_LUT4AB/FrameData[28] Tile_X3Y1_LUT4AB/FrameData[29]
+ Tile_X3Y1_LUT4AB/FrameData[2] Tile_X3Y1_LUT4AB/FrameData[30] Tile_X3Y1_LUT4AB/FrameData[31]
+ Tile_X3Y1_LUT4AB/FrameData[3] Tile_X3Y1_LUT4AB/FrameData[4] Tile_X3Y1_LUT4AB/FrameData[5]
+ Tile_X3Y1_LUT4AB/FrameData[6] Tile_X3Y1_LUT4AB/FrameData[7] Tile_X3Y1_LUT4AB/FrameData[8]
+ Tile_X3Y1_LUT4AB/FrameData[9] Tile_X2Y1_LUT4AB/FrameStrobe[0] Tile_X2Y1_LUT4AB/FrameStrobe[10]
+ Tile_X2Y1_LUT4AB/FrameStrobe[11] Tile_X2Y1_LUT4AB/FrameStrobe[12] Tile_X2Y1_LUT4AB/FrameStrobe[13]
+ Tile_X2Y1_LUT4AB/FrameStrobe[14] Tile_X2Y1_LUT4AB/FrameStrobe[15] Tile_X2Y1_LUT4AB/FrameStrobe[16]
+ Tile_X2Y1_LUT4AB/FrameStrobe[17] Tile_X2Y1_LUT4AB/FrameStrobe[18] Tile_X2Y1_LUT4AB/FrameStrobe[19]
+ Tile_X2Y1_LUT4AB/FrameStrobe[1] Tile_X2Y1_LUT4AB/FrameStrobe[2] Tile_X2Y1_LUT4AB/FrameStrobe[3]
+ Tile_X2Y1_LUT4AB/FrameStrobe[4] Tile_X2Y1_LUT4AB/FrameStrobe[5] Tile_X2Y1_LUT4AB/FrameStrobe[6]
+ Tile_X2Y1_LUT4AB/FrameStrobe[7] Tile_X2Y1_LUT4AB/FrameStrobe[8] Tile_X2Y1_LUT4AB/FrameStrobe[9]
+ Tile_X2Y0_N_IO4/FrameStrobe[0] Tile_X2Y0_N_IO4/FrameStrobe[10] Tile_X2Y0_N_IO4/FrameStrobe[11]
+ Tile_X2Y0_N_IO4/FrameStrobe[12] Tile_X2Y0_N_IO4/FrameStrobe[13] Tile_X2Y0_N_IO4/FrameStrobe[14]
+ Tile_X2Y0_N_IO4/FrameStrobe[15] Tile_X2Y0_N_IO4/FrameStrobe[16] Tile_X2Y0_N_IO4/FrameStrobe[17]
+ Tile_X2Y0_N_IO4/FrameStrobe[18] Tile_X2Y0_N_IO4/FrameStrobe[19] Tile_X2Y0_N_IO4/FrameStrobe[1]
+ Tile_X2Y0_N_IO4/FrameStrobe[2] Tile_X2Y0_N_IO4/FrameStrobe[3] Tile_X2Y0_N_IO4/FrameStrobe[4]
+ Tile_X2Y0_N_IO4/FrameStrobe[5] Tile_X2Y0_N_IO4/FrameStrobe[6] Tile_X2Y0_N_IO4/FrameStrobe[7]
+ Tile_X2Y0_N_IO4/FrameStrobe[8] Tile_X2Y0_N_IO4/FrameStrobe[9] Tile_X2Y0_N_IO4/N1END[0]
+ Tile_X2Y0_N_IO4/N1END[1] Tile_X2Y0_N_IO4/N1END[2] Tile_X2Y0_N_IO4/N1END[3] Tile_X2Y2_LUT4AB/N1BEG[0]
+ Tile_X2Y2_LUT4AB/N1BEG[1] Tile_X2Y2_LUT4AB/N1BEG[2] Tile_X2Y2_LUT4AB/N1BEG[3] Tile_X2Y0_N_IO4/N2MID[0]
+ Tile_X2Y0_N_IO4/N2MID[1] Tile_X2Y0_N_IO4/N2MID[2] Tile_X2Y0_N_IO4/N2MID[3] Tile_X2Y0_N_IO4/N2MID[4]
+ Tile_X2Y0_N_IO4/N2MID[5] Tile_X2Y0_N_IO4/N2MID[6] Tile_X2Y0_N_IO4/N2MID[7] Tile_X2Y0_N_IO4/N2END[0]
+ Tile_X2Y0_N_IO4/N2END[1] Tile_X2Y0_N_IO4/N2END[2] Tile_X2Y0_N_IO4/N2END[3] Tile_X2Y0_N_IO4/N2END[4]
+ Tile_X2Y0_N_IO4/N2END[5] Tile_X2Y0_N_IO4/N2END[6] Tile_X2Y0_N_IO4/N2END[7] Tile_X2Y1_LUT4AB/N2END[0]
+ Tile_X2Y1_LUT4AB/N2END[1] Tile_X2Y1_LUT4AB/N2END[2] Tile_X2Y1_LUT4AB/N2END[3] Tile_X2Y1_LUT4AB/N2END[4]
+ Tile_X2Y1_LUT4AB/N2END[5] Tile_X2Y1_LUT4AB/N2END[6] Tile_X2Y1_LUT4AB/N2END[7] Tile_X2Y2_LUT4AB/N2BEG[0]
+ Tile_X2Y2_LUT4AB/N2BEG[1] Tile_X2Y2_LUT4AB/N2BEG[2] Tile_X2Y2_LUT4AB/N2BEG[3] Tile_X2Y2_LUT4AB/N2BEG[4]
+ Tile_X2Y2_LUT4AB/N2BEG[5] Tile_X2Y2_LUT4AB/N2BEG[6] Tile_X2Y2_LUT4AB/N2BEG[7] Tile_X2Y0_N_IO4/N4END[0]
+ Tile_X2Y0_N_IO4/N4END[10] Tile_X2Y0_N_IO4/N4END[11] Tile_X2Y0_N_IO4/N4END[12] Tile_X2Y0_N_IO4/N4END[13]
+ Tile_X2Y0_N_IO4/N4END[14] Tile_X2Y0_N_IO4/N4END[15] Tile_X2Y0_N_IO4/N4END[1] Tile_X2Y0_N_IO4/N4END[2]
+ Tile_X2Y0_N_IO4/N4END[3] Tile_X2Y0_N_IO4/N4END[4] Tile_X2Y0_N_IO4/N4END[5] Tile_X2Y0_N_IO4/N4END[6]
+ Tile_X2Y0_N_IO4/N4END[7] Tile_X2Y0_N_IO4/N4END[8] Tile_X2Y0_N_IO4/N4END[9] Tile_X2Y2_LUT4AB/N4BEG[0]
+ Tile_X2Y2_LUT4AB/N4BEG[10] Tile_X2Y2_LUT4AB/N4BEG[11] Tile_X2Y2_LUT4AB/N4BEG[12]
+ Tile_X2Y2_LUT4AB/N4BEG[13] Tile_X2Y2_LUT4AB/N4BEG[14] Tile_X2Y2_LUT4AB/N4BEG[15]
+ Tile_X2Y2_LUT4AB/N4BEG[1] Tile_X2Y2_LUT4AB/N4BEG[2] Tile_X2Y2_LUT4AB/N4BEG[3] Tile_X2Y2_LUT4AB/N4BEG[4]
+ Tile_X2Y2_LUT4AB/N4BEG[5] Tile_X2Y2_LUT4AB/N4BEG[6] Tile_X2Y2_LUT4AB/N4BEG[7] Tile_X2Y2_LUT4AB/N4BEG[8]
+ Tile_X2Y2_LUT4AB/N4BEG[9] Tile_X2Y0_N_IO4/NN4END[0] Tile_X2Y0_N_IO4/NN4END[10] Tile_X2Y0_N_IO4/NN4END[11]
+ Tile_X2Y0_N_IO4/NN4END[12] Tile_X2Y0_N_IO4/NN4END[13] Tile_X2Y0_N_IO4/NN4END[14]
+ Tile_X2Y0_N_IO4/NN4END[15] Tile_X2Y0_N_IO4/NN4END[1] Tile_X2Y0_N_IO4/NN4END[2] Tile_X2Y0_N_IO4/NN4END[3]
+ Tile_X2Y0_N_IO4/NN4END[4] Tile_X2Y0_N_IO4/NN4END[5] Tile_X2Y0_N_IO4/NN4END[6] Tile_X2Y0_N_IO4/NN4END[7]
+ Tile_X2Y0_N_IO4/NN4END[8] Tile_X2Y0_N_IO4/NN4END[9] Tile_X2Y2_LUT4AB/NN4BEG[0] Tile_X2Y2_LUT4AB/NN4BEG[10]
+ Tile_X2Y2_LUT4AB/NN4BEG[11] Tile_X2Y2_LUT4AB/NN4BEG[12] Tile_X2Y2_LUT4AB/NN4BEG[13]
+ Tile_X2Y2_LUT4AB/NN4BEG[14] Tile_X2Y2_LUT4AB/NN4BEG[15] Tile_X2Y2_LUT4AB/NN4BEG[1]
+ Tile_X2Y2_LUT4AB/NN4BEG[2] Tile_X2Y2_LUT4AB/NN4BEG[3] Tile_X2Y2_LUT4AB/NN4BEG[4]
+ Tile_X2Y2_LUT4AB/NN4BEG[5] Tile_X2Y2_LUT4AB/NN4BEG[6] Tile_X2Y2_LUT4AB/NN4BEG[7]
+ Tile_X2Y2_LUT4AB/NN4BEG[8] Tile_X2Y2_LUT4AB/NN4BEG[9] Tile_X2Y2_LUT4AB/S1END[0]
+ Tile_X2Y2_LUT4AB/S1END[1] Tile_X2Y2_LUT4AB/S1END[2] Tile_X2Y2_LUT4AB/S1END[3] Tile_X2Y0_N_IO4/S1BEG[0]
+ Tile_X2Y0_N_IO4/S1BEG[1] Tile_X2Y0_N_IO4/S1BEG[2] Tile_X2Y0_N_IO4/S1BEG[3] Tile_X2Y2_LUT4AB/S2MID[0]
+ Tile_X2Y2_LUT4AB/S2MID[1] Tile_X2Y2_LUT4AB/S2MID[2] Tile_X2Y2_LUT4AB/S2MID[3] Tile_X2Y2_LUT4AB/S2MID[4]
+ Tile_X2Y2_LUT4AB/S2MID[5] Tile_X2Y2_LUT4AB/S2MID[6] Tile_X2Y2_LUT4AB/S2MID[7] Tile_X2Y2_LUT4AB/S2END[0]
+ Tile_X2Y2_LUT4AB/S2END[1] Tile_X2Y2_LUT4AB/S2END[2] Tile_X2Y2_LUT4AB/S2END[3] Tile_X2Y2_LUT4AB/S2END[4]
+ Tile_X2Y2_LUT4AB/S2END[5] Tile_X2Y2_LUT4AB/S2END[6] Tile_X2Y2_LUT4AB/S2END[7] Tile_X2Y1_LUT4AB/S2END[0]
+ Tile_X2Y1_LUT4AB/S2END[1] Tile_X2Y1_LUT4AB/S2END[2] Tile_X2Y1_LUT4AB/S2END[3] Tile_X2Y1_LUT4AB/S2END[4]
+ Tile_X2Y1_LUT4AB/S2END[5] Tile_X2Y1_LUT4AB/S2END[6] Tile_X2Y1_LUT4AB/S2END[7] Tile_X2Y0_N_IO4/S2BEG[0]
+ Tile_X2Y0_N_IO4/S2BEG[1] Tile_X2Y0_N_IO4/S2BEG[2] Tile_X2Y0_N_IO4/S2BEG[3] Tile_X2Y0_N_IO4/S2BEG[4]
+ Tile_X2Y0_N_IO4/S2BEG[5] Tile_X2Y0_N_IO4/S2BEG[6] Tile_X2Y0_N_IO4/S2BEG[7] Tile_X2Y2_LUT4AB/S4END[0]
+ Tile_X2Y2_LUT4AB/S4END[10] Tile_X2Y2_LUT4AB/S4END[11] Tile_X2Y2_LUT4AB/S4END[12]
+ Tile_X2Y2_LUT4AB/S4END[13] Tile_X2Y2_LUT4AB/S4END[14] Tile_X2Y2_LUT4AB/S4END[15]
+ Tile_X2Y2_LUT4AB/S4END[1] Tile_X2Y2_LUT4AB/S4END[2] Tile_X2Y2_LUT4AB/S4END[3] Tile_X2Y2_LUT4AB/S4END[4]
+ Tile_X2Y2_LUT4AB/S4END[5] Tile_X2Y2_LUT4AB/S4END[6] Tile_X2Y2_LUT4AB/S4END[7] Tile_X2Y2_LUT4AB/S4END[8]
+ Tile_X2Y2_LUT4AB/S4END[9] Tile_X2Y0_N_IO4/S4BEG[0] Tile_X2Y0_N_IO4/S4BEG[10] Tile_X2Y0_N_IO4/S4BEG[11]
+ Tile_X2Y0_N_IO4/S4BEG[12] Tile_X2Y0_N_IO4/S4BEG[13] Tile_X2Y0_N_IO4/S4BEG[14] Tile_X2Y0_N_IO4/S4BEG[15]
+ Tile_X2Y0_N_IO4/S4BEG[1] Tile_X2Y0_N_IO4/S4BEG[2] Tile_X2Y0_N_IO4/S4BEG[3] Tile_X2Y0_N_IO4/S4BEG[4]
+ Tile_X2Y0_N_IO4/S4BEG[5] Tile_X2Y0_N_IO4/S4BEG[6] Tile_X2Y0_N_IO4/S4BEG[7] Tile_X2Y0_N_IO4/S4BEG[8]
+ Tile_X2Y0_N_IO4/S4BEG[9] Tile_X2Y2_LUT4AB/SS4END[0] Tile_X2Y2_LUT4AB/SS4END[10]
+ Tile_X2Y2_LUT4AB/SS4END[11] Tile_X2Y2_LUT4AB/SS4END[12] Tile_X2Y2_LUT4AB/SS4END[13]
+ Tile_X2Y2_LUT4AB/SS4END[14] Tile_X2Y2_LUT4AB/SS4END[15] Tile_X2Y2_LUT4AB/SS4END[1]
+ Tile_X2Y2_LUT4AB/SS4END[2] Tile_X2Y2_LUT4AB/SS4END[3] Tile_X2Y2_LUT4AB/SS4END[4]
+ Tile_X2Y2_LUT4AB/SS4END[5] Tile_X2Y2_LUT4AB/SS4END[6] Tile_X2Y2_LUT4AB/SS4END[7]
+ Tile_X2Y2_LUT4AB/SS4END[8] Tile_X2Y2_LUT4AB/SS4END[9] Tile_X2Y0_N_IO4/SS4BEG[0]
+ Tile_X2Y0_N_IO4/SS4BEG[10] Tile_X2Y0_N_IO4/SS4BEG[11] Tile_X2Y0_N_IO4/SS4BEG[12]
+ Tile_X2Y0_N_IO4/SS4BEG[13] Tile_X2Y0_N_IO4/SS4BEG[14] Tile_X2Y0_N_IO4/SS4BEG[15]
+ Tile_X2Y0_N_IO4/SS4BEG[1] Tile_X2Y0_N_IO4/SS4BEG[2] Tile_X2Y0_N_IO4/SS4BEG[3] Tile_X2Y0_N_IO4/SS4BEG[4]
+ Tile_X2Y0_N_IO4/SS4BEG[5] Tile_X2Y0_N_IO4/SS4BEG[6] Tile_X2Y0_N_IO4/SS4BEG[7] Tile_X2Y0_N_IO4/SS4BEG[8]
+ Tile_X2Y0_N_IO4/SS4BEG[9] Tile_X2Y1_LUT4AB/UserCLK Tile_X2Y0_N_IO4/UserCLK VGND
+ VPWR Tile_X2Y1_LUT4AB/W1BEG[0] Tile_X2Y1_LUT4AB/W1BEG[1] Tile_X2Y1_LUT4AB/W1BEG[2]
+ Tile_X2Y1_LUT4AB/W1BEG[3] Tile_X3Y1_LUT4AB/W1BEG[0] Tile_X3Y1_LUT4AB/W1BEG[1] Tile_X3Y1_LUT4AB/W1BEG[2]
+ Tile_X3Y1_LUT4AB/W1BEG[3] Tile_X2Y1_LUT4AB/W2BEG[0] Tile_X2Y1_LUT4AB/W2BEG[1] Tile_X2Y1_LUT4AB/W2BEG[2]
+ Tile_X2Y1_LUT4AB/W2BEG[3] Tile_X2Y1_LUT4AB/W2BEG[4] Tile_X2Y1_LUT4AB/W2BEG[5] Tile_X2Y1_LUT4AB/W2BEG[6]
+ Tile_X2Y1_LUT4AB/W2BEG[7] Tile_X1Y1_LUT4AB/W2END[0] Tile_X1Y1_LUT4AB/W2END[1] Tile_X1Y1_LUT4AB/W2END[2]
+ Tile_X1Y1_LUT4AB/W2END[3] Tile_X1Y1_LUT4AB/W2END[4] Tile_X1Y1_LUT4AB/W2END[5] Tile_X1Y1_LUT4AB/W2END[6]
+ Tile_X1Y1_LUT4AB/W2END[7] Tile_X2Y1_LUT4AB/W2END[0] Tile_X2Y1_LUT4AB/W2END[1] Tile_X2Y1_LUT4AB/W2END[2]
+ Tile_X2Y1_LUT4AB/W2END[3] Tile_X2Y1_LUT4AB/W2END[4] Tile_X2Y1_LUT4AB/W2END[5] Tile_X2Y1_LUT4AB/W2END[6]
+ Tile_X2Y1_LUT4AB/W2END[7] Tile_X3Y1_LUT4AB/W2BEG[0] Tile_X3Y1_LUT4AB/W2BEG[1] Tile_X3Y1_LUT4AB/W2BEG[2]
+ Tile_X3Y1_LUT4AB/W2BEG[3] Tile_X3Y1_LUT4AB/W2BEG[4] Tile_X3Y1_LUT4AB/W2BEG[5] Tile_X3Y1_LUT4AB/W2BEG[6]
+ Tile_X3Y1_LUT4AB/W2BEG[7] Tile_X2Y1_LUT4AB/W6BEG[0] Tile_X2Y1_LUT4AB/W6BEG[10] Tile_X2Y1_LUT4AB/W6BEG[11]
+ Tile_X2Y1_LUT4AB/W6BEG[1] Tile_X2Y1_LUT4AB/W6BEG[2] Tile_X2Y1_LUT4AB/W6BEG[3] Tile_X2Y1_LUT4AB/W6BEG[4]
+ Tile_X2Y1_LUT4AB/W6BEG[5] Tile_X2Y1_LUT4AB/W6BEG[6] Tile_X2Y1_LUT4AB/W6BEG[7] Tile_X2Y1_LUT4AB/W6BEG[8]
+ Tile_X2Y1_LUT4AB/W6BEG[9] Tile_X3Y1_LUT4AB/W6BEG[0] Tile_X3Y1_LUT4AB/W6BEG[10] Tile_X3Y1_LUT4AB/W6BEG[11]
+ Tile_X3Y1_LUT4AB/W6BEG[1] Tile_X3Y1_LUT4AB/W6BEG[2] Tile_X3Y1_LUT4AB/W6BEG[3] Tile_X3Y1_LUT4AB/W6BEG[4]
+ Tile_X3Y1_LUT4AB/W6BEG[5] Tile_X3Y1_LUT4AB/W6BEG[6] Tile_X3Y1_LUT4AB/W6BEG[7] Tile_X3Y1_LUT4AB/W6BEG[8]
+ Tile_X3Y1_LUT4AB/W6BEG[9] Tile_X2Y1_LUT4AB/WW4BEG[0] Tile_X2Y1_LUT4AB/WW4BEG[10]
+ Tile_X2Y1_LUT4AB/WW4BEG[11] Tile_X2Y1_LUT4AB/WW4BEG[12] Tile_X2Y1_LUT4AB/WW4BEG[13]
+ Tile_X2Y1_LUT4AB/WW4BEG[14] Tile_X2Y1_LUT4AB/WW4BEG[15] Tile_X2Y1_LUT4AB/WW4BEG[1]
+ Tile_X2Y1_LUT4AB/WW4BEG[2] Tile_X2Y1_LUT4AB/WW4BEG[3] Tile_X2Y1_LUT4AB/WW4BEG[4]
+ Tile_X2Y1_LUT4AB/WW4BEG[5] Tile_X2Y1_LUT4AB/WW4BEG[6] Tile_X2Y1_LUT4AB/WW4BEG[7]
+ Tile_X2Y1_LUT4AB/WW4BEG[8] Tile_X2Y1_LUT4AB/WW4BEG[9] Tile_X3Y1_LUT4AB/WW4BEG[0]
+ Tile_X3Y1_LUT4AB/WW4BEG[10] Tile_X3Y1_LUT4AB/WW4BEG[11] Tile_X3Y1_LUT4AB/WW4BEG[12]
+ Tile_X3Y1_LUT4AB/WW4BEG[13] Tile_X3Y1_LUT4AB/WW4BEG[14] Tile_X3Y1_LUT4AB/WW4BEG[15]
+ Tile_X3Y1_LUT4AB/WW4BEG[1] Tile_X3Y1_LUT4AB/WW4BEG[2] Tile_X3Y1_LUT4AB/WW4BEG[3]
+ Tile_X3Y1_LUT4AB/WW4BEG[4] Tile_X3Y1_LUT4AB/WW4BEG[5] Tile_X3Y1_LUT4AB/WW4BEG[6]
+ Tile_X3Y1_LUT4AB/WW4BEG[7] Tile_X3Y1_LUT4AB/WW4BEG[8] Tile_X3Y1_LUT4AB/WW4BEG[9]
+ LUT4AB
XTile_X5Y4_E_TT_IF Tile_X5Y4_CLK_TT_PROJECT Tile_X4Y4_LUT4AB/E1BEG[0] Tile_X4Y4_LUT4AB/E1BEG[1]
+ Tile_X4Y4_LUT4AB/E1BEG[2] Tile_X4Y4_LUT4AB/E1BEG[3] Tile_X5Y4_E_TT_IF/E2END[0] Tile_X5Y4_E_TT_IF/E2END[1]
+ Tile_X5Y4_E_TT_IF/E2END[2] Tile_X5Y4_E_TT_IF/E2END[3] Tile_X5Y4_E_TT_IF/E2END[4]
+ Tile_X5Y4_E_TT_IF/E2END[5] Tile_X5Y4_E_TT_IF/E2END[6] Tile_X5Y4_E_TT_IF/E2END[7]
+ Tile_X4Y4_LUT4AB/E2BEG[0] Tile_X4Y4_LUT4AB/E2BEG[1] Tile_X4Y4_LUT4AB/E2BEG[2] Tile_X4Y4_LUT4AB/E2BEG[3]
+ Tile_X4Y4_LUT4AB/E2BEG[4] Tile_X4Y4_LUT4AB/E2BEG[5] Tile_X4Y4_LUT4AB/E2BEG[6] Tile_X4Y4_LUT4AB/E2BEG[7]
+ Tile_X4Y4_LUT4AB/E6BEG[0] Tile_X4Y4_LUT4AB/E6BEG[10] Tile_X4Y4_LUT4AB/E6BEG[11]
+ Tile_X4Y4_LUT4AB/E6BEG[1] Tile_X4Y4_LUT4AB/E6BEG[2] Tile_X4Y4_LUT4AB/E6BEG[3] Tile_X4Y4_LUT4AB/E6BEG[4]
+ Tile_X4Y4_LUT4AB/E6BEG[5] Tile_X4Y4_LUT4AB/E6BEG[6] Tile_X4Y4_LUT4AB/E6BEG[7] Tile_X4Y4_LUT4AB/E6BEG[8]
+ Tile_X4Y4_LUT4AB/E6BEG[9] Tile_X4Y4_LUT4AB/EE4BEG[0] Tile_X4Y4_LUT4AB/EE4BEG[10]
+ Tile_X4Y4_LUT4AB/EE4BEG[11] Tile_X4Y4_LUT4AB/EE4BEG[12] Tile_X4Y4_LUT4AB/EE4BEG[13]
+ Tile_X4Y4_LUT4AB/EE4BEG[14] Tile_X4Y4_LUT4AB/EE4BEG[15] Tile_X4Y4_LUT4AB/EE4BEG[1]
+ Tile_X4Y4_LUT4AB/EE4BEG[2] Tile_X4Y4_LUT4AB/EE4BEG[3] Tile_X4Y4_LUT4AB/EE4BEG[4]
+ Tile_X4Y4_LUT4AB/EE4BEG[5] Tile_X4Y4_LUT4AB/EE4BEG[6] Tile_X4Y4_LUT4AB/EE4BEG[7]
+ Tile_X4Y4_LUT4AB/EE4BEG[8] Tile_X4Y4_LUT4AB/EE4BEG[9] Tile_X5Y4_ENA_TT_PROJECT Tile_X5Y4_E_TT_IF/FrameData[0]
+ Tile_X5Y4_E_TT_IF/FrameData[10] Tile_X5Y4_E_TT_IF/FrameData[11] Tile_X5Y4_E_TT_IF/FrameData[12]
+ Tile_X5Y4_E_TT_IF/FrameData[13] Tile_X5Y4_E_TT_IF/FrameData[14] Tile_X5Y4_E_TT_IF/FrameData[15]
+ Tile_X5Y4_E_TT_IF/FrameData[16] Tile_X5Y4_E_TT_IF/FrameData[17] Tile_X5Y4_E_TT_IF/FrameData[18]
+ Tile_X5Y4_E_TT_IF/FrameData[19] Tile_X5Y4_E_TT_IF/FrameData[1] Tile_X5Y4_E_TT_IF/FrameData[20]
+ Tile_X5Y4_E_TT_IF/FrameData[21] Tile_X5Y4_E_TT_IF/FrameData[22] Tile_X5Y4_E_TT_IF/FrameData[23]
+ Tile_X5Y4_E_TT_IF/FrameData[24] Tile_X5Y4_E_TT_IF/FrameData[25] Tile_X5Y4_E_TT_IF/FrameData[26]
+ Tile_X5Y4_E_TT_IF/FrameData[27] Tile_X5Y4_E_TT_IF/FrameData[28] Tile_X5Y4_E_TT_IF/FrameData[29]
+ Tile_X5Y4_E_TT_IF/FrameData[2] Tile_X5Y4_E_TT_IF/FrameData[30] Tile_X5Y4_E_TT_IF/FrameData[31]
+ Tile_X5Y4_E_TT_IF/FrameData[3] Tile_X5Y4_E_TT_IF/FrameData[4] Tile_X5Y4_E_TT_IF/FrameData[5]
+ Tile_X5Y4_E_TT_IF/FrameData[6] Tile_X5Y4_E_TT_IF/FrameData[7] Tile_X5Y4_E_TT_IF/FrameData[8]
+ Tile_X5Y4_E_TT_IF/FrameData[9] Tile_X5Y4_E_TT_IF/FrameData_O[0] Tile_X5Y4_E_TT_IF/FrameData_O[10]
+ Tile_X5Y4_E_TT_IF/FrameData_O[11] Tile_X5Y4_E_TT_IF/FrameData_O[12] Tile_X5Y4_E_TT_IF/FrameData_O[13]
+ Tile_X5Y4_E_TT_IF/FrameData_O[14] Tile_X5Y4_E_TT_IF/FrameData_O[15] Tile_X5Y4_E_TT_IF/FrameData_O[16]
+ Tile_X5Y4_E_TT_IF/FrameData_O[17] Tile_X5Y4_E_TT_IF/FrameData_O[18] Tile_X5Y4_E_TT_IF/FrameData_O[19]
+ Tile_X5Y4_E_TT_IF/FrameData_O[1] Tile_X5Y4_E_TT_IF/FrameData_O[20] Tile_X5Y4_E_TT_IF/FrameData_O[21]
+ Tile_X5Y4_E_TT_IF/FrameData_O[22] Tile_X5Y4_E_TT_IF/FrameData_O[23] Tile_X5Y4_E_TT_IF/FrameData_O[24]
+ Tile_X5Y4_E_TT_IF/FrameData_O[25] Tile_X5Y4_E_TT_IF/FrameData_O[26] Tile_X5Y4_E_TT_IF/FrameData_O[27]
+ Tile_X5Y4_E_TT_IF/FrameData_O[28] Tile_X5Y4_E_TT_IF/FrameData_O[29] Tile_X5Y4_E_TT_IF/FrameData_O[2]
+ Tile_X5Y4_E_TT_IF/FrameData_O[30] Tile_X5Y4_E_TT_IF/FrameData_O[31] Tile_X5Y4_E_TT_IF/FrameData_O[3]
+ Tile_X5Y4_E_TT_IF/FrameData_O[4] Tile_X5Y4_E_TT_IF/FrameData_O[5] Tile_X5Y4_E_TT_IF/FrameData_O[6]
+ Tile_X5Y4_E_TT_IF/FrameData_O[7] Tile_X5Y4_E_TT_IF/FrameData_O[8] Tile_X5Y4_E_TT_IF/FrameData_O[9]
+ Tile_X5Y4_E_TT_IF/FrameStrobe[0] Tile_X5Y4_E_TT_IF/FrameStrobe[10] Tile_X5Y4_E_TT_IF/FrameStrobe[11]
+ Tile_X5Y4_E_TT_IF/FrameStrobe[12] Tile_X5Y4_E_TT_IF/FrameStrobe[13] Tile_X5Y4_E_TT_IF/FrameStrobe[14]
+ Tile_X5Y4_E_TT_IF/FrameStrobe[15] Tile_X5Y4_E_TT_IF/FrameStrobe[16] Tile_X5Y4_E_TT_IF/FrameStrobe[17]
+ Tile_X5Y4_E_TT_IF/FrameStrobe[18] Tile_X5Y4_E_TT_IF/FrameStrobe[19] Tile_X5Y4_E_TT_IF/FrameStrobe[1]
+ Tile_X5Y4_E_TT_IF/FrameStrobe[2] Tile_X5Y4_E_TT_IF/FrameStrobe[3] Tile_X5Y4_E_TT_IF/FrameStrobe[4]
+ Tile_X5Y4_E_TT_IF/FrameStrobe[5] Tile_X5Y4_E_TT_IF/FrameStrobe[6] Tile_X5Y4_E_TT_IF/FrameStrobe[7]
+ Tile_X5Y4_E_TT_IF/FrameStrobe[8] Tile_X5Y4_E_TT_IF/FrameStrobe[9] Tile_X5Y3_E_TT_IF/FrameStrobe[0]
+ Tile_X5Y3_E_TT_IF/FrameStrobe[10] Tile_X5Y3_E_TT_IF/FrameStrobe[11] Tile_X5Y3_E_TT_IF/FrameStrobe[12]
+ Tile_X5Y3_E_TT_IF/FrameStrobe[13] Tile_X5Y3_E_TT_IF/FrameStrobe[14] Tile_X5Y3_E_TT_IF/FrameStrobe[15]
+ Tile_X5Y3_E_TT_IF/FrameStrobe[16] Tile_X5Y3_E_TT_IF/FrameStrobe[17] Tile_X5Y3_E_TT_IF/FrameStrobe[18]
+ Tile_X5Y3_E_TT_IF/FrameStrobe[19] Tile_X5Y3_E_TT_IF/FrameStrobe[1] Tile_X5Y3_E_TT_IF/FrameStrobe[2]
+ Tile_X5Y3_E_TT_IF/FrameStrobe[3] Tile_X5Y3_E_TT_IF/FrameStrobe[4] Tile_X5Y3_E_TT_IF/FrameStrobe[5]
+ Tile_X5Y3_E_TT_IF/FrameStrobe[6] Tile_X5Y3_E_TT_IF/FrameStrobe[7] Tile_X5Y3_E_TT_IF/FrameStrobe[8]
+ Tile_X5Y3_E_TT_IF/FrameStrobe[9] Tile_X5Y4_E_TT_IF/N1BEG[0] Tile_X5Y4_E_TT_IF/N1BEG[1]
+ Tile_X5Y4_E_TT_IF/N1BEG[2] Tile_X5Y4_E_TT_IF/N1BEG[3] Tile_X5Y5_E_TT_IF/N1BEG[0]
+ Tile_X5Y5_E_TT_IF/N1BEG[1] Tile_X5Y5_E_TT_IF/N1BEG[2] Tile_X5Y5_E_TT_IF/N1BEG[3]
+ Tile_X5Y4_E_TT_IF/N2BEG[0] Tile_X5Y4_E_TT_IF/N2BEG[1] Tile_X5Y4_E_TT_IF/N2BEG[2]
+ Tile_X5Y4_E_TT_IF/N2BEG[3] Tile_X5Y4_E_TT_IF/N2BEG[4] Tile_X5Y4_E_TT_IF/N2BEG[5]
+ Tile_X5Y4_E_TT_IF/N2BEG[6] Tile_X5Y4_E_TT_IF/N2BEG[7] Tile_X5Y3_E_TT_IF/N2END[0]
+ Tile_X5Y3_E_TT_IF/N2END[1] Tile_X5Y3_E_TT_IF/N2END[2] Tile_X5Y3_E_TT_IF/N2END[3]
+ Tile_X5Y3_E_TT_IF/N2END[4] Tile_X5Y3_E_TT_IF/N2END[5] Tile_X5Y3_E_TT_IF/N2END[6]
+ Tile_X5Y3_E_TT_IF/N2END[7] Tile_X5Y4_E_TT_IF/N2END[0] Tile_X5Y4_E_TT_IF/N2END[1]
+ Tile_X5Y4_E_TT_IF/N2END[2] Tile_X5Y4_E_TT_IF/N2END[3] Tile_X5Y4_E_TT_IF/N2END[4]
+ Tile_X5Y4_E_TT_IF/N2END[5] Tile_X5Y4_E_TT_IF/N2END[6] Tile_X5Y4_E_TT_IF/N2END[7]
+ Tile_X5Y5_E_TT_IF/N2BEG[0] Tile_X5Y5_E_TT_IF/N2BEG[1] Tile_X5Y5_E_TT_IF/N2BEG[2]
+ Tile_X5Y5_E_TT_IF/N2BEG[3] Tile_X5Y5_E_TT_IF/N2BEG[4] Tile_X5Y5_E_TT_IF/N2BEG[5]
+ Tile_X5Y5_E_TT_IF/N2BEG[6] Tile_X5Y5_E_TT_IF/N2BEG[7] Tile_X5Y4_E_TT_IF/N4BEG[0]
+ Tile_X5Y4_E_TT_IF/N4BEG[10] Tile_X5Y4_E_TT_IF/N4BEG[11] Tile_X5Y4_E_TT_IF/N4BEG[12]
+ Tile_X5Y4_E_TT_IF/N4BEG[13] Tile_X5Y4_E_TT_IF/N4BEG[14] Tile_X5Y4_E_TT_IF/N4BEG[15]
+ Tile_X5Y4_E_TT_IF/N4BEG[1] Tile_X5Y4_E_TT_IF/N4BEG[2] Tile_X5Y4_E_TT_IF/N4BEG[3]
+ Tile_X5Y4_E_TT_IF/N4BEG[4] Tile_X5Y4_E_TT_IF/N4BEG[5] Tile_X5Y4_E_TT_IF/N4BEG[6]
+ Tile_X5Y4_E_TT_IF/N4BEG[7] Tile_X5Y4_E_TT_IF/N4BEG[8] Tile_X5Y4_E_TT_IF/N4BEG[9]
+ Tile_X5Y5_E_TT_IF/N4BEG[0] Tile_X5Y5_E_TT_IF/N4BEG[10] Tile_X5Y5_E_TT_IF/N4BEG[11]
+ Tile_X5Y5_E_TT_IF/N4BEG[12] Tile_X5Y5_E_TT_IF/N4BEG[13] Tile_X5Y5_E_TT_IF/N4BEG[14]
+ Tile_X5Y5_E_TT_IF/N4BEG[15] Tile_X5Y5_E_TT_IF/N4BEG[1] Tile_X5Y5_E_TT_IF/N4BEG[2]
+ Tile_X5Y5_E_TT_IF/N4BEG[3] Tile_X5Y5_E_TT_IF/N4BEG[4] Tile_X5Y5_E_TT_IF/N4BEG[5]
+ Tile_X5Y5_E_TT_IF/N4BEG[6] Tile_X5Y5_E_TT_IF/N4BEG[7] Tile_X5Y5_E_TT_IF/N4BEG[8]
+ Tile_X5Y5_E_TT_IF/N4BEG[9] Tile_X5Y4_RST_N_TT_PROJECT Tile_X5Y5_E_TT_IF/S1END[0]
+ Tile_X5Y5_E_TT_IF/S1END[1] Tile_X5Y5_E_TT_IF/S1END[2] Tile_X5Y5_E_TT_IF/S1END[3]
+ Tile_X5Y4_E_TT_IF/S1END[0] Tile_X5Y4_E_TT_IF/S1END[1] Tile_X5Y4_E_TT_IF/S1END[2]
+ Tile_X5Y4_E_TT_IF/S1END[3] Tile_X5Y5_E_TT_IF/S2MID[0] Tile_X5Y5_E_TT_IF/S2MID[1]
+ Tile_X5Y5_E_TT_IF/S2MID[2] Tile_X5Y5_E_TT_IF/S2MID[3] Tile_X5Y5_E_TT_IF/S2MID[4]
+ Tile_X5Y5_E_TT_IF/S2MID[5] Tile_X5Y5_E_TT_IF/S2MID[6] Tile_X5Y5_E_TT_IF/S2MID[7]
+ Tile_X5Y5_E_TT_IF/S2END[0] Tile_X5Y5_E_TT_IF/S2END[1] Tile_X5Y5_E_TT_IF/S2END[2]
+ Tile_X5Y5_E_TT_IF/S2END[3] Tile_X5Y5_E_TT_IF/S2END[4] Tile_X5Y5_E_TT_IF/S2END[5]
+ Tile_X5Y5_E_TT_IF/S2END[6] Tile_X5Y5_E_TT_IF/S2END[7] Tile_X5Y4_E_TT_IF/S2END[0]
+ Tile_X5Y4_E_TT_IF/S2END[1] Tile_X5Y4_E_TT_IF/S2END[2] Tile_X5Y4_E_TT_IF/S2END[3]
+ Tile_X5Y4_E_TT_IF/S2END[4] Tile_X5Y4_E_TT_IF/S2END[5] Tile_X5Y4_E_TT_IF/S2END[6]
+ Tile_X5Y4_E_TT_IF/S2END[7] Tile_X5Y4_E_TT_IF/S2MID[0] Tile_X5Y4_E_TT_IF/S2MID[1]
+ Tile_X5Y4_E_TT_IF/S2MID[2] Tile_X5Y4_E_TT_IF/S2MID[3] Tile_X5Y4_E_TT_IF/S2MID[4]
+ Tile_X5Y4_E_TT_IF/S2MID[5] Tile_X5Y4_E_TT_IF/S2MID[6] Tile_X5Y4_E_TT_IF/S2MID[7]
+ Tile_X5Y5_E_TT_IF/S4END[0] Tile_X5Y5_E_TT_IF/S4END[10] Tile_X5Y5_E_TT_IF/S4END[11]
+ Tile_X5Y5_E_TT_IF/S4END[12] Tile_X5Y5_E_TT_IF/S4END[13] Tile_X5Y5_E_TT_IF/S4END[14]
+ Tile_X5Y5_E_TT_IF/S4END[15] Tile_X5Y5_E_TT_IF/S4END[1] Tile_X5Y5_E_TT_IF/S4END[2]
+ Tile_X5Y5_E_TT_IF/S4END[3] Tile_X5Y5_E_TT_IF/S4END[4] Tile_X5Y5_E_TT_IF/S4END[5]
+ Tile_X5Y5_E_TT_IF/S4END[6] Tile_X5Y5_E_TT_IF/S4END[7] Tile_X5Y5_E_TT_IF/S4END[8]
+ Tile_X5Y5_E_TT_IF/S4END[9] Tile_X5Y4_E_TT_IF/S4END[0] Tile_X5Y4_E_TT_IF/S4END[10]
+ Tile_X5Y4_E_TT_IF/S4END[11] Tile_X5Y4_E_TT_IF/S4END[12] Tile_X5Y4_E_TT_IF/S4END[13]
+ Tile_X5Y4_E_TT_IF/S4END[14] Tile_X5Y4_E_TT_IF/S4END[15] Tile_X5Y4_E_TT_IF/S4END[1]
+ Tile_X5Y4_E_TT_IF/S4END[2] Tile_X5Y4_E_TT_IF/S4END[3] Tile_X5Y4_E_TT_IF/S4END[4]
+ Tile_X5Y4_E_TT_IF/S4END[5] Tile_X5Y4_E_TT_IF/S4END[6] Tile_X5Y4_E_TT_IF/S4END[7]
+ Tile_X5Y4_E_TT_IF/S4END[8] Tile_X5Y4_E_TT_IF/S4END[9] Tile_X5Y4_UIO_IN_TT_PROJECT0
+ Tile_X5Y4_UIO_IN_TT_PROJECT1 Tile_X5Y4_UIO_IN_TT_PROJECT2 Tile_X5Y4_UIO_IN_TT_PROJECT3
+ Tile_X5Y4_UIO_IN_TT_PROJECT4 Tile_X5Y4_UIO_IN_TT_PROJECT5 Tile_X5Y4_UIO_IN_TT_PROJECT6
+ Tile_X5Y4_UIO_IN_TT_PROJECT7 Tile_X5Y4_UIO_OE_TT_PROJECT0 Tile_X5Y4_UIO_OE_TT_PROJECT1
+ Tile_X5Y4_UIO_OE_TT_PROJECT2 Tile_X5Y4_UIO_OE_TT_PROJECT3 Tile_X5Y4_UIO_OE_TT_PROJECT4
+ Tile_X5Y4_UIO_OE_TT_PROJECT5 Tile_X5Y4_UIO_OE_TT_PROJECT6 Tile_X5Y4_UIO_OE_TT_PROJECT7
+ Tile_X5Y4_UIO_OUT_TT_PROJECT0 Tile_X5Y4_UIO_OUT_TT_PROJECT1 Tile_X5Y4_UIO_OUT_TT_PROJECT2
+ Tile_X5Y4_UIO_OUT_TT_PROJECT3 Tile_X5Y4_UIO_OUT_TT_PROJECT4 Tile_X5Y4_UIO_OUT_TT_PROJECT5
+ Tile_X5Y4_UIO_OUT_TT_PROJECT6 Tile_X5Y4_UIO_OUT_TT_PROJECT7 Tile_X5Y4_UI_IN_TT_PROJECT0
+ Tile_X5Y4_UI_IN_TT_PROJECT1 Tile_X5Y4_UI_IN_TT_PROJECT2 Tile_X5Y4_UI_IN_TT_PROJECT3
+ Tile_X5Y4_UI_IN_TT_PROJECT4 Tile_X5Y4_UI_IN_TT_PROJECT5 Tile_X5Y4_UI_IN_TT_PROJECT6
+ Tile_X5Y4_UI_IN_TT_PROJECT7 Tile_X5Y4_UO_OUT_TT_PROJECT0 Tile_X5Y4_UO_OUT_TT_PROJECT1
+ Tile_X5Y4_UO_OUT_TT_PROJECT2 Tile_X5Y4_UO_OUT_TT_PROJECT3 Tile_X5Y4_UO_OUT_TT_PROJECT4
+ Tile_X5Y4_UO_OUT_TT_PROJECT5 Tile_X5Y4_UO_OUT_TT_PROJECT6 Tile_X5Y4_UO_OUT_TT_PROJECT7
+ Tile_X5Y4_E_TT_IF/UserCLK Tile_X5Y3_E_TT_IF/UserCLK VGND VPWR Tile_X4Y4_LUT4AB/W1END[0]
+ Tile_X4Y4_LUT4AB/W1END[1] Tile_X4Y4_LUT4AB/W1END[2] Tile_X4Y4_LUT4AB/W1END[3] Tile_X4Y4_LUT4AB/W2MID[0]
+ Tile_X4Y4_LUT4AB/W2MID[1] Tile_X4Y4_LUT4AB/W2MID[2] Tile_X4Y4_LUT4AB/W2MID[3] Tile_X4Y4_LUT4AB/W2MID[4]
+ Tile_X4Y4_LUT4AB/W2MID[5] Tile_X4Y4_LUT4AB/W2MID[6] Tile_X4Y4_LUT4AB/W2MID[7] Tile_X4Y4_LUT4AB/W2END[0]
+ Tile_X4Y4_LUT4AB/W2END[1] Tile_X4Y4_LUT4AB/W2END[2] Tile_X4Y4_LUT4AB/W2END[3] Tile_X4Y4_LUT4AB/W2END[4]
+ Tile_X4Y4_LUT4AB/W2END[5] Tile_X4Y4_LUT4AB/W2END[6] Tile_X4Y4_LUT4AB/W2END[7] Tile_X4Y4_LUT4AB/W6END[0]
+ Tile_X4Y4_LUT4AB/W6END[10] Tile_X4Y4_LUT4AB/W6END[11] Tile_X4Y4_LUT4AB/W6END[1]
+ Tile_X4Y4_LUT4AB/W6END[2] Tile_X4Y4_LUT4AB/W6END[3] Tile_X4Y4_LUT4AB/W6END[4] Tile_X4Y4_LUT4AB/W6END[5]
+ Tile_X4Y4_LUT4AB/W6END[6] Tile_X4Y4_LUT4AB/W6END[7] Tile_X4Y4_LUT4AB/W6END[8] Tile_X4Y4_LUT4AB/W6END[9]
+ Tile_X4Y4_LUT4AB/WW4END[0] Tile_X4Y4_LUT4AB/WW4END[10] Tile_X4Y4_LUT4AB/WW4END[11]
+ Tile_X4Y4_LUT4AB/WW4END[12] Tile_X4Y4_LUT4AB/WW4END[13] Tile_X4Y4_LUT4AB/WW4END[14]
+ Tile_X4Y4_LUT4AB/WW4END[15] Tile_X4Y4_LUT4AB/WW4END[1] Tile_X4Y4_LUT4AB/WW4END[2]
+ Tile_X4Y4_LUT4AB/WW4END[3] Tile_X4Y4_LUT4AB/WW4END[4] Tile_X4Y4_LUT4AB/WW4END[5]
+ Tile_X4Y4_LUT4AB/WW4END[6] Tile_X4Y4_LUT4AB/WW4END[7] Tile_X4Y4_LUT4AB/WW4END[8]
+ Tile_X4Y4_LUT4AB/WW4END[9] E_TT_IF
XTile_X1Y5_LUT4AB Tile_X1Y6_LUT4AB/Co Tile_X1Y5_LUT4AB/Co Tile_X2Y5_LUT4AB/E1END[0]
+ Tile_X2Y5_LUT4AB/E1END[1] Tile_X2Y5_LUT4AB/E1END[2] Tile_X2Y5_LUT4AB/E1END[3] Tile_X1Y5_LUT4AB/E1END[0]
+ Tile_X1Y5_LUT4AB/E1END[1] Tile_X1Y5_LUT4AB/E1END[2] Tile_X1Y5_LUT4AB/E1END[3] Tile_X2Y5_LUT4AB/E2MID[0]
+ Tile_X2Y5_LUT4AB/E2MID[1] Tile_X2Y5_LUT4AB/E2MID[2] Tile_X2Y5_LUT4AB/E2MID[3] Tile_X2Y5_LUT4AB/E2MID[4]
+ Tile_X2Y5_LUT4AB/E2MID[5] Tile_X2Y5_LUT4AB/E2MID[6] Tile_X2Y5_LUT4AB/E2MID[7] Tile_X2Y5_LUT4AB/E2END[0]
+ Tile_X2Y5_LUT4AB/E2END[1] Tile_X2Y5_LUT4AB/E2END[2] Tile_X2Y5_LUT4AB/E2END[3] Tile_X2Y5_LUT4AB/E2END[4]
+ Tile_X2Y5_LUT4AB/E2END[5] Tile_X2Y5_LUT4AB/E2END[6] Tile_X2Y5_LUT4AB/E2END[7] Tile_X1Y5_LUT4AB/E2END[0]
+ Tile_X1Y5_LUT4AB/E2END[1] Tile_X1Y5_LUT4AB/E2END[2] Tile_X1Y5_LUT4AB/E2END[3] Tile_X1Y5_LUT4AB/E2END[4]
+ Tile_X1Y5_LUT4AB/E2END[5] Tile_X1Y5_LUT4AB/E2END[6] Tile_X1Y5_LUT4AB/E2END[7] Tile_X1Y5_LUT4AB/E2MID[0]
+ Tile_X1Y5_LUT4AB/E2MID[1] Tile_X1Y5_LUT4AB/E2MID[2] Tile_X1Y5_LUT4AB/E2MID[3] Tile_X1Y5_LUT4AB/E2MID[4]
+ Tile_X1Y5_LUT4AB/E2MID[5] Tile_X1Y5_LUT4AB/E2MID[6] Tile_X1Y5_LUT4AB/E2MID[7] Tile_X2Y5_LUT4AB/E6END[0]
+ Tile_X2Y5_LUT4AB/E6END[10] Tile_X2Y5_LUT4AB/E6END[11] Tile_X2Y5_LUT4AB/E6END[1]
+ Tile_X2Y5_LUT4AB/E6END[2] Tile_X2Y5_LUT4AB/E6END[3] Tile_X2Y5_LUT4AB/E6END[4] Tile_X2Y5_LUT4AB/E6END[5]
+ Tile_X2Y5_LUT4AB/E6END[6] Tile_X2Y5_LUT4AB/E6END[7] Tile_X2Y5_LUT4AB/E6END[8] Tile_X2Y5_LUT4AB/E6END[9]
+ Tile_X1Y5_LUT4AB/E6END[0] Tile_X1Y5_LUT4AB/E6END[10] Tile_X1Y5_LUT4AB/E6END[11]
+ Tile_X1Y5_LUT4AB/E6END[1] Tile_X1Y5_LUT4AB/E6END[2] Tile_X1Y5_LUT4AB/E6END[3] Tile_X1Y5_LUT4AB/E6END[4]
+ Tile_X1Y5_LUT4AB/E6END[5] Tile_X1Y5_LUT4AB/E6END[6] Tile_X1Y5_LUT4AB/E6END[7] Tile_X1Y5_LUT4AB/E6END[8]
+ Tile_X1Y5_LUT4AB/E6END[9] Tile_X2Y5_LUT4AB/EE4END[0] Tile_X2Y5_LUT4AB/EE4END[10]
+ Tile_X2Y5_LUT4AB/EE4END[11] Tile_X2Y5_LUT4AB/EE4END[12] Tile_X2Y5_LUT4AB/EE4END[13]
+ Tile_X2Y5_LUT4AB/EE4END[14] Tile_X2Y5_LUT4AB/EE4END[15] Tile_X2Y5_LUT4AB/EE4END[1]
+ Tile_X2Y5_LUT4AB/EE4END[2] Tile_X2Y5_LUT4AB/EE4END[3] Tile_X2Y5_LUT4AB/EE4END[4]
+ Tile_X2Y5_LUT4AB/EE4END[5] Tile_X2Y5_LUT4AB/EE4END[6] Tile_X2Y5_LUT4AB/EE4END[7]
+ Tile_X2Y5_LUT4AB/EE4END[8] Tile_X2Y5_LUT4AB/EE4END[9] Tile_X1Y5_LUT4AB/EE4END[0]
+ Tile_X1Y5_LUT4AB/EE4END[10] Tile_X1Y5_LUT4AB/EE4END[11] Tile_X1Y5_LUT4AB/EE4END[12]
+ Tile_X1Y5_LUT4AB/EE4END[13] Tile_X1Y5_LUT4AB/EE4END[14] Tile_X1Y5_LUT4AB/EE4END[15]
+ Tile_X1Y5_LUT4AB/EE4END[1] Tile_X1Y5_LUT4AB/EE4END[2] Tile_X1Y5_LUT4AB/EE4END[3]
+ Tile_X1Y5_LUT4AB/EE4END[4] Tile_X1Y5_LUT4AB/EE4END[5] Tile_X1Y5_LUT4AB/EE4END[6]
+ Tile_X1Y5_LUT4AB/EE4END[7] Tile_X1Y5_LUT4AB/EE4END[8] Tile_X1Y5_LUT4AB/EE4END[9]
+ Tile_X1Y5_LUT4AB/FrameData[0] Tile_X1Y5_LUT4AB/FrameData[10] Tile_X1Y5_LUT4AB/FrameData[11]
+ Tile_X1Y5_LUT4AB/FrameData[12] Tile_X1Y5_LUT4AB/FrameData[13] Tile_X1Y5_LUT4AB/FrameData[14]
+ Tile_X1Y5_LUT4AB/FrameData[15] Tile_X1Y5_LUT4AB/FrameData[16] Tile_X1Y5_LUT4AB/FrameData[17]
+ Tile_X1Y5_LUT4AB/FrameData[18] Tile_X1Y5_LUT4AB/FrameData[19] Tile_X1Y5_LUT4AB/FrameData[1]
+ Tile_X1Y5_LUT4AB/FrameData[20] Tile_X1Y5_LUT4AB/FrameData[21] Tile_X1Y5_LUT4AB/FrameData[22]
+ Tile_X1Y5_LUT4AB/FrameData[23] Tile_X1Y5_LUT4AB/FrameData[24] Tile_X1Y5_LUT4AB/FrameData[25]
+ Tile_X1Y5_LUT4AB/FrameData[26] Tile_X1Y5_LUT4AB/FrameData[27] Tile_X1Y5_LUT4AB/FrameData[28]
+ Tile_X1Y5_LUT4AB/FrameData[29] Tile_X1Y5_LUT4AB/FrameData[2] Tile_X1Y5_LUT4AB/FrameData[30]
+ Tile_X1Y5_LUT4AB/FrameData[31] Tile_X1Y5_LUT4AB/FrameData[3] Tile_X1Y5_LUT4AB/FrameData[4]
+ Tile_X1Y5_LUT4AB/FrameData[5] Tile_X1Y5_LUT4AB/FrameData[6] Tile_X1Y5_LUT4AB/FrameData[7]
+ Tile_X1Y5_LUT4AB/FrameData[8] Tile_X1Y5_LUT4AB/FrameData[9] Tile_X2Y5_LUT4AB/FrameData[0]
+ Tile_X2Y5_LUT4AB/FrameData[10] Tile_X2Y5_LUT4AB/FrameData[11] Tile_X2Y5_LUT4AB/FrameData[12]
+ Tile_X2Y5_LUT4AB/FrameData[13] Tile_X2Y5_LUT4AB/FrameData[14] Tile_X2Y5_LUT4AB/FrameData[15]
+ Tile_X2Y5_LUT4AB/FrameData[16] Tile_X2Y5_LUT4AB/FrameData[17] Tile_X2Y5_LUT4AB/FrameData[18]
+ Tile_X2Y5_LUT4AB/FrameData[19] Tile_X2Y5_LUT4AB/FrameData[1] Tile_X2Y5_LUT4AB/FrameData[20]
+ Tile_X2Y5_LUT4AB/FrameData[21] Tile_X2Y5_LUT4AB/FrameData[22] Tile_X2Y5_LUT4AB/FrameData[23]
+ Tile_X2Y5_LUT4AB/FrameData[24] Tile_X2Y5_LUT4AB/FrameData[25] Tile_X2Y5_LUT4AB/FrameData[26]
+ Tile_X2Y5_LUT4AB/FrameData[27] Tile_X2Y5_LUT4AB/FrameData[28] Tile_X2Y5_LUT4AB/FrameData[29]
+ Tile_X2Y5_LUT4AB/FrameData[2] Tile_X2Y5_LUT4AB/FrameData[30] Tile_X2Y5_LUT4AB/FrameData[31]
+ Tile_X2Y5_LUT4AB/FrameData[3] Tile_X2Y5_LUT4AB/FrameData[4] Tile_X2Y5_LUT4AB/FrameData[5]
+ Tile_X2Y5_LUT4AB/FrameData[6] Tile_X2Y5_LUT4AB/FrameData[7] Tile_X2Y5_LUT4AB/FrameData[8]
+ Tile_X2Y5_LUT4AB/FrameData[9] Tile_X1Y5_LUT4AB/FrameStrobe[0] Tile_X1Y5_LUT4AB/FrameStrobe[10]
+ Tile_X1Y5_LUT4AB/FrameStrobe[11] Tile_X1Y5_LUT4AB/FrameStrobe[12] Tile_X1Y5_LUT4AB/FrameStrobe[13]
+ Tile_X1Y5_LUT4AB/FrameStrobe[14] Tile_X1Y5_LUT4AB/FrameStrobe[15] Tile_X1Y5_LUT4AB/FrameStrobe[16]
+ Tile_X1Y5_LUT4AB/FrameStrobe[17] Tile_X1Y5_LUT4AB/FrameStrobe[18] Tile_X1Y5_LUT4AB/FrameStrobe[19]
+ Tile_X1Y5_LUT4AB/FrameStrobe[1] Tile_X1Y5_LUT4AB/FrameStrobe[2] Tile_X1Y5_LUT4AB/FrameStrobe[3]
+ Tile_X1Y5_LUT4AB/FrameStrobe[4] Tile_X1Y5_LUT4AB/FrameStrobe[5] Tile_X1Y5_LUT4AB/FrameStrobe[6]
+ Tile_X1Y5_LUT4AB/FrameStrobe[7] Tile_X1Y5_LUT4AB/FrameStrobe[8] Tile_X1Y5_LUT4AB/FrameStrobe[9]
+ Tile_X1Y4_LUT4AB/FrameStrobe[0] Tile_X1Y4_LUT4AB/FrameStrobe[10] Tile_X1Y4_LUT4AB/FrameStrobe[11]
+ Tile_X1Y4_LUT4AB/FrameStrobe[12] Tile_X1Y4_LUT4AB/FrameStrobe[13] Tile_X1Y4_LUT4AB/FrameStrobe[14]
+ Tile_X1Y4_LUT4AB/FrameStrobe[15] Tile_X1Y4_LUT4AB/FrameStrobe[16] Tile_X1Y4_LUT4AB/FrameStrobe[17]
+ Tile_X1Y4_LUT4AB/FrameStrobe[18] Tile_X1Y4_LUT4AB/FrameStrobe[19] Tile_X1Y4_LUT4AB/FrameStrobe[1]
+ Tile_X1Y4_LUT4AB/FrameStrobe[2] Tile_X1Y4_LUT4AB/FrameStrobe[3] Tile_X1Y4_LUT4AB/FrameStrobe[4]
+ Tile_X1Y4_LUT4AB/FrameStrobe[5] Tile_X1Y4_LUT4AB/FrameStrobe[6] Tile_X1Y4_LUT4AB/FrameStrobe[7]
+ Tile_X1Y4_LUT4AB/FrameStrobe[8] Tile_X1Y4_LUT4AB/FrameStrobe[9] Tile_X1Y5_LUT4AB/N1BEG[0]
+ Tile_X1Y5_LUT4AB/N1BEG[1] Tile_X1Y5_LUT4AB/N1BEG[2] Tile_X1Y5_LUT4AB/N1BEG[3] Tile_X1Y6_LUT4AB/N1BEG[0]
+ Tile_X1Y6_LUT4AB/N1BEG[1] Tile_X1Y6_LUT4AB/N1BEG[2] Tile_X1Y6_LUT4AB/N1BEG[3] Tile_X1Y5_LUT4AB/N2BEG[0]
+ Tile_X1Y5_LUT4AB/N2BEG[1] Tile_X1Y5_LUT4AB/N2BEG[2] Tile_X1Y5_LUT4AB/N2BEG[3] Tile_X1Y5_LUT4AB/N2BEG[4]
+ Tile_X1Y5_LUT4AB/N2BEG[5] Tile_X1Y5_LUT4AB/N2BEG[6] Tile_X1Y5_LUT4AB/N2BEG[7] Tile_X1Y4_LUT4AB/N2END[0]
+ Tile_X1Y4_LUT4AB/N2END[1] Tile_X1Y4_LUT4AB/N2END[2] Tile_X1Y4_LUT4AB/N2END[3] Tile_X1Y4_LUT4AB/N2END[4]
+ Tile_X1Y4_LUT4AB/N2END[5] Tile_X1Y4_LUT4AB/N2END[6] Tile_X1Y4_LUT4AB/N2END[7] Tile_X1Y5_LUT4AB/N2END[0]
+ Tile_X1Y5_LUT4AB/N2END[1] Tile_X1Y5_LUT4AB/N2END[2] Tile_X1Y5_LUT4AB/N2END[3] Tile_X1Y5_LUT4AB/N2END[4]
+ Tile_X1Y5_LUT4AB/N2END[5] Tile_X1Y5_LUT4AB/N2END[6] Tile_X1Y5_LUT4AB/N2END[7] Tile_X1Y6_LUT4AB/N2BEG[0]
+ Tile_X1Y6_LUT4AB/N2BEG[1] Tile_X1Y6_LUT4AB/N2BEG[2] Tile_X1Y6_LUT4AB/N2BEG[3] Tile_X1Y6_LUT4AB/N2BEG[4]
+ Tile_X1Y6_LUT4AB/N2BEG[5] Tile_X1Y6_LUT4AB/N2BEG[6] Tile_X1Y6_LUT4AB/N2BEG[7] Tile_X1Y5_LUT4AB/N4BEG[0]
+ Tile_X1Y5_LUT4AB/N4BEG[10] Tile_X1Y5_LUT4AB/N4BEG[11] Tile_X1Y5_LUT4AB/N4BEG[12]
+ Tile_X1Y5_LUT4AB/N4BEG[13] Tile_X1Y5_LUT4AB/N4BEG[14] Tile_X1Y5_LUT4AB/N4BEG[15]
+ Tile_X1Y5_LUT4AB/N4BEG[1] Tile_X1Y5_LUT4AB/N4BEG[2] Tile_X1Y5_LUT4AB/N4BEG[3] Tile_X1Y5_LUT4AB/N4BEG[4]
+ Tile_X1Y5_LUT4AB/N4BEG[5] Tile_X1Y5_LUT4AB/N4BEG[6] Tile_X1Y5_LUT4AB/N4BEG[7] Tile_X1Y5_LUT4AB/N4BEG[8]
+ Tile_X1Y5_LUT4AB/N4BEG[9] Tile_X1Y6_LUT4AB/N4BEG[0] Tile_X1Y6_LUT4AB/N4BEG[10] Tile_X1Y6_LUT4AB/N4BEG[11]
+ Tile_X1Y6_LUT4AB/N4BEG[12] Tile_X1Y6_LUT4AB/N4BEG[13] Tile_X1Y6_LUT4AB/N4BEG[14]
+ Tile_X1Y6_LUT4AB/N4BEG[15] Tile_X1Y6_LUT4AB/N4BEG[1] Tile_X1Y6_LUT4AB/N4BEG[2] Tile_X1Y6_LUT4AB/N4BEG[3]
+ Tile_X1Y6_LUT4AB/N4BEG[4] Tile_X1Y6_LUT4AB/N4BEG[5] Tile_X1Y6_LUT4AB/N4BEG[6] Tile_X1Y6_LUT4AB/N4BEG[7]
+ Tile_X1Y6_LUT4AB/N4BEG[8] Tile_X1Y6_LUT4AB/N4BEG[9] Tile_X1Y5_LUT4AB/NN4BEG[0] Tile_X1Y5_LUT4AB/NN4BEG[10]
+ Tile_X1Y5_LUT4AB/NN4BEG[11] Tile_X1Y5_LUT4AB/NN4BEG[12] Tile_X1Y5_LUT4AB/NN4BEG[13]
+ Tile_X1Y5_LUT4AB/NN4BEG[14] Tile_X1Y5_LUT4AB/NN4BEG[15] Tile_X1Y5_LUT4AB/NN4BEG[1]
+ Tile_X1Y5_LUT4AB/NN4BEG[2] Tile_X1Y5_LUT4AB/NN4BEG[3] Tile_X1Y5_LUT4AB/NN4BEG[4]
+ Tile_X1Y5_LUT4AB/NN4BEG[5] Tile_X1Y5_LUT4AB/NN4BEG[6] Tile_X1Y5_LUT4AB/NN4BEG[7]
+ Tile_X1Y5_LUT4AB/NN4BEG[8] Tile_X1Y5_LUT4AB/NN4BEG[9] Tile_X1Y6_LUT4AB/NN4BEG[0]
+ Tile_X1Y6_LUT4AB/NN4BEG[10] Tile_X1Y6_LUT4AB/NN4BEG[11] Tile_X1Y6_LUT4AB/NN4BEG[12]
+ Tile_X1Y6_LUT4AB/NN4BEG[13] Tile_X1Y6_LUT4AB/NN4BEG[14] Tile_X1Y6_LUT4AB/NN4BEG[15]
+ Tile_X1Y6_LUT4AB/NN4BEG[1] Tile_X1Y6_LUT4AB/NN4BEG[2] Tile_X1Y6_LUT4AB/NN4BEG[3]
+ Tile_X1Y6_LUT4AB/NN4BEG[4] Tile_X1Y6_LUT4AB/NN4BEG[5] Tile_X1Y6_LUT4AB/NN4BEG[6]
+ Tile_X1Y6_LUT4AB/NN4BEG[7] Tile_X1Y6_LUT4AB/NN4BEG[8] Tile_X1Y6_LUT4AB/NN4BEG[9]
+ Tile_X1Y6_LUT4AB/S1END[0] Tile_X1Y6_LUT4AB/S1END[1] Tile_X1Y6_LUT4AB/S1END[2] Tile_X1Y6_LUT4AB/S1END[3]
+ Tile_X1Y5_LUT4AB/S1END[0] Tile_X1Y5_LUT4AB/S1END[1] Tile_X1Y5_LUT4AB/S1END[2] Tile_X1Y5_LUT4AB/S1END[3]
+ Tile_X1Y6_LUT4AB/S2MID[0] Tile_X1Y6_LUT4AB/S2MID[1] Tile_X1Y6_LUT4AB/S2MID[2] Tile_X1Y6_LUT4AB/S2MID[3]
+ Tile_X1Y6_LUT4AB/S2MID[4] Tile_X1Y6_LUT4AB/S2MID[5] Tile_X1Y6_LUT4AB/S2MID[6] Tile_X1Y6_LUT4AB/S2MID[7]
+ Tile_X1Y6_LUT4AB/S2END[0] Tile_X1Y6_LUT4AB/S2END[1] Tile_X1Y6_LUT4AB/S2END[2] Tile_X1Y6_LUT4AB/S2END[3]
+ Tile_X1Y6_LUT4AB/S2END[4] Tile_X1Y6_LUT4AB/S2END[5] Tile_X1Y6_LUT4AB/S2END[6] Tile_X1Y6_LUT4AB/S2END[7]
+ Tile_X1Y5_LUT4AB/S2END[0] Tile_X1Y5_LUT4AB/S2END[1] Tile_X1Y5_LUT4AB/S2END[2] Tile_X1Y5_LUT4AB/S2END[3]
+ Tile_X1Y5_LUT4AB/S2END[4] Tile_X1Y5_LUT4AB/S2END[5] Tile_X1Y5_LUT4AB/S2END[6] Tile_X1Y5_LUT4AB/S2END[7]
+ Tile_X1Y5_LUT4AB/S2MID[0] Tile_X1Y5_LUT4AB/S2MID[1] Tile_X1Y5_LUT4AB/S2MID[2] Tile_X1Y5_LUT4AB/S2MID[3]
+ Tile_X1Y5_LUT4AB/S2MID[4] Tile_X1Y5_LUT4AB/S2MID[5] Tile_X1Y5_LUT4AB/S2MID[6] Tile_X1Y5_LUT4AB/S2MID[7]
+ Tile_X1Y6_LUT4AB/S4END[0] Tile_X1Y6_LUT4AB/S4END[10] Tile_X1Y6_LUT4AB/S4END[11]
+ Tile_X1Y6_LUT4AB/S4END[12] Tile_X1Y6_LUT4AB/S4END[13] Tile_X1Y6_LUT4AB/S4END[14]
+ Tile_X1Y6_LUT4AB/S4END[15] Tile_X1Y6_LUT4AB/S4END[1] Tile_X1Y6_LUT4AB/S4END[2] Tile_X1Y6_LUT4AB/S4END[3]
+ Tile_X1Y6_LUT4AB/S4END[4] Tile_X1Y6_LUT4AB/S4END[5] Tile_X1Y6_LUT4AB/S4END[6] Tile_X1Y6_LUT4AB/S4END[7]
+ Tile_X1Y6_LUT4AB/S4END[8] Tile_X1Y6_LUT4AB/S4END[9] Tile_X1Y5_LUT4AB/S4END[0] Tile_X1Y5_LUT4AB/S4END[10]
+ Tile_X1Y5_LUT4AB/S4END[11] Tile_X1Y5_LUT4AB/S4END[12] Tile_X1Y5_LUT4AB/S4END[13]
+ Tile_X1Y5_LUT4AB/S4END[14] Tile_X1Y5_LUT4AB/S4END[15] Tile_X1Y5_LUT4AB/S4END[1]
+ Tile_X1Y5_LUT4AB/S4END[2] Tile_X1Y5_LUT4AB/S4END[3] Tile_X1Y5_LUT4AB/S4END[4] Tile_X1Y5_LUT4AB/S4END[5]
+ Tile_X1Y5_LUT4AB/S4END[6] Tile_X1Y5_LUT4AB/S4END[7] Tile_X1Y5_LUT4AB/S4END[8] Tile_X1Y5_LUT4AB/S4END[9]
+ Tile_X1Y6_LUT4AB/SS4END[0] Tile_X1Y6_LUT4AB/SS4END[10] Tile_X1Y6_LUT4AB/SS4END[11]
+ Tile_X1Y6_LUT4AB/SS4END[12] Tile_X1Y6_LUT4AB/SS4END[13] Tile_X1Y6_LUT4AB/SS4END[14]
+ Tile_X1Y6_LUT4AB/SS4END[15] Tile_X1Y6_LUT4AB/SS4END[1] Tile_X1Y6_LUT4AB/SS4END[2]
+ Tile_X1Y6_LUT4AB/SS4END[3] Tile_X1Y6_LUT4AB/SS4END[4] Tile_X1Y6_LUT4AB/SS4END[5]
+ Tile_X1Y6_LUT4AB/SS4END[6] Tile_X1Y6_LUT4AB/SS4END[7] Tile_X1Y6_LUT4AB/SS4END[8]
+ Tile_X1Y6_LUT4AB/SS4END[9] Tile_X1Y5_LUT4AB/SS4END[0] Tile_X1Y5_LUT4AB/SS4END[10]
+ Tile_X1Y5_LUT4AB/SS4END[11] Tile_X1Y5_LUT4AB/SS4END[12] Tile_X1Y5_LUT4AB/SS4END[13]
+ Tile_X1Y5_LUT4AB/SS4END[14] Tile_X1Y5_LUT4AB/SS4END[15] Tile_X1Y5_LUT4AB/SS4END[1]
+ Tile_X1Y5_LUT4AB/SS4END[2] Tile_X1Y5_LUT4AB/SS4END[3] Tile_X1Y5_LUT4AB/SS4END[4]
+ Tile_X1Y5_LUT4AB/SS4END[5] Tile_X1Y5_LUT4AB/SS4END[6] Tile_X1Y5_LUT4AB/SS4END[7]
+ Tile_X1Y5_LUT4AB/SS4END[8] Tile_X1Y5_LUT4AB/SS4END[9] Tile_X1Y5_LUT4AB/UserCLK Tile_X1Y4_LUT4AB/UserCLK
+ VGND VPWR Tile_X1Y5_LUT4AB/W1BEG[0] Tile_X1Y5_LUT4AB/W1BEG[1] Tile_X1Y5_LUT4AB/W1BEG[2]
+ Tile_X1Y5_LUT4AB/W1BEG[3] Tile_X2Y5_LUT4AB/W1BEG[0] Tile_X2Y5_LUT4AB/W1BEG[1] Tile_X2Y5_LUT4AB/W1BEG[2]
+ Tile_X2Y5_LUT4AB/W1BEG[3] Tile_X1Y5_LUT4AB/W2BEG[0] Tile_X1Y5_LUT4AB/W2BEG[1] Tile_X1Y5_LUT4AB/W2BEG[2]
+ Tile_X1Y5_LUT4AB/W2BEG[3] Tile_X1Y5_LUT4AB/W2BEG[4] Tile_X1Y5_LUT4AB/W2BEG[5] Tile_X1Y5_LUT4AB/W2BEG[6]
+ Tile_X1Y5_LUT4AB/W2BEG[7] Tile_X1Y5_LUT4AB/W2BEGb[0] Tile_X1Y5_LUT4AB/W2BEGb[1]
+ Tile_X1Y5_LUT4AB/W2BEGb[2] Tile_X1Y5_LUT4AB/W2BEGb[3] Tile_X1Y5_LUT4AB/W2BEGb[4]
+ Tile_X1Y5_LUT4AB/W2BEGb[5] Tile_X1Y5_LUT4AB/W2BEGb[6] Tile_X1Y5_LUT4AB/W2BEGb[7]
+ Tile_X1Y5_LUT4AB/W2END[0] Tile_X1Y5_LUT4AB/W2END[1] Tile_X1Y5_LUT4AB/W2END[2] Tile_X1Y5_LUT4AB/W2END[3]
+ Tile_X1Y5_LUT4AB/W2END[4] Tile_X1Y5_LUT4AB/W2END[5] Tile_X1Y5_LUT4AB/W2END[6] Tile_X1Y5_LUT4AB/W2END[7]
+ Tile_X2Y5_LUT4AB/W2BEG[0] Tile_X2Y5_LUT4AB/W2BEG[1] Tile_X2Y5_LUT4AB/W2BEG[2] Tile_X2Y5_LUT4AB/W2BEG[3]
+ Tile_X2Y5_LUT4AB/W2BEG[4] Tile_X2Y5_LUT4AB/W2BEG[5] Tile_X2Y5_LUT4AB/W2BEG[6] Tile_X2Y5_LUT4AB/W2BEG[7]
+ Tile_X1Y5_LUT4AB/W6BEG[0] Tile_X1Y5_LUT4AB/W6BEG[10] Tile_X1Y5_LUT4AB/W6BEG[11]
+ Tile_X1Y5_LUT4AB/W6BEG[1] Tile_X1Y5_LUT4AB/W6BEG[2] Tile_X1Y5_LUT4AB/W6BEG[3] Tile_X1Y5_LUT4AB/W6BEG[4]
+ Tile_X1Y5_LUT4AB/W6BEG[5] Tile_X1Y5_LUT4AB/W6BEG[6] Tile_X1Y5_LUT4AB/W6BEG[7] Tile_X1Y5_LUT4AB/W6BEG[8]
+ Tile_X1Y5_LUT4AB/W6BEG[9] Tile_X2Y5_LUT4AB/W6BEG[0] Tile_X2Y5_LUT4AB/W6BEG[10] Tile_X2Y5_LUT4AB/W6BEG[11]
+ Tile_X2Y5_LUT4AB/W6BEG[1] Tile_X2Y5_LUT4AB/W6BEG[2] Tile_X2Y5_LUT4AB/W6BEG[3] Tile_X2Y5_LUT4AB/W6BEG[4]
+ Tile_X2Y5_LUT4AB/W6BEG[5] Tile_X2Y5_LUT4AB/W6BEG[6] Tile_X2Y5_LUT4AB/W6BEG[7] Tile_X2Y5_LUT4AB/W6BEG[8]
+ Tile_X2Y5_LUT4AB/W6BEG[9] Tile_X1Y5_LUT4AB/WW4BEG[0] Tile_X1Y5_LUT4AB/WW4BEG[10]
+ Tile_X1Y5_LUT4AB/WW4BEG[11] Tile_X1Y5_LUT4AB/WW4BEG[12] Tile_X1Y5_LUT4AB/WW4BEG[13]
+ Tile_X1Y5_LUT4AB/WW4BEG[14] Tile_X1Y5_LUT4AB/WW4BEG[15] Tile_X1Y5_LUT4AB/WW4BEG[1]
+ Tile_X1Y5_LUT4AB/WW4BEG[2] Tile_X1Y5_LUT4AB/WW4BEG[3] Tile_X1Y5_LUT4AB/WW4BEG[4]
+ Tile_X1Y5_LUT4AB/WW4BEG[5] Tile_X1Y5_LUT4AB/WW4BEG[6] Tile_X1Y5_LUT4AB/WW4BEG[7]
+ Tile_X1Y5_LUT4AB/WW4BEG[8] Tile_X1Y5_LUT4AB/WW4BEG[9] Tile_X2Y5_LUT4AB/WW4BEG[0]
+ Tile_X2Y5_LUT4AB/WW4BEG[10] Tile_X2Y5_LUT4AB/WW4BEG[11] Tile_X2Y5_LUT4AB/WW4BEG[12]
+ Tile_X2Y5_LUT4AB/WW4BEG[13] Tile_X2Y5_LUT4AB/WW4BEG[14] Tile_X2Y5_LUT4AB/WW4BEG[15]
+ Tile_X2Y5_LUT4AB/WW4BEG[1] Tile_X2Y5_LUT4AB/WW4BEG[2] Tile_X2Y5_LUT4AB/WW4BEG[3]
+ Tile_X2Y5_LUT4AB/WW4BEG[4] Tile_X2Y5_LUT4AB/WW4BEG[5] Tile_X2Y5_LUT4AB/WW4BEG[6]
+ Tile_X2Y5_LUT4AB/WW4BEG[7] Tile_X2Y5_LUT4AB/WW4BEG[8] Tile_X2Y5_LUT4AB/WW4BEG[9]
+ LUT4AB
XTile_X5Y8_E_TT_IF Tile_X5Y8_CLK_TT_PROJECT Tile_X4Y8_LUT4AB/E1BEG[0] Tile_X4Y8_LUT4AB/E1BEG[1]
+ Tile_X4Y8_LUT4AB/E1BEG[2] Tile_X4Y8_LUT4AB/E1BEG[3] Tile_X5Y8_E_TT_IF/E2END[0] Tile_X5Y8_E_TT_IF/E2END[1]
+ Tile_X5Y8_E_TT_IF/E2END[2] Tile_X5Y8_E_TT_IF/E2END[3] Tile_X5Y8_E_TT_IF/E2END[4]
+ Tile_X5Y8_E_TT_IF/E2END[5] Tile_X5Y8_E_TT_IF/E2END[6] Tile_X5Y8_E_TT_IF/E2END[7]
+ Tile_X4Y8_LUT4AB/E2BEG[0] Tile_X4Y8_LUT4AB/E2BEG[1] Tile_X4Y8_LUT4AB/E2BEG[2] Tile_X4Y8_LUT4AB/E2BEG[3]
+ Tile_X4Y8_LUT4AB/E2BEG[4] Tile_X4Y8_LUT4AB/E2BEG[5] Tile_X4Y8_LUT4AB/E2BEG[6] Tile_X4Y8_LUT4AB/E2BEG[7]
+ Tile_X4Y8_LUT4AB/E6BEG[0] Tile_X4Y8_LUT4AB/E6BEG[10] Tile_X4Y8_LUT4AB/E6BEG[11]
+ Tile_X4Y8_LUT4AB/E6BEG[1] Tile_X4Y8_LUT4AB/E6BEG[2] Tile_X4Y8_LUT4AB/E6BEG[3] Tile_X4Y8_LUT4AB/E6BEG[4]
+ Tile_X4Y8_LUT4AB/E6BEG[5] Tile_X4Y8_LUT4AB/E6BEG[6] Tile_X4Y8_LUT4AB/E6BEG[7] Tile_X4Y8_LUT4AB/E6BEG[8]
+ Tile_X4Y8_LUT4AB/E6BEG[9] Tile_X4Y8_LUT4AB/EE4BEG[0] Tile_X4Y8_LUT4AB/EE4BEG[10]
+ Tile_X4Y8_LUT4AB/EE4BEG[11] Tile_X4Y8_LUT4AB/EE4BEG[12] Tile_X4Y8_LUT4AB/EE4BEG[13]
+ Tile_X4Y8_LUT4AB/EE4BEG[14] Tile_X4Y8_LUT4AB/EE4BEG[15] Tile_X4Y8_LUT4AB/EE4BEG[1]
+ Tile_X4Y8_LUT4AB/EE4BEG[2] Tile_X4Y8_LUT4AB/EE4BEG[3] Tile_X4Y8_LUT4AB/EE4BEG[4]
+ Tile_X4Y8_LUT4AB/EE4BEG[5] Tile_X4Y8_LUT4AB/EE4BEG[6] Tile_X4Y8_LUT4AB/EE4BEG[7]
+ Tile_X4Y8_LUT4AB/EE4BEG[8] Tile_X4Y8_LUT4AB/EE4BEG[9] Tile_X5Y8_ENA_TT_PROJECT Tile_X5Y8_E_TT_IF/FrameData[0]
+ Tile_X5Y8_E_TT_IF/FrameData[10] Tile_X5Y8_E_TT_IF/FrameData[11] Tile_X5Y8_E_TT_IF/FrameData[12]
+ Tile_X5Y8_E_TT_IF/FrameData[13] Tile_X5Y8_E_TT_IF/FrameData[14] Tile_X5Y8_E_TT_IF/FrameData[15]
+ Tile_X5Y8_E_TT_IF/FrameData[16] Tile_X5Y8_E_TT_IF/FrameData[17] Tile_X5Y8_E_TT_IF/FrameData[18]
+ Tile_X5Y8_E_TT_IF/FrameData[19] Tile_X5Y8_E_TT_IF/FrameData[1] Tile_X5Y8_E_TT_IF/FrameData[20]
+ Tile_X5Y8_E_TT_IF/FrameData[21] Tile_X5Y8_E_TT_IF/FrameData[22] Tile_X5Y8_E_TT_IF/FrameData[23]
+ Tile_X5Y8_E_TT_IF/FrameData[24] Tile_X5Y8_E_TT_IF/FrameData[25] Tile_X5Y8_E_TT_IF/FrameData[26]
+ Tile_X5Y8_E_TT_IF/FrameData[27] Tile_X5Y8_E_TT_IF/FrameData[28] Tile_X5Y8_E_TT_IF/FrameData[29]
+ Tile_X5Y8_E_TT_IF/FrameData[2] Tile_X5Y8_E_TT_IF/FrameData[30] Tile_X5Y8_E_TT_IF/FrameData[31]
+ Tile_X5Y8_E_TT_IF/FrameData[3] Tile_X5Y8_E_TT_IF/FrameData[4] Tile_X5Y8_E_TT_IF/FrameData[5]
+ Tile_X5Y8_E_TT_IF/FrameData[6] Tile_X5Y8_E_TT_IF/FrameData[7] Tile_X5Y8_E_TT_IF/FrameData[8]
+ Tile_X5Y8_E_TT_IF/FrameData[9] Tile_X5Y8_E_TT_IF/FrameData_O[0] Tile_X5Y8_E_TT_IF/FrameData_O[10]
+ Tile_X5Y8_E_TT_IF/FrameData_O[11] Tile_X5Y8_E_TT_IF/FrameData_O[12] Tile_X5Y8_E_TT_IF/FrameData_O[13]
+ Tile_X5Y8_E_TT_IF/FrameData_O[14] Tile_X5Y8_E_TT_IF/FrameData_O[15] Tile_X5Y8_E_TT_IF/FrameData_O[16]
+ Tile_X5Y8_E_TT_IF/FrameData_O[17] Tile_X5Y8_E_TT_IF/FrameData_O[18] Tile_X5Y8_E_TT_IF/FrameData_O[19]
+ Tile_X5Y8_E_TT_IF/FrameData_O[1] Tile_X5Y8_E_TT_IF/FrameData_O[20] Tile_X5Y8_E_TT_IF/FrameData_O[21]
+ Tile_X5Y8_E_TT_IF/FrameData_O[22] Tile_X5Y8_E_TT_IF/FrameData_O[23] Tile_X5Y8_E_TT_IF/FrameData_O[24]
+ Tile_X5Y8_E_TT_IF/FrameData_O[25] Tile_X5Y8_E_TT_IF/FrameData_O[26] Tile_X5Y8_E_TT_IF/FrameData_O[27]
+ Tile_X5Y8_E_TT_IF/FrameData_O[28] Tile_X5Y8_E_TT_IF/FrameData_O[29] Tile_X5Y8_E_TT_IF/FrameData_O[2]
+ Tile_X5Y8_E_TT_IF/FrameData_O[30] Tile_X5Y8_E_TT_IF/FrameData_O[31] Tile_X5Y8_E_TT_IF/FrameData_O[3]
+ Tile_X5Y8_E_TT_IF/FrameData_O[4] Tile_X5Y8_E_TT_IF/FrameData_O[5] Tile_X5Y8_E_TT_IF/FrameData_O[6]
+ Tile_X5Y8_E_TT_IF/FrameData_O[7] Tile_X5Y8_E_TT_IF/FrameData_O[8] Tile_X5Y8_E_TT_IF/FrameData_O[9]
+ Tile_X5Y8_E_TT_IF/FrameStrobe[0] Tile_X5Y8_E_TT_IF/FrameStrobe[10] Tile_X5Y8_E_TT_IF/FrameStrobe[11]
+ Tile_X5Y8_E_TT_IF/FrameStrobe[12] Tile_X5Y8_E_TT_IF/FrameStrobe[13] Tile_X5Y8_E_TT_IF/FrameStrobe[14]
+ Tile_X5Y8_E_TT_IF/FrameStrobe[15] Tile_X5Y8_E_TT_IF/FrameStrobe[16] Tile_X5Y8_E_TT_IF/FrameStrobe[17]
+ Tile_X5Y8_E_TT_IF/FrameStrobe[18] Tile_X5Y8_E_TT_IF/FrameStrobe[19] Tile_X5Y8_E_TT_IF/FrameStrobe[1]
+ Tile_X5Y8_E_TT_IF/FrameStrobe[2] Tile_X5Y8_E_TT_IF/FrameStrobe[3] Tile_X5Y8_E_TT_IF/FrameStrobe[4]
+ Tile_X5Y8_E_TT_IF/FrameStrobe[5] Tile_X5Y8_E_TT_IF/FrameStrobe[6] Tile_X5Y8_E_TT_IF/FrameStrobe[7]
+ Tile_X5Y8_E_TT_IF/FrameStrobe[8] Tile_X5Y8_E_TT_IF/FrameStrobe[9] Tile_X5Y7_E_TT_IF/FrameStrobe[0]
+ Tile_X5Y7_E_TT_IF/FrameStrobe[10] Tile_X5Y7_E_TT_IF/FrameStrobe[11] Tile_X5Y7_E_TT_IF/FrameStrobe[12]
+ Tile_X5Y7_E_TT_IF/FrameStrobe[13] Tile_X5Y7_E_TT_IF/FrameStrobe[14] Tile_X5Y7_E_TT_IF/FrameStrobe[15]
+ Tile_X5Y7_E_TT_IF/FrameStrobe[16] Tile_X5Y7_E_TT_IF/FrameStrobe[17] Tile_X5Y7_E_TT_IF/FrameStrobe[18]
+ Tile_X5Y7_E_TT_IF/FrameStrobe[19] Tile_X5Y7_E_TT_IF/FrameStrobe[1] Tile_X5Y7_E_TT_IF/FrameStrobe[2]
+ Tile_X5Y7_E_TT_IF/FrameStrobe[3] Tile_X5Y7_E_TT_IF/FrameStrobe[4] Tile_X5Y7_E_TT_IF/FrameStrobe[5]
+ Tile_X5Y7_E_TT_IF/FrameStrobe[6] Tile_X5Y7_E_TT_IF/FrameStrobe[7] Tile_X5Y7_E_TT_IF/FrameStrobe[8]
+ Tile_X5Y7_E_TT_IF/FrameStrobe[9] Tile_X5Y8_E_TT_IF/N1BEG[0] Tile_X5Y8_E_TT_IF/N1BEG[1]
+ Tile_X5Y8_E_TT_IF/N1BEG[2] Tile_X5Y8_E_TT_IF/N1BEG[3] Tile_X5Y9_SE_term/N1BEG[0]
+ Tile_X5Y9_SE_term/N1BEG[1] Tile_X5Y9_SE_term/N1BEG[2] Tile_X5Y9_SE_term/N1BEG[3]
+ Tile_X5Y8_E_TT_IF/N2BEG[0] Tile_X5Y8_E_TT_IF/N2BEG[1] Tile_X5Y8_E_TT_IF/N2BEG[2]
+ Tile_X5Y8_E_TT_IF/N2BEG[3] Tile_X5Y8_E_TT_IF/N2BEG[4] Tile_X5Y8_E_TT_IF/N2BEG[5]
+ Tile_X5Y8_E_TT_IF/N2BEG[6] Tile_X5Y8_E_TT_IF/N2BEG[7] Tile_X5Y7_E_TT_IF/N2END[0]
+ Tile_X5Y7_E_TT_IF/N2END[1] Tile_X5Y7_E_TT_IF/N2END[2] Tile_X5Y7_E_TT_IF/N2END[3]
+ Tile_X5Y7_E_TT_IF/N2END[4] Tile_X5Y7_E_TT_IF/N2END[5] Tile_X5Y7_E_TT_IF/N2END[6]
+ Tile_X5Y7_E_TT_IF/N2END[7] Tile_X5Y8_E_TT_IF/N2END[0] Tile_X5Y8_E_TT_IF/N2END[1]
+ Tile_X5Y8_E_TT_IF/N2END[2] Tile_X5Y8_E_TT_IF/N2END[3] Tile_X5Y8_E_TT_IF/N2END[4]
+ Tile_X5Y8_E_TT_IF/N2END[5] Tile_X5Y8_E_TT_IF/N2END[6] Tile_X5Y8_E_TT_IF/N2END[7]
+ Tile_X5Y9_SE_term/N2BEG[0] Tile_X5Y9_SE_term/N2BEG[1] Tile_X5Y9_SE_term/N2BEG[2]
+ Tile_X5Y9_SE_term/N2BEG[3] Tile_X5Y9_SE_term/N2BEG[4] Tile_X5Y9_SE_term/N2BEG[5]
+ Tile_X5Y9_SE_term/N2BEG[6] Tile_X5Y9_SE_term/N2BEG[7] Tile_X5Y8_E_TT_IF/N4BEG[0]
+ Tile_X5Y8_E_TT_IF/N4BEG[10] Tile_X5Y8_E_TT_IF/N4BEG[11] Tile_X5Y8_E_TT_IF/N4BEG[12]
+ Tile_X5Y8_E_TT_IF/N4BEG[13] Tile_X5Y8_E_TT_IF/N4BEG[14] Tile_X5Y8_E_TT_IF/N4BEG[15]
+ Tile_X5Y8_E_TT_IF/N4BEG[1] Tile_X5Y8_E_TT_IF/N4BEG[2] Tile_X5Y8_E_TT_IF/N4BEG[3]
+ Tile_X5Y8_E_TT_IF/N4BEG[4] Tile_X5Y8_E_TT_IF/N4BEG[5] Tile_X5Y8_E_TT_IF/N4BEG[6]
+ Tile_X5Y8_E_TT_IF/N4BEG[7] Tile_X5Y8_E_TT_IF/N4BEG[8] Tile_X5Y8_E_TT_IF/N4BEG[9]
+ Tile_X5Y9_SE_term/N4BEG[0] Tile_X5Y9_SE_term/N4BEG[10] Tile_X5Y9_SE_term/N4BEG[11]
+ Tile_X5Y9_SE_term/N4BEG[12] Tile_X5Y9_SE_term/N4BEG[13] Tile_X5Y9_SE_term/N4BEG[14]
+ Tile_X5Y9_SE_term/N4BEG[15] Tile_X5Y9_SE_term/N4BEG[1] Tile_X5Y9_SE_term/N4BEG[2]
+ Tile_X5Y9_SE_term/N4BEG[3] Tile_X5Y9_SE_term/N4BEG[4] Tile_X5Y9_SE_term/N4BEG[5]
+ Tile_X5Y9_SE_term/N4BEG[6] Tile_X5Y9_SE_term/N4BEG[7] Tile_X5Y9_SE_term/N4BEG[8]
+ Tile_X5Y9_SE_term/N4BEG[9] Tile_X5Y8_RST_N_TT_PROJECT Tile_X5Y9_SE_term/S1END[0]
+ Tile_X5Y9_SE_term/S1END[1] Tile_X5Y9_SE_term/S1END[2] Tile_X5Y9_SE_term/S1END[3]
+ Tile_X5Y8_E_TT_IF/S1END[0] Tile_X5Y8_E_TT_IF/S1END[1] Tile_X5Y8_E_TT_IF/S1END[2]
+ Tile_X5Y8_E_TT_IF/S1END[3] Tile_X5Y9_SE_term/S2MID[0] Tile_X5Y9_SE_term/S2MID[1]
+ Tile_X5Y9_SE_term/S2MID[2] Tile_X5Y9_SE_term/S2MID[3] Tile_X5Y9_SE_term/S2MID[4]
+ Tile_X5Y9_SE_term/S2MID[5] Tile_X5Y9_SE_term/S2MID[6] Tile_X5Y9_SE_term/S2MID[7]
+ Tile_X5Y9_SE_term/S2END[0] Tile_X5Y9_SE_term/S2END[1] Tile_X5Y9_SE_term/S2END[2]
+ Tile_X5Y9_SE_term/S2END[3] Tile_X5Y9_SE_term/S2END[4] Tile_X5Y9_SE_term/S2END[5]
+ Tile_X5Y9_SE_term/S2END[6] Tile_X5Y9_SE_term/S2END[7] Tile_X5Y8_E_TT_IF/S2END[0]
+ Tile_X5Y8_E_TT_IF/S2END[1] Tile_X5Y8_E_TT_IF/S2END[2] Tile_X5Y8_E_TT_IF/S2END[3]
+ Tile_X5Y8_E_TT_IF/S2END[4] Tile_X5Y8_E_TT_IF/S2END[5] Tile_X5Y8_E_TT_IF/S2END[6]
+ Tile_X5Y8_E_TT_IF/S2END[7] Tile_X5Y8_E_TT_IF/S2MID[0] Tile_X5Y8_E_TT_IF/S2MID[1]
+ Tile_X5Y8_E_TT_IF/S2MID[2] Tile_X5Y8_E_TT_IF/S2MID[3] Tile_X5Y8_E_TT_IF/S2MID[4]
+ Tile_X5Y8_E_TT_IF/S2MID[5] Tile_X5Y8_E_TT_IF/S2MID[6] Tile_X5Y8_E_TT_IF/S2MID[7]
+ Tile_X5Y9_SE_term/S4END[0] Tile_X5Y9_SE_term/S4END[10] Tile_X5Y9_SE_term/S4END[11]
+ Tile_X5Y9_SE_term/S4END[12] Tile_X5Y9_SE_term/S4END[13] Tile_X5Y9_SE_term/S4END[14]
+ Tile_X5Y9_SE_term/S4END[15] Tile_X5Y9_SE_term/S4END[1] Tile_X5Y9_SE_term/S4END[2]
+ Tile_X5Y9_SE_term/S4END[3] Tile_X5Y9_SE_term/S4END[4] Tile_X5Y9_SE_term/S4END[5]
+ Tile_X5Y9_SE_term/S4END[6] Tile_X5Y9_SE_term/S4END[7] Tile_X5Y9_SE_term/S4END[8]
+ Tile_X5Y9_SE_term/S4END[9] Tile_X5Y8_E_TT_IF/S4END[0] Tile_X5Y8_E_TT_IF/S4END[10]
+ Tile_X5Y8_E_TT_IF/S4END[11] Tile_X5Y8_E_TT_IF/S4END[12] Tile_X5Y8_E_TT_IF/S4END[13]
+ Tile_X5Y8_E_TT_IF/S4END[14] Tile_X5Y8_E_TT_IF/S4END[15] Tile_X5Y8_E_TT_IF/S4END[1]
+ Tile_X5Y8_E_TT_IF/S4END[2] Tile_X5Y8_E_TT_IF/S4END[3] Tile_X5Y8_E_TT_IF/S4END[4]
+ Tile_X5Y8_E_TT_IF/S4END[5] Tile_X5Y8_E_TT_IF/S4END[6] Tile_X5Y8_E_TT_IF/S4END[7]
+ Tile_X5Y8_E_TT_IF/S4END[8] Tile_X5Y8_E_TT_IF/S4END[9] Tile_X5Y8_UIO_IN_TT_PROJECT0
+ Tile_X5Y8_UIO_IN_TT_PROJECT1 Tile_X5Y8_UIO_IN_TT_PROJECT2 Tile_X5Y8_UIO_IN_TT_PROJECT3
+ Tile_X5Y8_UIO_IN_TT_PROJECT4 Tile_X5Y8_UIO_IN_TT_PROJECT5 Tile_X5Y8_UIO_IN_TT_PROJECT6
+ Tile_X5Y8_UIO_IN_TT_PROJECT7 Tile_X5Y8_UIO_OE_TT_PROJECT0 Tile_X5Y8_UIO_OE_TT_PROJECT1
+ Tile_X5Y8_UIO_OE_TT_PROJECT2 Tile_X5Y8_UIO_OE_TT_PROJECT3 Tile_X5Y8_UIO_OE_TT_PROJECT4
+ Tile_X5Y8_UIO_OE_TT_PROJECT5 Tile_X5Y8_UIO_OE_TT_PROJECT6 Tile_X5Y8_UIO_OE_TT_PROJECT7
+ Tile_X5Y8_UIO_OUT_TT_PROJECT0 Tile_X5Y8_UIO_OUT_TT_PROJECT1 Tile_X5Y8_UIO_OUT_TT_PROJECT2
+ Tile_X5Y8_UIO_OUT_TT_PROJECT3 Tile_X5Y8_UIO_OUT_TT_PROJECT4 Tile_X5Y8_UIO_OUT_TT_PROJECT5
+ Tile_X5Y8_UIO_OUT_TT_PROJECT6 Tile_X5Y8_UIO_OUT_TT_PROJECT7 Tile_X5Y8_UI_IN_TT_PROJECT0
+ Tile_X5Y8_UI_IN_TT_PROJECT1 Tile_X5Y8_UI_IN_TT_PROJECT2 Tile_X5Y8_UI_IN_TT_PROJECT3
+ Tile_X5Y8_UI_IN_TT_PROJECT4 Tile_X5Y8_UI_IN_TT_PROJECT5 Tile_X5Y8_UI_IN_TT_PROJECT6
+ Tile_X5Y8_UI_IN_TT_PROJECT7 Tile_X5Y8_UO_OUT_TT_PROJECT0 Tile_X5Y8_UO_OUT_TT_PROJECT1
+ Tile_X5Y8_UO_OUT_TT_PROJECT2 Tile_X5Y8_UO_OUT_TT_PROJECT3 Tile_X5Y8_UO_OUT_TT_PROJECT4
+ Tile_X5Y8_UO_OUT_TT_PROJECT5 Tile_X5Y8_UO_OUT_TT_PROJECT6 Tile_X5Y8_UO_OUT_TT_PROJECT7
+ Tile_X5Y8_E_TT_IF/UserCLK Tile_X5Y7_E_TT_IF/UserCLK VGND VPWR Tile_X4Y8_LUT4AB/W1END[0]
+ Tile_X4Y8_LUT4AB/W1END[1] Tile_X4Y8_LUT4AB/W1END[2] Tile_X4Y8_LUT4AB/W1END[3] Tile_X4Y8_LUT4AB/W2MID[0]
+ Tile_X4Y8_LUT4AB/W2MID[1] Tile_X4Y8_LUT4AB/W2MID[2] Tile_X4Y8_LUT4AB/W2MID[3] Tile_X4Y8_LUT4AB/W2MID[4]
+ Tile_X4Y8_LUT4AB/W2MID[5] Tile_X4Y8_LUT4AB/W2MID[6] Tile_X4Y8_LUT4AB/W2MID[7] Tile_X4Y8_LUT4AB/W2END[0]
+ Tile_X4Y8_LUT4AB/W2END[1] Tile_X4Y8_LUT4AB/W2END[2] Tile_X4Y8_LUT4AB/W2END[3] Tile_X4Y8_LUT4AB/W2END[4]
+ Tile_X4Y8_LUT4AB/W2END[5] Tile_X4Y8_LUT4AB/W2END[6] Tile_X4Y8_LUT4AB/W2END[7] Tile_X4Y8_LUT4AB/W6END[0]
+ Tile_X4Y8_LUT4AB/W6END[10] Tile_X4Y8_LUT4AB/W6END[11] Tile_X4Y8_LUT4AB/W6END[1]
+ Tile_X4Y8_LUT4AB/W6END[2] Tile_X4Y8_LUT4AB/W6END[3] Tile_X4Y8_LUT4AB/W6END[4] Tile_X4Y8_LUT4AB/W6END[5]
+ Tile_X4Y8_LUT4AB/W6END[6] Tile_X4Y8_LUT4AB/W6END[7] Tile_X4Y8_LUT4AB/W6END[8] Tile_X4Y8_LUT4AB/W6END[9]
+ Tile_X4Y8_LUT4AB/WW4END[0] Tile_X4Y8_LUT4AB/WW4END[10] Tile_X4Y8_LUT4AB/WW4END[11]
+ Tile_X4Y8_LUT4AB/WW4END[12] Tile_X4Y8_LUT4AB/WW4END[13] Tile_X4Y8_LUT4AB/WW4END[14]
+ Tile_X4Y8_LUT4AB/WW4END[15] Tile_X4Y8_LUT4AB/WW4END[1] Tile_X4Y8_LUT4AB/WW4END[2]
+ Tile_X4Y8_LUT4AB/WW4END[3] Tile_X4Y8_LUT4AB/WW4END[4] Tile_X4Y8_LUT4AB/WW4END[5]
+ Tile_X4Y8_LUT4AB/WW4END[6] Tile_X4Y8_LUT4AB/WW4END[7] Tile_X4Y8_LUT4AB/WW4END[8]
+ Tile_X4Y8_LUT4AB/WW4END[9] E_TT_IF
.ends

