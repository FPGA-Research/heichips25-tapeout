module eFPGA (Tile_X0Y2_CLK_TT_PROJECT,
    Tile_X0Y2_ENA_TT_PROJECT,
    Tile_X0Y2_RST_N_TT_PROJECT,
    Tile_X0Y2_UIO_IN_TT_PROJECT0,
    Tile_X0Y2_UIO_IN_TT_PROJECT1,
    Tile_X0Y2_UIO_IN_TT_PROJECT2,
    Tile_X0Y2_UIO_IN_TT_PROJECT3,
    Tile_X0Y2_UIO_IN_TT_PROJECT4,
    Tile_X0Y2_UIO_IN_TT_PROJECT5,
    Tile_X0Y2_UIO_IN_TT_PROJECT6,
    Tile_X0Y2_UIO_IN_TT_PROJECT7,
    Tile_X0Y2_UIO_OE_TT_PROJECT0,
    Tile_X0Y2_UIO_OE_TT_PROJECT1,
    Tile_X0Y2_UIO_OE_TT_PROJECT2,
    Tile_X0Y2_UIO_OE_TT_PROJECT3,
    Tile_X0Y2_UIO_OE_TT_PROJECT4,
    Tile_X0Y2_UIO_OE_TT_PROJECT5,
    Tile_X0Y2_UIO_OE_TT_PROJECT6,
    Tile_X0Y2_UIO_OE_TT_PROJECT7,
    Tile_X0Y2_UIO_OUT_TT_PROJECT0,
    Tile_X0Y2_UIO_OUT_TT_PROJECT1,
    Tile_X0Y2_UIO_OUT_TT_PROJECT2,
    Tile_X0Y2_UIO_OUT_TT_PROJECT3,
    Tile_X0Y2_UIO_OUT_TT_PROJECT4,
    Tile_X0Y2_UIO_OUT_TT_PROJECT5,
    Tile_X0Y2_UIO_OUT_TT_PROJECT6,
    Tile_X0Y2_UIO_OUT_TT_PROJECT7,
    Tile_X0Y2_UI_IN_TT_PROJECT0,
    Tile_X0Y2_UI_IN_TT_PROJECT1,
    Tile_X0Y2_UI_IN_TT_PROJECT2,
    Tile_X0Y2_UI_IN_TT_PROJECT3,
    Tile_X0Y2_UI_IN_TT_PROJECT4,
    Tile_X0Y2_UI_IN_TT_PROJECT5,
    Tile_X0Y2_UI_IN_TT_PROJECT6,
    Tile_X0Y2_UI_IN_TT_PROJECT7,
    Tile_X0Y2_UO_OUT_TT_PROJECT0,
    Tile_X0Y2_UO_OUT_TT_PROJECT1,
    Tile_X0Y2_UO_OUT_TT_PROJECT2,
    Tile_X0Y2_UO_OUT_TT_PROJECT3,
    Tile_X0Y2_UO_OUT_TT_PROJECT4,
    Tile_X0Y2_UO_OUT_TT_PROJECT5,
    Tile_X0Y2_UO_OUT_TT_PROJECT6,
    Tile_X0Y2_UO_OUT_TT_PROJECT7,
    Tile_X0Y3_CLK_TT_PROJECT,
    Tile_X0Y3_ENA_TT_PROJECT,
    Tile_X0Y3_RST_N_TT_PROJECT,
    Tile_X0Y3_UIO_IN_TT_PROJECT0,
    Tile_X0Y3_UIO_IN_TT_PROJECT1,
    Tile_X0Y3_UIO_IN_TT_PROJECT2,
    Tile_X0Y3_UIO_IN_TT_PROJECT3,
    Tile_X0Y3_UIO_IN_TT_PROJECT4,
    Tile_X0Y3_UIO_IN_TT_PROJECT5,
    Tile_X0Y3_UIO_IN_TT_PROJECT6,
    Tile_X0Y3_UIO_IN_TT_PROJECT7,
    Tile_X0Y3_UIO_OE_TT_PROJECT0,
    Tile_X0Y3_UIO_OE_TT_PROJECT1,
    Tile_X0Y3_UIO_OE_TT_PROJECT2,
    Tile_X0Y3_UIO_OE_TT_PROJECT3,
    Tile_X0Y3_UIO_OE_TT_PROJECT4,
    Tile_X0Y3_UIO_OE_TT_PROJECT5,
    Tile_X0Y3_UIO_OE_TT_PROJECT6,
    Tile_X0Y3_UIO_OE_TT_PROJECT7,
    Tile_X0Y3_UIO_OUT_TT_PROJECT0,
    Tile_X0Y3_UIO_OUT_TT_PROJECT1,
    Tile_X0Y3_UIO_OUT_TT_PROJECT2,
    Tile_X0Y3_UIO_OUT_TT_PROJECT3,
    Tile_X0Y3_UIO_OUT_TT_PROJECT4,
    Tile_X0Y3_UIO_OUT_TT_PROJECT5,
    Tile_X0Y3_UIO_OUT_TT_PROJECT6,
    Tile_X0Y3_UIO_OUT_TT_PROJECT7,
    Tile_X0Y3_UI_IN_TT_PROJECT0,
    Tile_X0Y3_UI_IN_TT_PROJECT1,
    Tile_X0Y3_UI_IN_TT_PROJECT2,
    Tile_X0Y3_UI_IN_TT_PROJECT3,
    Tile_X0Y3_UI_IN_TT_PROJECT4,
    Tile_X0Y3_UI_IN_TT_PROJECT5,
    Tile_X0Y3_UI_IN_TT_PROJECT6,
    Tile_X0Y3_UI_IN_TT_PROJECT7,
    Tile_X0Y3_UO_OUT_TT_PROJECT0,
    Tile_X0Y3_UO_OUT_TT_PROJECT1,
    Tile_X0Y3_UO_OUT_TT_PROJECT2,
    Tile_X0Y3_UO_OUT_TT_PROJECT3,
    Tile_X0Y3_UO_OUT_TT_PROJECT4,
    Tile_X0Y3_UO_OUT_TT_PROJECT5,
    Tile_X0Y3_UO_OUT_TT_PROJECT6,
    Tile_X0Y3_UO_OUT_TT_PROJECT7,
    Tile_X0Y4_CLK_TT_PROJECT,
    Tile_X0Y4_ENA_TT_PROJECT,
    Tile_X0Y4_RST_N_TT_PROJECT,
    Tile_X0Y4_UIO_IN_TT_PROJECT0,
    Tile_X0Y4_UIO_IN_TT_PROJECT1,
    Tile_X0Y4_UIO_IN_TT_PROJECT2,
    Tile_X0Y4_UIO_IN_TT_PROJECT3,
    Tile_X0Y4_UIO_IN_TT_PROJECT4,
    Tile_X0Y4_UIO_IN_TT_PROJECT5,
    Tile_X0Y4_UIO_IN_TT_PROJECT6,
    Tile_X0Y4_UIO_IN_TT_PROJECT7,
    Tile_X0Y4_UIO_OE_TT_PROJECT0,
    Tile_X0Y4_UIO_OE_TT_PROJECT1,
    Tile_X0Y4_UIO_OE_TT_PROJECT2,
    Tile_X0Y4_UIO_OE_TT_PROJECT3,
    Tile_X0Y4_UIO_OE_TT_PROJECT4,
    Tile_X0Y4_UIO_OE_TT_PROJECT5,
    Tile_X0Y4_UIO_OE_TT_PROJECT6,
    Tile_X0Y4_UIO_OE_TT_PROJECT7,
    Tile_X0Y4_UIO_OUT_TT_PROJECT0,
    Tile_X0Y4_UIO_OUT_TT_PROJECT1,
    Tile_X0Y4_UIO_OUT_TT_PROJECT2,
    Tile_X0Y4_UIO_OUT_TT_PROJECT3,
    Tile_X0Y4_UIO_OUT_TT_PROJECT4,
    Tile_X0Y4_UIO_OUT_TT_PROJECT5,
    Tile_X0Y4_UIO_OUT_TT_PROJECT6,
    Tile_X0Y4_UIO_OUT_TT_PROJECT7,
    Tile_X0Y4_UI_IN_TT_PROJECT0,
    Tile_X0Y4_UI_IN_TT_PROJECT1,
    Tile_X0Y4_UI_IN_TT_PROJECT2,
    Tile_X0Y4_UI_IN_TT_PROJECT3,
    Tile_X0Y4_UI_IN_TT_PROJECT4,
    Tile_X0Y4_UI_IN_TT_PROJECT5,
    Tile_X0Y4_UI_IN_TT_PROJECT6,
    Tile_X0Y4_UI_IN_TT_PROJECT7,
    Tile_X0Y4_UO_OUT_TT_PROJECT0,
    Tile_X0Y4_UO_OUT_TT_PROJECT1,
    Tile_X0Y4_UO_OUT_TT_PROJECT2,
    Tile_X0Y4_UO_OUT_TT_PROJECT3,
    Tile_X0Y4_UO_OUT_TT_PROJECT4,
    Tile_X0Y4_UO_OUT_TT_PROJECT5,
    Tile_X0Y4_UO_OUT_TT_PROJECT6,
    Tile_X0Y4_UO_OUT_TT_PROJECT7,
    Tile_X0Y5_CLK_TT_PROJECT,
    Tile_X0Y5_ENA_TT_PROJECT,
    Tile_X0Y5_RST_N_TT_PROJECT,
    Tile_X0Y5_UIO_IN_TT_PROJECT0,
    Tile_X0Y5_UIO_IN_TT_PROJECT1,
    Tile_X0Y5_UIO_IN_TT_PROJECT2,
    Tile_X0Y5_UIO_IN_TT_PROJECT3,
    Tile_X0Y5_UIO_IN_TT_PROJECT4,
    Tile_X0Y5_UIO_IN_TT_PROJECT5,
    Tile_X0Y5_UIO_IN_TT_PROJECT6,
    Tile_X0Y5_UIO_IN_TT_PROJECT7,
    Tile_X0Y5_UIO_OE_TT_PROJECT0,
    Tile_X0Y5_UIO_OE_TT_PROJECT1,
    Tile_X0Y5_UIO_OE_TT_PROJECT2,
    Tile_X0Y5_UIO_OE_TT_PROJECT3,
    Tile_X0Y5_UIO_OE_TT_PROJECT4,
    Tile_X0Y5_UIO_OE_TT_PROJECT5,
    Tile_X0Y5_UIO_OE_TT_PROJECT6,
    Tile_X0Y5_UIO_OE_TT_PROJECT7,
    Tile_X0Y5_UIO_OUT_TT_PROJECT0,
    Tile_X0Y5_UIO_OUT_TT_PROJECT1,
    Tile_X0Y5_UIO_OUT_TT_PROJECT2,
    Tile_X0Y5_UIO_OUT_TT_PROJECT3,
    Tile_X0Y5_UIO_OUT_TT_PROJECT4,
    Tile_X0Y5_UIO_OUT_TT_PROJECT5,
    Tile_X0Y5_UIO_OUT_TT_PROJECT6,
    Tile_X0Y5_UIO_OUT_TT_PROJECT7,
    Tile_X0Y5_UI_IN_TT_PROJECT0,
    Tile_X0Y5_UI_IN_TT_PROJECT1,
    Tile_X0Y5_UI_IN_TT_PROJECT2,
    Tile_X0Y5_UI_IN_TT_PROJECT3,
    Tile_X0Y5_UI_IN_TT_PROJECT4,
    Tile_X0Y5_UI_IN_TT_PROJECT5,
    Tile_X0Y5_UI_IN_TT_PROJECT6,
    Tile_X0Y5_UI_IN_TT_PROJECT7,
    Tile_X0Y5_UO_OUT_TT_PROJECT0,
    Tile_X0Y5_UO_OUT_TT_PROJECT1,
    Tile_X0Y5_UO_OUT_TT_PROJECT2,
    Tile_X0Y5_UO_OUT_TT_PROJECT3,
    Tile_X0Y5_UO_OUT_TT_PROJECT4,
    Tile_X0Y5_UO_OUT_TT_PROJECT5,
    Tile_X0Y5_UO_OUT_TT_PROJECT6,
    Tile_X0Y5_UO_OUT_TT_PROJECT7,
    Tile_X0Y6_CLK_TT_PROJECT,
    Tile_X0Y6_ENA_TT_PROJECT,
    Tile_X0Y6_RST_N_TT_PROJECT,
    Tile_X0Y6_UIO_IN_TT_PROJECT0,
    Tile_X0Y6_UIO_IN_TT_PROJECT1,
    Tile_X0Y6_UIO_IN_TT_PROJECT2,
    Tile_X0Y6_UIO_IN_TT_PROJECT3,
    Tile_X0Y6_UIO_IN_TT_PROJECT4,
    Tile_X0Y6_UIO_IN_TT_PROJECT5,
    Tile_X0Y6_UIO_IN_TT_PROJECT6,
    Tile_X0Y6_UIO_IN_TT_PROJECT7,
    Tile_X0Y6_UIO_OE_TT_PROJECT0,
    Tile_X0Y6_UIO_OE_TT_PROJECT1,
    Tile_X0Y6_UIO_OE_TT_PROJECT2,
    Tile_X0Y6_UIO_OE_TT_PROJECT3,
    Tile_X0Y6_UIO_OE_TT_PROJECT4,
    Tile_X0Y6_UIO_OE_TT_PROJECT5,
    Tile_X0Y6_UIO_OE_TT_PROJECT6,
    Tile_X0Y6_UIO_OE_TT_PROJECT7,
    Tile_X0Y6_UIO_OUT_TT_PROJECT0,
    Tile_X0Y6_UIO_OUT_TT_PROJECT1,
    Tile_X0Y6_UIO_OUT_TT_PROJECT2,
    Tile_X0Y6_UIO_OUT_TT_PROJECT3,
    Tile_X0Y6_UIO_OUT_TT_PROJECT4,
    Tile_X0Y6_UIO_OUT_TT_PROJECT5,
    Tile_X0Y6_UIO_OUT_TT_PROJECT6,
    Tile_X0Y6_UIO_OUT_TT_PROJECT7,
    Tile_X0Y6_UI_IN_TT_PROJECT0,
    Tile_X0Y6_UI_IN_TT_PROJECT1,
    Tile_X0Y6_UI_IN_TT_PROJECT2,
    Tile_X0Y6_UI_IN_TT_PROJECT3,
    Tile_X0Y6_UI_IN_TT_PROJECT4,
    Tile_X0Y6_UI_IN_TT_PROJECT5,
    Tile_X0Y6_UI_IN_TT_PROJECT6,
    Tile_X0Y6_UI_IN_TT_PROJECT7,
    Tile_X0Y6_UO_OUT_TT_PROJECT0,
    Tile_X0Y6_UO_OUT_TT_PROJECT1,
    Tile_X0Y6_UO_OUT_TT_PROJECT2,
    Tile_X0Y6_UO_OUT_TT_PROJECT3,
    Tile_X0Y6_UO_OUT_TT_PROJECT4,
    Tile_X0Y6_UO_OUT_TT_PROJECT5,
    Tile_X0Y6_UO_OUT_TT_PROJECT6,
    Tile_X0Y6_UO_OUT_TT_PROJECT7,
    Tile_X0Y7_CLK_TT_PROJECT,
    Tile_X0Y7_ENA_TT_PROJECT,
    Tile_X0Y7_RST_N_TT_PROJECT,
    Tile_X0Y7_UIO_IN_TT_PROJECT0,
    Tile_X0Y7_UIO_IN_TT_PROJECT1,
    Tile_X0Y7_UIO_IN_TT_PROJECT2,
    Tile_X0Y7_UIO_IN_TT_PROJECT3,
    Tile_X0Y7_UIO_IN_TT_PROJECT4,
    Tile_X0Y7_UIO_IN_TT_PROJECT5,
    Tile_X0Y7_UIO_IN_TT_PROJECT6,
    Tile_X0Y7_UIO_IN_TT_PROJECT7,
    Tile_X0Y7_UIO_OE_TT_PROJECT0,
    Tile_X0Y7_UIO_OE_TT_PROJECT1,
    Tile_X0Y7_UIO_OE_TT_PROJECT2,
    Tile_X0Y7_UIO_OE_TT_PROJECT3,
    Tile_X0Y7_UIO_OE_TT_PROJECT4,
    Tile_X0Y7_UIO_OE_TT_PROJECT5,
    Tile_X0Y7_UIO_OE_TT_PROJECT6,
    Tile_X0Y7_UIO_OE_TT_PROJECT7,
    Tile_X0Y7_UIO_OUT_TT_PROJECT0,
    Tile_X0Y7_UIO_OUT_TT_PROJECT1,
    Tile_X0Y7_UIO_OUT_TT_PROJECT2,
    Tile_X0Y7_UIO_OUT_TT_PROJECT3,
    Tile_X0Y7_UIO_OUT_TT_PROJECT4,
    Tile_X0Y7_UIO_OUT_TT_PROJECT5,
    Tile_X0Y7_UIO_OUT_TT_PROJECT6,
    Tile_X0Y7_UIO_OUT_TT_PROJECT7,
    Tile_X0Y7_UI_IN_TT_PROJECT0,
    Tile_X0Y7_UI_IN_TT_PROJECT1,
    Tile_X0Y7_UI_IN_TT_PROJECT2,
    Tile_X0Y7_UI_IN_TT_PROJECT3,
    Tile_X0Y7_UI_IN_TT_PROJECT4,
    Tile_X0Y7_UI_IN_TT_PROJECT5,
    Tile_X0Y7_UI_IN_TT_PROJECT6,
    Tile_X0Y7_UI_IN_TT_PROJECT7,
    Tile_X0Y7_UO_OUT_TT_PROJECT0,
    Tile_X0Y7_UO_OUT_TT_PROJECT1,
    Tile_X0Y7_UO_OUT_TT_PROJECT2,
    Tile_X0Y7_UO_OUT_TT_PROJECT3,
    Tile_X0Y7_UO_OUT_TT_PROJECT4,
    Tile_X0Y7_UO_OUT_TT_PROJECT5,
    Tile_X0Y7_UO_OUT_TT_PROJECT6,
    Tile_X0Y7_UO_OUT_TT_PROJECT7,
    Tile_X0Y8_CLK_TT_PROJECT,
    Tile_X0Y8_ENA_TT_PROJECT,
    Tile_X0Y8_RST_N_TT_PROJECT,
    Tile_X0Y8_UIO_IN_TT_PROJECT0,
    Tile_X0Y8_UIO_IN_TT_PROJECT1,
    Tile_X0Y8_UIO_IN_TT_PROJECT2,
    Tile_X0Y8_UIO_IN_TT_PROJECT3,
    Tile_X0Y8_UIO_IN_TT_PROJECT4,
    Tile_X0Y8_UIO_IN_TT_PROJECT5,
    Tile_X0Y8_UIO_IN_TT_PROJECT6,
    Tile_X0Y8_UIO_IN_TT_PROJECT7,
    Tile_X0Y8_UIO_OE_TT_PROJECT0,
    Tile_X0Y8_UIO_OE_TT_PROJECT1,
    Tile_X0Y8_UIO_OE_TT_PROJECT2,
    Tile_X0Y8_UIO_OE_TT_PROJECT3,
    Tile_X0Y8_UIO_OE_TT_PROJECT4,
    Tile_X0Y8_UIO_OE_TT_PROJECT5,
    Tile_X0Y8_UIO_OE_TT_PROJECT6,
    Tile_X0Y8_UIO_OE_TT_PROJECT7,
    Tile_X0Y8_UIO_OUT_TT_PROJECT0,
    Tile_X0Y8_UIO_OUT_TT_PROJECT1,
    Tile_X0Y8_UIO_OUT_TT_PROJECT2,
    Tile_X0Y8_UIO_OUT_TT_PROJECT3,
    Tile_X0Y8_UIO_OUT_TT_PROJECT4,
    Tile_X0Y8_UIO_OUT_TT_PROJECT5,
    Tile_X0Y8_UIO_OUT_TT_PROJECT6,
    Tile_X0Y8_UIO_OUT_TT_PROJECT7,
    Tile_X0Y8_UI_IN_TT_PROJECT0,
    Tile_X0Y8_UI_IN_TT_PROJECT1,
    Tile_X0Y8_UI_IN_TT_PROJECT2,
    Tile_X0Y8_UI_IN_TT_PROJECT3,
    Tile_X0Y8_UI_IN_TT_PROJECT4,
    Tile_X0Y8_UI_IN_TT_PROJECT5,
    Tile_X0Y8_UI_IN_TT_PROJECT6,
    Tile_X0Y8_UI_IN_TT_PROJECT7,
    Tile_X0Y8_UO_OUT_TT_PROJECT0,
    Tile_X0Y8_UO_OUT_TT_PROJECT1,
    Tile_X0Y8_UO_OUT_TT_PROJECT2,
    Tile_X0Y8_UO_OUT_TT_PROJECT3,
    Tile_X0Y8_UO_OUT_TT_PROJECT4,
    Tile_X0Y8_UO_OUT_TT_PROJECT5,
    Tile_X0Y8_UO_OUT_TT_PROJECT6,
    Tile_X0Y8_UO_OUT_TT_PROJECT7,
    Tile_X1Y0_A_I_top,
    Tile_X1Y0_A_O_top,
    Tile_X1Y0_A_T_top,
    Tile_X1Y0_B_I_top,
    Tile_X1Y0_B_O_top,
    Tile_X1Y0_B_T_top,
    Tile_X1Y0_C_I_top,
    Tile_X1Y0_C_O_top,
    Tile_X1Y0_C_T_top,
    Tile_X1Y0_D_I_top,
    Tile_X1Y0_D_O_top,
    Tile_X1Y0_D_T_top,
    Tile_X1Y9_A_I_top,
    Tile_X1Y9_A_O_top,
    Tile_X1Y9_A_T_top,
    Tile_X1Y9_B_I_top,
    Tile_X1Y9_B_O_top,
    Tile_X1Y9_B_T_top,
    Tile_X1Y9_C_I_top,
    Tile_X1Y9_C_O_top,
    Tile_X1Y9_C_T_top,
    Tile_X1Y9_D_I_top,
    Tile_X1Y9_D_O_top,
    Tile_X1Y9_D_T_top,
    Tile_X2Y0_A_I_top,
    Tile_X2Y0_A_O_top,
    Tile_X2Y0_A_T_top,
    Tile_X2Y0_B_I_top,
    Tile_X2Y0_B_O_top,
    Tile_X2Y0_B_T_top,
    Tile_X2Y0_C_I_top,
    Tile_X2Y0_C_O_top,
    Tile_X2Y0_C_T_top,
    Tile_X2Y0_D_I_top,
    Tile_X2Y0_D_O_top,
    Tile_X2Y0_D_T_top,
    Tile_X2Y9_A_I_top,
    Tile_X2Y9_A_O_top,
    Tile_X2Y9_A_T_top,
    Tile_X2Y9_B_I_top,
    Tile_X2Y9_B_O_top,
    Tile_X2Y9_B_T_top,
    Tile_X2Y9_C_I_top,
    Tile_X2Y9_C_O_top,
    Tile_X2Y9_C_T_top,
    Tile_X2Y9_D_I_top,
    Tile_X2Y9_D_O_top,
    Tile_X2Y9_D_T_top,
    Tile_X3Y0_A_I_top,
    Tile_X3Y0_A_O_top,
    Tile_X3Y0_A_T_top,
    Tile_X3Y0_B_I_top,
    Tile_X3Y0_B_O_top,
    Tile_X3Y0_B_T_top,
    Tile_X3Y0_C_I_top,
    Tile_X3Y0_C_O_top,
    Tile_X3Y0_C_T_top,
    Tile_X3Y0_D_I_top,
    Tile_X3Y0_D_O_top,
    Tile_X3Y0_D_T_top,
    Tile_X3Y9_A_I_top,
    Tile_X3Y9_A_O_top,
    Tile_X3Y9_A_T_top,
    Tile_X3Y9_B_I_top,
    Tile_X3Y9_B_O_top,
    Tile_X3Y9_B_T_top,
    Tile_X3Y9_C_I_top,
    Tile_X3Y9_C_O_top,
    Tile_X3Y9_C_T_top,
    Tile_X3Y9_D_I_top,
    Tile_X3Y9_D_O_top,
    Tile_X3Y9_D_T_top,
    Tile_X4Y0_A_I_top,
    Tile_X4Y0_A_O_top,
    Tile_X4Y0_A_T_top,
    Tile_X4Y0_B_I_top,
    Tile_X4Y0_B_O_top,
    Tile_X4Y0_B_T_top,
    Tile_X4Y0_C_I_top,
    Tile_X4Y0_C_O_top,
    Tile_X4Y0_C_T_top,
    Tile_X4Y0_D_I_top,
    Tile_X4Y0_D_O_top,
    Tile_X4Y0_D_T_top,
    Tile_X4Y9_A_I_top,
    Tile_X4Y9_A_O_top,
    Tile_X4Y9_A_T_top,
    Tile_X4Y9_B_I_top,
    Tile_X4Y9_B_O_top,
    Tile_X4Y9_B_T_top,
    Tile_X4Y9_C_I_top,
    Tile_X4Y9_C_O_top,
    Tile_X4Y9_C_T_top,
    Tile_X4Y9_D_I_top,
    Tile_X4Y9_D_O_top,
    Tile_X4Y9_D_T_top,
    Tile_X5Y2_ADDR_SRAM0,
    Tile_X5Y2_ADDR_SRAM1,
    Tile_X5Y2_ADDR_SRAM2,
    Tile_X5Y2_ADDR_SRAM3,
    Tile_X5Y2_ADDR_SRAM4,
    Tile_X5Y2_ADDR_SRAM5,
    Tile_X5Y2_ADDR_SRAM6,
    Tile_X5Y2_ADDR_SRAM7,
    Tile_X5Y2_ADDR_SRAM8,
    Tile_X5Y2_ADDR_SRAM9,
    Tile_X5Y2_BM_SRAM0,
    Tile_X5Y2_BM_SRAM1,
    Tile_X5Y2_BM_SRAM10,
    Tile_X5Y2_BM_SRAM11,
    Tile_X5Y2_BM_SRAM12,
    Tile_X5Y2_BM_SRAM13,
    Tile_X5Y2_BM_SRAM14,
    Tile_X5Y2_BM_SRAM15,
    Tile_X5Y2_BM_SRAM16,
    Tile_X5Y2_BM_SRAM17,
    Tile_X5Y2_BM_SRAM18,
    Tile_X5Y2_BM_SRAM19,
    Tile_X5Y2_BM_SRAM2,
    Tile_X5Y2_BM_SRAM20,
    Tile_X5Y2_BM_SRAM21,
    Tile_X5Y2_BM_SRAM22,
    Tile_X5Y2_BM_SRAM23,
    Tile_X5Y2_BM_SRAM24,
    Tile_X5Y2_BM_SRAM25,
    Tile_X5Y2_BM_SRAM26,
    Tile_X5Y2_BM_SRAM27,
    Tile_X5Y2_BM_SRAM28,
    Tile_X5Y2_BM_SRAM29,
    Tile_X5Y2_BM_SRAM3,
    Tile_X5Y2_BM_SRAM30,
    Tile_X5Y2_BM_SRAM31,
    Tile_X5Y2_BM_SRAM4,
    Tile_X5Y2_BM_SRAM5,
    Tile_X5Y2_BM_SRAM6,
    Tile_X5Y2_BM_SRAM7,
    Tile_X5Y2_BM_SRAM8,
    Tile_X5Y2_BM_SRAM9,
    Tile_X5Y2_CLK_SRAM,
    Tile_X5Y2_CONFIGURED_top,
    Tile_X5Y2_DIN_SRAM0,
    Tile_X5Y2_DIN_SRAM1,
    Tile_X5Y2_DIN_SRAM10,
    Tile_X5Y2_DIN_SRAM11,
    Tile_X5Y2_DIN_SRAM12,
    Tile_X5Y2_DIN_SRAM13,
    Tile_X5Y2_DIN_SRAM14,
    Tile_X5Y2_DIN_SRAM15,
    Tile_X5Y2_DIN_SRAM16,
    Tile_X5Y2_DIN_SRAM17,
    Tile_X5Y2_DIN_SRAM18,
    Tile_X5Y2_DIN_SRAM19,
    Tile_X5Y2_DIN_SRAM2,
    Tile_X5Y2_DIN_SRAM20,
    Tile_X5Y2_DIN_SRAM21,
    Tile_X5Y2_DIN_SRAM22,
    Tile_X5Y2_DIN_SRAM23,
    Tile_X5Y2_DIN_SRAM24,
    Tile_X5Y2_DIN_SRAM25,
    Tile_X5Y2_DIN_SRAM26,
    Tile_X5Y2_DIN_SRAM27,
    Tile_X5Y2_DIN_SRAM28,
    Tile_X5Y2_DIN_SRAM29,
    Tile_X5Y2_DIN_SRAM3,
    Tile_X5Y2_DIN_SRAM30,
    Tile_X5Y2_DIN_SRAM31,
    Tile_X5Y2_DIN_SRAM4,
    Tile_X5Y2_DIN_SRAM5,
    Tile_X5Y2_DIN_SRAM6,
    Tile_X5Y2_DIN_SRAM7,
    Tile_X5Y2_DIN_SRAM8,
    Tile_X5Y2_DIN_SRAM9,
    Tile_X5Y2_DOUT_SRAM0,
    Tile_X5Y2_DOUT_SRAM1,
    Tile_X5Y2_DOUT_SRAM10,
    Tile_X5Y2_DOUT_SRAM11,
    Tile_X5Y2_DOUT_SRAM12,
    Tile_X5Y2_DOUT_SRAM13,
    Tile_X5Y2_DOUT_SRAM14,
    Tile_X5Y2_DOUT_SRAM15,
    Tile_X5Y2_DOUT_SRAM16,
    Tile_X5Y2_DOUT_SRAM17,
    Tile_X5Y2_DOUT_SRAM18,
    Tile_X5Y2_DOUT_SRAM19,
    Tile_X5Y2_DOUT_SRAM2,
    Tile_X5Y2_DOUT_SRAM20,
    Tile_X5Y2_DOUT_SRAM21,
    Tile_X5Y2_DOUT_SRAM22,
    Tile_X5Y2_DOUT_SRAM23,
    Tile_X5Y2_DOUT_SRAM24,
    Tile_X5Y2_DOUT_SRAM25,
    Tile_X5Y2_DOUT_SRAM26,
    Tile_X5Y2_DOUT_SRAM27,
    Tile_X5Y2_DOUT_SRAM28,
    Tile_X5Y2_DOUT_SRAM29,
    Tile_X5Y2_DOUT_SRAM3,
    Tile_X5Y2_DOUT_SRAM30,
    Tile_X5Y2_DOUT_SRAM31,
    Tile_X5Y2_DOUT_SRAM4,
    Tile_X5Y2_DOUT_SRAM5,
    Tile_X5Y2_DOUT_SRAM6,
    Tile_X5Y2_DOUT_SRAM7,
    Tile_X5Y2_DOUT_SRAM8,
    Tile_X5Y2_DOUT_SRAM9,
    Tile_X5Y2_MEN_SRAM,
    Tile_X5Y2_REN_SRAM,
    Tile_X5Y2_TIE_HIGH_SRAM,
    Tile_X5Y2_TIE_LOW_SRAM,
    Tile_X5Y2_WEN_SRAM,
    Tile_X5Y4_CLK_TT_PROJECT,
    Tile_X5Y4_ENA_TT_PROJECT,
    Tile_X5Y4_RST_N_TT_PROJECT,
    Tile_X5Y4_UIO_IN_TT_PROJECT0,
    Tile_X5Y4_UIO_IN_TT_PROJECT1,
    Tile_X5Y4_UIO_IN_TT_PROJECT2,
    Tile_X5Y4_UIO_IN_TT_PROJECT3,
    Tile_X5Y4_UIO_IN_TT_PROJECT4,
    Tile_X5Y4_UIO_IN_TT_PROJECT5,
    Tile_X5Y4_UIO_IN_TT_PROJECT6,
    Tile_X5Y4_UIO_IN_TT_PROJECT7,
    Tile_X5Y4_UIO_OE_TT_PROJECT0,
    Tile_X5Y4_UIO_OE_TT_PROJECT1,
    Tile_X5Y4_UIO_OE_TT_PROJECT2,
    Tile_X5Y4_UIO_OE_TT_PROJECT3,
    Tile_X5Y4_UIO_OE_TT_PROJECT4,
    Tile_X5Y4_UIO_OE_TT_PROJECT5,
    Tile_X5Y4_UIO_OE_TT_PROJECT6,
    Tile_X5Y4_UIO_OE_TT_PROJECT7,
    Tile_X5Y4_UIO_OUT_TT_PROJECT0,
    Tile_X5Y4_UIO_OUT_TT_PROJECT1,
    Tile_X5Y4_UIO_OUT_TT_PROJECT2,
    Tile_X5Y4_UIO_OUT_TT_PROJECT3,
    Tile_X5Y4_UIO_OUT_TT_PROJECT4,
    Tile_X5Y4_UIO_OUT_TT_PROJECT5,
    Tile_X5Y4_UIO_OUT_TT_PROJECT6,
    Tile_X5Y4_UIO_OUT_TT_PROJECT7,
    Tile_X5Y4_UI_IN_TT_PROJECT0,
    Tile_X5Y4_UI_IN_TT_PROJECT1,
    Tile_X5Y4_UI_IN_TT_PROJECT2,
    Tile_X5Y4_UI_IN_TT_PROJECT3,
    Tile_X5Y4_UI_IN_TT_PROJECT4,
    Tile_X5Y4_UI_IN_TT_PROJECT5,
    Tile_X5Y4_UI_IN_TT_PROJECT6,
    Tile_X5Y4_UI_IN_TT_PROJECT7,
    Tile_X5Y4_UO_OUT_TT_PROJECT0,
    Tile_X5Y4_UO_OUT_TT_PROJECT1,
    Tile_X5Y4_UO_OUT_TT_PROJECT2,
    Tile_X5Y4_UO_OUT_TT_PROJECT3,
    Tile_X5Y4_UO_OUT_TT_PROJECT4,
    Tile_X5Y4_UO_OUT_TT_PROJECT5,
    Tile_X5Y4_UO_OUT_TT_PROJECT6,
    Tile_X5Y4_UO_OUT_TT_PROJECT7,
    Tile_X5Y5_CLK_TT_PROJECT,
    Tile_X5Y5_ENA_TT_PROJECT,
    Tile_X5Y5_RST_N_TT_PROJECT,
    Tile_X5Y5_UIO_IN_TT_PROJECT0,
    Tile_X5Y5_UIO_IN_TT_PROJECT1,
    Tile_X5Y5_UIO_IN_TT_PROJECT2,
    Tile_X5Y5_UIO_IN_TT_PROJECT3,
    Tile_X5Y5_UIO_IN_TT_PROJECT4,
    Tile_X5Y5_UIO_IN_TT_PROJECT5,
    Tile_X5Y5_UIO_IN_TT_PROJECT6,
    Tile_X5Y5_UIO_IN_TT_PROJECT7,
    Tile_X5Y5_UIO_OE_TT_PROJECT0,
    Tile_X5Y5_UIO_OE_TT_PROJECT1,
    Tile_X5Y5_UIO_OE_TT_PROJECT2,
    Tile_X5Y5_UIO_OE_TT_PROJECT3,
    Tile_X5Y5_UIO_OE_TT_PROJECT4,
    Tile_X5Y5_UIO_OE_TT_PROJECT5,
    Tile_X5Y5_UIO_OE_TT_PROJECT6,
    Tile_X5Y5_UIO_OE_TT_PROJECT7,
    Tile_X5Y5_UIO_OUT_TT_PROJECT0,
    Tile_X5Y5_UIO_OUT_TT_PROJECT1,
    Tile_X5Y5_UIO_OUT_TT_PROJECT2,
    Tile_X5Y5_UIO_OUT_TT_PROJECT3,
    Tile_X5Y5_UIO_OUT_TT_PROJECT4,
    Tile_X5Y5_UIO_OUT_TT_PROJECT5,
    Tile_X5Y5_UIO_OUT_TT_PROJECT6,
    Tile_X5Y5_UIO_OUT_TT_PROJECT7,
    Tile_X5Y5_UI_IN_TT_PROJECT0,
    Tile_X5Y5_UI_IN_TT_PROJECT1,
    Tile_X5Y5_UI_IN_TT_PROJECT2,
    Tile_X5Y5_UI_IN_TT_PROJECT3,
    Tile_X5Y5_UI_IN_TT_PROJECT4,
    Tile_X5Y5_UI_IN_TT_PROJECT5,
    Tile_X5Y5_UI_IN_TT_PROJECT6,
    Tile_X5Y5_UI_IN_TT_PROJECT7,
    Tile_X5Y5_UO_OUT_TT_PROJECT0,
    Tile_X5Y5_UO_OUT_TT_PROJECT1,
    Tile_X5Y5_UO_OUT_TT_PROJECT2,
    Tile_X5Y5_UO_OUT_TT_PROJECT3,
    Tile_X5Y5_UO_OUT_TT_PROJECT4,
    Tile_X5Y5_UO_OUT_TT_PROJECT5,
    Tile_X5Y5_UO_OUT_TT_PROJECT6,
    Tile_X5Y5_UO_OUT_TT_PROJECT7,
    Tile_X5Y6_CLK_TT_PROJECT,
    Tile_X5Y6_ENA_TT_PROJECT,
    Tile_X5Y6_RST_N_TT_PROJECT,
    Tile_X5Y6_UIO_IN_TT_PROJECT0,
    Tile_X5Y6_UIO_IN_TT_PROJECT1,
    Tile_X5Y6_UIO_IN_TT_PROJECT2,
    Tile_X5Y6_UIO_IN_TT_PROJECT3,
    Tile_X5Y6_UIO_IN_TT_PROJECT4,
    Tile_X5Y6_UIO_IN_TT_PROJECT5,
    Tile_X5Y6_UIO_IN_TT_PROJECT6,
    Tile_X5Y6_UIO_IN_TT_PROJECT7,
    Tile_X5Y6_UIO_OE_TT_PROJECT0,
    Tile_X5Y6_UIO_OE_TT_PROJECT1,
    Tile_X5Y6_UIO_OE_TT_PROJECT2,
    Tile_X5Y6_UIO_OE_TT_PROJECT3,
    Tile_X5Y6_UIO_OE_TT_PROJECT4,
    Tile_X5Y6_UIO_OE_TT_PROJECT5,
    Tile_X5Y6_UIO_OE_TT_PROJECT6,
    Tile_X5Y6_UIO_OE_TT_PROJECT7,
    Tile_X5Y6_UIO_OUT_TT_PROJECT0,
    Tile_X5Y6_UIO_OUT_TT_PROJECT1,
    Tile_X5Y6_UIO_OUT_TT_PROJECT2,
    Tile_X5Y6_UIO_OUT_TT_PROJECT3,
    Tile_X5Y6_UIO_OUT_TT_PROJECT4,
    Tile_X5Y6_UIO_OUT_TT_PROJECT5,
    Tile_X5Y6_UIO_OUT_TT_PROJECT6,
    Tile_X5Y6_UIO_OUT_TT_PROJECT7,
    Tile_X5Y6_UI_IN_TT_PROJECT0,
    Tile_X5Y6_UI_IN_TT_PROJECT1,
    Tile_X5Y6_UI_IN_TT_PROJECT2,
    Tile_X5Y6_UI_IN_TT_PROJECT3,
    Tile_X5Y6_UI_IN_TT_PROJECT4,
    Tile_X5Y6_UI_IN_TT_PROJECT5,
    Tile_X5Y6_UI_IN_TT_PROJECT6,
    Tile_X5Y6_UI_IN_TT_PROJECT7,
    Tile_X5Y6_UO_OUT_TT_PROJECT0,
    Tile_X5Y6_UO_OUT_TT_PROJECT1,
    Tile_X5Y6_UO_OUT_TT_PROJECT2,
    Tile_X5Y6_UO_OUT_TT_PROJECT3,
    Tile_X5Y6_UO_OUT_TT_PROJECT4,
    Tile_X5Y6_UO_OUT_TT_PROJECT5,
    Tile_X5Y6_UO_OUT_TT_PROJECT6,
    Tile_X5Y6_UO_OUT_TT_PROJECT7,
    Tile_X5Y7_CLK_TT_PROJECT,
    Tile_X5Y7_ENA_TT_PROJECT,
    Tile_X5Y7_RST_N_TT_PROJECT,
    Tile_X5Y7_UIO_IN_TT_PROJECT0,
    Tile_X5Y7_UIO_IN_TT_PROJECT1,
    Tile_X5Y7_UIO_IN_TT_PROJECT2,
    Tile_X5Y7_UIO_IN_TT_PROJECT3,
    Tile_X5Y7_UIO_IN_TT_PROJECT4,
    Tile_X5Y7_UIO_IN_TT_PROJECT5,
    Tile_X5Y7_UIO_IN_TT_PROJECT6,
    Tile_X5Y7_UIO_IN_TT_PROJECT7,
    Tile_X5Y7_UIO_OE_TT_PROJECT0,
    Tile_X5Y7_UIO_OE_TT_PROJECT1,
    Tile_X5Y7_UIO_OE_TT_PROJECT2,
    Tile_X5Y7_UIO_OE_TT_PROJECT3,
    Tile_X5Y7_UIO_OE_TT_PROJECT4,
    Tile_X5Y7_UIO_OE_TT_PROJECT5,
    Tile_X5Y7_UIO_OE_TT_PROJECT6,
    Tile_X5Y7_UIO_OE_TT_PROJECT7,
    Tile_X5Y7_UIO_OUT_TT_PROJECT0,
    Tile_X5Y7_UIO_OUT_TT_PROJECT1,
    Tile_X5Y7_UIO_OUT_TT_PROJECT2,
    Tile_X5Y7_UIO_OUT_TT_PROJECT3,
    Tile_X5Y7_UIO_OUT_TT_PROJECT4,
    Tile_X5Y7_UIO_OUT_TT_PROJECT5,
    Tile_X5Y7_UIO_OUT_TT_PROJECT6,
    Tile_X5Y7_UIO_OUT_TT_PROJECT7,
    Tile_X5Y7_UI_IN_TT_PROJECT0,
    Tile_X5Y7_UI_IN_TT_PROJECT1,
    Tile_X5Y7_UI_IN_TT_PROJECT2,
    Tile_X5Y7_UI_IN_TT_PROJECT3,
    Tile_X5Y7_UI_IN_TT_PROJECT4,
    Tile_X5Y7_UI_IN_TT_PROJECT5,
    Tile_X5Y7_UI_IN_TT_PROJECT6,
    Tile_X5Y7_UI_IN_TT_PROJECT7,
    Tile_X5Y7_UO_OUT_TT_PROJECT0,
    Tile_X5Y7_UO_OUT_TT_PROJECT1,
    Tile_X5Y7_UO_OUT_TT_PROJECT2,
    Tile_X5Y7_UO_OUT_TT_PROJECT3,
    Tile_X5Y7_UO_OUT_TT_PROJECT4,
    Tile_X5Y7_UO_OUT_TT_PROJECT5,
    Tile_X5Y7_UO_OUT_TT_PROJECT6,
    Tile_X5Y7_UO_OUT_TT_PROJECT7,
    Tile_X5Y8_CLK_TT_PROJECT,
    Tile_X5Y8_ENA_TT_PROJECT,
    Tile_X5Y8_RST_N_TT_PROJECT,
    Tile_X5Y8_UIO_IN_TT_PROJECT0,
    Tile_X5Y8_UIO_IN_TT_PROJECT1,
    Tile_X5Y8_UIO_IN_TT_PROJECT2,
    Tile_X5Y8_UIO_IN_TT_PROJECT3,
    Tile_X5Y8_UIO_IN_TT_PROJECT4,
    Tile_X5Y8_UIO_IN_TT_PROJECT5,
    Tile_X5Y8_UIO_IN_TT_PROJECT6,
    Tile_X5Y8_UIO_IN_TT_PROJECT7,
    Tile_X5Y8_UIO_OE_TT_PROJECT0,
    Tile_X5Y8_UIO_OE_TT_PROJECT1,
    Tile_X5Y8_UIO_OE_TT_PROJECT2,
    Tile_X5Y8_UIO_OE_TT_PROJECT3,
    Tile_X5Y8_UIO_OE_TT_PROJECT4,
    Tile_X5Y8_UIO_OE_TT_PROJECT5,
    Tile_X5Y8_UIO_OE_TT_PROJECT6,
    Tile_X5Y8_UIO_OE_TT_PROJECT7,
    Tile_X5Y8_UIO_OUT_TT_PROJECT0,
    Tile_X5Y8_UIO_OUT_TT_PROJECT1,
    Tile_X5Y8_UIO_OUT_TT_PROJECT2,
    Tile_X5Y8_UIO_OUT_TT_PROJECT3,
    Tile_X5Y8_UIO_OUT_TT_PROJECT4,
    Tile_X5Y8_UIO_OUT_TT_PROJECT5,
    Tile_X5Y8_UIO_OUT_TT_PROJECT6,
    Tile_X5Y8_UIO_OUT_TT_PROJECT7,
    Tile_X5Y8_UI_IN_TT_PROJECT0,
    Tile_X5Y8_UI_IN_TT_PROJECT1,
    Tile_X5Y8_UI_IN_TT_PROJECT2,
    Tile_X5Y8_UI_IN_TT_PROJECT3,
    Tile_X5Y8_UI_IN_TT_PROJECT4,
    Tile_X5Y8_UI_IN_TT_PROJECT5,
    Tile_X5Y8_UI_IN_TT_PROJECT6,
    Tile_X5Y8_UI_IN_TT_PROJECT7,
    Tile_X5Y8_UO_OUT_TT_PROJECT0,
    Tile_X5Y8_UO_OUT_TT_PROJECT1,
    Tile_X5Y8_UO_OUT_TT_PROJECT2,
    Tile_X5Y8_UO_OUT_TT_PROJECT3,
    Tile_X5Y8_UO_OUT_TT_PROJECT4,
    Tile_X5Y8_UO_OUT_TT_PROJECT5,
    Tile_X5Y8_UO_OUT_TT_PROJECT6,
    Tile_X5Y8_UO_OUT_TT_PROJECT7,
    UserCLK,
    VPWR,
    VGND,
    FrameData,
    FrameStrobe);
 output Tile_X0Y2_CLK_TT_PROJECT;
 output Tile_X0Y2_ENA_TT_PROJECT;
 output Tile_X0Y2_RST_N_TT_PROJECT;
 output Tile_X0Y2_UIO_IN_TT_PROJECT0;
 output Tile_X0Y2_UIO_IN_TT_PROJECT1;
 output Tile_X0Y2_UIO_IN_TT_PROJECT2;
 output Tile_X0Y2_UIO_IN_TT_PROJECT3;
 output Tile_X0Y2_UIO_IN_TT_PROJECT4;
 output Tile_X0Y2_UIO_IN_TT_PROJECT5;
 output Tile_X0Y2_UIO_IN_TT_PROJECT6;
 output Tile_X0Y2_UIO_IN_TT_PROJECT7;
 input Tile_X0Y2_UIO_OE_TT_PROJECT0;
 input Tile_X0Y2_UIO_OE_TT_PROJECT1;
 input Tile_X0Y2_UIO_OE_TT_PROJECT2;
 input Tile_X0Y2_UIO_OE_TT_PROJECT3;
 input Tile_X0Y2_UIO_OE_TT_PROJECT4;
 input Tile_X0Y2_UIO_OE_TT_PROJECT5;
 input Tile_X0Y2_UIO_OE_TT_PROJECT6;
 input Tile_X0Y2_UIO_OE_TT_PROJECT7;
 input Tile_X0Y2_UIO_OUT_TT_PROJECT0;
 input Tile_X0Y2_UIO_OUT_TT_PROJECT1;
 input Tile_X0Y2_UIO_OUT_TT_PROJECT2;
 input Tile_X0Y2_UIO_OUT_TT_PROJECT3;
 input Tile_X0Y2_UIO_OUT_TT_PROJECT4;
 input Tile_X0Y2_UIO_OUT_TT_PROJECT5;
 input Tile_X0Y2_UIO_OUT_TT_PROJECT6;
 input Tile_X0Y2_UIO_OUT_TT_PROJECT7;
 output Tile_X0Y2_UI_IN_TT_PROJECT0;
 output Tile_X0Y2_UI_IN_TT_PROJECT1;
 output Tile_X0Y2_UI_IN_TT_PROJECT2;
 output Tile_X0Y2_UI_IN_TT_PROJECT3;
 output Tile_X0Y2_UI_IN_TT_PROJECT4;
 output Tile_X0Y2_UI_IN_TT_PROJECT5;
 output Tile_X0Y2_UI_IN_TT_PROJECT6;
 output Tile_X0Y2_UI_IN_TT_PROJECT7;
 input Tile_X0Y2_UO_OUT_TT_PROJECT0;
 input Tile_X0Y2_UO_OUT_TT_PROJECT1;
 input Tile_X0Y2_UO_OUT_TT_PROJECT2;
 input Tile_X0Y2_UO_OUT_TT_PROJECT3;
 input Tile_X0Y2_UO_OUT_TT_PROJECT4;
 input Tile_X0Y2_UO_OUT_TT_PROJECT5;
 input Tile_X0Y2_UO_OUT_TT_PROJECT6;
 input Tile_X0Y2_UO_OUT_TT_PROJECT7;
 output Tile_X0Y3_CLK_TT_PROJECT;
 output Tile_X0Y3_ENA_TT_PROJECT;
 output Tile_X0Y3_RST_N_TT_PROJECT;
 output Tile_X0Y3_UIO_IN_TT_PROJECT0;
 output Tile_X0Y3_UIO_IN_TT_PROJECT1;
 output Tile_X0Y3_UIO_IN_TT_PROJECT2;
 output Tile_X0Y3_UIO_IN_TT_PROJECT3;
 output Tile_X0Y3_UIO_IN_TT_PROJECT4;
 output Tile_X0Y3_UIO_IN_TT_PROJECT5;
 output Tile_X0Y3_UIO_IN_TT_PROJECT6;
 output Tile_X0Y3_UIO_IN_TT_PROJECT7;
 input Tile_X0Y3_UIO_OE_TT_PROJECT0;
 input Tile_X0Y3_UIO_OE_TT_PROJECT1;
 input Tile_X0Y3_UIO_OE_TT_PROJECT2;
 input Tile_X0Y3_UIO_OE_TT_PROJECT3;
 input Tile_X0Y3_UIO_OE_TT_PROJECT4;
 input Tile_X0Y3_UIO_OE_TT_PROJECT5;
 input Tile_X0Y3_UIO_OE_TT_PROJECT6;
 input Tile_X0Y3_UIO_OE_TT_PROJECT7;
 input Tile_X0Y3_UIO_OUT_TT_PROJECT0;
 input Tile_X0Y3_UIO_OUT_TT_PROJECT1;
 input Tile_X0Y3_UIO_OUT_TT_PROJECT2;
 input Tile_X0Y3_UIO_OUT_TT_PROJECT3;
 input Tile_X0Y3_UIO_OUT_TT_PROJECT4;
 input Tile_X0Y3_UIO_OUT_TT_PROJECT5;
 input Tile_X0Y3_UIO_OUT_TT_PROJECT6;
 input Tile_X0Y3_UIO_OUT_TT_PROJECT7;
 output Tile_X0Y3_UI_IN_TT_PROJECT0;
 output Tile_X0Y3_UI_IN_TT_PROJECT1;
 output Tile_X0Y3_UI_IN_TT_PROJECT2;
 output Tile_X0Y3_UI_IN_TT_PROJECT3;
 output Tile_X0Y3_UI_IN_TT_PROJECT4;
 output Tile_X0Y3_UI_IN_TT_PROJECT5;
 output Tile_X0Y3_UI_IN_TT_PROJECT6;
 output Tile_X0Y3_UI_IN_TT_PROJECT7;
 input Tile_X0Y3_UO_OUT_TT_PROJECT0;
 input Tile_X0Y3_UO_OUT_TT_PROJECT1;
 input Tile_X0Y3_UO_OUT_TT_PROJECT2;
 input Tile_X0Y3_UO_OUT_TT_PROJECT3;
 input Tile_X0Y3_UO_OUT_TT_PROJECT4;
 input Tile_X0Y3_UO_OUT_TT_PROJECT5;
 input Tile_X0Y3_UO_OUT_TT_PROJECT6;
 input Tile_X0Y3_UO_OUT_TT_PROJECT7;
 output Tile_X0Y4_CLK_TT_PROJECT;
 output Tile_X0Y4_ENA_TT_PROJECT;
 output Tile_X0Y4_RST_N_TT_PROJECT;
 output Tile_X0Y4_UIO_IN_TT_PROJECT0;
 output Tile_X0Y4_UIO_IN_TT_PROJECT1;
 output Tile_X0Y4_UIO_IN_TT_PROJECT2;
 output Tile_X0Y4_UIO_IN_TT_PROJECT3;
 output Tile_X0Y4_UIO_IN_TT_PROJECT4;
 output Tile_X0Y4_UIO_IN_TT_PROJECT5;
 output Tile_X0Y4_UIO_IN_TT_PROJECT6;
 output Tile_X0Y4_UIO_IN_TT_PROJECT7;
 input Tile_X0Y4_UIO_OE_TT_PROJECT0;
 input Tile_X0Y4_UIO_OE_TT_PROJECT1;
 input Tile_X0Y4_UIO_OE_TT_PROJECT2;
 input Tile_X0Y4_UIO_OE_TT_PROJECT3;
 input Tile_X0Y4_UIO_OE_TT_PROJECT4;
 input Tile_X0Y4_UIO_OE_TT_PROJECT5;
 input Tile_X0Y4_UIO_OE_TT_PROJECT6;
 input Tile_X0Y4_UIO_OE_TT_PROJECT7;
 input Tile_X0Y4_UIO_OUT_TT_PROJECT0;
 input Tile_X0Y4_UIO_OUT_TT_PROJECT1;
 input Tile_X0Y4_UIO_OUT_TT_PROJECT2;
 input Tile_X0Y4_UIO_OUT_TT_PROJECT3;
 input Tile_X0Y4_UIO_OUT_TT_PROJECT4;
 input Tile_X0Y4_UIO_OUT_TT_PROJECT5;
 input Tile_X0Y4_UIO_OUT_TT_PROJECT6;
 input Tile_X0Y4_UIO_OUT_TT_PROJECT7;
 output Tile_X0Y4_UI_IN_TT_PROJECT0;
 output Tile_X0Y4_UI_IN_TT_PROJECT1;
 output Tile_X0Y4_UI_IN_TT_PROJECT2;
 output Tile_X0Y4_UI_IN_TT_PROJECT3;
 output Tile_X0Y4_UI_IN_TT_PROJECT4;
 output Tile_X0Y4_UI_IN_TT_PROJECT5;
 output Tile_X0Y4_UI_IN_TT_PROJECT6;
 output Tile_X0Y4_UI_IN_TT_PROJECT7;
 input Tile_X0Y4_UO_OUT_TT_PROJECT0;
 input Tile_X0Y4_UO_OUT_TT_PROJECT1;
 input Tile_X0Y4_UO_OUT_TT_PROJECT2;
 input Tile_X0Y4_UO_OUT_TT_PROJECT3;
 input Tile_X0Y4_UO_OUT_TT_PROJECT4;
 input Tile_X0Y4_UO_OUT_TT_PROJECT5;
 input Tile_X0Y4_UO_OUT_TT_PROJECT6;
 input Tile_X0Y4_UO_OUT_TT_PROJECT7;
 output Tile_X0Y5_CLK_TT_PROJECT;
 output Tile_X0Y5_ENA_TT_PROJECT;
 output Tile_X0Y5_RST_N_TT_PROJECT;
 output Tile_X0Y5_UIO_IN_TT_PROJECT0;
 output Tile_X0Y5_UIO_IN_TT_PROJECT1;
 output Tile_X0Y5_UIO_IN_TT_PROJECT2;
 output Tile_X0Y5_UIO_IN_TT_PROJECT3;
 output Tile_X0Y5_UIO_IN_TT_PROJECT4;
 output Tile_X0Y5_UIO_IN_TT_PROJECT5;
 output Tile_X0Y5_UIO_IN_TT_PROJECT6;
 output Tile_X0Y5_UIO_IN_TT_PROJECT7;
 input Tile_X0Y5_UIO_OE_TT_PROJECT0;
 input Tile_X0Y5_UIO_OE_TT_PROJECT1;
 input Tile_X0Y5_UIO_OE_TT_PROJECT2;
 input Tile_X0Y5_UIO_OE_TT_PROJECT3;
 input Tile_X0Y5_UIO_OE_TT_PROJECT4;
 input Tile_X0Y5_UIO_OE_TT_PROJECT5;
 input Tile_X0Y5_UIO_OE_TT_PROJECT6;
 input Tile_X0Y5_UIO_OE_TT_PROJECT7;
 input Tile_X0Y5_UIO_OUT_TT_PROJECT0;
 input Tile_X0Y5_UIO_OUT_TT_PROJECT1;
 input Tile_X0Y5_UIO_OUT_TT_PROJECT2;
 input Tile_X0Y5_UIO_OUT_TT_PROJECT3;
 input Tile_X0Y5_UIO_OUT_TT_PROJECT4;
 input Tile_X0Y5_UIO_OUT_TT_PROJECT5;
 input Tile_X0Y5_UIO_OUT_TT_PROJECT6;
 input Tile_X0Y5_UIO_OUT_TT_PROJECT7;
 output Tile_X0Y5_UI_IN_TT_PROJECT0;
 output Tile_X0Y5_UI_IN_TT_PROJECT1;
 output Tile_X0Y5_UI_IN_TT_PROJECT2;
 output Tile_X0Y5_UI_IN_TT_PROJECT3;
 output Tile_X0Y5_UI_IN_TT_PROJECT4;
 output Tile_X0Y5_UI_IN_TT_PROJECT5;
 output Tile_X0Y5_UI_IN_TT_PROJECT6;
 output Tile_X0Y5_UI_IN_TT_PROJECT7;
 input Tile_X0Y5_UO_OUT_TT_PROJECT0;
 input Tile_X0Y5_UO_OUT_TT_PROJECT1;
 input Tile_X0Y5_UO_OUT_TT_PROJECT2;
 input Tile_X0Y5_UO_OUT_TT_PROJECT3;
 input Tile_X0Y5_UO_OUT_TT_PROJECT4;
 input Tile_X0Y5_UO_OUT_TT_PROJECT5;
 input Tile_X0Y5_UO_OUT_TT_PROJECT6;
 input Tile_X0Y5_UO_OUT_TT_PROJECT7;
 output Tile_X0Y6_CLK_TT_PROJECT;
 output Tile_X0Y6_ENA_TT_PROJECT;
 output Tile_X0Y6_RST_N_TT_PROJECT;
 output Tile_X0Y6_UIO_IN_TT_PROJECT0;
 output Tile_X0Y6_UIO_IN_TT_PROJECT1;
 output Tile_X0Y6_UIO_IN_TT_PROJECT2;
 output Tile_X0Y6_UIO_IN_TT_PROJECT3;
 output Tile_X0Y6_UIO_IN_TT_PROJECT4;
 output Tile_X0Y6_UIO_IN_TT_PROJECT5;
 output Tile_X0Y6_UIO_IN_TT_PROJECT6;
 output Tile_X0Y6_UIO_IN_TT_PROJECT7;
 input Tile_X0Y6_UIO_OE_TT_PROJECT0;
 input Tile_X0Y6_UIO_OE_TT_PROJECT1;
 input Tile_X0Y6_UIO_OE_TT_PROJECT2;
 input Tile_X0Y6_UIO_OE_TT_PROJECT3;
 input Tile_X0Y6_UIO_OE_TT_PROJECT4;
 input Tile_X0Y6_UIO_OE_TT_PROJECT5;
 input Tile_X0Y6_UIO_OE_TT_PROJECT6;
 input Tile_X0Y6_UIO_OE_TT_PROJECT7;
 input Tile_X0Y6_UIO_OUT_TT_PROJECT0;
 input Tile_X0Y6_UIO_OUT_TT_PROJECT1;
 input Tile_X0Y6_UIO_OUT_TT_PROJECT2;
 input Tile_X0Y6_UIO_OUT_TT_PROJECT3;
 input Tile_X0Y6_UIO_OUT_TT_PROJECT4;
 input Tile_X0Y6_UIO_OUT_TT_PROJECT5;
 input Tile_X0Y6_UIO_OUT_TT_PROJECT6;
 input Tile_X0Y6_UIO_OUT_TT_PROJECT7;
 output Tile_X0Y6_UI_IN_TT_PROJECT0;
 output Tile_X0Y6_UI_IN_TT_PROJECT1;
 output Tile_X0Y6_UI_IN_TT_PROJECT2;
 output Tile_X0Y6_UI_IN_TT_PROJECT3;
 output Tile_X0Y6_UI_IN_TT_PROJECT4;
 output Tile_X0Y6_UI_IN_TT_PROJECT5;
 output Tile_X0Y6_UI_IN_TT_PROJECT6;
 output Tile_X0Y6_UI_IN_TT_PROJECT7;
 input Tile_X0Y6_UO_OUT_TT_PROJECT0;
 input Tile_X0Y6_UO_OUT_TT_PROJECT1;
 input Tile_X0Y6_UO_OUT_TT_PROJECT2;
 input Tile_X0Y6_UO_OUT_TT_PROJECT3;
 input Tile_X0Y6_UO_OUT_TT_PROJECT4;
 input Tile_X0Y6_UO_OUT_TT_PROJECT5;
 input Tile_X0Y6_UO_OUT_TT_PROJECT6;
 input Tile_X0Y6_UO_OUT_TT_PROJECT7;
 output Tile_X0Y7_CLK_TT_PROJECT;
 output Tile_X0Y7_ENA_TT_PROJECT;
 output Tile_X0Y7_RST_N_TT_PROJECT;
 output Tile_X0Y7_UIO_IN_TT_PROJECT0;
 output Tile_X0Y7_UIO_IN_TT_PROJECT1;
 output Tile_X0Y7_UIO_IN_TT_PROJECT2;
 output Tile_X0Y7_UIO_IN_TT_PROJECT3;
 output Tile_X0Y7_UIO_IN_TT_PROJECT4;
 output Tile_X0Y7_UIO_IN_TT_PROJECT5;
 output Tile_X0Y7_UIO_IN_TT_PROJECT6;
 output Tile_X0Y7_UIO_IN_TT_PROJECT7;
 input Tile_X0Y7_UIO_OE_TT_PROJECT0;
 input Tile_X0Y7_UIO_OE_TT_PROJECT1;
 input Tile_X0Y7_UIO_OE_TT_PROJECT2;
 input Tile_X0Y7_UIO_OE_TT_PROJECT3;
 input Tile_X0Y7_UIO_OE_TT_PROJECT4;
 input Tile_X0Y7_UIO_OE_TT_PROJECT5;
 input Tile_X0Y7_UIO_OE_TT_PROJECT6;
 input Tile_X0Y7_UIO_OE_TT_PROJECT7;
 input Tile_X0Y7_UIO_OUT_TT_PROJECT0;
 input Tile_X0Y7_UIO_OUT_TT_PROJECT1;
 input Tile_X0Y7_UIO_OUT_TT_PROJECT2;
 input Tile_X0Y7_UIO_OUT_TT_PROJECT3;
 input Tile_X0Y7_UIO_OUT_TT_PROJECT4;
 input Tile_X0Y7_UIO_OUT_TT_PROJECT5;
 input Tile_X0Y7_UIO_OUT_TT_PROJECT6;
 input Tile_X0Y7_UIO_OUT_TT_PROJECT7;
 output Tile_X0Y7_UI_IN_TT_PROJECT0;
 output Tile_X0Y7_UI_IN_TT_PROJECT1;
 output Tile_X0Y7_UI_IN_TT_PROJECT2;
 output Tile_X0Y7_UI_IN_TT_PROJECT3;
 output Tile_X0Y7_UI_IN_TT_PROJECT4;
 output Tile_X0Y7_UI_IN_TT_PROJECT5;
 output Tile_X0Y7_UI_IN_TT_PROJECT6;
 output Tile_X0Y7_UI_IN_TT_PROJECT7;
 input Tile_X0Y7_UO_OUT_TT_PROJECT0;
 input Tile_X0Y7_UO_OUT_TT_PROJECT1;
 input Tile_X0Y7_UO_OUT_TT_PROJECT2;
 input Tile_X0Y7_UO_OUT_TT_PROJECT3;
 input Tile_X0Y7_UO_OUT_TT_PROJECT4;
 input Tile_X0Y7_UO_OUT_TT_PROJECT5;
 input Tile_X0Y7_UO_OUT_TT_PROJECT6;
 input Tile_X0Y7_UO_OUT_TT_PROJECT7;
 output Tile_X0Y8_CLK_TT_PROJECT;
 output Tile_X0Y8_ENA_TT_PROJECT;
 output Tile_X0Y8_RST_N_TT_PROJECT;
 output Tile_X0Y8_UIO_IN_TT_PROJECT0;
 output Tile_X0Y8_UIO_IN_TT_PROJECT1;
 output Tile_X0Y8_UIO_IN_TT_PROJECT2;
 output Tile_X0Y8_UIO_IN_TT_PROJECT3;
 output Tile_X0Y8_UIO_IN_TT_PROJECT4;
 output Tile_X0Y8_UIO_IN_TT_PROJECT5;
 output Tile_X0Y8_UIO_IN_TT_PROJECT6;
 output Tile_X0Y8_UIO_IN_TT_PROJECT7;
 input Tile_X0Y8_UIO_OE_TT_PROJECT0;
 input Tile_X0Y8_UIO_OE_TT_PROJECT1;
 input Tile_X0Y8_UIO_OE_TT_PROJECT2;
 input Tile_X0Y8_UIO_OE_TT_PROJECT3;
 input Tile_X0Y8_UIO_OE_TT_PROJECT4;
 input Tile_X0Y8_UIO_OE_TT_PROJECT5;
 input Tile_X0Y8_UIO_OE_TT_PROJECT6;
 input Tile_X0Y8_UIO_OE_TT_PROJECT7;
 input Tile_X0Y8_UIO_OUT_TT_PROJECT0;
 input Tile_X0Y8_UIO_OUT_TT_PROJECT1;
 input Tile_X0Y8_UIO_OUT_TT_PROJECT2;
 input Tile_X0Y8_UIO_OUT_TT_PROJECT3;
 input Tile_X0Y8_UIO_OUT_TT_PROJECT4;
 input Tile_X0Y8_UIO_OUT_TT_PROJECT5;
 input Tile_X0Y8_UIO_OUT_TT_PROJECT6;
 input Tile_X0Y8_UIO_OUT_TT_PROJECT7;
 output Tile_X0Y8_UI_IN_TT_PROJECT0;
 output Tile_X0Y8_UI_IN_TT_PROJECT1;
 output Tile_X0Y8_UI_IN_TT_PROJECT2;
 output Tile_X0Y8_UI_IN_TT_PROJECT3;
 output Tile_X0Y8_UI_IN_TT_PROJECT4;
 output Tile_X0Y8_UI_IN_TT_PROJECT5;
 output Tile_X0Y8_UI_IN_TT_PROJECT6;
 output Tile_X0Y8_UI_IN_TT_PROJECT7;
 input Tile_X0Y8_UO_OUT_TT_PROJECT0;
 input Tile_X0Y8_UO_OUT_TT_PROJECT1;
 input Tile_X0Y8_UO_OUT_TT_PROJECT2;
 input Tile_X0Y8_UO_OUT_TT_PROJECT3;
 input Tile_X0Y8_UO_OUT_TT_PROJECT4;
 input Tile_X0Y8_UO_OUT_TT_PROJECT5;
 input Tile_X0Y8_UO_OUT_TT_PROJECT6;
 input Tile_X0Y8_UO_OUT_TT_PROJECT7;
 output Tile_X1Y0_A_I_top;
 input Tile_X1Y0_A_O_top;
 output Tile_X1Y0_A_T_top;
 output Tile_X1Y0_B_I_top;
 input Tile_X1Y0_B_O_top;
 output Tile_X1Y0_B_T_top;
 output Tile_X1Y0_C_I_top;
 input Tile_X1Y0_C_O_top;
 output Tile_X1Y0_C_T_top;
 output Tile_X1Y0_D_I_top;
 input Tile_X1Y0_D_O_top;
 output Tile_X1Y0_D_T_top;
 output Tile_X1Y9_A_I_top;
 input Tile_X1Y9_A_O_top;
 output Tile_X1Y9_A_T_top;
 output Tile_X1Y9_B_I_top;
 input Tile_X1Y9_B_O_top;
 output Tile_X1Y9_B_T_top;
 output Tile_X1Y9_C_I_top;
 input Tile_X1Y9_C_O_top;
 output Tile_X1Y9_C_T_top;
 output Tile_X1Y9_D_I_top;
 input Tile_X1Y9_D_O_top;
 output Tile_X1Y9_D_T_top;
 output Tile_X2Y0_A_I_top;
 input Tile_X2Y0_A_O_top;
 output Tile_X2Y0_A_T_top;
 output Tile_X2Y0_B_I_top;
 input Tile_X2Y0_B_O_top;
 output Tile_X2Y0_B_T_top;
 output Tile_X2Y0_C_I_top;
 input Tile_X2Y0_C_O_top;
 output Tile_X2Y0_C_T_top;
 output Tile_X2Y0_D_I_top;
 input Tile_X2Y0_D_O_top;
 output Tile_X2Y0_D_T_top;
 output Tile_X2Y9_A_I_top;
 input Tile_X2Y9_A_O_top;
 output Tile_X2Y9_A_T_top;
 output Tile_X2Y9_B_I_top;
 input Tile_X2Y9_B_O_top;
 output Tile_X2Y9_B_T_top;
 output Tile_X2Y9_C_I_top;
 input Tile_X2Y9_C_O_top;
 output Tile_X2Y9_C_T_top;
 output Tile_X2Y9_D_I_top;
 input Tile_X2Y9_D_O_top;
 output Tile_X2Y9_D_T_top;
 output Tile_X3Y0_A_I_top;
 input Tile_X3Y0_A_O_top;
 output Tile_X3Y0_A_T_top;
 output Tile_X3Y0_B_I_top;
 input Tile_X3Y0_B_O_top;
 output Tile_X3Y0_B_T_top;
 output Tile_X3Y0_C_I_top;
 input Tile_X3Y0_C_O_top;
 output Tile_X3Y0_C_T_top;
 output Tile_X3Y0_D_I_top;
 input Tile_X3Y0_D_O_top;
 output Tile_X3Y0_D_T_top;
 output Tile_X3Y9_A_I_top;
 input Tile_X3Y9_A_O_top;
 output Tile_X3Y9_A_T_top;
 output Tile_X3Y9_B_I_top;
 input Tile_X3Y9_B_O_top;
 output Tile_X3Y9_B_T_top;
 output Tile_X3Y9_C_I_top;
 input Tile_X3Y9_C_O_top;
 output Tile_X3Y9_C_T_top;
 output Tile_X3Y9_D_I_top;
 input Tile_X3Y9_D_O_top;
 output Tile_X3Y9_D_T_top;
 output Tile_X4Y0_A_I_top;
 input Tile_X4Y0_A_O_top;
 output Tile_X4Y0_A_T_top;
 output Tile_X4Y0_B_I_top;
 input Tile_X4Y0_B_O_top;
 output Tile_X4Y0_B_T_top;
 output Tile_X4Y0_C_I_top;
 input Tile_X4Y0_C_O_top;
 output Tile_X4Y0_C_T_top;
 output Tile_X4Y0_D_I_top;
 input Tile_X4Y0_D_O_top;
 output Tile_X4Y0_D_T_top;
 output Tile_X4Y9_A_I_top;
 input Tile_X4Y9_A_O_top;
 output Tile_X4Y9_A_T_top;
 output Tile_X4Y9_B_I_top;
 input Tile_X4Y9_B_O_top;
 output Tile_X4Y9_B_T_top;
 output Tile_X4Y9_C_I_top;
 input Tile_X4Y9_C_O_top;
 output Tile_X4Y9_C_T_top;
 output Tile_X4Y9_D_I_top;
 input Tile_X4Y9_D_O_top;
 output Tile_X4Y9_D_T_top;
 output Tile_X5Y2_ADDR_SRAM0;
 output Tile_X5Y2_ADDR_SRAM1;
 output Tile_X5Y2_ADDR_SRAM2;
 output Tile_X5Y2_ADDR_SRAM3;
 output Tile_X5Y2_ADDR_SRAM4;
 output Tile_X5Y2_ADDR_SRAM5;
 output Tile_X5Y2_ADDR_SRAM6;
 output Tile_X5Y2_ADDR_SRAM7;
 output Tile_X5Y2_ADDR_SRAM8;
 output Tile_X5Y2_ADDR_SRAM9;
 output Tile_X5Y2_BM_SRAM0;
 output Tile_X5Y2_BM_SRAM1;
 output Tile_X5Y2_BM_SRAM10;
 output Tile_X5Y2_BM_SRAM11;
 output Tile_X5Y2_BM_SRAM12;
 output Tile_X5Y2_BM_SRAM13;
 output Tile_X5Y2_BM_SRAM14;
 output Tile_X5Y2_BM_SRAM15;
 output Tile_X5Y2_BM_SRAM16;
 output Tile_X5Y2_BM_SRAM17;
 output Tile_X5Y2_BM_SRAM18;
 output Tile_X5Y2_BM_SRAM19;
 output Tile_X5Y2_BM_SRAM2;
 output Tile_X5Y2_BM_SRAM20;
 output Tile_X5Y2_BM_SRAM21;
 output Tile_X5Y2_BM_SRAM22;
 output Tile_X5Y2_BM_SRAM23;
 output Tile_X5Y2_BM_SRAM24;
 output Tile_X5Y2_BM_SRAM25;
 output Tile_X5Y2_BM_SRAM26;
 output Tile_X5Y2_BM_SRAM27;
 output Tile_X5Y2_BM_SRAM28;
 output Tile_X5Y2_BM_SRAM29;
 output Tile_X5Y2_BM_SRAM3;
 output Tile_X5Y2_BM_SRAM30;
 output Tile_X5Y2_BM_SRAM31;
 output Tile_X5Y2_BM_SRAM4;
 output Tile_X5Y2_BM_SRAM5;
 output Tile_X5Y2_BM_SRAM6;
 output Tile_X5Y2_BM_SRAM7;
 output Tile_X5Y2_BM_SRAM8;
 output Tile_X5Y2_BM_SRAM9;
 output Tile_X5Y2_CLK_SRAM;
 input Tile_X5Y2_CONFIGURED_top;
 output Tile_X5Y2_DIN_SRAM0;
 output Tile_X5Y2_DIN_SRAM1;
 output Tile_X5Y2_DIN_SRAM10;
 output Tile_X5Y2_DIN_SRAM11;
 output Tile_X5Y2_DIN_SRAM12;
 output Tile_X5Y2_DIN_SRAM13;
 output Tile_X5Y2_DIN_SRAM14;
 output Tile_X5Y2_DIN_SRAM15;
 output Tile_X5Y2_DIN_SRAM16;
 output Tile_X5Y2_DIN_SRAM17;
 output Tile_X5Y2_DIN_SRAM18;
 output Tile_X5Y2_DIN_SRAM19;
 output Tile_X5Y2_DIN_SRAM2;
 output Tile_X5Y2_DIN_SRAM20;
 output Tile_X5Y2_DIN_SRAM21;
 output Tile_X5Y2_DIN_SRAM22;
 output Tile_X5Y2_DIN_SRAM23;
 output Tile_X5Y2_DIN_SRAM24;
 output Tile_X5Y2_DIN_SRAM25;
 output Tile_X5Y2_DIN_SRAM26;
 output Tile_X5Y2_DIN_SRAM27;
 output Tile_X5Y2_DIN_SRAM28;
 output Tile_X5Y2_DIN_SRAM29;
 output Tile_X5Y2_DIN_SRAM3;
 output Tile_X5Y2_DIN_SRAM30;
 output Tile_X5Y2_DIN_SRAM31;
 output Tile_X5Y2_DIN_SRAM4;
 output Tile_X5Y2_DIN_SRAM5;
 output Tile_X5Y2_DIN_SRAM6;
 output Tile_X5Y2_DIN_SRAM7;
 output Tile_X5Y2_DIN_SRAM8;
 output Tile_X5Y2_DIN_SRAM9;
 input Tile_X5Y2_DOUT_SRAM0;
 input Tile_X5Y2_DOUT_SRAM1;
 input Tile_X5Y2_DOUT_SRAM10;
 input Tile_X5Y2_DOUT_SRAM11;
 input Tile_X5Y2_DOUT_SRAM12;
 input Tile_X5Y2_DOUT_SRAM13;
 input Tile_X5Y2_DOUT_SRAM14;
 input Tile_X5Y2_DOUT_SRAM15;
 input Tile_X5Y2_DOUT_SRAM16;
 input Tile_X5Y2_DOUT_SRAM17;
 input Tile_X5Y2_DOUT_SRAM18;
 input Tile_X5Y2_DOUT_SRAM19;
 input Tile_X5Y2_DOUT_SRAM2;
 input Tile_X5Y2_DOUT_SRAM20;
 input Tile_X5Y2_DOUT_SRAM21;
 input Tile_X5Y2_DOUT_SRAM22;
 input Tile_X5Y2_DOUT_SRAM23;
 input Tile_X5Y2_DOUT_SRAM24;
 input Tile_X5Y2_DOUT_SRAM25;
 input Tile_X5Y2_DOUT_SRAM26;
 input Tile_X5Y2_DOUT_SRAM27;
 input Tile_X5Y2_DOUT_SRAM28;
 input Tile_X5Y2_DOUT_SRAM29;
 input Tile_X5Y2_DOUT_SRAM3;
 input Tile_X5Y2_DOUT_SRAM30;
 input Tile_X5Y2_DOUT_SRAM31;
 input Tile_X5Y2_DOUT_SRAM4;
 input Tile_X5Y2_DOUT_SRAM5;
 input Tile_X5Y2_DOUT_SRAM6;
 input Tile_X5Y2_DOUT_SRAM7;
 input Tile_X5Y2_DOUT_SRAM8;
 input Tile_X5Y2_DOUT_SRAM9;
 output Tile_X5Y2_MEN_SRAM;
 output Tile_X5Y2_REN_SRAM;
 output Tile_X5Y2_TIE_HIGH_SRAM;
 output Tile_X5Y2_TIE_LOW_SRAM;
 output Tile_X5Y2_WEN_SRAM;
 output Tile_X5Y4_CLK_TT_PROJECT;
 output Tile_X5Y4_ENA_TT_PROJECT;
 output Tile_X5Y4_RST_N_TT_PROJECT;
 output Tile_X5Y4_UIO_IN_TT_PROJECT0;
 output Tile_X5Y4_UIO_IN_TT_PROJECT1;
 output Tile_X5Y4_UIO_IN_TT_PROJECT2;
 output Tile_X5Y4_UIO_IN_TT_PROJECT3;
 output Tile_X5Y4_UIO_IN_TT_PROJECT4;
 output Tile_X5Y4_UIO_IN_TT_PROJECT5;
 output Tile_X5Y4_UIO_IN_TT_PROJECT6;
 output Tile_X5Y4_UIO_IN_TT_PROJECT7;
 input Tile_X5Y4_UIO_OE_TT_PROJECT0;
 input Tile_X5Y4_UIO_OE_TT_PROJECT1;
 input Tile_X5Y4_UIO_OE_TT_PROJECT2;
 input Tile_X5Y4_UIO_OE_TT_PROJECT3;
 input Tile_X5Y4_UIO_OE_TT_PROJECT4;
 input Tile_X5Y4_UIO_OE_TT_PROJECT5;
 input Tile_X5Y4_UIO_OE_TT_PROJECT6;
 input Tile_X5Y4_UIO_OE_TT_PROJECT7;
 input Tile_X5Y4_UIO_OUT_TT_PROJECT0;
 input Tile_X5Y4_UIO_OUT_TT_PROJECT1;
 input Tile_X5Y4_UIO_OUT_TT_PROJECT2;
 input Tile_X5Y4_UIO_OUT_TT_PROJECT3;
 input Tile_X5Y4_UIO_OUT_TT_PROJECT4;
 input Tile_X5Y4_UIO_OUT_TT_PROJECT5;
 input Tile_X5Y4_UIO_OUT_TT_PROJECT6;
 input Tile_X5Y4_UIO_OUT_TT_PROJECT7;
 output Tile_X5Y4_UI_IN_TT_PROJECT0;
 output Tile_X5Y4_UI_IN_TT_PROJECT1;
 output Tile_X5Y4_UI_IN_TT_PROJECT2;
 output Tile_X5Y4_UI_IN_TT_PROJECT3;
 output Tile_X5Y4_UI_IN_TT_PROJECT4;
 output Tile_X5Y4_UI_IN_TT_PROJECT5;
 output Tile_X5Y4_UI_IN_TT_PROJECT6;
 output Tile_X5Y4_UI_IN_TT_PROJECT7;
 input Tile_X5Y4_UO_OUT_TT_PROJECT0;
 input Tile_X5Y4_UO_OUT_TT_PROJECT1;
 input Tile_X5Y4_UO_OUT_TT_PROJECT2;
 input Tile_X5Y4_UO_OUT_TT_PROJECT3;
 input Tile_X5Y4_UO_OUT_TT_PROJECT4;
 input Tile_X5Y4_UO_OUT_TT_PROJECT5;
 input Tile_X5Y4_UO_OUT_TT_PROJECT6;
 input Tile_X5Y4_UO_OUT_TT_PROJECT7;
 output Tile_X5Y5_CLK_TT_PROJECT;
 output Tile_X5Y5_ENA_TT_PROJECT;
 output Tile_X5Y5_RST_N_TT_PROJECT;
 output Tile_X5Y5_UIO_IN_TT_PROJECT0;
 output Tile_X5Y5_UIO_IN_TT_PROJECT1;
 output Tile_X5Y5_UIO_IN_TT_PROJECT2;
 output Tile_X5Y5_UIO_IN_TT_PROJECT3;
 output Tile_X5Y5_UIO_IN_TT_PROJECT4;
 output Tile_X5Y5_UIO_IN_TT_PROJECT5;
 output Tile_X5Y5_UIO_IN_TT_PROJECT6;
 output Tile_X5Y5_UIO_IN_TT_PROJECT7;
 input Tile_X5Y5_UIO_OE_TT_PROJECT0;
 input Tile_X5Y5_UIO_OE_TT_PROJECT1;
 input Tile_X5Y5_UIO_OE_TT_PROJECT2;
 input Tile_X5Y5_UIO_OE_TT_PROJECT3;
 input Tile_X5Y5_UIO_OE_TT_PROJECT4;
 input Tile_X5Y5_UIO_OE_TT_PROJECT5;
 input Tile_X5Y5_UIO_OE_TT_PROJECT6;
 input Tile_X5Y5_UIO_OE_TT_PROJECT7;
 input Tile_X5Y5_UIO_OUT_TT_PROJECT0;
 input Tile_X5Y5_UIO_OUT_TT_PROJECT1;
 input Tile_X5Y5_UIO_OUT_TT_PROJECT2;
 input Tile_X5Y5_UIO_OUT_TT_PROJECT3;
 input Tile_X5Y5_UIO_OUT_TT_PROJECT4;
 input Tile_X5Y5_UIO_OUT_TT_PROJECT5;
 input Tile_X5Y5_UIO_OUT_TT_PROJECT6;
 input Tile_X5Y5_UIO_OUT_TT_PROJECT7;
 output Tile_X5Y5_UI_IN_TT_PROJECT0;
 output Tile_X5Y5_UI_IN_TT_PROJECT1;
 output Tile_X5Y5_UI_IN_TT_PROJECT2;
 output Tile_X5Y5_UI_IN_TT_PROJECT3;
 output Tile_X5Y5_UI_IN_TT_PROJECT4;
 output Tile_X5Y5_UI_IN_TT_PROJECT5;
 output Tile_X5Y5_UI_IN_TT_PROJECT6;
 output Tile_X5Y5_UI_IN_TT_PROJECT7;
 input Tile_X5Y5_UO_OUT_TT_PROJECT0;
 input Tile_X5Y5_UO_OUT_TT_PROJECT1;
 input Tile_X5Y5_UO_OUT_TT_PROJECT2;
 input Tile_X5Y5_UO_OUT_TT_PROJECT3;
 input Tile_X5Y5_UO_OUT_TT_PROJECT4;
 input Tile_X5Y5_UO_OUT_TT_PROJECT5;
 input Tile_X5Y5_UO_OUT_TT_PROJECT6;
 input Tile_X5Y5_UO_OUT_TT_PROJECT7;
 output Tile_X5Y6_CLK_TT_PROJECT;
 output Tile_X5Y6_ENA_TT_PROJECT;
 output Tile_X5Y6_RST_N_TT_PROJECT;
 output Tile_X5Y6_UIO_IN_TT_PROJECT0;
 output Tile_X5Y6_UIO_IN_TT_PROJECT1;
 output Tile_X5Y6_UIO_IN_TT_PROJECT2;
 output Tile_X5Y6_UIO_IN_TT_PROJECT3;
 output Tile_X5Y6_UIO_IN_TT_PROJECT4;
 output Tile_X5Y6_UIO_IN_TT_PROJECT5;
 output Tile_X5Y6_UIO_IN_TT_PROJECT6;
 output Tile_X5Y6_UIO_IN_TT_PROJECT7;
 input Tile_X5Y6_UIO_OE_TT_PROJECT0;
 input Tile_X5Y6_UIO_OE_TT_PROJECT1;
 input Tile_X5Y6_UIO_OE_TT_PROJECT2;
 input Tile_X5Y6_UIO_OE_TT_PROJECT3;
 input Tile_X5Y6_UIO_OE_TT_PROJECT4;
 input Tile_X5Y6_UIO_OE_TT_PROJECT5;
 input Tile_X5Y6_UIO_OE_TT_PROJECT6;
 input Tile_X5Y6_UIO_OE_TT_PROJECT7;
 input Tile_X5Y6_UIO_OUT_TT_PROJECT0;
 input Tile_X5Y6_UIO_OUT_TT_PROJECT1;
 input Tile_X5Y6_UIO_OUT_TT_PROJECT2;
 input Tile_X5Y6_UIO_OUT_TT_PROJECT3;
 input Tile_X5Y6_UIO_OUT_TT_PROJECT4;
 input Tile_X5Y6_UIO_OUT_TT_PROJECT5;
 input Tile_X5Y6_UIO_OUT_TT_PROJECT6;
 input Tile_X5Y6_UIO_OUT_TT_PROJECT7;
 output Tile_X5Y6_UI_IN_TT_PROJECT0;
 output Tile_X5Y6_UI_IN_TT_PROJECT1;
 output Tile_X5Y6_UI_IN_TT_PROJECT2;
 output Tile_X5Y6_UI_IN_TT_PROJECT3;
 output Tile_X5Y6_UI_IN_TT_PROJECT4;
 output Tile_X5Y6_UI_IN_TT_PROJECT5;
 output Tile_X5Y6_UI_IN_TT_PROJECT6;
 output Tile_X5Y6_UI_IN_TT_PROJECT7;
 input Tile_X5Y6_UO_OUT_TT_PROJECT0;
 input Tile_X5Y6_UO_OUT_TT_PROJECT1;
 input Tile_X5Y6_UO_OUT_TT_PROJECT2;
 input Tile_X5Y6_UO_OUT_TT_PROJECT3;
 input Tile_X5Y6_UO_OUT_TT_PROJECT4;
 input Tile_X5Y6_UO_OUT_TT_PROJECT5;
 input Tile_X5Y6_UO_OUT_TT_PROJECT6;
 input Tile_X5Y6_UO_OUT_TT_PROJECT7;
 output Tile_X5Y7_CLK_TT_PROJECT;
 output Tile_X5Y7_ENA_TT_PROJECT;
 output Tile_X5Y7_RST_N_TT_PROJECT;
 output Tile_X5Y7_UIO_IN_TT_PROJECT0;
 output Tile_X5Y7_UIO_IN_TT_PROJECT1;
 output Tile_X5Y7_UIO_IN_TT_PROJECT2;
 output Tile_X5Y7_UIO_IN_TT_PROJECT3;
 output Tile_X5Y7_UIO_IN_TT_PROJECT4;
 output Tile_X5Y7_UIO_IN_TT_PROJECT5;
 output Tile_X5Y7_UIO_IN_TT_PROJECT6;
 output Tile_X5Y7_UIO_IN_TT_PROJECT7;
 input Tile_X5Y7_UIO_OE_TT_PROJECT0;
 input Tile_X5Y7_UIO_OE_TT_PROJECT1;
 input Tile_X5Y7_UIO_OE_TT_PROJECT2;
 input Tile_X5Y7_UIO_OE_TT_PROJECT3;
 input Tile_X5Y7_UIO_OE_TT_PROJECT4;
 input Tile_X5Y7_UIO_OE_TT_PROJECT5;
 input Tile_X5Y7_UIO_OE_TT_PROJECT6;
 input Tile_X5Y7_UIO_OE_TT_PROJECT7;
 input Tile_X5Y7_UIO_OUT_TT_PROJECT0;
 input Tile_X5Y7_UIO_OUT_TT_PROJECT1;
 input Tile_X5Y7_UIO_OUT_TT_PROJECT2;
 input Tile_X5Y7_UIO_OUT_TT_PROJECT3;
 input Tile_X5Y7_UIO_OUT_TT_PROJECT4;
 input Tile_X5Y7_UIO_OUT_TT_PROJECT5;
 input Tile_X5Y7_UIO_OUT_TT_PROJECT6;
 input Tile_X5Y7_UIO_OUT_TT_PROJECT7;
 output Tile_X5Y7_UI_IN_TT_PROJECT0;
 output Tile_X5Y7_UI_IN_TT_PROJECT1;
 output Tile_X5Y7_UI_IN_TT_PROJECT2;
 output Tile_X5Y7_UI_IN_TT_PROJECT3;
 output Tile_X5Y7_UI_IN_TT_PROJECT4;
 output Tile_X5Y7_UI_IN_TT_PROJECT5;
 output Tile_X5Y7_UI_IN_TT_PROJECT6;
 output Tile_X5Y7_UI_IN_TT_PROJECT7;
 input Tile_X5Y7_UO_OUT_TT_PROJECT0;
 input Tile_X5Y7_UO_OUT_TT_PROJECT1;
 input Tile_X5Y7_UO_OUT_TT_PROJECT2;
 input Tile_X5Y7_UO_OUT_TT_PROJECT3;
 input Tile_X5Y7_UO_OUT_TT_PROJECT4;
 input Tile_X5Y7_UO_OUT_TT_PROJECT5;
 input Tile_X5Y7_UO_OUT_TT_PROJECT6;
 input Tile_X5Y7_UO_OUT_TT_PROJECT7;
 output Tile_X5Y8_CLK_TT_PROJECT;
 output Tile_X5Y8_ENA_TT_PROJECT;
 output Tile_X5Y8_RST_N_TT_PROJECT;
 output Tile_X5Y8_UIO_IN_TT_PROJECT0;
 output Tile_X5Y8_UIO_IN_TT_PROJECT1;
 output Tile_X5Y8_UIO_IN_TT_PROJECT2;
 output Tile_X5Y8_UIO_IN_TT_PROJECT3;
 output Tile_X5Y8_UIO_IN_TT_PROJECT4;
 output Tile_X5Y8_UIO_IN_TT_PROJECT5;
 output Tile_X5Y8_UIO_IN_TT_PROJECT6;
 output Tile_X5Y8_UIO_IN_TT_PROJECT7;
 input Tile_X5Y8_UIO_OE_TT_PROJECT0;
 input Tile_X5Y8_UIO_OE_TT_PROJECT1;
 input Tile_X5Y8_UIO_OE_TT_PROJECT2;
 input Tile_X5Y8_UIO_OE_TT_PROJECT3;
 input Tile_X5Y8_UIO_OE_TT_PROJECT4;
 input Tile_X5Y8_UIO_OE_TT_PROJECT5;
 input Tile_X5Y8_UIO_OE_TT_PROJECT6;
 input Tile_X5Y8_UIO_OE_TT_PROJECT7;
 input Tile_X5Y8_UIO_OUT_TT_PROJECT0;
 input Tile_X5Y8_UIO_OUT_TT_PROJECT1;
 input Tile_X5Y8_UIO_OUT_TT_PROJECT2;
 input Tile_X5Y8_UIO_OUT_TT_PROJECT3;
 input Tile_X5Y8_UIO_OUT_TT_PROJECT4;
 input Tile_X5Y8_UIO_OUT_TT_PROJECT5;
 input Tile_X5Y8_UIO_OUT_TT_PROJECT6;
 input Tile_X5Y8_UIO_OUT_TT_PROJECT7;
 output Tile_X5Y8_UI_IN_TT_PROJECT0;
 output Tile_X5Y8_UI_IN_TT_PROJECT1;
 output Tile_X5Y8_UI_IN_TT_PROJECT2;
 output Tile_X5Y8_UI_IN_TT_PROJECT3;
 output Tile_X5Y8_UI_IN_TT_PROJECT4;
 output Tile_X5Y8_UI_IN_TT_PROJECT5;
 output Tile_X5Y8_UI_IN_TT_PROJECT6;
 output Tile_X5Y8_UI_IN_TT_PROJECT7;
 input Tile_X5Y8_UO_OUT_TT_PROJECT0;
 input Tile_X5Y8_UO_OUT_TT_PROJECT1;
 input Tile_X5Y8_UO_OUT_TT_PROJECT2;
 input Tile_X5Y8_UO_OUT_TT_PROJECT3;
 input Tile_X5Y8_UO_OUT_TT_PROJECT4;
 input Tile_X5Y8_UO_OUT_TT_PROJECT5;
 input Tile_X5Y8_UO_OUT_TT_PROJECT6;
 input Tile_X5Y8_UO_OUT_TT_PROJECT7;
 input UserCLK;
 inout VPWR;
 inout VGND;
 input [319:0] FrameData;
 input [119:0] FrameStrobe;

 wire \Tile_X0Y0_FrameData_O[0] ;
 wire \Tile_X0Y0_FrameData_O[10] ;
 wire \Tile_X0Y0_FrameData_O[11] ;
 wire \Tile_X0Y0_FrameData_O[12] ;
 wire \Tile_X0Y0_FrameData_O[13] ;
 wire \Tile_X0Y0_FrameData_O[14] ;
 wire \Tile_X0Y0_FrameData_O[15] ;
 wire \Tile_X0Y0_FrameData_O[16] ;
 wire \Tile_X0Y0_FrameData_O[17] ;
 wire \Tile_X0Y0_FrameData_O[18] ;
 wire \Tile_X0Y0_FrameData_O[19] ;
 wire \Tile_X0Y0_FrameData_O[1] ;
 wire \Tile_X0Y0_FrameData_O[20] ;
 wire \Tile_X0Y0_FrameData_O[21] ;
 wire \Tile_X0Y0_FrameData_O[22] ;
 wire \Tile_X0Y0_FrameData_O[23] ;
 wire \Tile_X0Y0_FrameData_O[24] ;
 wire \Tile_X0Y0_FrameData_O[25] ;
 wire \Tile_X0Y0_FrameData_O[26] ;
 wire \Tile_X0Y0_FrameData_O[27] ;
 wire \Tile_X0Y0_FrameData_O[28] ;
 wire \Tile_X0Y0_FrameData_O[29] ;
 wire \Tile_X0Y0_FrameData_O[2] ;
 wire \Tile_X0Y0_FrameData_O[30] ;
 wire \Tile_X0Y0_FrameData_O[31] ;
 wire \Tile_X0Y0_FrameData_O[3] ;
 wire \Tile_X0Y0_FrameData_O[4] ;
 wire \Tile_X0Y0_FrameData_O[5] ;
 wire \Tile_X0Y0_FrameData_O[6] ;
 wire \Tile_X0Y0_FrameData_O[7] ;
 wire \Tile_X0Y0_FrameData_O[8] ;
 wire \Tile_X0Y0_FrameData_O[9] ;
 wire \Tile_X0Y0_FrameStrobe_O[0] ;
 wire \Tile_X0Y0_FrameStrobe_O[10] ;
 wire \Tile_X0Y0_FrameStrobe_O[11] ;
 wire \Tile_X0Y0_FrameStrobe_O[12] ;
 wire \Tile_X0Y0_FrameStrobe_O[13] ;
 wire \Tile_X0Y0_FrameStrobe_O[14] ;
 wire \Tile_X0Y0_FrameStrobe_O[15] ;
 wire \Tile_X0Y0_FrameStrobe_O[16] ;
 wire \Tile_X0Y0_FrameStrobe_O[17] ;
 wire \Tile_X0Y0_FrameStrobe_O[18] ;
 wire \Tile_X0Y0_FrameStrobe_O[19] ;
 wire \Tile_X0Y0_FrameStrobe_O[1] ;
 wire \Tile_X0Y0_FrameStrobe_O[2] ;
 wire \Tile_X0Y0_FrameStrobe_O[3] ;
 wire \Tile_X0Y0_FrameStrobe_O[4] ;
 wire \Tile_X0Y0_FrameStrobe_O[5] ;
 wire \Tile_X0Y0_FrameStrobe_O[6] ;
 wire \Tile_X0Y0_FrameStrobe_O[7] ;
 wire \Tile_X0Y0_FrameStrobe_O[8] ;
 wire \Tile_X0Y0_FrameStrobe_O[9] ;
 wire \Tile_X0Y0_S1BEG[0] ;
 wire \Tile_X0Y0_S1BEG[1] ;
 wire \Tile_X0Y0_S1BEG[2] ;
 wire \Tile_X0Y0_S1BEG[3] ;
 wire \Tile_X0Y0_S2BEG[0] ;
 wire \Tile_X0Y0_S2BEG[1] ;
 wire \Tile_X0Y0_S2BEG[2] ;
 wire \Tile_X0Y0_S2BEG[3] ;
 wire \Tile_X0Y0_S2BEG[4] ;
 wire \Tile_X0Y0_S2BEG[5] ;
 wire \Tile_X0Y0_S2BEG[6] ;
 wire \Tile_X0Y0_S2BEG[7] ;
 wire \Tile_X0Y0_S2BEGb[0] ;
 wire \Tile_X0Y0_S2BEGb[1] ;
 wire \Tile_X0Y0_S2BEGb[2] ;
 wire \Tile_X0Y0_S2BEGb[3] ;
 wire \Tile_X0Y0_S2BEGb[4] ;
 wire \Tile_X0Y0_S2BEGb[5] ;
 wire \Tile_X0Y0_S2BEGb[6] ;
 wire \Tile_X0Y0_S2BEGb[7] ;
 wire \Tile_X0Y0_S4BEG[0] ;
 wire \Tile_X0Y0_S4BEG[10] ;
 wire \Tile_X0Y0_S4BEG[11] ;
 wire \Tile_X0Y0_S4BEG[12] ;
 wire \Tile_X0Y0_S4BEG[13] ;
 wire \Tile_X0Y0_S4BEG[14] ;
 wire \Tile_X0Y0_S4BEG[15] ;
 wire \Tile_X0Y0_S4BEG[1] ;
 wire \Tile_X0Y0_S4BEG[2] ;
 wire \Tile_X0Y0_S4BEG[3] ;
 wire \Tile_X0Y0_S4BEG[4] ;
 wire \Tile_X0Y0_S4BEG[5] ;
 wire \Tile_X0Y0_S4BEG[6] ;
 wire \Tile_X0Y0_S4BEG[7] ;
 wire \Tile_X0Y0_S4BEG[8] ;
 wire \Tile_X0Y0_S4BEG[9] ;
 wire Tile_X0Y0_UserCLKo;
 wire \Tile_X0Y1_E1BEG[0] ;
 wire \Tile_X0Y1_E1BEG[1] ;
 wire \Tile_X0Y1_E1BEG[2] ;
 wire \Tile_X0Y1_E1BEG[3] ;
 wire \Tile_X0Y1_E2BEG[0] ;
 wire \Tile_X0Y1_E2BEG[1] ;
 wire \Tile_X0Y1_E2BEG[2] ;
 wire \Tile_X0Y1_E2BEG[3] ;
 wire \Tile_X0Y1_E2BEG[4] ;
 wire \Tile_X0Y1_E2BEG[5] ;
 wire \Tile_X0Y1_E2BEG[6] ;
 wire \Tile_X0Y1_E2BEG[7] ;
 wire \Tile_X0Y1_E2BEGb[0] ;
 wire \Tile_X0Y1_E2BEGb[1] ;
 wire \Tile_X0Y1_E2BEGb[2] ;
 wire \Tile_X0Y1_E2BEGb[3] ;
 wire \Tile_X0Y1_E2BEGb[4] ;
 wire \Tile_X0Y1_E2BEGb[5] ;
 wire \Tile_X0Y1_E2BEGb[6] ;
 wire \Tile_X0Y1_E2BEGb[7] ;
 wire \Tile_X0Y1_E6BEG[0] ;
 wire \Tile_X0Y1_E6BEG[10] ;
 wire \Tile_X0Y1_E6BEG[11] ;
 wire \Tile_X0Y1_E6BEG[1] ;
 wire \Tile_X0Y1_E6BEG[2] ;
 wire \Tile_X0Y1_E6BEG[3] ;
 wire \Tile_X0Y1_E6BEG[4] ;
 wire \Tile_X0Y1_E6BEG[5] ;
 wire \Tile_X0Y1_E6BEG[6] ;
 wire \Tile_X0Y1_E6BEG[7] ;
 wire \Tile_X0Y1_E6BEG[8] ;
 wire \Tile_X0Y1_E6BEG[9] ;
 wire \Tile_X0Y1_EE4BEG[0] ;
 wire \Tile_X0Y1_EE4BEG[10] ;
 wire \Tile_X0Y1_EE4BEG[11] ;
 wire \Tile_X0Y1_EE4BEG[12] ;
 wire \Tile_X0Y1_EE4BEG[13] ;
 wire \Tile_X0Y1_EE4BEG[14] ;
 wire \Tile_X0Y1_EE4BEG[15] ;
 wire \Tile_X0Y1_EE4BEG[1] ;
 wire \Tile_X0Y1_EE4BEG[2] ;
 wire \Tile_X0Y1_EE4BEG[3] ;
 wire \Tile_X0Y1_EE4BEG[4] ;
 wire \Tile_X0Y1_EE4BEG[5] ;
 wire \Tile_X0Y1_EE4BEG[6] ;
 wire \Tile_X0Y1_EE4BEG[7] ;
 wire \Tile_X0Y1_EE4BEG[8] ;
 wire \Tile_X0Y1_EE4BEG[9] ;
 wire \Tile_X0Y1_FrameData_O[0] ;
 wire \Tile_X0Y1_FrameData_O[10] ;
 wire \Tile_X0Y1_FrameData_O[11] ;
 wire \Tile_X0Y1_FrameData_O[12] ;
 wire \Tile_X0Y1_FrameData_O[13] ;
 wire \Tile_X0Y1_FrameData_O[14] ;
 wire \Tile_X0Y1_FrameData_O[15] ;
 wire \Tile_X0Y1_FrameData_O[16] ;
 wire \Tile_X0Y1_FrameData_O[17] ;
 wire \Tile_X0Y1_FrameData_O[18] ;
 wire \Tile_X0Y1_FrameData_O[19] ;
 wire \Tile_X0Y1_FrameData_O[1] ;
 wire \Tile_X0Y1_FrameData_O[20] ;
 wire \Tile_X0Y1_FrameData_O[21] ;
 wire \Tile_X0Y1_FrameData_O[22] ;
 wire \Tile_X0Y1_FrameData_O[23] ;
 wire \Tile_X0Y1_FrameData_O[24] ;
 wire \Tile_X0Y1_FrameData_O[25] ;
 wire \Tile_X0Y1_FrameData_O[26] ;
 wire \Tile_X0Y1_FrameData_O[27] ;
 wire \Tile_X0Y1_FrameData_O[28] ;
 wire \Tile_X0Y1_FrameData_O[29] ;
 wire \Tile_X0Y1_FrameData_O[2] ;
 wire \Tile_X0Y1_FrameData_O[30] ;
 wire \Tile_X0Y1_FrameData_O[31] ;
 wire \Tile_X0Y1_FrameData_O[3] ;
 wire \Tile_X0Y1_FrameData_O[4] ;
 wire \Tile_X0Y1_FrameData_O[5] ;
 wire \Tile_X0Y1_FrameData_O[6] ;
 wire \Tile_X0Y1_FrameData_O[7] ;
 wire \Tile_X0Y1_FrameData_O[8] ;
 wire \Tile_X0Y1_FrameData_O[9] ;
 wire \Tile_X0Y1_FrameStrobe_O[0] ;
 wire \Tile_X0Y1_FrameStrobe_O[10] ;
 wire \Tile_X0Y1_FrameStrobe_O[11] ;
 wire \Tile_X0Y1_FrameStrobe_O[12] ;
 wire \Tile_X0Y1_FrameStrobe_O[13] ;
 wire \Tile_X0Y1_FrameStrobe_O[14] ;
 wire \Tile_X0Y1_FrameStrobe_O[15] ;
 wire \Tile_X0Y1_FrameStrobe_O[16] ;
 wire \Tile_X0Y1_FrameStrobe_O[17] ;
 wire \Tile_X0Y1_FrameStrobe_O[18] ;
 wire \Tile_X0Y1_FrameStrobe_O[19] ;
 wire \Tile_X0Y1_FrameStrobe_O[1] ;
 wire \Tile_X0Y1_FrameStrobe_O[2] ;
 wire \Tile_X0Y1_FrameStrobe_O[3] ;
 wire \Tile_X0Y1_FrameStrobe_O[4] ;
 wire \Tile_X0Y1_FrameStrobe_O[5] ;
 wire \Tile_X0Y1_FrameStrobe_O[6] ;
 wire \Tile_X0Y1_FrameStrobe_O[7] ;
 wire \Tile_X0Y1_FrameStrobe_O[8] ;
 wire \Tile_X0Y1_FrameStrobe_O[9] ;
 wire \Tile_X0Y1_N1BEG[0] ;
 wire \Tile_X0Y1_N1BEG[1] ;
 wire \Tile_X0Y1_N1BEG[2] ;
 wire \Tile_X0Y1_N1BEG[3] ;
 wire \Tile_X0Y1_N2BEG[0] ;
 wire \Tile_X0Y1_N2BEG[1] ;
 wire \Tile_X0Y1_N2BEG[2] ;
 wire \Tile_X0Y1_N2BEG[3] ;
 wire \Tile_X0Y1_N2BEG[4] ;
 wire \Tile_X0Y1_N2BEG[5] ;
 wire \Tile_X0Y1_N2BEG[6] ;
 wire \Tile_X0Y1_N2BEG[7] ;
 wire \Tile_X0Y1_N2BEGb[0] ;
 wire \Tile_X0Y1_N2BEGb[1] ;
 wire \Tile_X0Y1_N2BEGb[2] ;
 wire \Tile_X0Y1_N2BEGb[3] ;
 wire \Tile_X0Y1_N2BEGb[4] ;
 wire \Tile_X0Y1_N2BEGb[5] ;
 wire \Tile_X0Y1_N2BEGb[6] ;
 wire \Tile_X0Y1_N2BEGb[7] ;
 wire \Tile_X0Y1_N4BEG[0] ;
 wire \Tile_X0Y1_N4BEG[10] ;
 wire \Tile_X0Y1_N4BEG[11] ;
 wire \Tile_X0Y1_N4BEG[12] ;
 wire \Tile_X0Y1_N4BEG[13] ;
 wire \Tile_X0Y1_N4BEG[14] ;
 wire \Tile_X0Y1_N4BEG[15] ;
 wire \Tile_X0Y1_N4BEG[1] ;
 wire \Tile_X0Y1_N4BEG[2] ;
 wire \Tile_X0Y1_N4BEG[3] ;
 wire \Tile_X0Y1_N4BEG[4] ;
 wire \Tile_X0Y1_N4BEG[5] ;
 wire \Tile_X0Y1_N4BEG[6] ;
 wire \Tile_X0Y1_N4BEG[7] ;
 wire \Tile_X0Y1_N4BEG[8] ;
 wire \Tile_X0Y1_N4BEG[9] ;
 wire Tile_X0Y1_UserCLKo;
 wire \Tile_X0Y2_E1BEG[0] ;
 wire \Tile_X0Y2_E1BEG[1] ;
 wire \Tile_X0Y2_E1BEG[2] ;
 wire \Tile_X0Y2_E1BEG[3] ;
 wire \Tile_X0Y2_E2BEG[0] ;
 wire \Tile_X0Y2_E2BEG[1] ;
 wire \Tile_X0Y2_E2BEG[2] ;
 wire \Tile_X0Y2_E2BEG[3] ;
 wire \Tile_X0Y2_E2BEG[4] ;
 wire \Tile_X0Y2_E2BEG[5] ;
 wire \Tile_X0Y2_E2BEG[6] ;
 wire \Tile_X0Y2_E2BEG[7] ;
 wire \Tile_X0Y2_E2BEGb[0] ;
 wire \Tile_X0Y2_E2BEGb[1] ;
 wire \Tile_X0Y2_E2BEGb[2] ;
 wire \Tile_X0Y2_E2BEGb[3] ;
 wire \Tile_X0Y2_E2BEGb[4] ;
 wire \Tile_X0Y2_E2BEGb[5] ;
 wire \Tile_X0Y2_E2BEGb[6] ;
 wire \Tile_X0Y2_E2BEGb[7] ;
 wire \Tile_X0Y2_E6BEG[0] ;
 wire \Tile_X0Y2_E6BEG[10] ;
 wire \Tile_X0Y2_E6BEG[11] ;
 wire \Tile_X0Y2_E6BEG[1] ;
 wire \Tile_X0Y2_E6BEG[2] ;
 wire \Tile_X0Y2_E6BEG[3] ;
 wire \Tile_X0Y2_E6BEG[4] ;
 wire \Tile_X0Y2_E6BEG[5] ;
 wire \Tile_X0Y2_E6BEG[6] ;
 wire \Tile_X0Y2_E6BEG[7] ;
 wire \Tile_X0Y2_E6BEG[8] ;
 wire \Tile_X0Y2_E6BEG[9] ;
 wire \Tile_X0Y2_EE4BEG[0] ;
 wire \Tile_X0Y2_EE4BEG[10] ;
 wire \Tile_X0Y2_EE4BEG[11] ;
 wire \Tile_X0Y2_EE4BEG[12] ;
 wire \Tile_X0Y2_EE4BEG[13] ;
 wire \Tile_X0Y2_EE4BEG[14] ;
 wire \Tile_X0Y2_EE4BEG[15] ;
 wire \Tile_X0Y2_EE4BEG[1] ;
 wire \Tile_X0Y2_EE4BEG[2] ;
 wire \Tile_X0Y2_EE4BEG[3] ;
 wire \Tile_X0Y2_EE4BEG[4] ;
 wire \Tile_X0Y2_EE4BEG[5] ;
 wire \Tile_X0Y2_EE4BEG[6] ;
 wire \Tile_X0Y2_EE4BEG[7] ;
 wire \Tile_X0Y2_EE4BEG[8] ;
 wire \Tile_X0Y2_EE4BEG[9] ;
 wire \Tile_X0Y2_FrameData_O[0] ;
 wire \Tile_X0Y2_FrameData_O[10] ;
 wire \Tile_X0Y2_FrameData_O[11] ;
 wire \Tile_X0Y2_FrameData_O[12] ;
 wire \Tile_X0Y2_FrameData_O[13] ;
 wire \Tile_X0Y2_FrameData_O[14] ;
 wire \Tile_X0Y2_FrameData_O[15] ;
 wire \Tile_X0Y2_FrameData_O[16] ;
 wire \Tile_X0Y2_FrameData_O[17] ;
 wire \Tile_X0Y2_FrameData_O[18] ;
 wire \Tile_X0Y2_FrameData_O[19] ;
 wire \Tile_X0Y2_FrameData_O[1] ;
 wire \Tile_X0Y2_FrameData_O[20] ;
 wire \Tile_X0Y2_FrameData_O[21] ;
 wire \Tile_X0Y2_FrameData_O[22] ;
 wire \Tile_X0Y2_FrameData_O[23] ;
 wire \Tile_X0Y2_FrameData_O[24] ;
 wire \Tile_X0Y2_FrameData_O[25] ;
 wire \Tile_X0Y2_FrameData_O[26] ;
 wire \Tile_X0Y2_FrameData_O[27] ;
 wire \Tile_X0Y2_FrameData_O[28] ;
 wire \Tile_X0Y2_FrameData_O[29] ;
 wire \Tile_X0Y2_FrameData_O[2] ;
 wire \Tile_X0Y2_FrameData_O[30] ;
 wire \Tile_X0Y2_FrameData_O[31] ;
 wire \Tile_X0Y2_FrameData_O[3] ;
 wire \Tile_X0Y2_FrameData_O[4] ;
 wire \Tile_X0Y2_FrameData_O[5] ;
 wire \Tile_X0Y2_FrameData_O[6] ;
 wire \Tile_X0Y2_FrameData_O[7] ;
 wire \Tile_X0Y2_FrameData_O[8] ;
 wire \Tile_X0Y2_FrameData_O[9] ;
 wire \Tile_X0Y2_S1BEG[0] ;
 wire \Tile_X0Y2_S1BEG[1] ;
 wire \Tile_X0Y2_S1BEG[2] ;
 wire \Tile_X0Y2_S1BEG[3] ;
 wire \Tile_X0Y2_S2BEG[0] ;
 wire \Tile_X0Y2_S2BEG[1] ;
 wire \Tile_X0Y2_S2BEG[2] ;
 wire \Tile_X0Y2_S2BEG[3] ;
 wire \Tile_X0Y2_S2BEG[4] ;
 wire \Tile_X0Y2_S2BEG[5] ;
 wire \Tile_X0Y2_S2BEG[6] ;
 wire \Tile_X0Y2_S2BEG[7] ;
 wire \Tile_X0Y2_S2BEGb[0] ;
 wire \Tile_X0Y2_S2BEGb[1] ;
 wire \Tile_X0Y2_S2BEGb[2] ;
 wire \Tile_X0Y2_S2BEGb[3] ;
 wire \Tile_X0Y2_S2BEGb[4] ;
 wire \Tile_X0Y2_S2BEGb[5] ;
 wire \Tile_X0Y2_S2BEGb[6] ;
 wire \Tile_X0Y2_S2BEGb[7] ;
 wire \Tile_X0Y2_S4BEG[0] ;
 wire \Tile_X0Y2_S4BEG[10] ;
 wire \Tile_X0Y2_S4BEG[11] ;
 wire \Tile_X0Y2_S4BEG[12] ;
 wire \Tile_X0Y2_S4BEG[13] ;
 wire \Tile_X0Y2_S4BEG[14] ;
 wire \Tile_X0Y2_S4BEG[15] ;
 wire \Tile_X0Y2_S4BEG[1] ;
 wire \Tile_X0Y2_S4BEG[2] ;
 wire \Tile_X0Y2_S4BEG[3] ;
 wire \Tile_X0Y2_S4BEG[4] ;
 wire \Tile_X0Y2_S4BEG[5] ;
 wire \Tile_X0Y2_S4BEG[6] ;
 wire \Tile_X0Y2_S4BEG[7] ;
 wire \Tile_X0Y2_S4BEG[8] ;
 wire \Tile_X0Y2_S4BEG[9] ;
 wire \Tile_X0Y3_E1BEG[0] ;
 wire \Tile_X0Y3_E1BEG[1] ;
 wire \Tile_X0Y3_E1BEG[2] ;
 wire \Tile_X0Y3_E1BEG[3] ;
 wire \Tile_X0Y3_E2BEG[0] ;
 wire \Tile_X0Y3_E2BEG[1] ;
 wire \Tile_X0Y3_E2BEG[2] ;
 wire \Tile_X0Y3_E2BEG[3] ;
 wire \Tile_X0Y3_E2BEG[4] ;
 wire \Tile_X0Y3_E2BEG[5] ;
 wire \Tile_X0Y3_E2BEG[6] ;
 wire \Tile_X0Y3_E2BEG[7] ;
 wire \Tile_X0Y3_E2BEGb[0] ;
 wire \Tile_X0Y3_E2BEGb[1] ;
 wire \Tile_X0Y3_E2BEGb[2] ;
 wire \Tile_X0Y3_E2BEGb[3] ;
 wire \Tile_X0Y3_E2BEGb[4] ;
 wire \Tile_X0Y3_E2BEGb[5] ;
 wire \Tile_X0Y3_E2BEGb[6] ;
 wire \Tile_X0Y3_E2BEGb[7] ;
 wire \Tile_X0Y3_E6BEG[0] ;
 wire \Tile_X0Y3_E6BEG[10] ;
 wire \Tile_X0Y3_E6BEG[11] ;
 wire \Tile_X0Y3_E6BEG[1] ;
 wire \Tile_X0Y3_E6BEG[2] ;
 wire \Tile_X0Y3_E6BEG[3] ;
 wire \Tile_X0Y3_E6BEG[4] ;
 wire \Tile_X0Y3_E6BEG[5] ;
 wire \Tile_X0Y3_E6BEG[6] ;
 wire \Tile_X0Y3_E6BEG[7] ;
 wire \Tile_X0Y3_E6BEG[8] ;
 wire \Tile_X0Y3_E6BEG[9] ;
 wire \Tile_X0Y3_EE4BEG[0] ;
 wire \Tile_X0Y3_EE4BEG[10] ;
 wire \Tile_X0Y3_EE4BEG[11] ;
 wire \Tile_X0Y3_EE4BEG[12] ;
 wire \Tile_X0Y3_EE4BEG[13] ;
 wire \Tile_X0Y3_EE4BEG[14] ;
 wire \Tile_X0Y3_EE4BEG[15] ;
 wire \Tile_X0Y3_EE4BEG[1] ;
 wire \Tile_X0Y3_EE4BEG[2] ;
 wire \Tile_X0Y3_EE4BEG[3] ;
 wire \Tile_X0Y3_EE4BEG[4] ;
 wire \Tile_X0Y3_EE4BEG[5] ;
 wire \Tile_X0Y3_EE4BEG[6] ;
 wire \Tile_X0Y3_EE4BEG[7] ;
 wire \Tile_X0Y3_EE4BEG[8] ;
 wire \Tile_X0Y3_EE4BEG[9] ;
 wire \Tile_X0Y3_FrameData_O[0] ;
 wire \Tile_X0Y3_FrameData_O[10] ;
 wire \Tile_X0Y3_FrameData_O[11] ;
 wire \Tile_X0Y3_FrameData_O[12] ;
 wire \Tile_X0Y3_FrameData_O[13] ;
 wire \Tile_X0Y3_FrameData_O[14] ;
 wire \Tile_X0Y3_FrameData_O[15] ;
 wire \Tile_X0Y3_FrameData_O[16] ;
 wire \Tile_X0Y3_FrameData_O[17] ;
 wire \Tile_X0Y3_FrameData_O[18] ;
 wire \Tile_X0Y3_FrameData_O[19] ;
 wire \Tile_X0Y3_FrameData_O[1] ;
 wire \Tile_X0Y3_FrameData_O[20] ;
 wire \Tile_X0Y3_FrameData_O[21] ;
 wire \Tile_X0Y3_FrameData_O[22] ;
 wire \Tile_X0Y3_FrameData_O[23] ;
 wire \Tile_X0Y3_FrameData_O[24] ;
 wire \Tile_X0Y3_FrameData_O[25] ;
 wire \Tile_X0Y3_FrameData_O[26] ;
 wire \Tile_X0Y3_FrameData_O[27] ;
 wire \Tile_X0Y3_FrameData_O[28] ;
 wire \Tile_X0Y3_FrameData_O[29] ;
 wire \Tile_X0Y3_FrameData_O[2] ;
 wire \Tile_X0Y3_FrameData_O[30] ;
 wire \Tile_X0Y3_FrameData_O[31] ;
 wire \Tile_X0Y3_FrameData_O[3] ;
 wire \Tile_X0Y3_FrameData_O[4] ;
 wire \Tile_X0Y3_FrameData_O[5] ;
 wire \Tile_X0Y3_FrameData_O[6] ;
 wire \Tile_X0Y3_FrameData_O[7] ;
 wire \Tile_X0Y3_FrameData_O[8] ;
 wire \Tile_X0Y3_FrameData_O[9] ;
 wire \Tile_X0Y3_FrameStrobe_O[0] ;
 wire \Tile_X0Y3_FrameStrobe_O[10] ;
 wire \Tile_X0Y3_FrameStrobe_O[11] ;
 wire \Tile_X0Y3_FrameStrobe_O[12] ;
 wire \Tile_X0Y3_FrameStrobe_O[13] ;
 wire \Tile_X0Y3_FrameStrobe_O[14] ;
 wire \Tile_X0Y3_FrameStrobe_O[15] ;
 wire \Tile_X0Y3_FrameStrobe_O[16] ;
 wire \Tile_X0Y3_FrameStrobe_O[17] ;
 wire \Tile_X0Y3_FrameStrobe_O[18] ;
 wire \Tile_X0Y3_FrameStrobe_O[19] ;
 wire \Tile_X0Y3_FrameStrobe_O[1] ;
 wire \Tile_X0Y3_FrameStrobe_O[2] ;
 wire \Tile_X0Y3_FrameStrobe_O[3] ;
 wire \Tile_X0Y3_FrameStrobe_O[4] ;
 wire \Tile_X0Y3_FrameStrobe_O[5] ;
 wire \Tile_X0Y3_FrameStrobe_O[6] ;
 wire \Tile_X0Y3_FrameStrobe_O[7] ;
 wire \Tile_X0Y3_FrameStrobe_O[8] ;
 wire \Tile_X0Y3_FrameStrobe_O[9] ;
 wire \Tile_X0Y3_N1BEG[0] ;
 wire \Tile_X0Y3_N1BEG[1] ;
 wire \Tile_X0Y3_N1BEG[2] ;
 wire \Tile_X0Y3_N1BEG[3] ;
 wire \Tile_X0Y3_N2BEG[0] ;
 wire \Tile_X0Y3_N2BEG[1] ;
 wire \Tile_X0Y3_N2BEG[2] ;
 wire \Tile_X0Y3_N2BEG[3] ;
 wire \Tile_X0Y3_N2BEG[4] ;
 wire \Tile_X0Y3_N2BEG[5] ;
 wire \Tile_X0Y3_N2BEG[6] ;
 wire \Tile_X0Y3_N2BEG[7] ;
 wire \Tile_X0Y3_N2BEGb[0] ;
 wire \Tile_X0Y3_N2BEGb[1] ;
 wire \Tile_X0Y3_N2BEGb[2] ;
 wire \Tile_X0Y3_N2BEGb[3] ;
 wire \Tile_X0Y3_N2BEGb[4] ;
 wire \Tile_X0Y3_N2BEGb[5] ;
 wire \Tile_X0Y3_N2BEGb[6] ;
 wire \Tile_X0Y3_N2BEGb[7] ;
 wire \Tile_X0Y3_N4BEG[0] ;
 wire \Tile_X0Y3_N4BEG[10] ;
 wire \Tile_X0Y3_N4BEG[11] ;
 wire \Tile_X0Y3_N4BEG[12] ;
 wire \Tile_X0Y3_N4BEG[13] ;
 wire \Tile_X0Y3_N4BEG[14] ;
 wire \Tile_X0Y3_N4BEG[15] ;
 wire \Tile_X0Y3_N4BEG[1] ;
 wire \Tile_X0Y3_N4BEG[2] ;
 wire \Tile_X0Y3_N4BEG[3] ;
 wire \Tile_X0Y3_N4BEG[4] ;
 wire \Tile_X0Y3_N4BEG[5] ;
 wire \Tile_X0Y3_N4BEG[6] ;
 wire \Tile_X0Y3_N4BEG[7] ;
 wire \Tile_X0Y3_N4BEG[8] ;
 wire \Tile_X0Y3_N4BEG[9] ;
 wire \Tile_X0Y3_S1BEG[0] ;
 wire \Tile_X0Y3_S1BEG[1] ;
 wire \Tile_X0Y3_S1BEG[2] ;
 wire \Tile_X0Y3_S1BEG[3] ;
 wire \Tile_X0Y3_S2BEG[0] ;
 wire \Tile_X0Y3_S2BEG[1] ;
 wire \Tile_X0Y3_S2BEG[2] ;
 wire \Tile_X0Y3_S2BEG[3] ;
 wire \Tile_X0Y3_S2BEG[4] ;
 wire \Tile_X0Y3_S2BEG[5] ;
 wire \Tile_X0Y3_S2BEG[6] ;
 wire \Tile_X0Y3_S2BEG[7] ;
 wire \Tile_X0Y3_S2BEGb[0] ;
 wire \Tile_X0Y3_S2BEGb[1] ;
 wire \Tile_X0Y3_S2BEGb[2] ;
 wire \Tile_X0Y3_S2BEGb[3] ;
 wire \Tile_X0Y3_S2BEGb[4] ;
 wire \Tile_X0Y3_S2BEGb[5] ;
 wire \Tile_X0Y3_S2BEGb[6] ;
 wire \Tile_X0Y3_S2BEGb[7] ;
 wire \Tile_X0Y3_S4BEG[0] ;
 wire \Tile_X0Y3_S4BEG[10] ;
 wire \Tile_X0Y3_S4BEG[11] ;
 wire \Tile_X0Y3_S4BEG[12] ;
 wire \Tile_X0Y3_S4BEG[13] ;
 wire \Tile_X0Y3_S4BEG[14] ;
 wire \Tile_X0Y3_S4BEG[15] ;
 wire \Tile_X0Y3_S4BEG[1] ;
 wire \Tile_X0Y3_S4BEG[2] ;
 wire \Tile_X0Y3_S4BEG[3] ;
 wire \Tile_X0Y3_S4BEG[4] ;
 wire \Tile_X0Y3_S4BEG[5] ;
 wire \Tile_X0Y3_S4BEG[6] ;
 wire \Tile_X0Y3_S4BEG[7] ;
 wire \Tile_X0Y3_S4BEG[8] ;
 wire \Tile_X0Y3_S4BEG[9] ;
 wire Tile_X0Y3_UserCLKo;
 wire \Tile_X0Y4_E1BEG[0] ;
 wire \Tile_X0Y4_E1BEG[1] ;
 wire \Tile_X0Y4_E1BEG[2] ;
 wire \Tile_X0Y4_E1BEG[3] ;
 wire \Tile_X0Y4_E2BEG[0] ;
 wire \Tile_X0Y4_E2BEG[1] ;
 wire \Tile_X0Y4_E2BEG[2] ;
 wire \Tile_X0Y4_E2BEG[3] ;
 wire \Tile_X0Y4_E2BEG[4] ;
 wire \Tile_X0Y4_E2BEG[5] ;
 wire \Tile_X0Y4_E2BEG[6] ;
 wire \Tile_X0Y4_E2BEG[7] ;
 wire \Tile_X0Y4_E2BEGb[0] ;
 wire \Tile_X0Y4_E2BEGb[1] ;
 wire \Tile_X0Y4_E2BEGb[2] ;
 wire \Tile_X0Y4_E2BEGb[3] ;
 wire \Tile_X0Y4_E2BEGb[4] ;
 wire \Tile_X0Y4_E2BEGb[5] ;
 wire \Tile_X0Y4_E2BEGb[6] ;
 wire \Tile_X0Y4_E2BEGb[7] ;
 wire \Tile_X0Y4_E6BEG[0] ;
 wire \Tile_X0Y4_E6BEG[10] ;
 wire \Tile_X0Y4_E6BEG[11] ;
 wire \Tile_X0Y4_E6BEG[1] ;
 wire \Tile_X0Y4_E6BEG[2] ;
 wire \Tile_X0Y4_E6BEG[3] ;
 wire \Tile_X0Y4_E6BEG[4] ;
 wire \Tile_X0Y4_E6BEG[5] ;
 wire \Tile_X0Y4_E6BEG[6] ;
 wire \Tile_X0Y4_E6BEG[7] ;
 wire \Tile_X0Y4_E6BEG[8] ;
 wire \Tile_X0Y4_E6BEG[9] ;
 wire \Tile_X0Y4_EE4BEG[0] ;
 wire \Tile_X0Y4_EE4BEG[10] ;
 wire \Tile_X0Y4_EE4BEG[11] ;
 wire \Tile_X0Y4_EE4BEG[12] ;
 wire \Tile_X0Y4_EE4BEG[13] ;
 wire \Tile_X0Y4_EE4BEG[14] ;
 wire \Tile_X0Y4_EE4BEG[15] ;
 wire \Tile_X0Y4_EE4BEG[1] ;
 wire \Tile_X0Y4_EE4BEG[2] ;
 wire \Tile_X0Y4_EE4BEG[3] ;
 wire \Tile_X0Y4_EE4BEG[4] ;
 wire \Tile_X0Y4_EE4BEG[5] ;
 wire \Tile_X0Y4_EE4BEG[6] ;
 wire \Tile_X0Y4_EE4BEG[7] ;
 wire \Tile_X0Y4_EE4BEG[8] ;
 wire \Tile_X0Y4_EE4BEG[9] ;
 wire \Tile_X0Y4_FrameData_O[0] ;
 wire \Tile_X0Y4_FrameData_O[10] ;
 wire \Tile_X0Y4_FrameData_O[11] ;
 wire \Tile_X0Y4_FrameData_O[12] ;
 wire \Tile_X0Y4_FrameData_O[13] ;
 wire \Tile_X0Y4_FrameData_O[14] ;
 wire \Tile_X0Y4_FrameData_O[15] ;
 wire \Tile_X0Y4_FrameData_O[16] ;
 wire \Tile_X0Y4_FrameData_O[17] ;
 wire \Tile_X0Y4_FrameData_O[18] ;
 wire \Tile_X0Y4_FrameData_O[19] ;
 wire \Tile_X0Y4_FrameData_O[1] ;
 wire \Tile_X0Y4_FrameData_O[20] ;
 wire \Tile_X0Y4_FrameData_O[21] ;
 wire \Tile_X0Y4_FrameData_O[22] ;
 wire \Tile_X0Y4_FrameData_O[23] ;
 wire \Tile_X0Y4_FrameData_O[24] ;
 wire \Tile_X0Y4_FrameData_O[25] ;
 wire \Tile_X0Y4_FrameData_O[26] ;
 wire \Tile_X0Y4_FrameData_O[27] ;
 wire \Tile_X0Y4_FrameData_O[28] ;
 wire \Tile_X0Y4_FrameData_O[29] ;
 wire \Tile_X0Y4_FrameData_O[2] ;
 wire \Tile_X0Y4_FrameData_O[30] ;
 wire \Tile_X0Y4_FrameData_O[31] ;
 wire \Tile_X0Y4_FrameData_O[3] ;
 wire \Tile_X0Y4_FrameData_O[4] ;
 wire \Tile_X0Y4_FrameData_O[5] ;
 wire \Tile_X0Y4_FrameData_O[6] ;
 wire \Tile_X0Y4_FrameData_O[7] ;
 wire \Tile_X0Y4_FrameData_O[8] ;
 wire \Tile_X0Y4_FrameData_O[9] ;
 wire \Tile_X0Y4_FrameStrobe_O[0] ;
 wire \Tile_X0Y4_FrameStrobe_O[10] ;
 wire \Tile_X0Y4_FrameStrobe_O[11] ;
 wire \Tile_X0Y4_FrameStrobe_O[12] ;
 wire \Tile_X0Y4_FrameStrobe_O[13] ;
 wire \Tile_X0Y4_FrameStrobe_O[14] ;
 wire \Tile_X0Y4_FrameStrobe_O[15] ;
 wire \Tile_X0Y4_FrameStrobe_O[16] ;
 wire \Tile_X0Y4_FrameStrobe_O[17] ;
 wire \Tile_X0Y4_FrameStrobe_O[18] ;
 wire \Tile_X0Y4_FrameStrobe_O[19] ;
 wire \Tile_X0Y4_FrameStrobe_O[1] ;
 wire \Tile_X0Y4_FrameStrobe_O[2] ;
 wire \Tile_X0Y4_FrameStrobe_O[3] ;
 wire \Tile_X0Y4_FrameStrobe_O[4] ;
 wire \Tile_X0Y4_FrameStrobe_O[5] ;
 wire \Tile_X0Y4_FrameStrobe_O[6] ;
 wire \Tile_X0Y4_FrameStrobe_O[7] ;
 wire \Tile_X0Y4_FrameStrobe_O[8] ;
 wire \Tile_X0Y4_FrameStrobe_O[9] ;
 wire \Tile_X0Y4_N1BEG[0] ;
 wire \Tile_X0Y4_N1BEG[1] ;
 wire \Tile_X0Y4_N1BEG[2] ;
 wire \Tile_X0Y4_N1BEG[3] ;
 wire \Tile_X0Y4_N2BEG[0] ;
 wire \Tile_X0Y4_N2BEG[1] ;
 wire \Tile_X0Y4_N2BEG[2] ;
 wire \Tile_X0Y4_N2BEG[3] ;
 wire \Tile_X0Y4_N2BEG[4] ;
 wire \Tile_X0Y4_N2BEG[5] ;
 wire \Tile_X0Y4_N2BEG[6] ;
 wire \Tile_X0Y4_N2BEG[7] ;
 wire \Tile_X0Y4_N2BEGb[0] ;
 wire \Tile_X0Y4_N2BEGb[1] ;
 wire \Tile_X0Y4_N2BEGb[2] ;
 wire \Tile_X0Y4_N2BEGb[3] ;
 wire \Tile_X0Y4_N2BEGb[4] ;
 wire \Tile_X0Y4_N2BEGb[5] ;
 wire \Tile_X0Y4_N2BEGb[6] ;
 wire \Tile_X0Y4_N2BEGb[7] ;
 wire \Tile_X0Y4_N4BEG[0] ;
 wire \Tile_X0Y4_N4BEG[10] ;
 wire \Tile_X0Y4_N4BEG[11] ;
 wire \Tile_X0Y4_N4BEG[12] ;
 wire \Tile_X0Y4_N4BEG[13] ;
 wire \Tile_X0Y4_N4BEG[14] ;
 wire \Tile_X0Y4_N4BEG[15] ;
 wire \Tile_X0Y4_N4BEG[1] ;
 wire \Tile_X0Y4_N4BEG[2] ;
 wire \Tile_X0Y4_N4BEG[3] ;
 wire \Tile_X0Y4_N4BEG[4] ;
 wire \Tile_X0Y4_N4BEG[5] ;
 wire \Tile_X0Y4_N4BEG[6] ;
 wire \Tile_X0Y4_N4BEG[7] ;
 wire \Tile_X0Y4_N4BEG[8] ;
 wire \Tile_X0Y4_N4BEG[9] ;
 wire \Tile_X0Y4_S1BEG[0] ;
 wire \Tile_X0Y4_S1BEG[1] ;
 wire \Tile_X0Y4_S1BEG[2] ;
 wire \Tile_X0Y4_S1BEG[3] ;
 wire \Tile_X0Y4_S2BEG[0] ;
 wire \Tile_X0Y4_S2BEG[1] ;
 wire \Tile_X0Y4_S2BEG[2] ;
 wire \Tile_X0Y4_S2BEG[3] ;
 wire \Tile_X0Y4_S2BEG[4] ;
 wire \Tile_X0Y4_S2BEG[5] ;
 wire \Tile_X0Y4_S2BEG[6] ;
 wire \Tile_X0Y4_S2BEG[7] ;
 wire \Tile_X0Y4_S2BEGb[0] ;
 wire \Tile_X0Y4_S2BEGb[1] ;
 wire \Tile_X0Y4_S2BEGb[2] ;
 wire \Tile_X0Y4_S2BEGb[3] ;
 wire \Tile_X0Y4_S2BEGb[4] ;
 wire \Tile_X0Y4_S2BEGb[5] ;
 wire \Tile_X0Y4_S2BEGb[6] ;
 wire \Tile_X0Y4_S2BEGb[7] ;
 wire \Tile_X0Y4_S4BEG[0] ;
 wire \Tile_X0Y4_S4BEG[10] ;
 wire \Tile_X0Y4_S4BEG[11] ;
 wire \Tile_X0Y4_S4BEG[12] ;
 wire \Tile_X0Y4_S4BEG[13] ;
 wire \Tile_X0Y4_S4BEG[14] ;
 wire \Tile_X0Y4_S4BEG[15] ;
 wire \Tile_X0Y4_S4BEG[1] ;
 wire \Tile_X0Y4_S4BEG[2] ;
 wire \Tile_X0Y4_S4BEG[3] ;
 wire \Tile_X0Y4_S4BEG[4] ;
 wire \Tile_X0Y4_S4BEG[5] ;
 wire \Tile_X0Y4_S4BEG[6] ;
 wire \Tile_X0Y4_S4BEG[7] ;
 wire \Tile_X0Y4_S4BEG[8] ;
 wire \Tile_X0Y4_S4BEG[9] ;
 wire Tile_X0Y4_UserCLKo;
 wire \Tile_X0Y5_E1BEG[0] ;
 wire \Tile_X0Y5_E1BEG[1] ;
 wire \Tile_X0Y5_E1BEG[2] ;
 wire \Tile_X0Y5_E1BEG[3] ;
 wire \Tile_X0Y5_E2BEG[0] ;
 wire \Tile_X0Y5_E2BEG[1] ;
 wire \Tile_X0Y5_E2BEG[2] ;
 wire \Tile_X0Y5_E2BEG[3] ;
 wire \Tile_X0Y5_E2BEG[4] ;
 wire \Tile_X0Y5_E2BEG[5] ;
 wire \Tile_X0Y5_E2BEG[6] ;
 wire \Tile_X0Y5_E2BEG[7] ;
 wire \Tile_X0Y5_E2BEGb[0] ;
 wire \Tile_X0Y5_E2BEGb[1] ;
 wire \Tile_X0Y5_E2BEGb[2] ;
 wire \Tile_X0Y5_E2BEGb[3] ;
 wire \Tile_X0Y5_E2BEGb[4] ;
 wire \Tile_X0Y5_E2BEGb[5] ;
 wire \Tile_X0Y5_E2BEGb[6] ;
 wire \Tile_X0Y5_E2BEGb[7] ;
 wire \Tile_X0Y5_E6BEG[0] ;
 wire \Tile_X0Y5_E6BEG[10] ;
 wire \Tile_X0Y5_E6BEG[11] ;
 wire \Tile_X0Y5_E6BEG[1] ;
 wire \Tile_X0Y5_E6BEG[2] ;
 wire \Tile_X0Y5_E6BEG[3] ;
 wire \Tile_X0Y5_E6BEG[4] ;
 wire \Tile_X0Y5_E6BEG[5] ;
 wire \Tile_X0Y5_E6BEG[6] ;
 wire \Tile_X0Y5_E6BEG[7] ;
 wire \Tile_X0Y5_E6BEG[8] ;
 wire \Tile_X0Y5_E6BEG[9] ;
 wire \Tile_X0Y5_EE4BEG[0] ;
 wire \Tile_X0Y5_EE4BEG[10] ;
 wire \Tile_X0Y5_EE4BEG[11] ;
 wire \Tile_X0Y5_EE4BEG[12] ;
 wire \Tile_X0Y5_EE4BEG[13] ;
 wire \Tile_X0Y5_EE4BEG[14] ;
 wire \Tile_X0Y5_EE4BEG[15] ;
 wire \Tile_X0Y5_EE4BEG[1] ;
 wire \Tile_X0Y5_EE4BEG[2] ;
 wire \Tile_X0Y5_EE4BEG[3] ;
 wire \Tile_X0Y5_EE4BEG[4] ;
 wire \Tile_X0Y5_EE4BEG[5] ;
 wire \Tile_X0Y5_EE4BEG[6] ;
 wire \Tile_X0Y5_EE4BEG[7] ;
 wire \Tile_X0Y5_EE4BEG[8] ;
 wire \Tile_X0Y5_EE4BEG[9] ;
 wire \Tile_X0Y5_FrameData_O[0] ;
 wire \Tile_X0Y5_FrameData_O[10] ;
 wire \Tile_X0Y5_FrameData_O[11] ;
 wire \Tile_X0Y5_FrameData_O[12] ;
 wire \Tile_X0Y5_FrameData_O[13] ;
 wire \Tile_X0Y5_FrameData_O[14] ;
 wire \Tile_X0Y5_FrameData_O[15] ;
 wire \Tile_X0Y5_FrameData_O[16] ;
 wire \Tile_X0Y5_FrameData_O[17] ;
 wire \Tile_X0Y5_FrameData_O[18] ;
 wire \Tile_X0Y5_FrameData_O[19] ;
 wire \Tile_X0Y5_FrameData_O[1] ;
 wire \Tile_X0Y5_FrameData_O[20] ;
 wire \Tile_X0Y5_FrameData_O[21] ;
 wire \Tile_X0Y5_FrameData_O[22] ;
 wire \Tile_X0Y5_FrameData_O[23] ;
 wire \Tile_X0Y5_FrameData_O[24] ;
 wire \Tile_X0Y5_FrameData_O[25] ;
 wire \Tile_X0Y5_FrameData_O[26] ;
 wire \Tile_X0Y5_FrameData_O[27] ;
 wire \Tile_X0Y5_FrameData_O[28] ;
 wire \Tile_X0Y5_FrameData_O[29] ;
 wire \Tile_X0Y5_FrameData_O[2] ;
 wire \Tile_X0Y5_FrameData_O[30] ;
 wire \Tile_X0Y5_FrameData_O[31] ;
 wire \Tile_X0Y5_FrameData_O[3] ;
 wire \Tile_X0Y5_FrameData_O[4] ;
 wire \Tile_X0Y5_FrameData_O[5] ;
 wire \Tile_X0Y5_FrameData_O[6] ;
 wire \Tile_X0Y5_FrameData_O[7] ;
 wire \Tile_X0Y5_FrameData_O[8] ;
 wire \Tile_X0Y5_FrameData_O[9] ;
 wire \Tile_X0Y5_FrameStrobe_O[0] ;
 wire \Tile_X0Y5_FrameStrobe_O[10] ;
 wire \Tile_X0Y5_FrameStrobe_O[11] ;
 wire \Tile_X0Y5_FrameStrobe_O[12] ;
 wire \Tile_X0Y5_FrameStrobe_O[13] ;
 wire \Tile_X0Y5_FrameStrobe_O[14] ;
 wire \Tile_X0Y5_FrameStrobe_O[15] ;
 wire \Tile_X0Y5_FrameStrobe_O[16] ;
 wire \Tile_X0Y5_FrameStrobe_O[17] ;
 wire \Tile_X0Y5_FrameStrobe_O[18] ;
 wire \Tile_X0Y5_FrameStrobe_O[19] ;
 wire \Tile_X0Y5_FrameStrobe_O[1] ;
 wire \Tile_X0Y5_FrameStrobe_O[2] ;
 wire \Tile_X0Y5_FrameStrobe_O[3] ;
 wire \Tile_X0Y5_FrameStrobe_O[4] ;
 wire \Tile_X0Y5_FrameStrobe_O[5] ;
 wire \Tile_X0Y5_FrameStrobe_O[6] ;
 wire \Tile_X0Y5_FrameStrobe_O[7] ;
 wire \Tile_X0Y5_FrameStrobe_O[8] ;
 wire \Tile_X0Y5_FrameStrobe_O[9] ;
 wire \Tile_X0Y5_N1BEG[0] ;
 wire \Tile_X0Y5_N1BEG[1] ;
 wire \Tile_X0Y5_N1BEG[2] ;
 wire \Tile_X0Y5_N1BEG[3] ;
 wire \Tile_X0Y5_N2BEG[0] ;
 wire \Tile_X0Y5_N2BEG[1] ;
 wire \Tile_X0Y5_N2BEG[2] ;
 wire \Tile_X0Y5_N2BEG[3] ;
 wire \Tile_X0Y5_N2BEG[4] ;
 wire \Tile_X0Y5_N2BEG[5] ;
 wire \Tile_X0Y5_N2BEG[6] ;
 wire \Tile_X0Y5_N2BEG[7] ;
 wire \Tile_X0Y5_N2BEGb[0] ;
 wire \Tile_X0Y5_N2BEGb[1] ;
 wire \Tile_X0Y5_N2BEGb[2] ;
 wire \Tile_X0Y5_N2BEGb[3] ;
 wire \Tile_X0Y5_N2BEGb[4] ;
 wire \Tile_X0Y5_N2BEGb[5] ;
 wire \Tile_X0Y5_N2BEGb[6] ;
 wire \Tile_X0Y5_N2BEGb[7] ;
 wire \Tile_X0Y5_N4BEG[0] ;
 wire \Tile_X0Y5_N4BEG[10] ;
 wire \Tile_X0Y5_N4BEG[11] ;
 wire \Tile_X0Y5_N4BEG[12] ;
 wire \Tile_X0Y5_N4BEG[13] ;
 wire \Tile_X0Y5_N4BEG[14] ;
 wire \Tile_X0Y5_N4BEG[15] ;
 wire \Tile_X0Y5_N4BEG[1] ;
 wire \Tile_X0Y5_N4BEG[2] ;
 wire \Tile_X0Y5_N4BEG[3] ;
 wire \Tile_X0Y5_N4BEG[4] ;
 wire \Tile_X0Y5_N4BEG[5] ;
 wire \Tile_X0Y5_N4BEG[6] ;
 wire \Tile_X0Y5_N4BEG[7] ;
 wire \Tile_X0Y5_N4BEG[8] ;
 wire \Tile_X0Y5_N4BEG[9] ;
 wire \Tile_X0Y5_S1BEG[0] ;
 wire \Tile_X0Y5_S1BEG[1] ;
 wire \Tile_X0Y5_S1BEG[2] ;
 wire \Tile_X0Y5_S1BEG[3] ;
 wire \Tile_X0Y5_S2BEG[0] ;
 wire \Tile_X0Y5_S2BEG[1] ;
 wire \Tile_X0Y5_S2BEG[2] ;
 wire \Tile_X0Y5_S2BEG[3] ;
 wire \Tile_X0Y5_S2BEG[4] ;
 wire \Tile_X0Y5_S2BEG[5] ;
 wire \Tile_X0Y5_S2BEG[6] ;
 wire \Tile_X0Y5_S2BEG[7] ;
 wire \Tile_X0Y5_S2BEGb[0] ;
 wire \Tile_X0Y5_S2BEGb[1] ;
 wire \Tile_X0Y5_S2BEGb[2] ;
 wire \Tile_X0Y5_S2BEGb[3] ;
 wire \Tile_X0Y5_S2BEGb[4] ;
 wire \Tile_X0Y5_S2BEGb[5] ;
 wire \Tile_X0Y5_S2BEGb[6] ;
 wire \Tile_X0Y5_S2BEGb[7] ;
 wire \Tile_X0Y5_S4BEG[0] ;
 wire \Tile_X0Y5_S4BEG[10] ;
 wire \Tile_X0Y5_S4BEG[11] ;
 wire \Tile_X0Y5_S4BEG[12] ;
 wire \Tile_X0Y5_S4BEG[13] ;
 wire \Tile_X0Y5_S4BEG[14] ;
 wire \Tile_X0Y5_S4BEG[15] ;
 wire \Tile_X0Y5_S4BEG[1] ;
 wire \Tile_X0Y5_S4BEG[2] ;
 wire \Tile_X0Y5_S4BEG[3] ;
 wire \Tile_X0Y5_S4BEG[4] ;
 wire \Tile_X0Y5_S4BEG[5] ;
 wire \Tile_X0Y5_S4BEG[6] ;
 wire \Tile_X0Y5_S4BEG[7] ;
 wire \Tile_X0Y5_S4BEG[8] ;
 wire \Tile_X0Y5_S4BEG[9] ;
 wire Tile_X0Y5_UserCLKo;
 wire \Tile_X0Y6_E1BEG[0] ;
 wire \Tile_X0Y6_E1BEG[1] ;
 wire \Tile_X0Y6_E1BEG[2] ;
 wire \Tile_X0Y6_E1BEG[3] ;
 wire \Tile_X0Y6_E2BEG[0] ;
 wire \Tile_X0Y6_E2BEG[1] ;
 wire \Tile_X0Y6_E2BEG[2] ;
 wire \Tile_X0Y6_E2BEG[3] ;
 wire \Tile_X0Y6_E2BEG[4] ;
 wire \Tile_X0Y6_E2BEG[5] ;
 wire \Tile_X0Y6_E2BEG[6] ;
 wire \Tile_X0Y6_E2BEG[7] ;
 wire \Tile_X0Y6_E2BEGb[0] ;
 wire \Tile_X0Y6_E2BEGb[1] ;
 wire \Tile_X0Y6_E2BEGb[2] ;
 wire \Tile_X0Y6_E2BEGb[3] ;
 wire \Tile_X0Y6_E2BEGb[4] ;
 wire \Tile_X0Y6_E2BEGb[5] ;
 wire \Tile_X0Y6_E2BEGb[6] ;
 wire \Tile_X0Y6_E2BEGb[7] ;
 wire \Tile_X0Y6_E6BEG[0] ;
 wire \Tile_X0Y6_E6BEG[10] ;
 wire \Tile_X0Y6_E6BEG[11] ;
 wire \Tile_X0Y6_E6BEG[1] ;
 wire \Tile_X0Y6_E6BEG[2] ;
 wire \Tile_X0Y6_E6BEG[3] ;
 wire \Tile_X0Y6_E6BEG[4] ;
 wire \Tile_X0Y6_E6BEG[5] ;
 wire \Tile_X0Y6_E6BEG[6] ;
 wire \Tile_X0Y6_E6BEG[7] ;
 wire \Tile_X0Y6_E6BEG[8] ;
 wire \Tile_X0Y6_E6BEG[9] ;
 wire \Tile_X0Y6_EE4BEG[0] ;
 wire \Tile_X0Y6_EE4BEG[10] ;
 wire \Tile_X0Y6_EE4BEG[11] ;
 wire \Tile_X0Y6_EE4BEG[12] ;
 wire \Tile_X0Y6_EE4BEG[13] ;
 wire \Tile_X0Y6_EE4BEG[14] ;
 wire \Tile_X0Y6_EE4BEG[15] ;
 wire \Tile_X0Y6_EE4BEG[1] ;
 wire \Tile_X0Y6_EE4BEG[2] ;
 wire \Tile_X0Y6_EE4BEG[3] ;
 wire \Tile_X0Y6_EE4BEG[4] ;
 wire \Tile_X0Y6_EE4BEG[5] ;
 wire \Tile_X0Y6_EE4BEG[6] ;
 wire \Tile_X0Y6_EE4BEG[7] ;
 wire \Tile_X0Y6_EE4BEG[8] ;
 wire \Tile_X0Y6_EE4BEG[9] ;
 wire \Tile_X0Y6_FrameData_O[0] ;
 wire \Tile_X0Y6_FrameData_O[10] ;
 wire \Tile_X0Y6_FrameData_O[11] ;
 wire \Tile_X0Y6_FrameData_O[12] ;
 wire \Tile_X0Y6_FrameData_O[13] ;
 wire \Tile_X0Y6_FrameData_O[14] ;
 wire \Tile_X0Y6_FrameData_O[15] ;
 wire \Tile_X0Y6_FrameData_O[16] ;
 wire \Tile_X0Y6_FrameData_O[17] ;
 wire \Tile_X0Y6_FrameData_O[18] ;
 wire \Tile_X0Y6_FrameData_O[19] ;
 wire \Tile_X0Y6_FrameData_O[1] ;
 wire \Tile_X0Y6_FrameData_O[20] ;
 wire \Tile_X0Y6_FrameData_O[21] ;
 wire \Tile_X0Y6_FrameData_O[22] ;
 wire \Tile_X0Y6_FrameData_O[23] ;
 wire \Tile_X0Y6_FrameData_O[24] ;
 wire \Tile_X0Y6_FrameData_O[25] ;
 wire \Tile_X0Y6_FrameData_O[26] ;
 wire \Tile_X0Y6_FrameData_O[27] ;
 wire \Tile_X0Y6_FrameData_O[28] ;
 wire \Tile_X0Y6_FrameData_O[29] ;
 wire \Tile_X0Y6_FrameData_O[2] ;
 wire \Tile_X0Y6_FrameData_O[30] ;
 wire \Tile_X0Y6_FrameData_O[31] ;
 wire \Tile_X0Y6_FrameData_O[3] ;
 wire \Tile_X0Y6_FrameData_O[4] ;
 wire \Tile_X0Y6_FrameData_O[5] ;
 wire \Tile_X0Y6_FrameData_O[6] ;
 wire \Tile_X0Y6_FrameData_O[7] ;
 wire \Tile_X0Y6_FrameData_O[8] ;
 wire \Tile_X0Y6_FrameData_O[9] ;
 wire \Tile_X0Y6_FrameStrobe_O[0] ;
 wire \Tile_X0Y6_FrameStrobe_O[10] ;
 wire \Tile_X0Y6_FrameStrobe_O[11] ;
 wire \Tile_X0Y6_FrameStrobe_O[12] ;
 wire \Tile_X0Y6_FrameStrobe_O[13] ;
 wire \Tile_X0Y6_FrameStrobe_O[14] ;
 wire \Tile_X0Y6_FrameStrobe_O[15] ;
 wire \Tile_X0Y6_FrameStrobe_O[16] ;
 wire \Tile_X0Y6_FrameStrobe_O[17] ;
 wire \Tile_X0Y6_FrameStrobe_O[18] ;
 wire \Tile_X0Y6_FrameStrobe_O[19] ;
 wire \Tile_X0Y6_FrameStrobe_O[1] ;
 wire \Tile_X0Y6_FrameStrobe_O[2] ;
 wire \Tile_X0Y6_FrameStrobe_O[3] ;
 wire \Tile_X0Y6_FrameStrobe_O[4] ;
 wire \Tile_X0Y6_FrameStrobe_O[5] ;
 wire \Tile_X0Y6_FrameStrobe_O[6] ;
 wire \Tile_X0Y6_FrameStrobe_O[7] ;
 wire \Tile_X0Y6_FrameStrobe_O[8] ;
 wire \Tile_X0Y6_FrameStrobe_O[9] ;
 wire \Tile_X0Y6_N1BEG[0] ;
 wire \Tile_X0Y6_N1BEG[1] ;
 wire \Tile_X0Y6_N1BEG[2] ;
 wire \Tile_X0Y6_N1BEG[3] ;
 wire \Tile_X0Y6_N2BEG[0] ;
 wire \Tile_X0Y6_N2BEG[1] ;
 wire \Tile_X0Y6_N2BEG[2] ;
 wire \Tile_X0Y6_N2BEG[3] ;
 wire \Tile_X0Y6_N2BEG[4] ;
 wire \Tile_X0Y6_N2BEG[5] ;
 wire \Tile_X0Y6_N2BEG[6] ;
 wire \Tile_X0Y6_N2BEG[7] ;
 wire \Tile_X0Y6_N2BEGb[0] ;
 wire \Tile_X0Y6_N2BEGb[1] ;
 wire \Tile_X0Y6_N2BEGb[2] ;
 wire \Tile_X0Y6_N2BEGb[3] ;
 wire \Tile_X0Y6_N2BEGb[4] ;
 wire \Tile_X0Y6_N2BEGb[5] ;
 wire \Tile_X0Y6_N2BEGb[6] ;
 wire \Tile_X0Y6_N2BEGb[7] ;
 wire \Tile_X0Y6_N4BEG[0] ;
 wire \Tile_X0Y6_N4BEG[10] ;
 wire \Tile_X0Y6_N4BEG[11] ;
 wire \Tile_X0Y6_N4BEG[12] ;
 wire \Tile_X0Y6_N4BEG[13] ;
 wire \Tile_X0Y6_N4BEG[14] ;
 wire \Tile_X0Y6_N4BEG[15] ;
 wire \Tile_X0Y6_N4BEG[1] ;
 wire \Tile_X0Y6_N4BEG[2] ;
 wire \Tile_X0Y6_N4BEG[3] ;
 wire \Tile_X0Y6_N4BEG[4] ;
 wire \Tile_X0Y6_N4BEG[5] ;
 wire \Tile_X0Y6_N4BEG[6] ;
 wire \Tile_X0Y6_N4BEG[7] ;
 wire \Tile_X0Y6_N4BEG[8] ;
 wire \Tile_X0Y6_N4BEG[9] ;
 wire \Tile_X0Y6_S1BEG[0] ;
 wire \Tile_X0Y6_S1BEG[1] ;
 wire \Tile_X0Y6_S1BEG[2] ;
 wire \Tile_X0Y6_S1BEG[3] ;
 wire \Tile_X0Y6_S2BEG[0] ;
 wire \Tile_X0Y6_S2BEG[1] ;
 wire \Tile_X0Y6_S2BEG[2] ;
 wire \Tile_X0Y6_S2BEG[3] ;
 wire \Tile_X0Y6_S2BEG[4] ;
 wire \Tile_X0Y6_S2BEG[5] ;
 wire \Tile_X0Y6_S2BEG[6] ;
 wire \Tile_X0Y6_S2BEG[7] ;
 wire \Tile_X0Y6_S2BEGb[0] ;
 wire \Tile_X0Y6_S2BEGb[1] ;
 wire \Tile_X0Y6_S2BEGb[2] ;
 wire \Tile_X0Y6_S2BEGb[3] ;
 wire \Tile_X0Y6_S2BEGb[4] ;
 wire \Tile_X0Y6_S2BEGb[5] ;
 wire \Tile_X0Y6_S2BEGb[6] ;
 wire \Tile_X0Y6_S2BEGb[7] ;
 wire \Tile_X0Y6_S4BEG[0] ;
 wire \Tile_X0Y6_S4BEG[10] ;
 wire \Tile_X0Y6_S4BEG[11] ;
 wire \Tile_X0Y6_S4BEG[12] ;
 wire \Tile_X0Y6_S4BEG[13] ;
 wire \Tile_X0Y6_S4BEG[14] ;
 wire \Tile_X0Y6_S4BEG[15] ;
 wire \Tile_X0Y6_S4BEG[1] ;
 wire \Tile_X0Y6_S4BEG[2] ;
 wire \Tile_X0Y6_S4BEG[3] ;
 wire \Tile_X0Y6_S4BEG[4] ;
 wire \Tile_X0Y6_S4BEG[5] ;
 wire \Tile_X0Y6_S4BEG[6] ;
 wire \Tile_X0Y6_S4BEG[7] ;
 wire \Tile_X0Y6_S4BEG[8] ;
 wire \Tile_X0Y6_S4BEG[9] ;
 wire Tile_X0Y6_UserCLKo;
 wire \Tile_X0Y7_E1BEG[0] ;
 wire \Tile_X0Y7_E1BEG[1] ;
 wire \Tile_X0Y7_E1BEG[2] ;
 wire \Tile_X0Y7_E1BEG[3] ;
 wire \Tile_X0Y7_E2BEG[0] ;
 wire \Tile_X0Y7_E2BEG[1] ;
 wire \Tile_X0Y7_E2BEG[2] ;
 wire \Tile_X0Y7_E2BEG[3] ;
 wire \Tile_X0Y7_E2BEG[4] ;
 wire \Tile_X0Y7_E2BEG[5] ;
 wire \Tile_X0Y7_E2BEG[6] ;
 wire \Tile_X0Y7_E2BEG[7] ;
 wire \Tile_X0Y7_E2BEGb[0] ;
 wire \Tile_X0Y7_E2BEGb[1] ;
 wire \Tile_X0Y7_E2BEGb[2] ;
 wire \Tile_X0Y7_E2BEGb[3] ;
 wire \Tile_X0Y7_E2BEGb[4] ;
 wire \Tile_X0Y7_E2BEGb[5] ;
 wire \Tile_X0Y7_E2BEGb[6] ;
 wire \Tile_X0Y7_E2BEGb[7] ;
 wire \Tile_X0Y7_E6BEG[0] ;
 wire \Tile_X0Y7_E6BEG[10] ;
 wire \Tile_X0Y7_E6BEG[11] ;
 wire \Tile_X0Y7_E6BEG[1] ;
 wire \Tile_X0Y7_E6BEG[2] ;
 wire \Tile_X0Y7_E6BEG[3] ;
 wire \Tile_X0Y7_E6BEG[4] ;
 wire \Tile_X0Y7_E6BEG[5] ;
 wire \Tile_X0Y7_E6BEG[6] ;
 wire \Tile_X0Y7_E6BEG[7] ;
 wire \Tile_X0Y7_E6BEG[8] ;
 wire \Tile_X0Y7_E6BEG[9] ;
 wire \Tile_X0Y7_EE4BEG[0] ;
 wire \Tile_X0Y7_EE4BEG[10] ;
 wire \Tile_X0Y7_EE4BEG[11] ;
 wire \Tile_X0Y7_EE4BEG[12] ;
 wire \Tile_X0Y7_EE4BEG[13] ;
 wire \Tile_X0Y7_EE4BEG[14] ;
 wire \Tile_X0Y7_EE4BEG[15] ;
 wire \Tile_X0Y7_EE4BEG[1] ;
 wire \Tile_X0Y7_EE4BEG[2] ;
 wire \Tile_X0Y7_EE4BEG[3] ;
 wire \Tile_X0Y7_EE4BEG[4] ;
 wire \Tile_X0Y7_EE4BEG[5] ;
 wire \Tile_X0Y7_EE4BEG[6] ;
 wire \Tile_X0Y7_EE4BEG[7] ;
 wire \Tile_X0Y7_EE4BEG[8] ;
 wire \Tile_X0Y7_EE4BEG[9] ;
 wire \Tile_X0Y7_FrameData_O[0] ;
 wire \Tile_X0Y7_FrameData_O[10] ;
 wire \Tile_X0Y7_FrameData_O[11] ;
 wire \Tile_X0Y7_FrameData_O[12] ;
 wire \Tile_X0Y7_FrameData_O[13] ;
 wire \Tile_X0Y7_FrameData_O[14] ;
 wire \Tile_X0Y7_FrameData_O[15] ;
 wire \Tile_X0Y7_FrameData_O[16] ;
 wire \Tile_X0Y7_FrameData_O[17] ;
 wire \Tile_X0Y7_FrameData_O[18] ;
 wire \Tile_X0Y7_FrameData_O[19] ;
 wire \Tile_X0Y7_FrameData_O[1] ;
 wire \Tile_X0Y7_FrameData_O[20] ;
 wire \Tile_X0Y7_FrameData_O[21] ;
 wire \Tile_X0Y7_FrameData_O[22] ;
 wire \Tile_X0Y7_FrameData_O[23] ;
 wire \Tile_X0Y7_FrameData_O[24] ;
 wire \Tile_X0Y7_FrameData_O[25] ;
 wire \Tile_X0Y7_FrameData_O[26] ;
 wire \Tile_X0Y7_FrameData_O[27] ;
 wire \Tile_X0Y7_FrameData_O[28] ;
 wire \Tile_X0Y7_FrameData_O[29] ;
 wire \Tile_X0Y7_FrameData_O[2] ;
 wire \Tile_X0Y7_FrameData_O[30] ;
 wire \Tile_X0Y7_FrameData_O[31] ;
 wire \Tile_X0Y7_FrameData_O[3] ;
 wire \Tile_X0Y7_FrameData_O[4] ;
 wire \Tile_X0Y7_FrameData_O[5] ;
 wire \Tile_X0Y7_FrameData_O[6] ;
 wire \Tile_X0Y7_FrameData_O[7] ;
 wire \Tile_X0Y7_FrameData_O[8] ;
 wire \Tile_X0Y7_FrameData_O[9] ;
 wire \Tile_X0Y7_FrameStrobe_O[0] ;
 wire \Tile_X0Y7_FrameStrobe_O[10] ;
 wire \Tile_X0Y7_FrameStrobe_O[11] ;
 wire \Tile_X0Y7_FrameStrobe_O[12] ;
 wire \Tile_X0Y7_FrameStrobe_O[13] ;
 wire \Tile_X0Y7_FrameStrobe_O[14] ;
 wire \Tile_X0Y7_FrameStrobe_O[15] ;
 wire \Tile_X0Y7_FrameStrobe_O[16] ;
 wire \Tile_X0Y7_FrameStrobe_O[17] ;
 wire \Tile_X0Y7_FrameStrobe_O[18] ;
 wire \Tile_X0Y7_FrameStrobe_O[19] ;
 wire \Tile_X0Y7_FrameStrobe_O[1] ;
 wire \Tile_X0Y7_FrameStrobe_O[2] ;
 wire \Tile_X0Y7_FrameStrobe_O[3] ;
 wire \Tile_X0Y7_FrameStrobe_O[4] ;
 wire \Tile_X0Y7_FrameStrobe_O[5] ;
 wire \Tile_X0Y7_FrameStrobe_O[6] ;
 wire \Tile_X0Y7_FrameStrobe_O[7] ;
 wire \Tile_X0Y7_FrameStrobe_O[8] ;
 wire \Tile_X0Y7_FrameStrobe_O[9] ;
 wire \Tile_X0Y7_N1BEG[0] ;
 wire \Tile_X0Y7_N1BEG[1] ;
 wire \Tile_X0Y7_N1BEG[2] ;
 wire \Tile_X0Y7_N1BEG[3] ;
 wire \Tile_X0Y7_N2BEG[0] ;
 wire \Tile_X0Y7_N2BEG[1] ;
 wire \Tile_X0Y7_N2BEG[2] ;
 wire \Tile_X0Y7_N2BEG[3] ;
 wire \Tile_X0Y7_N2BEG[4] ;
 wire \Tile_X0Y7_N2BEG[5] ;
 wire \Tile_X0Y7_N2BEG[6] ;
 wire \Tile_X0Y7_N2BEG[7] ;
 wire \Tile_X0Y7_N2BEGb[0] ;
 wire \Tile_X0Y7_N2BEGb[1] ;
 wire \Tile_X0Y7_N2BEGb[2] ;
 wire \Tile_X0Y7_N2BEGb[3] ;
 wire \Tile_X0Y7_N2BEGb[4] ;
 wire \Tile_X0Y7_N2BEGb[5] ;
 wire \Tile_X0Y7_N2BEGb[6] ;
 wire \Tile_X0Y7_N2BEGb[7] ;
 wire \Tile_X0Y7_N4BEG[0] ;
 wire \Tile_X0Y7_N4BEG[10] ;
 wire \Tile_X0Y7_N4BEG[11] ;
 wire \Tile_X0Y7_N4BEG[12] ;
 wire \Tile_X0Y7_N4BEG[13] ;
 wire \Tile_X0Y7_N4BEG[14] ;
 wire \Tile_X0Y7_N4BEG[15] ;
 wire \Tile_X0Y7_N4BEG[1] ;
 wire \Tile_X0Y7_N4BEG[2] ;
 wire \Tile_X0Y7_N4BEG[3] ;
 wire \Tile_X0Y7_N4BEG[4] ;
 wire \Tile_X0Y7_N4BEG[5] ;
 wire \Tile_X0Y7_N4BEG[6] ;
 wire \Tile_X0Y7_N4BEG[7] ;
 wire \Tile_X0Y7_N4BEG[8] ;
 wire \Tile_X0Y7_N4BEG[9] ;
 wire \Tile_X0Y7_S1BEG[0] ;
 wire \Tile_X0Y7_S1BEG[1] ;
 wire \Tile_X0Y7_S1BEG[2] ;
 wire \Tile_X0Y7_S1BEG[3] ;
 wire \Tile_X0Y7_S2BEG[0] ;
 wire \Tile_X0Y7_S2BEG[1] ;
 wire \Tile_X0Y7_S2BEG[2] ;
 wire \Tile_X0Y7_S2BEG[3] ;
 wire \Tile_X0Y7_S2BEG[4] ;
 wire \Tile_X0Y7_S2BEG[5] ;
 wire \Tile_X0Y7_S2BEG[6] ;
 wire \Tile_X0Y7_S2BEG[7] ;
 wire \Tile_X0Y7_S2BEGb[0] ;
 wire \Tile_X0Y7_S2BEGb[1] ;
 wire \Tile_X0Y7_S2BEGb[2] ;
 wire \Tile_X0Y7_S2BEGb[3] ;
 wire \Tile_X0Y7_S2BEGb[4] ;
 wire \Tile_X0Y7_S2BEGb[5] ;
 wire \Tile_X0Y7_S2BEGb[6] ;
 wire \Tile_X0Y7_S2BEGb[7] ;
 wire \Tile_X0Y7_S4BEG[0] ;
 wire \Tile_X0Y7_S4BEG[10] ;
 wire \Tile_X0Y7_S4BEG[11] ;
 wire \Tile_X0Y7_S4BEG[12] ;
 wire \Tile_X0Y7_S4BEG[13] ;
 wire \Tile_X0Y7_S4BEG[14] ;
 wire \Tile_X0Y7_S4BEG[15] ;
 wire \Tile_X0Y7_S4BEG[1] ;
 wire \Tile_X0Y7_S4BEG[2] ;
 wire \Tile_X0Y7_S4BEG[3] ;
 wire \Tile_X0Y7_S4BEG[4] ;
 wire \Tile_X0Y7_S4BEG[5] ;
 wire \Tile_X0Y7_S4BEG[6] ;
 wire \Tile_X0Y7_S4BEG[7] ;
 wire \Tile_X0Y7_S4BEG[8] ;
 wire \Tile_X0Y7_S4BEG[9] ;
 wire Tile_X0Y7_UserCLKo;
 wire \Tile_X0Y8_E1BEG[0] ;
 wire \Tile_X0Y8_E1BEG[1] ;
 wire \Tile_X0Y8_E1BEG[2] ;
 wire \Tile_X0Y8_E1BEG[3] ;
 wire \Tile_X0Y8_E2BEG[0] ;
 wire \Tile_X0Y8_E2BEG[1] ;
 wire \Tile_X0Y8_E2BEG[2] ;
 wire \Tile_X0Y8_E2BEG[3] ;
 wire \Tile_X0Y8_E2BEG[4] ;
 wire \Tile_X0Y8_E2BEG[5] ;
 wire \Tile_X0Y8_E2BEG[6] ;
 wire \Tile_X0Y8_E2BEG[7] ;
 wire \Tile_X0Y8_E2BEGb[0] ;
 wire \Tile_X0Y8_E2BEGb[1] ;
 wire \Tile_X0Y8_E2BEGb[2] ;
 wire \Tile_X0Y8_E2BEGb[3] ;
 wire \Tile_X0Y8_E2BEGb[4] ;
 wire \Tile_X0Y8_E2BEGb[5] ;
 wire \Tile_X0Y8_E2BEGb[6] ;
 wire \Tile_X0Y8_E2BEGb[7] ;
 wire \Tile_X0Y8_E6BEG[0] ;
 wire \Tile_X0Y8_E6BEG[10] ;
 wire \Tile_X0Y8_E6BEG[11] ;
 wire \Tile_X0Y8_E6BEG[1] ;
 wire \Tile_X0Y8_E6BEG[2] ;
 wire \Tile_X0Y8_E6BEG[3] ;
 wire \Tile_X0Y8_E6BEG[4] ;
 wire \Tile_X0Y8_E6BEG[5] ;
 wire \Tile_X0Y8_E6BEG[6] ;
 wire \Tile_X0Y8_E6BEG[7] ;
 wire \Tile_X0Y8_E6BEG[8] ;
 wire \Tile_X0Y8_E6BEG[9] ;
 wire \Tile_X0Y8_EE4BEG[0] ;
 wire \Tile_X0Y8_EE4BEG[10] ;
 wire \Tile_X0Y8_EE4BEG[11] ;
 wire \Tile_X0Y8_EE4BEG[12] ;
 wire \Tile_X0Y8_EE4BEG[13] ;
 wire \Tile_X0Y8_EE4BEG[14] ;
 wire \Tile_X0Y8_EE4BEG[15] ;
 wire \Tile_X0Y8_EE4BEG[1] ;
 wire \Tile_X0Y8_EE4BEG[2] ;
 wire \Tile_X0Y8_EE4BEG[3] ;
 wire \Tile_X0Y8_EE4BEG[4] ;
 wire \Tile_X0Y8_EE4BEG[5] ;
 wire \Tile_X0Y8_EE4BEG[6] ;
 wire \Tile_X0Y8_EE4BEG[7] ;
 wire \Tile_X0Y8_EE4BEG[8] ;
 wire \Tile_X0Y8_EE4BEG[9] ;
 wire \Tile_X0Y8_FrameData_O[0] ;
 wire \Tile_X0Y8_FrameData_O[10] ;
 wire \Tile_X0Y8_FrameData_O[11] ;
 wire \Tile_X0Y8_FrameData_O[12] ;
 wire \Tile_X0Y8_FrameData_O[13] ;
 wire \Tile_X0Y8_FrameData_O[14] ;
 wire \Tile_X0Y8_FrameData_O[15] ;
 wire \Tile_X0Y8_FrameData_O[16] ;
 wire \Tile_X0Y8_FrameData_O[17] ;
 wire \Tile_X0Y8_FrameData_O[18] ;
 wire \Tile_X0Y8_FrameData_O[19] ;
 wire \Tile_X0Y8_FrameData_O[1] ;
 wire \Tile_X0Y8_FrameData_O[20] ;
 wire \Tile_X0Y8_FrameData_O[21] ;
 wire \Tile_X0Y8_FrameData_O[22] ;
 wire \Tile_X0Y8_FrameData_O[23] ;
 wire \Tile_X0Y8_FrameData_O[24] ;
 wire \Tile_X0Y8_FrameData_O[25] ;
 wire \Tile_X0Y8_FrameData_O[26] ;
 wire \Tile_X0Y8_FrameData_O[27] ;
 wire \Tile_X0Y8_FrameData_O[28] ;
 wire \Tile_X0Y8_FrameData_O[29] ;
 wire \Tile_X0Y8_FrameData_O[2] ;
 wire \Tile_X0Y8_FrameData_O[30] ;
 wire \Tile_X0Y8_FrameData_O[31] ;
 wire \Tile_X0Y8_FrameData_O[3] ;
 wire \Tile_X0Y8_FrameData_O[4] ;
 wire \Tile_X0Y8_FrameData_O[5] ;
 wire \Tile_X0Y8_FrameData_O[6] ;
 wire \Tile_X0Y8_FrameData_O[7] ;
 wire \Tile_X0Y8_FrameData_O[8] ;
 wire \Tile_X0Y8_FrameData_O[9] ;
 wire \Tile_X0Y8_FrameStrobe_O[0] ;
 wire \Tile_X0Y8_FrameStrobe_O[10] ;
 wire \Tile_X0Y8_FrameStrobe_O[11] ;
 wire \Tile_X0Y8_FrameStrobe_O[12] ;
 wire \Tile_X0Y8_FrameStrobe_O[13] ;
 wire \Tile_X0Y8_FrameStrobe_O[14] ;
 wire \Tile_X0Y8_FrameStrobe_O[15] ;
 wire \Tile_X0Y8_FrameStrobe_O[16] ;
 wire \Tile_X0Y8_FrameStrobe_O[17] ;
 wire \Tile_X0Y8_FrameStrobe_O[18] ;
 wire \Tile_X0Y8_FrameStrobe_O[19] ;
 wire \Tile_X0Y8_FrameStrobe_O[1] ;
 wire \Tile_X0Y8_FrameStrobe_O[2] ;
 wire \Tile_X0Y8_FrameStrobe_O[3] ;
 wire \Tile_X0Y8_FrameStrobe_O[4] ;
 wire \Tile_X0Y8_FrameStrobe_O[5] ;
 wire \Tile_X0Y8_FrameStrobe_O[6] ;
 wire \Tile_X0Y8_FrameStrobe_O[7] ;
 wire \Tile_X0Y8_FrameStrobe_O[8] ;
 wire \Tile_X0Y8_FrameStrobe_O[9] ;
 wire \Tile_X0Y8_N1BEG[0] ;
 wire \Tile_X0Y8_N1BEG[1] ;
 wire \Tile_X0Y8_N1BEG[2] ;
 wire \Tile_X0Y8_N1BEG[3] ;
 wire \Tile_X0Y8_N2BEG[0] ;
 wire \Tile_X0Y8_N2BEG[1] ;
 wire \Tile_X0Y8_N2BEG[2] ;
 wire \Tile_X0Y8_N2BEG[3] ;
 wire \Tile_X0Y8_N2BEG[4] ;
 wire \Tile_X0Y8_N2BEG[5] ;
 wire \Tile_X0Y8_N2BEG[6] ;
 wire \Tile_X0Y8_N2BEG[7] ;
 wire \Tile_X0Y8_N2BEGb[0] ;
 wire \Tile_X0Y8_N2BEGb[1] ;
 wire \Tile_X0Y8_N2BEGb[2] ;
 wire \Tile_X0Y8_N2BEGb[3] ;
 wire \Tile_X0Y8_N2BEGb[4] ;
 wire \Tile_X0Y8_N2BEGb[5] ;
 wire \Tile_X0Y8_N2BEGb[6] ;
 wire \Tile_X0Y8_N2BEGb[7] ;
 wire \Tile_X0Y8_N4BEG[0] ;
 wire \Tile_X0Y8_N4BEG[10] ;
 wire \Tile_X0Y8_N4BEG[11] ;
 wire \Tile_X0Y8_N4BEG[12] ;
 wire \Tile_X0Y8_N4BEG[13] ;
 wire \Tile_X0Y8_N4BEG[14] ;
 wire \Tile_X0Y8_N4BEG[15] ;
 wire \Tile_X0Y8_N4BEG[1] ;
 wire \Tile_X0Y8_N4BEG[2] ;
 wire \Tile_X0Y8_N4BEG[3] ;
 wire \Tile_X0Y8_N4BEG[4] ;
 wire \Tile_X0Y8_N4BEG[5] ;
 wire \Tile_X0Y8_N4BEG[6] ;
 wire \Tile_X0Y8_N4BEG[7] ;
 wire \Tile_X0Y8_N4BEG[8] ;
 wire \Tile_X0Y8_N4BEG[9] ;
 wire \Tile_X0Y8_S1BEG[0] ;
 wire \Tile_X0Y8_S1BEG[1] ;
 wire \Tile_X0Y8_S1BEG[2] ;
 wire \Tile_X0Y8_S1BEG[3] ;
 wire \Tile_X0Y8_S2BEG[0] ;
 wire \Tile_X0Y8_S2BEG[1] ;
 wire \Tile_X0Y8_S2BEG[2] ;
 wire \Tile_X0Y8_S2BEG[3] ;
 wire \Tile_X0Y8_S2BEG[4] ;
 wire \Tile_X0Y8_S2BEG[5] ;
 wire \Tile_X0Y8_S2BEG[6] ;
 wire \Tile_X0Y8_S2BEG[7] ;
 wire \Tile_X0Y8_S2BEGb[0] ;
 wire \Tile_X0Y8_S2BEGb[1] ;
 wire \Tile_X0Y8_S2BEGb[2] ;
 wire \Tile_X0Y8_S2BEGb[3] ;
 wire \Tile_X0Y8_S2BEGb[4] ;
 wire \Tile_X0Y8_S2BEGb[5] ;
 wire \Tile_X0Y8_S2BEGb[6] ;
 wire \Tile_X0Y8_S2BEGb[7] ;
 wire \Tile_X0Y8_S4BEG[0] ;
 wire \Tile_X0Y8_S4BEG[10] ;
 wire \Tile_X0Y8_S4BEG[11] ;
 wire \Tile_X0Y8_S4BEG[12] ;
 wire \Tile_X0Y8_S4BEG[13] ;
 wire \Tile_X0Y8_S4BEG[14] ;
 wire \Tile_X0Y8_S4BEG[15] ;
 wire \Tile_X0Y8_S4BEG[1] ;
 wire \Tile_X0Y8_S4BEG[2] ;
 wire \Tile_X0Y8_S4BEG[3] ;
 wire \Tile_X0Y8_S4BEG[4] ;
 wire \Tile_X0Y8_S4BEG[5] ;
 wire \Tile_X0Y8_S4BEG[6] ;
 wire \Tile_X0Y8_S4BEG[7] ;
 wire \Tile_X0Y8_S4BEG[8] ;
 wire \Tile_X0Y8_S4BEG[9] ;
 wire Tile_X0Y8_UserCLKo;
 wire \Tile_X0Y9_FrameData_O[0] ;
 wire \Tile_X0Y9_FrameData_O[10] ;
 wire \Tile_X0Y9_FrameData_O[11] ;
 wire \Tile_X0Y9_FrameData_O[12] ;
 wire \Tile_X0Y9_FrameData_O[13] ;
 wire \Tile_X0Y9_FrameData_O[14] ;
 wire \Tile_X0Y9_FrameData_O[15] ;
 wire \Tile_X0Y9_FrameData_O[16] ;
 wire \Tile_X0Y9_FrameData_O[17] ;
 wire \Tile_X0Y9_FrameData_O[18] ;
 wire \Tile_X0Y9_FrameData_O[19] ;
 wire \Tile_X0Y9_FrameData_O[1] ;
 wire \Tile_X0Y9_FrameData_O[20] ;
 wire \Tile_X0Y9_FrameData_O[21] ;
 wire \Tile_X0Y9_FrameData_O[22] ;
 wire \Tile_X0Y9_FrameData_O[23] ;
 wire \Tile_X0Y9_FrameData_O[24] ;
 wire \Tile_X0Y9_FrameData_O[25] ;
 wire \Tile_X0Y9_FrameData_O[26] ;
 wire \Tile_X0Y9_FrameData_O[27] ;
 wire \Tile_X0Y9_FrameData_O[28] ;
 wire \Tile_X0Y9_FrameData_O[29] ;
 wire \Tile_X0Y9_FrameData_O[2] ;
 wire \Tile_X0Y9_FrameData_O[30] ;
 wire \Tile_X0Y9_FrameData_O[31] ;
 wire \Tile_X0Y9_FrameData_O[3] ;
 wire \Tile_X0Y9_FrameData_O[4] ;
 wire \Tile_X0Y9_FrameData_O[5] ;
 wire \Tile_X0Y9_FrameData_O[6] ;
 wire \Tile_X0Y9_FrameData_O[7] ;
 wire \Tile_X0Y9_FrameData_O[8] ;
 wire \Tile_X0Y9_FrameData_O[9] ;
 wire \Tile_X0Y9_FrameStrobe_O[0] ;
 wire \Tile_X0Y9_FrameStrobe_O[10] ;
 wire \Tile_X0Y9_FrameStrobe_O[11] ;
 wire \Tile_X0Y9_FrameStrobe_O[12] ;
 wire \Tile_X0Y9_FrameStrobe_O[13] ;
 wire \Tile_X0Y9_FrameStrobe_O[14] ;
 wire \Tile_X0Y9_FrameStrobe_O[15] ;
 wire \Tile_X0Y9_FrameStrobe_O[16] ;
 wire \Tile_X0Y9_FrameStrobe_O[17] ;
 wire \Tile_X0Y9_FrameStrobe_O[18] ;
 wire \Tile_X0Y9_FrameStrobe_O[19] ;
 wire \Tile_X0Y9_FrameStrobe_O[1] ;
 wire \Tile_X0Y9_FrameStrobe_O[2] ;
 wire \Tile_X0Y9_FrameStrobe_O[3] ;
 wire \Tile_X0Y9_FrameStrobe_O[4] ;
 wire \Tile_X0Y9_FrameStrobe_O[5] ;
 wire \Tile_X0Y9_FrameStrobe_O[6] ;
 wire \Tile_X0Y9_FrameStrobe_O[7] ;
 wire \Tile_X0Y9_FrameStrobe_O[8] ;
 wire \Tile_X0Y9_FrameStrobe_O[9] ;
 wire \Tile_X0Y9_N1BEG[0] ;
 wire \Tile_X0Y9_N1BEG[1] ;
 wire \Tile_X0Y9_N1BEG[2] ;
 wire \Tile_X0Y9_N1BEG[3] ;
 wire \Tile_X0Y9_N2BEG[0] ;
 wire \Tile_X0Y9_N2BEG[1] ;
 wire \Tile_X0Y9_N2BEG[2] ;
 wire \Tile_X0Y9_N2BEG[3] ;
 wire \Tile_X0Y9_N2BEG[4] ;
 wire \Tile_X0Y9_N2BEG[5] ;
 wire \Tile_X0Y9_N2BEG[6] ;
 wire \Tile_X0Y9_N2BEG[7] ;
 wire \Tile_X0Y9_N2BEGb[0] ;
 wire \Tile_X0Y9_N2BEGb[1] ;
 wire \Tile_X0Y9_N2BEGb[2] ;
 wire \Tile_X0Y9_N2BEGb[3] ;
 wire \Tile_X0Y9_N2BEGb[4] ;
 wire \Tile_X0Y9_N2BEGb[5] ;
 wire \Tile_X0Y9_N2BEGb[6] ;
 wire \Tile_X0Y9_N2BEGb[7] ;
 wire \Tile_X0Y9_N4BEG[0] ;
 wire \Tile_X0Y9_N4BEG[10] ;
 wire \Tile_X0Y9_N4BEG[11] ;
 wire \Tile_X0Y9_N4BEG[12] ;
 wire \Tile_X0Y9_N4BEG[13] ;
 wire \Tile_X0Y9_N4BEG[14] ;
 wire \Tile_X0Y9_N4BEG[15] ;
 wire \Tile_X0Y9_N4BEG[1] ;
 wire \Tile_X0Y9_N4BEG[2] ;
 wire \Tile_X0Y9_N4BEG[3] ;
 wire \Tile_X0Y9_N4BEG[4] ;
 wire \Tile_X0Y9_N4BEG[5] ;
 wire \Tile_X0Y9_N4BEG[6] ;
 wire \Tile_X0Y9_N4BEG[7] ;
 wire \Tile_X0Y9_N4BEG[8] ;
 wire \Tile_X0Y9_N4BEG[9] ;
 wire Tile_X0Y9_UserCLKo;
 wire \Tile_X1Y0_FrameData_O[0] ;
 wire \Tile_X1Y0_FrameData_O[10] ;
 wire \Tile_X1Y0_FrameData_O[11] ;
 wire \Tile_X1Y0_FrameData_O[12] ;
 wire \Tile_X1Y0_FrameData_O[13] ;
 wire \Tile_X1Y0_FrameData_O[14] ;
 wire \Tile_X1Y0_FrameData_O[15] ;
 wire \Tile_X1Y0_FrameData_O[16] ;
 wire \Tile_X1Y0_FrameData_O[17] ;
 wire \Tile_X1Y0_FrameData_O[18] ;
 wire \Tile_X1Y0_FrameData_O[19] ;
 wire \Tile_X1Y0_FrameData_O[1] ;
 wire \Tile_X1Y0_FrameData_O[20] ;
 wire \Tile_X1Y0_FrameData_O[21] ;
 wire \Tile_X1Y0_FrameData_O[22] ;
 wire \Tile_X1Y0_FrameData_O[23] ;
 wire \Tile_X1Y0_FrameData_O[24] ;
 wire \Tile_X1Y0_FrameData_O[25] ;
 wire \Tile_X1Y0_FrameData_O[26] ;
 wire \Tile_X1Y0_FrameData_O[27] ;
 wire \Tile_X1Y0_FrameData_O[28] ;
 wire \Tile_X1Y0_FrameData_O[29] ;
 wire \Tile_X1Y0_FrameData_O[2] ;
 wire \Tile_X1Y0_FrameData_O[30] ;
 wire \Tile_X1Y0_FrameData_O[31] ;
 wire \Tile_X1Y0_FrameData_O[3] ;
 wire \Tile_X1Y0_FrameData_O[4] ;
 wire \Tile_X1Y0_FrameData_O[5] ;
 wire \Tile_X1Y0_FrameData_O[6] ;
 wire \Tile_X1Y0_FrameData_O[7] ;
 wire \Tile_X1Y0_FrameData_O[8] ;
 wire \Tile_X1Y0_FrameData_O[9] ;
 wire \Tile_X1Y0_FrameStrobe_O[0] ;
 wire \Tile_X1Y0_FrameStrobe_O[10] ;
 wire \Tile_X1Y0_FrameStrobe_O[11] ;
 wire \Tile_X1Y0_FrameStrobe_O[12] ;
 wire \Tile_X1Y0_FrameStrobe_O[13] ;
 wire \Tile_X1Y0_FrameStrobe_O[14] ;
 wire \Tile_X1Y0_FrameStrobe_O[15] ;
 wire \Tile_X1Y0_FrameStrobe_O[16] ;
 wire \Tile_X1Y0_FrameStrobe_O[17] ;
 wire \Tile_X1Y0_FrameStrobe_O[18] ;
 wire \Tile_X1Y0_FrameStrobe_O[19] ;
 wire \Tile_X1Y0_FrameStrobe_O[1] ;
 wire \Tile_X1Y0_FrameStrobe_O[2] ;
 wire \Tile_X1Y0_FrameStrobe_O[3] ;
 wire \Tile_X1Y0_FrameStrobe_O[4] ;
 wire \Tile_X1Y0_FrameStrobe_O[5] ;
 wire \Tile_X1Y0_FrameStrobe_O[6] ;
 wire \Tile_X1Y0_FrameStrobe_O[7] ;
 wire \Tile_X1Y0_FrameStrobe_O[8] ;
 wire \Tile_X1Y0_FrameStrobe_O[9] ;
 wire \Tile_X1Y0_S1BEG[0] ;
 wire \Tile_X1Y0_S1BEG[1] ;
 wire \Tile_X1Y0_S1BEG[2] ;
 wire \Tile_X1Y0_S1BEG[3] ;
 wire \Tile_X1Y0_S2BEG[0] ;
 wire \Tile_X1Y0_S2BEG[1] ;
 wire \Tile_X1Y0_S2BEG[2] ;
 wire \Tile_X1Y0_S2BEG[3] ;
 wire \Tile_X1Y0_S2BEG[4] ;
 wire \Tile_X1Y0_S2BEG[5] ;
 wire \Tile_X1Y0_S2BEG[6] ;
 wire \Tile_X1Y0_S2BEG[7] ;
 wire \Tile_X1Y0_S2BEGb[0] ;
 wire \Tile_X1Y0_S2BEGb[1] ;
 wire \Tile_X1Y0_S2BEGb[2] ;
 wire \Tile_X1Y0_S2BEGb[3] ;
 wire \Tile_X1Y0_S2BEGb[4] ;
 wire \Tile_X1Y0_S2BEGb[5] ;
 wire \Tile_X1Y0_S2BEGb[6] ;
 wire \Tile_X1Y0_S2BEGb[7] ;
 wire \Tile_X1Y0_S4BEG[0] ;
 wire \Tile_X1Y0_S4BEG[10] ;
 wire \Tile_X1Y0_S4BEG[11] ;
 wire \Tile_X1Y0_S4BEG[12] ;
 wire \Tile_X1Y0_S4BEG[13] ;
 wire \Tile_X1Y0_S4BEG[14] ;
 wire \Tile_X1Y0_S4BEG[15] ;
 wire \Tile_X1Y0_S4BEG[1] ;
 wire \Tile_X1Y0_S4BEG[2] ;
 wire \Tile_X1Y0_S4BEG[3] ;
 wire \Tile_X1Y0_S4BEG[4] ;
 wire \Tile_X1Y0_S4BEG[5] ;
 wire \Tile_X1Y0_S4BEG[6] ;
 wire \Tile_X1Y0_S4BEG[7] ;
 wire \Tile_X1Y0_S4BEG[8] ;
 wire \Tile_X1Y0_S4BEG[9] ;
 wire \Tile_X1Y0_SS4BEG[0] ;
 wire \Tile_X1Y0_SS4BEG[10] ;
 wire \Tile_X1Y0_SS4BEG[11] ;
 wire \Tile_X1Y0_SS4BEG[12] ;
 wire \Tile_X1Y0_SS4BEG[13] ;
 wire \Tile_X1Y0_SS4BEG[14] ;
 wire \Tile_X1Y0_SS4BEG[15] ;
 wire \Tile_X1Y0_SS4BEG[1] ;
 wire \Tile_X1Y0_SS4BEG[2] ;
 wire \Tile_X1Y0_SS4BEG[3] ;
 wire \Tile_X1Y0_SS4BEG[4] ;
 wire \Tile_X1Y0_SS4BEG[5] ;
 wire \Tile_X1Y0_SS4BEG[6] ;
 wire \Tile_X1Y0_SS4BEG[7] ;
 wire \Tile_X1Y0_SS4BEG[8] ;
 wire \Tile_X1Y0_SS4BEG[9] ;
 wire Tile_X1Y0_UserCLKo;
 wire Tile_X1Y1_Co;
 wire \Tile_X1Y1_E1BEG[0] ;
 wire \Tile_X1Y1_E1BEG[1] ;
 wire \Tile_X1Y1_E1BEG[2] ;
 wire \Tile_X1Y1_E1BEG[3] ;
 wire \Tile_X1Y1_E2BEG[0] ;
 wire \Tile_X1Y1_E2BEG[1] ;
 wire \Tile_X1Y1_E2BEG[2] ;
 wire \Tile_X1Y1_E2BEG[3] ;
 wire \Tile_X1Y1_E2BEG[4] ;
 wire \Tile_X1Y1_E2BEG[5] ;
 wire \Tile_X1Y1_E2BEG[6] ;
 wire \Tile_X1Y1_E2BEG[7] ;
 wire \Tile_X1Y1_E2BEGb[0] ;
 wire \Tile_X1Y1_E2BEGb[1] ;
 wire \Tile_X1Y1_E2BEGb[2] ;
 wire \Tile_X1Y1_E2BEGb[3] ;
 wire \Tile_X1Y1_E2BEGb[4] ;
 wire \Tile_X1Y1_E2BEGb[5] ;
 wire \Tile_X1Y1_E2BEGb[6] ;
 wire \Tile_X1Y1_E2BEGb[7] ;
 wire \Tile_X1Y1_E6BEG[0] ;
 wire \Tile_X1Y1_E6BEG[10] ;
 wire \Tile_X1Y1_E6BEG[11] ;
 wire \Tile_X1Y1_E6BEG[1] ;
 wire \Tile_X1Y1_E6BEG[2] ;
 wire \Tile_X1Y1_E6BEG[3] ;
 wire \Tile_X1Y1_E6BEG[4] ;
 wire \Tile_X1Y1_E6BEG[5] ;
 wire \Tile_X1Y1_E6BEG[6] ;
 wire \Tile_X1Y1_E6BEG[7] ;
 wire \Tile_X1Y1_E6BEG[8] ;
 wire \Tile_X1Y1_E6BEG[9] ;
 wire \Tile_X1Y1_EE4BEG[0] ;
 wire \Tile_X1Y1_EE4BEG[10] ;
 wire \Tile_X1Y1_EE4BEG[11] ;
 wire \Tile_X1Y1_EE4BEG[12] ;
 wire \Tile_X1Y1_EE4BEG[13] ;
 wire \Tile_X1Y1_EE4BEG[14] ;
 wire \Tile_X1Y1_EE4BEG[15] ;
 wire \Tile_X1Y1_EE4BEG[1] ;
 wire \Tile_X1Y1_EE4BEG[2] ;
 wire \Tile_X1Y1_EE4BEG[3] ;
 wire \Tile_X1Y1_EE4BEG[4] ;
 wire \Tile_X1Y1_EE4BEG[5] ;
 wire \Tile_X1Y1_EE4BEG[6] ;
 wire \Tile_X1Y1_EE4BEG[7] ;
 wire \Tile_X1Y1_EE4BEG[8] ;
 wire \Tile_X1Y1_EE4BEG[9] ;
 wire \Tile_X1Y1_FrameData_O[0] ;
 wire \Tile_X1Y1_FrameData_O[10] ;
 wire \Tile_X1Y1_FrameData_O[11] ;
 wire \Tile_X1Y1_FrameData_O[12] ;
 wire \Tile_X1Y1_FrameData_O[13] ;
 wire \Tile_X1Y1_FrameData_O[14] ;
 wire \Tile_X1Y1_FrameData_O[15] ;
 wire \Tile_X1Y1_FrameData_O[16] ;
 wire \Tile_X1Y1_FrameData_O[17] ;
 wire \Tile_X1Y1_FrameData_O[18] ;
 wire \Tile_X1Y1_FrameData_O[19] ;
 wire \Tile_X1Y1_FrameData_O[1] ;
 wire \Tile_X1Y1_FrameData_O[20] ;
 wire \Tile_X1Y1_FrameData_O[21] ;
 wire \Tile_X1Y1_FrameData_O[22] ;
 wire \Tile_X1Y1_FrameData_O[23] ;
 wire \Tile_X1Y1_FrameData_O[24] ;
 wire \Tile_X1Y1_FrameData_O[25] ;
 wire \Tile_X1Y1_FrameData_O[26] ;
 wire \Tile_X1Y1_FrameData_O[27] ;
 wire \Tile_X1Y1_FrameData_O[28] ;
 wire \Tile_X1Y1_FrameData_O[29] ;
 wire \Tile_X1Y1_FrameData_O[2] ;
 wire \Tile_X1Y1_FrameData_O[30] ;
 wire \Tile_X1Y1_FrameData_O[31] ;
 wire \Tile_X1Y1_FrameData_O[3] ;
 wire \Tile_X1Y1_FrameData_O[4] ;
 wire \Tile_X1Y1_FrameData_O[5] ;
 wire \Tile_X1Y1_FrameData_O[6] ;
 wire \Tile_X1Y1_FrameData_O[7] ;
 wire \Tile_X1Y1_FrameData_O[8] ;
 wire \Tile_X1Y1_FrameData_O[9] ;
 wire \Tile_X1Y1_FrameStrobe_O[0] ;
 wire \Tile_X1Y1_FrameStrobe_O[10] ;
 wire \Tile_X1Y1_FrameStrobe_O[11] ;
 wire \Tile_X1Y1_FrameStrobe_O[12] ;
 wire \Tile_X1Y1_FrameStrobe_O[13] ;
 wire \Tile_X1Y1_FrameStrobe_O[14] ;
 wire \Tile_X1Y1_FrameStrobe_O[15] ;
 wire \Tile_X1Y1_FrameStrobe_O[16] ;
 wire \Tile_X1Y1_FrameStrobe_O[17] ;
 wire \Tile_X1Y1_FrameStrobe_O[18] ;
 wire \Tile_X1Y1_FrameStrobe_O[19] ;
 wire \Tile_X1Y1_FrameStrobe_O[1] ;
 wire \Tile_X1Y1_FrameStrobe_O[2] ;
 wire \Tile_X1Y1_FrameStrobe_O[3] ;
 wire \Tile_X1Y1_FrameStrobe_O[4] ;
 wire \Tile_X1Y1_FrameStrobe_O[5] ;
 wire \Tile_X1Y1_FrameStrobe_O[6] ;
 wire \Tile_X1Y1_FrameStrobe_O[7] ;
 wire \Tile_X1Y1_FrameStrobe_O[8] ;
 wire \Tile_X1Y1_FrameStrobe_O[9] ;
 wire \Tile_X1Y1_N1BEG[0] ;
 wire \Tile_X1Y1_N1BEG[1] ;
 wire \Tile_X1Y1_N1BEG[2] ;
 wire \Tile_X1Y1_N1BEG[3] ;
 wire \Tile_X1Y1_N2BEG[0] ;
 wire \Tile_X1Y1_N2BEG[1] ;
 wire \Tile_X1Y1_N2BEG[2] ;
 wire \Tile_X1Y1_N2BEG[3] ;
 wire \Tile_X1Y1_N2BEG[4] ;
 wire \Tile_X1Y1_N2BEG[5] ;
 wire \Tile_X1Y1_N2BEG[6] ;
 wire \Tile_X1Y1_N2BEG[7] ;
 wire \Tile_X1Y1_N2BEGb[0] ;
 wire \Tile_X1Y1_N2BEGb[1] ;
 wire \Tile_X1Y1_N2BEGb[2] ;
 wire \Tile_X1Y1_N2BEGb[3] ;
 wire \Tile_X1Y1_N2BEGb[4] ;
 wire \Tile_X1Y1_N2BEGb[5] ;
 wire \Tile_X1Y1_N2BEGb[6] ;
 wire \Tile_X1Y1_N2BEGb[7] ;
 wire \Tile_X1Y1_N4BEG[0] ;
 wire \Tile_X1Y1_N4BEG[10] ;
 wire \Tile_X1Y1_N4BEG[11] ;
 wire \Tile_X1Y1_N4BEG[12] ;
 wire \Tile_X1Y1_N4BEG[13] ;
 wire \Tile_X1Y1_N4BEG[14] ;
 wire \Tile_X1Y1_N4BEG[15] ;
 wire \Tile_X1Y1_N4BEG[1] ;
 wire \Tile_X1Y1_N4BEG[2] ;
 wire \Tile_X1Y1_N4BEG[3] ;
 wire \Tile_X1Y1_N4BEG[4] ;
 wire \Tile_X1Y1_N4BEG[5] ;
 wire \Tile_X1Y1_N4BEG[6] ;
 wire \Tile_X1Y1_N4BEG[7] ;
 wire \Tile_X1Y1_N4BEG[8] ;
 wire \Tile_X1Y1_N4BEG[9] ;
 wire \Tile_X1Y1_NN4BEG[0] ;
 wire \Tile_X1Y1_NN4BEG[10] ;
 wire \Tile_X1Y1_NN4BEG[11] ;
 wire \Tile_X1Y1_NN4BEG[12] ;
 wire \Tile_X1Y1_NN4BEG[13] ;
 wire \Tile_X1Y1_NN4BEG[14] ;
 wire \Tile_X1Y1_NN4BEG[15] ;
 wire \Tile_X1Y1_NN4BEG[1] ;
 wire \Tile_X1Y1_NN4BEG[2] ;
 wire \Tile_X1Y1_NN4BEG[3] ;
 wire \Tile_X1Y1_NN4BEG[4] ;
 wire \Tile_X1Y1_NN4BEG[5] ;
 wire \Tile_X1Y1_NN4BEG[6] ;
 wire \Tile_X1Y1_NN4BEG[7] ;
 wire \Tile_X1Y1_NN4BEG[8] ;
 wire \Tile_X1Y1_NN4BEG[9] ;
 wire \Tile_X1Y1_S1BEG[0] ;
 wire \Tile_X1Y1_S1BEG[1] ;
 wire \Tile_X1Y1_S1BEG[2] ;
 wire \Tile_X1Y1_S1BEG[3] ;
 wire \Tile_X1Y1_S2BEG[0] ;
 wire \Tile_X1Y1_S2BEG[1] ;
 wire \Tile_X1Y1_S2BEG[2] ;
 wire \Tile_X1Y1_S2BEG[3] ;
 wire \Tile_X1Y1_S2BEG[4] ;
 wire \Tile_X1Y1_S2BEG[5] ;
 wire \Tile_X1Y1_S2BEG[6] ;
 wire \Tile_X1Y1_S2BEG[7] ;
 wire \Tile_X1Y1_S2BEGb[0] ;
 wire \Tile_X1Y1_S2BEGb[1] ;
 wire \Tile_X1Y1_S2BEGb[2] ;
 wire \Tile_X1Y1_S2BEGb[3] ;
 wire \Tile_X1Y1_S2BEGb[4] ;
 wire \Tile_X1Y1_S2BEGb[5] ;
 wire \Tile_X1Y1_S2BEGb[6] ;
 wire \Tile_X1Y1_S2BEGb[7] ;
 wire \Tile_X1Y1_S4BEG[0] ;
 wire \Tile_X1Y1_S4BEG[10] ;
 wire \Tile_X1Y1_S4BEG[11] ;
 wire \Tile_X1Y1_S4BEG[12] ;
 wire \Tile_X1Y1_S4BEG[13] ;
 wire \Tile_X1Y1_S4BEG[14] ;
 wire \Tile_X1Y1_S4BEG[15] ;
 wire \Tile_X1Y1_S4BEG[1] ;
 wire \Tile_X1Y1_S4BEG[2] ;
 wire \Tile_X1Y1_S4BEG[3] ;
 wire \Tile_X1Y1_S4BEG[4] ;
 wire \Tile_X1Y1_S4BEG[5] ;
 wire \Tile_X1Y1_S4BEG[6] ;
 wire \Tile_X1Y1_S4BEG[7] ;
 wire \Tile_X1Y1_S4BEG[8] ;
 wire \Tile_X1Y1_S4BEG[9] ;
 wire \Tile_X1Y1_SS4BEG[0] ;
 wire \Tile_X1Y1_SS4BEG[10] ;
 wire \Tile_X1Y1_SS4BEG[11] ;
 wire \Tile_X1Y1_SS4BEG[12] ;
 wire \Tile_X1Y1_SS4BEG[13] ;
 wire \Tile_X1Y1_SS4BEG[14] ;
 wire \Tile_X1Y1_SS4BEG[15] ;
 wire \Tile_X1Y1_SS4BEG[1] ;
 wire \Tile_X1Y1_SS4BEG[2] ;
 wire \Tile_X1Y1_SS4BEG[3] ;
 wire \Tile_X1Y1_SS4BEG[4] ;
 wire \Tile_X1Y1_SS4BEG[5] ;
 wire \Tile_X1Y1_SS4BEG[6] ;
 wire \Tile_X1Y1_SS4BEG[7] ;
 wire \Tile_X1Y1_SS4BEG[8] ;
 wire \Tile_X1Y1_SS4BEG[9] ;
 wire Tile_X1Y1_UserCLKo;
 wire \Tile_X1Y1_W1BEG[0] ;
 wire \Tile_X1Y1_W1BEG[1] ;
 wire \Tile_X1Y1_W1BEG[2] ;
 wire \Tile_X1Y1_W1BEG[3] ;
 wire \Tile_X1Y1_W2BEG[0] ;
 wire \Tile_X1Y1_W2BEG[1] ;
 wire \Tile_X1Y1_W2BEG[2] ;
 wire \Tile_X1Y1_W2BEG[3] ;
 wire \Tile_X1Y1_W2BEG[4] ;
 wire \Tile_X1Y1_W2BEG[5] ;
 wire \Tile_X1Y1_W2BEG[6] ;
 wire \Tile_X1Y1_W2BEG[7] ;
 wire \Tile_X1Y1_W2BEGb[0] ;
 wire \Tile_X1Y1_W2BEGb[1] ;
 wire \Tile_X1Y1_W2BEGb[2] ;
 wire \Tile_X1Y1_W2BEGb[3] ;
 wire \Tile_X1Y1_W2BEGb[4] ;
 wire \Tile_X1Y1_W2BEGb[5] ;
 wire \Tile_X1Y1_W2BEGb[6] ;
 wire \Tile_X1Y1_W2BEGb[7] ;
 wire \Tile_X1Y1_W6BEG[0] ;
 wire \Tile_X1Y1_W6BEG[10] ;
 wire \Tile_X1Y1_W6BEG[11] ;
 wire \Tile_X1Y1_W6BEG[1] ;
 wire \Tile_X1Y1_W6BEG[2] ;
 wire \Tile_X1Y1_W6BEG[3] ;
 wire \Tile_X1Y1_W6BEG[4] ;
 wire \Tile_X1Y1_W6BEG[5] ;
 wire \Tile_X1Y1_W6BEG[6] ;
 wire \Tile_X1Y1_W6BEG[7] ;
 wire \Tile_X1Y1_W6BEG[8] ;
 wire \Tile_X1Y1_W6BEG[9] ;
 wire \Tile_X1Y1_WW4BEG[0] ;
 wire \Tile_X1Y1_WW4BEG[10] ;
 wire \Tile_X1Y1_WW4BEG[11] ;
 wire \Tile_X1Y1_WW4BEG[12] ;
 wire \Tile_X1Y1_WW4BEG[13] ;
 wire \Tile_X1Y1_WW4BEG[14] ;
 wire \Tile_X1Y1_WW4BEG[15] ;
 wire \Tile_X1Y1_WW4BEG[1] ;
 wire \Tile_X1Y1_WW4BEG[2] ;
 wire \Tile_X1Y1_WW4BEG[3] ;
 wire \Tile_X1Y1_WW4BEG[4] ;
 wire \Tile_X1Y1_WW4BEG[5] ;
 wire \Tile_X1Y1_WW4BEG[6] ;
 wire \Tile_X1Y1_WW4BEG[7] ;
 wire \Tile_X1Y1_WW4BEG[8] ;
 wire \Tile_X1Y1_WW4BEG[9] ;
 wire Tile_X1Y2_Co;
 wire \Tile_X1Y2_E1BEG[0] ;
 wire \Tile_X1Y2_E1BEG[1] ;
 wire \Tile_X1Y2_E1BEG[2] ;
 wire \Tile_X1Y2_E1BEG[3] ;
 wire \Tile_X1Y2_E2BEG[0] ;
 wire \Tile_X1Y2_E2BEG[1] ;
 wire \Tile_X1Y2_E2BEG[2] ;
 wire \Tile_X1Y2_E2BEG[3] ;
 wire \Tile_X1Y2_E2BEG[4] ;
 wire \Tile_X1Y2_E2BEG[5] ;
 wire \Tile_X1Y2_E2BEG[6] ;
 wire \Tile_X1Y2_E2BEG[7] ;
 wire \Tile_X1Y2_E2BEGb[0] ;
 wire \Tile_X1Y2_E2BEGb[1] ;
 wire \Tile_X1Y2_E2BEGb[2] ;
 wire \Tile_X1Y2_E2BEGb[3] ;
 wire \Tile_X1Y2_E2BEGb[4] ;
 wire \Tile_X1Y2_E2BEGb[5] ;
 wire \Tile_X1Y2_E2BEGb[6] ;
 wire \Tile_X1Y2_E2BEGb[7] ;
 wire \Tile_X1Y2_E6BEG[0] ;
 wire \Tile_X1Y2_E6BEG[10] ;
 wire \Tile_X1Y2_E6BEG[11] ;
 wire \Tile_X1Y2_E6BEG[1] ;
 wire \Tile_X1Y2_E6BEG[2] ;
 wire \Tile_X1Y2_E6BEG[3] ;
 wire \Tile_X1Y2_E6BEG[4] ;
 wire \Tile_X1Y2_E6BEG[5] ;
 wire \Tile_X1Y2_E6BEG[6] ;
 wire \Tile_X1Y2_E6BEG[7] ;
 wire \Tile_X1Y2_E6BEG[8] ;
 wire \Tile_X1Y2_E6BEG[9] ;
 wire \Tile_X1Y2_EE4BEG[0] ;
 wire \Tile_X1Y2_EE4BEG[10] ;
 wire \Tile_X1Y2_EE4BEG[11] ;
 wire \Tile_X1Y2_EE4BEG[12] ;
 wire \Tile_X1Y2_EE4BEG[13] ;
 wire \Tile_X1Y2_EE4BEG[14] ;
 wire \Tile_X1Y2_EE4BEG[15] ;
 wire \Tile_X1Y2_EE4BEG[1] ;
 wire \Tile_X1Y2_EE4BEG[2] ;
 wire \Tile_X1Y2_EE4BEG[3] ;
 wire \Tile_X1Y2_EE4BEG[4] ;
 wire \Tile_X1Y2_EE4BEG[5] ;
 wire \Tile_X1Y2_EE4BEG[6] ;
 wire \Tile_X1Y2_EE4BEG[7] ;
 wire \Tile_X1Y2_EE4BEG[8] ;
 wire \Tile_X1Y2_EE4BEG[9] ;
 wire \Tile_X1Y2_FrameData_O[0] ;
 wire \Tile_X1Y2_FrameData_O[10] ;
 wire \Tile_X1Y2_FrameData_O[11] ;
 wire \Tile_X1Y2_FrameData_O[12] ;
 wire \Tile_X1Y2_FrameData_O[13] ;
 wire \Tile_X1Y2_FrameData_O[14] ;
 wire \Tile_X1Y2_FrameData_O[15] ;
 wire \Tile_X1Y2_FrameData_O[16] ;
 wire \Tile_X1Y2_FrameData_O[17] ;
 wire \Tile_X1Y2_FrameData_O[18] ;
 wire \Tile_X1Y2_FrameData_O[19] ;
 wire \Tile_X1Y2_FrameData_O[1] ;
 wire \Tile_X1Y2_FrameData_O[20] ;
 wire \Tile_X1Y2_FrameData_O[21] ;
 wire \Tile_X1Y2_FrameData_O[22] ;
 wire \Tile_X1Y2_FrameData_O[23] ;
 wire \Tile_X1Y2_FrameData_O[24] ;
 wire \Tile_X1Y2_FrameData_O[25] ;
 wire \Tile_X1Y2_FrameData_O[26] ;
 wire \Tile_X1Y2_FrameData_O[27] ;
 wire \Tile_X1Y2_FrameData_O[28] ;
 wire \Tile_X1Y2_FrameData_O[29] ;
 wire \Tile_X1Y2_FrameData_O[2] ;
 wire \Tile_X1Y2_FrameData_O[30] ;
 wire \Tile_X1Y2_FrameData_O[31] ;
 wire \Tile_X1Y2_FrameData_O[3] ;
 wire \Tile_X1Y2_FrameData_O[4] ;
 wire \Tile_X1Y2_FrameData_O[5] ;
 wire \Tile_X1Y2_FrameData_O[6] ;
 wire \Tile_X1Y2_FrameData_O[7] ;
 wire \Tile_X1Y2_FrameData_O[8] ;
 wire \Tile_X1Y2_FrameData_O[9] ;
 wire \Tile_X1Y2_FrameStrobe_O[0] ;
 wire \Tile_X1Y2_FrameStrobe_O[10] ;
 wire \Tile_X1Y2_FrameStrobe_O[11] ;
 wire \Tile_X1Y2_FrameStrobe_O[12] ;
 wire \Tile_X1Y2_FrameStrobe_O[13] ;
 wire \Tile_X1Y2_FrameStrobe_O[14] ;
 wire \Tile_X1Y2_FrameStrobe_O[15] ;
 wire \Tile_X1Y2_FrameStrobe_O[16] ;
 wire \Tile_X1Y2_FrameStrobe_O[17] ;
 wire \Tile_X1Y2_FrameStrobe_O[18] ;
 wire \Tile_X1Y2_FrameStrobe_O[19] ;
 wire \Tile_X1Y2_FrameStrobe_O[1] ;
 wire \Tile_X1Y2_FrameStrobe_O[2] ;
 wire \Tile_X1Y2_FrameStrobe_O[3] ;
 wire \Tile_X1Y2_FrameStrobe_O[4] ;
 wire \Tile_X1Y2_FrameStrobe_O[5] ;
 wire \Tile_X1Y2_FrameStrobe_O[6] ;
 wire \Tile_X1Y2_FrameStrobe_O[7] ;
 wire \Tile_X1Y2_FrameStrobe_O[8] ;
 wire \Tile_X1Y2_FrameStrobe_O[9] ;
 wire \Tile_X1Y2_N1BEG[0] ;
 wire \Tile_X1Y2_N1BEG[1] ;
 wire \Tile_X1Y2_N1BEG[2] ;
 wire \Tile_X1Y2_N1BEG[3] ;
 wire \Tile_X1Y2_N2BEG[0] ;
 wire \Tile_X1Y2_N2BEG[1] ;
 wire \Tile_X1Y2_N2BEG[2] ;
 wire \Tile_X1Y2_N2BEG[3] ;
 wire \Tile_X1Y2_N2BEG[4] ;
 wire \Tile_X1Y2_N2BEG[5] ;
 wire \Tile_X1Y2_N2BEG[6] ;
 wire \Tile_X1Y2_N2BEG[7] ;
 wire \Tile_X1Y2_N2BEGb[0] ;
 wire \Tile_X1Y2_N2BEGb[1] ;
 wire \Tile_X1Y2_N2BEGb[2] ;
 wire \Tile_X1Y2_N2BEGb[3] ;
 wire \Tile_X1Y2_N2BEGb[4] ;
 wire \Tile_X1Y2_N2BEGb[5] ;
 wire \Tile_X1Y2_N2BEGb[6] ;
 wire \Tile_X1Y2_N2BEGb[7] ;
 wire \Tile_X1Y2_N4BEG[0] ;
 wire \Tile_X1Y2_N4BEG[10] ;
 wire \Tile_X1Y2_N4BEG[11] ;
 wire \Tile_X1Y2_N4BEG[12] ;
 wire \Tile_X1Y2_N4BEG[13] ;
 wire \Tile_X1Y2_N4BEG[14] ;
 wire \Tile_X1Y2_N4BEG[15] ;
 wire \Tile_X1Y2_N4BEG[1] ;
 wire \Tile_X1Y2_N4BEG[2] ;
 wire \Tile_X1Y2_N4BEG[3] ;
 wire \Tile_X1Y2_N4BEG[4] ;
 wire \Tile_X1Y2_N4BEG[5] ;
 wire \Tile_X1Y2_N4BEG[6] ;
 wire \Tile_X1Y2_N4BEG[7] ;
 wire \Tile_X1Y2_N4BEG[8] ;
 wire \Tile_X1Y2_N4BEG[9] ;
 wire \Tile_X1Y2_NN4BEG[0] ;
 wire \Tile_X1Y2_NN4BEG[10] ;
 wire \Tile_X1Y2_NN4BEG[11] ;
 wire \Tile_X1Y2_NN4BEG[12] ;
 wire \Tile_X1Y2_NN4BEG[13] ;
 wire \Tile_X1Y2_NN4BEG[14] ;
 wire \Tile_X1Y2_NN4BEG[15] ;
 wire \Tile_X1Y2_NN4BEG[1] ;
 wire \Tile_X1Y2_NN4BEG[2] ;
 wire \Tile_X1Y2_NN4BEG[3] ;
 wire \Tile_X1Y2_NN4BEG[4] ;
 wire \Tile_X1Y2_NN4BEG[5] ;
 wire \Tile_X1Y2_NN4BEG[6] ;
 wire \Tile_X1Y2_NN4BEG[7] ;
 wire \Tile_X1Y2_NN4BEG[8] ;
 wire \Tile_X1Y2_NN4BEG[9] ;
 wire \Tile_X1Y2_S1BEG[0] ;
 wire \Tile_X1Y2_S1BEG[1] ;
 wire \Tile_X1Y2_S1BEG[2] ;
 wire \Tile_X1Y2_S1BEG[3] ;
 wire \Tile_X1Y2_S2BEG[0] ;
 wire \Tile_X1Y2_S2BEG[1] ;
 wire \Tile_X1Y2_S2BEG[2] ;
 wire \Tile_X1Y2_S2BEG[3] ;
 wire \Tile_X1Y2_S2BEG[4] ;
 wire \Tile_X1Y2_S2BEG[5] ;
 wire \Tile_X1Y2_S2BEG[6] ;
 wire \Tile_X1Y2_S2BEG[7] ;
 wire \Tile_X1Y2_S2BEGb[0] ;
 wire \Tile_X1Y2_S2BEGb[1] ;
 wire \Tile_X1Y2_S2BEGb[2] ;
 wire \Tile_X1Y2_S2BEGb[3] ;
 wire \Tile_X1Y2_S2BEGb[4] ;
 wire \Tile_X1Y2_S2BEGb[5] ;
 wire \Tile_X1Y2_S2BEGb[6] ;
 wire \Tile_X1Y2_S2BEGb[7] ;
 wire \Tile_X1Y2_S4BEG[0] ;
 wire \Tile_X1Y2_S4BEG[10] ;
 wire \Tile_X1Y2_S4BEG[11] ;
 wire \Tile_X1Y2_S4BEG[12] ;
 wire \Tile_X1Y2_S4BEG[13] ;
 wire \Tile_X1Y2_S4BEG[14] ;
 wire \Tile_X1Y2_S4BEG[15] ;
 wire \Tile_X1Y2_S4BEG[1] ;
 wire \Tile_X1Y2_S4BEG[2] ;
 wire \Tile_X1Y2_S4BEG[3] ;
 wire \Tile_X1Y2_S4BEG[4] ;
 wire \Tile_X1Y2_S4BEG[5] ;
 wire \Tile_X1Y2_S4BEG[6] ;
 wire \Tile_X1Y2_S4BEG[7] ;
 wire \Tile_X1Y2_S4BEG[8] ;
 wire \Tile_X1Y2_S4BEG[9] ;
 wire \Tile_X1Y2_SS4BEG[0] ;
 wire \Tile_X1Y2_SS4BEG[10] ;
 wire \Tile_X1Y2_SS4BEG[11] ;
 wire \Tile_X1Y2_SS4BEG[12] ;
 wire \Tile_X1Y2_SS4BEG[13] ;
 wire \Tile_X1Y2_SS4BEG[14] ;
 wire \Tile_X1Y2_SS4BEG[15] ;
 wire \Tile_X1Y2_SS4BEG[1] ;
 wire \Tile_X1Y2_SS4BEG[2] ;
 wire \Tile_X1Y2_SS4BEG[3] ;
 wire \Tile_X1Y2_SS4BEG[4] ;
 wire \Tile_X1Y2_SS4BEG[5] ;
 wire \Tile_X1Y2_SS4BEG[6] ;
 wire \Tile_X1Y2_SS4BEG[7] ;
 wire \Tile_X1Y2_SS4BEG[8] ;
 wire \Tile_X1Y2_SS4BEG[9] ;
 wire Tile_X1Y2_UserCLKo;
 wire \Tile_X1Y2_W1BEG[0] ;
 wire \Tile_X1Y2_W1BEG[1] ;
 wire \Tile_X1Y2_W1BEG[2] ;
 wire \Tile_X1Y2_W1BEG[3] ;
 wire \Tile_X1Y2_W2BEG[0] ;
 wire \Tile_X1Y2_W2BEG[1] ;
 wire \Tile_X1Y2_W2BEG[2] ;
 wire \Tile_X1Y2_W2BEG[3] ;
 wire \Tile_X1Y2_W2BEG[4] ;
 wire \Tile_X1Y2_W2BEG[5] ;
 wire \Tile_X1Y2_W2BEG[6] ;
 wire \Tile_X1Y2_W2BEG[7] ;
 wire \Tile_X1Y2_W2BEGb[0] ;
 wire \Tile_X1Y2_W2BEGb[1] ;
 wire \Tile_X1Y2_W2BEGb[2] ;
 wire \Tile_X1Y2_W2BEGb[3] ;
 wire \Tile_X1Y2_W2BEGb[4] ;
 wire \Tile_X1Y2_W2BEGb[5] ;
 wire \Tile_X1Y2_W2BEGb[6] ;
 wire \Tile_X1Y2_W2BEGb[7] ;
 wire \Tile_X1Y2_W6BEG[0] ;
 wire \Tile_X1Y2_W6BEG[10] ;
 wire \Tile_X1Y2_W6BEG[11] ;
 wire \Tile_X1Y2_W6BEG[1] ;
 wire \Tile_X1Y2_W6BEG[2] ;
 wire \Tile_X1Y2_W6BEG[3] ;
 wire \Tile_X1Y2_W6BEG[4] ;
 wire \Tile_X1Y2_W6BEG[5] ;
 wire \Tile_X1Y2_W6BEG[6] ;
 wire \Tile_X1Y2_W6BEG[7] ;
 wire \Tile_X1Y2_W6BEG[8] ;
 wire \Tile_X1Y2_W6BEG[9] ;
 wire \Tile_X1Y2_WW4BEG[0] ;
 wire \Tile_X1Y2_WW4BEG[10] ;
 wire \Tile_X1Y2_WW4BEG[11] ;
 wire \Tile_X1Y2_WW4BEG[12] ;
 wire \Tile_X1Y2_WW4BEG[13] ;
 wire \Tile_X1Y2_WW4BEG[14] ;
 wire \Tile_X1Y2_WW4BEG[15] ;
 wire \Tile_X1Y2_WW4BEG[1] ;
 wire \Tile_X1Y2_WW4BEG[2] ;
 wire \Tile_X1Y2_WW4BEG[3] ;
 wire \Tile_X1Y2_WW4BEG[4] ;
 wire \Tile_X1Y2_WW4BEG[5] ;
 wire \Tile_X1Y2_WW4BEG[6] ;
 wire \Tile_X1Y2_WW4BEG[7] ;
 wire \Tile_X1Y2_WW4BEG[8] ;
 wire \Tile_X1Y2_WW4BEG[9] ;
 wire Tile_X1Y3_Co;
 wire \Tile_X1Y3_E1BEG[0] ;
 wire \Tile_X1Y3_E1BEG[1] ;
 wire \Tile_X1Y3_E1BEG[2] ;
 wire \Tile_X1Y3_E1BEG[3] ;
 wire \Tile_X1Y3_E2BEG[0] ;
 wire \Tile_X1Y3_E2BEG[1] ;
 wire \Tile_X1Y3_E2BEG[2] ;
 wire \Tile_X1Y3_E2BEG[3] ;
 wire \Tile_X1Y3_E2BEG[4] ;
 wire \Tile_X1Y3_E2BEG[5] ;
 wire \Tile_X1Y3_E2BEG[6] ;
 wire \Tile_X1Y3_E2BEG[7] ;
 wire \Tile_X1Y3_E2BEGb[0] ;
 wire \Tile_X1Y3_E2BEGb[1] ;
 wire \Tile_X1Y3_E2BEGb[2] ;
 wire \Tile_X1Y3_E2BEGb[3] ;
 wire \Tile_X1Y3_E2BEGb[4] ;
 wire \Tile_X1Y3_E2BEGb[5] ;
 wire \Tile_X1Y3_E2BEGb[6] ;
 wire \Tile_X1Y3_E2BEGb[7] ;
 wire \Tile_X1Y3_E6BEG[0] ;
 wire \Tile_X1Y3_E6BEG[10] ;
 wire \Tile_X1Y3_E6BEG[11] ;
 wire \Tile_X1Y3_E6BEG[1] ;
 wire \Tile_X1Y3_E6BEG[2] ;
 wire \Tile_X1Y3_E6BEG[3] ;
 wire \Tile_X1Y3_E6BEG[4] ;
 wire \Tile_X1Y3_E6BEG[5] ;
 wire \Tile_X1Y3_E6BEG[6] ;
 wire \Tile_X1Y3_E6BEG[7] ;
 wire \Tile_X1Y3_E6BEG[8] ;
 wire \Tile_X1Y3_E6BEG[9] ;
 wire \Tile_X1Y3_EE4BEG[0] ;
 wire \Tile_X1Y3_EE4BEG[10] ;
 wire \Tile_X1Y3_EE4BEG[11] ;
 wire \Tile_X1Y3_EE4BEG[12] ;
 wire \Tile_X1Y3_EE4BEG[13] ;
 wire \Tile_X1Y3_EE4BEG[14] ;
 wire \Tile_X1Y3_EE4BEG[15] ;
 wire \Tile_X1Y3_EE4BEG[1] ;
 wire \Tile_X1Y3_EE4BEG[2] ;
 wire \Tile_X1Y3_EE4BEG[3] ;
 wire \Tile_X1Y3_EE4BEG[4] ;
 wire \Tile_X1Y3_EE4BEG[5] ;
 wire \Tile_X1Y3_EE4BEG[6] ;
 wire \Tile_X1Y3_EE4BEG[7] ;
 wire \Tile_X1Y3_EE4BEG[8] ;
 wire \Tile_X1Y3_EE4BEG[9] ;
 wire \Tile_X1Y3_FrameData_O[0] ;
 wire \Tile_X1Y3_FrameData_O[10] ;
 wire \Tile_X1Y3_FrameData_O[11] ;
 wire \Tile_X1Y3_FrameData_O[12] ;
 wire \Tile_X1Y3_FrameData_O[13] ;
 wire \Tile_X1Y3_FrameData_O[14] ;
 wire \Tile_X1Y3_FrameData_O[15] ;
 wire \Tile_X1Y3_FrameData_O[16] ;
 wire \Tile_X1Y3_FrameData_O[17] ;
 wire \Tile_X1Y3_FrameData_O[18] ;
 wire \Tile_X1Y3_FrameData_O[19] ;
 wire \Tile_X1Y3_FrameData_O[1] ;
 wire \Tile_X1Y3_FrameData_O[20] ;
 wire \Tile_X1Y3_FrameData_O[21] ;
 wire \Tile_X1Y3_FrameData_O[22] ;
 wire \Tile_X1Y3_FrameData_O[23] ;
 wire \Tile_X1Y3_FrameData_O[24] ;
 wire \Tile_X1Y3_FrameData_O[25] ;
 wire \Tile_X1Y3_FrameData_O[26] ;
 wire \Tile_X1Y3_FrameData_O[27] ;
 wire \Tile_X1Y3_FrameData_O[28] ;
 wire \Tile_X1Y3_FrameData_O[29] ;
 wire \Tile_X1Y3_FrameData_O[2] ;
 wire \Tile_X1Y3_FrameData_O[30] ;
 wire \Tile_X1Y3_FrameData_O[31] ;
 wire \Tile_X1Y3_FrameData_O[3] ;
 wire \Tile_X1Y3_FrameData_O[4] ;
 wire \Tile_X1Y3_FrameData_O[5] ;
 wire \Tile_X1Y3_FrameData_O[6] ;
 wire \Tile_X1Y3_FrameData_O[7] ;
 wire \Tile_X1Y3_FrameData_O[8] ;
 wire \Tile_X1Y3_FrameData_O[9] ;
 wire \Tile_X1Y3_FrameStrobe_O[0] ;
 wire \Tile_X1Y3_FrameStrobe_O[10] ;
 wire \Tile_X1Y3_FrameStrobe_O[11] ;
 wire \Tile_X1Y3_FrameStrobe_O[12] ;
 wire \Tile_X1Y3_FrameStrobe_O[13] ;
 wire \Tile_X1Y3_FrameStrobe_O[14] ;
 wire \Tile_X1Y3_FrameStrobe_O[15] ;
 wire \Tile_X1Y3_FrameStrobe_O[16] ;
 wire \Tile_X1Y3_FrameStrobe_O[17] ;
 wire \Tile_X1Y3_FrameStrobe_O[18] ;
 wire \Tile_X1Y3_FrameStrobe_O[19] ;
 wire \Tile_X1Y3_FrameStrobe_O[1] ;
 wire \Tile_X1Y3_FrameStrobe_O[2] ;
 wire \Tile_X1Y3_FrameStrobe_O[3] ;
 wire \Tile_X1Y3_FrameStrobe_O[4] ;
 wire \Tile_X1Y3_FrameStrobe_O[5] ;
 wire \Tile_X1Y3_FrameStrobe_O[6] ;
 wire \Tile_X1Y3_FrameStrobe_O[7] ;
 wire \Tile_X1Y3_FrameStrobe_O[8] ;
 wire \Tile_X1Y3_FrameStrobe_O[9] ;
 wire \Tile_X1Y3_N1BEG[0] ;
 wire \Tile_X1Y3_N1BEG[1] ;
 wire \Tile_X1Y3_N1BEG[2] ;
 wire \Tile_X1Y3_N1BEG[3] ;
 wire \Tile_X1Y3_N2BEG[0] ;
 wire \Tile_X1Y3_N2BEG[1] ;
 wire \Tile_X1Y3_N2BEG[2] ;
 wire \Tile_X1Y3_N2BEG[3] ;
 wire \Tile_X1Y3_N2BEG[4] ;
 wire \Tile_X1Y3_N2BEG[5] ;
 wire \Tile_X1Y3_N2BEG[6] ;
 wire \Tile_X1Y3_N2BEG[7] ;
 wire \Tile_X1Y3_N2BEGb[0] ;
 wire \Tile_X1Y3_N2BEGb[1] ;
 wire \Tile_X1Y3_N2BEGb[2] ;
 wire \Tile_X1Y3_N2BEGb[3] ;
 wire \Tile_X1Y3_N2BEGb[4] ;
 wire \Tile_X1Y3_N2BEGb[5] ;
 wire \Tile_X1Y3_N2BEGb[6] ;
 wire \Tile_X1Y3_N2BEGb[7] ;
 wire \Tile_X1Y3_N4BEG[0] ;
 wire \Tile_X1Y3_N4BEG[10] ;
 wire \Tile_X1Y3_N4BEG[11] ;
 wire \Tile_X1Y3_N4BEG[12] ;
 wire \Tile_X1Y3_N4BEG[13] ;
 wire \Tile_X1Y3_N4BEG[14] ;
 wire \Tile_X1Y3_N4BEG[15] ;
 wire \Tile_X1Y3_N4BEG[1] ;
 wire \Tile_X1Y3_N4BEG[2] ;
 wire \Tile_X1Y3_N4BEG[3] ;
 wire \Tile_X1Y3_N4BEG[4] ;
 wire \Tile_X1Y3_N4BEG[5] ;
 wire \Tile_X1Y3_N4BEG[6] ;
 wire \Tile_X1Y3_N4BEG[7] ;
 wire \Tile_X1Y3_N4BEG[8] ;
 wire \Tile_X1Y3_N4BEG[9] ;
 wire \Tile_X1Y3_NN4BEG[0] ;
 wire \Tile_X1Y3_NN4BEG[10] ;
 wire \Tile_X1Y3_NN4BEG[11] ;
 wire \Tile_X1Y3_NN4BEG[12] ;
 wire \Tile_X1Y3_NN4BEG[13] ;
 wire \Tile_X1Y3_NN4BEG[14] ;
 wire \Tile_X1Y3_NN4BEG[15] ;
 wire \Tile_X1Y3_NN4BEG[1] ;
 wire \Tile_X1Y3_NN4BEG[2] ;
 wire \Tile_X1Y3_NN4BEG[3] ;
 wire \Tile_X1Y3_NN4BEG[4] ;
 wire \Tile_X1Y3_NN4BEG[5] ;
 wire \Tile_X1Y3_NN4BEG[6] ;
 wire \Tile_X1Y3_NN4BEG[7] ;
 wire \Tile_X1Y3_NN4BEG[8] ;
 wire \Tile_X1Y3_NN4BEG[9] ;
 wire \Tile_X1Y3_S1BEG[0] ;
 wire \Tile_X1Y3_S1BEG[1] ;
 wire \Tile_X1Y3_S1BEG[2] ;
 wire \Tile_X1Y3_S1BEG[3] ;
 wire \Tile_X1Y3_S2BEG[0] ;
 wire \Tile_X1Y3_S2BEG[1] ;
 wire \Tile_X1Y3_S2BEG[2] ;
 wire \Tile_X1Y3_S2BEG[3] ;
 wire \Tile_X1Y3_S2BEG[4] ;
 wire \Tile_X1Y3_S2BEG[5] ;
 wire \Tile_X1Y3_S2BEG[6] ;
 wire \Tile_X1Y3_S2BEG[7] ;
 wire \Tile_X1Y3_S2BEGb[0] ;
 wire \Tile_X1Y3_S2BEGb[1] ;
 wire \Tile_X1Y3_S2BEGb[2] ;
 wire \Tile_X1Y3_S2BEGb[3] ;
 wire \Tile_X1Y3_S2BEGb[4] ;
 wire \Tile_X1Y3_S2BEGb[5] ;
 wire \Tile_X1Y3_S2BEGb[6] ;
 wire \Tile_X1Y3_S2BEGb[7] ;
 wire \Tile_X1Y3_S4BEG[0] ;
 wire \Tile_X1Y3_S4BEG[10] ;
 wire \Tile_X1Y3_S4BEG[11] ;
 wire \Tile_X1Y3_S4BEG[12] ;
 wire \Tile_X1Y3_S4BEG[13] ;
 wire \Tile_X1Y3_S4BEG[14] ;
 wire \Tile_X1Y3_S4BEG[15] ;
 wire \Tile_X1Y3_S4BEG[1] ;
 wire \Tile_X1Y3_S4BEG[2] ;
 wire \Tile_X1Y3_S4BEG[3] ;
 wire \Tile_X1Y3_S4BEG[4] ;
 wire \Tile_X1Y3_S4BEG[5] ;
 wire \Tile_X1Y3_S4BEG[6] ;
 wire \Tile_X1Y3_S4BEG[7] ;
 wire \Tile_X1Y3_S4BEG[8] ;
 wire \Tile_X1Y3_S4BEG[9] ;
 wire \Tile_X1Y3_SS4BEG[0] ;
 wire \Tile_X1Y3_SS4BEG[10] ;
 wire \Tile_X1Y3_SS4BEG[11] ;
 wire \Tile_X1Y3_SS4BEG[12] ;
 wire \Tile_X1Y3_SS4BEG[13] ;
 wire \Tile_X1Y3_SS4BEG[14] ;
 wire \Tile_X1Y3_SS4BEG[15] ;
 wire \Tile_X1Y3_SS4BEG[1] ;
 wire \Tile_X1Y3_SS4BEG[2] ;
 wire \Tile_X1Y3_SS4BEG[3] ;
 wire \Tile_X1Y3_SS4BEG[4] ;
 wire \Tile_X1Y3_SS4BEG[5] ;
 wire \Tile_X1Y3_SS4BEG[6] ;
 wire \Tile_X1Y3_SS4BEG[7] ;
 wire \Tile_X1Y3_SS4BEG[8] ;
 wire \Tile_X1Y3_SS4BEG[9] ;
 wire Tile_X1Y3_UserCLKo;
 wire \Tile_X1Y3_W1BEG[0] ;
 wire \Tile_X1Y3_W1BEG[1] ;
 wire \Tile_X1Y3_W1BEG[2] ;
 wire \Tile_X1Y3_W1BEG[3] ;
 wire \Tile_X1Y3_W2BEG[0] ;
 wire \Tile_X1Y3_W2BEG[1] ;
 wire \Tile_X1Y3_W2BEG[2] ;
 wire \Tile_X1Y3_W2BEG[3] ;
 wire \Tile_X1Y3_W2BEG[4] ;
 wire \Tile_X1Y3_W2BEG[5] ;
 wire \Tile_X1Y3_W2BEG[6] ;
 wire \Tile_X1Y3_W2BEG[7] ;
 wire \Tile_X1Y3_W2BEGb[0] ;
 wire \Tile_X1Y3_W2BEGb[1] ;
 wire \Tile_X1Y3_W2BEGb[2] ;
 wire \Tile_X1Y3_W2BEGb[3] ;
 wire \Tile_X1Y3_W2BEGb[4] ;
 wire \Tile_X1Y3_W2BEGb[5] ;
 wire \Tile_X1Y3_W2BEGb[6] ;
 wire \Tile_X1Y3_W2BEGb[7] ;
 wire \Tile_X1Y3_W6BEG[0] ;
 wire \Tile_X1Y3_W6BEG[10] ;
 wire \Tile_X1Y3_W6BEG[11] ;
 wire \Tile_X1Y3_W6BEG[1] ;
 wire \Tile_X1Y3_W6BEG[2] ;
 wire \Tile_X1Y3_W6BEG[3] ;
 wire \Tile_X1Y3_W6BEG[4] ;
 wire \Tile_X1Y3_W6BEG[5] ;
 wire \Tile_X1Y3_W6BEG[6] ;
 wire \Tile_X1Y3_W6BEG[7] ;
 wire \Tile_X1Y3_W6BEG[8] ;
 wire \Tile_X1Y3_W6BEG[9] ;
 wire \Tile_X1Y3_WW4BEG[0] ;
 wire \Tile_X1Y3_WW4BEG[10] ;
 wire \Tile_X1Y3_WW4BEG[11] ;
 wire \Tile_X1Y3_WW4BEG[12] ;
 wire \Tile_X1Y3_WW4BEG[13] ;
 wire \Tile_X1Y3_WW4BEG[14] ;
 wire \Tile_X1Y3_WW4BEG[15] ;
 wire \Tile_X1Y3_WW4BEG[1] ;
 wire \Tile_X1Y3_WW4BEG[2] ;
 wire \Tile_X1Y3_WW4BEG[3] ;
 wire \Tile_X1Y3_WW4BEG[4] ;
 wire \Tile_X1Y3_WW4BEG[5] ;
 wire \Tile_X1Y3_WW4BEG[6] ;
 wire \Tile_X1Y3_WW4BEG[7] ;
 wire \Tile_X1Y3_WW4BEG[8] ;
 wire \Tile_X1Y3_WW4BEG[9] ;
 wire Tile_X1Y4_Co;
 wire \Tile_X1Y4_E1BEG[0] ;
 wire \Tile_X1Y4_E1BEG[1] ;
 wire \Tile_X1Y4_E1BEG[2] ;
 wire \Tile_X1Y4_E1BEG[3] ;
 wire \Tile_X1Y4_E2BEG[0] ;
 wire \Tile_X1Y4_E2BEG[1] ;
 wire \Tile_X1Y4_E2BEG[2] ;
 wire \Tile_X1Y4_E2BEG[3] ;
 wire \Tile_X1Y4_E2BEG[4] ;
 wire \Tile_X1Y4_E2BEG[5] ;
 wire \Tile_X1Y4_E2BEG[6] ;
 wire \Tile_X1Y4_E2BEG[7] ;
 wire \Tile_X1Y4_E2BEGb[0] ;
 wire \Tile_X1Y4_E2BEGb[1] ;
 wire \Tile_X1Y4_E2BEGb[2] ;
 wire \Tile_X1Y4_E2BEGb[3] ;
 wire \Tile_X1Y4_E2BEGb[4] ;
 wire \Tile_X1Y4_E2BEGb[5] ;
 wire \Tile_X1Y4_E2BEGb[6] ;
 wire \Tile_X1Y4_E2BEGb[7] ;
 wire \Tile_X1Y4_E6BEG[0] ;
 wire \Tile_X1Y4_E6BEG[10] ;
 wire \Tile_X1Y4_E6BEG[11] ;
 wire \Tile_X1Y4_E6BEG[1] ;
 wire \Tile_X1Y4_E6BEG[2] ;
 wire \Tile_X1Y4_E6BEG[3] ;
 wire \Tile_X1Y4_E6BEG[4] ;
 wire \Tile_X1Y4_E6BEG[5] ;
 wire \Tile_X1Y4_E6BEG[6] ;
 wire \Tile_X1Y4_E6BEG[7] ;
 wire \Tile_X1Y4_E6BEG[8] ;
 wire \Tile_X1Y4_E6BEG[9] ;
 wire \Tile_X1Y4_EE4BEG[0] ;
 wire \Tile_X1Y4_EE4BEG[10] ;
 wire \Tile_X1Y4_EE4BEG[11] ;
 wire \Tile_X1Y4_EE4BEG[12] ;
 wire \Tile_X1Y4_EE4BEG[13] ;
 wire \Tile_X1Y4_EE4BEG[14] ;
 wire \Tile_X1Y4_EE4BEG[15] ;
 wire \Tile_X1Y4_EE4BEG[1] ;
 wire \Tile_X1Y4_EE4BEG[2] ;
 wire \Tile_X1Y4_EE4BEG[3] ;
 wire \Tile_X1Y4_EE4BEG[4] ;
 wire \Tile_X1Y4_EE4BEG[5] ;
 wire \Tile_X1Y4_EE4BEG[6] ;
 wire \Tile_X1Y4_EE4BEG[7] ;
 wire \Tile_X1Y4_EE4BEG[8] ;
 wire \Tile_X1Y4_EE4BEG[9] ;
 wire \Tile_X1Y4_FrameData_O[0] ;
 wire \Tile_X1Y4_FrameData_O[10] ;
 wire \Tile_X1Y4_FrameData_O[11] ;
 wire \Tile_X1Y4_FrameData_O[12] ;
 wire \Tile_X1Y4_FrameData_O[13] ;
 wire \Tile_X1Y4_FrameData_O[14] ;
 wire \Tile_X1Y4_FrameData_O[15] ;
 wire \Tile_X1Y4_FrameData_O[16] ;
 wire \Tile_X1Y4_FrameData_O[17] ;
 wire \Tile_X1Y4_FrameData_O[18] ;
 wire \Tile_X1Y4_FrameData_O[19] ;
 wire \Tile_X1Y4_FrameData_O[1] ;
 wire \Tile_X1Y4_FrameData_O[20] ;
 wire \Tile_X1Y4_FrameData_O[21] ;
 wire \Tile_X1Y4_FrameData_O[22] ;
 wire \Tile_X1Y4_FrameData_O[23] ;
 wire \Tile_X1Y4_FrameData_O[24] ;
 wire \Tile_X1Y4_FrameData_O[25] ;
 wire \Tile_X1Y4_FrameData_O[26] ;
 wire \Tile_X1Y4_FrameData_O[27] ;
 wire \Tile_X1Y4_FrameData_O[28] ;
 wire \Tile_X1Y4_FrameData_O[29] ;
 wire \Tile_X1Y4_FrameData_O[2] ;
 wire \Tile_X1Y4_FrameData_O[30] ;
 wire \Tile_X1Y4_FrameData_O[31] ;
 wire \Tile_X1Y4_FrameData_O[3] ;
 wire \Tile_X1Y4_FrameData_O[4] ;
 wire \Tile_X1Y4_FrameData_O[5] ;
 wire \Tile_X1Y4_FrameData_O[6] ;
 wire \Tile_X1Y4_FrameData_O[7] ;
 wire \Tile_X1Y4_FrameData_O[8] ;
 wire \Tile_X1Y4_FrameData_O[9] ;
 wire \Tile_X1Y4_FrameStrobe_O[0] ;
 wire \Tile_X1Y4_FrameStrobe_O[10] ;
 wire \Tile_X1Y4_FrameStrobe_O[11] ;
 wire \Tile_X1Y4_FrameStrobe_O[12] ;
 wire \Tile_X1Y4_FrameStrobe_O[13] ;
 wire \Tile_X1Y4_FrameStrobe_O[14] ;
 wire \Tile_X1Y4_FrameStrobe_O[15] ;
 wire \Tile_X1Y4_FrameStrobe_O[16] ;
 wire \Tile_X1Y4_FrameStrobe_O[17] ;
 wire \Tile_X1Y4_FrameStrobe_O[18] ;
 wire \Tile_X1Y4_FrameStrobe_O[19] ;
 wire \Tile_X1Y4_FrameStrobe_O[1] ;
 wire \Tile_X1Y4_FrameStrobe_O[2] ;
 wire \Tile_X1Y4_FrameStrobe_O[3] ;
 wire \Tile_X1Y4_FrameStrobe_O[4] ;
 wire \Tile_X1Y4_FrameStrobe_O[5] ;
 wire \Tile_X1Y4_FrameStrobe_O[6] ;
 wire \Tile_X1Y4_FrameStrobe_O[7] ;
 wire \Tile_X1Y4_FrameStrobe_O[8] ;
 wire \Tile_X1Y4_FrameStrobe_O[9] ;
 wire \Tile_X1Y4_N1BEG[0] ;
 wire \Tile_X1Y4_N1BEG[1] ;
 wire \Tile_X1Y4_N1BEG[2] ;
 wire \Tile_X1Y4_N1BEG[3] ;
 wire \Tile_X1Y4_N2BEG[0] ;
 wire \Tile_X1Y4_N2BEG[1] ;
 wire \Tile_X1Y4_N2BEG[2] ;
 wire \Tile_X1Y4_N2BEG[3] ;
 wire \Tile_X1Y4_N2BEG[4] ;
 wire \Tile_X1Y4_N2BEG[5] ;
 wire \Tile_X1Y4_N2BEG[6] ;
 wire \Tile_X1Y4_N2BEG[7] ;
 wire \Tile_X1Y4_N2BEGb[0] ;
 wire \Tile_X1Y4_N2BEGb[1] ;
 wire \Tile_X1Y4_N2BEGb[2] ;
 wire \Tile_X1Y4_N2BEGb[3] ;
 wire \Tile_X1Y4_N2BEGb[4] ;
 wire \Tile_X1Y4_N2BEGb[5] ;
 wire \Tile_X1Y4_N2BEGb[6] ;
 wire \Tile_X1Y4_N2BEGb[7] ;
 wire \Tile_X1Y4_N4BEG[0] ;
 wire \Tile_X1Y4_N4BEG[10] ;
 wire \Tile_X1Y4_N4BEG[11] ;
 wire \Tile_X1Y4_N4BEG[12] ;
 wire \Tile_X1Y4_N4BEG[13] ;
 wire \Tile_X1Y4_N4BEG[14] ;
 wire \Tile_X1Y4_N4BEG[15] ;
 wire \Tile_X1Y4_N4BEG[1] ;
 wire \Tile_X1Y4_N4BEG[2] ;
 wire \Tile_X1Y4_N4BEG[3] ;
 wire \Tile_X1Y4_N4BEG[4] ;
 wire \Tile_X1Y4_N4BEG[5] ;
 wire \Tile_X1Y4_N4BEG[6] ;
 wire \Tile_X1Y4_N4BEG[7] ;
 wire \Tile_X1Y4_N4BEG[8] ;
 wire \Tile_X1Y4_N4BEG[9] ;
 wire \Tile_X1Y4_NN4BEG[0] ;
 wire \Tile_X1Y4_NN4BEG[10] ;
 wire \Tile_X1Y4_NN4BEG[11] ;
 wire \Tile_X1Y4_NN4BEG[12] ;
 wire \Tile_X1Y4_NN4BEG[13] ;
 wire \Tile_X1Y4_NN4BEG[14] ;
 wire \Tile_X1Y4_NN4BEG[15] ;
 wire \Tile_X1Y4_NN4BEG[1] ;
 wire \Tile_X1Y4_NN4BEG[2] ;
 wire \Tile_X1Y4_NN4BEG[3] ;
 wire \Tile_X1Y4_NN4BEG[4] ;
 wire \Tile_X1Y4_NN4BEG[5] ;
 wire \Tile_X1Y4_NN4BEG[6] ;
 wire \Tile_X1Y4_NN4BEG[7] ;
 wire \Tile_X1Y4_NN4BEG[8] ;
 wire \Tile_X1Y4_NN4BEG[9] ;
 wire \Tile_X1Y4_S1BEG[0] ;
 wire \Tile_X1Y4_S1BEG[1] ;
 wire \Tile_X1Y4_S1BEG[2] ;
 wire \Tile_X1Y4_S1BEG[3] ;
 wire \Tile_X1Y4_S2BEG[0] ;
 wire \Tile_X1Y4_S2BEG[1] ;
 wire \Tile_X1Y4_S2BEG[2] ;
 wire \Tile_X1Y4_S2BEG[3] ;
 wire \Tile_X1Y4_S2BEG[4] ;
 wire \Tile_X1Y4_S2BEG[5] ;
 wire \Tile_X1Y4_S2BEG[6] ;
 wire \Tile_X1Y4_S2BEG[7] ;
 wire \Tile_X1Y4_S2BEGb[0] ;
 wire \Tile_X1Y4_S2BEGb[1] ;
 wire \Tile_X1Y4_S2BEGb[2] ;
 wire \Tile_X1Y4_S2BEGb[3] ;
 wire \Tile_X1Y4_S2BEGb[4] ;
 wire \Tile_X1Y4_S2BEGb[5] ;
 wire \Tile_X1Y4_S2BEGb[6] ;
 wire \Tile_X1Y4_S2BEGb[7] ;
 wire \Tile_X1Y4_S4BEG[0] ;
 wire \Tile_X1Y4_S4BEG[10] ;
 wire \Tile_X1Y4_S4BEG[11] ;
 wire \Tile_X1Y4_S4BEG[12] ;
 wire \Tile_X1Y4_S4BEG[13] ;
 wire \Tile_X1Y4_S4BEG[14] ;
 wire \Tile_X1Y4_S4BEG[15] ;
 wire \Tile_X1Y4_S4BEG[1] ;
 wire \Tile_X1Y4_S4BEG[2] ;
 wire \Tile_X1Y4_S4BEG[3] ;
 wire \Tile_X1Y4_S4BEG[4] ;
 wire \Tile_X1Y4_S4BEG[5] ;
 wire \Tile_X1Y4_S4BEG[6] ;
 wire \Tile_X1Y4_S4BEG[7] ;
 wire \Tile_X1Y4_S4BEG[8] ;
 wire \Tile_X1Y4_S4BEG[9] ;
 wire \Tile_X1Y4_SS4BEG[0] ;
 wire \Tile_X1Y4_SS4BEG[10] ;
 wire \Tile_X1Y4_SS4BEG[11] ;
 wire \Tile_X1Y4_SS4BEG[12] ;
 wire \Tile_X1Y4_SS4BEG[13] ;
 wire \Tile_X1Y4_SS4BEG[14] ;
 wire \Tile_X1Y4_SS4BEG[15] ;
 wire \Tile_X1Y4_SS4BEG[1] ;
 wire \Tile_X1Y4_SS4BEG[2] ;
 wire \Tile_X1Y4_SS4BEG[3] ;
 wire \Tile_X1Y4_SS4BEG[4] ;
 wire \Tile_X1Y4_SS4BEG[5] ;
 wire \Tile_X1Y4_SS4BEG[6] ;
 wire \Tile_X1Y4_SS4BEG[7] ;
 wire \Tile_X1Y4_SS4BEG[8] ;
 wire \Tile_X1Y4_SS4BEG[9] ;
 wire Tile_X1Y4_UserCLKo;
 wire \Tile_X1Y4_W1BEG[0] ;
 wire \Tile_X1Y4_W1BEG[1] ;
 wire \Tile_X1Y4_W1BEG[2] ;
 wire \Tile_X1Y4_W1BEG[3] ;
 wire \Tile_X1Y4_W2BEG[0] ;
 wire \Tile_X1Y4_W2BEG[1] ;
 wire \Tile_X1Y4_W2BEG[2] ;
 wire \Tile_X1Y4_W2BEG[3] ;
 wire \Tile_X1Y4_W2BEG[4] ;
 wire \Tile_X1Y4_W2BEG[5] ;
 wire \Tile_X1Y4_W2BEG[6] ;
 wire \Tile_X1Y4_W2BEG[7] ;
 wire \Tile_X1Y4_W2BEGb[0] ;
 wire \Tile_X1Y4_W2BEGb[1] ;
 wire \Tile_X1Y4_W2BEGb[2] ;
 wire \Tile_X1Y4_W2BEGb[3] ;
 wire \Tile_X1Y4_W2BEGb[4] ;
 wire \Tile_X1Y4_W2BEGb[5] ;
 wire \Tile_X1Y4_W2BEGb[6] ;
 wire \Tile_X1Y4_W2BEGb[7] ;
 wire \Tile_X1Y4_W6BEG[0] ;
 wire \Tile_X1Y4_W6BEG[10] ;
 wire \Tile_X1Y4_W6BEG[11] ;
 wire \Tile_X1Y4_W6BEG[1] ;
 wire \Tile_X1Y4_W6BEG[2] ;
 wire \Tile_X1Y4_W6BEG[3] ;
 wire \Tile_X1Y4_W6BEG[4] ;
 wire \Tile_X1Y4_W6BEG[5] ;
 wire \Tile_X1Y4_W6BEG[6] ;
 wire \Tile_X1Y4_W6BEG[7] ;
 wire \Tile_X1Y4_W6BEG[8] ;
 wire \Tile_X1Y4_W6BEG[9] ;
 wire \Tile_X1Y4_WW4BEG[0] ;
 wire \Tile_X1Y4_WW4BEG[10] ;
 wire \Tile_X1Y4_WW4BEG[11] ;
 wire \Tile_X1Y4_WW4BEG[12] ;
 wire \Tile_X1Y4_WW4BEG[13] ;
 wire \Tile_X1Y4_WW4BEG[14] ;
 wire \Tile_X1Y4_WW4BEG[15] ;
 wire \Tile_X1Y4_WW4BEG[1] ;
 wire \Tile_X1Y4_WW4BEG[2] ;
 wire \Tile_X1Y4_WW4BEG[3] ;
 wire \Tile_X1Y4_WW4BEG[4] ;
 wire \Tile_X1Y4_WW4BEG[5] ;
 wire \Tile_X1Y4_WW4BEG[6] ;
 wire \Tile_X1Y4_WW4BEG[7] ;
 wire \Tile_X1Y4_WW4BEG[8] ;
 wire \Tile_X1Y4_WW4BEG[9] ;
 wire Tile_X1Y5_Co;
 wire \Tile_X1Y5_E1BEG[0] ;
 wire \Tile_X1Y5_E1BEG[1] ;
 wire \Tile_X1Y5_E1BEG[2] ;
 wire \Tile_X1Y5_E1BEG[3] ;
 wire \Tile_X1Y5_E2BEG[0] ;
 wire \Tile_X1Y5_E2BEG[1] ;
 wire \Tile_X1Y5_E2BEG[2] ;
 wire \Tile_X1Y5_E2BEG[3] ;
 wire \Tile_X1Y5_E2BEG[4] ;
 wire \Tile_X1Y5_E2BEG[5] ;
 wire \Tile_X1Y5_E2BEG[6] ;
 wire \Tile_X1Y5_E2BEG[7] ;
 wire \Tile_X1Y5_E2BEGb[0] ;
 wire \Tile_X1Y5_E2BEGb[1] ;
 wire \Tile_X1Y5_E2BEGb[2] ;
 wire \Tile_X1Y5_E2BEGb[3] ;
 wire \Tile_X1Y5_E2BEGb[4] ;
 wire \Tile_X1Y5_E2BEGb[5] ;
 wire \Tile_X1Y5_E2BEGb[6] ;
 wire \Tile_X1Y5_E2BEGb[7] ;
 wire \Tile_X1Y5_E6BEG[0] ;
 wire \Tile_X1Y5_E6BEG[10] ;
 wire \Tile_X1Y5_E6BEG[11] ;
 wire \Tile_X1Y5_E6BEG[1] ;
 wire \Tile_X1Y5_E6BEG[2] ;
 wire \Tile_X1Y5_E6BEG[3] ;
 wire \Tile_X1Y5_E6BEG[4] ;
 wire \Tile_X1Y5_E6BEG[5] ;
 wire \Tile_X1Y5_E6BEG[6] ;
 wire \Tile_X1Y5_E6BEG[7] ;
 wire \Tile_X1Y5_E6BEG[8] ;
 wire \Tile_X1Y5_E6BEG[9] ;
 wire \Tile_X1Y5_EE4BEG[0] ;
 wire \Tile_X1Y5_EE4BEG[10] ;
 wire \Tile_X1Y5_EE4BEG[11] ;
 wire \Tile_X1Y5_EE4BEG[12] ;
 wire \Tile_X1Y5_EE4BEG[13] ;
 wire \Tile_X1Y5_EE4BEG[14] ;
 wire \Tile_X1Y5_EE4BEG[15] ;
 wire \Tile_X1Y5_EE4BEG[1] ;
 wire \Tile_X1Y5_EE4BEG[2] ;
 wire \Tile_X1Y5_EE4BEG[3] ;
 wire \Tile_X1Y5_EE4BEG[4] ;
 wire \Tile_X1Y5_EE4BEG[5] ;
 wire \Tile_X1Y5_EE4BEG[6] ;
 wire \Tile_X1Y5_EE4BEG[7] ;
 wire \Tile_X1Y5_EE4BEG[8] ;
 wire \Tile_X1Y5_EE4BEG[9] ;
 wire \Tile_X1Y5_FrameData_O[0] ;
 wire \Tile_X1Y5_FrameData_O[10] ;
 wire \Tile_X1Y5_FrameData_O[11] ;
 wire \Tile_X1Y5_FrameData_O[12] ;
 wire \Tile_X1Y5_FrameData_O[13] ;
 wire \Tile_X1Y5_FrameData_O[14] ;
 wire \Tile_X1Y5_FrameData_O[15] ;
 wire \Tile_X1Y5_FrameData_O[16] ;
 wire \Tile_X1Y5_FrameData_O[17] ;
 wire \Tile_X1Y5_FrameData_O[18] ;
 wire \Tile_X1Y5_FrameData_O[19] ;
 wire \Tile_X1Y5_FrameData_O[1] ;
 wire \Tile_X1Y5_FrameData_O[20] ;
 wire \Tile_X1Y5_FrameData_O[21] ;
 wire \Tile_X1Y5_FrameData_O[22] ;
 wire \Tile_X1Y5_FrameData_O[23] ;
 wire \Tile_X1Y5_FrameData_O[24] ;
 wire \Tile_X1Y5_FrameData_O[25] ;
 wire \Tile_X1Y5_FrameData_O[26] ;
 wire \Tile_X1Y5_FrameData_O[27] ;
 wire \Tile_X1Y5_FrameData_O[28] ;
 wire \Tile_X1Y5_FrameData_O[29] ;
 wire \Tile_X1Y5_FrameData_O[2] ;
 wire \Tile_X1Y5_FrameData_O[30] ;
 wire \Tile_X1Y5_FrameData_O[31] ;
 wire \Tile_X1Y5_FrameData_O[3] ;
 wire \Tile_X1Y5_FrameData_O[4] ;
 wire \Tile_X1Y5_FrameData_O[5] ;
 wire \Tile_X1Y5_FrameData_O[6] ;
 wire \Tile_X1Y5_FrameData_O[7] ;
 wire \Tile_X1Y5_FrameData_O[8] ;
 wire \Tile_X1Y5_FrameData_O[9] ;
 wire \Tile_X1Y5_FrameStrobe_O[0] ;
 wire \Tile_X1Y5_FrameStrobe_O[10] ;
 wire \Tile_X1Y5_FrameStrobe_O[11] ;
 wire \Tile_X1Y5_FrameStrobe_O[12] ;
 wire \Tile_X1Y5_FrameStrobe_O[13] ;
 wire \Tile_X1Y5_FrameStrobe_O[14] ;
 wire \Tile_X1Y5_FrameStrobe_O[15] ;
 wire \Tile_X1Y5_FrameStrobe_O[16] ;
 wire \Tile_X1Y5_FrameStrobe_O[17] ;
 wire \Tile_X1Y5_FrameStrobe_O[18] ;
 wire \Tile_X1Y5_FrameStrobe_O[19] ;
 wire \Tile_X1Y5_FrameStrobe_O[1] ;
 wire \Tile_X1Y5_FrameStrobe_O[2] ;
 wire \Tile_X1Y5_FrameStrobe_O[3] ;
 wire \Tile_X1Y5_FrameStrobe_O[4] ;
 wire \Tile_X1Y5_FrameStrobe_O[5] ;
 wire \Tile_X1Y5_FrameStrobe_O[6] ;
 wire \Tile_X1Y5_FrameStrobe_O[7] ;
 wire \Tile_X1Y5_FrameStrobe_O[8] ;
 wire \Tile_X1Y5_FrameStrobe_O[9] ;
 wire \Tile_X1Y5_N1BEG[0] ;
 wire \Tile_X1Y5_N1BEG[1] ;
 wire \Tile_X1Y5_N1BEG[2] ;
 wire \Tile_X1Y5_N1BEG[3] ;
 wire \Tile_X1Y5_N2BEG[0] ;
 wire \Tile_X1Y5_N2BEG[1] ;
 wire \Tile_X1Y5_N2BEG[2] ;
 wire \Tile_X1Y5_N2BEG[3] ;
 wire \Tile_X1Y5_N2BEG[4] ;
 wire \Tile_X1Y5_N2BEG[5] ;
 wire \Tile_X1Y5_N2BEG[6] ;
 wire \Tile_X1Y5_N2BEG[7] ;
 wire \Tile_X1Y5_N2BEGb[0] ;
 wire \Tile_X1Y5_N2BEGb[1] ;
 wire \Tile_X1Y5_N2BEGb[2] ;
 wire \Tile_X1Y5_N2BEGb[3] ;
 wire \Tile_X1Y5_N2BEGb[4] ;
 wire \Tile_X1Y5_N2BEGb[5] ;
 wire \Tile_X1Y5_N2BEGb[6] ;
 wire \Tile_X1Y5_N2BEGb[7] ;
 wire \Tile_X1Y5_N4BEG[0] ;
 wire \Tile_X1Y5_N4BEG[10] ;
 wire \Tile_X1Y5_N4BEG[11] ;
 wire \Tile_X1Y5_N4BEG[12] ;
 wire \Tile_X1Y5_N4BEG[13] ;
 wire \Tile_X1Y5_N4BEG[14] ;
 wire \Tile_X1Y5_N4BEG[15] ;
 wire \Tile_X1Y5_N4BEG[1] ;
 wire \Tile_X1Y5_N4BEG[2] ;
 wire \Tile_X1Y5_N4BEG[3] ;
 wire \Tile_X1Y5_N4BEG[4] ;
 wire \Tile_X1Y5_N4BEG[5] ;
 wire \Tile_X1Y5_N4BEG[6] ;
 wire \Tile_X1Y5_N4BEG[7] ;
 wire \Tile_X1Y5_N4BEG[8] ;
 wire \Tile_X1Y5_N4BEG[9] ;
 wire \Tile_X1Y5_NN4BEG[0] ;
 wire \Tile_X1Y5_NN4BEG[10] ;
 wire \Tile_X1Y5_NN4BEG[11] ;
 wire \Tile_X1Y5_NN4BEG[12] ;
 wire \Tile_X1Y5_NN4BEG[13] ;
 wire \Tile_X1Y5_NN4BEG[14] ;
 wire \Tile_X1Y5_NN4BEG[15] ;
 wire \Tile_X1Y5_NN4BEG[1] ;
 wire \Tile_X1Y5_NN4BEG[2] ;
 wire \Tile_X1Y5_NN4BEG[3] ;
 wire \Tile_X1Y5_NN4BEG[4] ;
 wire \Tile_X1Y5_NN4BEG[5] ;
 wire \Tile_X1Y5_NN4BEG[6] ;
 wire \Tile_X1Y5_NN4BEG[7] ;
 wire \Tile_X1Y5_NN4BEG[8] ;
 wire \Tile_X1Y5_NN4BEG[9] ;
 wire \Tile_X1Y5_S1BEG[0] ;
 wire \Tile_X1Y5_S1BEG[1] ;
 wire \Tile_X1Y5_S1BEG[2] ;
 wire \Tile_X1Y5_S1BEG[3] ;
 wire \Tile_X1Y5_S2BEG[0] ;
 wire \Tile_X1Y5_S2BEG[1] ;
 wire \Tile_X1Y5_S2BEG[2] ;
 wire \Tile_X1Y5_S2BEG[3] ;
 wire \Tile_X1Y5_S2BEG[4] ;
 wire \Tile_X1Y5_S2BEG[5] ;
 wire \Tile_X1Y5_S2BEG[6] ;
 wire \Tile_X1Y5_S2BEG[7] ;
 wire \Tile_X1Y5_S2BEGb[0] ;
 wire \Tile_X1Y5_S2BEGb[1] ;
 wire \Tile_X1Y5_S2BEGb[2] ;
 wire \Tile_X1Y5_S2BEGb[3] ;
 wire \Tile_X1Y5_S2BEGb[4] ;
 wire \Tile_X1Y5_S2BEGb[5] ;
 wire \Tile_X1Y5_S2BEGb[6] ;
 wire \Tile_X1Y5_S2BEGb[7] ;
 wire \Tile_X1Y5_S4BEG[0] ;
 wire \Tile_X1Y5_S4BEG[10] ;
 wire \Tile_X1Y5_S4BEG[11] ;
 wire \Tile_X1Y5_S4BEG[12] ;
 wire \Tile_X1Y5_S4BEG[13] ;
 wire \Tile_X1Y5_S4BEG[14] ;
 wire \Tile_X1Y5_S4BEG[15] ;
 wire \Tile_X1Y5_S4BEG[1] ;
 wire \Tile_X1Y5_S4BEG[2] ;
 wire \Tile_X1Y5_S4BEG[3] ;
 wire \Tile_X1Y5_S4BEG[4] ;
 wire \Tile_X1Y5_S4BEG[5] ;
 wire \Tile_X1Y5_S4BEG[6] ;
 wire \Tile_X1Y5_S4BEG[7] ;
 wire \Tile_X1Y5_S4BEG[8] ;
 wire \Tile_X1Y5_S4BEG[9] ;
 wire \Tile_X1Y5_SS4BEG[0] ;
 wire \Tile_X1Y5_SS4BEG[10] ;
 wire \Tile_X1Y5_SS4BEG[11] ;
 wire \Tile_X1Y5_SS4BEG[12] ;
 wire \Tile_X1Y5_SS4BEG[13] ;
 wire \Tile_X1Y5_SS4BEG[14] ;
 wire \Tile_X1Y5_SS4BEG[15] ;
 wire \Tile_X1Y5_SS4BEG[1] ;
 wire \Tile_X1Y5_SS4BEG[2] ;
 wire \Tile_X1Y5_SS4BEG[3] ;
 wire \Tile_X1Y5_SS4BEG[4] ;
 wire \Tile_X1Y5_SS4BEG[5] ;
 wire \Tile_X1Y5_SS4BEG[6] ;
 wire \Tile_X1Y5_SS4BEG[7] ;
 wire \Tile_X1Y5_SS4BEG[8] ;
 wire \Tile_X1Y5_SS4BEG[9] ;
 wire Tile_X1Y5_UserCLKo;
 wire \Tile_X1Y5_W1BEG[0] ;
 wire \Tile_X1Y5_W1BEG[1] ;
 wire \Tile_X1Y5_W1BEG[2] ;
 wire \Tile_X1Y5_W1BEG[3] ;
 wire \Tile_X1Y5_W2BEG[0] ;
 wire \Tile_X1Y5_W2BEG[1] ;
 wire \Tile_X1Y5_W2BEG[2] ;
 wire \Tile_X1Y5_W2BEG[3] ;
 wire \Tile_X1Y5_W2BEG[4] ;
 wire \Tile_X1Y5_W2BEG[5] ;
 wire \Tile_X1Y5_W2BEG[6] ;
 wire \Tile_X1Y5_W2BEG[7] ;
 wire \Tile_X1Y5_W2BEGb[0] ;
 wire \Tile_X1Y5_W2BEGb[1] ;
 wire \Tile_X1Y5_W2BEGb[2] ;
 wire \Tile_X1Y5_W2BEGb[3] ;
 wire \Tile_X1Y5_W2BEGb[4] ;
 wire \Tile_X1Y5_W2BEGb[5] ;
 wire \Tile_X1Y5_W2BEGb[6] ;
 wire \Tile_X1Y5_W2BEGb[7] ;
 wire \Tile_X1Y5_W6BEG[0] ;
 wire \Tile_X1Y5_W6BEG[10] ;
 wire \Tile_X1Y5_W6BEG[11] ;
 wire \Tile_X1Y5_W6BEG[1] ;
 wire \Tile_X1Y5_W6BEG[2] ;
 wire \Tile_X1Y5_W6BEG[3] ;
 wire \Tile_X1Y5_W6BEG[4] ;
 wire \Tile_X1Y5_W6BEG[5] ;
 wire \Tile_X1Y5_W6BEG[6] ;
 wire \Tile_X1Y5_W6BEG[7] ;
 wire \Tile_X1Y5_W6BEG[8] ;
 wire \Tile_X1Y5_W6BEG[9] ;
 wire \Tile_X1Y5_WW4BEG[0] ;
 wire \Tile_X1Y5_WW4BEG[10] ;
 wire \Tile_X1Y5_WW4BEG[11] ;
 wire \Tile_X1Y5_WW4BEG[12] ;
 wire \Tile_X1Y5_WW4BEG[13] ;
 wire \Tile_X1Y5_WW4BEG[14] ;
 wire \Tile_X1Y5_WW4BEG[15] ;
 wire \Tile_X1Y5_WW4BEG[1] ;
 wire \Tile_X1Y5_WW4BEG[2] ;
 wire \Tile_X1Y5_WW4BEG[3] ;
 wire \Tile_X1Y5_WW4BEG[4] ;
 wire \Tile_X1Y5_WW4BEG[5] ;
 wire \Tile_X1Y5_WW4BEG[6] ;
 wire \Tile_X1Y5_WW4BEG[7] ;
 wire \Tile_X1Y5_WW4BEG[8] ;
 wire \Tile_X1Y5_WW4BEG[9] ;
 wire Tile_X1Y6_Co;
 wire \Tile_X1Y6_E1BEG[0] ;
 wire \Tile_X1Y6_E1BEG[1] ;
 wire \Tile_X1Y6_E1BEG[2] ;
 wire \Tile_X1Y6_E1BEG[3] ;
 wire \Tile_X1Y6_E2BEG[0] ;
 wire \Tile_X1Y6_E2BEG[1] ;
 wire \Tile_X1Y6_E2BEG[2] ;
 wire \Tile_X1Y6_E2BEG[3] ;
 wire \Tile_X1Y6_E2BEG[4] ;
 wire \Tile_X1Y6_E2BEG[5] ;
 wire \Tile_X1Y6_E2BEG[6] ;
 wire \Tile_X1Y6_E2BEG[7] ;
 wire \Tile_X1Y6_E2BEGb[0] ;
 wire \Tile_X1Y6_E2BEGb[1] ;
 wire \Tile_X1Y6_E2BEGb[2] ;
 wire \Tile_X1Y6_E2BEGb[3] ;
 wire \Tile_X1Y6_E2BEGb[4] ;
 wire \Tile_X1Y6_E2BEGb[5] ;
 wire \Tile_X1Y6_E2BEGb[6] ;
 wire \Tile_X1Y6_E2BEGb[7] ;
 wire \Tile_X1Y6_E6BEG[0] ;
 wire \Tile_X1Y6_E6BEG[10] ;
 wire \Tile_X1Y6_E6BEG[11] ;
 wire \Tile_X1Y6_E6BEG[1] ;
 wire \Tile_X1Y6_E6BEG[2] ;
 wire \Tile_X1Y6_E6BEG[3] ;
 wire \Tile_X1Y6_E6BEG[4] ;
 wire \Tile_X1Y6_E6BEG[5] ;
 wire \Tile_X1Y6_E6BEG[6] ;
 wire \Tile_X1Y6_E6BEG[7] ;
 wire \Tile_X1Y6_E6BEG[8] ;
 wire \Tile_X1Y6_E6BEG[9] ;
 wire \Tile_X1Y6_EE4BEG[0] ;
 wire \Tile_X1Y6_EE4BEG[10] ;
 wire \Tile_X1Y6_EE4BEG[11] ;
 wire \Tile_X1Y6_EE4BEG[12] ;
 wire \Tile_X1Y6_EE4BEG[13] ;
 wire \Tile_X1Y6_EE4BEG[14] ;
 wire \Tile_X1Y6_EE4BEG[15] ;
 wire \Tile_X1Y6_EE4BEG[1] ;
 wire \Tile_X1Y6_EE4BEG[2] ;
 wire \Tile_X1Y6_EE4BEG[3] ;
 wire \Tile_X1Y6_EE4BEG[4] ;
 wire \Tile_X1Y6_EE4BEG[5] ;
 wire \Tile_X1Y6_EE4BEG[6] ;
 wire \Tile_X1Y6_EE4BEG[7] ;
 wire \Tile_X1Y6_EE4BEG[8] ;
 wire \Tile_X1Y6_EE4BEG[9] ;
 wire \Tile_X1Y6_FrameData_O[0] ;
 wire \Tile_X1Y6_FrameData_O[10] ;
 wire \Tile_X1Y6_FrameData_O[11] ;
 wire \Tile_X1Y6_FrameData_O[12] ;
 wire \Tile_X1Y6_FrameData_O[13] ;
 wire \Tile_X1Y6_FrameData_O[14] ;
 wire \Tile_X1Y6_FrameData_O[15] ;
 wire \Tile_X1Y6_FrameData_O[16] ;
 wire \Tile_X1Y6_FrameData_O[17] ;
 wire \Tile_X1Y6_FrameData_O[18] ;
 wire \Tile_X1Y6_FrameData_O[19] ;
 wire \Tile_X1Y6_FrameData_O[1] ;
 wire \Tile_X1Y6_FrameData_O[20] ;
 wire \Tile_X1Y6_FrameData_O[21] ;
 wire \Tile_X1Y6_FrameData_O[22] ;
 wire \Tile_X1Y6_FrameData_O[23] ;
 wire \Tile_X1Y6_FrameData_O[24] ;
 wire \Tile_X1Y6_FrameData_O[25] ;
 wire \Tile_X1Y6_FrameData_O[26] ;
 wire \Tile_X1Y6_FrameData_O[27] ;
 wire \Tile_X1Y6_FrameData_O[28] ;
 wire \Tile_X1Y6_FrameData_O[29] ;
 wire \Tile_X1Y6_FrameData_O[2] ;
 wire \Tile_X1Y6_FrameData_O[30] ;
 wire \Tile_X1Y6_FrameData_O[31] ;
 wire \Tile_X1Y6_FrameData_O[3] ;
 wire \Tile_X1Y6_FrameData_O[4] ;
 wire \Tile_X1Y6_FrameData_O[5] ;
 wire \Tile_X1Y6_FrameData_O[6] ;
 wire \Tile_X1Y6_FrameData_O[7] ;
 wire \Tile_X1Y6_FrameData_O[8] ;
 wire \Tile_X1Y6_FrameData_O[9] ;
 wire \Tile_X1Y6_FrameStrobe_O[0] ;
 wire \Tile_X1Y6_FrameStrobe_O[10] ;
 wire \Tile_X1Y6_FrameStrobe_O[11] ;
 wire \Tile_X1Y6_FrameStrobe_O[12] ;
 wire \Tile_X1Y6_FrameStrobe_O[13] ;
 wire \Tile_X1Y6_FrameStrobe_O[14] ;
 wire \Tile_X1Y6_FrameStrobe_O[15] ;
 wire \Tile_X1Y6_FrameStrobe_O[16] ;
 wire \Tile_X1Y6_FrameStrobe_O[17] ;
 wire \Tile_X1Y6_FrameStrobe_O[18] ;
 wire \Tile_X1Y6_FrameStrobe_O[19] ;
 wire \Tile_X1Y6_FrameStrobe_O[1] ;
 wire \Tile_X1Y6_FrameStrobe_O[2] ;
 wire \Tile_X1Y6_FrameStrobe_O[3] ;
 wire \Tile_X1Y6_FrameStrobe_O[4] ;
 wire \Tile_X1Y6_FrameStrobe_O[5] ;
 wire \Tile_X1Y6_FrameStrobe_O[6] ;
 wire \Tile_X1Y6_FrameStrobe_O[7] ;
 wire \Tile_X1Y6_FrameStrobe_O[8] ;
 wire \Tile_X1Y6_FrameStrobe_O[9] ;
 wire \Tile_X1Y6_N1BEG[0] ;
 wire \Tile_X1Y6_N1BEG[1] ;
 wire \Tile_X1Y6_N1BEG[2] ;
 wire \Tile_X1Y6_N1BEG[3] ;
 wire \Tile_X1Y6_N2BEG[0] ;
 wire \Tile_X1Y6_N2BEG[1] ;
 wire \Tile_X1Y6_N2BEG[2] ;
 wire \Tile_X1Y6_N2BEG[3] ;
 wire \Tile_X1Y6_N2BEG[4] ;
 wire \Tile_X1Y6_N2BEG[5] ;
 wire \Tile_X1Y6_N2BEG[6] ;
 wire \Tile_X1Y6_N2BEG[7] ;
 wire \Tile_X1Y6_N2BEGb[0] ;
 wire \Tile_X1Y6_N2BEGb[1] ;
 wire \Tile_X1Y6_N2BEGb[2] ;
 wire \Tile_X1Y6_N2BEGb[3] ;
 wire \Tile_X1Y6_N2BEGb[4] ;
 wire \Tile_X1Y6_N2BEGb[5] ;
 wire \Tile_X1Y6_N2BEGb[6] ;
 wire \Tile_X1Y6_N2BEGb[7] ;
 wire \Tile_X1Y6_N4BEG[0] ;
 wire \Tile_X1Y6_N4BEG[10] ;
 wire \Tile_X1Y6_N4BEG[11] ;
 wire \Tile_X1Y6_N4BEG[12] ;
 wire \Tile_X1Y6_N4BEG[13] ;
 wire \Tile_X1Y6_N4BEG[14] ;
 wire \Tile_X1Y6_N4BEG[15] ;
 wire \Tile_X1Y6_N4BEG[1] ;
 wire \Tile_X1Y6_N4BEG[2] ;
 wire \Tile_X1Y6_N4BEG[3] ;
 wire \Tile_X1Y6_N4BEG[4] ;
 wire \Tile_X1Y6_N4BEG[5] ;
 wire \Tile_X1Y6_N4BEG[6] ;
 wire \Tile_X1Y6_N4BEG[7] ;
 wire \Tile_X1Y6_N4BEG[8] ;
 wire \Tile_X1Y6_N4BEG[9] ;
 wire \Tile_X1Y6_NN4BEG[0] ;
 wire \Tile_X1Y6_NN4BEG[10] ;
 wire \Tile_X1Y6_NN4BEG[11] ;
 wire \Tile_X1Y6_NN4BEG[12] ;
 wire \Tile_X1Y6_NN4BEG[13] ;
 wire \Tile_X1Y6_NN4BEG[14] ;
 wire \Tile_X1Y6_NN4BEG[15] ;
 wire \Tile_X1Y6_NN4BEG[1] ;
 wire \Tile_X1Y6_NN4BEG[2] ;
 wire \Tile_X1Y6_NN4BEG[3] ;
 wire \Tile_X1Y6_NN4BEG[4] ;
 wire \Tile_X1Y6_NN4BEG[5] ;
 wire \Tile_X1Y6_NN4BEG[6] ;
 wire \Tile_X1Y6_NN4BEG[7] ;
 wire \Tile_X1Y6_NN4BEG[8] ;
 wire \Tile_X1Y6_NN4BEG[9] ;
 wire \Tile_X1Y6_S1BEG[0] ;
 wire \Tile_X1Y6_S1BEG[1] ;
 wire \Tile_X1Y6_S1BEG[2] ;
 wire \Tile_X1Y6_S1BEG[3] ;
 wire \Tile_X1Y6_S2BEG[0] ;
 wire \Tile_X1Y6_S2BEG[1] ;
 wire \Tile_X1Y6_S2BEG[2] ;
 wire \Tile_X1Y6_S2BEG[3] ;
 wire \Tile_X1Y6_S2BEG[4] ;
 wire \Tile_X1Y6_S2BEG[5] ;
 wire \Tile_X1Y6_S2BEG[6] ;
 wire \Tile_X1Y6_S2BEG[7] ;
 wire \Tile_X1Y6_S2BEGb[0] ;
 wire \Tile_X1Y6_S2BEGb[1] ;
 wire \Tile_X1Y6_S2BEGb[2] ;
 wire \Tile_X1Y6_S2BEGb[3] ;
 wire \Tile_X1Y6_S2BEGb[4] ;
 wire \Tile_X1Y6_S2BEGb[5] ;
 wire \Tile_X1Y6_S2BEGb[6] ;
 wire \Tile_X1Y6_S2BEGb[7] ;
 wire \Tile_X1Y6_S4BEG[0] ;
 wire \Tile_X1Y6_S4BEG[10] ;
 wire \Tile_X1Y6_S4BEG[11] ;
 wire \Tile_X1Y6_S4BEG[12] ;
 wire \Tile_X1Y6_S4BEG[13] ;
 wire \Tile_X1Y6_S4BEG[14] ;
 wire \Tile_X1Y6_S4BEG[15] ;
 wire \Tile_X1Y6_S4BEG[1] ;
 wire \Tile_X1Y6_S4BEG[2] ;
 wire \Tile_X1Y6_S4BEG[3] ;
 wire \Tile_X1Y6_S4BEG[4] ;
 wire \Tile_X1Y6_S4BEG[5] ;
 wire \Tile_X1Y6_S4BEG[6] ;
 wire \Tile_X1Y6_S4BEG[7] ;
 wire \Tile_X1Y6_S4BEG[8] ;
 wire \Tile_X1Y6_S4BEG[9] ;
 wire \Tile_X1Y6_SS4BEG[0] ;
 wire \Tile_X1Y6_SS4BEG[10] ;
 wire \Tile_X1Y6_SS4BEG[11] ;
 wire \Tile_X1Y6_SS4BEG[12] ;
 wire \Tile_X1Y6_SS4BEG[13] ;
 wire \Tile_X1Y6_SS4BEG[14] ;
 wire \Tile_X1Y6_SS4BEG[15] ;
 wire \Tile_X1Y6_SS4BEG[1] ;
 wire \Tile_X1Y6_SS4BEG[2] ;
 wire \Tile_X1Y6_SS4BEG[3] ;
 wire \Tile_X1Y6_SS4BEG[4] ;
 wire \Tile_X1Y6_SS4BEG[5] ;
 wire \Tile_X1Y6_SS4BEG[6] ;
 wire \Tile_X1Y6_SS4BEG[7] ;
 wire \Tile_X1Y6_SS4BEG[8] ;
 wire \Tile_X1Y6_SS4BEG[9] ;
 wire Tile_X1Y6_UserCLKo;
 wire \Tile_X1Y6_W1BEG[0] ;
 wire \Tile_X1Y6_W1BEG[1] ;
 wire \Tile_X1Y6_W1BEG[2] ;
 wire \Tile_X1Y6_W1BEG[3] ;
 wire \Tile_X1Y6_W2BEG[0] ;
 wire \Tile_X1Y6_W2BEG[1] ;
 wire \Tile_X1Y6_W2BEG[2] ;
 wire \Tile_X1Y6_W2BEG[3] ;
 wire \Tile_X1Y6_W2BEG[4] ;
 wire \Tile_X1Y6_W2BEG[5] ;
 wire \Tile_X1Y6_W2BEG[6] ;
 wire \Tile_X1Y6_W2BEG[7] ;
 wire \Tile_X1Y6_W2BEGb[0] ;
 wire \Tile_X1Y6_W2BEGb[1] ;
 wire \Tile_X1Y6_W2BEGb[2] ;
 wire \Tile_X1Y6_W2BEGb[3] ;
 wire \Tile_X1Y6_W2BEGb[4] ;
 wire \Tile_X1Y6_W2BEGb[5] ;
 wire \Tile_X1Y6_W2BEGb[6] ;
 wire \Tile_X1Y6_W2BEGb[7] ;
 wire \Tile_X1Y6_W6BEG[0] ;
 wire \Tile_X1Y6_W6BEG[10] ;
 wire \Tile_X1Y6_W6BEG[11] ;
 wire \Tile_X1Y6_W6BEG[1] ;
 wire \Tile_X1Y6_W6BEG[2] ;
 wire \Tile_X1Y6_W6BEG[3] ;
 wire \Tile_X1Y6_W6BEG[4] ;
 wire \Tile_X1Y6_W6BEG[5] ;
 wire \Tile_X1Y6_W6BEG[6] ;
 wire \Tile_X1Y6_W6BEG[7] ;
 wire \Tile_X1Y6_W6BEG[8] ;
 wire \Tile_X1Y6_W6BEG[9] ;
 wire \Tile_X1Y6_WW4BEG[0] ;
 wire \Tile_X1Y6_WW4BEG[10] ;
 wire \Tile_X1Y6_WW4BEG[11] ;
 wire \Tile_X1Y6_WW4BEG[12] ;
 wire \Tile_X1Y6_WW4BEG[13] ;
 wire \Tile_X1Y6_WW4BEG[14] ;
 wire \Tile_X1Y6_WW4BEG[15] ;
 wire \Tile_X1Y6_WW4BEG[1] ;
 wire \Tile_X1Y6_WW4BEG[2] ;
 wire \Tile_X1Y6_WW4BEG[3] ;
 wire \Tile_X1Y6_WW4BEG[4] ;
 wire \Tile_X1Y6_WW4BEG[5] ;
 wire \Tile_X1Y6_WW4BEG[6] ;
 wire \Tile_X1Y6_WW4BEG[7] ;
 wire \Tile_X1Y6_WW4BEG[8] ;
 wire \Tile_X1Y6_WW4BEG[9] ;
 wire Tile_X1Y7_Co;
 wire \Tile_X1Y7_E1BEG[0] ;
 wire \Tile_X1Y7_E1BEG[1] ;
 wire \Tile_X1Y7_E1BEG[2] ;
 wire \Tile_X1Y7_E1BEG[3] ;
 wire \Tile_X1Y7_E2BEG[0] ;
 wire \Tile_X1Y7_E2BEG[1] ;
 wire \Tile_X1Y7_E2BEG[2] ;
 wire \Tile_X1Y7_E2BEG[3] ;
 wire \Tile_X1Y7_E2BEG[4] ;
 wire \Tile_X1Y7_E2BEG[5] ;
 wire \Tile_X1Y7_E2BEG[6] ;
 wire \Tile_X1Y7_E2BEG[7] ;
 wire \Tile_X1Y7_E2BEGb[0] ;
 wire \Tile_X1Y7_E2BEGb[1] ;
 wire \Tile_X1Y7_E2BEGb[2] ;
 wire \Tile_X1Y7_E2BEGb[3] ;
 wire \Tile_X1Y7_E2BEGb[4] ;
 wire \Tile_X1Y7_E2BEGb[5] ;
 wire \Tile_X1Y7_E2BEGb[6] ;
 wire \Tile_X1Y7_E2BEGb[7] ;
 wire \Tile_X1Y7_E6BEG[0] ;
 wire \Tile_X1Y7_E6BEG[10] ;
 wire \Tile_X1Y7_E6BEG[11] ;
 wire \Tile_X1Y7_E6BEG[1] ;
 wire \Tile_X1Y7_E6BEG[2] ;
 wire \Tile_X1Y7_E6BEG[3] ;
 wire \Tile_X1Y7_E6BEG[4] ;
 wire \Tile_X1Y7_E6BEG[5] ;
 wire \Tile_X1Y7_E6BEG[6] ;
 wire \Tile_X1Y7_E6BEG[7] ;
 wire \Tile_X1Y7_E6BEG[8] ;
 wire \Tile_X1Y7_E6BEG[9] ;
 wire \Tile_X1Y7_EE4BEG[0] ;
 wire \Tile_X1Y7_EE4BEG[10] ;
 wire \Tile_X1Y7_EE4BEG[11] ;
 wire \Tile_X1Y7_EE4BEG[12] ;
 wire \Tile_X1Y7_EE4BEG[13] ;
 wire \Tile_X1Y7_EE4BEG[14] ;
 wire \Tile_X1Y7_EE4BEG[15] ;
 wire \Tile_X1Y7_EE4BEG[1] ;
 wire \Tile_X1Y7_EE4BEG[2] ;
 wire \Tile_X1Y7_EE4BEG[3] ;
 wire \Tile_X1Y7_EE4BEG[4] ;
 wire \Tile_X1Y7_EE4BEG[5] ;
 wire \Tile_X1Y7_EE4BEG[6] ;
 wire \Tile_X1Y7_EE4BEG[7] ;
 wire \Tile_X1Y7_EE4BEG[8] ;
 wire \Tile_X1Y7_EE4BEG[9] ;
 wire \Tile_X1Y7_FrameData_O[0] ;
 wire \Tile_X1Y7_FrameData_O[10] ;
 wire \Tile_X1Y7_FrameData_O[11] ;
 wire \Tile_X1Y7_FrameData_O[12] ;
 wire \Tile_X1Y7_FrameData_O[13] ;
 wire \Tile_X1Y7_FrameData_O[14] ;
 wire \Tile_X1Y7_FrameData_O[15] ;
 wire \Tile_X1Y7_FrameData_O[16] ;
 wire \Tile_X1Y7_FrameData_O[17] ;
 wire \Tile_X1Y7_FrameData_O[18] ;
 wire \Tile_X1Y7_FrameData_O[19] ;
 wire \Tile_X1Y7_FrameData_O[1] ;
 wire \Tile_X1Y7_FrameData_O[20] ;
 wire \Tile_X1Y7_FrameData_O[21] ;
 wire \Tile_X1Y7_FrameData_O[22] ;
 wire \Tile_X1Y7_FrameData_O[23] ;
 wire \Tile_X1Y7_FrameData_O[24] ;
 wire \Tile_X1Y7_FrameData_O[25] ;
 wire \Tile_X1Y7_FrameData_O[26] ;
 wire \Tile_X1Y7_FrameData_O[27] ;
 wire \Tile_X1Y7_FrameData_O[28] ;
 wire \Tile_X1Y7_FrameData_O[29] ;
 wire \Tile_X1Y7_FrameData_O[2] ;
 wire \Tile_X1Y7_FrameData_O[30] ;
 wire \Tile_X1Y7_FrameData_O[31] ;
 wire \Tile_X1Y7_FrameData_O[3] ;
 wire \Tile_X1Y7_FrameData_O[4] ;
 wire \Tile_X1Y7_FrameData_O[5] ;
 wire \Tile_X1Y7_FrameData_O[6] ;
 wire \Tile_X1Y7_FrameData_O[7] ;
 wire \Tile_X1Y7_FrameData_O[8] ;
 wire \Tile_X1Y7_FrameData_O[9] ;
 wire \Tile_X1Y7_FrameStrobe_O[0] ;
 wire \Tile_X1Y7_FrameStrobe_O[10] ;
 wire \Tile_X1Y7_FrameStrobe_O[11] ;
 wire \Tile_X1Y7_FrameStrobe_O[12] ;
 wire \Tile_X1Y7_FrameStrobe_O[13] ;
 wire \Tile_X1Y7_FrameStrobe_O[14] ;
 wire \Tile_X1Y7_FrameStrobe_O[15] ;
 wire \Tile_X1Y7_FrameStrobe_O[16] ;
 wire \Tile_X1Y7_FrameStrobe_O[17] ;
 wire \Tile_X1Y7_FrameStrobe_O[18] ;
 wire \Tile_X1Y7_FrameStrobe_O[19] ;
 wire \Tile_X1Y7_FrameStrobe_O[1] ;
 wire \Tile_X1Y7_FrameStrobe_O[2] ;
 wire \Tile_X1Y7_FrameStrobe_O[3] ;
 wire \Tile_X1Y7_FrameStrobe_O[4] ;
 wire \Tile_X1Y7_FrameStrobe_O[5] ;
 wire \Tile_X1Y7_FrameStrobe_O[6] ;
 wire \Tile_X1Y7_FrameStrobe_O[7] ;
 wire \Tile_X1Y7_FrameStrobe_O[8] ;
 wire \Tile_X1Y7_FrameStrobe_O[9] ;
 wire \Tile_X1Y7_N1BEG[0] ;
 wire \Tile_X1Y7_N1BEG[1] ;
 wire \Tile_X1Y7_N1BEG[2] ;
 wire \Tile_X1Y7_N1BEG[3] ;
 wire \Tile_X1Y7_N2BEG[0] ;
 wire \Tile_X1Y7_N2BEG[1] ;
 wire \Tile_X1Y7_N2BEG[2] ;
 wire \Tile_X1Y7_N2BEG[3] ;
 wire \Tile_X1Y7_N2BEG[4] ;
 wire \Tile_X1Y7_N2BEG[5] ;
 wire \Tile_X1Y7_N2BEG[6] ;
 wire \Tile_X1Y7_N2BEG[7] ;
 wire \Tile_X1Y7_N2BEGb[0] ;
 wire \Tile_X1Y7_N2BEGb[1] ;
 wire \Tile_X1Y7_N2BEGb[2] ;
 wire \Tile_X1Y7_N2BEGb[3] ;
 wire \Tile_X1Y7_N2BEGb[4] ;
 wire \Tile_X1Y7_N2BEGb[5] ;
 wire \Tile_X1Y7_N2BEGb[6] ;
 wire \Tile_X1Y7_N2BEGb[7] ;
 wire \Tile_X1Y7_N4BEG[0] ;
 wire \Tile_X1Y7_N4BEG[10] ;
 wire \Tile_X1Y7_N4BEG[11] ;
 wire \Tile_X1Y7_N4BEG[12] ;
 wire \Tile_X1Y7_N4BEG[13] ;
 wire \Tile_X1Y7_N4BEG[14] ;
 wire \Tile_X1Y7_N4BEG[15] ;
 wire \Tile_X1Y7_N4BEG[1] ;
 wire \Tile_X1Y7_N4BEG[2] ;
 wire \Tile_X1Y7_N4BEG[3] ;
 wire \Tile_X1Y7_N4BEG[4] ;
 wire \Tile_X1Y7_N4BEG[5] ;
 wire \Tile_X1Y7_N4BEG[6] ;
 wire \Tile_X1Y7_N4BEG[7] ;
 wire \Tile_X1Y7_N4BEG[8] ;
 wire \Tile_X1Y7_N4BEG[9] ;
 wire \Tile_X1Y7_NN4BEG[0] ;
 wire \Tile_X1Y7_NN4BEG[10] ;
 wire \Tile_X1Y7_NN4BEG[11] ;
 wire \Tile_X1Y7_NN4BEG[12] ;
 wire \Tile_X1Y7_NN4BEG[13] ;
 wire \Tile_X1Y7_NN4BEG[14] ;
 wire \Tile_X1Y7_NN4BEG[15] ;
 wire \Tile_X1Y7_NN4BEG[1] ;
 wire \Tile_X1Y7_NN4BEG[2] ;
 wire \Tile_X1Y7_NN4BEG[3] ;
 wire \Tile_X1Y7_NN4BEG[4] ;
 wire \Tile_X1Y7_NN4BEG[5] ;
 wire \Tile_X1Y7_NN4BEG[6] ;
 wire \Tile_X1Y7_NN4BEG[7] ;
 wire \Tile_X1Y7_NN4BEG[8] ;
 wire \Tile_X1Y7_NN4BEG[9] ;
 wire \Tile_X1Y7_S1BEG[0] ;
 wire \Tile_X1Y7_S1BEG[1] ;
 wire \Tile_X1Y7_S1BEG[2] ;
 wire \Tile_X1Y7_S1BEG[3] ;
 wire \Tile_X1Y7_S2BEG[0] ;
 wire \Tile_X1Y7_S2BEG[1] ;
 wire \Tile_X1Y7_S2BEG[2] ;
 wire \Tile_X1Y7_S2BEG[3] ;
 wire \Tile_X1Y7_S2BEG[4] ;
 wire \Tile_X1Y7_S2BEG[5] ;
 wire \Tile_X1Y7_S2BEG[6] ;
 wire \Tile_X1Y7_S2BEG[7] ;
 wire \Tile_X1Y7_S2BEGb[0] ;
 wire \Tile_X1Y7_S2BEGb[1] ;
 wire \Tile_X1Y7_S2BEGb[2] ;
 wire \Tile_X1Y7_S2BEGb[3] ;
 wire \Tile_X1Y7_S2BEGb[4] ;
 wire \Tile_X1Y7_S2BEGb[5] ;
 wire \Tile_X1Y7_S2BEGb[6] ;
 wire \Tile_X1Y7_S2BEGb[7] ;
 wire \Tile_X1Y7_S4BEG[0] ;
 wire \Tile_X1Y7_S4BEG[10] ;
 wire \Tile_X1Y7_S4BEG[11] ;
 wire \Tile_X1Y7_S4BEG[12] ;
 wire \Tile_X1Y7_S4BEG[13] ;
 wire \Tile_X1Y7_S4BEG[14] ;
 wire \Tile_X1Y7_S4BEG[15] ;
 wire \Tile_X1Y7_S4BEG[1] ;
 wire \Tile_X1Y7_S4BEG[2] ;
 wire \Tile_X1Y7_S4BEG[3] ;
 wire \Tile_X1Y7_S4BEG[4] ;
 wire \Tile_X1Y7_S4BEG[5] ;
 wire \Tile_X1Y7_S4BEG[6] ;
 wire \Tile_X1Y7_S4BEG[7] ;
 wire \Tile_X1Y7_S4BEG[8] ;
 wire \Tile_X1Y7_S4BEG[9] ;
 wire \Tile_X1Y7_SS4BEG[0] ;
 wire \Tile_X1Y7_SS4BEG[10] ;
 wire \Tile_X1Y7_SS4BEG[11] ;
 wire \Tile_X1Y7_SS4BEG[12] ;
 wire \Tile_X1Y7_SS4BEG[13] ;
 wire \Tile_X1Y7_SS4BEG[14] ;
 wire \Tile_X1Y7_SS4BEG[15] ;
 wire \Tile_X1Y7_SS4BEG[1] ;
 wire \Tile_X1Y7_SS4BEG[2] ;
 wire \Tile_X1Y7_SS4BEG[3] ;
 wire \Tile_X1Y7_SS4BEG[4] ;
 wire \Tile_X1Y7_SS4BEG[5] ;
 wire \Tile_X1Y7_SS4BEG[6] ;
 wire \Tile_X1Y7_SS4BEG[7] ;
 wire \Tile_X1Y7_SS4BEG[8] ;
 wire \Tile_X1Y7_SS4BEG[9] ;
 wire Tile_X1Y7_UserCLKo;
 wire \Tile_X1Y7_W1BEG[0] ;
 wire \Tile_X1Y7_W1BEG[1] ;
 wire \Tile_X1Y7_W1BEG[2] ;
 wire \Tile_X1Y7_W1BEG[3] ;
 wire \Tile_X1Y7_W2BEG[0] ;
 wire \Tile_X1Y7_W2BEG[1] ;
 wire \Tile_X1Y7_W2BEG[2] ;
 wire \Tile_X1Y7_W2BEG[3] ;
 wire \Tile_X1Y7_W2BEG[4] ;
 wire \Tile_X1Y7_W2BEG[5] ;
 wire \Tile_X1Y7_W2BEG[6] ;
 wire \Tile_X1Y7_W2BEG[7] ;
 wire \Tile_X1Y7_W2BEGb[0] ;
 wire \Tile_X1Y7_W2BEGb[1] ;
 wire \Tile_X1Y7_W2BEGb[2] ;
 wire \Tile_X1Y7_W2BEGb[3] ;
 wire \Tile_X1Y7_W2BEGb[4] ;
 wire \Tile_X1Y7_W2BEGb[5] ;
 wire \Tile_X1Y7_W2BEGb[6] ;
 wire \Tile_X1Y7_W2BEGb[7] ;
 wire \Tile_X1Y7_W6BEG[0] ;
 wire \Tile_X1Y7_W6BEG[10] ;
 wire \Tile_X1Y7_W6BEG[11] ;
 wire \Tile_X1Y7_W6BEG[1] ;
 wire \Tile_X1Y7_W6BEG[2] ;
 wire \Tile_X1Y7_W6BEG[3] ;
 wire \Tile_X1Y7_W6BEG[4] ;
 wire \Tile_X1Y7_W6BEG[5] ;
 wire \Tile_X1Y7_W6BEG[6] ;
 wire \Tile_X1Y7_W6BEG[7] ;
 wire \Tile_X1Y7_W6BEG[8] ;
 wire \Tile_X1Y7_W6BEG[9] ;
 wire \Tile_X1Y7_WW4BEG[0] ;
 wire \Tile_X1Y7_WW4BEG[10] ;
 wire \Tile_X1Y7_WW4BEG[11] ;
 wire \Tile_X1Y7_WW4BEG[12] ;
 wire \Tile_X1Y7_WW4BEG[13] ;
 wire \Tile_X1Y7_WW4BEG[14] ;
 wire \Tile_X1Y7_WW4BEG[15] ;
 wire \Tile_X1Y7_WW4BEG[1] ;
 wire \Tile_X1Y7_WW4BEG[2] ;
 wire \Tile_X1Y7_WW4BEG[3] ;
 wire \Tile_X1Y7_WW4BEG[4] ;
 wire \Tile_X1Y7_WW4BEG[5] ;
 wire \Tile_X1Y7_WW4BEG[6] ;
 wire \Tile_X1Y7_WW4BEG[7] ;
 wire \Tile_X1Y7_WW4BEG[8] ;
 wire \Tile_X1Y7_WW4BEG[9] ;
 wire Tile_X1Y8_Co;
 wire \Tile_X1Y8_E1BEG[0] ;
 wire \Tile_X1Y8_E1BEG[1] ;
 wire \Tile_X1Y8_E1BEG[2] ;
 wire \Tile_X1Y8_E1BEG[3] ;
 wire \Tile_X1Y8_E2BEG[0] ;
 wire \Tile_X1Y8_E2BEG[1] ;
 wire \Tile_X1Y8_E2BEG[2] ;
 wire \Tile_X1Y8_E2BEG[3] ;
 wire \Tile_X1Y8_E2BEG[4] ;
 wire \Tile_X1Y8_E2BEG[5] ;
 wire \Tile_X1Y8_E2BEG[6] ;
 wire \Tile_X1Y8_E2BEG[7] ;
 wire \Tile_X1Y8_E2BEGb[0] ;
 wire \Tile_X1Y8_E2BEGb[1] ;
 wire \Tile_X1Y8_E2BEGb[2] ;
 wire \Tile_X1Y8_E2BEGb[3] ;
 wire \Tile_X1Y8_E2BEGb[4] ;
 wire \Tile_X1Y8_E2BEGb[5] ;
 wire \Tile_X1Y8_E2BEGb[6] ;
 wire \Tile_X1Y8_E2BEGb[7] ;
 wire \Tile_X1Y8_E6BEG[0] ;
 wire \Tile_X1Y8_E6BEG[10] ;
 wire \Tile_X1Y8_E6BEG[11] ;
 wire \Tile_X1Y8_E6BEG[1] ;
 wire \Tile_X1Y8_E6BEG[2] ;
 wire \Tile_X1Y8_E6BEG[3] ;
 wire \Tile_X1Y8_E6BEG[4] ;
 wire \Tile_X1Y8_E6BEG[5] ;
 wire \Tile_X1Y8_E6BEG[6] ;
 wire \Tile_X1Y8_E6BEG[7] ;
 wire \Tile_X1Y8_E6BEG[8] ;
 wire \Tile_X1Y8_E6BEG[9] ;
 wire \Tile_X1Y8_EE4BEG[0] ;
 wire \Tile_X1Y8_EE4BEG[10] ;
 wire \Tile_X1Y8_EE4BEG[11] ;
 wire \Tile_X1Y8_EE4BEG[12] ;
 wire \Tile_X1Y8_EE4BEG[13] ;
 wire \Tile_X1Y8_EE4BEG[14] ;
 wire \Tile_X1Y8_EE4BEG[15] ;
 wire \Tile_X1Y8_EE4BEG[1] ;
 wire \Tile_X1Y8_EE4BEG[2] ;
 wire \Tile_X1Y8_EE4BEG[3] ;
 wire \Tile_X1Y8_EE4BEG[4] ;
 wire \Tile_X1Y8_EE4BEG[5] ;
 wire \Tile_X1Y8_EE4BEG[6] ;
 wire \Tile_X1Y8_EE4BEG[7] ;
 wire \Tile_X1Y8_EE4BEG[8] ;
 wire \Tile_X1Y8_EE4BEG[9] ;
 wire \Tile_X1Y8_FrameData_O[0] ;
 wire \Tile_X1Y8_FrameData_O[10] ;
 wire \Tile_X1Y8_FrameData_O[11] ;
 wire \Tile_X1Y8_FrameData_O[12] ;
 wire \Tile_X1Y8_FrameData_O[13] ;
 wire \Tile_X1Y8_FrameData_O[14] ;
 wire \Tile_X1Y8_FrameData_O[15] ;
 wire \Tile_X1Y8_FrameData_O[16] ;
 wire \Tile_X1Y8_FrameData_O[17] ;
 wire \Tile_X1Y8_FrameData_O[18] ;
 wire \Tile_X1Y8_FrameData_O[19] ;
 wire \Tile_X1Y8_FrameData_O[1] ;
 wire \Tile_X1Y8_FrameData_O[20] ;
 wire \Tile_X1Y8_FrameData_O[21] ;
 wire \Tile_X1Y8_FrameData_O[22] ;
 wire \Tile_X1Y8_FrameData_O[23] ;
 wire \Tile_X1Y8_FrameData_O[24] ;
 wire \Tile_X1Y8_FrameData_O[25] ;
 wire \Tile_X1Y8_FrameData_O[26] ;
 wire \Tile_X1Y8_FrameData_O[27] ;
 wire \Tile_X1Y8_FrameData_O[28] ;
 wire \Tile_X1Y8_FrameData_O[29] ;
 wire \Tile_X1Y8_FrameData_O[2] ;
 wire \Tile_X1Y8_FrameData_O[30] ;
 wire \Tile_X1Y8_FrameData_O[31] ;
 wire \Tile_X1Y8_FrameData_O[3] ;
 wire \Tile_X1Y8_FrameData_O[4] ;
 wire \Tile_X1Y8_FrameData_O[5] ;
 wire \Tile_X1Y8_FrameData_O[6] ;
 wire \Tile_X1Y8_FrameData_O[7] ;
 wire \Tile_X1Y8_FrameData_O[8] ;
 wire \Tile_X1Y8_FrameData_O[9] ;
 wire \Tile_X1Y8_FrameStrobe_O[0] ;
 wire \Tile_X1Y8_FrameStrobe_O[10] ;
 wire \Tile_X1Y8_FrameStrobe_O[11] ;
 wire \Tile_X1Y8_FrameStrobe_O[12] ;
 wire \Tile_X1Y8_FrameStrobe_O[13] ;
 wire \Tile_X1Y8_FrameStrobe_O[14] ;
 wire \Tile_X1Y8_FrameStrobe_O[15] ;
 wire \Tile_X1Y8_FrameStrobe_O[16] ;
 wire \Tile_X1Y8_FrameStrobe_O[17] ;
 wire \Tile_X1Y8_FrameStrobe_O[18] ;
 wire \Tile_X1Y8_FrameStrobe_O[19] ;
 wire \Tile_X1Y8_FrameStrobe_O[1] ;
 wire \Tile_X1Y8_FrameStrobe_O[2] ;
 wire \Tile_X1Y8_FrameStrobe_O[3] ;
 wire \Tile_X1Y8_FrameStrobe_O[4] ;
 wire \Tile_X1Y8_FrameStrobe_O[5] ;
 wire \Tile_X1Y8_FrameStrobe_O[6] ;
 wire \Tile_X1Y8_FrameStrobe_O[7] ;
 wire \Tile_X1Y8_FrameStrobe_O[8] ;
 wire \Tile_X1Y8_FrameStrobe_O[9] ;
 wire \Tile_X1Y8_N1BEG[0] ;
 wire \Tile_X1Y8_N1BEG[1] ;
 wire \Tile_X1Y8_N1BEG[2] ;
 wire \Tile_X1Y8_N1BEG[3] ;
 wire \Tile_X1Y8_N2BEG[0] ;
 wire \Tile_X1Y8_N2BEG[1] ;
 wire \Tile_X1Y8_N2BEG[2] ;
 wire \Tile_X1Y8_N2BEG[3] ;
 wire \Tile_X1Y8_N2BEG[4] ;
 wire \Tile_X1Y8_N2BEG[5] ;
 wire \Tile_X1Y8_N2BEG[6] ;
 wire \Tile_X1Y8_N2BEG[7] ;
 wire \Tile_X1Y8_N2BEGb[0] ;
 wire \Tile_X1Y8_N2BEGb[1] ;
 wire \Tile_X1Y8_N2BEGb[2] ;
 wire \Tile_X1Y8_N2BEGb[3] ;
 wire \Tile_X1Y8_N2BEGb[4] ;
 wire \Tile_X1Y8_N2BEGb[5] ;
 wire \Tile_X1Y8_N2BEGb[6] ;
 wire \Tile_X1Y8_N2BEGb[7] ;
 wire \Tile_X1Y8_N4BEG[0] ;
 wire \Tile_X1Y8_N4BEG[10] ;
 wire \Tile_X1Y8_N4BEG[11] ;
 wire \Tile_X1Y8_N4BEG[12] ;
 wire \Tile_X1Y8_N4BEG[13] ;
 wire \Tile_X1Y8_N4BEG[14] ;
 wire \Tile_X1Y8_N4BEG[15] ;
 wire \Tile_X1Y8_N4BEG[1] ;
 wire \Tile_X1Y8_N4BEG[2] ;
 wire \Tile_X1Y8_N4BEG[3] ;
 wire \Tile_X1Y8_N4BEG[4] ;
 wire \Tile_X1Y8_N4BEG[5] ;
 wire \Tile_X1Y8_N4BEG[6] ;
 wire \Tile_X1Y8_N4BEG[7] ;
 wire \Tile_X1Y8_N4BEG[8] ;
 wire \Tile_X1Y8_N4BEG[9] ;
 wire \Tile_X1Y8_NN4BEG[0] ;
 wire \Tile_X1Y8_NN4BEG[10] ;
 wire \Tile_X1Y8_NN4BEG[11] ;
 wire \Tile_X1Y8_NN4BEG[12] ;
 wire \Tile_X1Y8_NN4BEG[13] ;
 wire \Tile_X1Y8_NN4BEG[14] ;
 wire \Tile_X1Y8_NN4BEG[15] ;
 wire \Tile_X1Y8_NN4BEG[1] ;
 wire \Tile_X1Y8_NN4BEG[2] ;
 wire \Tile_X1Y8_NN4BEG[3] ;
 wire \Tile_X1Y8_NN4BEG[4] ;
 wire \Tile_X1Y8_NN4BEG[5] ;
 wire \Tile_X1Y8_NN4BEG[6] ;
 wire \Tile_X1Y8_NN4BEG[7] ;
 wire \Tile_X1Y8_NN4BEG[8] ;
 wire \Tile_X1Y8_NN4BEG[9] ;
 wire \Tile_X1Y8_S1BEG[0] ;
 wire \Tile_X1Y8_S1BEG[1] ;
 wire \Tile_X1Y8_S1BEG[2] ;
 wire \Tile_X1Y8_S1BEG[3] ;
 wire \Tile_X1Y8_S2BEG[0] ;
 wire \Tile_X1Y8_S2BEG[1] ;
 wire \Tile_X1Y8_S2BEG[2] ;
 wire \Tile_X1Y8_S2BEG[3] ;
 wire \Tile_X1Y8_S2BEG[4] ;
 wire \Tile_X1Y8_S2BEG[5] ;
 wire \Tile_X1Y8_S2BEG[6] ;
 wire \Tile_X1Y8_S2BEG[7] ;
 wire \Tile_X1Y8_S2BEGb[0] ;
 wire \Tile_X1Y8_S2BEGb[1] ;
 wire \Tile_X1Y8_S2BEGb[2] ;
 wire \Tile_X1Y8_S2BEGb[3] ;
 wire \Tile_X1Y8_S2BEGb[4] ;
 wire \Tile_X1Y8_S2BEGb[5] ;
 wire \Tile_X1Y8_S2BEGb[6] ;
 wire \Tile_X1Y8_S2BEGb[7] ;
 wire \Tile_X1Y8_S4BEG[0] ;
 wire \Tile_X1Y8_S4BEG[10] ;
 wire \Tile_X1Y8_S4BEG[11] ;
 wire \Tile_X1Y8_S4BEG[12] ;
 wire \Tile_X1Y8_S4BEG[13] ;
 wire \Tile_X1Y8_S4BEG[14] ;
 wire \Tile_X1Y8_S4BEG[15] ;
 wire \Tile_X1Y8_S4BEG[1] ;
 wire \Tile_X1Y8_S4BEG[2] ;
 wire \Tile_X1Y8_S4BEG[3] ;
 wire \Tile_X1Y8_S4BEG[4] ;
 wire \Tile_X1Y8_S4BEG[5] ;
 wire \Tile_X1Y8_S4BEG[6] ;
 wire \Tile_X1Y8_S4BEG[7] ;
 wire \Tile_X1Y8_S4BEG[8] ;
 wire \Tile_X1Y8_S4BEG[9] ;
 wire \Tile_X1Y8_SS4BEG[0] ;
 wire \Tile_X1Y8_SS4BEG[10] ;
 wire \Tile_X1Y8_SS4BEG[11] ;
 wire \Tile_X1Y8_SS4BEG[12] ;
 wire \Tile_X1Y8_SS4BEG[13] ;
 wire \Tile_X1Y8_SS4BEG[14] ;
 wire \Tile_X1Y8_SS4BEG[15] ;
 wire \Tile_X1Y8_SS4BEG[1] ;
 wire \Tile_X1Y8_SS4BEG[2] ;
 wire \Tile_X1Y8_SS4BEG[3] ;
 wire \Tile_X1Y8_SS4BEG[4] ;
 wire \Tile_X1Y8_SS4BEG[5] ;
 wire \Tile_X1Y8_SS4BEG[6] ;
 wire \Tile_X1Y8_SS4BEG[7] ;
 wire \Tile_X1Y8_SS4BEG[8] ;
 wire \Tile_X1Y8_SS4BEG[9] ;
 wire Tile_X1Y8_UserCLKo;
 wire \Tile_X1Y8_W1BEG[0] ;
 wire \Tile_X1Y8_W1BEG[1] ;
 wire \Tile_X1Y8_W1BEG[2] ;
 wire \Tile_X1Y8_W1BEG[3] ;
 wire \Tile_X1Y8_W2BEG[0] ;
 wire \Tile_X1Y8_W2BEG[1] ;
 wire \Tile_X1Y8_W2BEG[2] ;
 wire \Tile_X1Y8_W2BEG[3] ;
 wire \Tile_X1Y8_W2BEG[4] ;
 wire \Tile_X1Y8_W2BEG[5] ;
 wire \Tile_X1Y8_W2BEG[6] ;
 wire \Tile_X1Y8_W2BEG[7] ;
 wire \Tile_X1Y8_W2BEGb[0] ;
 wire \Tile_X1Y8_W2BEGb[1] ;
 wire \Tile_X1Y8_W2BEGb[2] ;
 wire \Tile_X1Y8_W2BEGb[3] ;
 wire \Tile_X1Y8_W2BEGb[4] ;
 wire \Tile_X1Y8_W2BEGb[5] ;
 wire \Tile_X1Y8_W2BEGb[6] ;
 wire \Tile_X1Y8_W2BEGb[7] ;
 wire \Tile_X1Y8_W6BEG[0] ;
 wire \Tile_X1Y8_W6BEG[10] ;
 wire \Tile_X1Y8_W6BEG[11] ;
 wire \Tile_X1Y8_W6BEG[1] ;
 wire \Tile_X1Y8_W6BEG[2] ;
 wire \Tile_X1Y8_W6BEG[3] ;
 wire \Tile_X1Y8_W6BEG[4] ;
 wire \Tile_X1Y8_W6BEG[5] ;
 wire \Tile_X1Y8_W6BEG[6] ;
 wire \Tile_X1Y8_W6BEG[7] ;
 wire \Tile_X1Y8_W6BEG[8] ;
 wire \Tile_X1Y8_W6BEG[9] ;
 wire \Tile_X1Y8_WW4BEG[0] ;
 wire \Tile_X1Y8_WW4BEG[10] ;
 wire \Tile_X1Y8_WW4BEG[11] ;
 wire \Tile_X1Y8_WW4BEG[12] ;
 wire \Tile_X1Y8_WW4BEG[13] ;
 wire \Tile_X1Y8_WW4BEG[14] ;
 wire \Tile_X1Y8_WW4BEG[15] ;
 wire \Tile_X1Y8_WW4BEG[1] ;
 wire \Tile_X1Y8_WW4BEG[2] ;
 wire \Tile_X1Y8_WW4BEG[3] ;
 wire \Tile_X1Y8_WW4BEG[4] ;
 wire \Tile_X1Y8_WW4BEG[5] ;
 wire \Tile_X1Y8_WW4BEG[6] ;
 wire \Tile_X1Y8_WW4BEG[7] ;
 wire \Tile_X1Y8_WW4BEG[8] ;
 wire \Tile_X1Y8_WW4BEG[9] ;
 wire Tile_X1Y9_Co;
 wire \Tile_X1Y9_FrameData_O[0] ;
 wire \Tile_X1Y9_FrameData_O[10] ;
 wire \Tile_X1Y9_FrameData_O[11] ;
 wire \Tile_X1Y9_FrameData_O[12] ;
 wire \Tile_X1Y9_FrameData_O[13] ;
 wire \Tile_X1Y9_FrameData_O[14] ;
 wire \Tile_X1Y9_FrameData_O[15] ;
 wire \Tile_X1Y9_FrameData_O[16] ;
 wire \Tile_X1Y9_FrameData_O[17] ;
 wire \Tile_X1Y9_FrameData_O[18] ;
 wire \Tile_X1Y9_FrameData_O[19] ;
 wire \Tile_X1Y9_FrameData_O[1] ;
 wire \Tile_X1Y9_FrameData_O[20] ;
 wire \Tile_X1Y9_FrameData_O[21] ;
 wire \Tile_X1Y9_FrameData_O[22] ;
 wire \Tile_X1Y9_FrameData_O[23] ;
 wire \Tile_X1Y9_FrameData_O[24] ;
 wire \Tile_X1Y9_FrameData_O[25] ;
 wire \Tile_X1Y9_FrameData_O[26] ;
 wire \Tile_X1Y9_FrameData_O[27] ;
 wire \Tile_X1Y9_FrameData_O[28] ;
 wire \Tile_X1Y9_FrameData_O[29] ;
 wire \Tile_X1Y9_FrameData_O[2] ;
 wire \Tile_X1Y9_FrameData_O[30] ;
 wire \Tile_X1Y9_FrameData_O[31] ;
 wire \Tile_X1Y9_FrameData_O[3] ;
 wire \Tile_X1Y9_FrameData_O[4] ;
 wire \Tile_X1Y9_FrameData_O[5] ;
 wire \Tile_X1Y9_FrameData_O[6] ;
 wire \Tile_X1Y9_FrameData_O[7] ;
 wire \Tile_X1Y9_FrameData_O[8] ;
 wire \Tile_X1Y9_FrameData_O[9] ;
 wire \Tile_X1Y9_FrameStrobe_O[0] ;
 wire \Tile_X1Y9_FrameStrobe_O[10] ;
 wire \Tile_X1Y9_FrameStrobe_O[11] ;
 wire \Tile_X1Y9_FrameStrobe_O[12] ;
 wire \Tile_X1Y9_FrameStrobe_O[13] ;
 wire \Tile_X1Y9_FrameStrobe_O[14] ;
 wire \Tile_X1Y9_FrameStrobe_O[15] ;
 wire \Tile_X1Y9_FrameStrobe_O[16] ;
 wire \Tile_X1Y9_FrameStrobe_O[17] ;
 wire \Tile_X1Y9_FrameStrobe_O[18] ;
 wire \Tile_X1Y9_FrameStrobe_O[19] ;
 wire \Tile_X1Y9_FrameStrobe_O[1] ;
 wire \Tile_X1Y9_FrameStrobe_O[2] ;
 wire \Tile_X1Y9_FrameStrobe_O[3] ;
 wire \Tile_X1Y9_FrameStrobe_O[4] ;
 wire \Tile_X1Y9_FrameStrobe_O[5] ;
 wire \Tile_X1Y9_FrameStrobe_O[6] ;
 wire \Tile_X1Y9_FrameStrobe_O[7] ;
 wire \Tile_X1Y9_FrameStrobe_O[8] ;
 wire \Tile_X1Y9_FrameStrobe_O[9] ;
 wire \Tile_X1Y9_N1BEG[0] ;
 wire \Tile_X1Y9_N1BEG[1] ;
 wire \Tile_X1Y9_N1BEG[2] ;
 wire \Tile_X1Y9_N1BEG[3] ;
 wire \Tile_X1Y9_N2BEG[0] ;
 wire \Tile_X1Y9_N2BEG[1] ;
 wire \Tile_X1Y9_N2BEG[2] ;
 wire \Tile_X1Y9_N2BEG[3] ;
 wire \Tile_X1Y9_N2BEG[4] ;
 wire \Tile_X1Y9_N2BEG[5] ;
 wire \Tile_X1Y9_N2BEG[6] ;
 wire \Tile_X1Y9_N2BEG[7] ;
 wire \Tile_X1Y9_N2BEGb[0] ;
 wire \Tile_X1Y9_N2BEGb[1] ;
 wire \Tile_X1Y9_N2BEGb[2] ;
 wire \Tile_X1Y9_N2BEGb[3] ;
 wire \Tile_X1Y9_N2BEGb[4] ;
 wire \Tile_X1Y9_N2BEGb[5] ;
 wire \Tile_X1Y9_N2BEGb[6] ;
 wire \Tile_X1Y9_N2BEGb[7] ;
 wire \Tile_X1Y9_N4BEG[0] ;
 wire \Tile_X1Y9_N4BEG[10] ;
 wire \Tile_X1Y9_N4BEG[11] ;
 wire \Tile_X1Y9_N4BEG[12] ;
 wire \Tile_X1Y9_N4BEG[13] ;
 wire \Tile_X1Y9_N4BEG[14] ;
 wire \Tile_X1Y9_N4BEG[15] ;
 wire \Tile_X1Y9_N4BEG[1] ;
 wire \Tile_X1Y9_N4BEG[2] ;
 wire \Tile_X1Y9_N4BEG[3] ;
 wire \Tile_X1Y9_N4BEG[4] ;
 wire \Tile_X1Y9_N4BEG[5] ;
 wire \Tile_X1Y9_N4BEG[6] ;
 wire \Tile_X1Y9_N4BEG[7] ;
 wire \Tile_X1Y9_N4BEG[8] ;
 wire \Tile_X1Y9_N4BEG[9] ;
 wire \Tile_X1Y9_NN4BEG[0] ;
 wire \Tile_X1Y9_NN4BEG[10] ;
 wire \Tile_X1Y9_NN4BEG[11] ;
 wire \Tile_X1Y9_NN4BEG[12] ;
 wire \Tile_X1Y9_NN4BEG[13] ;
 wire \Tile_X1Y9_NN4BEG[14] ;
 wire \Tile_X1Y9_NN4BEG[15] ;
 wire \Tile_X1Y9_NN4BEG[1] ;
 wire \Tile_X1Y9_NN4BEG[2] ;
 wire \Tile_X1Y9_NN4BEG[3] ;
 wire \Tile_X1Y9_NN4BEG[4] ;
 wire \Tile_X1Y9_NN4BEG[5] ;
 wire \Tile_X1Y9_NN4BEG[6] ;
 wire \Tile_X1Y9_NN4BEG[7] ;
 wire \Tile_X1Y9_NN4BEG[8] ;
 wire \Tile_X1Y9_NN4BEG[9] ;
 wire Tile_X1Y9_UserCLKo;
 wire \Tile_X2Y0_FrameData_O[0] ;
 wire \Tile_X2Y0_FrameData_O[10] ;
 wire \Tile_X2Y0_FrameData_O[11] ;
 wire \Tile_X2Y0_FrameData_O[12] ;
 wire \Tile_X2Y0_FrameData_O[13] ;
 wire \Tile_X2Y0_FrameData_O[14] ;
 wire \Tile_X2Y0_FrameData_O[15] ;
 wire \Tile_X2Y0_FrameData_O[16] ;
 wire \Tile_X2Y0_FrameData_O[17] ;
 wire \Tile_X2Y0_FrameData_O[18] ;
 wire \Tile_X2Y0_FrameData_O[19] ;
 wire \Tile_X2Y0_FrameData_O[1] ;
 wire \Tile_X2Y0_FrameData_O[20] ;
 wire \Tile_X2Y0_FrameData_O[21] ;
 wire \Tile_X2Y0_FrameData_O[22] ;
 wire \Tile_X2Y0_FrameData_O[23] ;
 wire \Tile_X2Y0_FrameData_O[24] ;
 wire \Tile_X2Y0_FrameData_O[25] ;
 wire \Tile_X2Y0_FrameData_O[26] ;
 wire \Tile_X2Y0_FrameData_O[27] ;
 wire \Tile_X2Y0_FrameData_O[28] ;
 wire \Tile_X2Y0_FrameData_O[29] ;
 wire \Tile_X2Y0_FrameData_O[2] ;
 wire \Tile_X2Y0_FrameData_O[30] ;
 wire \Tile_X2Y0_FrameData_O[31] ;
 wire \Tile_X2Y0_FrameData_O[3] ;
 wire \Tile_X2Y0_FrameData_O[4] ;
 wire \Tile_X2Y0_FrameData_O[5] ;
 wire \Tile_X2Y0_FrameData_O[6] ;
 wire \Tile_X2Y0_FrameData_O[7] ;
 wire \Tile_X2Y0_FrameData_O[8] ;
 wire \Tile_X2Y0_FrameData_O[9] ;
 wire \Tile_X2Y0_FrameStrobe_O[0] ;
 wire \Tile_X2Y0_FrameStrobe_O[10] ;
 wire \Tile_X2Y0_FrameStrobe_O[11] ;
 wire \Tile_X2Y0_FrameStrobe_O[12] ;
 wire \Tile_X2Y0_FrameStrobe_O[13] ;
 wire \Tile_X2Y0_FrameStrobe_O[14] ;
 wire \Tile_X2Y0_FrameStrobe_O[15] ;
 wire \Tile_X2Y0_FrameStrobe_O[16] ;
 wire \Tile_X2Y0_FrameStrobe_O[17] ;
 wire \Tile_X2Y0_FrameStrobe_O[18] ;
 wire \Tile_X2Y0_FrameStrobe_O[19] ;
 wire \Tile_X2Y0_FrameStrobe_O[1] ;
 wire \Tile_X2Y0_FrameStrobe_O[2] ;
 wire \Tile_X2Y0_FrameStrobe_O[3] ;
 wire \Tile_X2Y0_FrameStrobe_O[4] ;
 wire \Tile_X2Y0_FrameStrobe_O[5] ;
 wire \Tile_X2Y0_FrameStrobe_O[6] ;
 wire \Tile_X2Y0_FrameStrobe_O[7] ;
 wire \Tile_X2Y0_FrameStrobe_O[8] ;
 wire \Tile_X2Y0_FrameStrobe_O[9] ;
 wire \Tile_X2Y0_S1BEG[0] ;
 wire \Tile_X2Y0_S1BEG[1] ;
 wire \Tile_X2Y0_S1BEG[2] ;
 wire \Tile_X2Y0_S1BEG[3] ;
 wire \Tile_X2Y0_S2BEG[0] ;
 wire \Tile_X2Y0_S2BEG[1] ;
 wire \Tile_X2Y0_S2BEG[2] ;
 wire \Tile_X2Y0_S2BEG[3] ;
 wire \Tile_X2Y0_S2BEG[4] ;
 wire \Tile_X2Y0_S2BEG[5] ;
 wire \Tile_X2Y0_S2BEG[6] ;
 wire \Tile_X2Y0_S2BEG[7] ;
 wire \Tile_X2Y0_S2BEGb[0] ;
 wire \Tile_X2Y0_S2BEGb[1] ;
 wire \Tile_X2Y0_S2BEGb[2] ;
 wire \Tile_X2Y0_S2BEGb[3] ;
 wire \Tile_X2Y0_S2BEGb[4] ;
 wire \Tile_X2Y0_S2BEGb[5] ;
 wire \Tile_X2Y0_S2BEGb[6] ;
 wire \Tile_X2Y0_S2BEGb[7] ;
 wire \Tile_X2Y0_S4BEG[0] ;
 wire \Tile_X2Y0_S4BEG[10] ;
 wire \Tile_X2Y0_S4BEG[11] ;
 wire \Tile_X2Y0_S4BEG[12] ;
 wire \Tile_X2Y0_S4BEG[13] ;
 wire \Tile_X2Y0_S4BEG[14] ;
 wire \Tile_X2Y0_S4BEG[15] ;
 wire \Tile_X2Y0_S4BEG[1] ;
 wire \Tile_X2Y0_S4BEG[2] ;
 wire \Tile_X2Y0_S4BEG[3] ;
 wire \Tile_X2Y0_S4BEG[4] ;
 wire \Tile_X2Y0_S4BEG[5] ;
 wire \Tile_X2Y0_S4BEG[6] ;
 wire \Tile_X2Y0_S4BEG[7] ;
 wire \Tile_X2Y0_S4BEG[8] ;
 wire \Tile_X2Y0_S4BEG[9] ;
 wire \Tile_X2Y0_SS4BEG[0] ;
 wire \Tile_X2Y0_SS4BEG[10] ;
 wire \Tile_X2Y0_SS4BEG[11] ;
 wire \Tile_X2Y0_SS4BEG[12] ;
 wire \Tile_X2Y0_SS4BEG[13] ;
 wire \Tile_X2Y0_SS4BEG[14] ;
 wire \Tile_X2Y0_SS4BEG[15] ;
 wire \Tile_X2Y0_SS4BEG[1] ;
 wire \Tile_X2Y0_SS4BEG[2] ;
 wire \Tile_X2Y0_SS4BEG[3] ;
 wire \Tile_X2Y0_SS4BEG[4] ;
 wire \Tile_X2Y0_SS4BEG[5] ;
 wire \Tile_X2Y0_SS4BEG[6] ;
 wire \Tile_X2Y0_SS4BEG[7] ;
 wire \Tile_X2Y0_SS4BEG[8] ;
 wire \Tile_X2Y0_SS4BEG[9] ;
 wire Tile_X2Y0_UserCLKo;
 wire Tile_X2Y1_Co;
 wire \Tile_X2Y1_E1BEG[0] ;
 wire \Tile_X2Y1_E1BEG[1] ;
 wire \Tile_X2Y1_E1BEG[2] ;
 wire \Tile_X2Y1_E1BEG[3] ;
 wire \Tile_X2Y1_E2BEG[0] ;
 wire \Tile_X2Y1_E2BEG[1] ;
 wire \Tile_X2Y1_E2BEG[2] ;
 wire \Tile_X2Y1_E2BEG[3] ;
 wire \Tile_X2Y1_E2BEG[4] ;
 wire \Tile_X2Y1_E2BEG[5] ;
 wire \Tile_X2Y1_E2BEG[6] ;
 wire \Tile_X2Y1_E2BEG[7] ;
 wire \Tile_X2Y1_E2BEGb[0] ;
 wire \Tile_X2Y1_E2BEGb[1] ;
 wire \Tile_X2Y1_E2BEGb[2] ;
 wire \Tile_X2Y1_E2BEGb[3] ;
 wire \Tile_X2Y1_E2BEGb[4] ;
 wire \Tile_X2Y1_E2BEGb[5] ;
 wire \Tile_X2Y1_E2BEGb[6] ;
 wire \Tile_X2Y1_E2BEGb[7] ;
 wire \Tile_X2Y1_E6BEG[0] ;
 wire \Tile_X2Y1_E6BEG[10] ;
 wire \Tile_X2Y1_E6BEG[11] ;
 wire \Tile_X2Y1_E6BEG[1] ;
 wire \Tile_X2Y1_E6BEG[2] ;
 wire \Tile_X2Y1_E6BEG[3] ;
 wire \Tile_X2Y1_E6BEG[4] ;
 wire \Tile_X2Y1_E6BEG[5] ;
 wire \Tile_X2Y1_E6BEG[6] ;
 wire \Tile_X2Y1_E6BEG[7] ;
 wire \Tile_X2Y1_E6BEG[8] ;
 wire \Tile_X2Y1_E6BEG[9] ;
 wire \Tile_X2Y1_EE4BEG[0] ;
 wire \Tile_X2Y1_EE4BEG[10] ;
 wire \Tile_X2Y1_EE4BEG[11] ;
 wire \Tile_X2Y1_EE4BEG[12] ;
 wire \Tile_X2Y1_EE4BEG[13] ;
 wire \Tile_X2Y1_EE4BEG[14] ;
 wire \Tile_X2Y1_EE4BEG[15] ;
 wire \Tile_X2Y1_EE4BEG[1] ;
 wire \Tile_X2Y1_EE4BEG[2] ;
 wire \Tile_X2Y1_EE4BEG[3] ;
 wire \Tile_X2Y1_EE4BEG[4] ;
 wire \Tile_X2Y1_EE4BEG[5] ;
 wire \Tile_X2Y1_EE4BEG[6] ;
 wire \Tile_X2Y1_EE4BEG[7] ;
 wire \Tile_X2Y1_EE4BEG[8] ;
 wire \Tile_X2Y1_EE4BEG[9] ;
 wire \Tile_X2Y1_FrameData_O[0] ;
 wire \Tile_X2Y1_FrameData_O[10] ;
 wire \Tile_X2Y1_FrameData_O[11] ;
 wire \Tile_X2Y1_FrameData_O[12] ;
 wire \Tile_X2Y1_FrameData_O[13] ;
 wire \Tile_X2Y1_FrameData_O[14] ;
 wire \Tile_X2Y1_FrameData_O[15] ;
 wire \Tile_X2Y1_FrameData_O[16] ;
 wire \Tile_X2Y1_FrameData_O[17] ;
 wire \Tile_X2Y1_FrameData_O[18] ;
 wire \Tile_X2Y1_FrameData_O[19] ;
 wire \Tile_X2Y1_FrameData_O[1] ;
 wire \Tile_X2Y1_FrameData_O[20] ;
 wire \Tile_X2Y1_FrameData_O[21] ;
 wire \Tile_X2Y1_FrameData_O[22] ;
 wire \Tile_X2Y1_FrameData_O[23] ;
 wire \Tile_X2Y1_FrameData_O[24] ;
 wire \Tile_X2Y1_FrameData_O[25] ;
 wire \Tile_X2Y1_FrameData_O[26] ;
 wire \Tile_X2Y1_FrameData_O[27] ;
 wire \Tile_X2Y1_FrameData_O[28] ;
 wire \Tile_X2Y1_FrameData_O[29] ;
 wire \Tile_X2Y1_FrameData_O[2] ;
 wire \Tile_X2Y1_FrameData_O[30] ;
 wire \Tile_X2Y1_FrameData_O[31] ;
 wire \Tile_X2Y1_FrameData_O[3] ;
 wire \Tile_X2Y1_FrameData_O[4] ;
 wire \Tile_X2Y1_FrameData_O[5] ;
 wire \Tile_X2Y1_FrameData_O[6] ;
 wire \Tile_X2Y1_FrameData_O[7] ;
 wire \Tile_X2Y1_FrameData_O[8] ;
 wire \Tile_X2Y1_FrameData_O[9] ;
 wire \Tile_X2Y1_FrameStrobe_O[0] ;
 wire \Tile_X2Y1_FrameStrobe_O[10] ;
 wire \Tile_X2Y1_FrameStrobe_O[11] ;
 wire \Tile_X2Y1_FrameStrobe_O[12] ;
 wire \Tile_X2Y1_FrameStrobe_O[13] ;
 wire \Tile_X2Y1_FrameStrobe_O[14] ;
 wire \Tile_X2Y1_FrameStrobe_O[15] ;
 wire \Tile_X2Y1_FrameStrobe_O[16] ;
 wire \Tile_X2Y1_FrameStrobe_O[17] ;
 wire \Tile_X2Y1_FrameStrobe_O[18] ;
 wire \Tile_X2Y1_FrameStrobe_O[19] ;
 wire \Tile_X2Y1_FrameStrobe_O[1] ;
 wire \Tile_X2Y1_FrameStrobe_O[2] ;
 wire \Tile_X2Y1_FrameStrobe_O[3] ;
 wire \Tile_X2Y1_FrameStrobe_O[4] ;
 wire \Tile_X2Y1_FrameStrobe_O[5] ;
 wire \Tile_X2Y1_FrameStrobe_O[6] ;
 wire \Tile_X2Y1_FrameStrobe_O[7] ;
 wire \Tile_X2Y1_FrameStrobe_O[8] ;
 wire \Tile_X2Y1_FrameStrobe_O[9] ;
 wire \Tile_X2Y1_N1BEG[0] ;
 wire \Tile_X2Y1_N1BEG[1] ;
 wire \Tile_X2Y1_N1BEG[2] ;
 wire \Tile_X2Y1_N1BEG[3] ;
 wire \Tile_X2Y1_N2BEG[0] ;
 wire \Tile_X2Y1_N2BEG[1] ;
 wire \Tile_X2Y1_N2BEG[2] ;
 wire \Tile_X2Y1_N2BEG[3] ;
 wire \Tile_X2Y1_N2BEG[4] ;
 wire \Tile_X2Y1_N2BEG[5] ;
 wire \Tile_X2Y1_N2BEG[6] ;
 wire \Tile_X2Y1_N2BEG[7] ;
 wire \Tile_X2Y1_N2BEGb[0] ;
 wire \Tile_X2Y1_N2BEGb[1] ;
 wire \Tile_X2Y1_N2BEGb[2] ;
 wire \Tile_X2Y1_N2BEGb[3] ;
 wire \Tile_X2Y1_N2BEGb[4] ;
 wire \Tile_X2Y1_N2BEGb[5] ;
 wire \Tile_X2Y1_N2BEGb[6] ;
 wire \Tile_X2Y1_N2BEGb[7] ;
 wire \Tile_X2Y1_N4BEG[0] ;
 wire \Tile_X2Y1_N4BEG[10] ;
 wire \Tile_X2Y1_N4BEG[11] ;
 wire \Tile_X2Y1_N4BEG[12] ;
 wire \Tile_X2Y1_N4BEG[13] ;
 wire \Tile_X2Y1_N4BEG[14] ;
 wire \Tile_X2Y1_N4BEG[15] ;
 wire \Tile_X2Y1_N4BEG[1] ;
 wire \Tile_X2Y1_N4BEG[2] ;
 wire \Tile_X2Y1_N4BEG[3] ;
 wire \Tile_X2Y1_N4BEG[4] ;
 wire \Tile_X2Y1_N4BEG[5] ;
 wire \Tile_X2Y1_N4BEG[6] ;
 wire \Tile_X2Y1_N4BEG[7] ;
 wire \Tile_X2Y1_N4BEG[8] ;
 wire \Tile_X2Y1_N4BEG[9] ;
 wire \Tile_X2Y1_NN4BEG[0] ;
 wire \Tile_X2Y1_NN4BEG[10] ;
 wire \Tile_X2Y1_NN4BEG[11] ;
 wire \Tile_X2Y1_NN4BEG[12] ;
 wire \Tile_X2Y1_NN4BEG[13] ;
 wire \Tile_X2Y1_NN4BEG[14] ;
 wire \Tile_X2Y1_NN4BEG[15] ;
 wire \Tile_X2Y1_NN4BEG[1] ;
 wire \Tile_X2Y1_NN4BEG[2] ;
 wire \Tile_X2Y1_NN4BEG[3] ;
 wire \Tile_X2Y1_NN4BEG[4] ;
 wire \Tile_X2Y1_NN4BEG[5] ;
 wire \Tile_X2Y1_NN4BEG[6] ;
 wire \Tile_X2Y1_NN4BEG[7] ;
 wire \Tile_X2Y1_NN4BEG[8] ;
 wire \Tile_X2Y1_NN4BEG[9] ;
 wire \Tile_X2Y1_S1BEG[0] ;
 wire \Tile_X2Y1_S1BEG[1] ;
 wire \Tile_X2Y1_S1BEG[2] ;
 wire \Tile_X2Y1_S1BEG[3] ;
 wire \Tile_X2Y1_S2BEG[0] ;
 wire \Tile_X2Y1_S2BEG[1] ;
 wire \Tile_X2Y1_S2BEG[2] ;
 wire \Tile_X2Y1_S2BEG[3] ;
 wire \Tile_X2Y1_S2BEG[4] ;
 wire \Tile_X2Y1_S2BEG[5] ;
 wire \Tile_X2Y1_S2BEG[6] ;
 wire \Tile_X2Y1_S2BEG[7] ;
 wire \Tile_X2Y1_S2BEGb[0] ;
 wire \Tile_X2Y1_S2BEGb[1] ;
 wire \Tile_X2Y1_S2BEGb[2] ;
 wire \Tile_X2Y1_S2BEGb[3] ;
 wire \Tile_X2Y1_S2BEGb[4] ;
 wire \Tile_X2Y1_S2BEGb[5] ;
 wire \Tile_X2Y1_S2BEGb[6] ;
 wire \Tile_X2Y1_S2BEGb[7] ;
 wire \Tile_X2Y1_S4BEG[0] ;
 wire \Tile_X2Y1_S4BEG[10] ;
 wire \Tile_X2Y1_S4BEG[11] ;
 wire \Tile_X2Y1_S4BEG[12] ;
 wire \Tile_X2Y1_S4BEG[13] ;
 wire \Tile_X2Y1_S4BEG[14] ;
 wire \Tile_X2Y1_S4BEG[15] ;
 wire \Tile_X2Y1_S4BEG[1] ;
 wire \Tile_X2Y1_S4BEG[2] ;
 wire \Tile_X2Y1_S4BEG[3] ;
 wire \Tile_X2Y1_S4BEG[4] ;
 wire \Tile_X2Y1_S4BEG[5] ;
 wire \Tile_X2Y1_S4BEG[6] ;
 wire \Tile_X2Y1_S4BEG[7] ;
 wire \Tile_X2Y1_S4BEG[8] ;
 wire \Tile_X2Y1_S4BEG[9] ;
 wire \Tile_X2Y1_SS4BEG[0] ;
 wire \Tile_X2Y1_SS4BEG[10] ;
 wire \Tile_X2Y1_SS4BEG[11] ;
 wire \Tile_X2Y1_SS4BEG[12] ;
 wire \Tile_X2Y1_SS4BEG[13] ;
 wire \Tile_X2Y1_SS4BEG[14] ;
 wire \Tile_X2Y1_SS4BEG[15] ;
 wire \Tile_X2Y1_SS4BEG[1] ;
 wire \Tile_X2Y1_SS4BEG[2] ;
 wire \Tile_X2Y1_SS4BEG[3] ;
 wire \Tile_X2Y1_SS4BEG[4] ;
 wire \Tile_X2Y1_SS4BEG[5] ;
 wire \Tile_X2Y1_SS4BEG[6] ;
 wire \Tile_X2Y1_SS4BEG[7] ;
 wire \Tile_X2Y1_SS4BEG[8] ;
 wire \Tile_X2Y1_SS4BEG[9] ;
 wire Tile_X2Y1_UserCLKo;
 wire \Tile_X2Y1_W1BEG[0] ;
 wire \Tile_X2Y1_W1BEG[1] ;
 wire \Tile_X2Y1_W1BEG[2] ;
 wire \Tile_X2Y1_W1BEG[3] ;
 wire \Tile_X2Y1_W2BEG[0] ;
 wire \Tile_X2Y1_W2BEG[1] ;
 wire \Tile_X2Y1_W2BEG[2] ;
 wire \Tile_X2Y1_W2BEG[3] ;
 wire \Tile_X2Y1_W2BEG[4] ;
 wire \Tile_X2Y1_W2BEG[5] ;
 wire \Tile_X2Y1_W2BEG[6] ;
 wire \Tile_X2Y1_W2BEG[7] ;
 wire \Tile_X2Y1_W2BEGb[0] ;
 wire \Tile_X2Y1_W2BEGb[1] ;
 wire \Tile_X2Y1_W2BEGb[2] ;
 wire \Tile_X2Y1_W2BEGb[3] ;
 wire \Tile_X2Y1_W2BEGb[4] ;
 wire \Tile_X2Y1_W2BEGb[5] ;
 wire \Tile_X2Y1_W2BEGb[6] ;
 wire \Tile_X2Y1_W2BEGb[7] ;
 wire \Tile_X2Y1_W6BEG[0] ;
 wire \Tile_X2Y1_W6BEG[10] ;
 wire \Tile_X2Y1_W6BEG[11] ;
 wire \Tile_X2Y1_W6BEG[1] ;
 wire \Tile_X2Y1_W6BEG[2] ;
 wire \Tile_X2Y1_W6BEG[3] ;
 wire \Tile_X2Y1_W6BEG[4] ;
 wire \Tile_X2Y1_W6BEG[5] ;
 wire \Tile_X2Y1_W6BEG[6] ;
 wire \Tile_X2Y1_W6BEG[7] ;
 wire \Tile_X2Y1_W6BEG[8] ;
 wire \Tile_X2Y1_W6BEG[9] ;
 wire \Tile_X2Y1_WW4BEG[0] ;
 wire \Tile_X2Y1_WW4BEG[10] ;
 wire \Tile_X2Y1_WW4BEG[11] ;
 wire \Tile_X2Y1_WW4BEG[12] ;
 wire \Tile_X2Y1_WW4BEG[13] ;
 wire \Tile_X2Y1_WW4BEG[14] ;
 wire \Tile_X2Y1_WW4BEG[15] ;
 wire \Tile_X2Y1_WW4BEG[1] ;
 wire \Tile_X2Y1_WW4BEG[2] ;
 wire \Tile_X2Y1_WW4BEG[3] ;
 wire \Tile_X2Y1_WW4BEG[4] ;
 wire \Tile_X2Y1_WW4BEG[5] ;
 wire \Tile_X2Y1_WW4BEG[6] ;
 wire \Tile_X2Y1_WW4BEG[7] ;
 wire \Tile_X2Y1_WW4BEG[8] ;
 wire \Tile_X2Y1_WW4BEG[9] ;
 wire Tile_X2Y2_Co;
 wire \Tile_X2Y2_E1BEG[0] ;
 wire \Tile_X2Y2_E1BEG[1] ;
 wire \Tile_X2Y2_E1BEG[2] ;
 wire \Tile_X2Y2_E1BEG[3] ;
 wire \Tile_X2Y2_E2BEG[0] ;
 wire \Tile_X2Y2_E2BEG[1] ;
 wire \Tile_X2Y2_E2BEG[2] ;
 wire \Tile_X2Y2_E2BEG[3] ;
 wire \Tile_X2Y2_E2BEG[4] ;
 wire \Tile_X2Y2_E2BEG[5] ;
 wire \Tile_X2Y2_E2BEG[6] ;
 wire \Tile_X2Y2_E2BEG[7] ;
 wire \Tile_X2Y2_E2BEGb[0] ;
 wire \Tile_X2Y2_E2BEGb[1] ;
 wire \Tile_X2Y2_E2BEGb[2] ;
 wire \Tile_X2Y2_E2BEGb[3] ;
 wire \Tile_X2Y2_E2BEGb[4] ;
 wire \Tile_X2Y2_E2BEGb[5] ;
 wire \Tile_X2Y2_E2BEGb[6] ;
 wire \Tile_X2Y2_E2BEGb[7] ;
 wire \Tile_X2Y2_E6BEG[0] ;
 wire \Tile_X2Y2_E6BEG[10] ;
 wire \Tile_X2Y2_E6BEG[11] ;
 wire \Tile_X2Y2_E6BEG[1] ;
 wire \Tile_X2Y2_E6BEG[2] ;
 wire \Tile_X2Y2_E6BEG[3] ;
 wire \Tile_X2Y2_E6BEG[4] ;
 wire \Tile_X2Y2_E6BEG[5] ;
 wire \Tile_X2Y2_E6BEG[6] ;
 wire \Tile_X2Y2_E6BEG[7] ;
 wire \Tile_X2Y2_E6BEG[8] ;
 wire \Tile_X2Y2_E6BEG[9] ;
 wire \Tile_X2Y2_EE4BEG[0] ;
 wire \Tile_X2Y2_EE4BEG[10] ;
 wire \Tile_X2Y2_EE4BEG[11] ;
 wire \Tile_X2Y2_EE4BEG[12] ;
 wire \Tile_X2Y2_EE4BEG[13] ;
 wire \Tile_X2Y2_EE4BEG[14] ;
 wire \Tile_X2Y2_EE4BEG[15] ;
 wire \Tile_X2Y2_EE4BEG[1] ;
 wire \Tile_X2Y2_EE4BEG[2] ;
 wire \Tile_X2Y2_EE4BEG[3] ;
 wire \Tile_X2Y2_EE4BEG[4] ;
 wire \Tile_X2Y2_EE4BEG[5] ;
 wire \Tile_X2Y2_EE4BEG[6] ;
 wire \Tile_X2Y2_EE4BEG[7] ;
 wire \Tile_X2Y2_EE4BEG[8] ;
 wire \Tile_X2Y2_EE4BEG[9] ;
 wire \Tile_X2Y2_FrameData_O[0] ;
 wire \Tile_X2Y2_FrameData_O[10] ;
 wire \Tile_X2Y2_FrameData_O[11] ;
 wire \Tile_X2Y2_FrameData_O[12] ;
 wire \Tile_X2Y2_FrameData_O[13] ;
 wire \Tile_X2Y2_FrameData_O[14] ;
 wire \Tile_X2Y2_FrameData_O[15] ;
 wire \Tile_X2Y2_FrameData_O[16] ;
 wire \Tile_X2Y2_FrameData_O[17] ;
 wire \Tile_X2Y2_FrameData_O[18] ;
 wire \Tile_X2Y2_FrameData_O[19] ;
 wire \Tile_X2Y2_FrameData_O[1] ;
 wire \Tile_X2Y2_FrameData_O[20] ;
 wire \Tile_X2Y2_FrameData_O[21] ;
 wire \Tile_X2Y2_FrameData_O[22] ;
 wire \Tile_X2Y2_FrameData_O[23] ;
 wire \Tile_X2Y2_FrameData_O[24] ;
 wire \Tile_X2Y2_FrameData_O[25] ;
 wire \Tile_X2Y2_FrameData_O[26] ;
 wire \Tile_X2Y2_FrameData_O[27] ;
 wire \Tile_X2Y2_FrameData_O[28] ;
 wire \Tile_X2Y2_FrameData_O[29] ;
 wire \Tile_X2Y2_FrameData_O[2] ;
 wire \Tile_X2Y2_FrameData_O[30] ;
 wire \Tile_X2Y2_FrameData_O[31] ;
 wire \Tile_X2Y2_FrameData_O[3] ;
 wire \Tile_X2Y2_FrameData_O[4] ;
 wire \Tile_X2Y2_FrameData_O[5] ;
 wire \Tile_X2Y2_FrameData_O[6] ;
 wire \Tile_X2Y2_FrameData_O[7] ;
 wire \Tile_X2Y2_FrameData_O[8] ;
 wire \Tile_X2Y2_FrameData_O[9] ;
 wire \Tile_X2Y2_FrameStrobe_O[0] ;
 wire \Tile_X2Y2_FrameStrobe_O[10] ;
 wire \Tile_X2Y2_FrameStrobe_O[11] ;
 wire \Tile_X2Y2_FrameStrobe_O[12] ;
 wire \Tile_X2Y2_FrameStrobe_O[13] ;
 wire \Tile_X2Y2_FrameStrobe_O[14] ;
 wire \Tile_X2Y2_FrameStrobe_O[15] ;
 wire \Tile_X2Y2_FrameStrobe_O[16] ;
 wire \Tile_X2Y2_FrameStrobe_O[17] ;
 wire \Tile_X2Y2_FrameStrobe_O[18] ;
 wire \Tile_X2Y2_FrameStrobe_O[19] ;
 wire \Tile_X2Y2_FrameStrobe_O[1] ;
 wire \Tile_X2Y2_FrameStrobe_O[2] ;
 wire \Tile_X2Y2_FrameStrobe_O[3] ;
 wire \Tile_X2Y2_FrameStrobe_O[4] ;
 wire \Tile_X2Y2_FrameStrobe_O[5] ;
 wire \Tile_X2Y2_FrameStrobe_O[6] ;
 wire \Tile_X2Y2_FrameStrobe_O[7] ;
 wire \Tile_X2Y2_FrameStrobe_O[8] ;
 wire \Tile_X2Y2_FrameStrobe_O[9] ;
 wire \Tile_X2Y2_N1BEG[0] ;
 wire \Tile_X2Y2_N1BEG[1] ;
 wire \Tile_X2Y2_N1BEG[2] ;
 wire \Tile_X2Y2_N1BEG[3] ;
 wire \Tile_X2Y2_N2BEG[0] ;
 wire \Tile_X2Y2_N2BEG[1] ;
 wire \Tile_X2Y2_N2BEG[2] ;
 wire \Tile_X2Y2_N2BEG[3] ;
 wire \Tile_X2Y2_N2BEG[4] ;
 wire \Tile_X2Y2_N2BEG[5] ;
 wire \Tile_X2Y2_N2BEG[6] ;
 wire \Tile_X2Y2_N2BEG[7] ;
 wire \Tile_X2Y2_N2BEGb[0] ;
 wire \Tile_X2Y2_N2BEGb[1] ;
 wire \Tile_X2Y2_N2BEGb[2] ;
 wire \Tile_X2Y2_N2BEGb[3] ;
 wire \Tile_X2Y2_N2BEGb[4] ;
 wire \Tile_X2Y2_N2BEGb[5] ;
 wire \Tile_X2Y2_N2BEGb[6] ;
 wire \Tile_X2Y2_N2BEGb[7] ;
 wire \Tile_X2Y2_N4BEG[0] ;
 wire \Tile_X2Y2_N4BEG[10] ;
 wire \Tile_X2Y2_N4BEG[11] ;
 wire \Tile_X2Y2_N4BEG[12] ;
 wire \Tile_X2Y2_N4BEG[13] ;
 wire \Tile_X2Y2_N4BEG[14] ;
 wire \Tile_X2Y2_N4BEG[15] ;
 wire \Tile_X2Y2_N4BEG[1] ;
 wire \Tile_X2Y2_N4BEG[2] ;
 wire \Tile_X2Y2_N4BEG[3] ;
 wire \Tile_X2Y2_N4BEG[4] ;
 wire \Tile_X2Y2_N4BEG[5] ;
 wire \Tile_X2Y2_N4BEG[6] ;
 wire \Tile_X2Y2_N4BEG[7] ;
 wire \Tile_X2Y2_N4BEG[8] ;
 wire \Tile_X2Y2_N4BEG[9] ;
 wire \Tile_X2Y2_NN4BEG[0] ;
 wire \Tile_X2Y2_NN4BEG[10] ;
 wire \Tile_X2Y2_NN4BEG[11] ;
 wire \Tile_X2Y2_NN4BEG[12] ;
 wire \Tile_X2Y2_NN4BEG[13] ;
 wire \Tile_X2Y2_NN4BEG[14] ;
 wire \Tile_X2Y2_NN4BEG[15] ;
 wire \Tile_X2Y2_NN4BEG[1] ;
 wire \Tile_X2Y2_NN4BEG[2] ;
 wire \Tile_X2Y2_NN4BEG[3] ;
 wire \Tile_X2Y2_NN4BEG[4] ;
 wire \Tile_X2Y2_NN4BEG[5] ;
 wire \Tile_X2Y2_NN4BEG[6] ;
 wire \Tile_X2Y2_NN4BEG[7] ;
 wire \Tile_X2Y2_NN4BEG[8] ;
 wire \Tile_X2Y2_NN4BEG[9] ;
 wire \Tile_X2Y2_S1BEG[0] ;
 wire \Tile_X2Y2_S1BEG[1] ;
 wire \Tile_X2Y2_S1BEG[2] ;
 wire \Tile_X2Y2_S1BEG[3] ;
 wire \Tile_X2Y2_S2BEG[0] ;
 wire \Tile_X2Y2_S2BEG[1] ;
 wire \Tile_X2Y2_S2BEG[2] ;
 wire \Tile_X2Y2_S2BEG[3] ;
 wire \Tile_X2Y2_S2BEG[4] ;
 wire \Tile_X2Y2_S2BEG[5] ;
 wire \Tile_X2Y2_S2BEG[6] ;
 wire \Tile_X2Y2_S2BEG[7] ;
 wire \Tile_X2Y2_S2BEGb[0] ;
 wire \Tile_X2Y2_S2BEGb[1] ;
 wire \Tile_X2Y2_S2BEGb[2] ;
 wire \Tile_X2Y2_S2BEGb[3] ;
 wire \Tile_X2Y2_S2BEGb[4] ;
 wire \Tile_X2Y2_S2BEGb[5] ;
 wire \Tile_X2Y2_S2BEGb[6] ;
 wire \Tile_X2Y2_S2BEGb[7] ;
 wire \Tile_X2Y2_S4BEG[0] ;
 wire \Tile_X2Y2_S4BEG[10] ;
 wire \Tile_X2Y2_S4BEG[11] ;
 wire \Tile_X2Y2_S4BEG[12] ;
 wire \Tile_X2Y2_S4BEG[13] ;
 wire \Tile_X2Y2_S4BEG[14] ;
 wire \Tile_X2Y2_S4BEG[15] ;
 wire \Tile_X2Y2_S4BEG[1] ;
 wire \Tile_X2Y2_S4BEG[2] ;
 wire \Tile_X2Y2_S4BEG[3] ;
 wire \Tile_X2Y2_S4BEG[4] ;
 wire \Tile_X2Y2_S4BEG[5] ;
 wire \Tile_X2Y2_S4BEG[6] ;
 wire \Tile_X2Y2_S4BEG[7] ;
 wire \Tile_X2Y2_S4BEG[8] ;
 wire \Tile_X2Y2_S4BEG[9] ;
 wire \Tile_X2Y2_SS4BEG[0] ;
 wire \Tile_X2Y2_SS4BEG[10] ;
 wire \Tile_X2Y2_SS4BEG[11] ;
 wire \Tile_X2Y2_SS4BEG[12] ;
 wire \Tile_X2Y2_SS4BEG[13] ;
 wire \Tile_X2Y2_SS4BEG[14] ;
 wire \Tile_X2Y2_SS4BEG[15] ;
 wire \Tile_X2Y2_SS4BEG[1] ;
 wire \Tile_X2Y2_SS4BEG[2] ;
 wire \Tile_X2Y2_SS4BEG[3] ;
 wire \Tile_X2Y2_SS4BEG[4] ;
 wire \Tile_X2Y2_SS4BEG[5] ;
 wire \Tile_X2Y2_SS4BEG[6] ;
 wire \Tile_X2Y2_SS4BEG[7] ;
 wire \Tile_X2Y2_SS4BEG[8] ;
 wire \Tile_X2Y2_SS4BEG[9] ;
 wire Tile_X2Y2_UserCLKo;
 wire \Tile_X2Y2_W1BEG[0] ;
 wire \Tile_X2Y2_W1BEG[1] ;
 wire \Tile_X2Y2_W1BEG[2] ;
 wire \Tile_X2Y2_W1BEG[3] ;
 wire \Tile_X2Y2_W2BEG[0] ;
 wire \Tile_X2Y2_W2BEG[1] ;
 wire \Tile_X2Y2_W2BEG[2] ;
 wire \Tile_X2Y2_W2BEG[3] ;
 wire \Tile_X2Y2_W2BEG[4] ;
 wire \Tile_X2Y2_W2BEG[5] ;
 wire \Tile_X2Y2_W2BEG[6] ;
 wire \Tile_X2Y2_W2BEG[7] ;
 wire \Tile_X2Y2_W2BEGb[0] ;
 wire \Tile_X2Y2_W2BEGb[1] ;
 wire \Tile_X2Y2_W2BEGb[2] ;
 wire \Tile_X2Y2_W2BEGb[3] ;
 wire \Tile_X2Y2_W2BEGb[4] ;
 wire \Tile_X2Y2_W2BEGb[5] ;
 wire \Tile_X2Y2_W2BEGb[6] ;
 wire \Tile_X2Y2_W2BEGb[7] ;
 wire \Tile_X2Y2_W6BEG[0] ;
 wire \Tile_X2Y2_W6BEG[10] ;
 wire \Tile_X2Y2_W6BEG[11] ;
 wire \Tile_X2Y2_W6BEG[1] ;
 wire \Tile_X2Y2_W6BEG[2] ;
 wire \Tile_X2Y2_W6BEG[3] ;
 wire \Tile_X2Y2_W6BEG[4] ;
 wire \Tile_X2Y2_W6BEG[5] ;
 wire \Tile_X2Y2_W6BEG[6] ;
 wire \Tile_X2Y2_W6BEG[7] ;
 wire \Tile_X2Y2_W6BEG[8] ;
 wire \Tile_X2Y2_W6BEG[9] ;
 wire \Tile_X2Y2_WW4BEG[0] ;
 wire \Tile_X2Y2_WW4BEG[10] ;
 wire \Tile_X2Y2_WW4BEG[11] ;
 wire \Tile_X2Y2_WW4BEG[12] ;
 wire \Tile_X2Y2_WW4BEG[13] ;
 wire \Tile_X2Y2_WW4BEG[14] ;
 wire \Tile_X2Y2_WW4BEG[15] ;
 wire \Tile_X2Y2_WW4BEG[1] ;
 wire \Tile_X2Y2_WW4BEG[2] ;
 wire \Tile_X2Y2_WW4BEG[3] ;
 wire \Tile_X2Y2_WW4BEG[4] ;
 wire \Tile_X2Y2_WW4BEG[5] ;
 wire \Tile_X2Y2_WW4BEG[6] ;
 wire \Tile_X2Y2_WW4BEG[7] ;
 wire \Tile_X2Y2_WW4BEG[8] ;
 wire \Tile_X2Y2_WW4BEG[9] ;
 wire Tile_X2Y3_Co;
 wire \Tile_X2Y3_E1BEG[0] ;
 wire \Tile_X2Y3_E1BEG[1] ;
 wire \Tile_X2Y3_E1BEG[2] ;
 wire \Tile_X2Y3_E1BEG[3] ;
 wire \Tile_X2Y3_E2BEG[0] ;
 wire \Tile_X2Y3_E2BEG[1] ;
 wire \Tile_X2Y3_E2BEG[2] ;
 wire \Tile_X2Y3_E2BEG[3] ;
 wire \Tile_X2Y3_E2BEG[4] ;
 wire \Tile_X2Y3_E2BEG[5] ;
 wire \Tile_X2Y3_E2BEG[6] ;
 wire \Tile_X2Y3_E2BEG[7] ;
 wire \Tile_X2Y3_E2BEGb[0] ;
 wire \Tile_X2Y3_E2BEGb[1] ;
 wire \Tile_X2Y3_E2BEGb[2] ;
 wire \Tile_X2Y3_E2BEGb[3] ;
 wire \Tile_X2Y3_E2BEGb[4] ;
 wire \Tile_X2Y3_E2BEGb[5] ;
 wire \Tile_X2Y3_E2BEGb[6] ;
 wire \Tile_X2Y3_E2BEGb[7] ;
 wire \Tile_X2Y3_E6BEG[0] ;
 wire \Tile_X2Y3_E6BEG[10] ;
 wire \Tile_X2Y3_E6BEG[11] ;
 wire \Tile_X2Y3_E6BEG[1] ;
 wire \Tile_X2Y3_E6BEG[2] ;
 wire \Tile_X2Y3_E6BEG[3] ;
 wire \Tile_X2Y3_E6BEG[4] ;
 wire \Tile_X2Y3_E6BEG[5] ;
 wire \Tile_X2Y3_E6BEG[6] ;
 wire \Tile_X2Y3_E6BEG[7] ;
 wire \Tile_X2Y3_E6BEG[8] ;
 wire \Tile_X2Y3_E6BEG[9] ;
 wire \Tile_X2Y3_EE4BEG[0] ;
 wire \Tile_X2Y3_EE4BEG[10] ;
 wire \Tile_X2Y3_EE4BEG[11] ;
 wire \Tile_X2Y3_EE4BEG[12] ;
 wire \Tile_X2Y3_EE4BEG[13] ;
 wire \Tile_X2Y3_EE4BEG[14] ;
 wire \Tile_X2Y3_EE4BEG[15] ;
 wire \Tile_X2Y3_EE4BEG[1] ;
 wire \Tile_X2Y3_EE4BEG[2] ;
 wire \Tile_X2Y3_EE4BEG[3] ;
 wire \Tile_X2Y3_EE4BEG[4] ;
 wire \Tile_X2Y3_EE4BEG[5] ;
 wire \Tile_X2Y3_EE4BEG[6] ;
 wire \Tile_X2Y3_EE4BEG[7] ;
 wire \Tile_X2Y3_EE4BEG[8] ;
 wire \Tile_X2Y3_EE4BEG[9] ;
 wire \Tile_X2Y3_FrameData_O[0] ;
 wire \Tile_X2Y3_FrameData_O[10] ;
 wire \Tile_X2Y3_FrameData_O[11] ;
 wire \Tile_X2Y3_FrameData_O[12] ;
 wire \Tile_X2Y3_FrameData_O[13] ;
 wire \Tile_X2Y3_FrameData_O[14] ;
 wire \Tile_X2Y3_FrameData_O[15] ;
 wire \Tile_X2Y3_FrameData_O[16] ;
 wire \Tile_X2Y3_FrameData_O[17] ;
 wire \Tile_X2Y3_FrameData_O[18] ;
 wire \Tile_X2Y3_FrameData_O[19] ;
 wire \Tile_X2Y3_FrameData_O[1] ;
 wire \Tile_X2Y3_FrameData_O[20] ;
 wire \Tile_X2Y3_FrameData_O[21] ;
 wire \Tile_X2Y3_FrameData_O[22] ;
 wire \Tile_X2Y3_FrameData_O[23] ;
 wire \Tile_X2Y3_FrameData_O[24] ;
 wire \Tile_X2Y3_FrameData_O[25] ;
 wire \Tile_X2Y3_FrameData_O[26] ;
 wire \Tile_X2Y3_FrameData_O[27] ;
 wire \Tile_X2Y3_FrameData_O[28] ;
 wire \Tile_X2Y3_FrameData_O[29] ;
 wire \Tile_X2Y3_FrameData_O[2] ;
 wire \Tile_X2Y3_FrameData_O[30] ;
 wire \Tile_X2Y3_FrameData_O[31] ;
 wire \Tile_X2Y3_FrameData_O[3] ;
 wire \Tile_X2Y3_FrameData_O[4] ;
 wire \Tile_X2Y3_FrameData_O[5] ;
 wire \Tile_X2Y3_FrameData_O[6] ;
 wire \Tile_X2Y3_FrameData_O[7] ;
 wire \Tile_X2Y3_FrameData_O[8] ;
 wire \Tile_X2Y3_FrameData_O[9] ;
 wire \Tile_X2Y3_FrameStrobe_O[0] ;
 wire \Tile_X2Y3_FrameStrobe_O[10] ;
 wire \Tile_X2Y3_FrameStrobe_O[11] ;
 wire \Tile_X2Y3_FrameStrobe_O[12] ;
 wire \Tile_X2Y3_FrameStrobe_O[13] ;
 wire \Tile_X2Y3_FrameStrobe_O[14] ;
 wire \Tile_X2Y3_FrameStrobe_O[15] ;
 wire \Tile_X2Y3_FrameStrobe_O[16] ;
 wire \Tile_X2Y3_FrameStrobe_O[17] ;
 wire \Tile_X2Y3_FrameStrobe_O[18] ;
 wire \Tile_X2Y3_FrameStrobe_O[19] ;
 wire \Tile_X2Y3_FrameStrobe_O[1] ;
 wire \Tile_X2Y3_FrameStrobe_O[2] ;
 wire \Tile_X2Y3_FrameStrobe_O[3] ;
 wire \Tile_X2Y3_FrameStrobe_O[4] ;
 wire \Tile_X2Y3_FrameStrobe_O[5] ;
 wire \Tile_X2Y3_FrameStrobe_O[6] ;
 wire \Tile_X2Y3_FrameStrobe_O[7] ;
 wire \Tile_X2Y3_FrameStrobe_O[8] ;
 wire \Tile_X2Y3_FrameStrobe_O[9] ;
 wire \Tile_X2Y3_N1BEG[0] ;
 wire \Tile_X2Y3_N1BEG[1] ;
 wire \Tile_X2Y3_N1BEG[2] ;
 wire \Tile_X2Y3_N1BEG[3] ;
 wire \Tile_X2Y3_N2BEG[0] ;
 wire \Tile_X2Y3_N2BEG[1] ;
 wire \Tile_X2Y3_N2BEG[2] ;
 wire \Tile_X2Y3_N2BEG[3] ;
 wire \Tile_X2Y3_N2BEG[4] ;
 wire \Tile_X2Y3_N2BEG[5] ;
 wire \Tile_X2Y3_N2BEG[6] ;
 wire \Tile_X2Y3_N2BEG[7] ;
 wire \Tile_X2Y3_N2BEGb[0] ;
 wire \Tile_X2Y3_N2BEGb[1] ;
 wire \Tile_X2Y3_N2BEGb[2] ;
 wire \Tile_X2Y3_N2BEGb[3] ;
 wire \Tile_X2Y3_N2BEGb[4] ;
 wire \Tile_X2Y3_N2BEGb[5] ;
 wire \Tile_X2Y3_N2BEGb[6] ;
 wire \Tile_X2Y3_N2BEGb[7] ;
 wire \Tile_X2Y3_N4BEG[0] ;
 wire \Tile_X2Y3_N4BEG[10] ;
 wire \Tile_X2Y3_N4BEG[11] ;
 wire \Tile_X2Y3_N4BEG[12] ;
 wire \Tile_X2Y3_N4BEG[13] ;
 wire \Tile_X2Y3_N4BEG[14] ;
 wire \Tile_X2Y3_N4BEG[15] ;
 wire \Tile_X2Y3_N4BEG[1] ;
 wire \Tile_X2Y3_N4BEG[2] ;
 wire \Tile_X2Y3_N4BEG[3] ;
 wire \Tile_X2Y3_N4BEG[4] ;
 wire \Tile_X2Y3_N4BEG[5] ;
 wire \Tile_X2Y3_N4BEG[6] ;
 wire \Tile_X2Y3_N4BEG[7] ;
 wire \Tile_X2Y3_N4BEG[8] ;
 wire \Tile_X2Y3_N4BEG[9] ;
 wire \Tile_X2Y3_NN4BEG[0] ;
 wire \Tile_X2Y3_NN4BEG[10] ;
 wire \Tile_X2Y3_NN4BEG[11] ;
 wire \Tile_X2Y3_NN4BEG[12] ;
 wire \Tile_X2Y3_NN4BEG[13] ;
 wire \Tile_X2Y3_NN4BEG[14] ;
 wire \Tile_X2Y3_NN4BEG[15] ;
 wire \Tile_X2Y3_NN4BEG[1] ;
 wire \Tile_X2Y3_NN4BEG[2] ;
 wire \Tile_X2Y3_NN4BEG[3] ;
 wire \Tile_X2Y3_NN4BEG[4] ;
 wire \Tile_X2Y3_NN4BEG[5] ;
 wire \Tile_X2Y3_NN4BEG[6] ;
 wire \Tile_X2Y3_NN4BEG[7] ;
 wire \Tile_X2Y3_NN4BEG[8] ;
 wire \Tile_X2Y3_NN4BEG[9] ;
 wire \Tile_X2Y3_S1BEG[0] ;
 wire \Tile_X2Y3_S1BEG[1] ;
 wire \Tile_X2Y3_S1BEG[2] ;
 wire \Tile_X2Y3_S1BEG[3] ;
 wire \Tile_X2Y3_S2BEG[0] ;
 wire \Tile_X2Y3_S2BEG[1] ;
 wire \Tile_X2Y3_S2BEG[2] ;
 wire \Tile_X2Y3_S2BEG[3] ;
 wire \Tile_X2Y3_S2BEG[4] ;
 wire \Tile_X2Y3_S2BEG[5] ;
 wire \Tile_X2Y3_S2BEG[6] ;
 wire \Tile_X2Y3_S2BEG[7] ;
 wire \Tile_X2Y3_S2BEGb[0] ;
 wire \Tile_X2Y3_S2BEGb[1] ;
 wire \Tile_X2Y3_S2BEGb[2] ;
 wire \Tile_X2Y3_S2BEGb[3] ;
 wire \Tile_X2Y3_S2BEGb[4] ;
 wire \Tile_X2Y3_S2BEGb[5] ;
 wire \Tile_X2Y3_S2BEGb[6] ;
 wire \Tile_X2Y3_S2BEGb[7] ;
 wire \Tile_X2Y3_S4BEG[0] ;
 wire \Tile_X2Y3_S4BEG[10] ;
 wire \Tile_X2Y3_S4BEG[11] ;
 wire \Tile_X2Y3_S4BEG[12] ;
 wire \Tile_X2Y3_S4BEG[13] ;
 wire \Tile_X2Y3_S4BEG[14] ;
 wire \Tile_X2Y3_S4BEG[15] ;
 wire \Tile_X2Y3_S4BEG[1] ;
 wire \Tile_X2Y3_S4BEG[2] ;
 wire \Tile_X2Y3_S4BEG[3] ;
 wire \Tile_X2Y3_S4BEG[4] ;
 wire \Tile_X2Y3_S4BEG[5] ;
 wire \Tile_X2Y3_S4BEG[6] ;
 wire \Tile_X2Y3_S4BEG[7] ;
 wire \Tile_X2Y3_S4BEG[8] ;
 wire \Tile_X2Y3_S4BEG[9] ;
 wire \Tile_X2Y3_SS4BEG[0] ;
 wire \Tile_X2Y3_SS4BEG[10] ;
 wire \Tile_X2Y3_SS4BEG[11] ;
 wire \Tile_X2Y3_SS4BEG[12] ;
 wire \Tile_X2Y3_SS4BEG[13] ;
 wire \Tile_X2Y3_SS4BEG[14] ;
 wire \Tile_X2Y3_SS4BEG[15] ;
 wire \Tile_X2Y3_SS4BEG[1] ;
 wire \Tile_X2Y3_SS4BEG[2] ;
 wire \Tile_X2Y3_SS4BEG[3] ;
 wire \Tile_X2Y3_SS4BEG[4] ;
 wire \Tile_X2Y3_SS4BEG[5] ;
 wire \Tile_X2Y3_SS4BEG[6] ;
 wire \Tile_X2Y3_SS4BEG[7] ;
 wire \Tile_X2Y3_SS4BEG[8] ;
 wire \Tile_X2Y3_SS4BEG[9] ;
 wire Tile_X2Y3_UserCLKo;
 wire \Tile_X2Y3_W1BEG[0] ;
 wire \Tile_X2Y3_W1BEG[1] ;
 wire \Tile_X2Y3_W1BEG[2] ;
 wire \Tile_X2Y3_W1BEG[3] ;
 wire \Tile_X2Y3_W2BEG[0] ;
 wire \Tile_X2Y3_W2BEG[1] ;
 wire \Tile_X2Y3_W2BEG[2] ;
 wire \Tile_X2Y3_W2BEG[3] ;
 wire \Tile_X2Y3_W2BEG[4] ;
 wire \Tile_X2Y3_W2BEG[5] ;
 wire \Tile_X2Y3_W2BEG[6] ;
 wire \Tile_X2Y3_W2BEG[7] ;
 wire \Tile_X2Y3_W2BEGb[0] ;
 wire \Tile_X2Y3_W2BEGb[1] ;
 wire \Tile_X2Y3_W2BEGb[2] ;
 wire \Tile_X2Y3_W2BEGb[3] ;
 wire \Tile_X2Y3_W2BEGb[4] ;
 wire \Tile_X2Y3_W2BEGb[5] ;
 wire \Tile_X2Y3_W2BEGb[6] ;
 wire \Tile_X2Y3_W2BEGb[7] ;
 wire \Tile_X2Y3_W6BEG[0] ;
 wire \Tile_X2Y3_W6BEG[10] ;
 wire \Tile_X2Y3_W6BEG[11] ;
 wire \Tile_X2Y3_W6BEG[1] ;
 wire \Tile_X2Y3_W6BEG[2] ;
 wire \Tile_X2Y3_W6BEG[3] ;
 wire \Tile_X2Y3_W6BEG[4] ;
 wire \Tile_X2Y3_W6BEG[5] ;
 wire \Tile_X2Y3_W6BEG[6] ;
 wire \Tile_X2Y3_W6BEG[7] ;
 wire \Tile_X2Y3_W6BEG[8] ;
 wire \Tile_X2Y3_W6BEG[9] ;
 wire \Tile_X2Y3_WW4BEG[0] ;
 wire \Tile_X2Y3_WW4BEG[10] ;
 wire \Tile_X2Y3_WW4BEG[11] ;
 wire \Tile_X2Y3_WW4BEG[12] ;
 wire \Tile_X2Y3_WW4BEG[13] ;
 wire \Tile_X2Y3_WW4BEG[14] ;
 wire \Tile_X2Y3_WW4BEG[15] ;
 wire \Tile_X2Y3_WW4BEG[1] ;
 wire \Tile_X2Y3_WW4BEG[2] ;
 wire \Tile_X2Y3_WW4BEG[3] ;
 wire \Tile_X2Y3_WW4BEG[4] ;
 wire \Tile_X2Y3_WW4BEG[5] ;
 wire \Tile_X2Y3_WW4BEG[6] ;
 wire \Tile_X2Y3_WW4BEG[7] ;
 wire \Tile_X2Y3_WW4BEG[8] ;
 wire \Tile_X2Y3_WW4BEG[9] ;
 wire Tile_X2Y4_Co;
 wire \Tile_X2Y4_E1BEG[0] ;
 wire \Tile_X2Y4_E1BEG[1] ;
 wire \Tile_X2Y4_E1BEG[2] ;
 wire \Tile_X2Y4_E1BEG[3] ;
 wire \Tile_X2Y4_E2BEG[0] ;
 wire \Tile_X2Y4_E2BEG[1] ;
 wire \Tile_X2Y4_E2BEG[2] ;
 wire \Tile_X2Y4_E2BEG[3] ;
 wire \Tile_X2Y4_E2BEG[4] ;
 wire \Tile_X2Y4_E2BEG[5] ;
 wire \Tile_X2Y4_E2BEG[6] ;
 wire \Tile_X2Y4_E2BEG[7] ;
 wire \Tile_X2Y4_E2BEGb[0] ;
 wire \Tile_X2Y4_E2BEGb[1] ;
 wire \Tile_X2Y4_E2BEGb[2] ;
 wire \Tile_X2Y4_E2BEGb[3] ;
 wire \Tile_X2Y4_E2BEGb[4] ;
 wire \Tile_X2Y4_E2BEGb[5] ;
 wire \Tile_X2Y4_E2BEGb[6] ;
 wire \Tile_X2Y4_E2BEGb[7] ;
 wire \Tile_X2Y4_E6BEG[0] ;
 wire \Tile_X2Y4_E6BEG[10] ;
 wire \Tile_X2Y4_E6BEG[11] ;
 wire \Tile_X2Y4_E6BEG[1] ;
 wire \Tile_X2Y4_E6BEG[2] ;
 wire \Tile_X2Y4_E6BEG[3] ;
 wire \Tile_X2Y4_E6BEG[4] ;
 wire \Tile_X2Y4_E6BEG[5] ;
 wire \Tile_X2Y4_E6BEG[6] ;
 wire \Tile_X2Y4_E6BEG[7] ;
 wire \Tile_X2Y4_E6BEG[8] ;
 wire \Tile_X2Y4_E6BEG[9] ;
 wire \Tile_X2Y4_EE4BEG[0] ;
 wire \Tile_X2Y4_EE4BEG[10] ;
 wire \Tile_X2Y4_EE4BEG[11] ;
 wire \Tile_X2Y4_EE4BEG[12] ;
 wire \Tile_X2Y4_EE4BEG[13] ;
 wire \Tile_X2Y4_EE4BEG[14] ;
 wire \Tile_X2Y4_EE4BEG[15] ;
 wire \Tile_X2Y4_EE4BEG[1] ;
 wire \Tile_X2Y4_EE4BEG[2] ;
 wire \Tile_X2Y4_EE4BEG[3] ;
 wire \Tile_X2Y4_EE4BEG[4] ;
 wire \Tile_X2Y4_EE4BEG[5] ;
 wire \Tile_X2Y4_EE4BEG[6] ;
 wire \Tile_X2Y4_EE4BEG[7] ;
 wire \Tile_X2Y4_EE4BEG[8] ;
 wire \Tile_X2Y4_EE4BEG[9] ;
 wire \Tile_X2Y4_FrameData_O[0] ;
 wire \Tile_X2Y4_FrameData_O[10] ;
 wire \Tile_X2Y4_FrameData_O[11] ;
 wire \Tile_X2Y4_FrameData_O[12] ;
 wire \Tile_X2Y4_FrameData_O[13] ;
 wire \Tile_X2Y4_FrameData_O[14] ;
 wire \Tile_X2Y4_FrameData_O[15] ;
 wire \Tile_X2Y4_FrameData_O[16] ;
 wire \Tile_X2Y4_FrameData_O[17] ;
 wire \Tile_X2Y4_FrameData_O[18] ;
 wire \Tile_X2Y4_FrameData_O[19] ;
 wire \Tile_X2Y4_FrameData_O[1] ;
 wire \Tile_X2Y4_FrameData_O[20] ;
 wire \Tile_X2Y4_FrameData_O[21] ;
 wire \Tile_X2Y4_FrameData_O[22] ;
 wire \Tile_X2Y4_FrameData_O[23] ;
 wire \Tile_X2Y4_FrameData_O[24] ;
 wire \Tile_X2Y4_FrameData_O[25] ;
 wire \Tile_X2Y4_FrameData_O[26] ;
 wire \Tile_X2Y4_FrameData_O[27] ;
 wire \Tile_X2Y4_FrameData_O[28] ;
 wire \Tile_X2Y4_FrameData_O[29] ;
 wire \Tile_X2Y4_FrameData_O[2] ;
 wire \Tile_X2Y4_FrameData_O[30] ;
 wire \Tile_X2Y4_FrameData_O[31] ;
 wire \Tile_X2Y4_FrameData_O[3] ;
 wire \Tile_X2Y4_FrameData_O[4] ;
 wire \Tile_X2Y4_FrameData_O[5] ;
 wire \Tile_X2Y4_FrameData_O[6] ;
 wire \Tile_X2Y4_FrameData_O[7] ;
 wire \Tile_X2Y4_FrameData_O[8] ;
 wire \Tile_X2Y4_FrameData_O[9] ;
 wire \Tile_X2Y4_FrameStrobe_O[0] ;
 wire \Tile_X2Y4_FrameStrobe_O[10] ;
 wire \Tile_X2Y4_FrameStrobe_O[11] ;
 wire \Tile_X2Y4_FrameStrobe_O[12] ;
 wire \Tile_X2Y4_FrameStrobe_O[13] ;
 wire \Tile_X2Y4_FrameStrobe_O[14] ;
 wire \Tile_X2Y4_FrameStrobe_O[15] ;
 wire \Tile_X2Y4_FrameStrobe_O[16] ;
 wire \Tile_X2Y4_FrameStrobe_O[17] ;
 wire \Tile_X2Y4_FrameStrobe_O[18] ;
 wire \Tile_X2Y4_FrameStrobe_O[19] ;
 wire \Tile_X2Y4_FrameStrobe_O[1] ;
 wire \Tile_X2Y4_FrameStrobe_O[2] ;
 wire \Tile_X2Y4_FrameStrobe_O[3] ;
 wire \Tile_X2Y4_FrameStrobe_O[4] ;
 wire \Tile_X2Y4_FrameStrobe_O[5] ;
 wire \Tile_X2Y4_FrameStrobe_O[6] ;
 wire \Tile_X2Y4_FrameStrobe_O[7] ;
 wire \Tile_X2Y4_FrameStrobe_O[8] ;
 wire \Tile_X2Y4_FrameStrobe_O[9] ;
 wire \Tile_X2Y4_N1BEG[0] ;
 wire \Tile_X2Y4_N1BEG[1] ;
 wire \Tile_X2Y4_N1BEG[2] ;
 wire \Tile_X2Y4_N1BEG[3] ;
 wire \Tile_X2Y4_N2BEG[0] ;
 wire \Tile_X2Y4_N2BEG[1] ;
 wire \Tile_X2Y4_N2BEG[2] ;
 wire \Tile_X2Y4_N2BEG[3] ;
 wire \Tile_X2Y4_N2BEG[4] ;
 wire \Tile_X2Y4_N2BEG[5] ;
 wire \Tile_X2Y4_N2BEG[6] ;
 wire \Tile_X2Y4_N2BEG[7] ;
 wire \Tile_X2Y4_N2BEGb[0] ;
 wire \Tile_X2Y4_N2BEGb[1] ;
 wire \Tile_X2Y4_N2BEGb[2] ;
 wire \Tile_X2Y4_N2BEGb[3] ;
 wire \Tile_X2Y4_N2BEGb[4] ;
 wire \Tile_X2Y4_N2BEGb[5] ;
 wire \Tile_X2Y4_N2BEGb[6] ;
 wire \Tile_X2Y4_N2BEGb[7] ;
 wire \Tile_X2Y4_N4BEG[0] ;
 wire \Tile_X2Y4_N4BEG[10] ;
 wire \Tile_X2Y4_N4BEG[11] ;
 wire \Tile_X2Y4_N4BEG[12] ;
 wire \Tile_X2Y4_N4BEG[13] ;
 wire \Tile_X2Y4_N4BEG[14] ;
 wire \Tile_X2Y4_N4BEG[15] ;
 wire \Tile_X2Y4_N4BEG[1] ;
 wire \Tile_X2Y4_N4BEG[2] ;
 wire \Tile_X2Y4_N4BEG[3] ;
 wire \Tile_X2Y4_N4BEG[4] ;
 wire \Tile_X2Y4_N4BEG[5] ;
 wire \Tile_X2Y4_N4BEG[6] ;
 wire \Tile_X2Y4_N4BEG[7] ;
 wire \Tile_X2Y4_N4BEG[8] ;
 wire \Tile_X2Y4_N4BEG[9] ;
 wire \Tile_X2Y4_NN4BEG[0] ;
 wire \Tile_X2Y4_NN4BEG[10] ;
 wire \Tile_X2Y4_NN4BEG[11] ;
 wire \Tile_X2Y4_NN4BEG[12] ;
 wire \Tile_X2Y4_NN4BEG[13] ;
 wire \Tile_X2Y4_NN4BEG[14] ;
 wire \Tile_X2Y4_NN4BEG[15] ;
 wire \Tile_X2Y4_NN4BEG[1] ;
 wire \Tile_X2Y4_NN4BEG[2] ;
 wire \Tile_X2Y4_NN4BEG[3] ;
 wire \Tile_X2Y4_NN4BEG[4] ;
 wire \Tile_X2Y4_NN4BEG[5] ;
 wire \Tile_X2Y4_NN4BEG[6] ;
 wire \Tile_X2Y4_NN4BEG[7] ;
 wire \Tile_X2Y4_NN4BEG[8] ;
 wire \Tile_X2Y4_NN4BEG[9] ;
 wire \Tile_X2Y4_S1BEG[0] ;
 wire \Tile_X2Y4_S1BEG[1] ;
 wire \Tile_X2Y4_S1BEG[2] ;
 wire \Tile_X2Y4_S1BEG[3] ;
 wire \Tile_X2Y4_S2BEG[0] ;
 wire \Tile_X2Y4_S2BEG[1] ;
 wire \Tile_X2Y4_S2BEG[2] ;
 wire \Tile_X2Y4_S2BEG[3] ;
 wire \Tile_X2Y4_S2BEG[4] ;
 wire \Tile_X2Y4_S2BEG[5] ;
 wire \Tile_X2Y4_S2BEG[6] ;
 wire \Tile_X2Y4_S2BEG[7] ;
 wire \Tile_X2Y4_S2BEGb[0] ;
 wire \Tile_X2Y4_S2BEGb[1] ;
 wire \Tile_X2Y4_S2BEGb[2] ;
 wire \Tile_X2Y4_S2BEGb[3] ;
 wire \Tile_X2Y4_S2BEGb[4] ;
 wire \Tile_X2Y4_S2BEGb[5] ;
 wire \Tile_X2Y4_S2BEGb[6] ;
 wire \Tile_X2Y4_S2BEGb[7] ;
 wire \Tile_X2Y4_S4BEG[0] ;
 wire \Tile_X2Y4_S4BEG[10] ;
 wire \Tile_X2Y4_S4BEG[11] ;
 wire \Tile_X2Y4_S4BEG[12] ;
 wire \Tile_X2Y4_S4BEG[13] ;
 wire \Tile_X2Y4_S4BEG[14] ;
 wire \Tile_X2Y4_S4BEG[15] ;
 wire \Tile_X2Y4_S4BEG[1] ;
 wire \Tile_X2Y4_S4BEG[2] ;
 wire \Tile_X2Y4_S4BEG[3] ;
 wire \Tile_X2Y4_S4BEG[4] ;
 wire \Tile_X2Y4_S4BEG[5] ;
 wire \Tile_X2Y4_S4BEG[6] ;
 wire \Tile_X2Y4_S4BEG[7] ;
 wire \Tile_X2Y4_S4BEG[8] ;
 wire \Tile_X2Y4_S4BEG[9] ;
 wire \Tile_X2Y4_SS4BEG[0] ;
 wire \Tile_X2Y4_SS4BEG[10] ;
 wire \Tile_X2Y4_SS4BEG[11] ;
 wire \Tile_X2Y4_SS4BEG[12] ;
 wire \Tile_X2Y4_SS4BEG[13] ;
 wire \Tile_X2Y4_SS4BEG[14] ;
 wire \Tile_X2Y4_SS4BEG[15] ;
 wire \Tile_X2Y4_SS4BEG[1] ;
 wire \Tile_X2Y4_SS4BEG[2] ;
 wire \Tile_X2Y4_SS4BEG[3] ;
 wire \Tile_X2Y4_SS4BEG[4] ;
 wire \Tile_X2Y4_SS4BEG[5] ;
 wire \Tile_X2Y4_SS4BEG[6] ;
 wire \Tile_X2Y4_SS4BEG[7] ;
 wire \Tile_X2Y4_SS4BEG[8] ;
 wire \Tile_X2Y4_SS4BEG[9] ;
 wire Tile_X2Y4_UserCLKo;
 wire \Tile_X2Y4_W1BEG[0] ;
 wire \Tile_X2Y4_W1BEG[1] ;
 wire \Tile_X2Y4_W1BEG[2] ;
 wire \Tile_X2Y4_W1BEG[3] ;
 wire \Tile_X2Y4_W2BEG[0] ;
 wire \Tile_X2Y4_W2BEG[1] ;
 wire \Tile_X2Y4_W2BEG[2] ;
 wire \Tile_X2Y4_W2BEG[3] ;
 wire \Tile_X2Y4_W2BEG[4] ;
 wire \Tile_X2Y4_W2BEG[5] ;
 wire \Tile_X2Y4_W2BEG[6] ;
 wire \Tile_X2Y4_W2BEG[7] ;
 wire \Tile_X2Y4_W2BEGb[0] ;
 wire \Tile_X2Y4_W2BEGb[1] ;
 wire \Tile_X2Y4_W2BEGb[2] ;
 wire \Tile_X2Y4_W2BEGb[3] ;
 wire \Tile_X2Y4_W2BEGb[4] ;
 wire \Tile_X2Y4_W2BEGb[5] ;
 wire \Tile_X2Y4_W2BEGb[6] ;
 wire \Tile_X2Y4_W2BEGb[7] ;
 wire \Tile_X2Y4_W6BEG[0] ;
 wire \Tile_X2Y4_W6BEG[10] ;
 wire \Tile_X2Y4_W6BEG[11] ;
 wire \Tile_X2Y4_W6BEG[1] ;
 wire \Tile_X2Y4_W6BEG[2] ;
 wire \Tile_X2Y4_W6BEG[3] ;
 wire \Tile_X2Y4_W6BEG[4] ;
 wire \Tile_X2Y4_W6BEG[5] ;
 wire \Tile_X2Y4_W6BEG[6] ;
 wire \Tile_X2Y4_W6BEG[7] ;
 wire \Tile_X2Y4_W6BEG[8] ;
 wire \Tile_X2Y4_W6BEG[9] ;
 wire \Tile_X2Y4_WW4BEG[0] ;
 wire \Tile_X2Y4_WW4BEG[10] ;
 wire \Tile_X2Y4_WW4BEG[11] ;
 wire \Tile_X2Y4_WW4BEG[12] ;
 wire \Tile_X2Y4_WW4BEG[13] ;
 wire \Tile_X2Y4_WW4BEG[14] ;
 wire \Tile_X2Y4_WW4BEG[15] ;
 wire \Tile_X2Y4_WW4BEG[1] ;
 wire \Tile_X2Y4_WW4BEG[2] ;
 wire \Tile_X2Y4_WW4BEG[3] ;
 wire \Tile_X2Y4_WW4BEG[4] ;
 wire \Tile_X2Y4_WW4BEG[5] ;
 wire \Tile_X2Y4_WW4BEG[6] ;
 wire \Tile_X2Y4_WW4BEG[7] ;
 wire \Tile_X2Y4_WW4BEG[8] ;
 wire \Tile_X2Y4_WW4BEG[9] ;
 wire Tile_X2Y5_Co;
 wire \Tile_X2Y5_E1BEG[0] ;
 wire \Tile_X2Y5_E1BEG[1] ;
 wire \Tile_X2Y5_E1BEG[2] ;
 wire \Tile_X2Y5_E1BEG[3] ;
 wire \Tile_X2Y5_E2BEG[0] ;
 wire \Tile_X2Y5_E2BEG[1] ;
 wire \Tile_X2Y5_E2BEG[2] ;
 wire \Tile_X2Y5_E2BEG[3] ;
 wire \Tile_X2Y5_E2BEG[4] ;
 wire \Tile_X2Y5_E2BEG[5] ;
 wire \Tile_X2Y5_E2BEG[6] ;
 wire \Tile_X2Y5_E2BEG[7] ;
 wire \Tile_X2Y5_E2BEGb[0] ;
 wire \Tile_X2Y5_E2BEGb[1] ;
 wire \Tile_X2Y5_E2BEGb[2] ;
 wire \Tile_X2Y5_E2BEGb[3] ;
 wire \Tile_X2Y5_E2BEGb[4] ;
 wire \Tile_X2Y5_E2BEGb[5] ;
 wire \Tile_X2Y5_E2BEGb[6] ;
 wire \Tile_X2Y5_E2BEGb[7] ;
 wire \Tile_X2Y5_E6BEG[0] ;
 wire \Tile_X2Y5_E6BEG[10] ;
 wire \Tile_X2Y5_E6BEG[11] ;
 wire \Tile_X2Y5_E6BEG[1] ;
 wire \Tile_X2Y5_E6BEG[2] ;
 wire \Tile_X2Y5_E6BEG[3] ;
 wire \Tile_X2Y5_E6BEG[4] ;
 wire \Tile_X2Y5_E6BEG[5] ;
 wire \Tile_X2Y5_E6BEG[6] ;
 wire \Tile_X2Y5_E6BEG[7] ;
 wire \Tile_X2Y5_E6BEG[8] ;
 wire \Tile_X2Y5_E6BEG[9] ;
 wire \Tile_X2Y5_EE4BEG[0] ;
 wire \Tile_X2Y5_EE4BEG[10] ;
 wire \Tile_X2Y5_EE4BEG[11] ;
 wire \Tile_X2Y5_EE4BEG[12] ;
 wire \Tile_X2Y5_EE4BEG[13] ;
 wire \Tile_X2Y5_EE4BEG[14] ;
 wire \Tile_X2Y5_EE4BEG[15] ;
 wire \Tile_X2Y5_EE4BEG[1] ;
 wire \Tile_X2Y5_EE4BEG[2] ;
 wire \Tile_X2Y5_EE4BEG[3] ;
 wire \Tile_X2Y5_EE4BEG[4] ;
 wire \Tile_X2Y5_EE4BEG[5] ;
 wire \Tile_X2Y5_EE4BEG[6] ;
 wire \Tile_X2Y5_EE4BEG[7] ;
 wire \Tile_X2Y5_EE4BEG[8] ;
 wire \Tile_X2Y5_EE4BEG[9] ;
 wire \Tile_X2Y5_FrameData_O[0] ;
 wire \Tile_X2Y5_FrameData_O[10] ;
 wire \Tile_X2Y5_FrameData_O[11] ;
 wire \Tile_X2Y5_FrameData_O[12] ;
 wire \Tile_X2Y5_FrameData_O[13] ;
 wire \Tile_X2Y5_FrameData_O[14] ;
 wire \Tile_X2Y5_FrameData_O[15] ;
 wire \Tile_X2Y5_FrameData_O[16] ;
 wire \Tile_X2Y5_FrameData_O[17] ;
 wire \Tile_X2Y5_FrameData_O[18] ;
 wire \Tile_X2Y5_FrameData_O[19] ;
 wire \Tile_X2Y5_FrameData_O[1] ;
 wire \Tile_X2Y5_FrameData_O[20] ;
 wire \Tile_X2Y5_FrameData_O[21] ;
 wire \Tile_X2Y5_FrameData_O[22] ;
 wire \Tile_X2Y5_FrameData_O[23] ;
 wire \Tile_X2Y5_FrameData_O[24] ;
 wire \Tile_X2Y5_FrameData_O[25] ;
 wire \Tile_X2Y5_FrameData_O[26] ;
 wire \Tile_X2Y5_FrameData_O[27] ;
 wire \Tile_X2Y5_FrameData_O[28] ;
 wire \Tile_X2Y5_FrameData_O[29] ;
 wire \Tile_X2Y5_FrameData_O[2] ;
 wire \Tile_X2Y5_FrameData_O[30] ;
 wire \Tile_X2Y5_FrameData_O[31] ;
 wire \Tile_X2Y5_FrameData_O[3] ;
 wire \Tile_X2Y5_FrameData_O[4] ;
 wire \Tile_X2Y5_FrameData_O[5] ;
 wire \Tile_X2Y5_FrameData_O[6] ;
 wire \Tile_X2Y5_FrameData_O[7] ;
 wire \Tile_X2Y5_FrameData_O[8] ;
 wire \Tile_X2Y5_FrameData_O[9] ;
 wire \Tile_X2Y5_FrameStrobe_O[0] ;
 wire \Tile_X2Y5_FrameStrobe_O[10] ;
 wire \Tile_X2Y5_FrameStrobe_O[11] ;
 wire \Tile_X2Y5_FrameStrobe_O[12] ;
 wire \Tile_X2Y5_FrameStrobe_O[13] ;
 wire \Tile_X2Y5_FrameStrobe_O[14] ;
 wire \Tile_X2Y5_FrameStrobe_O[15] ;
 wire \Tile_X2Y5_FrameStrobe_O[16] ;
 wire \Tile_X2Y5_FrameStrobe_O[17] ;
 wire \Tile_X2Y5_FrameStrobe_O[18] ;
 wire \Tile_X2Y5_FrameStrobe_O[19] ;
 wire \Tile_X2Y5_FrameStrobe_O[1] ;
 wire \Tile_X2Y5_FrameStrobe_O[2] ;
 wire \Tile_X2Y5_FrameStrobe_O[3] ;
 wire \Tile_X2Y5_FrameStrobe_O[4] ;
 wire \Tile_X2Y5_FrameStrobe_O[5] ;
 wire \Tile_X2Y5_FrameStrobe_O[6] ;
 wire \Tile_X2Y5_FrameStrobe_O[7] ;
 wire \Tile_X2Y5_FrameStrobe_O[8] ;
 wire \Tile_X2Y5_FrameStrobe_O[9] ;
 wire \Tile_X2Y5_N1BEG[0] ;
 wire \Tile_X2Y5_N1BEG[1] ;
 wire \Tile_X2Y5_N1BEG[2] ;
 wire \Tile_X2Y5_N1BEG[3] ;
 wire \Tile_X2Y5_N2BEG[0] ;
 wire \Tile_X2Y5_N2BEG[1] ;
 wire \Tile_X2Y5_N2BEG[2] ;
 wire \Tile_X2Y5_N2BEG[3] ;
 wire \Tile_X2Y5_N2BEG[4] ;
 wire \Tile_X2Y5_N2BEG[5] ;
 wire \Tile_X2Y5_N2BEG[6] ;
 wire \Tile_X2Y5_N2BEG[7] ;
 wire \Tile_X2Y5_N2BEGb[0] ;
 wire \Tile_X2Y5_N2BEGb[1] ;
 wire \Tile_X2Y5_N2BEGb[2] ;
 wire \Tile_X2Y5_N2BEGb[3] ;
 wire \Tile_X2Y5_N2BEGb[4] ;
 wire \Tile_X2Y5_N2BEGb[5] ;
 wire \Tile_X2Y5_N2BEGb[6] ;
 wire \Tile_X2Y5_N2BEGb[7] ;
 wire \Tile_X2Y5_N4BEG[0] ;
 wire \Tile_X2Y5_N4BEG[10] ;
 wire \Tile_X2Y5_N4BEG[11] ;
 wire \Tile_X2Y5_N4BEG[12] ;
 wire \Tile_X2Y5_N4BEG[13] ;
 wire \Tile_X2Y5_N4BEG[14] ;
 wire \Tile_X2Y5_N4BEG[15] ;
 wire \Tile_X2Y5_N4BEG[1] ;
 wire \Tile_X2Y5_N4BEG[2] ;
 wire \Tile_X2Y5_N4BEG[3] ;
 wire \Tile_X2Y5_N4BEG[4] ;
 wire \Tile_X2Y5_N4BEG[5] ;
 wire \Tile_X2Y5_N4BEG[6] ;
 wire \Tile_X2Y5_N4BEG[7] ;
 wire \Tile_X2Y5_N4BEG[8] ;
 wire \Tile_X2Y5_N4BEG[9] ;
 wire \Tile_X2Y5_NN4BEG[0] ;
 wire \Tile_X2Y5_NN4BEG[10] ;
 wire \Tile_X2Y5_NN4BEG[11] ;
 wire \Tile_X2Y5_NN4BEG[12] ;
 wire \Tile_X2Y5_NN4BEG[13] ;
 wire \Tile_X2Y5_NN4BEG[14] ;
 wire \Tile_X2Y5_NN4BEG[15] ;
 wire \Tile_X2Y5_NN4BEG[1] ;
 wire \Tile_X2Y5_NN4BEG[2] ;
 wire \Tile_X2Y5_NN4BEG[3] ;
 wire \Tile_X2Y5_NN4BEG[4] ;
 wire \Tile_X2Y5_NN4BEG[5] ;
 wire \Tile_X2Y5_NN4BEG[6] ;
 wire \Tile_X2Y5_NN4BEG[7] ;
 wire \Tile_X2Y5_NN4BEG[8] ;
 wire \Tile_X2Y5_NN4BEG[9] ;
 wire \Tile_X2Y5_S1BEG[0] ;
 wire \Tile_X2Y5_S1BEG[1] ;
 wire \Tile_X2Y5_S1BEG[2] ;
 wire \Tile_X2Y5_S1BEG[3] ;
 wire \Tile_X2Y5_S2BEG[0] ;
 wire \Tile_X2Y5_S2BEG[1] ;
 wire \Tile_X2Y5_S2BEG[2] ;
 wire \Tile_X2Y5_S2BEG[3] ;
 wire \Tile_X2Y5_S2BEG[4] ;
 wire \Tile_X2Y5_S2BEG[5] ;
 wire \Tile_X2Y5_S2BEG[6] ;
 wire \Tile_X2Y5_S2BEG[7] ;
 wire \Tile_X2Y5_S2BEGb[0] ;
 wire \Tile_X2Y5_S2BEGb[1] ;
 wire \Tile_X2Y5_S2BEGb[2] ;
 wire \Tile_X2Y5_S2BEGb[3] ;
 wire \Tile_X2Y5_S2BEGb[4] ;
 wire \Tile_X2Y5_S2BEGb[5] ;
 wire \Tile_X2Y5_S2BEGb[6] ;
 wire \Tile_X2Y5_S2BEGb[7] ;
 wire \Tile_X2Y5_S4BEG[0] ;
 wire \Tile_X2Y5_S4BEG[10] ;
 wire \Tile_X2Y5_S4BEG[11] ;
 wire \Tile_X2Y5_S4BEG[12] ;
 wire \Tile_X2Y5_S4BEG[13] ;
 wire \Tile_X2Y5_S4BEG[14] ;
 wire \Tile_X2Y5_S4BEG[15] ;
 wire \Tile_X2Y5_S4BEG[1] ;
 wire \Tile_X2Y5_S4BEG[2] ;
 wire \Tile_X2Y5_S4BEG[3] ;
 wire \Tile_X2Y5_S4BEG[4] ;
 wire \Tile_X2Y5_S4BEG[5] ;
 wire \Tile_X2Y5_S4BEG[6] ;
 wire \Tile_X2Y5_S4BEG[7] ;
 wire \Tile_X2Y5_S4BEG[8] ;
 wire \Tile_X2Y5_S4BEG[9] ;
 wire \Tile_X2Y5_SS4BEG[0] ;
 wire \Tile_X2Y5_SS4BEG[10] ;
 wire \Tile_X2Y5_SS4BEG[11] ;
 wire \Tile_X2Y5_SS4BEG[12] ;
 wire \Tile_X2Y5_SS4BEG[13] ;
 wire \Tile_X2Y5_SS4BEG[14] ;
 wire \Tile_X2Y5_SS4BEG[15] ;
 wire \Tile_X2Y5_SS4BEG[1] ;
 wire \Tile_X2Y5_SS4BEG[2] ;
 wire \Tile_X2Y5_SS4BEG[3] ;
 wire \Tile_X2Y5_SS4BEG[4] ;
 wire \Tile_X2Y5_SS4BEG[5] ;
 wire \Tile_X2Y5_SS4BEG[6] ;
 wire \Tile_X2Y5_SS4BEG[7] ;
 wire \Tile_X2Y5_SS4BEG[8] ;
 wire \Tile_X2Y5_SS4BEG[9] ;
 wire Tile_X2Y5_UserCLKo;
 wire \Tile_X2Y5_W1BEG[0] ;
 wire \Tile_X2Y5_W1BEG[1] ;
 wire \Tile_X2Y5_W1BEG[2] ;
 wire \Tile_X2Y5_W1BEG[3] ;
 wire \Tile_X2Y5_W2BEG[0] ;
 wire \Tile_X2Y5_W2BEG[1] ;
 wire \Tile_X2Y5_W2BEG[2] ;
 wire \Tile_X2Y5_W2BEG[3] ;
 wire \Tile_X2Y5_W2BEG[4] ;
 wire \Tile_X2Y5_W2BEG[5] ;
 wire \Tile_X2Y5_W2BEG[6] ;
 wire \Tile_X2Y5_W2BEG[7] ;
 wire \Tile_X2Y5_W2BEGb[0] ;
 wire \Tile_X2Y5_W2BEGb[1] ;
 wire \Tile_X2Y5_W2BEGb[2] ;
 wire \Tile_X2Y5_W2BEGb[3] ;
 wire \Tile_X2Y5_W2BEGb[4] ;
 wire \Tile_X2Y5_W2BEGb[5] ;
 wire \Tile_X2Y5_W2BEGb[6] ;
 wire \Tile_X2Y5_W2BEGb[7] ;
 wire \Tile_X2Y5_W6BEG[0] ;
 wire \Tile_X2Y5_W6BEG[10] ;
 wire \Tile_X2Y5_W6BEG[11] ;
 wire \Tile_X2Y5_W6BEG[1] ;
 wire \Tile_X2Y5_W6BEG[2] ;
 wire \Tile_X2Y5_W6BEG[3] ;
 wire \Tile_X2Y5_W6BEG[4] ;
 wire \Tile_X2Y5_W6BEG[5] ;
 wire \Tile_X2Y5_W6BEG[6] ;
 wire \Tile_X2Y5_W6BEG[7] ;
 wire \Tile_X2Y5_W6BEG[8] ;
 wire \Tile_X2Y5_W6BEG[9] ;
 wire \Tile_X2Y5_WW4BEG[0] ;
 wire \Tile_X2Y5_WW4BEG[10] ;
 wire \Tile_X2Y5_WW4BEG[11] ;
 wire \Tile_X2Y5_WW4BEG[12] ;
 wire \Tile_X2Y5_WW4BEG[13] ;
 wire \Tile_X2Y5_WW4BEG[14] ;
 wire \Tile_X2Y5_WW4BEG[15] ;
 wire \Tile_X2Y5_WW4BEG[1] ;
 wire \Tile_X2Y5_WW4BEG[2] ;
 wire \Tile_X2Y5_WW4BEG[3] ;
 wire \Tile_X2Y5_WW4BEG[4] ;
 wire \Tile_X2Y5_WW4BEG[5] ;
 wire \Tile_X2Y5_WW4BEG[6] ;
 wire \Tile_X2Y5_WW4BEG[7] ;
 wire \Tile_X2Y5_WW4BEG[8] ;
 wire \Tile_X2Y5_WW4BEG[9] ;
 wire Tile_X2Y6_Co;
 wire \Tile_X2Y6_E1BEG[0] ;
 wire \Tile_X2Y6_E1BEG[1] ;
 wire \Tile_X2Y6_E1BEG[2] ;
 wire \Tile_X2Y6_E1BEG[3] ;
 wire \Tile_X2Y6_E2BEG[0] ;
 wire \Tile_X2Y6_E2BEG[1] ;
 wire \Tile_X2Y6_E2BEG[2] ;
 wire \Tile_X2Y6_E2BEG[3] ;
 wire \Tile_X2Y6_E2BEG[4] ;
 wire \Tile_X2Y6_E2BEG[5] ;
 wire \Tile_X2Y6_E2BEG[6] ;
 wire \Tile_X2Y6_E2BEG[7] ;
 wire \Tile_X2Y6_E2BEGb[0] ;
 wire \Tile_X2Y6_E2BEGb[1] ;
 wire \Tile_X2Y6_E2BEGb[2] ;
 wire \Tile_X2Y6_E2BEGb[3] ;
 wire \Tile_X2Y6_E2BEGb[4] ;
 wire \Tile_X2Y6_E2BEGb[5] ;
 wire \Tile_X2Y6_E2BEGb[6] ;
 wire \Tile_X2Y6_E2BEGb[7] ;
 wire \Tile_X2Y6_E6BEG[0] ;
 wire \Tile_X2Y6_E6BEG[10] ;
 wire \Tile_X2Y6_E6BEG[11] ;
 wire \Tile_X2Y6_E6BEG[1] ;
 wire \Tile_X2Y6_E6BEG[2] ;
 wire \Tile_X2Y6_E6BEG[3] ;
 wire \Tile_X2Y6_E6BEG[4] ;
 wire \Tile_X2Y6_E6BEG[5] ;
 wire \Tile_X2Y6_E6BEG[6] ;
 wire \Tile_X2Y6_E6BEG[7] ;
 wire \Tile_X2Y6_E6BEG[8] ;
 wire \Tile_X2Y6_E6BEG[9] ;
 wire \Tile_X2Y6_EE4BEG[0] ;
 wire \Tile_X2Y6_EE4BEG[10] ;
 wire \Tile_X2Y6_EE4BEG[11] ;
 wire \Tile_X2Y6_EE4BEG[12] ;
 wire \Tile_X2Y6_EE4BEG[13] ;
 wire \Tile_X2Y6_EE4BEG[14] ;
 wire \Tile_X2Y6_EE4BEG[15] ;
 wire \Tile_X2Y6_EE4BEG[1] ;
 wire \Tile_X2Y6_EE4BEG[2] ;
 wire \Tile_X2Y6_EE4BEG[3] ;
 wire \Tile_X2Y6_EE4BEG[4] ;
 wire \Tile_X2Y6_EE4BEG[5] ;
 wire \Tile_X2Y6_EE4BEG[6] ;
 wire \Tile_X2Y6_EE4BEG[7] ;
 wire \Tile_X2Y6_EE4BEG[8] ;
 wire \Tile_X2Y6_EE4BEG[9] ;
 wire \Tile_X2Y6_FrameData_O[0] ;
 wire \Tile_X2Y6_FrameData_O[10] ;
 wire \Tile_X2Y6_FrameData_O[11] ;
 wire \Tile_X2Y6_FrameData_O[12] ;
 wire \Tile_X2Y6_FrameData_O[13] ;
 wire \Tile_X2Y6_FrameData_O[14] ;
 wire \Tile_X2Y6_FrameData_O[15] ;
 wire \Tile_X2Y6_FrameData_O[16] ;
 wire \Tile_X2Y6_FrameData_O[17] ;
 wire \Tile_X2Y6_FrameData_O[18] ;
 wire \Tile_X2Y6_FrameData_O[19] ;
 wire \Tile_X2Y6_FrameData_O[1] ;
 wire \Tile_X2Y6_FrameData_O[20] ;
 wire \Tile_X2Y6_FrameData_O[21] ;
 wire \Tile_X2Y6_FrameData_O[22] ;
 wire \Tile_X2Y6_FrameData_O[23] ;
 wire \Tile_X2Y6_FrameData_O[24] ;
 wire \Tile_X2Y6_FrameData_O[25] ;
 wire \Tile_X2Y6_FrameData_O[26] ;
 wire \Tile_X2Y6_FrameData_O[27] ;
 wire \Tile_X2Y6_FrameData_O[28] ;
 wire \Tile_X2Y6_FrameData_O[29] ;
 wire \Tile_X2Y6_FrameData_O[2] ;
 wire \Tile_X2Y6_FrameData_O[30] ;
 wire \Tile_X2Y6_FrameData_O[31] ;
 wire \Tile_X2Y6_FrameData_O[3] ;
 wire \Tile_X2Y6_FrameData_O[4] ;
 wire \Tile_X2Y6_FrameData_O[5] ;
 wire \Tile_X2Y6_FrameData_O[6] ;
 wire \Tile_X2Y6_FrameData_O[7] ;
 wire \Tile_X2Y6_FrameData_O[8] ;
 wire \Tile_X2Y6_FrameData_O[9] ;
 wire \Tile_X2Y6_FrameStrobe_O[0] ;
 wire \Tile_X2Y6_FrameStrobe_O[10] ;
 wire \Tile_X2Y6_FrameStrobe_O[11] ;
 wire \Tile_X2Y6_FrameStrobe_O[12] ;
 wire \Tile_X2Y6_FrameStrobe_O[13] ;
 wire \Tile_X2Y6_FrameStrobe_O[14] ;
 wire \Tile_X2Y6_FrameStrobe_O[15] ;
 wire \Tile_X2Y6_FrameStrobe_O[16] ;
 wire \Tile_X2Y6_FrameStrobe_O[17] ;
 wire \Tile_X2Y6_FrameStrobe_O[18] ;
 wire \Tile_X2Y6_FrameStrobe_O[19] ;
 wire \Tile_X2Y6_FrameStrobe_O[1] ;
 wire \Tile_X2Y6_FrameStrobe_O[2] ;
 wire \Tile_X2Y6_FrameStrobe_O[3] ;
 wire \Tile_X2Y6_FrameStrobe_O[4] ;
 wire \Tile_X2Y6_FrameStrobe_O[5] ;
 wire \Tile_X2Y6_FrameStrobe_O[6] ;
 wire \Tile_X2Y6_FrameStrobe_O[7] ;
 wire \Tile_X2Y6_FrameStrobe_O[8] ;
 wire \Tile_X2Y6_FrameStrobe_O[9] ;
 wire \Tile_X2Y6_N1BEG[0] ;
 wire \Tile_X2Y6_N1BEG[1] ;
 wire \Tile_X2Y6_N1BEG[2] ;
 wire \Tile_X2Y6_N1BEG[3] ;
 wire \Tile_X2Y6_N2BEG[0] ;
 wire \Tile_X2Y6_N2BEG[1] ;
 wire \Tile_X2Y6_N2BEG[2] ;
 wire \Tile_X2Y6_N2BEG[3] ;
 wire \Tile_X2Y6_N2BEG[4] ;
 wire \Tile_X2Y6_N2BEG[5] ;
 wire \Tile_X2Y6_N2BEG[6] ;
 wire \Tile_X2Y6_N2BEG[7] ;
 wire \Tile_X2Y6_N2BEGb[0] ;
 wire \Tile_X2Y6_N2BEGb[1] ;
 wire \Tile_X2Y6_N2BEGb[2] ;
 wire \Tile_X2Y6_N2BEGb[3] ;
 wire \Tile_X2Y6_N2BEGb[4] ;
 wire \Tile_X2Y6_N2BEGb[5] ;
 wire \Tile_X2Y6_N2BEGb[6] ;
 wire \Tile_X2Y6_N2BEGb[7] ;
 wire \Tile_X2Y6_N4BEG[0] ;
 wire \Tile_X2Y6_N4BEG[10] ;
 wire \Tile_X2Y6_N4BEG[11] ;
 wire \Tile_X2Y6_N4BEG[12] ;
 wire \Tile_X2Y6_N4BEG[13] ;
 wire \Tile_X2Y6_N4BEG[14] ;
 wire \Tile_X2Y6_N4BEG[15] ;
 wire \Tile_X2Y6_N4BEG[1] ;
 wire \Tile_X2Y6_N4BEG[2] ;
 wire \Tile_X2Y6_N4BEG[3] ;
 wire \Tile_X2Y6_N4BEG[4] ;
 wire \Tile_X2Y6_N4BEG[5] ;
 wire \Tile_X2Y6_N4BEG[6] ;
 wire \Tile_X2Y6_N4BEG[7] ;
 wire \Tile_X2Y6_N4BEG[8] ;
 wire \Tile_X2Y6_N4BEG[9] ;
 wire \Tile_X2Y6_NN4BEG[0] ;
 wire \Tile_X2Y6_NN4BEG[10] ;
 wire \Tile_X2Y6_NN4BEG[11] ;
 wire \Tile_X2Y6_NN4BEG[12] ;
 wire \Tile_X2Y6_NN4BEG[13] ;
 wire \Tile_X2Y6_NN4BEG[14] ;
 wire \Tile_X2Y6_NN4BEG[15] ;
 wire \Tile_X2Y6_NN4BEG[1] ;
 wire \Tile_X2Y6_NN4BEG[2] ;
 wire \Tile_X2Y6_NN4BEG[3] ;
 wire \Tile_X2Y6_NN4BEG[4] ;
 wire \Tile_X2Y6_NN4BEG[5] ;
 wire \Tile_X2Y6_NN4BEG[6] ;
 wire \Tile_X2Y6_NN4BEG[7] ;
 wire \Tile_X2Y6_NN4BEG[8] ;
 wire \Tile_X2Y6_NN4BEG[9] ;
 wire \Tile_X2Y6_S1BEG[0] ;
 wire \Tile_X2Y6_S1BEG[1] ;
 wire \Tile_X2Y6_S1BEG[2] ;
 wire \Tile_X2Y6_S1BEG[3] ;
 wire \Tile_X2Y6_S2BEG[0] ;
 wire \Tile_X2Y6_S2BEG[1] ;
 wire \Tile_X2Y6_S2BEG[2] ;
 wire \Tile_X2Y6_S2BEG[3] ;
 wire \Tile_X2Y6_S2BEG[4] ;
 wire \Tile_X2Y6_S2BEG[5] ;
 wire \Tile_X2Y6_S2BEG[6] ;
 wire \Tile_X2Y6_S2BEG[7] ;
 wire \Tile_X2Y6_S2BEGb[0] ;
 wire \Tile_X2Y6_S2BEGb[1] ;
 wire \Tile_X2Y6_S2BEGb[2] ;
 wire \Tile_X2Y6_S2BEGb[3] ;
 wire \Tile_X2Y6_S2BEGb[4] ;
 wire \Tile_X2Y6_S2BEGb[5] ;
 wire \Tile_X2Y6_S2BEGb[6] ;
 wire \Tile_X2Y6_S2BEGb[7] ;
 wire \Tile_X2Y6_S4BEG[0] ;
 wire \Tile_X2Y6_S4BEG[10] ;
 wire \Tile_X2Y6_S4BEG[11] ;
 wire \Tile_X2Y6_S4BEG[12] ;
 wire \Tile_X2Y6_S4BEG[13] ;
 wire \Tile_X2Y6_S4BEG[14] ;
 wire \Tile_X2Y6_S4BEG[15] ;
 wire \Tile_X2Y6_S4BEG[1] ;
 wire \Tile_X2Y6_S4BEG[2] ;
 wire \Tile_X2Y6_S4BEG[3] ;
 wire \Tile_X2Y6_S4BEG[4] ;
 wire \Tile_X2Y6_S4BEG[5] ;
 wire \Tile_X2Y6_S4BEG[6] ;
 wire \Tile_X2Y6_S4BEG[7] ;
 wire \Tile_X2Y6_S4BEG[8] ;
 wire \Tile_X2Y6_S4BEG[9] ;
 wire \Tile_X2Y6_SS4BEG[0] ;
 wire \Tile_X2Y6_SS4BEG[10] ;
 wire \Tile_X2Y6_SS4BEG[11] ;
 wire \Tile_X2Y6_SS4BEG[12] ;
 wire \Tile_X2Y6_SS4BEG[13] ;
 wire \Tile_X2Y6_SS4BEG[14] ;
 wire \Tile_X2Y6_SS4BEG[15] ;
 wire \Tile_X2Y6_SS4BEG[1] ;
 wire \Tile_X2Y6_SS4BEG[2] ;
 wire \Tile_X2Y6_SS4BEG[3] ;
 wire \Tile_X2Y6_SS4BEG[4] ;
 wire \Tile_X2Y6_SS4BEG[5] ;
 wire \Tile_X2Y6_SS4BEG[6] ;
 wire \Tile_X2Y6_SS4BEG[7] ;
 wire \Tile_X2Y6_SS4BEG[8] ;
 wire \Tile_X2Y6_SS4BEG[9] ;
 wire Tile_X2Y6_UserCLKo;
 wire \Tile_X2Y6_W1BEG[0] ;
 wire \Tile_X2Y6_W1BEG[1] ;
 wire \Tile_X2Y6_W1BEG[2] ;
 wire \Tile_X2Y6_W1BEG[3] ;
 wire \Tile_X2Y6_W2BEG[0] ;
 wire \Tile_X2Y6_W2BEG[1] ;
 wire \Tile_X2Y6_W2BEG[2] ;
 wire \Tile_X2Y6_W2BEG[3] ;
 wire \Tile_X2Y6_W2BEG[4] ;
 wire \Tile_X2Y6_W2BEG[5] ;
 wire \Tile_X2Y6_W2BEG[6] ;
 wire \Tile_X2Y6_W2BEG[7] ;
 wire \Tile_X2Y6_W2BEGb[0] ;
 wire \Tile_X2Y6_W2BEGb[1] ;
 wire \Tile_X2Y6_W2BEGb[2] ;
 wire \Tile_X2Y6_W2BEGb[3] ;
 wire \Tile_X2Y6_W2BEGb[4] ;
 wire \Tile_X2Y6_W2BEGb[5] ;
 wire \Tile_X2Y6_W2BEGb[6] ;
 wire \Tile_X2Y6_W2BEGb[7] ;
 wire \Tile_X2Y6_W6BEG[0] ;
 wire \Tile_X2Y6_W6BEG[10] ;
 wire \Tile_X2Y6_W6BEG[11] ;
 wire \Tile_X2Y6_W6BEG[1] ;
 wire \Tile_X2Y6_W6BEG[2] ;
 wire \Tile_X2Y6_W6BEG[3] ;
 wire \Tile_X2Y6_W6BEG[4] ;
 wire \Tile_X2Y6_W6BEG[5] ;
 wire \Tile_X2Y6_W6BEG[6] ;
 wire \Tile_X2Y6_W6BEG[7] ;
 wire \Tile_X2Y6_W6BEG[8] ;
 wire \Tile_X2Y6_W6BEG[9] ;
 wire \Tile_X2Y6_WW4BEG[0] ;
 wire \Tile_X2Y6_WW4BEG[10] ;
 wire \Tile_X2Y6_WW4BEG[11] ;
 wire \Tile_X2Y6_WW4BEG[12] ;
 wire \Tile_X2Y6_WW4BEG[13] ;
 wire \Tile_X2Y6_WW4BEG[14] ;
 wire \Tile_X2Y6_WW4BEG[15] ;
 wire \Tile_X2Y6_WW4BEG[1] ;
 wire \Tile_X2Y6_WW4BEG[2] ;
 wire \Tile_X2Y6_WW4BEG[3] ;
 wire \Tile_X2Y6_WW4BEG[4] ;
 wire \Tile_X2Y6_WW4BEG[5] ;
 wire \Tile_X2Y6_WW4BEG[6] ;
 wire \Tile_X2Y6_WW4BEG[7] ;
 wire \Tile_X2Y6_WW4BEG[8] ;
 wire \Tile_X2Y6_WW4BEG[9] ;
 wire Tile_X2Y7_Co;
 wire \Tile_X2Y7_E1BEG[0] ;
 wire \Tile_X2Y7_E1BEG[1] ;
 wire \Tile_X2Y7_E1BEG[2] ;
 wire \Tile_X2Y7_E1BEG[3] ;
 wire \Tile_X2Y7_E2BEG[0] ;
 wire \Tile_X2Y7_E2BEG[1] ;
 wire \Tile_X2Y7_E2BEG[2] ;
 wire \Tile_X2Y7_E2BEG[3] ;
 wire \Tile_X2Y7_E2BEG[4] ;
 wire \Tile_X2Y7_E2BEG[5] ;
 wire \Tile_X2Y7_E2BEG[6] ;
 wire \Tile_X2Y7_E2BEG[7] ;
 wire \Tile_X2Y7_E2BEGb[0] ;
 wire \Tile_X2Y7_E2BEGb[1] ;
 wire \Tile_X2Y7_E2BEGb[2] ;
 wire \Tile_X2Y7_E2BEGb[3] ;
 wire \Tile_X2Y7_E2BEGb[4] ;
 wire \Tile_X2Y7_E2BEGb[5] ;
 wire \Tile_X2Y7_E2BEGb[6] ;
 wire \Tile_X2Y7_E2BEGb[7] ;
 wire \Tile_X2Y7_E6BEG[0] ;
 wire \Tile_X2Y7_E6BEG[10] ;
 wire \Tile_X2Y7_E6BEG[11] ;
 wire \Tile_X2Y7_E6BEG[1] ;
 wire \Tile_X2Y7_E6BEG[2] ;
 wire \Tile_X2Y7_E6BEG[3] ;
 wire \Tile_X2Y7_E6BEG[4] ;
 wire \Tile_X2Y7_E6BEG[5] ;
 wire \Tile_X2Y7_E6BEG[6] ;
 wire \Tile_X2Y7_E6BEG[7] ;
 wire \Tile_X2Y7_E6BEG[8] ;
 wire \Tile_X2Y7_E6BEG[9] ;
 wire \Tile_X2Y7_EE4BEG[0] ;
 wire \Tile_X2Y7_EE4BEG[10] ;
 wire \Tile_X2Y7_EE4BEG[11] ;
 wire \Tile_X2Y7_EE4BEG[12] ;
 wire \Tile_X2Y7_EE4BEG[13] ;
 wire \Tile_X2Y7_EE4BEG[14] ;
 wire \Tile_X2Y7_EE4BEG[15] ;
 wire \Tile_X2Y7_EE4BEG[1] ;
 wire \Tile_X2Y7_EE4BEG[2] ;
 wire \Tile_X2Y7_EE4BEG[3] ;
 wire \Tile_X2Y7_EE4BEG[4] ;
 wire \Tile_X2Y7_EE4BEG[5] ;
 wire \Tile_X2Y7_EE4BEG[6] ;
 wire \Tile_X2Y7_EE4BEG[7] ;
 wire \Tile_X2Y7_EE4BEG[8] ;
 wire \Tile_X2Y7_EE4BEG[9] ;
 wire \Tile_X2Y7_FrameData_O[0] ;
 wire \Tile_X2Y7_FrameData_O[10] ;
 wire \Tile_X2Y7_FrameData_O[11] ;
 wire \Tile_X2Y7_FrameData_O[12] ;
 wire \Tile_X2Y7_FrameData_O[13] ;
 wire \Tile_X2Y7_FrameData_O[14] ;
 wire \Tile_X2Y7_FrameData_O[15] ;
 wire \Tile_X2Y7_FrameData_O[16] ;
 wire \Tile_X2Y7_FrameData_O[17] ;
 wire \Tile_X2Y7_FrameData_O[18] ;
 wire \Tile_X2Y7_FrameData_O[19] ;
 wire \Tile_X2Y7_FrameData_O[1] ;
 wire \Tile_X2Y7_FrameData_O[20] ;
 wire \Tile_X2Y7_FrameData_O[21] ;
 wire \Tile_X2Y7_FrameData_O[22] ;
 wire \Tile_X2Y7_FrameData_O[23] ;
 wire \Tile_X2Y7_FrameData_O[24] ;
 wire \Tile_X2Y7_FrameData_O[25] ;
 wire \Tile_X2Y7_FrameData_O[26] ;
 wire \Tile_X2Y7_FrameData_O[27] ;
 wire \Tile_X2Y7_FrameData_O[28] ;
 wire \Tile_X2Y7_FrameData_O[29] ;
 wire \Tile_X2Y7_FrameData_O[2] ;
 wire \Tile_X2Y7_FrameData_O[30] ;
 wire \Tile_X2Y7_FrameData_O[31] ;
 wire \Tile_X2Y7_FrameData_O[3] ;
 wire \Tile_X2Y7_FrameData_O[4] ;
 wire \Tile_X2Y7_FrameData_O[5] ;
 wire \Tile_X2Y7_FrameData_O[6] ;
 wire \Tile_X2Y7_FrameData_O[7] ;
 wire \Tile_X2Y7_FrameData_O[8] ;
 wire \Tile_X2Y7_FrameData_O[9] ;
 wire \Tile_X2Y7_FrameStrobe_O[0] ;
 wire \Tile_X2Y7_FrameStrobe_O[10] ;
 wire \Tile_X2Y7_FrameStrobe_O[11] ;
 wire \Tile_X2Y7_FrameStrobe_O[12] ;
 wire \Tile_X2Y7_FrameStrobe_O[13] ;
 wire \Tile_X2Y7_FrameStrobe_O[14] ;
 wire \Tile_X2Y7_FrameStrobe_O[15] ;
 wire \Tile_X2Y7_FrameStrobe_O[16] ;
 wire \Tile_X2Y7_FrameStrobe_O[17] ;
 wire \Tile_X2Y7_FrameStrobe_O[18] ;
 wire \Tile_X2Y7_FrameStrobe_O[19] ;
 wire \Tile_X2Y7_FrameStrobe_O[1] ;
 wire \Tile_X2Y7_FrameStrobe_O[2] ;
 wire \Tile_X2Y7_FrameStrobe_O[3] ;
 wire \Tile_X2Y7_FrameStrobe_O[4] ;
 wire \Tile_X2Y7_FrameStrobe_O[5] ;
 wire \Tile_X2Y7_FrameStrobe_O[6] ;
 wire \Tile_X2Y7_FrameStrobe_O[7] ;
 wire \Tile_X2Y7_FrameStrobe_O[8] ;
 wire \Tile_X2Y7_FrameStrobe_O[9] ;
 wire \Tile_X2Y7_N1BEG[0] ;
 wire \Tile_X2Y7_N1BEG[1] ;
 wire \Tile_X2Y7_N1BEG[2] ;
 wire \Tile_X2Y7_N1BEG[3] ;
 wire \Tile_X2Y7_N2BEG[0] ;
 wire \Tile_X2Y7_N2BEG[1] ;
 wire \Tile_X2Y7_N2BEG[2] ;
 wire \Tile_X2Y7_N2BEG[3] ;
 wire \Tile_X2Y7_N2BEG[4] ;
 wire \Tile_X2Y7_N2BEG[5] ;
 wire \Tile_X2Y7_N2BEG[6] ;
 wire \Tile_X2Y7_N2BEG[7] ;
 wire \Tile_X2Y7_N2BEGb[0] ;
 wire \Tile_X2Y7_N2BEGb[1] ;
 wire \Tile_X2Y7_N2BEGb[2] ;
 wire \Tile_X2Y7_N2BEGb[3] ;
 wire \Tile_X2Y7_N2BEGb[4] ;
 wire \Tile_X2Y7_N2BEGb[5] ;
 wire \Tile_X2Y7_N2BEGb[6] ;
 wire \Tile_X2Y7_N2BEGb[7] ;
 wire \Tile_X2Y7_N4BEG[0] ;
 wire \Tile_X2Y7_N4BEG[10] ;
 wire \Tile_X2Y7_N4BEG[11] ;
 wire \Tile_X2Y7_N4BEG[12] ;
 wire \Tile_X2Y7_N4BEG[13] ;
 wire \Tile_X2Y7_N4BEG[14] ;
 wire \Tile_X2Y7_N4BEG[15] ;
 wire \Tile_X2Y7_N4BEG[1] ;
 wire \Tile_X2Y7_N4BEG[2] ;
 wire \Tile_X2Y7_N4BEG[3] ;
 wire \Tile_X2Y7_N4BEG[4] ;
 wire \Tile_X2Y7_N4BEG[5] ;
 wire \Tile_X2Y7_N4BEG[6] ;
 wire \Tile_X2Y7_N4BEG[7] ;
 wire \Tile_X2Y7_N4BEG[8] ;
 wire \Tile_X2Y7_N4BEG[9] ;
 wire \Tile_X2Y7_NN4BEG[0] ;
 wire \Tile_X2Y7_NN4BEG[10] ;
 wire \Tile_X2Y7_NN4BEG[11] ;
 wire \Tile_X2Y7_NN4BEG[12] ;
 wire \Tile_X2Y7_NN4BEG[13] ;
 wire \Tile_X2Y7_NN4BEG[14] ;
 wire \Tile_X2Y7_NN4BEG[15] ;
 wire \Tile_X2Y7_NN4BEG[1] ;
 wire \Tile_X2Y7_NN4BEG[2] ;
 wire \Tile_X2Y7_NN4BEG[3] ;
 wire \Tile_X2Y7_NN4BEG[4] ;
 wire \Tile_X2Y7_NN4BEG[5] ;
 wire \Tile_X2Y7_NN4BEG[6] ;
 wire \Tile_X2Y7_NN4BEG[7] ;
 wire \Tile_X2Y7_NN4BEG[8] ;
 wire \Tile_X2Y7_NN4BEG[9] ;
 wire \Tile_X2Y7_S1BEG[0] ;
 wire \Tile_X2Y7_S1BEG[1] ;
 wire \Tile_X2Y7_S1BEG[2] ;
 wire \Tile_X2Y7_S1BEG[3] ;
 wire \Tile_X2Y7_S2BEG[0] ;
 wire \Tile_X2Y7_S2BEG[1] ;
 wire \Tile_X2Y7_S2BEG[2] ;
 wire \Tile_X2Y7_S2BEG[3] ;
 wire \Tile_X2Y7_S2BEG[4] ;
 wire \Tile_X2Y7_S2BEG[5] ;
 wire \Tile_X2Y7_S2BEG[6] ;
 wire \Tile_X2Y7_S2BEG[7] ;
 wire \Tile_X2Y7_S2BEGb[0] ;
 wire \Tile_X2Y7_S2BEGb[1] ;
 wire \Tile_X2Y7_S2BEGb[2] ;
 wire \Tile_X2Y7_S2BEGb[3] ;
 wire \Tile_X2Y7_S2BEGb[4] ;
 wire \Tile_X2Y7_S2BEGb[5] ;
 wire \Tile_X2Y7_S2BEGb[6] ;
 wire \Tile_X2Y7_S2BEGb[7] ;
 wire \Tile_X2Y7_S4BEG[0] ;
 wire \Tile_X2Y7_S4BEG[10] ;
 wire \Tile_X2Y7_S4BEG[11] ;
 wire \Tile_X2Y7_S4BEG[12] ;
 wire \Tile_X2Y7_S4BEG[13] ;
 wire \Tile_X2Y7_S4BEG[14] ;
 wire \Tile_X2Y7_S4BEG[15] ;
 wire \Tile_X2Y7_S4BEG[1] ;
 wire \Tile_X2Y7_S4BEG[2] ;
 wire \Tile_X2Y7_S4BEG[3] ;
 wire \Tile_X2Y7_S4BEG[4] ;
 wire \Tile_X2Y7_S4BEG[5] ;
 wire \Tile_X2Y7_S4BEG[6] ;
 wire \Tile_X2Y7_S4BEG[7] ;
 wire \Tile_X2Y7_S4BEG[8] ;
 wire \Tile_X2Y7_S4BEG[9] ;
 wire \Tile_X2Y7_SS4BEG[0] ;
 wire \Tile_X2Y7_SS4BEG[10] ;
 wire \Tile_X2Y7_SS4BEG[11] ;
 wire \Tile_X2Y7_SS4BEG[12] ;
 wire \Tile_X2Y7_SS4BEG[13] ;
 wire \Tile_X2Y7_SS4BEG[14] ;
 wire \Tile_X2Y7_SS4BEG[15] ;
 wire \Tile_X2Y7_SS4BEG[1] ;
 wire \Tile_X2Y7_SS4BEG[2] ;
 wire \Tile_X2Y7_SS4BEG[3] ;
 wire \Tile_X2Y7_SS4BEG[4] ;
 wire \Tile_X2Y7_SS4BEG[5] ;
 wire \Tile_X2Y7_SS4BEG[6] ;
 wire \Tile_X2Y7_SS4BEG[7] ;
 wire \Tile_X2Y7_SS4BEG[8] ;
 wire \Tile_X2Y7_SS4BEG[9] ;
 wire Tile_X2Y7_UserCLKo;
 wire \Tile_X2Y7_W1BEG[0] ;
 wire \Tile_X2Y7_W1BEG[1] ;
 wire \Tile_X2Y7_W1BEG[2] ;
 wire \Tile_X2Y7_W1BEG[3] ;
 wire \Tile_X2Y7_W2BEG[0] ;
 wire \Tile_X2Y7_W2BEG[1] ;
 wire \Tile_X2Y7_W2BEG[2] ;
 wire \Tile_X2Y7_W2BEG[3] ;
 wire \Tile_X2Y7_W2BEG[4] ;
 wire \Tile_X2Y7_W2BEG[5] ;
 wire \Tile_X2Y7_W2BEG[6] ;
 wire \Tile_X2Y7_W2BEG[7] ;
 wire \Tile_X2Y7_W2BEGb[0] ;
 wire \Tile_X2Y7_W2BEGb[1] ;
 wire \Tile_X2Y7_W2BEGb[2] ;
 wire \Tile_X2Y7_W2BEGb[3] ;
 wire \Tile_X2Y7_W2BEGb[4] ;
 wire \Tile_X2Y7_W2BEGb[5] ;
 wire \Tile_X2Y7_W2BEGb[6] ;
 wire \Tile_X2Y7_W2BEGb[7] ;
 wire \Tile_X2Y7_W6BEG[0] ;
 wire \Tile_X2Y7_W6BEG[10] ;
 wire \Tile_X2Y7_W6BEG[11] ;
 wire \Tile_X2Y7_W6BEG[1] ;
 wire \Tile_X2Y7_W6BEG[2] ;
 wire \Tile_X2Y7_W6BEG[3] ;
 wire \Tile_X2Y7_W6BEG[4] ;
 wire \Tile_X2Y7_W6BEG[5] ;
 wire \Tile_X2Y7_W6BEG[6] ;
 wire \Tile_X2Y7_W6BEG[7] ;
 wire \Tile_X2Y7_W6BEG[8] ;
 wire \Tile_X2Y7_W6BEG[9] ;
 wire \Tile_X2Y7_WW4BEG[0] ;
 wire \Tile_X2Y7_WW4BEG[10] ;
 wire \Tile_X2Y7_WW4BEG[11] ;
 wire \Tile_X2Y7_WW4BEG[12] ;
 wire \Tile_X2Y7_WW4BEG[13] ;
 wire \Tile_X2Y7_WW4BEG[14] ;
 wire \Tile_X2Y7_WW4BEG[15] ;
 wire \Tile_X2Y7_WW4BEG[1] ;
 wire \Tile_X2Y7_WW4BEG[2] ;
 wire \Tile_X2Y7_WW4BEG[3] ;
 wire \Tile_X2Y7_WW4BEG[4] ;
 wire \Tile_X2Y7_WW4BEG[5] ;
 wire \Tile_X2Y7_WW4BEG[6] ;
 wire \Tile_X2Y7_WW4BEG[7] ;
 wire \Tile_X2Y7_WW4BEG[8] ;
 wire \Tile_X2Y7_WW4BEG[9] ;
 wire Tile_X2Y8_Co;
 wire \Tile_X2Y8_E1BEG[0] ;
 wire \Tile_X2Y8_E1BEG[1] ;
 wire \Tile_X2Y8_E1BEG[2] ;
 wire \Tile_X2Y8_E1BEG[3] ;
 wire \Tile_X2Y8_E2BEG[0] ;
 wire \Tile_X2Y8_E2BEG[1] ;
 wire \Tile_X2Y8_E2BEG[2] ;
 wire \Tile_X2Y8_E2BEG[3] ;
 wire \Tile_X2Y8_E2BEG[4] ;
 wire \Tile_X2Y8_E2BEG[5] ;
 wire \Tile_X2Y8_E2BEG[6] ;
 wire \Tile_X2Y8_E2BEG[7] ;
 wire \Tile_X2Y8_E2BEGb[0] ;
 wire \Tile_X2Y8_E2BEGb[1] ;
 wire \Tile_X2Y8_E2BEGb[2] ;
 wire \Tile_X2Y8_E2BEGb[3] ;
 wire \Tile_X2Y8_E2BEGb[4] ;
 wire \Tile_X2Y8_E2BEGb[5] ;
 wire \Tile_X2Y8_E2BEGb[6] ;
 wire \Tile_X2Y8_E2BEGb[7] ;
 wire \Tile_X2Y8_E6BEG[0] ;
 wire \Tile_X2Y8_E6BEG[10] ;
 wire \Tile_X2Y8_E6BEG[11] ;
 wire \Tile_X2Y8_E6BEG[1] ;
 wire \Tile_X2Y8_E6BEG[2] ;
 wire \Tile_X2Y8_E6BEG[3] ;
 wire \Tile_X2Y8_E6BEG[4] ;
 wire \Tile_X2Y8_E6BEG[5] ;
 wire \Tile_X2Y8_E6BEG[6] ;
 wire \Tile_X2Y8_E6BEG[7] ;
 wire \Tile_X2Y8_E6BEG[8] ;
 wire \Tile_X2Y8_E6BEG[9] ;
 wire \Tile_X2Y8_EE4BEG[0] ;
 wire \Tile_X2Y8_EE4BEG[10] ;
 wire \Tile_X2Y8_EE4BEG[11] ;
 wire \Tile_X2Y8_EE4BEG[12] ;
 wire \Tile_X2Y8_EE4BEG[13] ;
 wire \Tile_X2Y8_EE4BEG[14] ;
 wire \Tile_X2Y8_EE4BEG[15] ;
 wire \Tile_X2Y8_EE4BEG[1] ;
 wire \Tile_X2Y8_EE4BEG[2] ;
 wire \Tile_X2Y8_EE4BEG[3] ;
 wire \Tile_X2Y8_EE4BEG[4] ;
 wire \Tile_X2Y8_EE4BEG[5] ;
 wire \Tile_X2Y8_EE4BEG[6] ;
 wire \Tile_X2Y8_EE4BEG[7] ;
 wire \Tile_X2Y8_EE4BEG[8] ;
 wire \Tile_X2Y8_EE4BEG[9] ;
 wire \Tile_X2Y8_FrameData_O[0] ;
 wire \Tile_X2Y8_FrameData_O[10] ;
 wire \Tile_X2Y8_FrameData_O[11] ;
 wire \Tile_X2Y8_FrameData_O[12] ;
 wire \Tile_X2Y8_FrameData_O[13] ;
 wire \Tile_X2Y8_FrameData_O[14] ;
 wire \Tile_X2Y8_FrameData_O[15] ;
 wire \Tile_X2Y8_FrameData_O[16] ;
 wire \Tile_X2Y8_FrameData_O[17] ;
 wire \Tile_X2Y8_FrameData_O[18] ;
 wire \Tile_X2Y8_FrameData_O[19] ;
 wire \Tile_X2Y8_FrameData_O[1] ;
 wire \Tile_X2Y8_FrameData_O[20] ;
 wire \Tile_X2Y8_FrameData_O[21] ;
 wire \Tile_X2Y8_FrameData_O[22] ;
 wire \Tile_X2Y8_FrameData_O[23] ;
 wire \Tile_X2Y8_FrameData_O[24] ;
 wire \Tile_X2Y8_FrameData_O[25] ;
 wire \Tile_X2Y8_FrameData_O[26] ;
 wire \Tile_X2Y8_FrameData_O[27] ;
 wire \Tile_X2Y8_FrameData_O[28] ;
 wire \Tile_X2Y8_FrameData_O[29] ;
 wire \Tile_X2Y8_FrameData_O[2] ;
 wire \Tile_X2Y8_FrameData_O[30] ;
 wire \Tile_X2Y8_FrameData_O[31] ;
 wire \Tile_X2Y8_FrameData_O[3] ;
 wire \Tile_X2Y8_FrameData_O[4] ;
 wire \Tile_X2Y8_FrameData_O[5] ;
 wire \Tile_X2Y8_FrameData_O[6] ;
 wire \Tile_X2Y8_FrameData_O[7] ;
 wire \Tile_X2Y8_FrameData_O[8] ;
 wire \Tile_X2Y8_FrameData_O[9] ;
 wire \Tile_X2Y8_FrameStrobe_O[0] ;
 wire \Tile_X2Y8_FrameStrobe_O[10] ;
 wire \Tile_X2Y8_FrameStrobe_O[11] ;
 wire \Tile_X2Y8_FrameStrobe_O[12] ;
 wire \Tile_X2Y8_FrameStrobe_O[13] ;
 wire \Tile_X2Y8_FrameStrobe_O[14] ;
 wire \Tile_X2Y8_FrameStrobe_O[15] ;
 wire \Tile_X2Y8_FrameStrobe_O[16] ;
 wire \Tile_X2Y8_FrameStrobe_O[17] ;
 wire \Tile_X2Y8_FrameStrobe_O[18] ;
 wire \Tile_X2Y8_FrameStrobe_O[19] ;
 wire \Tile_X2Y8_FrameStrobe_O[1] ;
 wire \Tile_X2Y8_FrameStrobe_O[2] ;
 wire \Tile_X2Y8_FrameStrobe_O[3] ;
 wire \Tile_X2Y8_FrameStrobe_O[4] ;
 wire \Tile_X2Y8_FrameStrobe_O[5] ;
 wire \Tile_X2Y8_FrameStrobe_O[6] ;
 wire \Tile_X2Y8_FrameStrobe_O[7] ;
 wire \Tile_X2Y8_FrameStrobe_O[8] ;
 wire \Tile_X2Y8_FrameStrobe_O[9] ;
 wire \Tile_X2Y8_N1BEG[0] ;
 wire \Tile_X2Y8_N1BEG[1] ;
 wire \Tile_X2Y8_N1BEG[2] ;
 wire \Tile_X2Y8_N1BEG[3] ;
 wire \Tile_X2Y8_N2BEG[0] ;
 wire \Tile_X2Y8_N2BEG[1] ;
 wire \Tile_X2Y8_N2BEG[2] ;
 wire \Tile_X2Y8_N2BEG[3] ;
 wire \Tile_X2Y8_N2BEG[4] ;
 wire \Tile_X2Y8_N2BEG[5] ;
 wire \Tile_X2Y8_N2BEG[6] ;
 wire \Tile_X2Y8_N2BEG[7] ;
 wire \Tile_X2Y8_N2BEGb[0] ;
 wire \Tile_X2Y8_N2BEGb[1] ;
 wire \Tile_X2Y8_N2BEGb[2] ;
 wire \Tile_X2Y8_N2BEGb[3] ;
 wire \Tile_X2Y8_N2BEGb[4] ;
 wire \Tile_X2Y8_N2BEGb[5] ;
 wire \Tile_X2Y8_N2BEGb[6] ;
 wire \Tile_X2Y8_N2BEGb[7] ;
 wire \Tile_X2Y8_N4BEG[0] ;
 wire \Tile_X2Y8_N4BEG[10] ;
 wire \Tile_X2Y8_N4BEG[11] ;
 wire \Tile_X2Y8_N4BEG[12] ;
 wire \Tile_X2Y8_N4BEG[13] ;
 wire \Tile_X2Y8_N4BEG[14] ;
 wire \Tile_X2Y8_N4BEG[15] ;
 wire \Tile_X2Y8_N4BEG[1] ;
 wire \Tile_X2Y8_N4BEG[2] ;
 wire \Tile_X2Y8_N4BEG[3] ;
 wire \Tile_X2Y8_N4BEG[4] ;
 wire \Tile_X2Y8_N4BEG[5] ;
 wire \Tile_X2Y8_N4BEG[6] ;
 wire \Tile_X2Y8_N4BEG[7] ;
 wire \Tile_X2Y8_N4BEG[8] ;
 wire \Tile_X2Y8_N4BEG[9] ;
 wire \Tile_X2Y8_NN4BEG[0] ;
 wire \Tile_X2Y8_NN4BEG[10] ;
 wire \Tile_X2Y8_NN4BEG[11] ;
 wire \Tile_X2Y8_NN4BEG[12] ;
 wire \Tile_X2Y8_NN4BEG[13] ;
 wire \Tile_X2Y8_NN4BEG[14] ;
 wire \Tile_X2Y8_NN4BEG[15] ;
 wire \Tile_X2Y8_NN4BEG[1] ;
 wire \Tile_X2Y8_NN4BEG[2] ;
 wire \Tile_X2Y8_NN4BEG[3] ;
 wire \Tile_X2Y8_NN4BEG[4] ;
 wire \Tile_X2Y8_NN4BEG[5] ;
 wire \Tile_X2Y8_NN4BEG[6] ;
 wire \Tile_X2Y8_NN4BEG[7] ;
 wire \Tile_X2Y8_NN4BEG[8] ;
 wire \Tile_X2Y8_NN4BEG[9] ;
 wire \Tile_X2Y8_S1BEG[0] ;
 wire \Tile_X2Y8_S1BEG[1] ;
 wire \Tile_X2Y8_S1BEG[2] ;
 wire \Tile_X2Y8_S1BEG[3] ;
 wire \Tile_X2Y8_S2BEG[0] ;
 wire \Tile_X2Y8_S2BEG[1] ;
 wire \Tile_X2Y8_S2BEG[2] ;
 wire \Tile_X2Y8_S2BEG[3] ;
 wire \Tile_X2Y8_S2BEG[4] ;
 wire \Tile_X2Y8_S2BEG[5] ;
 wire \Tile_X2Y8_S2BEG[6] ;
 wire \Tile_X2Y8_S2BEG[7] ;
 wire \Tile_X2Y8_S2BEGb[0] ;
 wire \Tile_X2Y8_S2BEGb[1] ;
 wire \Tile_X2Y8_S2BEGb[2] ;
 wire \Tile_X2Y8_S2BEGb[3] ;
 wire \Tile_X2Y8_S2BEGb[4] ;
 wire \Tile_X2Y8_S2BEGb[5] ;
 wire \Tile_X2Y8_S2BEGb[6] ;
 wire \Tile_X2Y8_S2BEGb[7] ;
 wire \Tile_X2Y8_S4BEG[0] ;
 wire \Tile_X2Y8_S4BEG[10] ;
 wire \Tile_X2Y8_S4BEG[11] ;
 wire \Tile_X2Y8_S4BEG[12] ;
 wire \Tile_X2Y8_S4BEG[13] ;
 wire \Tile_X2Y8_S4BEG[14] ;
 wire \Tile_X2Y8_S4BEG[15] ;
 wire \Tile_X2Y8_S4BEG[1] ;
 wire \Tile_X2Y8_S4BEG[2] ;
 wire \Tile_X2Y8_S4BEG[3] ;
 wire \Tile_X2Y8_S4BEG[4] ;
 wire \Tile_X2Y8_S4BEG[5] ;
 wire \Tile_X2Y8_S4BEG[6] ;
 wire \Tile_X2Y8_S4BEG[7] ;
 wire \Tile_X2Y8_S4BEG[8] ;
 wire \Tile_X2Y8_S4BEG[9] ;
 wire \Tile_X2Y8_SS4BEG[0] ;
 wire \Tile_X2Y8_SS4BEG[10] ;
 wire \Tile_X2Y8_SS4BEG[11] ;
 wire \Tile_X2Y8_SS4BEG[12] ;
 wire \Tile_X2Y8_SS4BEG[13] ;
 wire \Tile_X2Y8_SS4BEG[14] ;
 wire \Tile_X2Y8_SS4BEG[15] ;
 wire \Tile_X2Y8_SS4BEG[1] ;
 wire \Tile_X2Y8_SS4BEG[2] ;
 wire \Tile_X2Y8_SS4BEG[3] ;
 wire \Tile_X2Y8_SS4BEG[4] ;
 wire \Tile_X2Y8_SS4BEG[5] ;
 wire \Tile_X2Y8_SS4BEG[6] ;
 wire \Tile_X2Y8_SS4BEG[7] ;
 wire \Tile_X2Y8_SS4BEG[8] ;
 wire \Tile_X2Y8_SS4BEG[9] ;
 wire Tile_X2Y8_UserCLKo;
 wire \Tile_X2Y8_W1BEG[0] ;
 wire \Tile_X2Y8_W1BEG[1] ;
 wire \Tile_X2Y8_W1BEG[2] ;
 wire \Tile_X2Y8_W1BEG[3] ;
 wire \Tile_X2Y8_W2BEG[0] ;
 wire \Tile_X2Y8_W2BEG[1] ;
 wire \Tile_X2Y8_W2BEG[2] ;
 wire \Tile_X2Y8_W2BEG[3] ;
 wire \Tile_X2Y8_W2BEG[4] ;
 wire \Tile_X2Y8_W2BEG[5] ;
 wire \Tile_X2Y8_W2BEG[6] ;
 wire \Tile_X2Y8_W2BEG[7] ;
 wire \Tile_X2Y8_W2BEGb[0] ;
 wire \Tile_X2Y8_W2BEGb[1] ;
 wire \Tile_X2Y8_W2BEGb[2] ;
 wire \Tile_X2Y8_W2BEGb[3] ;
 wire \Tile_X2Y8_W2BEGb[4] ;
 wire \Tile_X2Y8_W2BEGb[5] ;
 wire \Tile_X2Y8_W2BEGb[6] ;
 wire \Tile_X2Y8_W2BEGb[7] ;
 wire \Tile_X2Y8_W6BEG[0] ;
 wire \Tile_X2Y8_W6BEG[10] ;
 wire \Tile_X2Y8_W6BEG[11] ;
 wire \Tile_X2Y8_W6BEG[1] ;
 wire \Tile_X2Y8_W6BEG[2] ;
 wire \Tile_X2Y8_W6BEG[3] ;
 wire \Tile_X2Y8_W6BEG[4] ;
 wire \Tile_X2Y8_W6BEG[5] ;
 wire \Tile_X2Y8_W6BEG[6] ;
 wire \Tile_X2Y8_W6BEG[7] ;
 wire \Tile_X2Y8_W6BEG[8] ;
 wire \Tile_X2Y8_W6BEG[9] ;
 wire \Tile_X2Y8_WW4BEG[0] ;
 wire \Tile_X2Y8_WW4BEG[10] ;
 wire \Tile_X2Y8_WW4BEG[11] ;
 wire \Tile_X2Y8_WW4BEG[12] ;
 wire \Tile_X2Y8_WW4BEG[13] ;
 wire \Tile_X2Y8_WW4BEG[14] ;
 wire \Tile_X2Y8_WW4BEG[15] ;
 wire \Tile_X2Y8_WW4BEG[1] ;
 wire \Tile_X2Y8_WW4BEG[2] ;
 wire \Tile_X2Y8_WW4BEG[3] ;
 wire \Tile_X2Y8_WW4BEG[4] ;
 wire \Tile_X2Y8_WW4BEG[5] ;
 wire \Tile_X2Y8_WW4BEG[6] ;
 wire \Tile_X2Y8_WW4BEG[7] ;
 wire \Tile_X2Y8_WW4BEG[8] ;
 wire \Tile_X2Y8_WW4BEG[9] ;
 wire Tile_X2Y9_Co;
 wire \Tile_X2Y9_FrameData_O[0] ;
 wire \Tile_X2Y9_FrameData_O[10] ;
 wire \Tile_X2Y9_FrameData_O[11] ;
 wire \Tile_X2Y9_FrameData_O[12] ;
 wire \Tile_X2Y9_FrameData_O[13] ;
 wire \Tile_X2Y9_FrameData_O[14] ;
 wire \Tile_X2Y9_FrameData_O[15] ;
 wire \Tile_X2Y9_FrameData_O[16] ;
 wire \Tile_X2Y9_FrameData_O[17] ;
 wire \Tile_X2Y9_FrameData_O[18] ;
 wire \Tile_X2Y9_FrameData_O[19] ;
 wire \Tile_X2Y9_FrameData_O[1] ;
 wire \Tile_X2Y9_FrameData_O[20] ;
 wire \Tile_X2Y9_FrameData_O[21] ;
 wire \Tile_X2Y9_FrameData_O[22] ;
 wire \Tile_X2Y9_FrameData_O[23] ;
 wire \Tile_X2Y9_FrameData_O[24] ;
 wire \Tile_X2Y9_FrameData_O[25] ;
 wire \Tile_X2Y9_FrameData_O[26] ;
 wire \Tile_X2Y9_FrameData_O[27] ;
 wire \Tile_X2Y9_FrameData_O[28] ;
 wire \Tile_X2Y9_FrameData_O[29] ;
 wire \Tile_X2Y9_FrameData_O[2] ;
 wire \Tile_X2Y9_FrameData_O[30] ;
 wire \Tile_X2Y9_FrameData_O[31] ;
 wire \Tile_X2Y9_FrameData_O[3] ;
 wire \Tile_X2Y9_FrameData_O[4] ;
 wire \Tile_X2Y9_FrameData_O[5] ;
 wire \Tile_X2Y9_FrameData_O[6] ;
 wire \Tile_X2Y9_FrameData_O[7] ;
 wire \Tile_X2Y9_FrameData_O[8] ;
 wire \Tile_X2Y9_FrameData_O[9] ;
 wire \Tile_X2Y9_FrameStrobe_O[0] ;
 wire \Tile_X2Y9_FrameStrobe_O[10] ;
 wire \Tile_X2Y9_FrameStrobe_O[11] ;
 wire \Tile_X2Y9_FrameStrobe_O[12] ;
 wire \Tile_X2Y9_FrameStrobe_O[13] ;
 wire \Tile_X2Y9_FrameStrobe_O[14] ;
 wire \Tile_X2Y9_FrameStrobe_O[15] ;
 wire \Tile_X2Y9_FrameStrobe_O[16] ;
 wire \Tile_X2Y9_FrameStrobe_O[17] ;
 wire \Tile_X2Y9_FrameStrobe_O[18] ;
 wire \Tile_X2Y9_FrameStrobe_O[19] ;
 wire \Tile_X2Y9_FrameStrobe_O[1] ;
 wire \Tile_X2Y9_FrameStrobe_O[2] ;
 wire \Tile_X2Y9_FrameStrobe_O[3] ;
 wire \Tile_X2Y9_FrameStrobe_O[4] ;
 wire \Tile_X2Y9_FrameStrobe_O[5] ;
 wire \Tile_X2Y9_FrameStrobe_O[6] ;
 wire \Tile_X2Y9_FrameStrobe_O[7] ;
 wire \Tile_X2Y9_FrameStrobe_O[8] ;
 wire \Tile_X2Y9_FrameStrobe_O[9] ;
 wire \Tile_X2Y9_N1BEG[0] ;
 wire \Tile_X2Y9_N1BEG[1] ;
 wire \Tile_X2Y9_N1BEG[2] ;
 wire \Tile_X2Y9_N1BEG[3] ;
 wire \Tile_X2Y9_N2BEG[0] ;
 wire \Tile_X2Y9_N2BEG[1] ;
 wire \Tile_X2Y9_N2BEG[2] ;
 wire \Tile_X2Y9_N2BEG[3] ;
 wire \Tile_X2Y9_N2BEG[4] ;
 wire \Tile_X2Y9_N2BEG[5] ;
 wire \Tile_X2Y9_N2BEG[6] ;
 wire \Tile_X2Y9_N2BEG[7] ;
 wire \Tile_X2Y9_N2BEGb[0] ;
 wire \Tile_X2Y9_N2BEGb[1] ;
 wire \Tile_X2Y9_N2BEGb[2] ;
 wire \Tile_X2Y9_N2BEGb[3] ;
 wire \Tile_X2Y9_N2BEGb[4] ;
 wire \Tile_X2Y9_N2BEGb[5] ;
 wire \Tile_X2Y9_N2BEGb[6] ;
 wire \Tile_X2Y9_N2BEGb[7] ;
 wire \Tile_X2Y9_N4BEG[0] ;
 wire \Tile_X2Y9_N4BEG[10] ;
 wire \Tile_X2Y9_N4BEG[11] ;
 wire \Tile_X2Y9_N4BEG[12] ;
 wire \Tile_X2Y9_N4BEG[13] ;
 wire \Tile_X2Y9_N4BEG[14] ;
 wire \Tile_X2Y9_N4BEG[15] ;
 wire \Tile_X2Y9_N4BEG[1] ;
 wire \Tile_X2Y9_N4BEG[2] ;
 wire \Tile_X2Y9_N4BEG[3] ;
 wire \Tile_X2Y9_N4BEG[4] ;
 wire \Tile_X2Y9_N4BEG[5] ;
 wire \Tile_X2Y9_N4BEG[6] ;
 wire \Tile_X2Y9_N4BEG[7] ;
 wire \Tile_X2Y9_N4BEG[8] ;
 wire \Tile_X2Y9_N4BEG[9] ;
 wire \Tile_X2Y9_NN4BEG[0] ;
 wire \Tile_X2Y9_NN4BEG[10] ;
 wire \Tile_X2Y9_NN4BEG[11] ;
 wire \Tile_X2Y9_NN4BEG[12] ;
 wire \Tile_X2Y9_NN4BEG[13] ;
 wire \Tile_X2Y9_NN4BEG[14] ;
 wire \Tile_X2Y9_NN4BEG[15] ;
 wire \Tile_X2Y9_NN4BEG[1] ;
 wire \Tile_X2Y9_NN4BEG[2] ;
 wire \Tile_X2Y9_NN4BEG[3] ;
 wire \Tile_X2Y9_NN4BEG[4] ;
 wire \Tile_X2Y9_NN4BEG[5] ;
 wire \Tile_X2Y9_NN4BEG[6] ;
 wire \Tile_X2Y9_NN4BEG[7] ;
 wire \Tile_X2Y9_NN4BEG[8] ;
 wire \Tile_X2Y9_NN4BEG[9] ;
 wire Tile_X2Y9_UserCLKo;
 wire \Tile_X3Y0_FrameData_O[0] ;
 wire \Tile_X3Y0_FrameData_O[10] ;
 wire \Tile_X3Y0_FrameData_O[11] ;
 wire \Tile_X3Y0_FrameData_O[12] ;
 wire \Tile_X3Y0_FrameData_O[13] ;
 wire \Tile_X3Y0_FrameData_O[14] ;
 wire \Tile_X3Y0_FrameData_O[15] ;
 wire \Tile_X3Y0_FrameData_O[16] ;
 wire \Tile_X3Y0_FrameData_O[17] ;
 wire \Tile_X3Y0_FrameData_O[18] ;
 wire \Tile_X3Y0_FrameData_O[19] ;
 wire \Tile_X3Y0_FrameData_O[1] ;
 wire \Tile_X3Y0_FrameData_O[20] ;
 wire \Tile_X3Y0_FrameData_O[21] ;
 wire \Tile_X3Y0_FrameData_O[22] ;
 wire \Tile_X3Y0_FrameData_O[23] ;
 wire \Tile_X3Y0_FrameData_O[24] ;
 wire \Tile_X3Y0_FrameData_O[25] ;
 wire \Tile_X3Y0_FrameData_O[26] ;
 wire \Tile_X3Y0_FrameData_O[27] ;
 wire \Tile_X3Y0_FrameData_O[28] ;
 wire \Tile_X3Y0_FrameData_O[29] ;
 wire \Tile_X3Y0_FrameData_O[2] ;
 wire \Tile_X3Y0_FrameData_O[30] ;
 wire \Tile_X3Y0_FrameData_O[31] ;
 wire \Tile_X3Y0_FrameData_O[3] ;
 wire \Tile_X3Y0_FrameData_O[4] ;
 wire \Tile_X3Y0_FrameData_O[5] ;
 wire \Tile_X3Y0_FrameData_O[6] ;
 wire \Tile_X3Y0_FrameData_O[7] ;
 wire \Tile_X3Y0_FrameData_O[8] ;
 wire \Tile_X3Y0_FrameData_O[9] ;
 wire \Tile_X3Y0_FrameStrobe_O[0] ;
 wire \Tile_X3Y0_FrameStrobe_O[10] ;
 wire \Tile_X3Y0_FrameStrobe_O[11] ;
 wire \Tile_X3Y0_FrameStrobe_O[12] ;
 wire \Tile_X3Y0_FrameStrobe_O[13] ;
 wire \Tile_X3Y0_FrameStrobe_O[14] ;
 wire \Tile_X3Y0_FrameStrobe_O[15] ;
 wire \Tile_X3Y0_FrameStrobe_O[16] ;
 wire \Tile_X3Y0_FrameStrobe_O[17] ;
 wire \Tile_X3Y0_FrameStrobe_O[18] ;
 wire \Tile_X3Y0_FrameStrobe_O[19] ;
 wire \Tile_X3Y0_FrameStrobe_O[1] ;
 wire \Tile_X3Y0_FrameStrobe_O[2] ;
 wire \Tile_X3Y0_FrameStrobe_O[3] ;
 wire \Tile_X3Y0_FrameStrobe_O[4] ;
 wire \Tile_X3Y0_FrameStrobe_O[5] ;
 wire \Tile_X3Y0_FrameStrobe_O[6] ;
 wire \Tile_X3Y0_FrameStrobe_O[7] ;
 wire \Tile_X3Y0_FrameStrobe_O[8] ;
 wire \Tile_X3Y0_FrameStrobe_O[9] ;
 wire \Tile_X3Y0_S1BEG[0] ;
 wire \Tile_X3Y0_S1BEG[1] ;
 wire \Tile_X3Y0_S1BEG[2] ;
 wire \Tile_X3Y0_S1BEG[3] ;
 wire \Tile_X3Y0_S2BEG[0] ;
 wire \Tile_X3Y0_S2BEG[1] ;
 wire \Tile_X3Y0_S2BEG[2] ;
 wire \Tile_X3Y0_S2BEG[3] ;
 wire \Tile_X3Y0_S2BEG[4] ;
 wire \Tile_X3Y0_S2BEG[5] ;
 wire \Tile_X3Y0_S2BEG[6] ;
 wire \Tile_X3Y0_S2BEG[7] ;
 wire \Tile_X3Y0_S2BEGb[0] ;
 wire \Tile_X3Y0_S2BEGb[1] ;
 wire \Tile_X3Y0_S2BEGb[2] ;
 wire \Tile_X3Y0_S2BEGb[3] ;
 wire \Tile_X3Y0_S2BEGb[4] ;
 wire \Tile_X3Y0_S2BEGb[5] ;
 wire \Tile_X3Y0_S2BEGb[6] ;
 wire \Tile_X3Y0_S2BEGb[7] ;
 wire \Tile_X3Y0_S4BEG[0] ;
 wire \Tile_X3Y0_S4BEG[10] ;
 wire \Tile_X3Y0_S4BEG[11] ;
 wire \Tile_X3Y0_S4BEG[12] ;
 wire \Tile_X3Y0_S4BEG[13] ;
 wire \Tile_X3Y0_S4BEG[14] ;
 wire \Tile_X3Y0_S4BEG[15] ;
 wire \Tile_X3Y0_S4BEG[1] ;
 wire \Tile_X3Y0_S4BEG[2] ;
 wire \Tile_X3Y0_S4BEG[3] ;
 wire \Tile_X3Y0_S4BEG[4] ;
 wire \Tile_X3Y0_S4BEG[5] ;
 wire \Tile_X3Y0_S4BEG[6] ;
 wire \Tile_X3Y0_S4BEG[7] ;
 wire \Tile_X3Y0_S4BEG[8] ;
 wire \Tile_X3Y0_S4BEG[9] ;
 wire \Tile_X3Y0_SS4BEG[0] ;
 wire \Tile_X3Y0_SS4BEG[10] ;
 wire \Tile_X3Y0_SS4BEG[11] ;
 wire \Tile_X3Y0_SS4BEG[12] ;
 wire \Tile_X3Y0_SS4BEG[13] ;
 wire \Tile_X3Y0_SS4BEG[14] ;
 wire \Tile_X3Y0_SS4BEG[15] ;
 wire \Tile_X3Y0_SS4BEG[1] ;
 wire \Tile_X3Y0_SS4BEG[2] ;
 wire \Tile_X3Y0_SS4BEG[3] ;
 wire \Tile_X3Y0_SS4BEG[4] ;
 wire \Tile_X3Y0_SS4BEG[5] ;
 wire \Tile_X3Y0_SS4BEG[6] ;
 wire \Tile_X3Y0_SS4BEG[7] ;
 wire \Tile_X3Y0_SS4BEG[8] ;
 wire \Tile_X3Y0_SS4BEG[9] ;
 wire Tile_X3Y0_UserCLKo;
 wire Tile_X3Y1_Co;
 wire \Tile_X3Y1_E1BEG[0] ;
 wire \Tile_X3Y1_E1BEG[1] ;
 wire \Tile_X3Y1_E1BEG[2] ;
 wire \Tile_X3Y1_E1BEG[3] ;
 wire \Tile_X3Y1_E2BEG[0] ;
 wire \Tile_X3Y1_E2BEG[1] ;
 wire \Tile_X3Y1_E2BEG[2] ;
 wire \Tile_X3Y1_E2BEG[3] ;
 wire \Tile_X3Y1_E2BEG[4] ;
 wire \Tile_X3Y1_E2BEG[5] ;
 wire \Tile_X3Y1_E2BEG[6] ;
 wire \Tile_X3Y1_E2BEG[7] ;
 wire \Tile_X3Y1_E2BEGb[0] ;
 wire \Tile_X3Y1_E2BEGb[1] ;
 wire \Tile_X3Y1_E2BEGb[2] ;
 wire \Tile_X3Y1_E2BEGb[3] ;
 wire \Tile_X3Y1_E2BEGb[4] ;
 wire \Tile_X3Y1_E2BEGb[5] ;
 wire \Tile_X3Y1_E2BEGb[6] ;
 wire \Tile_X3Y1_E2BEGb[7] ;
 wire \Tile_X3Y1_E6BEG[0] ;
 wire \Tile_X3Y1_E6BEG[10] ;
 wire \Tile_X3Y1_E6BEG[11] ;
 wire \Tile_X3Y1_E6BEG[1] ;
 wire \Tile_X3Y1_E6BEG[2] ;
 wire \Tile_X3Y1_E6BEG[3] ;
 wire \Tile_X3Y1_E6BEG[4] ;
 wire \Tile_X3Y1_E6BEG[5] ;
 wire \Tile_X3Y1_E6BEG[6] ;
 wire \Tile_X3Y1_E6BEG[7] ;
 wire \Tile_X3Y1_E6BEG[8] ;
 wire \Tile_X3Y1_E6BEG[9] ;
 wire \Tile_X3Y1_EE4BEG[0] ;
 wire \Tile_X3Y1_EE4BEG[10] ;
 wire \Tile_X3Y1_EE4BEG[11] ;
 wire \Tile_X3Y1_EE4BEG[12] ;
 wire \Tile_X3Y1_EE4BEG[13] ;
 wire \Tile_X3Y1_EE4BEG[14] ;
 wire \Tile_X3Y1_EE4BEG[15] ;
 wire \Tile_X3Y1_EE4BEG[1] ;
 wire \Tile_X3Y1_EE4BEG[2] ;
 wire \Tile_X3Y1_EE4BEG[3] ;
 wire \Tile_X3Y1_EE4BEG[4] ;
 wire \Tile_X3Y1_EE4BEG[5] ;
 wire \Tile_X3Y1_EE4BEG[6] ;
 wire \Tile_X3Y1_EE4BEG[7] ;
 wire \Tile_X3Y1_EE4BEG[8] ;
 wire \Tile_X3Y1_EE4BEG[9] ;
 wire \Tile_X3Y1_FrameData_O[0] ;
 wire \Tile_X3Y1_FrameData_O[10] ;
 wire \Tile_X3Y1_FrameData_O[11] ;
 wire \Tile_X3Y1_FrameData_O[12] ;
 wire \Tile_X3Y1_FrameData_O[13] ;
 wire \Tile_X3Y1_FrameData_O[14] ;
 wire \Tile_X3Y1_FrameData_O[15] ;
 wire \Tile_X3Y1_FrameData_O[16] ;
 wire \Tile_X3Y1_FrameData_O[17] ;
 wire \Tile_X3Y1_FrameData_O[18] ;
 wire \Tile_X3Y1_FrameData_O[19] ;
 wire \Tile_X3Y1_FrameData_O[1] ;
 wire \Tile_X3Y1_FrameData_O[20] ;
 wire \Tile_X3Y1_FrameData_O[21] ;
 wire \Tile_X3Y1_FrameData_O[22] ;
 wire \Tile_X3Y1_FrameData_O[23] ;
 wire \Tile_X3Y1_FrameData_O[24] ;
 wire \Tile_X3Y1_FrameData_O[25] ;
 wire \Tile_X3Y1_FrameData_O[26] ;
 wire \Tile_X3Y1_FrameData_O[27] ;
 wire \Tile_X3Y1_FrameData_O[28] ;
 wire \Tile_X3Y1_FrameData_O[29] ;
 wire \Tile_X3Y1_FrameData_O[2] ;
 wire \Tile_X3Y1_FrameData_O[30] ;
 wire \Tile_X3Y1_FrameData_O[31] ;
 wire \Tile_X3Y1_FrameData_O[3] ;
 wire \Tile_X3Y1_FrameData_O[4] ;
 wire \Tile_X3Y1_FrameData_O[5] ;
 wire \Tile_X3Y1_FrameData_O[6] ;
 wire \Tile_X3Y1_FrameData_O[7] ;
 wire \Tile_X3Y1_FrameData_O[8] ;
 wire \Tile_X3Y1_FrameData_O[9] ;
 wire \Tile_X3Y1_FrameStrobe_O[0] ;
 wire \Tile_X3Y1_FrameStrobe_O[10] ;
 wire \Tile_X3Y1_FrameStrobe_O[11] ;
 wire \Tile_X3Y1_FrameStrobe_O[12] ;
 wire \Tile_X3Y1_FrameStrobe_O[13] ;
 wire \Tile_X3Y1_FrameStrobe_O[14] ;
 wire \Tile_X3Y1_FrameStrobe_O[15] ;
 wire \Tile_X3Y1_FrameStrobe_O[16] ;
 wire \Tile_X3Y1_FrameStrobe_O[17] ;
 wire \Tile_X3Y1_FrameStrobe_O[18] ;
 wire \Tile_X3Y1_FrameStrobe_O[19] ;
 wire \Tile_X3Y1_FrameStrobe_O[1] ;
 wire \Tile_X3Y1_FrameStrobe_O[2] ;
 wire \Tile_X3Y1_FrameStrobe_O[3] ;
 wire \Tile_X3Y1_FrameStrobe_O[4] ;
 wire \Tile_X3Y1_FrameStrobe_O[5] ;
 wire \Tile_X3Y1_FrameStrobe_O[6] ;
 wire \Tile_X3Y1_FrameStrobe_O[7] ;
 wire \Tile_X3Y1_FrameStrobe_O[8] ;
 wire \Tile_X3Y1_FrameStrobe_O[9] ;
 wire \Tile_X3Y1_N1BEG[0] ;
 wire \Tile_X3Y1_N1BEG[1] ;
 wire \Tile_X3Y1_N1BEG[2] ;
 wire \Tile_X3Y1_N1BEG[3] ;
 wire \Tile_X3Y1_N2BEG[0] ;
 wire \Tile_X3Y1_N2BEG[1] ;
 wire \Tile_X3Y1_N2BEG[2] ;
 wire \Tile_X3Y1_N2BEG[3] ;
 wire \Tile_X3Y1_N2BEG[4] ;
 wire \Tile_X3Y1_N2BEG[5] ;
 wire \Tile_X3Y1_N2BEG[6] ;
 wire \Tile_X3Y1_N2BEG[7] ;
 wire \Tile_X3Y1_N2BEGb[0] ;
 wire \Tile_X3Y1_N2BEGb[1] ;
 wire \Tile_X3Y1_N2BEGb[2] ;
 wire \Tile_X3Y1_N2BEGb[3] ;
 wire \Tile_X3Y1_N2BEGb[4] ;
 wire \Tile_X3Y1_N2BEGb[5] ;
 wire \Tile_X3Y1_N2BEGb[6] ;
 wire \Tile_X3Y1_N2BEGb[7] ;
 wire \Tile_X3Y1_N4BEG[0] ;
 wire \Tile_X3Y1_N4BEG[10] ;
 wire \Tile_X3Y1_N4BEG[11] ;
 wire \Tile_X3Y1_N4BEG[12] ;
 wire \Tile_X3Y1_N4BEG[13] ;
 wire \Tile_X3Y1_N4BEG[14] ;
 wire \Tile_X3Y1_N4BEG[15] ;
 wire \Tile_X3Y1_N4BEG[1] ;
 wire \Tile_X3Y1_N4BEG[2] ;
 wire \Tile_X3Y1_N4BEG[3] ;
 wire \Tile_X3Y1_N4BEG[4] ;
 wire \Tile_X3Y1_N4BEG[5] ;
 wire \Tile_X3Y1_N4BEG[6] ;
 wire \Tile_X3Y1_N4BEG[7] ;
 wire \Tile_X3Y1_N4BEG[8] ;
 wire \Tile_X3Y1_N4BEG[9] ;
 wire \Tile_X3Y1_NN4BEG[0] ;
 wire \Tile_X3Y1_NN4BEG[10] ;
 wire \Tile_X3Y1_NN4BEG[11] ;
 wire \Tile_X3Y1_NN4BEG[12] ;
 wire \Tile_X3Y1_NN4BEG[13] ;
 wire \Tile_X3Y1_NN4BEG[14] ;
 wire \Tile_X3Y1_NN4BEG[15] ;
 wire \Tile_X3Y1_NN4BEG[1] ;
 wire \Tile_X3Y1_NN4BEG[2] ;
 wire \Tile_X3Y1_NN4BEG[3] ;
 wire \Tile_X3Y1_NN4BEG[4] ;
 wire \Tile_X3Y1_NN4BEG[5] ;
 wire \Tile_X3Y1_NN4BEG[6] ;
 wire \Tile_X3Y1_NN4BEG[7] ;
 wire \Tile_X3Y1_NN4BEG[8] ;
 wire \Tile_X3Y1_NN4BEG[9] ;
 wire \Tile_X3Y1_S1BEG[0] ;
 wire \Tile_X3Y1_S1BEG[1] ;
 wire \Tile_X3Y1_S1BEG[2] ;
 wire \Tile_X3Y1_S1BEG[3] ;
 wire \Tile_X3Y1_S2BEG[0] ;
 wire \Tile_X3Y1_S2BEG[1] ;
 wire \Tile_X3Y1_S2BEG[2] ;
 wire \Tile_X3Y1_S2BEG[3] ;
 wire \Tile_X3Y1_S2BEG[4] ;
 wire \Tile_X3Y1_S2BEG[5] ;
 wire \Tile_X3Y1_S2BEG[6] ;
 wire \Tile_X3Y1_S2BEG[7] ;
 wire \Tile_X3Y1_S2BEGb[0] ;
 wire \Tile_X3Y1_S2BEGb[1] ;
 wire \Tile_X3Y1_S2BEGb[2] ;
 wire \Tile_X3Y1_S2BEGb[3] ;
 wire \Tile_X3Y1_S2BEGb[4] ;
 wire \Tile_X3Y1_S2BEGb[5] ;
 wire \Tile_X3Y1_S2BEGb[6] ;
 wire \Tile_X3Y1_S2BEGb[7] ;
 wire \Tile_X3Y1_S4BEG[0] ;
 wire \Tile_X3Y1_S4BEG[10] ;
 wire \Tile_X3Y1_S4BEG[11] ;
 wire \Tile_X3Y1_S4BEG[12] ;
 wire \Tile_X3Y1_S4BEG[13] ;
 wire \Tile_X3Y1_S4BEG[14] ;
 wire \Tile_X3Y1_S4BEG[15] ;
 wire \Tile_X3Y1_S4BEG[1] ;
 wire \Tile_X3Y1_S4BEG[2] ;
 wire \Tile_X3Y1_S4BEG[3] ;
 wire \Tile_X3Y1_S4BEG[4] ;
 wire \Tile_X3Y1_S4BEG[5] ;
 wire \Tile_X3Y1_S4BEG[6] ;
 wire \Tile_X3Y1_S4BEG[7] ;
 wire \Tile_X3Y1_S4BEG[8] ;
 wire \Tile_X3Y1_S4BEG[9] ;
 wire \Tile_X3Y1_SS4BEG[0] ;
 wire \Tile_X3Y1_SS4BEG[10] ;
 wire \Tile_X3Y1_SS4BEG[11] ;
 wire \Tile_X3Y1_SS4BEG[12] ;
 wire \Tile_X3Y1_SS4BEG[13] ;
 wire \Tile_X3Y1_SS4BEG[14] ;
 wire \Tile_X3Y1_SS4BEG[15] ;
 wire \Tile_X3Y1_SS4BEG[1] ;
 wire \Tile_X3Y1_SS4BEG[2] ;
 wire \Tile_X3Y1_SS4BEG[3] ;
 wire \Tile_X3Y1_SS4BEG[4] ;
 wire \Tile_X3Y1_SS4BEG[5] ;
 wire \Tile_X3Y1_SS4BEG[6] ;
 wire \Tile_X3Y1_SS4BEG[7] ;
 wire \Tile_X3Y1_SS4BEG[8] ;
 wire \Tile_X3Y1_SS4BEG[9] ;
 wire Tile_X3Y1_UserCLKo;
 wire \Tile_X3Y1_W1BEG[0] ;
 wire \Tile_X3Y1_W1BEG[1] ;
 wire \Tile_X3Y1_W1BEG[2] ;
 wire \Tile_X3Y1_W1BEG[3] ;
 wire \Tile_X3Y1_W2BEG[0] ;
 wire \Tile_X3Y1_W2BEG[1] ;
 wire \Tile_X3Y1_W2BEG[2] ;
 wire \Tile_X3Y1_W2BEG[3] ;
 wire \Tile_X3Y1_W2BEG[4] ;
 wire \Tile_X3Y1_W2BEG[5] ;
 wire \Tile_X3Y1_W2BEG[6] ;
 wire \Tile_X3Y1_W2BEG[7] ;
 wire \Tile_X3Y1_W2BEGb[0] ;
 wire \Tile_X3Y1_W2BEGb[1] ;
 wire \Tile_X3Y1_W2BEGb[2] ;
 wire \Tile_X3Y1_W2BEGb[3] ;
 wire \Tile_X3Y1_W2BEGb[4] ;
 wire \Tile_X3Y1_W2BEGb[5] ;
 wire \Tile_X3Y1_W2BEGb[6] ;
 wire \Tile_X3Y1_W2BEGb[7] ;
 wire \Tile_X3Y1_W6BEG[0] ;
 wire \Tile_X3Y1_W6BEG[10] ;
 wire \Tile_X3Y1_W6BEG[11] ;
 wire \Tile_X3Y1_W6BEG[1] ;
 wire \Tile_X3Y1_W6BEG[2] ;
 wire \Tile_X3Y1_W6BEG[3] ;
 wire \Tile_X3Y1_W6BEG[4] ;
 wire \Tile_X3Y1_W6BEG[5] ;
 wire \Tile_X3Y1_W6BEG[6] ;
 wire \Tile_X3Y1_W6BEG[7] ;
 wire \Tile_X3Y1_W6BEG[8] ;
 wire \Tile_X3Y1_W6BEG[9] ;
 wire \Tile_X3Y1_WW4BEG[0] ;
 wire \Tile_X3Y1_WW4BEG[10] ;
 wire \Tile_X3Y1_WW4BEG[11] ;
 wire \Tile_X3Y1_WW4BEG[12] ;
 wire \Tile_X3Y1_WW4BEG[13] ;
 wire \Tile_X3Y1_WW4BEG[14] ;
 wire \Tile_X3Y1_WW4BEG[15] ;
 wire \Tile_X3Y1_WW4BEG[1] ;
 wire \Tile_X3Y1_WW4BEG[2] ;
 wire \Tile_X3Y1_WW4BEG[3] ;
 wire \Tile_X3Y1_WW4BEG[4] ;
 wire \Tile_X3Y1_WW4BEG[5] ;
 wire \Tile_X3Y1_WW4BEG[6] ;
 wire \Tile_X3Y1_WW4BEG[7] ;
 wire \Tile_X3Y1_WW4BEG[8] ;
 wire \Tile_X3Y1_WW4BEG[9] ;
 wire Tile_X3Y2_Co;
 wire \Tile_X3Y2_E1BEG[0] ;
 wire \Tile_X3Y2_E1BEG[1] ;
 wire \Tile_X3Y2_E1BEG[2] ;
 wire \Tile_X3Y2_E1BEG[3] ;
 wire \Tile_X3Y2_E2BEG[0] ;
 wire \Tile_X3Y2_E2BEG[1] ;
 wire \Tile_X3Y2_E2BEG[2] ;
 wire \Tile_X3Y2_E2BEG[3] ;
 wire \Tile_X3Y2_E2BEG[4] ;
 wire \Tile_X3Y2_E2BEG[5] ;
 wire \Tile_X3Y2_E2BEG[6] ;
 wire \Tile_X3Y2_E2BEG[7] ;
 wire \Tile_X3Y2_E2BEGb[0] ;
 wire \Tile_X3Y2_E2BEGb[1] ;
 wire \Tile_X3Y2_E2BEGb[2] ;
 wire \Tile_X3Y2_E2BEGb[3] ;
 wire \Tile_X3Y2_E2BEGb[4] ;
 wire \Tile_X3Y2_E2BEGb[5] ;
 wire \Tile_X3Y2_E2BEGb[6] ;
 wire \Tile_X3Y2_E2BEGb[7] ;
 wire \Tile_X3Y2_E6BEG[0] ;
 wire \Tile_X3Y2_E6BEG[10] ;
 wire \Tile_X3Y2_E6BEG[11] ;
 wire \Tile_X3Y2_E6BEG[1] ;
 wire \Tile_X3Y2_E6BEG[2] ;
 wire \Tile_X3Y2_E6BEG[3] ;
 wire \Tile_X3Y2_E6BEG[4] ;
 wire \Tile_X3Y2_E6BEG[5] ;
 wire \Tile_X3Y2_E6BEG[6] ;
 wire \Tile_X3Y2_E6BEG[7] ;
 wire \Tile_X3Y2_E6BEG[8] ;
 wire \Tile_X3Y2_E6BEG[9] ;
 wire \Tile_X3Y2_EE4BEG[0] ;
 wire \Tile_X3Y2_EE4BEG[10] ;
 wire \Tile_X3Y2_EE4BEG[11] ;
 wire \Tile_X3Y2_EE4BEG[12] ;
 wire \Tile_X3Y2_EE4BEG[13] ;
 wire \Tile_X3Y2_EE4BEG[14] ;
 wire \Tile_X3Y2_EE4BEG[15] ;
 wire \Tile_X3Y2_EE4BEG[1] ;
 wire \Tile_X3Y2_EE4BEG[2] ;
 wire \Tile_X3Y2_EE4BEG[3] ;
 wire \Tile_X3Y2_EE4BEG[4] ;
 wire \Tile_X3Y2_EE4BEG[5] ;
 wire \Tile_X3Y2_EE4BEG[6] ;
 wire \Tile_X3Y2_EE4BEG[7] ;
 wire \Tile_X3Y2_EE4BEG[8] ;
 wire \Tile_X3Y2_EE4BEG[9] ;
 wire \Tile_X3Y2_FrameData_O[0] ;
 wire \Tile_X3Y2_FrameData_O[10] ;
 wire \Tile_X3Y2_FrameData_O[11] ;
 wire \Tile_X3Y2_FrameData_O[12] ;
 wire \Tile_X3Y2_FrameData_O[13] ;
 wire \Tile_X3Y2_FrameData_O[14] ;
 wire \Tile_X3Y2_FrameData_O[15] ;
 wire \Tile_X3Y2_FrameData_O[16] ;
 wire \Tile_X3Y2_FrameData_O[17] ;
 wire \Tile_X3Y2_FrameData_O[18] ;
 wire \Tile_X3Y2_FrameData_O[19] ;
 wire \Tile_X3Y2_FrameData_O[1] ;
 wire \Tile_X3Y2_FrameData_O[20] ;
 wire \Tile_X3Y2_FrameData_O[21] ;
 wire \Tile_X3Y2_FrameData_O[22] ;
 wire \Tile_X3Y2_FrameData_O[23] ;
 wire \Tile_X3Y2_FrameData_O[24] ;
 wire \Tile_X3Y2_FrameData_O[25] ;
 wire \Tile_X3Y2_FrameData_O[26] ;
 wire \Tile_X3Y2_FrameData_O[27] ;
 wire \Tile_X3Y2_FrameData_O[28] ;
 wire \Tile_X3Y2_FrameData_O[29] ;
 wire \Tile_X3Y2_FrameData_O[2] ;
 wire \Tile_X3Y2_FrameData_O[30] ;
 wire \Tile_X3Y2_FrameData_O[31] ;
 wire \Tile_X3Y2_FrameData_O[3] ;
 wire \Tile_X3Y2_FrameData_O[4] ;
 wire \Tile_X3Y2_FrameData_O[5] ;
 wire \Tile_X3Y2_FrameData_O[6] ;
 wire \Tile_X3Y2_FrameData_O[7] ;
 wire \Tile_X3Y2_FrameData_O[8] ;
 wire \Tile_X3Y2_FrameData_O[9] ;
 wire \Tile_X3Y2_FrameStrobe_O[0] ;
 wire \Tile_X3Y2_FrameStrobe_O[10] ;
 wire \Tile_X3Y2_FrameStrobe_O[11] ;
 wire \Tile_X3Y2_FrameStrobe_O[12] ;
 wire \Tile_X3Y2_FrameStrobe_O[13] ;
 wire \Tile_X3Y2_FrameStrobe_O[14] ;
 wire \Tile_X3Y2_FrameStrobe_O[15] ;
 wire \Tile_X3Y2_FrameStrobe_O[16] ;
 wire \Tile_X3Y2_FrameStrobe_O[17] ;
 wire \Tile_X3Y2_FrameStrobe_O[18] ;
 wire \Tile_X3Y2_FrameStrobe_O[19] ;
 wire \Tile_X3Y2_FrameStrobe_O[1] ;
 wire \Tile_X3Y2_FrameStrobe_O[2] ;
 wire \Tile_X3Y2_FrameStrobe_O[3] ;
 wire \Tile_X3Y2_FrameStrobe_O[4] ;
 wire \Tile_X3Y2_FrameStrobe_O[5] ;
 wire \Tile_X3Y2_FrameStrobe_O[6] ;
 wire \Tile_X3Y2_FrameStrobe_O[7] ;
 wire \Tile_X3Y2_FrameStrobe_O[8] ;
 wire \Tile_X3Y2_FrameStrobe_O[9] ;
 wire \Tile_X3Y2_N1BEG[0] ;
 wire \Tile_X3Y2_N1BEG[1] ;
 wire \Tile_X3Y2_N1BEG[2] ;
 wire \Tile_X3Y2_N1BEG[3] ;
 wire \Tile_X3Y2_N2BEG[0] ;
 wire \Tile_X3Y2_N2BEG[1] ;
 wire \Tile_X3Y2_N2BEG[2] ;
 wire \Tile_X3Y2_N2BEG[3] ;
 wire \Tile_X3Y2_N2BEG[4] ;
 wire \Tile_X3Y2_N2BEG[5] ;
 wire \Tile_X3Y2_N2BEG[6] ;
 wire \Tile_X3Y2_N2BEG[7] ;
 wire \Tile_X3Y2_N2BEGb[0] ;
 wire \Tile_X3Y2_N2BEGb[1] ;
 wire \Tile_X3Y2_N2BEGb[2] ;
 wire \Tile_X3Y2_N2BEGb[3] ;
 wire \Tile_X3Y2_N2BEGb[4] ;
 wire \Tile_X3Y2_N2BEGb[5] ;
 wire \Tile_X3Y2_N2BEGb[6] ;
 wire \Tile_X3Y2_N2BEGb[7] ;
 wire \Tile_X3Y2_N4BEG[0] ;
 wire \Tile_X3Y2_N4BEG[10] ;
 wire \Tile_X3Y2_N4BEG[11] ;
 wire \Tile_X3Y2_N4BEG[12] ;
 wire \Tile_X3Y2_N4BEG[13] ;
 wire \Tile_X3Y2_N4BEG[14] ;
 wire \Tile_X3Y2_N4BEG[15] ;
 wire \Tile_X3Y2_N4BEG[1] ;
 wire \Tile_X3Y2_N4BEG[2] ;
 wire \Tile_X3Y2_N4BEG[3] ;
 wire \Tile_X3Y2_N4BEG[4] ;
 wire \Tile_X3Y2_N4BEG[5] ;
 wire \Tile_X3Y2_N4BEG[6] ;
 wire \Tile_X3Y2_N4BEG[7] ;
 wire \Tile_X3Y2_N4BEG[8] ;
 wire \Tile_X3Y2_N4BEG[9] ;
 wire \Tile_X3Y2_NN4BEG[0] ;
 wire \Tile_X3Y2_NN4BEG[10] ;
 wire \Tile_X3Y2_NN4BEG[11] ;
 wire \Tile_X3Y2_NN4BEG[12] ;
 wire \Tile_X3Y2_NN4BEG[13] ;
 wire \Tile_X3Y2_NN4BEG[14] ;
 wire \Tile_X3Y2_NN4BEG[15] ;
 wire \Tile_X3Y2_NN4BEG[1] ;
 wire \Tile_X3Y2_NN4BEG[2] ;
 wire \Tile_X3Y2_NN4BEG[3] ;
 wire \Tile_X3Y2_NN4BEG[4] ;
 wire \Tile_X3Y2_NN4BEG[5] ;
 wire \Tile_X3Y2_NN4BEG[6] ;
 wire \Tile_X3Y2_NN4BEG[7] ;
 wire \Tile_X3Y2_NN4BEG[8] ;
 wire \Tile_X3Y2_NN4BEG[9] ;
 wire \Tile_X3Y2_S1BEG[0] ;
 wire \Tile_X3Y2_S1BEG[1] ;
 wire \Tile_X3Y2_S1BEG[2] ;
 wire \Tile_X3Y2_S1BEG[3] ;
 wire \Tile_X3Y2_S2BEG[0] ;
 wire \Tile_X3Y2_S2BEG[1] ;
 wire \Tile_X3Y2_S2BEG[2] ;
 wire \Tile_X3Y2_S2BEG[3] ;
 wire \Tile_X3Y2_S2BEG[4] ;
 wire \Tile_X3Y2_S2BEG[5] ;
 wire \Tile_X3Y2_S2BEG[6] ;
 wire \Tile_X3Y2_S2BEG[7] ;
 wire \Tile_X3Y2_S2BEGb[0] ;
 wire \Tile_X3Y2_S2BEGb[1] ;
 wire \Tile_X3Y2_S2BEGb[2] ;
 wire \Tile_X3Y2_S2BEGb[3] ;
 wire \Tile_X3Y2_S2BEGb[4] ;
 wire \Tile_X3Y2_S2BEGb[5] ;
 wire \Tile_X3Y2_S2BEGb[6] ;
 wire \Tile_X3Y2_S2BEGb[7] ;
 wire \Tile_X3Y2_S4BEG[0] ;
 wire \Tile_X3Y2_S4BEG[10] ;
 wire \Tile_X3Y2_S4BEG[11] ;
 wire \Tile_X3Y2_S4BEG[12] ;
 wire \Tile_X3Y2_S4BEG[13] ;
 wire \Tile_X3Y2_S4BEG[14] ;
 wire \Tile_X3Y2_S4BEG[15] ;
 wire \Tile_X3Y2_S4BEG[1] ;
 wire \Tile_X3Y2_S4BEG[2] ;
 wire \Tile_X3Y2_S4BEG[3] ;
 wire \Tile_X3Y2_S4BEG[4] ;
 wire \Tile_X3Y2_S4BEG[5] ;
 wire \Tile_X3Y2_S4BEG[6] ;
 wire \Tile_X3Y2_S4BEG[7] ;
 wire \Tile_X3Y2_S4BEG[8] ;
 wire \Tile_X3Y2_S4BEG[9] ;
 wire \Tile_X3Y2_SS4BEG[0] ;
 wire \Tile_X3Y2_SS4BEG[10] ;
 wire \Tile_X3Y2_SS4BEG[11] ;
 wire \Tile_X3Y2_SS4BEG[12] ;
 wire \Tile_X3Y2_SS4BEG[13] ;
 wire \Tile_X3Y2_SS4BEG[14] ;
 wire \Tile_X3Y2_SS4BEG[15] ;
 wire \Tile_X3Y2_SS4BEG[1] ;
 wire \Tile_X3Y2_SS4BEG[2] ;
 wire \Tile_X3Y2_SS4BEG[3] ;
 wire \Tile_X3Y2_SS4BEG[4] ;
 wire \Tile_X3Y2_SS4BEG[5] ;
 wire \Tile_X3Y2_SS4BEG[6] ;
 wire \Tile_X3Y2_SS4BEG[7] ;
 wire \Tile_X3Y2_SS4BEG[8] ;
 wire \Tile_X3Y2_SS4BEG[9] ;
 wire Tile_X3Y2_UserCLKo;
 wire \Tile_X3Y2_W1BEG[0] ;
 wire \Tile_X3Y2_W1BEG[1] ;
 wire \Tile_X3Y2_W1BEG[2] ;
 wire \Tile_X3Y2_W1BEG[3] ;
 wire \Tile_X3Y2_W2BEG[0] ;
 wire \Tile_X3Y2_W2BEG[1] ;
 wire \Tile_X3Y2_W2BEG[2] ;
 wire \Tile_X3Y2_W2BEG[3] ;
 wire \Tile_X3Y2_W2BEG[4] ;
 wire \Tile_X3Y2_W2BEG[5] ;
 wire \Tile_X3Y2_W2BEG[6] ;
 wire \Tile_X3Y2_W2BEG[7] ;
 wire \Tile_X3Y2_W2BEGb[0] ;
 wire \Tile_X3Y2_W2BEGb[1] ;
 wire \Tile_X3Y2_W2BEGb[2] ;
 wire \Tile_X3Y2_W2BEGb[3] ;
 wire \Tile_X3Y2_W2BEGb[4] ;
 wire \Tile_X3Y2_W2BEGb[5] ;
 wire \Tile_X3Y2_W2BEGb[6] ;
 wire \Tile_X3Y2_W2BEGb[7] ;
 wire \Tile_X3Y2_W6BEG[0] ;
 wire \Tile_X3Y2_W6BEG[10] ;
 wire \Tile_X3Y2_W6BEG[11] ;
 wire \Tile_X3Y2_W6BEG[1] ;
 wire \Tile_X3Y2_W6BEG[2] ;
 wire \Tile_X3Y2_W6BEG[3] ;
 wire \Tile_X3Y2_W6BEG[4] ;
 wire \Tile_X3Y2_W6BEG[5] ;
 wire \Tile_X3Y2_W6BEG[6] ;
 wire \Tile_X3Y2_W6BEG[7] ;
 wire \Tile_X3Y2_W6BEG[8] ;
 wire \Tile_X3Y2_W6BEG[9] ;
 wire \Tile_X3Y2_WW4BEG[0] ;
 wire \Tile_X3Y2_WW4BEG[10] ;
 wire \Tile_X3Y2_WW4BEG[11] ;
 wire \Tile_X3Y2_WW4BEG[12] ;
 wire \Tile_X3Y2_WW4BEG[13] ;
 wire \Tile_X3Y2_WW4BEG[14] ;
 wire \Tile_X3Y2_WW4BEG[15] ;
 wire \Tile_X3Y2_WW4BEG[1] ;
 wire \Tile_X3Y2_WW4BEG[2] ;
 wire \Tile_X3Y2_WW4BEG[3] ;
 wire \Tile_X3Y2_WW4BEG[4] ;
 wire \Tile_X3Y2_WW4BEG[5] ;
 wire \Tile_X3Y2_WW4BEG[6] ;
 wire \Tile_X3Y2_WW4BEG[7] ;
 wire \Tile_X3Y2_WW4BEG[8] ;
 wire \Tile_X3Y2_WW4BEG[9] ;
 wire Tile_X3Y3_Co;
 wire \Tile_X3Y3_E1BEG[0] ;
 wire \Tile_X3Y3_E1BEG[1] ;
 wire \Tile_X3Y3_E1BEG[2] ;
 wire \Tile_X3Y3_E1BEG[3] ;
 wire \Tile_X3Y3_E2BEG[0] ;
 wire \Tile_X3Y3_E2BEG[1] ;
 wire \Tile_X3Y3_E2BEG[2] ;
 wire \Tile_X3Y3_E2BEG[3] ;
 wire \Tile_X3Y3_E2BEG[4] ;
 wire \Tile_X3Y3_E2BEG[5] ;
 wire \Tile_X3Y3_E2BEG[6] ;
 wire \Tile_X3Y3_E2BEG[7] ;
 wire \Tile_X3Y3_E2BEGb[0] ;
 wire \Tile_X3Y3_E2BEGb[1] ;
 wire \Tile_X3Y3_E2BEGb[2] ;
 wire \Tile_X3Y3_E2BEGb[3] ;
 wire \Tile_X3Y3_E2BEGb[4] ;
 wire \Tile_X3Y3_E2BEGb[5] ;
 wire \Tile_X3Y3_E2BEGb[6] ;
 wire \Tile_X3Y3_E2BEGb[7] ;
 wire \Tile_X3Y3_E6BEG[0] ;
 wire \Tile_X3Y3_E6BEG[10] ;
 wire \Tile_X3Y3_E6BEG[11] ;
 wire \Tile_X3Y3_E6BEG[1] ;
 wire \Tile_X3Y3_E6BEG[2] ;
 wire \Tile_X3Y3_E6BEG[3] ;
 wire \Tile_X3Y3_E6BEG[4] ;
 wire \Tile_X3Y3_E6BEG[5] ;
 wire \Tile_X3Y3_E6BEG[6] ;
 wire \Tile_X3Y3_E6BEG[7] ;
 wire \Tile_X3Y3_E6BEG[8] ;
 wire \Tile_X3Y3_E6BEG[9] ;
 wire \Tile_X3Y3_EE4BEG[0] ;
 wire \Tile_X3Y3_EE4BEG[10] ;
 wire \Tile_X3Y3_EE4BEG[11] ;
 wire \Tile_X3Y3_EE4BEG[12] ;
 wire \Tile_X3Y3_EE4BEG[13] ;
 wire \Tile_X3Y3_EE4BEG[14] ;
 wire \Tile_X3Y3_EE4BEG[15] ;
 wire \Tile_X3Y3_EE4BEG[1] ;
 wire \Tile_X3Y3_EE4BEG[2] ;
 wire \Tile_X3Y3_EE4BEG[3] ;
 wire \Tile_X3Y3_EE4BEG[4] ;
 wire \Tile_X3Y3_EE4BEG[5] ;
 wire \Tile_X3Y3_EE4BEG[6] ;
 wire \Tile_X3Y3_EE4BEG[7] ;
 wire \Tile_X3Y3_EE4BEG[8] ;
 wire \Tile_X3Y3_EE4BEG[9] ;
 wire \Tile_X3Y3_FrameData_O[0] ;
 wire \Tile_X3Y3_FrameData_O[10] ;
 wire \Tile_X3Y3_FrameData_O[11] ;
 wire \Tile_X3Y3_FrameData_O[12] ;
 wire \Tile_X3Y3_FrameData_O[13] ;
 wire \Tile_X3Y3_FrameData_O[14] ;
 wire \Tile_X3Y3_FrameData_O[15] ;
 wire \Tile_X3Y3_FrameData_O[16] ;
 wire \Tile_X3Y3_FrameData_O[17] ;
 wire \Tile_X3Y3_FrameData_O[18] ;
 wire \Tile_X3Y3_FrameData_O[19] ;
 wire \Tile_X3Y3_FrameData_O[1] ;
 wire \Tile_X3Y3_FrameData_O[20] ;
 wire \Tile_X3Y3_FrameData_O[21] ;
 wire \Tile_X3Y3_FrameData_O[22] ;
 wire \Tile_X3Y3_FrameData_O[23] ;
 wire \Tile_X3Y3_FrameData_O[24] ;
 wire \Tile_X3Y3_FrameData_O[25] ;
 wire \Tile_X3Y3_FrameData_O[26] ;
 wire \Tile_X3Y3_FrameData_O[27] ;
 wire \Tile_X3Y3_FrameData_O[28] ;
 wire \Tile_X3Y3_FrameData_O[29] ;
 wire \Tile_X3Y3_FrameData_O[2] ;
 wire \Tile_X3Y3_FrameData_O[30] ;
 wire \Tile_X3Y3_FrameData_O[31] ;
 wire \Tile_X3Y3_FrameData_O[3] ;
 wire \Tile_X3Y3_FrameData_O[4] ;
 wire \Tile_X3Y3_FrameData_O[5] ;
 wire \Tile_X3Y3_FrameData_O[6] ;
 wire \Tile_X3Y3_FrameData_O[7] ;
 wire \Tile_X3Y3_FrameData_O[8] ;
 wire \Tile_X3Y3_FrameData_O[9] ;
 wire \Tile_X3Y3_FrameStrobe_O[0] ;
 wire \Tile_X3Y3_FrameStrobe_O[10] ;
 wire \Tile_X3Y3_FrameStrobe_O[11] ;
 wire \Tile_X3Y3_FrameStrobe_O[12] ;
 wire \Tile_X3Y3_FrameStrobe_O[13] ;
 wire \Tile_X3Y3_FrameStrobe_O[14] ;
 wire \Tile_X3Y3_FrameStrobe_O[15] ;
 wire \Tile_X3Y3_FrameStrobe_O[16] ;
 wire \Tile_X3Y3_FrameStrobe_O[17] ;
 wire \Tile_X3Y3_FrameStrobe_O[18] ;
 wire \Tile_X3Y3_FrameStrobe_O[19] ;
 wire \Tile_X3Y3_FrameStrobe_O[1] ;
 wire \Tile_X3Y3_FrameStrobe_O[2] ;
 wire \Tile_X3Y3_FrameStrobe_O[3] ;
 wire \Tile_X3Y3_FrameStrobe_O[4] ;
 wire \Tile_X3Y3_FrameStrobe_O[5] ;
 wire \Tile_X3Y3_FrameStrobe_O[6] ;
 wire \Tile_X3Y3_FrameStrobe_O[7] ;
 wire \Tile_X3Y3_FrameStrobe_O[8] ;
 wire \Tile_X3Y3_FrameStrobe_O[9] ;
 wire \Tile_X3Y3_N1BEG[0] ;
 wire \Tile_X3Y3_N1BEG[1] ;
 wire \Tile_X3Y3_N1BEG[2] ;
 wire \Tile_X3Y3_N1BEG[3] ;
 wire \Tile_X3Y3_N2BEG[0] ;
 wire \Tile_X3Y3_N2BEG[1] ;
 wire \Tile_X3Y3_N2BEG[2] ;
 wire \Tile_X3Y3_N2BEG[3] ;
 wire \Tile_X3Y3_N2BEG[4] ;
 wire \Tile_X3Y3_N2BEG[5] ;
 wire \Tile_X3Y3_N2BEG[6] ;
 wire \Tile_X3Y3_N2BEG[7] ;
 wire \Tile_X3Y3_N2BEGb[0] ;
 wire \Tile_X3Y3_N2BEGb[1] ;
 wire \Tile_X3Y3_N2BEGb[2] ;
 wire \Tile_X3Y3_N2BEGb[3] ;
 wire \Tile_X3Y3_N2BEGb[4] ;
 wire \Tile_X3Y3_N2BEGb[5] ;
 wire \Tile_X3Y3_N2BEGb[6] ;
 wire \Tile_X3Y3_N2BEGb[7] ;
 wire \Tile_X3Y3_N4BEG[0] ;
 wire \Tile_X3Y3_N4BEG[10] ;
 wire \Tile_X3Y3_N4BEG[11] ;
 wire \Tile_X3Y3_N4BEG[12] ;
 wire \Tile_X3Y3_N4BEG[13] ;
 wire \Tile_X3Y3_N4BEG[14] ;
 wire \Tile_X3Y3_N4BEG[15] ;
 wire \Tile_X3Y3_N4BEG[1] ;
 wire \Tile_X3Y3_N4BEG[2] ;
 wire \Tile_X3Y3_N4BEG[3] ;
 wire \Tile_X3Y3_N4BEG[4] ;
 wire \Tile_X3Y3_N4BEG[5] ;
 wire \Tile_X3Y3_N4BEG[6] ;
 wire \Tile_X3Y3_N4BEG[7] ;
 wire \Tile_X3Y3_N4BEG[8] ;
 wire \Tile_X3Y3_N4BEG[9] ;
 wire \Tile_X3Y3_NN4BEG[0] ;
 wire \Tile_X3Y3_NN4BEG[10] ;
 wire \Tile_X3Y3_NN4BEG[11] ;
 wire \Tile_X3Y3_NN4BEG[12] ;
 wire \Tile_X3Y3_NN4BEG[13] ;
 wire \Tile_X3Y3_NN4BEG[14] ;
 wire \Tile_X3Y3_NN4BEG[15] ;
 wire \Tile_X3Y3_NN4BEG[1] ;
 wire \Tile_X3Y3_NN4BEG[2] ;
 wire \Tile_X3Y3_NN4BEG[3] ;
 wire \Tile_X3Y3_NN4BEG[4] ;
 wire \Tile_X3Y3_NN4BEG[5] ;
 wire \Tile_X3Y3_NN4BEG[6] ;
 wire \Tile_X3Y3_NN4BEG[7] ;
 wire \Tile_X3Y3_NN4BEG[8] ;
 wire \Tile_X3Y3_NN4BEG[9] ;
 wire \Tile_X3Y3_S1BEG[0] ;
 wire \Tile_X3Y3_S1BEG[1] ;
 wire \Tile_X3Y3_S1BEG[2] ;
 wire \Tile_X3Y3_S1BEG[3] ;
 wire \Tile_X3Y3_S2BEG[0] ;
 wire \Tile_X3Y3_S2BEG[1] ;
 wire \Tile_X3Y3_S2BEG[2] ;
 wire \Tile_X3Y3_S2BEG[3] ;
 wire \Tile_X3Y3_S2BEG[4] ;
 wire \Tile_X3Y3_S2BEG[5] ;
 wire \Tile_X3Y3_S2BEG[6] ;
 wire \Tile_X3Y3_S2BEG[7] ;
 wire \Tile_X3Y3_S2BEGb[0] ;
 wire \Tile_X3Y3_S2BEGb[1] ;
 wire \Tile_X3Y3_S2BEGb[2] ;
 wire \Tile_X3Y3_S2BEGb[3] ;
 wire \Tile_X3Y3_S2BEGb[4] ;
 wire \Tile_X3Y3_S2BEGb[5] ;
 wire \Tile_X3Y3_S2BEGb[6] ;
 wire \Tile_X3Y3_S2BEGb[7] ;
 wire \Tile_X3Y3_S4BEG[0] ;
 wire \Tile_X3Y3_S4BEG[10] ;
 wire \Tile_X3Y3_S4BEG[11] ;
 wire \Tile_X3Y3_S4BEG[12] ;
 wire \Tile_X3Y3_S4BEG[13] ;
 wire \Tile_X3Y3_S4BEG[14] ;
 wire \Tile_X3Y3_S4BEG[15] ;
 wire \Tile_X3Y3_S4BEG[1] ;
 wire \Tile_X3Y3_S4BEG[2] ;
 wire \Tile_X3Y3_S4BEG[3] ;
 wire \Tile_X3Y3_S4BEG[4] ;
 wire \Tile_X3Y3_S4BEG[5] ;
 wire \Tile_X3Y3_S4BEG[6] ;
 wire \Tile_X3Y3_S4BEG[7] ;
 wire \Tile_X3Y3_S4BEG[8] ;
 wire \Tile_X3Y3_S4BEG[9] ;
 wire \Tile_X3Y3_SS4BEG[0] ;
 wire \Tile_X3Y3_SS4BEG[10] ;
 wire \Tile_X3Y3_SS4BEG[11] ;
 wire \Tile_X3Y3_SS4BEG[12] ;
 wire \Tile_X3Y3_SS4BEG[13] ;
 wire \Tile_X3Y3_SS4BEG[14] ;
 wire \Tile_X3Y3_SS4BEG[15] ;
 wire \Tile_X3Y3_SS4BEG[1] ;
 wire \Tile_X3Y3_SS4BEG[2] ;
 wire \Tile_X3Y3_SS4BEG[3] ;
 wire \Tile_X3Y3_SS4BEG[4] ;
 wire \Tile_X3Y3_SS4BEG[5] ;
 wire \Tile_X3Y3_SS4BEG[6] ;
 wire \Tile_X3Y3_SS4BEG[7] ;
 wire \Tile_X3Y3_SS4BEG[8] ;
 wire \Tile_X3Y3_SS4BEG[9] ;
 wire Tile_X3Y3_UserCLKo;
 wire \Tile_X3Y3_W1BEG[0] ;
 wire \Tile_X3Y3_W1BEG[1] ;
 wire \Tile_X3Y3_W1BEG[2] ;
 wire \Tile_X3Y3_W1BEG[3] ;
 wire \Tile_X3Y3_W2BEG[0] ;
 wire \Tile_X3Y3_W2BEG[1] ;
 wire \Tile_X3Y3_W2BEG[2] ;
 wire \Tile_X3Y3_W2BEG[3] ;
 wire \Tile_X3Y3_W2BEG[4] ;
 wire \Tile_X3Y3_W2BEG[5] ;
 wire \Tile_X3Y3_W2BEG[6] ;
 wire \Tile_X3Y3_W2BEG[7] ;
 wire \Tile_X3Y3_W2BEGb[0] ;
 wire \Tile_X3Y3_W2BEGb[1] ;
 wire \Tile_X3Y3_W2BEGb[2] ;
 wire \Tile_X3Y3_W2BEGb[3] ;
 wire \Tile_X3Y3_W2BEGb[4] ;
 wire \Tile_X3Y3_W2BEGb[5] ;
 wire \Tile_X3Y3_W2BEGb[6] ;
 wire \Tile_X3Y3_W2BEGb[7] ;
 wire \Tile_X3Y3_W6BEG[0] ;
 wire \Tile_X3Y3_W6BEG[10] ;
 wire \Tile_X3Y3_W6BEG[11] ;
 wire \Tile_X3Y3_W6BEG[1] ;
 wire \Tile_X3Y3_W6BEG[2] ;
 wire \Tile_X3Y3_W6BEG[3] ;
 wire \Tile_X3Y3_W6BEG[4] ;
 wire \Tile_X3Y3_W6BEG[5] ;
 wire \Tile_X3Y3_W6BEG[6] ;
 wire \Tile_X3Y3_W6BEG[7] ;
 wire \Tile_X3Y3_W6BEG[8] ;
 wire \Tile_X3Y3_W6BEG[9] ;
 wire \Tile_X3Y3_WW4BEG[0] ;
 wire \Tile_X3Y3_WW4BEG[10] ;
 wire \Tile_X3Y3_WW4BEG[11] ;
 wire \Tile_X3Y3_WW4BEG[12] ;
 wire \Tile_X3Y3_WW4BEG[13] ;
 wire \Tile_X3Y3_WW4BEG[14] ;
 wire \Tile_X3Y3_WW4BEG[15] ;
 wire \Tile_X3Y3_WW4BEG[1] ;
 wire \Tile_X3Y3_WW4BEG[2] ;
 wire \Tile_X3Y3_WW4BEG[3] ;
 wire \Tile_X3Y3_WW4BEG[4] ;
 wire \Tile_X3Y3_WW4BEG[5] ;
 wire \Tile_X3Y3_WW4BEG[6] ;
 wire \Tile_X3Y3_WW4BEG[7] ;
 wire \Tile_X3Y3_WW4BEG[8] ;
 wire \Tile_X3Y3_WW4BEG[9] ;
 wire Tile_X3Y4_Co;
 wire \Tile_X3Y4_E1BEG[0] ;
 wire \Tile_X3Y4_E1BEG[1] ;
 wire \Tile_X3Y4_E1BEG[2] ;
 wire \Tile_X3Y4_E1BEG[3] ;
 wire \Tile_X3Y4_E2BEG[0] ;
 wire \Tile_X3Y4_E2BEG[1] ;
 wire \Tile_X3Y4_E2BEG[2] ;
 wire \Tile_X3Y4_E2BEG[3] ;
 wire \Tile_X3Y4_E2BEG[4] ;
 wire \Tile_X3Y4_E2BEG[5] ;
 wire \Tile_X3Y4_E2BEG[6] ;
 wire \Tile_X3Y4_E2BEG[7] ;
 wire \Tile_X3Y4_E2BEGb[0] ;
 wire \Tile_X3Y4_E2BEGb[1] ;
 wire \Tile_X3Y4_E2BEGb[2] ;
 wire \Tile_X3Y4_E2BEGb[3] ;
 wire \Tile_X3Y4_E2BEGb[4] ;
 wire \Tile_X3Y4_E2BEGb[5] ;
 wire \Tile_X3Y4_E2BEGb[6] ;
 wire \Tile_X3Y4_E2BEGb[7] ;
 wire \Tile_X3Y4_E6BEG[0] ;
 wire \Tile_X3Y4_E6BEG[10] ;
 wire \Tile_X3Y4_E6BEG[11] ;
 wire \Tile_X3Y4_E6BEG[1] ;
 wire \Tile_X3Y4_E6BEG[2] ;
 wire \Tile_X3Y4_E6BEG[3] ;
 wire \Tile_X3Y4_E6BEG[4] ;
 wire \Tile_X3Y4_E6BEG[5] ;
 wire \Tile_X3Y4_E6BEG[6] ;
 wire \Tile_X3Y4_E6BEG[7] ;
 wire \Tile_X3Y4_E6BEG[8] ;
 wire \Tile_X3Y4_E6BEG[9] ;
 wire \Tile_X3Y4_EE4BEG[0] ;
 wire \Tile_X3Y4_EE4BEG[10] ;
 wire \Tile_X3Y4_EE4BEG[11] ;
 wire \Tile_X3Y4_EE4BEG[12] ;
 wire \Tile_X3Y4_EE4BEG[13] ;
 wire \Tile_X3Y4_EE4BEG[14] ;
 wire \Tile_X3Y4_EE4BEG[15] ;
 wire \Tile_X3Y4_EE4BEG[1] ;
 wire \Tile_X3Y4_EE4BEG[2] ;
 wire \Tile_X3Y4_EE4BEG[3] ;
 wire \Tile_X3Y4_EE4BEG[4] ;
 wire \Tile_X3Y4_EE4BEG[5] ;
 wire \Tile_X3Y4_EE4BEG[6] ;
 wire \Tile_X3Y4_EE4BEG[7] ;
 wire \Tile_X3Y4_EE4BEG[8] ;
 wire \Tile_X3Y4_EE4BEG[9] ;
 wire \Tile_X3Y4_FrameData_O[0] ;
 wire \Tile_X3Y4_FrameData_O[10] ;
 wire \Tile_X3Y4_FrameData_O[11] ;
 wire \Tile_X3Y4_FrameData_O[12] ;
 wire \Tile_X3Y4_FrameData_O[13] ;
 wire \Tile_X3Y4_FrameData_O[14] ;
 wire \Tile_X3Y4_FrameData_O[15] ;
 wire \Tile_X3Y4_FrameData_O[16] ;
 wire \Tile_X3Y4_FrameData_O[17] ;
 wire \Tile_X3Y4_FrameData_O[18] ;
 wire \Tile_X3Y4_FrameData_O[19] ;
 wire \Tile_X3Y4_FrameData_O[1] ;
 wire \Tile_X3Y4_FrameData_O[20] ;
 wire \Tile_X3Y4_FrameData_O[21] ;
 wire \Tile_X3Y4_FrameData_O[22] ;
 wire \Tile_X3Y4_FrameData_O[23] ;
 wire \Tile_X3Y4_FrameData_O[24] ;
 wire \Tile_X3Y4_FrameData_O[25] ;
 wire \Tile_X3Y4_FrameData_O[26] ;
 wire \Tile_X3Y4_FrameData_O[27] ;
 wire \Tile_X3Y4_FrameData_O[28] ;
 wire \Tile_X3Y4_FrameData_O[29] ;
 wire \Tile_X3Y4_FrameData_O[2] ;
 wire \Tile_X3Y4_FrameData_O[30] ;
 wire \Tile_X3Y4_FrameData_O[31] ;
 wire \Tile_X3Y4_FrameData_O[3] ;
 wire \Tile_X3Y4_FrameData_O[4] ;
 wire \Tile_X3Y4_FrameData_O[5] ;
 wire \Tile_X3Y4_FrameData_O[6] ;
 wire \Tile_X3Y4_FrameData_O[7] ;
 wire \Tile_X3Y4_FrameData_O[8] ;
 wire \Tile_X3Y4_FrameData_O[9] ;
 wire \Tile_X3Y4_FrameStrobe_O[0] ;
 wire \Tile_X3Y4_FrameStrobe_O[10] ;
 wire \Tile_X3Y4_FrameStrobe_O[11] ;
 wire \Tile_X3Y4_FrameStrobe_O[12] ;
 wire \Tile_X3Y4_FrameStrobe_O[13] ;
 wire \Tile_X3Y4_FrameStrobe_O[14] ;
 wire \Tile_X3Y4_FrameStrobe_O[15] ;
 wire \Tile_X3Y4_FrameStrobe_O[16] ;
 wire \Tile_X3Y4_FrameStrobe_O[17] ;
 wire \Tile_X3Y4_FrameStrobe_O[18] ;
 wire \Tile_X3Y4_FrameStrobe_O[19] ;
 wire \Tile_X3Y4_FrameStrobe_O[1] ;
 wire \Tile_X3Y4_FrameStrobe_O[2] ;
 wire \Tile_X3Y4_FrameStrobe_O[3] ;
 wire \Tile_X3Y4_FrameStrobe_O[4] ;
 wire \Tile_X3Y4_FrameStrobe_O[5] ;
 wire \Tile_X3Y4_FrameStrobe_O[6] ;
 wire \Tile_X3Y4_FrameStrobe_O[7] ;
 wire \Tile_X3Y4_FrameStrobe_O[8] ;
 wire \Tile_X3Y4_FrameStrobe_O[9] ;
 wire \Tile_X3Y4_N1BEG[0] ;
 wire \Tile_X3Y4_N1BEG[1] ;
 wire \Tile_X3Y4_N1BEG[2] ;
 wire \Tile_X3Y4_N1BEG[3] ;
 wire \Tile_X3Y4_N2BEG[0] ;
 wire \Tile_X3Y4_N2BEG[1] ;
 wire \Tile_X3Y4_N2BEG[2] ;
 wire \Tile_X3Y4_N2BEG[3] ;
 wire \Tile_X3Y4_N2BEG[4] ;
 wire \Tile_X3Y4_N2BEG[5] ;
 wire \Tile_X3Y4_N2BEG[6] ;
 wire \Tile_X3Y4_N2BEG[7] ;
 wire \Tile_X3Y4_N2BEGb[0] ;
 wire \Tile_X3Y4_N2BEGb[1] ;
 wire \Tile_X3Y4_N2BEGb[2] ;
 wire \Tile_X3Y4_N2BEGb[3] ;
 wire \Tile_X3Y4_N2BEGb[4] ;
 wire \Tile_X3Y4_N2BEGb[5] ;
 wire \Tile_X3Y4_N2BEGb[6] ;
 wire \Tile_X3Y4_N2BEGb[7] ;
 wire \Tile_X3Y4_N4BEG[0] ;
 wire \Tile_X3Y4_N4BEG[10] ;
 wire \Tile_X3Y4_N4BEG[11] ;
 wire \Tile_X3Y4_N4BEG[12] ;
 wire \Tile_X3Y4_N4BEG[13] ;
 wire \Tile_X3Y4_N4BEG[14] ;
 wire \Tile_X3Y4_N4BEG[15] ;
 wire \Tile_X3Y4_N4BEG[1] ;
 wire \Tile_X3Y4_N4BEG[2] ;
 wire \Tile_X3Y4_N4BEG[3] ;
 wire \Tile_X3Y4_N4BEG[4] ;
 wire \Tile_X3Y4_N4BEG[5] ;
 wire \Tile_X3Y4_N4BEG[6] ;
 wire \Tile_X3Y4_N4BEG[7] ;
 wire \Tile_X3Y4_N4BEG[8] ;
 wire \Tile_X3Y4_N4BEG[9] ;
 wire \Tile_X3Y4_NN4BEG[0] ;
 wire \Tile_X3Y4_NN4BEG[10] ;
 wire \Tile_X3Y4_NN4BEG[11] ;
 wire \Tile_X3Y4_NN4BEG[12] ;
 wire \Tile_X3Y4_NN4BEG[13] ;
 wire \Tile_X3Y4_NN4BEG[14] ;
 wire \Tile_X3Y4_NN4BEG[15] ;
 wire \Tile_X3Y4_NN4BEG[1] ;
 wire \Tile_X3Y4_NN4BEG[2] ;
 wire \Tile_X3Y4_NN4BEG[3] ;
 wire \Tile_X3Y4_NN4BEG[4] ;
 wire \Tile_X3Y4_NN4BEG[5] ;
 wire \Tile_X3Y4_NN4BEG[6] ;
 wire \Tile_X3Y4_NN4BEG[7] ;
 wire \Tile_X3Y4_NN4BEG[8] ;
 wire \Tile_X3Y4_NN4BEG[9] ;
 wire \Tile_X3Y4_S1BEG[0] ;
 wire \Tile_X3Y4_S1BEG[1] ;
 wire \Tile_X3Y4_S1BEG[2] ;
 wire \Tile_X3Y4_S1BEG[3] ;
 wire \Tile_X3Y4_S2BEG[0] ;
 wire \Tile_X3Y4_S2BEG[1] ;
 wire \Tile_X3Y4_S2BEG[2] ;
 wire \Tile_X3Y4_S2BEG[3] ;
 wire \Tile_X3Y4_S2BEG[4] ;
 wire \Tile_X3Y4_S2BEG[5] ;
 wire \Tile_X3Y4_S2BEG[6] ;
 wire \Tile_X3Y4_S2BEG[7] ;
 wire \Tile_X3Y4_S2BEGb[0] ;
 wire \Tile_X3Y4_S2BEGb[1] ;
 wire \Tile_X3Y4_S2BEGb[2] ;
 wire \Tile_X3Y4_S2BEGb[3] ;
 wire \Tile_X3Y4_S2BEGb[4] ;
 wire \Tile_X3Y4_S2BEGb[5] ;
 wire \Tile_X3Y4_S2BEGb[6] ;
 wire \Tile_X3Y4_S2BEGb[7] ;
 wire \Tile_X3Y4_S4BEG[0] ;
 wire \Tile_X3Y4_S4BEG[10] ;
 wire \Tile_X3Y4_S4BEG[11] ;
 wire \Tile_X3Y4_S4BEG[12] ;
 wire \Tile_X3Y4_S4BEG[13] ;
 wire \Tile_X3Y4_S4BEG[14] ;
 wire \Tile_X3Y4_S4BEG[15] ;
 wire \Tile_X3Y4_S4BEG[1] ;
 wire \Tile_X3Y4_S4BEG[2] ;
 wire \Tile_X3Y4_S4BEG[3] ;
 wire \Tile_X3Y4_S4BEG[4] ;
 wire \Tile_X3Y4_S4BEG[5] ;
 wire \Tile_X3Y4_S4BEG[6] ;
 wire \Tile_X3Y4_S4BEG[7] ;
 wire \Tile_X3Y4_S4BEG[8] ;
 wire \Tile_X3Y4_S4BEG[9] ;
 wire \Tile_X3Y4_SS4BEG[0] ;
 wire \Tile_X3Y4_SS4BEG[10] ;
 wire \Tile_X3Y4_SS4BEG[11] ;
 wire \Tile_X3Y4_SS4BEG[12] ;
 wire \Tile_X3Y4_SS4BEG[13] ;
 wire \Tile_X3Y4_SS4BEG[14] ;
 wire \Tile_X3Y4_SS4BEG[15] ;
 wire \Tile_X3Y4_SS4BEG[1] ;
 wire \Tile_X3Y4_SS4BEG[2] ;
 wire \Tile_X3Y4_SS4BEG[3] ;
 wire \Tile_X3Y4_SS4BEG[4] ;
 wire \Tile_X3Y4_SS4BEG[5] ;
 wire \Tile_X3Y4_SS4BEG[6] ;
 wire \Tile_X3Y4_SS4BEG[7] ;
 wire \Tile_X3Y4_SS4BEG[8] ;
 wire \Tile_X3Y4_SS4BEG[9] ;
 wire Tile_X3Y4_UserCLKo;
 wire \Tile_X3Y4_W1BEG[0] ;
 wire \Tile_X3Y4_W1BEG[1] ;
 wire \Tile_X3Y4_W1BEG[2] ;
 wire \Tile_X3Y4_W1BEG[3] ;
 wire \Tile_X3Y4_W2BEG[0] ;
 wire \Tile_X3Y4_W2BEG[1] ;
 wire \Tile_X3Y4_W2BEG[2] ;
 wire \Tile_X3Y4_W2BEG[3] ;
 wire \Tile_X3Y4_W2BEG[4] ;
 wire \Tile_X3Y4_W2BEG[5] ;
 wire \Tile_X3Y4_W2BEG[6] ;
 wire \Tile_X3Y4_W2BEG[7] ;
 wire \Tile_X3Y4_W2BEGb[0] ;
 wire \Tile_X3Y4_W2BEGb[1] ;
 wire \Tile_X3Y4_W2BEGb[2] ;
 wire \Tile_X3Y4_W2BEGb[3] ;
 wire \Tile_X3Y4_W2BEGb[4] ;
 wire \Tile_X3Y4_W2BEGb[5] ;
 wire \Tile_X3Y4_W2BEGb[6] ;
 wire \Tile_X3Y4_W2BEGb[7] ;
 wire \Tile_X3Y4_W6BEG[0] ;
 wire \Tile_X3Y4_W6BEG[10] ;
 wire \Tile_X3Y4_W6BEG[11] ;
 wire \Tile_X3Y4_W6BEG[1] ;
 wire \Tile_X3Y4_W6BEG[2] ;
 wire \Tile_X3Y4_W6BEG[3] ;
 wire \Tile_X3Y4_W6BEG[4] ;
 wire \Tile_X3Y4_W6BEG[5] ;
 wire \Tile_X3Y4_W6BEG[6] ;
 wire \Tile_X3Y4_W6BEG[7] ;
 wire \Tile_X3Y4_W6BEG[8] ;
 wire \Tile_X3Y4_W6BEG[9] ;
 wire \Tile_X3Y4_WW4BEG[0] ;
 wire \Tile_X3Y4_WW4BEG[10] ;
 wire \Tile_X3Y4_WW4BEG[11] ;
 wire \Tile_X3Y4_WW4BEG[12] ;
 wire \Tile_X3Y4_WW4BEG[13] ;
 wire \Tile_X3Y4_WW4BEG[14] ;
 wire \Tile_X3Y4_WW4BEG[15] ;
 wire \Tile_X3Y4_WW4BEG[1] ;
 wire \Tile_X3Y4_WW4BEG[2] ;
 wire \Tile_X3Y4_WW4BEG[3] ;
 wire \Tile_X3Y4_WW4BEG[4] ;
 wire \Tile_X3Y4_WW4BEG[5] ;
 wire \Tile_X3Y4_WW4BEG[6] ;
 wire \Tile_X3Y4_WW4BEG[7] ;
 wire \Tile_X3Y4_WW4BEG[8] ;
 wire \Tile_X3Y4_WW4BEG[9] ;
 wire Tile_X3Y5_Co;
 wire \Tile_X3Y5_E1BEG[0] ;
 wire \Tile_X3Y5_E1BEG[1] ;
 wire \Tile_X3Y5_E1BEG[2] ;
 wire \Tile_X3Y5_E1BEG[3] ;
 wire \Tile_X3Y5_E2BEG[0] ;
 wire \Tile_X3Y5_E2BEG[1] ;
 wire \Tile_X3Y5_E2BEG[2] ;
 wire \Tile_X3Y5_E2BEG[3] ;
 wire \Tile_X3Y5_E2BEG[4] ;
 wire \Tile_X3Y5_E2BEG[5] ;
 wire \Tile_X3Y5_E2BEG[6] ;
 wire \Tile_X3Y5_E2BEG[7] ;
 wire \Tile_X3Y5_E2BEGb[0] ;
 wire \Tile_X3Y5_E2BEGb[1] ;
 wire \Tile_X3Y5_E2BEGb[2] ;
 wire \Tile_X3Y5_E2BEGb[3] ;
 wire \Tile_X3Y5_E2BEGb[4] ;
 wire \Tile_X3Y5_E2BEGb[5] ;
 wire \Tile_X3Y5_E2BEGb[6] ;
 wire \Tile_X3Y5_E2BEGb[7] ;
 wire \Tile_X3Y5_E6BEG[0] ;
 wire \Tile_X3Y5_E6BEG[10] ;
 wire \Tile_X3Y5_E6BEG[11] ;
 wire \Tile_X3Y5_E6BEG[1] ;
 wire \Tile_X3Y5_E6BEG[2] ;
 wire \Tile_X3Y5_E6BEG[3] ;
 wire \Tile_X3Y5_E6BEG[4] ;
 wire \Tile_X3Y5_E6BEG[5] ;
 wire \Tile_X3Y5_E6BEG[6] ;
 wire \Tile_X3Y5_E6BEG[7] ;
 wire \Tile_X3Y5_E6BEG[8] ;
 wire \Tile_X3Y5_E6BEG[9] ;
 wire \Tile_X3Y5_EE4BEG[0] ;
 wire \Tile_X3Y5_EE4BEG[10] ;
 wire \Tile_X3Y5_EE4BEG[11] ;
 wire \Tile_X3Y5_EE4BEG[12] ;
 wire \Tile_X3Y5_EE4BEG[13] ;
 wire \Tile_X3Y5_EE4BEG[14] ;
 wire \Tile_X3Y5_EE4BEG[15] ;
 wire \Tile_X3Y5_EE4BEG[1] ;
 wire \Tile_X3Y5_EE4BEG[2] ;
 wire \Tile_X3Y5_EE4BEG[3] ;
 wire \Tile_X3Y5_EE4BEG[4] ;
 wire \Tile_X3Y5_EE4BEG[5] ;
 wire \Tile_X3Y5_EE4BEG[6] ;
 wire \Tile_X3Y5_EE4BEG[7] ;
 wire \Tile_X3Y5_EE4BEG[8] ;
 wire \Tile_X3Y5_EE4BEG[9] ;
 wire \Tile_X3Y5_FrameData_O[0] ;
 wire \Tile_X3Y5_FrameData_O[10] ;
 wire \Tile_X3Y5_FrameData_O[11] ;
 wire \Tile_X3Y5_FrameData_O[12] ;
 wire \Tile_X3Y5_FrameData_O[13] ;
 wire \Tile_X3Y5_FrameData_O[14] ;
 wire \Tile_X3Y5_FrameData_O[15] ;
 wire \Tile_X3Y5_FrameData_O[16] ;
 wire \Tile_X3Y5_FrameData_O[17] ;
 wire \Tile_X3Y5_FrameData_O[18] ;
 wire \Tile_X3Y5_FrameData_O[19] ;
 wire \Tile_X3Y5_FrameData_O[1] ;
 wire \Tile_X3Y5_FrameData_O[20] ;
 wire \Tile_X3Y5_FrameData_O[21] ;
 wire \Tile_X3Y5_FrameData_O[22] ;
 wire \Tile_X3Y5_FrameData_O[23] ;
 wire \Tile_X3Y5_FrameData_O[24] ;
 wire \Tile_X3Y5_FrameData_O[25] ;
 wire \Tile_X3Y5_FrameData_O[26] ;
 wire \Tile_X3Y5_FrameData_O[27] ;
 wire \Tile_X3Y5_FrameData_O[28] ;
 wire \Tile_X3Y5_FrameData_O[29] ;
 wire \Tile_X3Y5_FrameData_O[2] ;
 wire \Tile_X3Y5_FrameData_O[30] ;
 wire \Tile_X3Y5_FrameData_O[31] ;
 wire \Tile_X3Y5_FrameData_O[3] ;
 wire \Tile_X3Y5_FrameData_O[4] ;
 wire \Tile_X3Y5_FrameData_O[5] ;
 wire \Tile_X3Y5_FrameData_O[6] ;
 wire \Tile_X3Y5_FrameData_O[7] ;
 wire \Tile_X3Y5_FrameData_O[8] ;
 wire \Tile_X3Y5_FrameData_O[9] ;
 wire \Tile_X3Y5_FrameStrobe_O[0] ;
 wire \Tile_X3Y5_FrameStrobe_O[10] ;
 wire \Tile_X3Y5_FrameStrobe_O[11] ;
 wire \Tile_X3Y5_FrameStrobe_O[12] ;
 wire \Tile_X3Y5_FrameStrobe_O[13] ;
 wire \Tile_X3Y5_FrameStrobe_O[14] ;
 wire \Tile_X3Y5_FrameStrobe_O[15] ;
 wire \Tile_X3Y5_FrameStrobe_O[16] ;
 wire \Tile_X3Y5_FrameStrobe_O[17] ;
 wire \Tile_X3Y5_FrameStrobe_O[18] ;
 wire \Tile_X3Y5_FrameStrobe_O[19] ;
 wire \Tile_X3Y5_FrameStrobe_O[1] ;
 wire \Tile_X3Y5_FrameStrobe_O[2] ;
 wire \Tile_X3Y5_FrameStrobe_O[3] ;
 wire \Tile_X3Y5_FrameStrobe_O[4] ;
 wire \Tile_X3Y5_FrameStrobe_O[5] ;
 wire \Tile_X3Y5_FrameStrobe_O[6] ;
 wire \Tile_X3Y5_FrameStrobe_O[7] ;
 wire \Tile_X3Y5_FrameStrobe_O[8] ;
 wire \Tile_X3Y5_FrameStrobe_O[9] ;
 wire \Tile_X3Y5_N1BEG[0] ;
 wire \Tile_X3Y5_N1BEG[1] ;
 wire \Tile_X3Y5_N1BEG[2] ;
 wire \Tile_X3Y5_N1BEG[3] ;
 wire \Tile_X3Y5_N2BEG[0] ;
 wire \Tile_X3Y5_N2BEG[1] ;
 wire \Tile_X3Y5_N2BEG[2] ;
 wire \Tile_X3Y5_N2BEG[3] ;
 wire \Tile_X3Y5_N2BEG[4] ;
 wire \Tile_X3Y5_N2BEG[5] ;
 wire \Tile_X3Y5_N2BEG[6] ;
 wire \Tile_X3Y5_N2BEG[7] ;
 wire \Tile_X3Y5_N2BEGb[0] ;
 wire \Tile_X3Y5_N2BEGb[1] ;
 wire \Tile_X3Y5_N2BEGb[2] ;
 wire \Tile_X3Y5_N2BEGb[3] ;
 wire \Tile_X3Y5_N2BEGb[4] ;
 wire \Tile_X3Y5_N2BEGb[5] ;
 wire \Tile_X3Y5_N2BEGb[6] ;
 wire \Tile_X3Y5_N2BEGb[7] ;
 wire \Tile_X3Y5_N4BEG[0] ;
 wire \Tile_X3Y5_N4BEG[10] ;
 wire \Tile_X3Y5_N4BEG[11] ;
 wire \Tile_X3Y5_N4BEG[12] ;
 wire \Tile_X3Y5_N4BEG[13] ;
 wire \Tile_X3Y5_N4BEG[14] ;
 wire \Tile_X3Y5_N4BEG[15] ;
 wire \Tile_X3Y5_N4BEG[1] ;
 wire \Tile_X3Y5_N4BEG[2] ;
 wire \Tile_X3Y5_N4BEG[3] ;
 wire \Tile_X3Y5_N4BEG[4] ;
 wire \Tile_X3Y5_N4BEG[5] ;
 wire \Tile_X3Y5_N4BEG[6] ;
 wire \Tile_X3Y5_N4BEG[7] ;
 wire \Tile_X3Y5_N4BEG[8] ;
 wire \Tile_X3Y5_N4BEG[9] ;
 wire \Tile_X3Y5_NN4BEG[0] ;
 wire \Tile_X3Y5_NN4BEG[10] ;
 wire \Tile_X3Y5_NN4BEG[11] ;
 wire \Tile_X3Y5_NN4BEG[12] ;
 wire \Tile_X3Y5_NN4BEG[13] ;
 wire \Tile_X3Y5_NN4BEG[14] ;
 wire \Tile_X3Y5_NN4BEG[15] ;
 wire \Tile_X3Y5_NN4BEG[1] ;
 wire \Tile_X3Y5_NN4BEG[2] ;
 wire \Tile_X3Y5_NN4BEG[3] ;
 wire \Tile_X3Y5_NN4BEG[4] ;
 wire \Tile_X3Y5_NN4BEG[5] ;
 wire \Tile_X3Y5_NN4BEG[6] ;
 wire \Tile_X3Y5_NN4BEG[7] ;
 wire \Tile_X3Y5_NN4BEG[8] ;
 wire \Tile_X3Y5_NN4BEG[9] ;
 wire \Tile_X3Y5_S1BEG[0] ;
 wire \Tile_X3Y5_S1BEG[1] ;
 wire \Tile_X3Y5_S1BEG[2] ;
 wire \Tile_X3Y5_S1BEG[3] ;
 wire \Tile_X3Y5_S2BEG[0] ;
 wire \Tile_X3Y5_S2BEG[1] ;
 wire \Tile_X3Y5_S2BEG[2] ;
 wire \Tile_X3Y5_S2BEG[3] ;
 wire \Tile_X3Y5_S2BEG[4] ;
 wire \Tile_X3Y5_S2BEG[5] ;
 wire \Tile_X3Y5_S2BEG[6] ;
 wire \Tile_X3Y5_S2BEG[7] ;
 wire \Tile_X3Y5_S2BEGb[0] ;
 wire \Tile_X3Y5_S2BEGb[1] ;
 wire \Tile_X3Y5_S2BEGb[2] ;
 wire \Tile_X3Y5_S2BEGb[3] ;
 wire \Tile_X3Y5_S2BEGb[4] ;
 wire \Tile_X3Y5_S2BEGb[5] ;
 wire \Tile_X3Y5_S2BEGb[6] ;
 wire \Tile_X3Y5_S2BEGb[7] ;
 wire \Tile_X3Y5_S4BEG[0] ;
 wire \Tile_X3Y5_S4BEG[10] ;
 wire \Tile_X3Y5_S4BEG[11] ;
 wire \Tile_X3Y5_S4BEG[12] ;
 wire \Tile_X3Y5_S4BEG[13] ;
 wire \Tile_X3Y5_S4BEG[14] ;
 wire \Tile_X3Y5_S4BEG[15] ;
 wire \Tile_X3Y5_S4BEG[1] ;
 wire \Tile_X3Y5_S4BEG[2] ;
 wire \Tile_X3Y5_S4BEG[3] ;
 wire \Tile_X3Y5_S4BEG[4] ;
 wire \Tile_X3Y5_S4BEG[5] ;
 wire \Tile_X3Y5_S4BEG[6] ;
 wire \Tile_X3Y5_S4BEG[7] ;
 wire \Tile_X3Y5_S4BEG[8] ;
 wire \Tile_X3Y5_S4BEG[9] ;
 wire \Tile_X3Y5_SS4BEG[0] ;
 wire \Tile_X3Y5_SS4BEG[10] ;
 wire \Tile_X3Y5_SS4BEG[11] ;
 wire \Tile_X3Y5_SS4BEG[12] ;
 wire \Tile_X3Y5_SS4BEG[13] ;
 wire \Tile_X3Y5_SS4BEG[14] ;
 wire \Tile_X3Y5_SS4BEG[15] ;
 wire \Tile_X3Y5_SS4BEG[1] ;
 wire \Tile_X3Y5_SS4BEG[2] ;
 wire \Tile_X3Y5_SS4BEG[3] ;
 wire \Tile_X3Y5_SS4BEG[4] ;
 wire \Tile_X3Y5_SS4BEG[5] ;
 wire \Tile_X3Y5_SS4BEG[6] ;
 wire \Tile_X3Y5_SS4BEG[7] ;
 wire \Tile_X3Y5_SS4BEG[8] ;
 wire \Tile_X3Y5_SS4BEG[9] ;
 wire Tile_X3Y5_UserCLKo;
 wire \Tile_X3Y5_W1BEG[0] ;
 wire \Tile_X3Y5_W1BEG[1] ;
 wire \Tile_X3Y5_W1BEG[2] ;
 wire \Tile_X3Y5_W1BEG[3] ;
 wire \Tile_X3Y5_W2BEG[0] ;
 wire \Tile_X3Y5_W2BEG[1] ;
 wire \Tile_X3Y5_W2BEG[2] ;
 wire \Tile_X3Y5_W2BEG[3] ;
 wire \Tile_X3Y5_W2BEG[4] ;
 wire \Tile_X3Y5_W2BEG[5] ;
 wire \Tile_X3Y5_W2BEG[6] ;
 wire \Tile_X3Y5_W2BEG[7] ;
 wire \Tile_X3Y5_W2BEGb[0] ;
 wire \Tile_X3Y5_W2BEGb[1] ;
 wire \Tile_X3Y5_W2BEGb[2] ;
 wire \Tile_X3Y5_W2BEGb[3] ;
 wire \Tile_X3Y5_W2BEGb[4] ;
 wire \Tile_X3Y5_W2BEGb[5] ;
 wire \Tile_X3Y5_W2BEGb[6] ;
 wire \Tile_X3Y5_W2BEGb[7] ;
 wire \Tile_X3Y5_W6BEG[0] ;
 wire \Tile_X3Y5_W6BEG[10] ;
 wire \Tile_X3Y5_W6BEG[11] ;
 wire \Tile_X3Y5_W6BEG[1] ;
 wire \Tile_X3Y5_W6BEG[2] ;
 wire \Tile_X3Y5_W6BEG[3] ;
 wire \Tile_X3Y5_W6BEG[4] ;
 wire \Tile_X3Y5_W6BEG[5] ;
 wire \Tile_X3Y5_W6BEG[6] ;
 wire \Tile_X3Y5_W6BEG[7] ;
 wire \Tile_X3Y5_W6BEG[8] ;
 wire \Tile_X3Y5_W6BEG[9] ;
 wire \Tile_X3Y5_WW4BEG[0] ;
 wire \Tile_X3Y5_WW4BEG[10] ;
 wire \Tile_X3Y5_WW4BEG[11] ;
 wire \Tile_X3Y5_WW4BEG[12] ;
 wire \Tile_X3Y5_WW4BEG[13] ;
 wire \Tile_X3Y5_WW4BEG[14] ;
 wire \Tile_X3Y5_WW4BEG[15] ;
 wire \Tile_X3Y5_WW4BEG[1] ;
 wire \Tile_X3Y5_WW4BEG[2] ;
 wire \Tile_X3Y5_WW4BEG[3] ;
 wire \Tile_X3Y5_WW4BEG[4] ;
 wire \Tile_X3Y5_WW4BEG[5] ;
 wire \Tile_X3Y5_WW4BEG[6] ;
 wire \Tile_X3Y5_WW4BEG[7] ;
 wire \Tile_X3Y5_WW4BEG[8] ;
 wire \Tile_X3Y5_WW4BEG[9] ;
 wire Tile_X3Y6_Co;
 wire \Tile_X3Y6_E1BEG[0] ;
 wire \Tile_X3Y6_E1BEG[1] ;
 wire \Tile_X3Y6_E1BEG[2] ;
 wire \Tile_X3Y6_E1BEG[3] ;
 wire \Tile_X3Y6_E2BEG[0] ;
 wire \Tile_X3Y6_E2BEG[1] ;
 wire \Tile_X3Y6_E2BEG[2] ;
 wire \Tile_X3Y6_E2BEG[3] ;
 wire \Tile_X3Y6_E2BEG[4] ;
 wire \Tile_X3Y6_E2BEG[5] ;
 wire \Tile_X3Y6_E2BEG[6] ;
 wire \Tile_X3Y6_E2BEG[7] ;
 wire \Tile_X3Y6_E2BEGb[0] ;
 wire \Tile_X3Y6_E2BEGb[1] ;
 wire \Tile_X3Y6_E2BEGb[2] ;
 wire \Tile_X3Y6_E2BEGb[3] ;
 wire \Tile_X3Y6_E2BEGb[4] ;
 wire \Tile_X3Y6_E2BEGb[5] ;
 wire \Tile_X3Y6_E2BEGb[6] ;
 wire \Tile_X3Y6_E2BEGb[7] ;
 wire \Tile_X3Y6_E6BEG[0] ;
 wire \Tile_X3Y6_E6BEG[10] ;
 wire \Tile_X3Y6_E6BEG[11] ;
 wire \Tile_X3Y6_E6BEG[1] ;
 wire \Tile_X3Y6_E6BEG[2] ;
 wire \Tile_X3Y6_E6BEG[3] ;
 wire \Tile_X3Y6_E6BEG[4] ;
 wire \Tile_X3Y6_E6BEG[5] ;
 wire \Tile_X3Y6_E6BEG[6] ;
 wire \Tile_X3Y6_E6BEG[7] ;
 wire \Tile_X3Y6_E6BEG[8] ;
 wire \Tile_X3Y6_E6BEG[9] ;
 wire \Tile_X3Y6_EE4BEG[0] ;
 wire \Tile_X3Y6_EE4BEG[10] ;
 wire \Tile_X3Y6_EE4BEG[11] ;
 wire \Tile_X3Y6_EE4BEG[12] ;
 wire \Tile_X3Y6_EE4BEG[13] ;
 wire \Tile_X3Y6_EE4BEG[14] ;
 wire \Tile_X3Y6_EE4BEG[15] ;
 wire \Tile_X3Y6_EE4BEG[1] ;
 wire \Tile_X3Y6_EE4BEG[2] ;
 wire \Tile_X3Y6_EE4BEG[3] ;
 wire \Tile_X3Y6_EE4BEG[4] ;
 wire \Tile_X3Y6_EE4BEG[5] ;
 wire \Tile_X3Y6_EE4BEG[6] ;
 wire \Tile_X3Y6_EE4BEG[7] ;
 wire \Tile_X3Y6_EE4BEG[8] ;
 wire \Tile_X3Y6_EE4BEG[9] ;
 wire \Tile_X3Y6_FrameData_O[0] ;
 wire \Tile_X3Y6_FrameData_O[10] ;
 wire \Tile_X3Y6_FrameData_O[11] ;
 wire \Tile_X3Y6_FrameData_O[12] ;
 wire \Tile_X3Y6_FrameData_O[13] ;
 wire \Tile_X3Y6_FrameData_O[14] ;
 wire \Tile_X3Y6_FrameData_O[15] ;
 wire \Tile_X3Y6_FrameData_O[16] ;
 wire \Tile_X3Y6_FrameData_O[17] ;
 wire \Tile_X3Y6_FrameData_O[18] ;
 wire \Tile_X3Y6_FrameData_O[19] ;
 wire \Tile_X3Y6_FrameData_O[1] ;
 wire \Tile_X3Y6_FrameData_O[20] ;
 wire \Tile_X3Y6_FrameData_O[21] ;
 wire \Tile_X3Y6_FrameData_O[22] ;
 wire \Tile_X3Y6_FrameData_O[23] ;
 wire \Tile_X3Y6_FrameData_O[24] ;
 wire \Tile_X3Y6_FrameData_O[25] ;
 wire \Tile_X3Y6_FrameData_O[26] ;
 wire \Tile_X3Y6_FrameData_O[27] ;
 wire \Tile_X3Y6_FrameData_O[28] ;
 wire \Tile_X3Y6_FrameData_O[29] ;
 wire \Tile_X3Y6_FrameData_O[2] ;
 wire \Tile_X3Y6_FrameData_O[30] ;
 wire \Tile_X3Y6_FrameData_O[31] ;
 wire \Tile_X3Y6_FrameData_O[3] ;
 wire \Tile_X3Y6_FrameData_O[4] ;
 wire \Tile_X3Y6_FrameData_O[5] ;
 wire \Tile_X3Y6_FrameData_O[6] ;
 wire \Tile_X3Y6_FrameData_O[7] ;
 wire \Tile_X3Y6_FrameData_O[8] ;
 wire \Tile_X3Y6_FrameData_O[9] ;
 wire \Tile_X3Y6_FrameStrobe_O[0] ;
 wire \Tile_X3Y6_FrameStrobe_O[10] ;
 wire \Tile_X3Y6_FrameStrobe_O[11] ;
 wire \Tile_X3Y6_FrameStrobe_O[12] ;
 wire \Tile_X3Y6_FrameStrobe_O[13] ;
 wire \Tile_X3Y6_FrameStrobe_O[14] ;
 wire \Tile_X3Y6_FrameStrobe_O[15] ;
 wire \Tile_X3Y6_FrameStrobe_O[16] ;
 wire \Tile_X3Y6_FrameStrobe_O[17] ;
 wire \Tile_X3Y6_FrameStrobe_O[18] ;
 wire \Tile_X3Y6_FrameStrobe_O[19] ;
 wire \Tile_X3Y6_FrameStrobe_O[1] ;
 wire \Tile_X3Y6_FrameStrobe_O[2] ;
 wire \Tile_X3Y6_FrameStrobe_O[3] ;
 wire \Tile_X3Y6_FrameStrobe_O[4] ;
 wire \Tile_X3Y6_FrameStrobe_O[5] ;
 wire \Tile_X3Y6_FrameStrobe_O[6] ;
 wire \Tile_X3Y6_FrameStrobe_O[7] ;
 wire \Tile_X3Y6_FrameStrobe_O[8] ;
 wire \Tile_X3Y6_FrameStrobe_O[9] ;
 wire \Tile_X3Y6_N1BEG[0] ;
 wire \Tile_X3Y6_N1BEG[1] ;
 wire \Tile_X3Y6_N1BEG[2] ;
 wire \Tile_X3Y6_N1BEG[3] ;
 wire \Tile_X3Y6_N2BEG[0] ;
 wire \Tile_X3Y6_N2BEG[1] ;
 wire \Tile_X3Y6_N2BEG[2] ;
 wire \Tile_X3Y6_N2BEG[3] ;
 wire \Tile_X3Y6_N2BEG[4] ;
 wire \Tile_X3Y6_N2BEG[5] ;
 wire \Tile_X3Y6_N2BEG[6] ;
 wire \Tile_X3Y6_N2BEG[7] ;
 wire \Tile_X3Y6_N2BEGb[0] ;
 wire \Tile_X3Y6_N2BEGb[1] ;
 wire \Tile_X3Y6_N2BEGb[2] ;
 wire \Tile_X3Y6_N2BEGb[3] ;
 wire \Tile_X3Y6_N2BEGb[4] ;
 wire \Tile_X3Y6_N2BEGb[5] ;
 wire \Tile_X3Y6_N2BEGb[6] ;
 wire \Tile_X3Y6_N2BEGb[7] ;
 wire \Tile_X3Y6_N4BEG[0] ;
 wire \Tile_X3Y6_N4BEG[10] ;
 wire \Tile_X3Y6_N4BEG[11] ;
 wire \Tile_X3Y6_N4BEG[12] ;
 wire \Tile_X3Y6_N4BEG[13] ;
 wire \Tile_X3Y6_N4BEG[14] ;
 wire \Tile_X3Y6_N4BEG[15] ;
 wire \Tile_X3Y6_N4BEG[1] ;
 wire \Tile_X3Y6_N4BEG[2] ;
 wire \Tile_X3Y6_N4BEG[3] ;
 wire \Tile_X3Y6_N4BEG[4] ;
 wire \Tile_X3Y6_N4BEG[5] ;
 wire \Tile_X3Y6_N4BEG[6] ;
 wire \Tile_X3Y6_N4BEG[7] ;
 wire \Tile_X3Y6_N4BEG[8] ;
 wire \Tile_X3Y6_N4BEG[9] ;
 wire \Tile_X3Y6_NN4BEG[0] ;
 wire \Tile_X3Y6_NN4BEG[10] ;
 wire \Tile_X3Y6_NN4BEG[11] ;
 wire \Tile_X3Y6_NN4BEG[12] ;
 wire \Tile_X3Y6_NN4BEG[13] ;
 wire \Tile_X3Y6_NN4BEG[14] ;
 wire \Tile_X3Y6_NN4BEG[15] ;
 wire \Tile_X3Y6_NN4BEG[1] ;
 wire \Tile_X3Y6_NN4BEG[2] ;
 wire \Tile_X3Y6_NN4BEG[3] ;
 wire \Tile_X3Y6_NN4BEG[4] ;
 wire \Tile_X3Y6_NN4BEG[5] ;
 wire \Tile_X3Y6_NN4BEG[6] ;
 wire \Tile_X3Y6_NN4BEG[7] ;
 wire \Tile_X3Y6_NN4BEG[8] ;
 wire \Tile_X3Y6_NN4BEG[9] ;
 wire \Tile_X3Y6_S1BEG[0] ;
 wire \Tile_X3Y6_S1BEG[1] ;
 wire \Tile_X3Y6_S1BEG[2] ;
 wire \Tile_X3Y6_S1BEG[3] ;
 wire \Tile_X3Y6_S2BEG[0] ;
 wire \Tile_X3Y6_S2BEG[1] ;
 wire \Tile_X3Y6_S2BEG[2] ;
 wire \Tile_X3Y6_S2BEG[3] ;
 wire \Tile_X3Y6_S2BEG[4] ;
 wire \Tile_X3Y6_S2BEG[5] ;
 wire \Tile_X3Y6_S2BEG[6] ;
 wire \Tile_X3Y6_S2BEG[7] ;
 wire \Tile_X3Y6_S2BEGb[0] ;
 wire \Tile_X3Y6_S2BEGb[1] ;
 wire \Tile_X3Y6_S2BEGb[2] ;
 wire \Tile_X3Y6_S2BEGb[3] ;
 wire \Tile_X3Y6_S2BEGb[4] ;
 wire \Tile_X3Y6_S2BEGb[5] ;
 wire \Tile_X3Y6_S2BEGb[6] ;
 wire \Tile_X3Y6_S2BEGb[7] ;
 wire \Tile_X3Y6_S4BEG[0] ;
 wire \Tile_X3Y6_S4BEG[10] ;
 wire \Tile_X3Y6_S4BEG[11] ;
 wire \Tile_X3Y6_S4BEG[12] ;
 wire \Tile_X3Y6_S4BEG[13] ;
 wire \Tile_X3Y6_S4BEG[14] ;
 wire \Tile_X3Y6_S4BEG[15] ;
 wire \Tile_X3Y6_S4BEG[1] ;
 wire \Tile_X3Y6_S4BEG[2] ;
 wire \Tile_X3Y6_S4BEG[3] ;
 wire \Tile_X3Y6_S4BEG[4] ;
 wire \Tile_X3Y6_S4BEG[5] ;
 wire \Tile_X3Y6_S4BEG[6] ;
 wire \Tile_X3Y6_S4BEG[7] ;
 wire \Tile_X3Y6_S4BEG[8] ;
 wire \Tile_X3Y6_S4BEG[9] ;
 wire \Tile_X3Y6_SS4BEG[0] ;
 wire \Tile_X3Y6_SS4BEG[10] ;
 wire \Tile_X3Y6_SS4BEG[11] ;
 wire \Tile_X3Y6_SS4BEG[12] ;
 wire \Tile_X3Y6_SS4BEG[13] ;
 wire \Tile_X3Y6_SS4BEG[14] ;
 wire \Tile_X3Y6_SS4BEG[15] ;
 wire \Tile_X3Y6_SS4BEG[1] ;
 wire \Tile_X3Y6_SS4BEG[2] ;
 wire \Tile_X3Y6_SS4BEG[3] ;
 wire \Tile_X3Y6_SS4BEG[4] ;
 wire \Tile_X3Y6_SS4BEG[5] ;
 wire \Tile_X3Y6_SS4BEG[6] ;
 wire \Tile_X3Y6_SS4BEG[7] ;
 wire \Tile_X3Y6_SS4BEG[8] ;
 wire \Tile_X3Y6_SS4BEG[9] ;
 wire Tile_X3Y6_UserCLKo;
 wire \Tile_X3Y6_W1BEG[0] ;
 wire \Tile_X3Y6_W1BEG[1] ;
 wire \Tile_X3Y6_W1BEG[2] ;
 wire \Tile_X3Y6_W1BEG[3] ;
 wire \Tile_X3Y6_W2BEG[0] ;
 wire \Tile_X3Y6_W2BEG[1] ;
 wire \Tile_X3Y6_W2BEG[2] ;
 wire \Tile_X3Y6_W2BEG[3] ;
 wire \Tile_X3Y6_W2BEG[4] ;
 wire \Tile_X3Y6_W2BEG[5] ;
 wire \Tile_X3Y6_W2BEG[6] ;
 wire \Tile_X3Y6_W2BEG[7] ;
 wire \Tile_X3Y6_W2BEGb[0] ;
 wire \Tile_X3Y6_W2BEGb[1] ;
 wire \Tile_X3Y6_W2BEGb[2] ;
 wire \Tile_X3Y6_W2BEGb[3] ;
 wire \Tile_X3Y6_W2BEGb[4] ;
 wire \Tile_X3Y6_W2BEGb[5] ;
 wire \Tile_X3Y6_W2BEGb[6] ;
 wire \Tile_X3Y6_W2BEGb[7] ;
 wire \Tile_X3Y6_W6BEG[0] ;
 wire \Tile_X3Y6_W6BEG[10] ;
 wire \Tile_X3Y6_W6BEG[11] ;
 wire \Tile_X3Y6_W6BEG[1] ;
 wire \Tile_X3Y6_W6BEG[2] ;
 wire \Tile_X3Y6_W6BEG[3] ;
 wire \Tile_X3Y6_W6BEG[4] ;
 wire \Tile_X3Y6_W6BEG[5] ;
 wire \Tile_X3Y6_W6BEG[6] ;
 wire \Tile_X3Y6_W6BEG[7] ;
 wire \Tile_X3Y6_W6BEG[8] ;
 wire \Tile_X3Y6_W6BEG[9] ;
 wire \Tile_X3Y6_WW4BEG[0] ;
 wire \Tile_X3Y6_WW4BEG[10] ;
 wire \Tile_X3Y6_WW4BEG[11] ;
 wire \Tile_X3Y6_WW4BEG[12] ;
 wire \Tile_X3Y6_WW4BEG[13] ;
 wire \Tile_X3Y6_WW4BEG[14] ;
 wire \Tile_X3Y6_WW4BEG[15] ;
 wire \Tile_X3Y6_WW4BEG[1] ;
 wire \Tile_X3Y6_WW4BEG[2] ;
 wire \Tile_X3Y6_WW4BEG[3] ;
 wire \Tile_X3Y6_WW4BEG[4] ;
 wire \Tile_X3Y6_WW4BEG[5] ;
 wire \Tile_X3Y6_WW4BEG[6] ;
 wire \Tile_X3Y6_WW4BEG[7] ;
 wire \Tile_X3Y6_WW4BEG[8] ;
 wire \Tile_X3Y6_WW4BEG[9] ;
 wire Tile_X3Y7_Co;
 wire \Tile_X3Y7_E1BEG[0] ;
 wire \Tile_X3Y7_E1BEG[1] ;
 wire \Tile_X3Y7_E1BEG[2] ;
 wire \Tile_X3Y7_E1BEG[3] ;
 wire \Tile_X3Y7_E2BEG[0] ;
 wire \Tile_X3Y7_E2BEG[1] ;
 wire \Tile_X3Y7_E2BEG[2] ;
 wire \Tile_X3Y7_E2BEG[3] ;
 wire \Tile_X3Y7_E2BEG[4] ;
 wire \Tile_X3Y7_E2BEG[5] ;
 wire \Tile_X3Y7_E2BEG[6] ;
 wire \Tile_X3Y7_E2BEG[7] ;
 wire \Tile_X3Y7_E2BEGb[0] ;
 wire \Tile_X3Y7_E2BEGb[1] ;
 wire \Tile_X3Y7_E2BEGb[2] ;
 wire \Tile_X3Y7_E2BEGb[3] ;
 wire \Tile_X3Y7_E2BEGb[4] ;
 wire \Tile_X3Y7_E2BEGb[5] ;
 wire \Tile_X3Y7_E2BEGb[6] ;
 wire \Tile_X3Y7_E2BEGb[7] ;
 wire \Tile_X3Y7_E6BEG[0] ;
 wire \Tile_X3Y7_E6BEG[10] ;
 wire \Tile_X3Y7_E6BEG[11] ;
 wire \Tile_X3Y7_E6BEG[1] ;
 wire \Tile_X3Y7_E6BEG[2] ;
 wire \Tile_X3Y7_E6BEG[3] ;
 wire \Tile_X3Y7_E6BEG[4] ;
 wire \Tile_X3Y7_E6BEG[5] ;
 wire \Tile_X3Y7_E6BEG[6] ;
 wire \Tile_X3Y7_E6BEG[7] ;
 wire \Tile_X3Y7_E6BEG[8] ;
 wire \Tile_X3Y7_E6BEG[9] ;
 wire \Tile_X3Y7_EE4BEG[0] ;
 wire \Tile_X3Y7_EE4BEG[10] ;
 wire \Tile_X3Y7_EE4BEG[11] ;
 wire \Tile_X3Y7_EE4BEG[12] ;
 wire \Tile_X3Y7_EE4BEG[13] ;
 wire \Tile_X3Y7_EE4BEG[14] ;
 wire \Tile_X3Y7_EE4BEG[15] ;
 wire \Tile_X3Y7_EE4BEG[1] ;
 wire \Tile_X3Y7_EE4BEG[2] ;
 wire \Tile_X3Y7_EE4BEG[3] ;
 wire \Tile_X3Y7_EE4BEG[4] ;
 wire \Tile_X3Y7_EE4BEG[5] ;
 wire \Tile_X3Y7_EE4BEG[6] ;
 wire \Tile_X3Y7_EE4BEG[7] ;
 wire \Tile_X3Y7_EE4BEG[8] ;
 wire \Tile_X3Y7_EE4BEG[9] ;
 wire \Tile_X3Y7_FrameData_O[0] ;
 wire \Tile_X3Y7_FrameData_O[10] ;
 wire \Tile_X3Y7_FrameData_O[11] ;
 wire \Tile_X3Y7_FrameData_O[12] ;
 wire \Tile_X3Y7_FrameData_O[13] ;
 wire \Tile_X3Y7_FrameData_O[14] ;
 wire \Tile_X3Y7_FrameData_O[15] ;
 wire \Tile_X3Y7_FrameData_O[16] ;
 wire \Tile_X3Y7_FrameData_O[17] ;
 wire \Tile_X3Y7_FrameData_O[18] ;
 wire \Tile_X3Y7_FrameData_O[19] ;
 wire \Tile_X3Y7_FrameData_O[1] ;
 wire \Tile_X3Y7_FrameData_O[20] ;
 wire \Tile_X3Y7_FrameData_O[21] ;
 wire \Tile_X3Y7_FrameData_O[22] ;
 wire \Tile_X3Y7_FrameData_O[23] ;
 wire \Tile_X3Y7_FrameData_O[24] ;
 wire \Tile_X3Y7_FrameData_O[25] ;
 wire \Tile_X3Y7_FrameData_O[26] ;
 wire \Tile_X3Y7_FrameData_O[27] ;
 wire \Tile_X3Y7_FrameData_O[28] ;
 wire \Tile_X3Y7_FrameData_O[29] ;
 wire \Tile_X3Y7_FrameData_O[2] ;
 wire \Tile_X3Y7_FrameData_O[30] ;
 wire \Tile_X3Y7_FrameData_O[31] ;
 wire \Tile_X3Y7_FrameData_O[3] ;
 wire \Tile_X3Y7_FrameData_O[4] ;
 wire \Tile_X3Y7_FrameData_O[5] ;
 wire \Tile_X3Y7_FrameData_O[6] ;
 wire \Tile_X3Y7_FrameData_O[7] ;
 wire \Tile_X3Y7_FrameData_O[8] ;
 wire \Tile_X3Y7_FrameData_O[9] ;
 wire \Tile_X3Y7_FrameStrobe_O[0] ;
 wire \Tile_X3Y7_FrameStrobe_O[10] ;
 wire \Tile_X3Y7_FrameStrobe_O[11] ;
 wire \Tile_X3Y7_FrameStrobe_O[12] ;
 wire \Tile_X3Y7_FrameStrobe_O[13] ;
 wire \Tile_X3Y7_FrameStrobe_O[14] ;
 wire \Tile_X3Y7_FrameStrobe_O[15] ;
 wire \Tile_X3Y7_FrameStrobe_O[16] ;
 wire \Tile_X3Y7_FrameStrobe_O[17] ;
 wire \Tile_X3Y7_FrameStrobe_O[18] ;
 wire \Tile_X3Y7_FrameStrobe_O[19] ;
 wire \Tile_X3Y7_FrameStrobe_O[1] ;
 wire \Tile_X3Y7_FrameStrobe_O[2] ;
 wire \Tile_X3Y7_FrameStrobe_O[3] ;
 wire \Tile_X3Y7_FrameStrobe_O[4] ;
 wire \Tile_X3Y7_FrameStrobe_O[5] ;
 wire \Tile_X3Y7_FrameStrobe_O[6] ;
 wire \Tile_X3Y7_FrameStrobe_O[7] ;
 wire \Tile_X3Y7_FrameStrobe_O[8] ;
 wire \Tile_X3Y7_FrameStrobe_O[9] ;
 wire \Tile_X3Y7_N1BEG[0] ;
 wire \Tile_X3Y7_N1BEG[1] ;
 wire \Tile_X3Y7_N1BEG[2] ;
 wire \Tile_X3Y7_N1BEG[3] ;
 wire \Tile_X3Y7_N2BEG[0] ;
 wire \Tile_X3Y7_N2BEG[1] ;
 wire \Tile_X3Y7_N2BEG[2] ;
 wire \Tile_X3Y7_N2BEG[3] ;
 wire \Tile_X3Y7_N2BEG[4] ;
 wire \Tile_X3Y7_N2BEG[5] ;
 wire \Tile_X3Y7_N2BEG[6] ;
 wire \Tile_X3Y7_N2BEG[7] ;
 wire \Tile_X3Y7_N2BEGb[0] ;
 wire \Tile_X3Y7_N2BEGb[1] ;
 wire \Tile_X3Y7_N2BEGb[2] ;
 wire \Tile_X3Y7_N2BEGb[3] ;
 wire \Tile_X3Y7_N2BEGb[4] ;
 wire \Tile_X3Y7_N2BEGb[5] ;
 wire \Tile_X3Y7_N2BEGb[6] ;
 wire \Tile_X3Y7_N2BEGb[7] ;
 wire \Tile_X3Y7_N4BEG[0] ;
 wire \Tile_X3Y7_N4BEG[10] ;
 wire \Tile_X3Y7_N4BEG[11] ;
 wire \Tile_X3Y7_N4BEG[12] ;
 wire \Tile_X3Y7_N4BEG[13] ;
 wire \Tile_X3Y7_N4BEG[14] ;
 wire \Tile_X3Y7_N4BEG[15] ;
 wire \Tile_X3Y7_N4BEG[1] ;
 wire \Tile_X3Y7_N4BEG[2] ;
 wire \Tile_X3Y7_N4BEG[3] ;
 wire \Tile_X3Y7_N4BEG[4] ;
 wire \Tile_X3Y7_N4BEG[5] ;
 wire \Tile_X3Y7_N4BEG[6] ;
 wire \Tile_X3Y7_N4BEG[7] ;
 wire \Tile_X3Y7_N4BEG[8] ;
 wire \Tile_X3Y7_N4BEG[9] ;
 wire \Tile_X3Y7_NN4BEG[0] ;
 wire \Tile_X3Y7_NN4BEG[10] ;
 wire \Tile_X3Y7_NN4BEG[11] ;
 wire \Tile_X3Y7_NN4BEG[12] ;
 wire \Tile_X3Y7_NN4BEG[13] ;
 wire \Tile_X3Y7_NN4BEG[14] ;
 wire \Tile_X3Y7_NN4BEG[15] ;
 wire \Tile_X3Y7_NN4BEG[1] ;
 wire \Tile_X3Y7_NN4BEG[2] ;
 wire \Tile_X3Y7_NN4BEG[3] ;
 wire \Tile_X3Y7_NN4BEG[4] ;
 wire \Tile_X3Y7_NN4BEG[5] ;
 wire \Tile_X3Y7_NN4BEG[6] ;
 wire \Tile_X3Y7_NN4BEG[7] ;
 wire \Tile_X3Y7_NN4BEG[8] ;
 wire \Tile_X3Y7_NN4BEG[9] ;
 wire \Tile_X3Y7_S1BEG[0] ;
 wire \Tile_X3Y7_S1BEG[1] ;
 wire \Tile_X3Y7_S1BEG[2] ;
 wire \Tile_X3Y7_S1BEG[3] ;
 wire \Tile_X3Y7_S2BEG[0] ;
 wire \Tile_X3Y7_S2BEG[1] ;
 wire \Tile_X3Y7_S2BEG[2] ;
 wire \Tile_X3Y7_S2BEG[3] ;
 wire \Tile_X3Y7_S2BEG[4] ;
 wire \Tile_X3Y7_S2BEG[5] ;
 wire \Tile_X3Y7_S2BEG[6] ;
 wire \Tile_X3Y7_S2BEG[7] ;
 wire \Tile_X3Y7_S2BEGb[0] ;
 wire \Tile_X3Y7_S2BEGb[1] ;
 wire \Tile_X3Y7_S2BEGb[2] ;
 wire \Tile_X3Y7_S2BEGb[3] ;
 wire \Tile_X3Y7_S2BEGb[4] ;
 wire \Tile_X3Y7_S2BEGb[5] ;
 wire \Tile_X3Y7_S2BEGb[6] ;
 wire \Tile_X3Y7_S2BEGb[7] ;
 wire \Tile_X3Y7_S4BEG[0] ;
 wire \Tile_X3Y7_S4BEG[10] ;
 wire \Tile_X3Y7_S4BEG[11] ;
 wire \Tile_X3Y7_S4BEG[12] ;
 wire \Tile_X3Y7_S4BEG[13] ;
 wire \Tile_X3Y7_S4BEG[14] ;
 wire \Tile_X3Y7_S4BEG[15] ;
 wire \Tile_X3Y7_S4BEG[1] ;
 wire \Tile_X3Y7_S4BEG[2] ;
 wire \Tile_X3Y7_S4BEG[3] ;
 wire \Tile_X3Y7_S4BEG[4] ;
 wire \Tile_X3Y7_S4BEG[5] ;
 wire \Tile_X3Y7_S4BEG[6] ;
 wire \Tile_X3Y7_S4BEG[7] ;
 wire \Tile_X3Y7_S4BEG[8] ;
 wire \Tile_X3Y7_S4BEG[9] ;
 wire \Tile_X3Y7_SS4BEG[0] ;
 wire \Tile_X3Y7_SS4BEG[10] ;
 wire \Tile_X3Y7_SS4BEG[11] ;
 wire \Tile_X3Y7_SS4BEG[12] ;
 wire \Tile_X3Y7_SS4BEG[13] ;
 wire \Tile_X3Y7_SS4BEG[14] ;
 wire \Tile_X3Y7_SS4BEG[15] ;
 wire \Tile_X3Y7_SS4BEG[1] ;
 wire \Tile_X3Y7_SS4BEG[2] ;
 wire \Tile_X3Y7_SS4BEG[3] ;
 wire \Tile_X3Y7_SS4BEG[4] ;
 wire \Tile_X3Y7_SS4BEG[5] ;
 wire \Tile_X3Y7_SS4BEG[6] ;
 wire \Tile_X3Y7_SS4BEG[7] ;
 wire \Tile_X3Y7_SS4BEG[8] ;
 wire \Tile_X3Y7_SS4BEG[9] ;
 wire Tile_X3Y7_UserCLKo;
 wire \Tile_X3Y7_W1BEG[0] ;
 wire \Tile_X3Y7_W1BEG[1] ;
 wire \Tile_X3Y7_W1BEG[2] ;
 wire \Tile_X3Y7_W1BEG[3] ;
 wire \Tile_X3Y7_W2BEG[0] ;
 wire \Tile_X3Y7_W2BEG[1] ;
 wire \Tile_X3Y7_W2BEG[2] ;
 wire \Tile_X3Y7_W2BEG[3] ;
 wire \Tile_X3Y7_W2BEG[4] ;
 wire \Tile_X3Y7_W2BEG[5] ;
 wire \Tile_X3Y7_W2BEG[6] ;
 wire \Tile_X3Y7_W2BEG[7] ;
 wire \Tile_X3Y7_W2BEGb[0] ;
 wire \Tile_X3Y7_W2BEGb[1] ;
 wire \Tile_X3Y7_W2BEGb[2] ;
 wire \Tile_X3Y7_W2BEGb[3] ;
 wire \Tile_X3Y7_W2BEGb[4] ;
 wire \Tile_X3Y7_W2BEGb[5] ;
 wire \Tile_X3Y7_W2BEGb[6] ;
 wire \Tile_X3Y7_W2BEGb[7] ;
 wire \Tile_X3Y7_W6BEG[0] ;
 wire \Tile_X3Y7_W6BEG[10] ;
 wire \Tile_X3Y7_W6BEG[11] ;
 wire \Tile_X3Y7_W6BEG[1] ;
 wire \Tile_X3Y7_W6BEG[2] ;
 wire \Tile_X3Y7_W6BEG[3] ;
 wire \Tile_X3Y7_W6BEG[4] ;
 wire \Tile_X3Y7_W6BEG[5] ;
 wire \Tile_X3Y7_W6BEG[6] ;
 wire \Tile_X3Y7_W6BEG[7] ;
 wire \Tile_X3Y7_W6BEG[8] ;
 wire \Tile_X3Y7_W6BEG[9] ;
 wire \Tile_X3Y7_WW4BEG[0] ;
 wire \Tile_X3Y7_WW4BEG[10] ;
 wire \Tile_X3Y7_WW4BEG[11] ;
 wire \Tile_X3Y7_WW4BEG[12] ;
 wire \Tile_X3Y7_WW4BEG[13] ;
 wire \Tile_X3Y7_WW4BEG[14] ;
 wire \Tile_X3Y7_WW4BEG[15] ;
 wire \Tile_X3Y7_WW4BEG[1] ;
 wire \Tile_X3Y7_WW4BEG[2] ;
 wire \Tile_X3Y7_WW4BEG[3] ;
 wire \Tile_X3Y7_WW4BEG[4] ;
 wire \Tile_X3Y7_WW4BEG[5] ;
 wire \Tile_X3Y7_WW4BEG[6] ;
 wire \Tile_X3Y7_WW4BEG[7] ;
 wire \Tile_X3Y7_WW4BEG[8] ;
 wire \Tile_X3Y7_WW4BEG[9] ;
 wire Tile_X3Y8_Co;
 wire \Tile_X3Y8_E1BEG[0] ;
 wire \Tile_X3Y8_E1BEG[1] ;
 wire \Tile_X3Y8_E1BEG[2] ;
 wire \Tile_X3Y8_E1BEG[3] ;
 wire \Tile_X3Y8_E2BEG[0] ;
 wire \Tile_X3Y8_E2BEG[1] ;
 wire \Tile_X3Y8_E2BEG[2] ;
 wire \Tile_X3Y8_E2BEG[3] ;
 wire \Tile_X3Y8_E2BEG[4] ;
 wire \Tile_X3Y8_E2BEG[5] ;
 wire \Tile_X3Y8_E2BEG[6] ;
 wire \Tile_X3Y8_E2BEG[7] ;
 wire \Tile_X3Y8_E2BEGb[0] ;
 wire \Tile_X3Y8_E2BEGb[1] ;
 wire \Tile_X3Y8_E2BEGb[2] ;
 wire \Tile_X3Y8_E2BEGb[3] ;
 wire \Tile_X3Y8_E2BEGb[4] ;
 wire \Tile_X3Y8_E2BEGb[5] ;
 wire \Tile_X3Y8_E2BEGb[6] ;
 wire \Tile_X3Y8_E2BEGb[7] ;
 wire \Tile_X3Y8_E6BEG[0] ;
 wire \Tile_X3Y8_E6BEG[10] ;
 wire \Tile_X3Y8_E6BEG[11] ;
 wire \Tile_X3Y8_E6BEG[1] ;
 wire \Tile_X3Y8_E6BEG[2] ;
 wire \Tile_X3Y8_E6BEG[3] ;
 wire \Tile_X3Y8_E6BEG[4] ;
 wire \Tile_X3Y8_E6BEG[5] ;
 wire \Tile_X3Y8_E6BEG[6] ;
 wire \Tile_X3Y8_E6BEG[7] ;
 wire \Tile_X3Y8_E6BEG[8] ;
 wire \Tile_X3Y8_E6BEG[9] ;
 wire \Tile_X3Y8_EE4BEG[0] ;
 wire \Tile_X3Y8_EE4BEG[10] ;
 wire \Tile_X3Y8_EE4BEG[11] ;
 wire \Tile_X3Y8_EE4BEG[12] ;
 wire \Tile_X3Y8_EE4BEG[13] ;
 wire \Tile_X3Y8_EE4BEG[14] ;
 wire \Tile_X3Y8_EE4BEG[15] ;
 wire \Tile_X3Y8_EE4BEG[1] ;
 wire \Tile_X3Y8_EE4BEG[2] ;
 wire \Tile_X3Y8_EE4BEG[3] ;
 wire \Tile_X3Y8_EE4BEG[4] ;
 wire \Tile_X3Y8_EE4BEG[5] ;
 wire \Tile_X3Y8_EE4BEG[6] ;
 wire \Tile_X3Y8_EE4BEG[7] ;
 wire \Tile_X3Y8_EE4BEG[8] ;
 wire \Tile_X3Y8_EE4BEG[9] ;
 wire \Tile_X3Y8_FrameData_O[0] ;
 wire \Tile_X3Y8_FrameData_O[10] ;
 wire \Tile_X3Y8_FrameData_O[11] ;
 wire \Tile_X3Y8_FrameData_O[12] ;
 wire \Tile_X3Y8_FrameData_O[13] ;
 wire \Tile_X3Y8_FrameData_O[14] ;
 wire \Tile_X3Y8_FrameData_O[15] ;
 wire \Tile_X3Y8_FrameData_O[16] ;
 wire \Tile_X3Y8_FrameData_O[17] ;
 wire \Tile_X3Y8_FrameData_O[18] ;
 wire \Tile_X3Y8_FrameData_O[19] ;
 wire \Tile_X3Y8_FrameData_O[1] ;
 wire \Tile_X3Y8_FrameData_O[20] ;
 wire \Tile_X3Y8_FrameData_O[21] ;
 wire \Tile_X3Y8_FrameData_O[22] ;
 wire \Tile_X3Y8_FrameData_O[23] ;
 wire \Tile_X3Y8_FrameData_O[24] ;
 wire \Tile_X3Y8_FrameData_O[25] ;
 wire \Tile_X3Y8_FrameData_O[26] ;
 wire \Tile_X3Y8_FrameData_O[27] ;
 wire \Tile_X3Y8_FrameData_O[28] ;
 wire \Tile_X3Y8_FrameData_O[29] ;
 wire \Tile_X3Y8_FrameData_O[2] ;
 wire \Tile_X3Y8_FrameData_O[30] ;
 wire \Tile_X3Y8_FrameData_O[31] ;
 wire \Tile_X3Y8_FrameData_O[3] ;
 wire \Tile_X3Y8_FrameData_O[4] ;
 wire \Tile_X3Y8_FrameData_O[5] ;
 wire \Tile_X3Y8_FrameData_O[6] ;
 wire \Tile_X3Y8_FrameData_O[7] ;
 wire \Tile_X3Y8_FrameData_O[8] ;
 wire \Tile_X3Y8_FrameData_O[9] ;
 wire \Tile_X3Y8_FrameStrobe_O[0] ;
 wire \Tile_X3Y8_FrameStrobe_O[10] ;
 wire \Tile_X3Y8_FrameStrobe_O[11] ;
 wire \Tile_X3Y8_FrameStrobe_O[12] ;
 wire \Tile_X3Y8_FrameStrobe_O[13] ;
 wire \Tile_X3Y8_FrameStrobe_O[14] ;
 wire \Tile_X3Y8_FrameStrobe_O[15] ;
 wire \Tile_X3Y8_FrameStrobe_O[16] ;
 wire \Tile_X3Y8_FrameStrobe_O[17] ;
 wire \Tile_X3Y8_FrameStrobe_O[18] ;
 wire \Tile_X3Y8_FrameStrobe_O[19] ;
 wire \Tile_X3Y8_FrameStrobe_O[1] ;
 wire \Tile_X3Y8_FrameStrobe_O[2] ;
 wire \Tile_X3Y8_FrameStrobe_O[3] ;
 wire \Tile_X3Y8_FrameStrobe_O[4] ;
 wire \Tile_X3Y8_FrameStrobe_O[5] ;
 wire \Tile_X3Y8_FrameStrobe_O[6] ;
 wire \Tile_X3Y8_FrameStrobe_O[7] ;
 wire \Tile_X3Y8_FrameStrobe_O[8] ;
 wire \Tile_X3Y8_FrameStrobe_O[9] ;
 wire \Tile_X3Y8_N1BEG[0] ;
 wire \Tile_X3Y8_N1BEG[1] ;
 wire \Tile_X3Y8_N1BEG[2] ;
 wire \Tile_X3Y8_N1BEG[3] ;
 wire \Tile_X3Y8_N2BEG[0] ;
 wire \Tile_X3Y8_N2BEG[1] ;
 wire \Tile_X3Y8_N2BEG[2] ;
 wire \Tile_X3Y8_N2BEG[3] ;
 wire \Tile_X3Y8_N2BEG[4] ;
 wire \Tile_X3Y8_N2BEG[5] ;
 wire \Tile_X3Y8_N2BEG[6] ;
 wire \Tile_X3Y8_N2BEG[7] ;
 wire \Tile_X3Y8_N2BEGb[0] ;
 wire \Tile_X3Y8_N2BEGb[1] ;
 wire \Tile_X3Y8_N2BEGb[2] ;
 wire \Tile_X3Y8_N2BEGb[3] ;
 wire \Tile_X3Y8_N2BEGb[4] ;
 wire \Tile_X3Y8_N2BEGb[5] ;
 wire \Tile_X3Y8_N2BEGb[6] ;
 wire \Tile_X3Y8_N2BEGb[7] ;
 wire \Tile_X3Y8_N4BEG[0] ;
 wire \Tile_X3Y8_N4BEG[10] ;
 wire \Tile_X3Y8_N4BEG[11] ;
 wire \Tile_X3Y8_N4BEG[12] ;
 wire \Tile_X3Y8_N4BEG[13] ;
 wire \Tile_X3Y8_N4BEG[14] ;
 wire \Tile_X3Y8_N4BEG[15] ;
 wire \Tile_X3Y8_N4BEG[1] ;
 wire \Tile_X3Y8_N4BEG[2] ;
 wire \Tile_X3Y8_N4BEG[3] ;
 wire \Tile_X3Y8_N4BEG[4] ;
 wire \Tile_X3Y8_N4BEG[5] ;
 wire \Tile_X3Y8_N4BEG[6] ;
 wire \Tile_X3Y8_N4BEG[7] ;
 wire \Tile_X3Y8_N4BEG[8] ;
 wire \Tile_X3Y8_N4BEG[9] ;
 wire \Tile_X3Y8_NN4BEG[0] ;
 wire \Tile_X3Y8_NN4BEG[10] ;
 wire \Tile_X3Y8_NN4BEG[11] ;
 wire \Tile_X3Y8_NN4BEG[12] ;
 wire \Tile_X3Y8_NN4BEG[13] ;
 wire \Tile_X3Y8_NN4BEG[14] ;
 wire \Tile_X3Y8_NN4BEG[15] ;
 wire \Tile_X3Y8_NN4BEG[1] ;
 wire \Tile_X3Y8_NN4BEG[2] ;
 wire \Tile_X3Y8_NN4BEG[3] ;
 wire \Tile_X3Y8_NN4BEG[4] ;
 wire \Tile_X3Y8_NN4BEG[5] ;
 wire \Tile_X3Y8_NN4BEG[6] ;
 wire \Tile_X3Y8_NN4BEG[7] ;
 wire \Tile_X3Y8_NN4BEG[8] ;
 wire \Tile_X3Y8_NN4BEG[9] ;
 wire \Tile_X3Y8_S1BEG[0] ;
 wire \Tile_X3Y8_S1BEG[1] ;
 wire \Tile_X3Y8_S1BEG[2] ;
 wire \Tile_X3Y8_S1BEG[3] ;
 wire \Tile_X3Y8_S2BEG[0] ;
 wire \Tile_X3Y8_S2BEG[1] ;
 wire \Tile_X3Y8_S2BEG[2] ;
 wire \Tile_X3Y8_S2BEG[3] ;
 wire \Tile_X3Y8_S2BEG[4] ;
 wire \Tile_X3Y8_S2BEG[5] ;
 wire \Tile_X3Y8_S2BEG[6] ;
 wire \Tile_X3Y8_S2BEG[7] ;
 wire \Tile_X3Y8_S2BEGb[0] ;
 wire \Tile_X3Y8_S2BEGb[1] ;
 wire \Tile_X3Y8_S2BEGb[2] ;
 wire \Tile_X3Y8_S2BEGb[3] ;
 wire \Tile_X3Y8_S2BEGb[4] ;
 wire \Tile_X3Y8_S2BEGb[5] ;
 wire \Tile_X3Y8_S2BEGb[6] ;
 wire \Tile_X3Y8_S2BEGb[7] ;
 wire \Tile_X3Y8_S4BEG[0] ;
 wire \Tile_X3Y8_S4BEG[10] ;
 wire \Tile_X3Y8_S4BEG[11] ;
 wire \Tile_X3Y8_S4BEG[12] ;
 wire \Tile_X3Y8_S4BEG[13] ;
 wire \Tile_X3Y8_S4BEG[14] ;
 wire \Tile_X3Y8_S4BEG[15] ;
 wire \Tile_X3Y8_S4BEG[1] ;
 wire \Tile_X3Y8_S4BEG[2] ;
 wire \Tile_X3Y8_S4BEG[3] ;
 wire \Tile_X3Y8_S4BEG[4] ;
 wire \Tile_X3Y8_S4BEG[5] ;
 wire \Tile_X3Y8_S4BEG[6] ;
 wire \Tile_X3Y8_S4BEG[7] ;
 wire \Tile_X3Y8_S4BEG[8] ;
 wire \Tile_X3Y8_S4BEG[9] ;
 wire \Tile_X3Y8_SS4BEG[0] ;
 wire \Tile_X3Y8_SS4BEG[10] ;
 wire \Tile_X3Y8_SS4BEG[11] ;
 wire \Tile_X3Y8_SS4BEG[12] ;
 wire \Tile_X3Y8_SS4BEG[13] ;
 wire \Tile_X3Y8_SS4BEG[14] ;
 wire \Tile_X3Y8_SS4BEG[15] ;
 wire \Tile_X3Y8_SS4BEG[1] ;
 wire \Tile_X3Y8_SS4BEG[2] ;
 wire \Tile_X3Y8_SS4BEG[3] ;
 wire \Tile_X3Y8_SS4BEG[4] ;
 wire \Tile_X3Y8_SS4BEG[5] ;
 wire \Tile_X3Y8_SS4BEG[6] ;
 wire \Tile_X3Y8_SS4BEG[7] ;
 wire \Tile_X3Y8_SS4BEG[8] ;
 wire \Tile_X3Y8_SS4BEG[9] ;
 wire Tile_X3Y8_UserCLKo;
 wire \Tile_X3Y8_W1BEG[0] ;
 wire \Tile_X3Y8_W1BEG[1] ;
 wire \Tile_X3Y8_W1BEG[2] ;
 wire \Tile_X3Y8_W1BEG[3] ;
 wire \Tile_X3Y8_W2BEG[0] ;
 wire \Tile_X3Y8_W2BEG[1] ;
 wire \Tile_X3Y8_W2BEG[2] ;
 wire \Tile_X3Y8_W2BEG[3] ;
 wire \Tile_X3Y8_W2BEG[4] ;
 wire \Tile_X3Y8_W2BEG[5] ;
 wire \Tile_X3Y8_W2BEG[6] ;
 wire \Tile_X3Y8_W2BEG[7] ;
 wire \Tile_X3Y8_W2BEGb[0] ;
 wire \Tile_X3Y8_W2BEGb[1] ;
 wire \Tile_X3Y8_W2BEGb[2] ;
 wire \Tile_X3Y8_W2BEGb[3] ;
 wire \Tile_X3Y8_W2BEGb[4] ;
 wire \Tile_X3Y8_W2BEGb[5] ;
 wire \Tile_X3Y8_W2BEGb[6] ;
 wire \Tile_X3Y8_W2BEGb[7] ;
 wire \Tile_X3Y8_W6BEG[0] ;
 wire \Tile_X3Y8_W6BEG[10] ;
 wire \Tile_X3Y8_W6BEG[11] ;
 wire \Tile_X3Y8_W6BEG[1] ;
 wire \Tile_X3Y8_W6BEG[2] ;
 wire \Tile_X3Y8_W6BEG[3] ;
 wire \Tile_X3Y8_W6BEG[4] ;
 wire \Tile_X3Y8_W6BEG[5] ;
 wire \Tile_X3Y8_W6BEG[6] ;
 wire \Tile_X3Y8_W6BEG[7] ;
 wire \Tile_X3Y8_W6BEG[8] ;
 wire \Tile_X3Y8_W6BEG[9] ;
 wire \Tile_X3Y8_WW4BEG[0] ;
 wire \Tile_X3Y8_WW4BEG[10] ;
 wire \Tile_X3Y8_WW4BEG[11] ;
 wire \Tile_X3Y8_WW4BEG[12] ;
 wire \Tile_X3Y8_WW4BEG[13] ;
 wire \Tile_X3Y8_WW4BEG[14] ;
 wire \Tile_X3Y8_WW4BEG[15] ;
 wire \Tile_X3Y8_WW4BEG[1] ;
 wire \Tile_X3Y8_WW4BEG[2] ;
 wire \Tile_X3Y8_WW4BEG[3] ;
 wire \Tile_X3Y8_WW4BEG[4] ;
 wire \Tile_X3Y8_WW4BEG[5] ;
 wire \Tile_X3Y8_WW4BEG[6] ;
 wire \Tile_X3Y8_WW4BEG[7] ;
 wire \Tile_X3Y8_WW4BEG[8] ;
 wire \Tile_X3Y8_WW4BEG[9] ;
 wire Tile_X3Y9_Co;
 wire \Tile_X3Y9_FrameData_O[0] ;
 wire \Tile_X3Y9_FrameData_O[10] ;
 wire \Tile_X3Y9_FrameData_O[11] ;
 wire \Tile_X3Y9_FrameData_O[12] ;
 wire \Tile_X3Y9_FrameData_O[13] ;
 wire \Tile_X3Y9_FrameData_O[14] ;
 wire \Tile_X3Y9_FrameData_O[15] ;
 wire \Tile_X3Y9_FrameData_O[16] ;
 wire \Tile_X3Y9_FrameData_O[17] ;
 wire \Tile_X3Y9_FrameData_O[18] ;
 wire \Tile_X3Y9_FrameData_O[19] ;
 wire \Tile_X3Y9_FrameData_O[1] ;
 wire \Tile_X3Y9_FrameData_O[20] ;
 wire \Tile_X3Y9_FrameData_O[21] ;
 wire \Tile_X3Y9_FrameData_O[22] ;
 wire \Tile_X3Y9_FrameData_O[23] ;
 wire \Tile_X3Y9_FrameData_O[24] ;
 wire \Tile_X3Y9_FrameData_O[25] ;
 wire \Tile_X3Y9_FrameData_O[26] ;
 wire \Tile_X3Y9_FrameData_O[27] ;
 wire \Tile_X3Y9_FrameData_O[28] ;
 wire \Tile_X3Y9_FrameData_O[29] ;
 wire \Tile_X3Y9_FrameData_O[2] ;
 wire \Tile_X3Y9_FrameData_O[30] ;
 wire \Tile_X3Y9_FrameData_O[31] ;
 wire \Tile_X3Y9_FrameData_O[3] ;
 wire \Tile_X3Y9_FrameData_O[4] ;
 wire \Tile_X3Y9_FrameData_O[5] ;
 wire \Tile_X3Y9_FrameData_O[6] ;
 wire \Tile_X3Y9_FrameData_O[7] ;
 wire \Tile_X3Y9_FrameData_O[8] ;
 wire \Tile_X3Y9_FrameData_O[9] ;
 wire \Tile_X3Y9_FrameStrobe_O[0] ;
 wire \Tile_X3Y9_FrameStrobe_O[10] ;
 wire \Tile_X3Y9_FrameStrobe_O[11] ;
 wire \Tile_X3Y9_FrameStrobe_O[12] ;
 wire \Tile_X3Y9_FrameStrobe_O[13] ;
 wire \Tile_X3Y9_FrameStrobe_O[14] ;
 wire \Tile_X3Y9_FrameStrobe_O[15] ;
 wire \Tile_X3Y9_FrameStrobe_O[16] ;
 wire \Tile_X3Y9_FrameStrobe_O[17] ;
 wire \Tile_X3Y9_FrameStrobe_O[18] ;
 wire \Tile_X3Y9_FrameStrobe_O[19] ;
 wire \Tile_X3Y9_FrameStrobe_O[1] ;
 wire \Tile_X3Y9_FrameStrobe_O[2] ;
 wire \Tile_X3Y9_FrameStrobe_O[3] ;
 wire \Tile_X3Y9_FrameStrobe_O[4] ;
 wire \Tile_X3Y9_FrameStrobe_O[5] ;
 wire \Tile_X3Y9_FrameStrobe_O[6] ;
 wire \Tile_X3Y9_FrameStrobe_O[7] ;
 wire \Tile_X3Y9_FrameStrobe_O[8] ;
 wire \Tile_X3Y9_FrameStrobe_O[9] ;
 wire \Tile_X3Y9_N1BEG[0] ;
 wire \Tile_X3Y9_N1BEG[1] ;
 wire \Tile_X3Y9_N1BEG[2] ;
 wire \Tile_X3Y9_N1BEG[3] ;
 wire \Tile_X3Y9_N2BEG[0] ;
 wire \Tile_X3Y9_N2BEG[1] ;
 wire \Tile_X3Y9_N2BEG[2] ;
 wire \Tile_X3Y9_N2BEG[3] ;
 wire \Tile_X3Y9_N2BEG[4] ;
 wire \Tile_X3Y9_N2BEG[5] ;
 wire \Tile_X3Y9_N2BEG[6] ;
 wire \Tile_X3Y9_N2BEG[7] ;
 wire \Tile_X3Y9_N2BEGb[0] ;
 wire \Tile_X3Y9_N2BEGb[1] ;
 wire \Tile_X3Y9_N2BEGb[2] ;
 wire \Tile_X3Y9_N2BEGb[3] ;
 wire \Tile_X3Y9_N2BEGb[4] ;
 wire \Tile_X3Y9_N2BEGb[5] ;
 wire \Tile_X3Y9_N2BEGb[6] ;
 wire \Tile_X3Y9_N2BEGb[7] ;
 wire \Tile_X3Y9_N4BEG[0] ;
 wire \Tile_X3Y9_N4BEG[10] ;
 wire \Tile_X3Y9_N4BEG[11] ;
 wire \Tile_X3Y9_N4BEG[12] ;
 wire \Tile_X3Y9_N4BEG[13] ;
 wire \Tile_X3Y9_N4BEG[14] ;
 wire \Tile_X3Y9_N4BEG[15] ;
 wire \Tile_X3Y9_N4BEG[1] ;
 wire \Tile_X3Y9_N4BEG[2] ;
 wire \Tile_X3Y9_N4BEG[3] ;
 wire \Tile_X3Y9_N4BEG[4] ;
 wire \Tile_X3Y9_N4BEG[5] ;
 wire \Tile_X3Y9_N4BEG[6] ;
 wire \Tile_X3Y9_N4BEG[7] ;
 wire \Tile_X3Y9_N4BEG[8] ;
 wire \Tile_X3Y9_N4BEG[9] ;
 wire \Tile_X3Y9_NN4BEG[0] ;
 wire \Tile_X3Y9_NN4BEG[10] ;
 wire \Tile_X3Y9_NN4BEG[11] ;
 wire \Tile_X3Y9_NN4BEG[12] ;
 wire \Tile_X3Y9_NN4BEG[13] ;
 wire \Tile_X3Y9_NN4BEG[14] ;
 wire \Tile_X3Y9_NN4BEG[15] ;
 wire \Tile_X3Y9_NN4BEG[1] ;
 wire \Tile_X3Y9_NN4BEG[2] ;
 wire \Tile_X3Y9_NN4BEG[3] ;
 wire \Tile_X3Y9_NN4BEG[4] ;
 wire \Tile_X3Y9_NN4BEG[5] ;
 wire \Tile_X3Y9_NN4BEG[6] ;
 wire \Tile_X3Y9_NN4BEG[7] ;
 wire \Tile_X3Y9_NN4BEG[8] ;
 wire \Tile_X3Y9_NN4BEG[9] ;
 wire Tile_X3Y9_UserCLKo;
 wire \Tile_X4Y0_FrameData_O[0] ;
 wire \Tile_X4Y0_FrameData_O[10] ;
 wire \Tile_X4Y0_FrameData_O[11] ;
 wire \Tile_X4Y0_FrameData_O[12] ;
 wire \Tile_X4Y0_FrameData_O[13] ;
 wire \Tile_X4Y0_FrameData_O[14] ;
 wire \Tile_X4Y0_FrameData_O[15] ;
 wire \Tile_X4Y0_FrameData_O[16] ;
 wire \Tile_X4Y0_FrameData_O[17] ;
 wire \Tile_X4Y0_FrameData_O[18] ;
 wire \Tile_X4Y0_FrameData_O[19] ;
 wire \Tile_X4Y0_FrameData_O[1] ;
 wire \Tile_X4Y0_FrameData_O[20] ;
 wire \Tile_X4Y0_FrameData_O[21] ;
 wire \Tile_X4Y0_FrameData_O[22] ;
 wire \Tile_X4Y0_FrameData_O[23] ;
 wire \Tile_X4Y0_FrameData_O[24] ;
 wire \Tile_X4Y0_FrameData_O[25] ;
 wire \Tile_X4Y0_FrameData_O[26] ;
 wire \Tile_X4Y0_FrameData_O[27] ;
 wire \Tile_X4Y0_FrameData_O[28] ;
 wire \Tile_X4Y0_FrameData_O[29] ;
 wire \Tile_X4Y0_FrameData_O[2] ;
 wire \Tile_X4Y0_FrameData_O[30] ;
 wire \Tile_X4Y0_FrameData_O[31] ;
 wire \Tile_X4Y0_FrameData_O[3] ;
 wire \Tile_X4Y0_FrameData_O[4] ;
 wire \Tile_X4Y0_FrameData_O[5] ;
 wire \Tile_X4Y0_FrameData_O[6] ;
 wire \Tile_X4Y0_FrameData_O[7] ;
 wire \Tile_X4Y0_FrameData_O[8] ;
 wire \Tile_X4Y0_FrameData_O[9] ;
 wire \Tile_X4Y0_FrameStrobe_O[0] ;
 wire \Tile_X4Y0_FrameStrobe_O[10] ;
 wire \Tile_X4Y0_FrameStrobe_O[11] ;
 wire \Tile_X4Y0_FrameStrobe_O[12] ;
 wire \Tile_X4Y0_FrameStrobe_O[13] ;
 wire \Tile_X4Y0_FrameStrobe_O[14] ;
 wire \Tile_X4Y0_FrameStrobe_O[15] ;
 wire \Tile_X4Y0_FrameStrobe_O[16] ;
 wire \Tile_X4Y0_FrameStrobe_O[17] ;
 wire \Tile_X4Y0_FrameStrobe_O[18] ;
 wire \Tile_X4Y0_FrameStrobe_O[19] ;
 wire \Tile_X4Y0_FrameStrobe_O[1] ;
 wire \Tile_X4Y0_FrameStrobe_O[2] ;
 wire \Tile_X4Y0_FrameStrobe_O[3] ;
 wire \Tile_X4Y0_FrameStrobe_O[4] ;
 wire \Tile_X4Y0_FrameStrobe_O[5] ;
 wire \Tile_X4Y0_FrameStrobe_O[6] ;
 wire \Tile_X4Y0_FrameStrobe_O[7] ;
 wire \Tile_X4Y0_FrameStrobe_O[8] ;
 wire \Tile_X4Y0_FrameStrobe_O[9] ;
 wire \Tile_X4Y0_S1BEG[0] ;
 wire \Tile_X4Y0_S1BEG[1] ;
 wire \Tile_X4Y0_S1BEG[2] ;
 wire \Tile_X4Y0_S1BEG[3] ;
 wire \Tile_X4Y0_S2BEG[0] ;
 wire \Tile_X4Y0_S2BEG[1] ;
 wire \Tile_X4Y0_S2BEG[2] ;
 wire \Tile_X4Y0_S2BEG[3] ;
 wire \Tile_X4Y0_S2BEG[4] ;
 wire \Tile_X4Y0_S2BEG[5] ;
 wire \Tile_X4Y0_S2BEG[6] ;
 wire \Tile_X4Y0_S2BEG[7] ;
 wire \Tile_X4Y0_S2BEGb[0] ;
 wire \Tile_X4Y0_S2BEGb[1] ;
 wire \Tile_X4Y0_S2BEGb[2] ;
 wire \Tile_X4Y0_S2BEGb[3] ;
 wire \Tile_X4Y0_S2BEGb[4] ;
 wire \Tile_X4Y0_S2BEGb[5] ;
 wire \Tile_X4Y0_S2BEGb[6] ;
 wire \Tile_X4Y0_S2BEGb[7] ;
 wire \Tile_X4Y0_S4BEG[0] ;
 wire \Tile_X4Y0_S4BEG[10] ;
 wire \Tile_X4Y0_S4BEG[11] ;
 wire \Tile_X4Y0_S4BEG[12] ;
 wire \Tile_X4Y0_S4BEG[13] ;
 wire \Tile_X4Y0_S4BEG[14] ;
 wire \Tile_X4Y0_S4BEG[15] ;
 wire \Tile_X4Y0_S4BEG[1] ;
 wire \Tile_X4Y0_S4BEG[2] ;
 wire \Tile_X4Y0_S4BEG[3] ;
 wire \Tile_X4Y0_S4BEG[4] ;
 wire \Tile_X4Y0_S4BEG[5] ;
 wire \Tile_X4Y0_S4BEG[6] ;
 wire \Tile_X4Y0_S4BEG[7] ;
 wire \Tile_X4Y0_S4BEG[8] ;
 wire \Tile_X4Y0_S4BEG[9] ;
 wire \Tile_X4Y0_SS4BEG[0] ;
 wire \Tile_X4Y0_SS4BEG[10] ;
 wire \Tile_X4Y0_SS4BEG[11] ;
 wire \Tile_X4Y0_SS4BEG[12] ;
 wire \Tile_X4Y0_SS4BEG[13] ;
 wire \Tile_X4Y0_SS4BEG[14] ;
 wire \Tile_X4Y0_SS4BEG[15] ;
 wire \Tile_X4Y0_SS4BEG[1] ;
 wire \Tile_X4Y0_SS4BEG[2] ;
 wire \Tile_X4Y0_SS4BEG[3] ;
 wire \Tile_X4Y0_SS4BEG[4] ;
 wire \Tile_X4Y0_SS4BEG[5] ;
 wire \Tile_X4Y0_SS4BEG[6] ;
 wire \Tile_X4Y0_SS4BEG[7] ;
 wire \Tile_X4Y0_SS4BEG[8] ;
 wire \Tile_X4Y0_SS4BEG[9] ;
 wire Tile_X4Y0_UserCLKo;
 wire Tile_X4Y1_Co;
 wire \Tile_X4Y1_E1BEG[0] ;
 wire \Tile_X4Y1_E1BEG[1] ;
 wire \Tile_X4Y1_E1BEG[2] ;
 wire \Tile_X4Y1_E1BEG[3] ;
 wire \Tile_X4Y1_E2BEG[0] ;
 wire \Tile_X4Y1_E2BEG[1] ;
 wire \Tile_X4Y1_E2BEG[2] ;
 wire \Tile_X4Y1_E2BEG[3] ;
 wire \Tile_X4Y1_E2BEG[4] ;
 wire \Tile_X4Y1_E2BEG[5] ;
 wire \Tile_X4Y1_E2BEG[6] ;
 wire \Tile_X4Y1_E2BEG[7] ;
 wire \Tile_X4Y1_E2BEGb[0] ;
 wire \Tile_X4Y1_E2BEGb[1] ;
 wire \Tile_X4Y1_E2BEGb[2] ;
 wire \Tile_X4Y1_E2BEGb[3] ;
 wire \Tile_X4Y1_E2BEGb[4] ;
 wire \Tile_X4Y1_E2BEGb[5] ;
 wire \Tile_X4Y1_E2BEGb[6] ;
 wire \Tile_X4Y1_E2BEGb[7] ;
 wire \Tile_X4Y1_E6BEG[0] ;
 wire \Tile_X4Y1_E6BEG[10] ;
 wire \Tile_X4Y1_E6BEG[11] ;
 wire \Tile_X4Y1_E6BEG[1] ;
 wire \Tile_X4Y1_E6BEG[2] ;
 wire \Tile_X4Y1_E6BEG[3] ;
 wire \Tile_X4Y1_E6BEG[4] ;
 wire \Tile_X4Y1_E6BEG[5] ;
 wire \Tile_X4Y1_E6BEG[6] ;
 wire \Tile_X4Y1_E6BEG[7] ;
 wire \Tile_X4Y1_E6BEG[8] ;
 wire \Tile_X4Y1_E6BEG[9] ;
 wire \Tile_X4Y1_EE4BEG[0] ;
 wire \Tile_X4Y1_EE4BEG[10] ;
 wire \Tile_X4Y1_EE4BEG[11] ;
 wire \Tile_X4Y1_EE4BEG[12] ;
 wire \Tile_X4Y1_EE4BEG[13] ;
 wire \Tile_X4Y1_EE4BEG[14] ;
 wire \Tile_X4Y1_EE4BEG[15] ;
 wire \Tile_X4Y1_EE4BEG[1] ;
 wire \Tile_X4Y1_EE4BEG[2] ;
 wire \Tile_X4Y1_EE4BEG[3] ;
 wire \Tile_X4Y1_EE4BEG[4] ;
 wire \Tile_X4Y1_EE4BEG[5] ;
 wire \Tile_X4Y1_EE4BEG[6] ;
 wire \Tile_X4Y1_EE4BEG[7] ;
 wire \Tile_X4Y1_EE4BEG[8] ;
 wire \Tile_X4Y1_EE4BEG[9] ;
 wire \Tile_X4Y1_FrameData_O[0] ;
 wire \Tile_X4Y1_FrameData_O[10] ;
 wire \Tile_X4Y1_FrameData_O[11] ;
 wire \Tile_X4Y1_FrameData_O[12] ;
 wire \Tile_X4Y1_FrameData_O[13] ;
 wire \Tile_X4Y1_FrameData_O[14] ;
 wire \Tile_X4Y1_FrameData_O[15] ;
 wire \Tile_X4Y1_FrameData_O[16] ;
 wire \Tile_X4Y1_FrameData_O[17] ;
 wire \Tile_X4Y1_FrameData_O[18] ;
 wire \Tile_X4Y1_FrameData_O[19] ;
 wire \Tile_X4Y1_FrameData_O[1] ;
 wire \Tile_X4Y1_FrameData_O[20] ;
 wire \Tile_X4Y1_FrameData_O[21] ;
 wire \Tile_X4Y1_FrameData_O[22] ;
 wire \Tile_X4Y1_FrameData_O[23] ;
 wire \Tile_X4Y1_FrameData_O[24] ;
 wire \Tile_X4Y1_FrameData_O[25] ;
 wire \Tile_X4Y1_FrameData_O[26] ;
 wire \Tile_X4Y1_FrameData_O[27] ;
 wire \Tile_X4Y1_FrameData_O[28] ;
 wire \Tile_X4Y1_FrameData_O[29] ;
 wire \Tile_X4Y1_FrameData_O[2] ;
 wire \Tile_X4Y1_FrameData_O[30] ;
 wire \Tile_X4Y1_FrameData_O[31] ;
 wire \Tile_X4Y1_FrameData_O[3] ;
 wire \Tile_X4Y1_FrameData_O[4] ;
 wire \Tile_X4Y1_FrameData_O[5] ;
 wire \Tile_X4Y1_FrameData_O[6] ;
 wire \Tile_X4Y1_FrameData_O[7] ;
 wire \Tile_X4Y1_FrameData_O[8] ;
 wire \Tile_X4Y1_FrameData_O[9] ;
 wire \Tile_X4Y1_FrameStrobe_O[0] ;
 wire \Tile_X4Y1_FrameStrobe_O[10] ;
 wire \Tile_X4Y1_FrameStrobe_O[11] ;
 wire \Tile_X4Y1_FrameStrobe_O[12] ;
 wire \Tile_X4Y1_FrameStrobe_O[13] ;
 wire \Tile_X4Y1_FrameStrobe_O[14] ;
 wire \Tile_X4Y1_FrameStrobe_O[15] ;
 wire \Tile_X4Y1_FrameStrobe_O[16] ;
 wire \Tile_X4Y1_FrameStrobe_O[17] ;
 wire \Tile_X4Y1_FrameStrobe_O[18] ;
 wire \Tile_X4Y1_FrameStrobe_O[19] ;
 wire \Tile_X4Y1_FrameStrobe_O[1] ;
 wire \Tile_X4Y1_FrameStrobe_O[2] ;
 wire \Tile_X4Y1_FrameStrobe_O[3] ;
 wire \Tile_X4Y1_FrameStrobe_O[4] ;
 wire \Tile_X4Y1_FrameStrobe_O[5] ;
 wire \Tile_X4Y1_FrameStrobe_O[6] ;
 wire \Tile_X4Y1_FrameStrobe_O[7] ;
 wire \Tile_X4Y1_FrameStrobe_O[8] ;
 wire \Tile_X4Y1_FrameStrobe_O[9] ;
 wire \Tile_X4Y1_N1BEG[0] ;
 wire \Tile_X4Y1_N1BEG[1] ;
 wire \Tile_X4Y1_N1BEG[2] ;
 wire \Tile_X4Y1_N1BEG[3] ;
 wire \Tile_X4Y1_N2BEG[0] ;
 wire \Tile_X4Y1_N2BEG[1] ;
 wire \Tile_X4Y1_N2BEG[2] ;
 wire \Tile_X4Y1_N2BEG[3] ;
 wire \Tile_X4Y1_N2BEG[4] ;
 wire \Tile_X4Y1_N2BEG[5] ;
 wire \Tile_X4Y1_N2BEG[6] ;
 wire \Tile_X4Y1_N2BEG[7] ;
 wire \Tile_X4Y1_N2BEGb[0] ;
 wire \Tile_X4Y1_N2BEGb[1] ;
 wire \Tile_X4Y1_N2BEGb[2] ;
 wire \Tile_X4Y1_N2BEGb[3] ;
 wire \Tile_X4Y1_N2BEGb[4] ;
 wire \Tile_X4Y1_N2BEGb[5] ;
 wire \Tile_X4Y1_N2BEGb[6] ;
 wire \Tile_X4Y1_N2BEGb[7] ;
 wire \Tile_X4Y1_N4BEG[0] ;
 wire \Tile_X4Y1_N4BEG[10] ;
 wire \Tile_X4Y1_N4BEG[11] ;
 wire \Tile_X4Y1_N4BEG[12] ;
 wire \Tile_X4Y1_N4BEG[13] ;
 wire \Tile_X4Y1_N4BEG[14] ;
 wire \Tile_X4Y1_N4BEG[15] ;
 wire \Tile_X4Y1_N4BEG[1] ;
 wire \Tile_X4Y1_N4BEG[2] ;
 wire \Tile_X4Y1_N4BEG[3] ;
 wire \Tile_X4Y1_N4BEG[4] ;
 wire \Tile_X4Y1_N4BEG[5] ;
 wire \Tile_X4Y1_N4BEG[6] ;
 wire \Tile_X4Y1_N4BEG[7] ;
 wire \Tile_X4Y1_N4BEG[8] ;
 wire \Tile_X4Y1_N4BEG[9] ;
 wire \Tile_X4Y1_NN4BEG[0] ;
 wire \Tile_X4Y1_NN4BEG[10] ;
 wire \Tile_X4Y1_NN4BEG[11] ;
 wire \Tile_X4Y1_NN4BEG[12] ;
 wire \Tile_X4Y1_NN4BEG[13] ;
 wire \Tile_X4Y1_NN4BEG[14] ;
 wire \Tile_X4Y1_NN4BEG[15] ;
 wire \Tile_X4Y1_NN4BEG[1] ;
 wire \Tile_X4Y1_NN4BEG[2] ;
 wire \Tile_X4Y1_NN4BEG[3] ;
 wire \Tile_X4Y1_NN4BEG[4] ;
 wire \Tile_X4Y1_NN4BEG[5] ;
 wire \Tile_X4Y1_NN4BEG[6] ;
 wire \Tile_X4Y1_NN4BEG[7] ;
 wire \Tile_X4Y1_NN4BEG[8] ;
 wire \Tile_X4Y1_NN4BEG[9] ;
 wire \Tile_X4Y1_S1BEG[0] ;
 wire \Tile_X4Y1_S1BEG[1] ;
 wire \Tile_X4Y1_S1BEG[2] ;
 wire \Tile_X4Y1_S1BEG[3] ;
 wire \Tile_X4Y1_S2BEG[0] ;
 wire \Tile_X4Y1_S2BEG[1] ;
 wire \Tile_X4Y1_S2BEG[2] ;
 wire \Tile_X4Y1_S2BEG[3] ;
 wire \Tile_X4Y1_S2BEG[4] ;
 wire \Tile_X4Y1_S2BEG[5] ;
 wire \Tile_X4Y1_S2BEG[6] ;
 wire \Tile_X4Y1_S2BEG[7] ;
 wire \Tile_X4Y1_S2BEGb[0] ;
 wire \Tile_X4Y1_S2BEGb[1] ;
 wire \Tile_X4Y1_S2BEGb[2] ;
 wire \Tile_X4Y1_S2BEGb[3] ;
 wire \Tile_X4Y1_S2BEGb[4] ;
 wire \Tile_X4Y1_S2BEGb[5] ;
 wire \Tile_X4Y1_S2BEGb[6] ;
 wire \Tile_X4Y1_S2BEGb[7] ;
 wire \Tile_X4Y1_S4BEG[0] ;
 wire \Tile_X4Y1_S4BEG[10] ;
 wire \Tile_X4Y1_S4BEG[11] ;
 wire \Tile_X4Y1_S4BEG[12] ;
 wire \Tile_X4Y1_S4BEG[13] ;
 wire \Tile_X4Y1_S4BEG[14] ;
 wire \Tile_X4Y1_S4BEG[15] ;
 wire \Tile_X4Y1_S4BEG[1] ;
 wire \Tile_X4Y1_S4BEG[2] ;
 wire \Tile_X4Y1_S4BEG[3] ;
 wire \Tile_X4Y1_S4BEG[4] ;
 wire \Tile_X4Y1_S4BEG[5] ;
 wire \Tile_X4Y1_S4BEG[6] ;
 wire \Tile_X4Y1_S4BEG[7] ;
 wire \Tile_X4Y1_S4BEG[8] ;
 wire \Tile_X4Y1_S4BEG[9] ;
 wire \Tile_X4Y1_SS4BEG[0] ;
 wire \Tile_X4Y1_SS4BEG[10] ;
 wire \Tile_X4Y1_SS4BEG[11] ;
 wire \Tile_X4Y1_SS4BEG[12] ;
 wire \Tile_X4Y1_SS4BEG[13] ;
 wire \Tile_X4Y1_SS4BEG[14] ;
 wire \Tile_X4Y1_SS4BEG[15] ;
 wire \Tile_X4Y1_SS4BEG[1] ;
 wire \Tile_X4Y1_SS4BEG[2] ;
 wire \Tile_X4Y1_SS4BEG[3] ;
 wire \Tile_X4Y1_SS4BEG[4] ;
 wire \Tile_X4Y1_SS4BEG[5] ;
 wire \Tile_X4Y1_SS4BEG[6] ;
 wire \Tile_X4Y1_SS4BEG[7] ;
 wire \Tile_X4Y1_SS4BEG[8] ;
 wire \Tile_X4Y1_SS4BEG[9] ;
 wire Tile_X4Y1_UserCLKo;
 wire \Tile_X4Y1_W1BEG[0] ;
 wire \Tile_X4Y1_W1BEG[1] ;
 wire \Tile_X4Y1_W1BEG[2] ;
 wire \Tile_X4Y1_W1BEG[3] ;
 wire \Tile_X4Y1_W2BEG[0] ;
 wire \Tile_X4Y1_W2BEG[1] ;
 wire \Tile_X4Y1_W2BEG[2] ;
 wire \Tile_X4Y1_W2BEG[3] ;
 wire \Tile_X4Y1_W2BEG[4] ;
 wire \Tile_X4Y1_W2BEG[5] ;
 wire \Tile_X4Y1_W2BEG[6] ;
 wire \Tile_X4Y1_W2BEG[7] ;
 wire \Tile_X4Y1_W2BEGb[0] ;
 wire \Tile_X4Y1_W2BEGb[1] ;
 wire \Tile_X4Y1_W2BEGb[2] ;
 wire \Tile_X4Y1_W2BEGb[3] ;
 wire \Tile_X4Y1_W2BEGb[4] ;
 wire \Tile_X4Y1_W2BEGb[5] ;
 wire \Tile_X4Y1_W2BEGb[6] ;
 wire \Tile_X4Y1_W2BEGb[7] ;
 wire \Tile_X4Y1_W6BEG[0] ;
 wire \Tile_X4Y1_W6BEG[10] ;
 wire \Tile_X4Y1_W6BEG[11] ;
 wire \Tile_X4Y1_W6BEG[1] ;
 wire \Tile_X4Y1_W6BEG[2] ;
 wire \Tile_X4Y1_W6BEG[3] ;
 wire \Tile_X4Y1_W6BEG[4] ;
 wire \Tile_X4Y1_W6BEG[5] ;
 wire \Tile_X4Y1_W6BEG[6] ;
 wire \Tile_X4Y1_W6BEG[7] ;
 wire \Tile_X4Y1_W6BEG[8] ;
 wire \Tile_X4Y1_W6BEG[9] ;
 wire \Tile_X4Y1_WW4BEG[0] ;
 wire \Tile_X4Y1_WW4BEG[10] ;
 wire \Tile_X4Y1_WW4BEG[11] ;
 wire \Tile_X4Y1_WW4BEG[12] ;
 wire \Tile_X4Y1_WW4BEG[13] ;
 wire \Tile_X4Y1_WW4BEG[14] ;
 wire \Tile_X4Y1_WW4BEG[15] ;
 wire \Tile_X4Y1_WW4BEG[1] ;
 wire \Tile_X4Y1_WW4BEG[2] ;
 wire \Tile_X4Y1_WW4BEG[3] ;
 wire \Tile_X4Y1_WW4BEG[4] ;
 wire \Tile_X4Y1_WW4BEG[5] ;
 wire \Tile_X4Y1_WW4BEG[6] ;
 wire \Tile_X4Y1_WW4BEG[7] ;
 wire \Tile_X4Y1_WW4BEG[8] ;
 wire \Tile_X4Y1_WW4BEG[9] ;
 wire Tile_X4Y2_Co;
 wire \Tile_X4Y2_E1BEG[0] ;
 wire \Tile_X4Y2_E1BEG[1] ;
 wire \Tile_X4Y2_E1BEG[2] ;
 wire \Tile_X4Y2_E1BEG[3] ;
 wire \Tile_X4Y2_E2BEG[0] ;
 wire \Tile_X4Y2_E2BEG[1] ;
 wire \Tile_X4Y2_E2BEG[2] ;
 wire \Tile_X4Y2_E2BEG[3] ;
 wire \Tile_X4Y2_E2BEG[4] ;
 wire \Tile_X4Y2_E2BEG[5] ;
 wire \Tile_X4Y2_E2BEG[6] ;
 wire \Tile_X4Y2_E2BEG[7] ;
 wire \Tile_X4Y2_E2BEGb[0] ;
 wire \Tile_X4Y2_E2BEGb[1] ;
 wire \Tile_X4Y2_E2BEGb[2] ;
 wire \Tile_X4Y2_E2BEGb[3] ;
 wire \Tile_X4Y2_E2BEGb[4] ;
 wire \Tile_X4Y2_E2BEGb[5] ;
 wire \Tile_X4Y2_E2BEGb[6] ;
 wire \Tile_X4Y2_E2BEGb[7] ;
 wire \Tile_X4Y2_E6BEG[0] ;
 wire \Tile_X4Y2_E6BEG[10] ;
 wire \Tile_X4Y2_E6BEG[11] ;
 wire \Tile_X4Y2_E6BEG[1] ;
 wire \Tile_X4Y2_E6BEG[2] ;
 wire \Tile_X4Y2_E6BEG[3] ;
 wire \Tile_X4Y2_E6BEG[4] ;
 wire \Tile_X4Y2_E6BEG[5] ;
 wire \Tile_X4Y2_E6BEG[6] ;
 wire \Tile_X4Y2_E6BEG[7] ;
 wire \Tile_X4Y2_E6BEG[8] ;
 wire \Tile_X4Y2_E6BEG[9] ;
 wire \Tile_X4Y2_EE4BEG[0] ;
 wire \Tile_X4Y2_EE4BEG[10] ;
 wire \Tile_X4Y2_EE4BEG[11] ;
 wire \Tile_X4Y2_EE4BEG[12] ;
 wire \Tile_X4Y2_EE4BEG[13] ;
 wire \Tile_X4Y2_EE4BEG[14] ;
 wire \Tile_X4Y2_EE4BEG[15] ;
 wire \Tile_X4Y2_EE4BEG[1] ;
 wire \Tile_X4Y2_EE4BEG[2] ;
 wire \Tile_X4Y2_EE4BEG[3] ;
 wire \Tile_X4Y2_EE4BEG[4] ;
 wire \Tile_X4Y2_EE4BEG[5] ;
 wire \Tile_X4Y2_EE4BEG[6] ;
 wire \Tile_X4Y2_EE4BEG[7] ;
 wire \Tile_X4Y2_EE4BEG[8] ;
 wire \Tile_X4Y2_EE4BEG[9] ;
 wire \Tile_X4Y2_FrameData_O[0] ;
 wire \Tile_X4Y2_FrameData_O[10] ;
 wire \Tile_X4Y2_FrameData_O[11] ;
 wire \Tile_X4Y2_FrameData_O[12] ;
 wire \Tile_X4Y2_FrameData_O[13] ;
 wire \Tile_X4Y2_FrameData_O[14] ;
 wire \Tile_X4Y2_FrameData_O[15] ;
 wire \Tile_X4Y2_FrameData_O[16] ;
 wire \Tile_X4Y2_FrameData_O[17] ;
 wire \Tile_X4Y2_FrameData_O[18] ;
 wire \Tile_X4Y2_FrameData_O[19] ;
 wire \Tile_X4Y2_FrameData_O[1] ;
 wire \Tile_X4Y2_FrameData_O[20] ;
 wire \Tile_X4Y2_FrameData_O[21] ;
 wire \Tile_X4Y2_FrameData_O[22] ;
 wire \Tile_X4Y2_FrameData_O[23] ;
 wire \Tile_X4Y2_FrameData_O[24] ;
 wire \Tile_X4Y2_FrameData_O[25] ;
 wire \Tile_X4Y2_FrameData_O[26] ;
 wire \Tile_X4Y2_FrameData_O[27] ;
 wire \Tile_X4Y2_FrameData_O[28] ;
 wire \Tile_X4Y2_FrameData_O[29] ;
 wire \Tile_X4Y2_FrameData_O[2] ;
 wire \Tile_X4Y2_FrameData_O[30] ;
 wire \Tile_X4Y2_FrameData_O[31] ;
 wire \Tile_X4Y2_FrameData_O[3] ;
 wire \Tile_X4Y2_FrameData_O[4] ;
 wire \Tile_X4Y2_FrameData_O[5] ;
 wire \Tile_X4Y2_FrameData_O[6] ;
 wire \Tile_X4Y2_FrameData_O[7] ;
 wire \Tile_X4Y2_FrameData_O[8] ;
 wire \Tile_X4Y2_FrameData_O[9] ;
 wire \Tile_X4Y2_FrameStrobe_O[0] ;
 wire \Tile_X4Y2_FrameStrobe_O[10] ;
 wire \Tile_X4Y2_FrameStrobe_O[11] ;
 wire \Tile_X4Y2_FrameStrobe_O[12] ;
 wire \Tile_X4Y2_FrameStrobe_O[13] ;
 wire \Tile_X4Y2_FrameStrobe_O[14] ;
 wire \Tile_X4Y2_FrameStrobe_O[15] ;
 wire \Tile_X4Y2_FrameStrobe_O[16] ;
 wire \Tile_X4Y2_FrameStrobe_O[17] ;
 wire \Tile_X4Y2_FrameStrobe_O[18] ;
 wire \Tile_X4Y2_FrameStrobe_O[19] ;
 wire \Tile_X4Y2_FrameStrobe_O[1] ;
 wire \Tile_X4Y2_FrameStrobe_O[2] ;
 wire \Tile_X4Y2_FrameStrobe_O[3] ;
 wire \Tile_X4Y2_FrameStrobe_O[4] ;
 wire \Tile_X4Y2_FrameStrobe_O[5] ;
 wire \Tile_X4Y2_FrameStrobe_O[6] ;
 wire \Tile_X4Y2_FrameStrobe_O[7] ;
 wire \Tile_X4Y2_FrameStrobe_O[8] ;
 wire \Tile_X4Y2_FrameStrobe_O[9] ;
 wire \Tile_X4Y2_N1BEG[0] ;
 wire \Tile_X4Y2_N1BEG[1] ;
 wire \Tile_X4Y2_N1BEG[2] ;
 wire \Tile_X4Y2_N1BEG[3] ;
 wire \Tile_X4Y2_N2BEG[0] ;
 wire \Tile_X4Y2_N2BEG[1] ;
 wire \Tile_X4Y2_N2BEG[2] ;
 wire \Tile_X4Y2_N2BEG[3] ;
 wire \Tile_X4Y2_N2BEG[4] ;
 wire \Tile_X4Y2_N2BEG[5] ;
 wire \Tile_X4Y2_N2BEG[6] ;
 wire \Tile_X4Y2_N2BEG[7] ;
 wire \Tile_X4Y2_N2BEGb[0] ;
 wire \Tile_X4Y2_N2BEGb[1] ;
 wire \Tile_X4Y2_N2BEGb[2] ;
 wire \Tile_X4Y2_N2BEGb[3] ;
 wire \Tile_X4Y2_N2BEGb[4] ;
 wire \Tile_X4Y2_N2BEGb[5] ;
 wire \Tile_X4Y2_N2BEGb[6] ;
 wire \Tile_X4Y2_N2BEGb[7] ;
 wire \Tile_X4Y2_N4BEG[0] ;
 wire \Tile_X4Y2_N4BEG[10] ;
 wire \Tile_X4Y2_N4BEG[11] ;
 wire \Tile_X4Y2_N4BEG[12] ;
 wire \Tile_X4Y2_N4BEG[13] ;
 wire \Tile_X4Y2_N4BEG[14] ;
 wire \Tile_X4Y2_N4BEG[15] ;
 wire \Tile_X4Y2_N4BEG[1] ;
 wire \Tile_X4Y2_N4BEG[2] ;
 wire \Tile_X4Y2_N4BEG[3] ;
 wire \Tile_X4Y2_N4BEG[4] ;
 wire \Tile_X4Y2_N4BEG[5] ;
 wire \Tile_X4Y2_N4BEG[6] ;
 wire \Tile_X4Y2_N4BEG[7] ;
 wire \Tile_X4Y2_N4BEG[8] ;
 wire \Tile_X4Y2_N4BEG[9] ;
 wire \Tile_X4Y2_NN4BEG[0] ;
 wire \Tile_X4Y2_NN4BEG[10] ;
 wire \Tile_X4Y2_NN4BEG[11] ;
 wire \Tile_X4Y2_NN4BEG[12] ;
 wire \Tile_X4Y2_NN4BEG[13] ;
 wire \Tile_X4Y2_NN4BEG[14] ;
 wire \Tile_X4Y2_NN4BEG[15] ;
 wire \Tile_X4Y2_NN4BEG[1] ;
 wire \Tile_X4Y2_NN4BEG[2] ;
 wire \Tile_X4Y2_NN4BEG[3] ;
 wire \Tile_X4Y2_NN4BEG[4] ;
 wire \Tile_X4Y2_NN4BEG[5] ;
 wire \Tile_X4Y2_NN4BEG[6] ;
 wire \Tile_X4Y2_NN4BEG[7] ;
 wire \Tile_X4Y2_NN4BEG[8] ;
 wire \Tile_X4Y2_NN4BEG[9] ;
 wire \Tile_X4Y2_S1BEG[0] ;
 wire \Tile_X4Y2_S1BEG[1] ;
 wire \Tile_X4Y2_S1BEG[2] ;
 wire \Tile_X4Y2_S1BEG[3] ;
 wire \Tile_X4Y2_S2BEG[0] ;
 wire \Tile_X4Y2_S2BEG[1] ;
 wire \Tile_X4Y2_S2BEG[2] ;
 wire \Tile_X4Y2_S2BEG[3] ;
 wire \Tile_X4Y2_S2BEG[4] ;
 wire \Tile_X4Y2_S2BEG[5] ;
 wire \Tile_X4Y2_S2BEG[6] ;
 wire \Tile_X4Y2_S2BEG[7] ;
 wire \Tile_X4Y2_S2BEGb[0] ;
 wire \Tile_X4Y2_S2BEGb[1] ;
 wire \Tile_X4Y2_S2BEGb[2] ;
 wire \Tile_X4Y2_S2BEGb[3] ;
 wire \Tile_X4Y2_S2BEGb[4] ;
 wire \Tile_X4Y2_S2BEGb[5] ;
 wire \Tile_X4Y2_S2BEGb[6] ;
 wire \Tile_X4Y2_S2BEGb[7] ;
 wire \Tile_X4Y2_S4BEG[0] ;
 wire \Tile_X4Y2_S4BEG[10] ;
 wire \Tile_X4Y2_S4BEG[11] ;
 wire \Tile_X4Y2_S4BEG[12] ;
 wire \Tile_X4Y2_S4BEG[13] ;
 wire \Tile_X4Y2_S4BEG[14] ;
 wire \Tile_X4Y2_S4BEG[15] ;
 wire \Tile_X4Y2_S4BEG[1] ;
 wire \Tile_X4Y2_S4BEG[2] ;
 wire \Tile_X4Y2_S4BEG[3] ;
 wire \Tile_X4Y2_S4BEG[4] ;
 wire \Tile_X4Y2_S4BEG[5] ;
 wire \Tile_X4Y2_S4BEG[6] ;
 wire \Tile_X4Y2_S4BEG[7] ;
 wire \Tile_X4Y2_S4BEG[8] ;
 wire \Tile_X4Y2_S4BEG[9] ;
 wire \Tile_X4Y2_SS4BEG[0] ;
 wire \Tile_X4Y2_SS4BEG[10] ;
 wire \Tile_X4Y2_SS4BEG[11] ;
 wire \Tile_X4Y2_SS4BEG[12] ;
 wire \Tile_X4Y2_SS4BEG[13] ;
 wire \Tile_X4Y2_SS4BEG[14] ;
 wire \Tile_X4Y2_SS4BEG[15] ;
 wire \Tile_X4Y2_SS4BEG[1] ;
 wire \Tile_X4Y2_SS4BEG[2] ;
 wire \Tile_X4Y2_SS4BEG[3] ;
 wire \Tile_X4Y2_SS4BEG[4] ;
 wire \Tile_X4Y2_SS4BEG[5] ;
 wire \Tile_X4Y2_SS4BEG[6] ;
 wire \Tile_X4Y2_SS4BEG[7] ;
 wire \Tile_X4Y2_SS4BEG[8] ;
 wire \Tile_X4Y2_SS4BEG[9] ;
 wire Tile_X4Y2_UserCLKo;
 wire \Tile_X4Y2_W1BEG[0] ;
 wire \Tile_X4Y2_W1BEG[1] ;
 wire \Tile_X4Y2_W1BEG[2] ;
 wire \Tile_X4Y2_W1BEG[3] ;
 wire \Tile_X4Y2_W2BEG[0] ;
 wire \Tile_X4Y2_W2BEG[1] ;
 wire \Tile_X4Y2_W2BEG[2] ;
 wire \Tile_X4Y2_W2BEG[3] ;
 wire \Tile_X4Y2_W2BEG[4] ;
 wire \Tile_X4Y2_W2BEG[5] ;
 wire \Tile_X4Y2_W2BEG[6] ;
 wire \Tile_X4Y2_W2BEG[7] ;
 wire \Tile_X4Y2_W2BEGb[0] ;
 wire \Tile_X4Y2_W2BEGb[1] ;
 wire \Tile_X4Y2_W2BEGb[2] ;
 wire \Tile_X4Y2_W2BEGb[3] ;
 wire \Tile_X4Y2_W2BEGb[4] ;
 wire \Tile_X4Y2_W2BEGb[5] ;
 wire \Tile_X4Y2_W2BEGb[6] ;
 wire \Tile_X4Y2_W2BEGb[7] ;
 wire \Tile_X4Y2_W6BEG[0] ;
 wire \Tile_X4Y2_W6BEG[10] ;
 wire \Tile_X4Y2_W6BEG[11] ;
 wire \Tile_X4Y2_W6BEG[1] ;
 wire \Tile_X4Y2_W6BEG[2] ;
 wire \Tile_X4Y2_W6BEG[3] ;
 wire \Tile_X4Y2_W6BEG[4] ;
 wire \Tile_X4Y2_W6BEG[5] ;
 wire \Tile_X4Y2_W6BEG[6] ;
 wire \Tile_X4Y2_W6BEG[7] ;
 wire \Tile_X4Y2_W6BEG[8] ;
 wire \Tile_X4Y2_W6BEG[9] ;
 wire \Tile_X4Y2_WW4BEG[0] ;
 wire \Tile_X4Y2_WW4BEG[10] ;
 wire \Tile_X4Y2_WW4BEG[11] ;
 wire \Tile_X4Y2_WW4BEG[12] ;
 wire \Tile_X4Y2_WW4BEG[13] ;
 wire \Tile_X4Y2_WW4BEG[14] ;
 wire \Tile_X4Y2_WW4BEG[15] ;
 wire \Tile_X4Y2_WW4BEG[1] ;
 wire \Tile_X4Y2_WW4BEG[2] ;
 wire \Tile_X4Y2_WW4BEG[3] ;
 wire \Tile_X4Y2_WW4BEG[4] ;
 wire \Tile_X4Y2_WW4BEG[5] ;
 wire \Tile_X4Y2_WW4BEG[6] ;
 wire \Tile_X4Y2_WW4BEG[7] ;
 wire \Tile_X4Y2_WW4BEG[8] ;
 wire \Tile_X4Y2_WW4BEG[9] ;
 wire Tile_X4Y3_Co;
 wire \Tile_X4Y3_E1BEG[0] ;
 wire \Tile_X4Y3_E1BEG[1] ;
 wire \Tile_X4Y3_E1BEG[2] ;
 wire \Tile_X4Y3_E1BEG[3] ;
 wire \Tile_X4Y3_E2BEG[0] ;
 wire \Tile_X4Y3_E2BEG[1] ;
 wire \Tile_X4Y3_E2BEG[2] ;
 wire \Tile_X4Y3_E2BEG[3] ;
 wire \Tile_X4Y3_E2BEG[4] ;
 wire \Tile_X4Y3_E2BEG[5] ;
 wire \Tile_X4Y3_E2BEG[6] ;
 wire \Tile_X4Y3_E2BEG[7] ;
 wire \Tile_X4Y3_E2BEGb[0] ;
 wire \Tile_X4Y3_E2BEGb[1] ;
 wire \Tile_X4Y3_E2BEGb[2] ;
 wire \Tile_X4Y3_E2BEGb[3] ;
 wire \Tile_X4Y3_E2BEGb[4] ;
 wire \Tile_X4Y3_E2BEGb[5] ;
 wire \Tile_X4Y3_E2BEGb[6] ;
 wire \Tile_X4Y3_E2BEGb[7] ;
 wire \Tile_X4Y3_E6BEG[0] ;
 wire \Tile_X4Y3_E6BEG[10] ;
 wire \Tile_X4Y3_E6BEG[11] ;
 wire \Tile_X4Y3_E6BEG[1] ;
 wire \Tile_X4Y3_E6BEG[2] ;
 wire \Tile_X4Y3_E6BEG[3] ;
 wire \Tile_X4Y3_E6BEG[4] ;
 wire \Tile_X4Y3_E6BEG[5] ;
 wire \Tile_X4Y3_E6BEG[6] ;
 wire \Tile_X4Y3_E6BEG[7] ;
 wire \Tile_X4Y3_E6BEG[8] ;
 wire \Tile_X4Y3_E6BEG[9] ;
 wire \Tile_X4Y3_EE4BEG[0] ;
 wire \Tile_X4Y3_EE4BEG[10] ;
 wire \Tile_X4Y3_EE4BEG[11] ;
 wire \Tile_X4Y3_EE4BEG[12] ;
 wire \Tile_X4Y3_EE4BEG[13] ;
 wire \Tile_X4Y3_EE4BEG[14] ;
 wire \Tile_X4Y3_EE4BEG[15] ;
 wire \Tile_X4Y3_EE4BEG[1] ;
 wire \Tile_X4Y3_EE4BEG[2] ;
 wire \Tile_X4Y3_EE4BEG[3] ;
 wire \Tile_X4Y3_EE4BEG[4] ;
 wire \Tile_X4Y3_EE4BEG[5] ;
 wire \Tile_X4Y3_EE4BEG[6] ;
 wire \Tile_X4Y3_EE4BEG[7] ;
 wire \Tile_X4Y3_EE4BEG[8] ;
 wire \Tile_X4Y3_EE4BEG[9] ;
 wire \Tile_X4Y3_FrameData_O[0] ;
 wire \Tile_X4Y3_FrameData_O[10] ;
 wire \Tile_X4Y3_FrameData_O[11] ;
 wire \Tile_X4Y3_FrameData_O[12] ;
 wire \Tile_X4Y3_FrameData_O[13] ;
 wire \Tile_X4Y3_FrameData_O[14] ;
 wire \Tile_X4Y3_FrameData_O[15] ;
 wire \Tile_X4Y3_FrameData_O[16] ;
 wire \Tile_X4Y3_FrameData_O[17] ;
 wire \Tile_X4Y3_FrameData_O[18] ;
 wire \Tile_X4Y3_FrameData_O[19] ;
 wire \Tile_X4Y3_FrameData_O[1] ;
 wire \Tile_X4Y3_FrameData_O[20] ;
 wire \Tile_X4Y3_FrameData_O[21] ;
 wire \Tile_X4Y3_FrameData_O[22] ;
 wire \Tile_X4Y3_FrameData_O[23] ;
 wire \Tile_X4Y3_FrameData_O[24] ;
 wire \Tile_X4Y3_FrameData_O[25] ;
 wire \Tile_X4Y3_FrameData_O[26] ;
 wire \Tile_X4Y3_FrameData_O[27] ;
 wire \Tile_X4Y3_FrameData_O[28] ;
 wire \Tile_X4Y3_FrameData_O[29] ;
 wire \Tile_X4Y3_FrameData_O[2] ;
 wire \Tile_X4Y3_FrameData_O[30] ;
 wire \Tile_X4Y3_FrameData_O[31] ;
 wire \Tile_X4Y3_FrameData_O[3] ;
 wire \Tile_X4Y3_FrameData_O[4] ;
 wire \Tile_X4Y3_FrameData_O[5] ;
 wire \Tile_X4Y3_FrameData_O[6] ;
 wire \Tile_X4Y3_FrameData_O[7] ;
 wire \Tile_X4Y3_FrameData_O[8] ;
 wire \Tile_X4Y3_FrameData_O[9] ;
 wire \Tile_X4Y3_FrameStrobe_O[0] ;
 wire \Tile_X4Y3_FrameStrobe_O[10] ;
 wire \Tile_X4Y3_FrameStrobe_O[11] ;
 wire \Tile_X4Y3_FrameStrobe_O[12] ;
 wire \Tile_X4Y3_FrameStrobe_O[13] ;
 wire \Tile_X4Y3_FrameStrobe_O[14] ;
 wire \Tile_X4Y3_FrameStrobe_O[15] ;
 wire \Tile_X4Y3_FrameStrobe_O[16] ;
 wire \Tile_X4Y3_FrameStrobe_O[17] ;
 wire \Tile_X4Y3_FrameStrobe_O[18] ;
 wire \Tile_X4Y3_FrameStrobe_O[19] ;
 wire \Tile_X4Y3_FrameStrobe_O[1] ;
 wire \Tile_X4Y3_FrameStrobe_O[2] ;
 wire \Tile_X4Y3_FrameStrobe_O[3] ;
 wire \Tile_X4Y3_FrameStrobe_O[4] ;
 wire \Tile_X4Y3_FrameStrobe_O[5] ;
 wire \Tile_X4Y3_FrameStrobe_O[6] ;
 wire \Tile_X4Y3_FrameStrobe_O[7] ;
 wire \Tile_X4Y3_FrameStrobe_O[8] ;
 wire \Tile_X4Y3_FrameStrobe_O[9] ;
 wire \Tile_X4Y3_N1BEG[0] ;
 wire \Tile_X4Y3_N1BEG[1] ;
 wire \Tile_X4Y3_N1BEG[2] ;
 wire \Tile_X4Y3_N1BEG[3] ;
 wire \Tile_X4Y3_N2BEG[0] ;
 wire \Tile_X4Y3_N2BEG[1] ;
 wire \Tile_X4Y3_N2BEG[2] ;
 wire \Tile_X4Y3_N2BEG[3] ;
 wire \Tile_X4Y3_N2BEG[4] ;
 wire \Tile_X4Y3_N2BEG[5] ;
 wire \Tile_X4Y3_N2BEG[6] ;
 wire \Tile_X4Y3_N2BEG[7] ;
 wire \Tile_X4Y3_N2BEGb[0] ;
 wire \Tile_X4Y3_N2BEGb[1] ;
 wire \Tile_X4Y3_N2BEGb[2] ;
 wire \Tile_X4Y3_N2BEGb[3] ;
 wire \Tile_X4Y3_N2BEGb[4] ;
 wire \Tile_X4Y3_N2BEGb[5] ;
 wire \Tile_X4Y3_N2BEGb[6] ;
 wire \Tile_X4Y3_N2BEGb[7] ;
 wire \Tile_X4Y3_N4BEG[0] ;
 wire \Tile_X4Y3_N4BEG[10] ;
 wire \Tile_X4Y3_N4BEG[11] ;
 wire \Tile_X4Y3_N4BEG[12] ;
 wire \Tile_X4Y3_N4BEG[13] ;
 wire \Tile_X4Y3_N4BEG[14] ;
 wire \Tile_X4Y3_N4BEG[15] ;
 wire \Tile_X4Y3_N4BEG[1] ;
 wire \Tile_X4Y3_N4BEG[2] ;
 wire \Tile_X4Y3_N4BEG[3] ;
 wire \Tile_X4Y3_N4BEG[4] ;
 wire \Tile_X4Y3_N4BEG[5] ;
 wire \Tile_X4Y3_N4BEG[6] ;
 wire \Tile_X4Y3_N4BEG[7] ;
 wire \Tile_X4Y3_N4BEG[8] ;
 wire \Tile_X4Y3_N4BEG[9] ;
 wire \Tile_X4Y3_NN4BEG[0] ;
 wire \Tile_X4Y3_NN4BEG[10] ;
 wire \Tile_X4Y3_NN4BEG[11] ;
 wire \Tile_X4Y3_NN4BEG[12] ;
 wire \Tile_X4Y3_NN4BEG[13] ;
 wire \Tile_X4Y3_NN4BEG[14] ;
 wire \Tile_X4Y3_NN4BEG[15] ;
 wire \Tile_X4Y3_NN4BEG[1] ;
 wire \Tile_X4Y3_NN4BEG[2] ;
 wire \Tile_X4Y3_NN4BEG[3] ;
 wire \Tile_X4Y3_NN4BEG[4] ;
 wire \Tile_X4Y3_NN4BEG[5] ;
 wire \Tile_X4Y3_NN4BEG[6] ;
 wire \Tile_X4Y3_NN4BEG[7] ;
 wire \Tile_X4Y3_NN4BEG[8] ;
 wire \Tile_X4Y3_NN4BEG[9] ;
 wire \Tile_X4Y3_S1BEG[0] ;
 wire \Tile_X4Y3_S1BEG[1] ;
 wire \Tile_X4Y3_S1BEG[2] ;
 wire \Tile_X4Y3_S1BEG[3] ;
 wire \Tile_X4Y3_S2BEG[0] ;
 wire \Tile_X4Y3_S2BEG[1] ;
 wire \Tile_X4Y3_S2BEG[2] ;
 wire \Tile_X4Y3_S2BEG[3] ;
 wire \Tile_X4Y3_S2BEG[4] ;
 wire \Tile_X4Y3_S2BEG[5] ;
 wire \Tile_X4Y3_S2BEG[6] ;
 wire \Tile_X4Y3_S2BEG[7] ;
 wire \Tile_X4Y3_S2BEGb[0] ;
 wire \Tile_X4Y3_S2BEGb[1] ;
 wire \Tile_X4Y3_S2BEGb[2] ;
 wire \Tile_X4Y3_S2BEGb[3] ;
 wire \Tile_X4Y3_S2BEGb[4] ;
 wire \Tile_X4Y3_S2BEGb[5] ;
 wire \Tile_X4Y3_S2BEGb[6] ;
 wire \Tile_X4Y3_S2BEGb[7] ;
 wire \Tile_X4Y3_S4BEG[0] ;
 wire \Tile_X4Y3_S4BEG[10] ;
 wire \Tile_X4Y3_S4BEG[11] ;
 wire \Tile_X4Y3_S4BEG[12] ;
 wire \Tile_X4Y3_S4BEG[13] ;
 wire \Tile_X4Y3_S4BEG[14] ;
 wire \Tile_X4Y3_S4BEG[15] ;
 wire \Tile_X4Y3_S4BEG[1] ;
 wire \Tile_X4Y3_S4BEG[2] ;
 wire \Tile_X4Y3_S4BEG[3] ;
 wire \Tile_X4Y3_S4BEG[4] ;
 wire \Tile_X4Y3_S4BEG[5] ;
 wire \Tile_X4Y3_S4BEG[6] ;
 wire \Tile_X4Y3_S4BEG[7] ;
 wire \Tile_X4Y3_S4BEG[8] ;
 wire \Tile_X4Y3_S4BEG[9] ;
 wire \Tile_X4Y3_SS4BEG[0] ;
 wire \Tile_X4Y3_SS4BEG[10] ;
 wire \Tile_X4Y3_SS4BEG[11] ;
 wire \Tile_X4Y3_SS4BEG[12] ;
 wire \Tile_X4Y3_SS4BEG[13] ;
 wire \Tile_X4Y3_SS4BEG[14] ;
 wire \Tile_X4Y3_SS4BEG[15] ;
 wire \Tile_X4Y3_SS4BEG[1] ;
 wire \Tile_X4Y3_SS4BEG[2] ;
 wire \Tile_X4Y3_SS4BEG[3] ;
 wire \Tile_X4Y3_SS4BEG[4] ;
 wire \Tile_X4Y3_SS4BEG[5] ;
 wire \Tile_X4Y3_SS4BEG[6] ;
 wire \Tile_X4Y3_SS4BEG[7] ;
 wire \Tile_X4Y3_SS4BEG[8] ;
 wire \Tile_X4Y3_SS4BEG[9] ;
 wire Tile_X4Y3_UserCLKo;
 wire \Tile_X4Y3_W1BEG[0] ;
 wire \Tile_X4Y3_W1BEG[1] ;
 wire \Tile_X4Y3_W1BEG[2] ;
 wire \Tile_X4Y3_W1BEG[3] ;
 wire \Tile_X4Y3_W2BEG[0] ;
 wire \Tile_X4Y3_W2BEG[1] ;
 wire \Tile_X4Y3_W2BEG[2] ;
 wire \Tile_X4Y3_W2BEG[3] ;
 wire \Tile_X4Y3_W2BEG[4] ;
 wire \Tile_X4Y3_W2BEG[5] ;
 wire \Tile_X4Y3_W2BEG[6] ;
 wire \Tile_X4Y3_W2BEG[7] ;
 wire \Tile_X4Y3_W2BEGb[0] ;
 wire \Tile_X4Y3_W2BEGb[1] ;
 wire \Tile_X4Y3_W2BEGb[2] ;
 wire \Tile_X4Y3_W2BEGb[3] ;
 wire \Tile_X4Y3_W2BEGb[4] ;
 wire \Tile_X4Y3_W2BEGb[5] ;
 wire \Tile_X4Y3_W2BEGb[6] ;
 wire \Tile_X4Y3_W2BEGb[7] ;
 wire \Tile_X4Y3_W6BEG[0] ;
 wire \Tile_X4Y3_W6BEG[10] ;
 wire \Tile_X4Y3_W6BEG[11] ;
 wire \Tile_X4Y3_W6BEG[1] ;
 wire \Tile_X4Y3_W6BEG[2] ;
 wire \Tile_X4Y3_W6BEG[3] ;
 wire \Tile_X4Y3_W6BEG[4] ;
 wire \Tile_X4Y3_W6BEG[5] ;
 wire \Tile_X4Y3_W6BEG[6] ;
 wire \Tile_X4Y3_W6BEG[7] ;
 wire \Tile_X4Y3_W6BEG[8] ;
 wire \Tile_X4Y3_W6BEG[9] ;
 wire \Tile_X4Y3_WW4BEG[0] ;
 wire \Tile_X4Y3_WW4BEG[10] ;
 wire \Tile_X4Y3_WW4BEG[11] ;
 wire \Tile_X4Y3_WW4BEG[12] ;
 wire \Tile_X4Y3_WW4BEG[13] ;
 wire \Tile_X4Y3_WW4BEG[14] ;
 wire \Tile_X4Y3_WW4BEG[15] ;
 wire \Tile_X4Y3_WW4BEG[1] ;
 wire \Tile_X4Y3_WW4BEG[2] ;
 wire \Tile_X4Y3_WW4BEG[3] ;
 wire \Tile_X4Y3_WW4BEG[4] ;
 wire \Tile_X4Y3_WW4BEG[5] ;
 wire \Tile_X4Y3_WW4BEG[6] ;
 wire \Tile_X4Y3_WW4BEG[7] ;
 wire \Tile_X4Y3_WW4BEG[8] ;
 wire \Tile_X4Y3_WW4BEG[9] ;
 wire Tile_X4Y4_Co;
 wire \Tile_X4Y4_E1BEG[0] ;
 wire \Tile_X4Y4_E1BEG[1] ;
 wire \Tile_X4Y4_E1BEG[2] ;
 wire \Tile_X4Y4_E1BEG[3] ;
 wire \Tile_X4Y4_E2BEG[0] ;
 wire \Tile_X4Y4_E2BEG[1] ;
 wire \Tile_X4Y4_E2BEG[2] ;
 wire \Tile_X4Y4_E2BEG[3] ;
 wire \Tile_X4Y4_E2BEG[4] ;
 wire \Tile_X4Y4_E2BEG[5] ;
 wire \Tile_X4Y4_E2BEG[6] ;
 wire \Tile_X4Y4_E2BEG[7] ;
 wire \Tile_X4Y4_E2BEGb[0] ;
 wire \Tile_X4Y4_E2BEGb[1] ;
 wire \Tile_X4Y4_E2BEGb[2] ;
 wire \Tile_X4Y4_E2BEGb[3] ;
 wire \Tile_X4Y4_E2BEGb[4] ;
 wire \Tile_X4Y4_E2BEGb[5] ;
 wire \Tile_X4Y4_E2BEGb[6] ;
 wire \Tile_X4Y4_E2BEGb[7] ;
 wire \Tile_X4Y4_E6BEG[0] ;
 wire \Tile_X4Y4_E6BEG[10] ;
 wire \Tile_X4Y4_E6BEG[11] ;
 wire \Tile_X4Y4_E6BEG[1] ;
 wire \Tile_X4Y4_E6BEG[2] ;
 wire \Tile_X4Y4_E6BEG[3] ;
 wire \Tile_X4Y4_E6BEG[4] ;
 wire \Tile_X4Y4_E6BEG[5] ;
 wire \Tile_X4Y4_E6BEG[6] ;
 wire \Tile_X4Y4_E6BEG[7] ;
 wire \Tile_X4Y4_E6BEG[8] ;
 wire \Tile_X4Y4_E6BEG[9] ;
 wire \Tile_X4Y4_EE4BEG[0] ;
 wire \Tile_X4Y4_EE4BEG[10] ;
 wire \Tile_X4Y4_EE4BEG[11] ;
 wire \Tile_X4Y4_EE4BEG[12] ;
 wire \Tile_X4Y4_EE4BEG[13] ;
 wire \Tile_X4Y4_EE4BEG[14] ;
 wire \Tile_X4Y4_EE4BEG[15] ;
 wire \Tile_X4Y4_EE4BEG[1] ;
 wire \Tile_X4Y4_EE4BEG[2] ;
 wire \Tile_X4Y4_EE4BEG[3] ;
 wire \Tile_X4Y4_EE4BEG[4] ;
 wire \Tile_X4Y4_EE4BEG[5] ;
 wire \Tile_X4Y4_EE4BEG[6] ;
 wire \Tile_X4Y4_EE4BEG[7] ;
 wire \Tile_X4Y4_EE4BEG[8] ;
 wire \Tile_X4Y4_EE4BEG[9] ;
 wire \Tile_X4Y4_FrameData_O[0] ;
 wire \Tile_X4Y4_FrameData_O[10] ;
 wire \Tile_X4Y4_FrameData_O[11] ;
 wire \Tile_X4Y4_FrameData_O[12] ;
 wire \Tile_X4Y4_FrameData_O[13] ;
 wire \Tile_X4Y4_FrameData_O[14] ;
 wire \Tile_X4Y4_FrameData_O[15] ;
 wire \Tile_X4Y4_FrameData_O[16] ;
 wire \Tile_X4Y4_FrameData_O[17] ;
 wire \Tile_X4Y4_FrameData_O[18] ;
 wire \Tile_X4Y4_FrameData_O[19] ;
 wire \Tile_X4Y4_FrameData_O[1] ;
 wire \Tile_X4Y4_FrameData_O[20] ;
 wire \Tile_X4Y4_FrameData_O[21] ;
 wire \Tile_X4Y4_FrameData_O[22] ;
 wire \Tile_X4Y4_FrameData_O[23] ;
 wire \Tile_X4Y4_FrameData_O[24] ;
 wire \Tile_X4Y4_FrameData_O[25] ;
 wire \Tile_X4Y4_FrameData_O[26] ;
 wire \Tile_X4Y4_FrameData_O[27] ;
 wire \Tile_X4Y4_FrameData_O[28] ;
 wire \Tile_X4Y4_FrameData_O[29] ;
 wire \Tile_X4Y4_FrameData_O[2] ;
 wire \Tile_X4Y4_FrameData_O[30] ;
 wire \Tile_X4Y4_FrameData_O[31] ;
 wire \Tile_X4Y4_FrameData_O[3] ;
 wire \Tile_X4Y4_FrameData_O[4] ;
 wire \Tile_X4Y4_FrameData_O[5] ;
 wire \Tile_X4Y4_FrameData_O[6] ;
 wire \Tile_X4Y4_FrameData_O[7] ;
 wire \Tile_X4Y4_FrameData_O[8] ;
 wire \Tile_X4Y4_FrameData_O[9] ;
 wire \Tile_X4Y4_FrameStrobe_O[0] ;
 wire \Tile_X4Y4_FrameStrobe_O[10] ;
 wire \Tile_X4Y4_FrameStrobe_O[11] ;
 wire \Tile_X4Y4_FrameStrobe_O[12] ;
 wire \Tile_X4Y4_FrameStrobe_O[13] ;
 wire \Tile_X4Y4_FrameStrobe_O[14] ;
 wire \Tile_X4Y4_FrameStrobe_O[15] ;
 wire \Tile_X4Y4_FrameStrobe_O[16] ;
 wire \Tile_X4Y4_FrameStrobe_O[17] ;
 wire \Tile_X4Y4_FrameStrobe_O[18] ;
 wire \Tile_X4Y4_FrameStrobe_O[19] ;
 wire \Tile_X4Y4_FrameStrobe_O[1] ;
 wire \Tile_X4Y4_FrameStrobe_O[2] ;
 wire \Tile_X4Y4_FrameStrobe_O[3] ;
 wire \Tile_X4Y4_FrameStrobe_O[4] ;
 wire \Tile_X4Y4_FrameStrobe_O[5] ;
 wire \Tile_X4Y4_FrameStrobe_O[6] ;
 wire \Tile_X4Y4_FrameStrobe_O[7] ;
 wire \Tile_X4Y4_FrameStrobe_O[8] ;
 wire \Tile_X4Y4_FrameStrobe_O[9] ;
 wire \Tile_X4Y4_N1BEG[0] ;
 wire \Tile_X4Y4_N1BEG[1] ;
 wire \Tile_X4Y4_N1BEG[2] ;
 wire \Tile_X4Y4_N1BEG[3] ;
 wire \Tile_X4Y4_N2BEG[0] ;
 wire \Tile_X4Y4_N2BEG[1] ;
 wire \Tile_X4Y4_N2BEG[2] ;
 wire \Tile_X4Y4_N2BEG[3] ;
 wire \Tile_X4Y4_N2BEG[4] ;
 wire \Tile_X4Y4_N2BEG[5] ;
 wire \Tile_X4Y4_N2BEG[6] ;
 wire \Tile_X4Y4_N2BEG[7] ;
 wire \Tile_X4Y4_N2BEGb[0] ;
 wire \Tile_X4Y4_N2BEGb[1] ;
 wire \Tile_X4Y4_N2BEGb[2] ;
 wire \Tile_X4Y4_N2BEGb[3] ;
 wire \Tile_X4Y4_N2BEGb[4] ;
 wire \Tile_X4Y4_N2BEGb[5] ;
 wire \Tile_X4Y4_N2BEGb[6] ;
 wire \Tile_X4Y4_N2BEGb[7] ;
 wire \Tile_X4Y4_N4BEG[0] ;
 wire \Tile_X4Y4_N4BEG[10] ;
 wire \Tile_X4Y4_N4BEG[11] ;
 wire \Tile_X4Y4_N4BEG[12] ;
 wire \Tile_X4Y4_N4BEG[13] ;
 wire \Tile_X4Y4_N4BEG[14] ;
 wire \Tile_X4Y4_N4BEG[15] ;
 wire \Tile_X4Y4_N4BEG[1] ;
 wire \Tile_X4Y4_N4BEG[2] ;
 wire \Tile_X4Y4_N4BEG[3] ;
 wire \Tile_X4Y4_N4BEG[4] ;
 wire \Tile_X4Y4_N4BEG[5] ;
 wire \Tile_X4Y4_N4BEG[6] ;
 wire \Tile_X4Y4_N4BEG[7] ;
 wire \Tile_X4Y4_N4BEG[8] ;
 wire \Tile_X4Y4_N4BEG[9] ;
 wire \Tile_X4Y4_NN4BEG[0] ;
 wire \Tile_X4Y4_NN4BEG[10] ;
 wire \Tile_X4Y4_NN4BEG[11] ;
 wire \Tile_X4Y4_NN4BEG[12] ;
 wire \Tile_X4Y4_NN4BEG[13] ;
 wire \Tile_X4Y4_NN4BEG[14] ;
 wire \Tile_X4Y4_NN4BEG[15] ;
 wire \Tile_X4Y4_NN4BEG[1] ;
 wire \Tile_X4Y4_NN4BEG[2] ;
 wire \Tile_X4Y4_NN4BEG[3] ;
 wire \Tile_X4Y4_NN4BEG[4] ;
 wire \Tile_X4Y4_NN4BEG[5] ;
 wire \Tile_X4Y4_NN4BEG[6] ;
 wire \Tile_X4Y4_NN4BEG[7] ;
 wire \Tile_X4Y4_NN4BEG[8] ;
 wire \Tile_X4Y4_NN4BEG[9] ;
 wire \Tile_X4Y4_S1BEG[0] ;
 wire \Tile_X4Y4_S1BEG[1] ;
 wire \Tile_X4Y4_S1BEG[2] ;
 wire \Tile_X4Y4_S1BEG[3] ;
 wire \Tile_X4Y4_S2BEG[0] ;
 wire \Tile_X4Y4_S2BEG[1] ;
 wire \Tile_X4Y4_S2BEG[2] ;
 wire \Tile_X4Y4_S2BEG[3] ;
 wire \Tile_X4Y4_S2BEG[4] ;
 wire \Tile_X4Y4_S2BEG[5] ;
 wire \Tile_X4Y4_S2BEG[6] ;
 wire \Tile_X4Y4_S2BEG[7] ;
 wire \Tile_X4Y4_S2BEGb[0] ;
 wire \Tile_X4Y4_S2BEGb[1] ;
 wire \Tile_X4Y4_S2BEGb[2] ;
 wire \Tile_X4Y4_S2BEGb[3] ;
 wire \Tile_X4Y4_S2BEGb[4] ;
 wire \Tile_X4Y4_S2BEGb[5] ;
 wire \Tile_X4Y4_S2BEGb[6] ;
 wire \Tile_X4Y4_S2BEGb[7] ;
 wire \Tile_X4Y4_S4BEG[0] ;
 wire \Tile_X4Y4_S4BEG[10] ;
 wire \Tile_X4Y4_S4BEG[11] ;
 wire \Tile_X4Y4_S4BEG[12] ;
 wire \Tile_X4Y4_S4BEG[13] ;
 wire \Tile_X4Y4_S4BEG[14] ;
 wire \Tile_X4Y4_S4BEG[15] ;
 wire \Tile_X4Y4_S4BEG[1] ;
 wire \Tile_X4Y4_S4BEG[2] ;
 wire \Tile_X4Y4_S4BEG[3] ;
 wire \Tile_X4Y4_S4BEG[4] ;
 wire \Tile_X4Y4_S4BEG[5] ;
 wire \Tile_X4Y4_S4BEG[6] ;
 wire \Tile_X4Y4_S4BEG[7] ;
 wire \Tile_X4Y4_S4BEG[8] ;
 wire \Tile_X4Y4_S4BEG[9] ;
 wire \Tile_X4Y4_SS4BEG[0] ;
 wire \Tile_X4Y4_SS4BEG[10] ;
 wire \Tile_X4Y4_SS4BEG[11] ;
 wire \Tile_X4Y4_SS4BEG[12] ;
 wire \Tile_X4Y4_SS4BEG[13] ;
 wire \Tile_X4Y4_SS4BEG[14] ;
 wire \Tile_X4Y4_SS4BEG[15] ;
 wire \Tile_X4Y4_SS4BEG[1] ;
 wire \Tile_X4Y4_SS4BEG[2] ;
 wire \Tile_X4Y4_SS4BEG[3] ;
 wire \Tile_X4Y4_SS4BEG[4] ;
 wire \Tile_X4Y4_SS4BEG[5] ;
 wire \Tile_X4Y4_SS4BEG[6] ;
 wire \Tile_X4Y4_SS4BEG[7] ;
 wire \Tile_X4Y4_SS4BEG[8] ;
 wire \Tile_X4Y4_SS4BEG[9] ;
 wire Tile_X4Y4_UserCLKo;
 wire \Tile_X4Y4_W1BEG[0] ;
 wire \Tile_X4Y4_W1BEG[1] ;
 wire \Tile_X4Y4_W1BEG[2] ;
 wire \Tile_X4Y4_W1BEG[3] ;
 wire \Tile_X4Y4_W2BEG[0] ;
 wire \Tile_X4Y4_W2BEG[1] ;
 wire \Tile_X4Y4_W2BEG[2] ;
 wire \Tile_X4Y4_W2BEG[3] ;
 wire \Tile_X4Y4_W2BEG[4] ;
 wire \Tile_X4Y4_W2BEG[5] ;
 wire \Tile_X4Y4_W2BEG[6] ;
 wire \Tile_X4Y4_W2BEG[7] ;
 wire \Tile_X4Y4_W2BEGb[0] ;
 wire \Tile_X4Y4_W2BEGb[1] ;
 wire \Tile_X4Y4_W2BEGb[2] ;
 wire \Tile_X4Y4_W2BEGb[3] ;
 wire \Tile_X4Y4_W2BEGb[4] ;
 wire \Tile_X4Y4_W2BEGb[5] ;
 wire \Tile_X4Y4_W2BEGb[6] ;
 wire \Tile_X4Y4_W2BEGb[7] ;
 wire \Tile_X4Y4_W6BEG[0] ;
 wire \Tile_X4Y4_W6BEG[10] ;
 wire \Tile_X4Y4_W6BEG[11] ;
 wire \Tile_X4Y4_W6BEG[1] ;
 wire \Tile_X4Y4_W6BEG[2] ;
 wire \Tile_X4Y4_W6BEG[3] ;
 wire \Tile_X4Y4_W6BEG[4] ;
 wire \Tile_X4Y4_W6BEG[5] ;
 wire \Tile_X4Y4_W6BEG[6] ;
 wire \Tile_X4Y4_W6BEG[7] ;
 wire \Tile_X4Y4_W6BEG[8] ;
 wire \Tile_X4Y4_W6BEG[9] ;
 wire \Tile_X4Y4_WW4BEG[0] ;
 wire \Tile_X4Y4_WW4BEG[10] ;
 wire \Tile_X4Y4_WW4BEG[11] ;
 wire \Tile_X4Y4_WW4BEG[12] ;
 wire \Tile_X4Y4_WW4BEG[13] ;
 wire \Tile_X4Y4_WW4BEG[14] ;
 wire \Tile_X4Y4_WW4BEG[15] ;
 wire \Tile_X4Y4_WW4BEG[1] ;
 wire \Tile_X4Y4_WW4BEG[2] ;
 wire \Tile_X4Y4_WW4BEG[3] ;
 wire \Tile_X4Y4_WW4BEG[4] ;
 wire \Tile_X4Y4_WW4BEG[5] ;
 wire \Tile_X4Y4_WW4BEG[6] ;
 wire \Tile_X4Y4_WW4BEG[7] ;
 wire \Tile_X4Y4_WW4BEG[8] ;
 wire \Tile_X4Y4_WW4BEG[9] ;
 wire Tile_X4Y5_Co;
 wire \Tile_X4Y5_E1BEG[0] ;
 wire \Tile_X4Y5_E1BEG[1] ;
 wire \Tile_X4Y5_E1BEG[2] ;
 wire \Tile_X4Y5_E1BEG[3] ;
 wire \Tile_X4Y5_E2BEG[0] ;
 wire \Tile_X4Y5_E2BEG[1] ;
 wire \Tile_X4Y5_E2BEG[2] ;
 wire \Tile_X4Y5_E2BEG[3] ;
 wire \Tile_X4Y5_E2BEG[4] ;
 wire \Tile_X4Y5_E2BEG[5] ;
 wire \Tile_X4Y5_E2BEG[6] ;
 wire \Tile_X4Y5_E2BEG[7] ;
 wire \Tile_X4Y5_E2BEGb[0] ;
 wire \Tile_X4Y5_E2BEGb[1] ;
 wire \Tile_X4Y5_E2BEGb[2] ;
 wire \Tile_X4Y5_E2BEGb[3] ;
 wire \Tile_X4Y5_E2BEGb[4] ;
 wire \Tile_X4Y5_E2BEGb[5] ;
 wire \Tile_X4Y5_E2BEGb[6] ;
 wire \Tile_X4Y5_E2BEGb[7] ;
 wire \Tile_X4Y5_E6BEG[0] ;
 wire \Tile_X4Y5_E6BEG[10] ;
 wire \Tile_X4Y5_E6BEG[11] ;
 wire \Tile_X4Y5_E6BEG[1] ;
 wire \Tile_X4Y5_E6BEG[2] ;
 wire \Tile_X4Y5_E6BEG[3] ;
 wire \Tile_X4Y5_E6BEG[4] ;
 wire \Tile_X4Y5_E6BEG[5] ;
 wire \Tile_X4Y5_E6BEG[6] ;
 wire \Tile_X4Y5_E6BEG[7] ;
 wire \Tile_X4Y5_E6BEG[8] ;
 wire \Tile_X4Y5_E6BEG[9] ;
 wire \Tile_X4Y5_EE4BEG[0] ;
 wire \Tile_X4Y5_EE4BEG[10] ;
 wire \Tile_X4Y5_EE4BEG[11] ;
 wire \Tile_X4Y5_EE4BEG[12] ;
 wire \Tile_X4Y5_EE4BEG[13] ;
 wire \Tile_X4Y5_EE4BEG[14] ;
 wire \Tile_X4Y5_EE4BEG[15] ;
 wire \Tile_X4Y5_EE4BEG[1] ;
 wire \Tile_X4Y5_EE4BEG[2] ;
 wire \Tile_X4Y5_EE4BEG[3] ;
 wire \Tile_X4Y5_EE4BEG[4] ;
 wire \Tile_X4Y5_EE4BEG[5] ;
 wire \Tile_X4Y5_EE4BEG[6] ;
 wire \Tile_X4Y5_EE4BEG[7] ;
 wire \Tile_X4Y5_EE4BEG[8] ;
 wire \Tile_X4Y5_EE4BEG[9] ;
 wire \Tile_X4Y5_FrameData_O[0] ;
 wire \Tile_X4Y5_FrameData_O[10] ;
 wire \Tile_X4Y5_FrameData_O[11] ;
 wire \Tile_X4Y5_FrameData_O[12] ;
 wire \Tile_X4Y5_FrameData_O[13] ;
 wire \Tile_X4Y5_FrameData_O[14] ;
 wire \Tile_X4Y5_FrameData_O[15] ;
 wire \Tile_X4Y5_FrameData_O[16] ;
 wire \Tile_X4Y5_FrameData_O[17] ;
 wire \Tile_X4Y5_FrameData_O[18] ;
 wire \Tile_X4Y5_FrameData_O[19] ;
 wire \Tile_X4Y5_FrameData_O[1] ;
 wire \Tile_X4Y5_FrameData_O[20] ;
 wire \Tile_X4Y5_FrameData_O[21] ;
 wire \Tile_X4Y5_FrameData_O[22] ;
 wire \Tile_X4Y5_FrameData_O[23] ;
 wire \Tile_X4Y5_FrameData_O[24] ;
 wire \Tile_X4Y5_FrameData_O[25] ;
 wire \Tile_X4Y5_FrameData_O[26] ;
 wire \Tile_X4Y5_FrameData_O[27] ;
 wire \Tile_X4Y5_FrameData_O[28] ;
 wire \Tile_X4Y5_FrameData_O[29] ;
 wire \Tile_X4Y5_FrameData_O[2] ;
 wire \Tile_X4Y5_FrameData_O[30] ;
 wire \Tile_X4Y5_FrameData_O[31] ;
 wire \Tile_X4Y5_FrameData_O[3] ;
 wire \Tile_X4Y5_FrameData_O[4] ;
 wire \Tile_X4Y5_FrameData_O[5] ;
 wire \Tile_X4Y5_FrameData_O[6] ;
 wire \Tile_X4Y5_FrameData_O[7] ;
 wire \Tile_X4Y5_FrameData_O[8] ;
 wire \Tile_X4Y5_FrameData_O[9] ;
 wire \Tile_X4Y5_FrameStrobe_O[0] ;
 wire \Tile_X4Y5_FrameStrobe_O[10] ;
 wire \Tile_X4Y5_FrameStrobe_O[11] ;
 wire \Tile_X4Y5_FrameStrobe_O[12] ;
 wire \Tile_X4Y5_FrameStrobe_O[13] ;
 wire \Tile_X4Y5_FrameStrobe_O[14] ;
 wire \Tile_X4Y5_FrameStrobe_O[15] ;
 wire \Tile_X4Y5_FrameStrobe_O[16] ;
 wire \Tile_X4Y5_FrameStrobe_O[17] ;
 wire \Tile_X4Y5_FrameStrobe_O[18] ;
 wire \Tile_X4Y5_FrameStrobe_O[19] ;
 wire \Tile_X4Y5_FrameStrobe_O[1] ;
 wire \Tile_X4Y5_FrameStrobe_O[2] ;
 wire \Tile_X4Y5_FrameStrobe_O[3] ;
 wire \Tile_X4Y5_FrameStrobe_O[4] ;
 wire \Tile_X4Y5_FrameStrobe_O[5] ;
 wire \Tile_X4Y5_FrameStrobe_O[6] ;
 wire \Tile_X4Y5_FrameStrobe_O[7] ;
 wire \Tile_X4Y5_FrameStrobe_O[8] ;
 wire \Tile_X4Y5_FrameStrobe_O[9] ;
 wire \Tile_X4Y5_N1BEG[0] ;
 wire \Tile_X4Y5_N1BEG[1] ;
 wire \Tile_X4Y5_N1BEG[2] ;
 wire \Tile_X4Y5_N1BEG[3] ;
 wire \Tile_X4Y5_N2BEG[0] ;
 wire \Tile_X4Y5_N2BEG[1] ;
 wire \Tile_X4Y5_N2BEG[2] ;
 wire \Tile_X4Y5_N2BEG[3] ;
 wire \Tile_X4Y5_N2BEG[4] ;
 wire \Tile_X4Y5_N2BEG[5] ;
 wire \Tile_X4Y5_N2BEG[6] ;
 wire \Tile_X4Y5_N2BEG[7] ;
 wire \Tile_X4Y5_N2BEGb[0] ;
 wire \Tile_X4Y5_N2BEGb[1] ;
 wire \Tile_X4Y5_N2BEGb[2] ;
 wire \Tile_X4Y5_N2BEGb[3] ;
 wire \Tile_X4Y5_N2BEGb[4] ;
 wire \Tile_X4Y5_N2BEGb[5] ;
 wire \Tile_X4Y5_N2BEGb[6] ;
 wire \Tile_X4Y5_N2BEGb[7] ;
 wire \Tile_X4Y5_N4BEG[0] ;
 wire \Tile_X4Y5_N4BEG[10] ;
 wire \Tile_X4Y5_N4BEG[11] ;
 wire \Tile_X4Y5_N4BEG[12] ;
 wire \Tile_X4Y5_N4BEG[13] ;
 wire \Tile_X4Y5_N4BEG[14] ;
 wire \Tile_X4Y5_N4BEG[15] ;
 wire \Tile_X4Y5_N4BEG[1] ;
 wire \Tile_X4Y5_N4BEG[2] ;
 wire \Tile_X4Y5_N4BEG[3] ;
 wire \Tile_X4Y5_N4BEG[4] ;
 wire \Tile_X4Y5_N4BEG[5] ;
 wire \Tile_X4Y5_N4BEG[6] ;
 wire \Tile_X4Y5_N4BEG[7] ;
 wire \Tile_X4Y5_N4BEG[8] ;
 wire \Tile_X4Y5_N4BEG[9] ;
 wire \Tile_X4Y5_NN4BEG[0] ;
 wire \Tile_X4Y5_NN4BEG[10] ;
 wire \Tile_X4Y5_NN4BEG[11] ;
 wire \Tile_X4Y5_NN4BEG[12] ;
 wire \Tile_X4Y5_NN4BEG[13] ;
 wire \Tile_X4Y5_NN4BEG[14] ;
 wire \Tile_X4Y5_NN4BEG[15] ;
 wire \Tile_X4Y5_NN4BEG[1] ;
 wire \Tile_X4Y5_NN4BEG[2] ;
 wire \Tile_X4Y5_NN4BEG[3] ;
 wire \Tile_X4Y5_NN4BEG[4] ;
 wire \Tile_X4Y5_NN4BEG[5] ;
 wire \Tile_X4Y5_NN4BEG[6] ;
 wire \Tile_X4Y5_NN4BEG[7] ;
 wire \Tile_X4Y5_NN4BEG[8] ;
 wire \Tile_X4Y5_NN4BEG[9] ;
 wire \Tile_X4Y5_S1BEG[0] ;
 wire \Tile_X4Y5_S1BEG[1] ;
 wire \Tile_X4Y5_S1BEG[2] ;
 wire \Tile_X4Y5_S1BEG[3] ;
 wire \Tile_X4Y5_S2BEG[0] ;
 wire \Tile_X4Y5_S2BEG[1] ;
 wire \Tile_X4Y5_S2BEG[2] ;
 wire \Tile_X4Y5_S2BEG[3] ;
 wire \Tile_X4Y5_S2BEG[4] ;
 wire \Tile_X4Y5_S2BEG[5] ;
 wire \Tile_X4Y5_S2BEG[6] ;
 wire \Tile_X4Y5_S2BEG[7] ;
 wire \Tile_X4Y5_S2BEGb[0] ;
 wire \Tile_X4Y5_S2BEGb[1] ;
 wire \Tile_X4Y5_S2BEGb[2] ;
 wire \Tile_X4Y5_S2BEGb[3] ;
 wire \Tile_X4Y5_S2BEGb[4] ;
 wire \Tile_X4Y5_S2BEGb[5] ;
 wire \Tile_X4Y5_S2BEGb[6] ;
 wire \Tile_X4Y5_S2BEGb[7] ;
 wire \Tile_X4Y5_S4BEG[0] ;
 wire \Tile_X4Y5_S4BEG[10] ;
 wire \Tile_X4Y5_S4BEG[11] ;
 wire \Tile_X4Y5_S4BEG[12] ;
 wire \Tile_X4Y5_S4BEG[13] ;
 wire \Tile_X4Y5_S4BEG[14] ;
 wire \Tile_X4Y5_S4BEG[15] ;
 wire \Tile_X4Y5_S4BEG[1] ;
 wire \Tile_X4Y5_S4BEG[2] ;
 wire \Tile_X4Y5_S4BEG[3] ;
 wire \Tile_X4Y5_S4BEG[4] ;
 wire \Tile_X4Y5_S4BEG[5] ;
 wire \Tile_X4Y5_S4BEG[6] ;
 wire \Tile_X4Y5_S4BEG[7] ;
 wire \Tile_X4Y5_S4BEG[8] ;
 wire \Tile_X4Y5_S4BEG[9] ;
 wire \Tile_X4Y5_SS4BEG[0] ;
 wire \Tile_X4Y5_SS4BEG[10] ;
 wire \Tile_X4Y5_SS4BEG[11] ;
 wire \Tile_X4Y5_SS4BEG[12] ;
 wire \Tile_X4Y5_SS4BEG[13] ;
 wire \Tile_X4Y5_SS4BEG[14] ;
 wire \Tile_X4Y5_SS4BEG[15] ;
 wire \Tile_X4Y5_SS4BEG[1] ;
 wire \Tile_X4Y5_SS4BEG[2] ;
 wire \Tile_X4Y5_SS4BEG[3] ;
 wire \Tile_X4Y5_SS4BEG[4] ;
 wire \Tile_X4Y5_SS4BEG[5] ;
 wire \Tile_X4Y5_SS4BEG[6] ;
 wire \Tile_X4Y5_SS4BEG[7] ;
 wire \Tile_X4Y5_SS4BEG[8] ;
 wire \Tile_X4Y5_SS4BEG[9] ;
 wire Tile_X4Y5_UserCLKo;
 wire \Tile_X4Y5_W1BEG[0] ;
 wire \Tile_X4Y5_W1BEG[1] ;
 wire \Tile_X4Y5_W1BEG[2] ;
 wire \Tile_X4Y5_W1BEG[3] ;
 wire \Tile_X4Y5_W2BEG[0] ;
 wire \Tile_X4Y5_W2BEG[1] ;
 wire \Tile_X4Y5_W2BEG[2] ;
 wire \Tile_X4Y5_W2BEG[3] ;
 wire \Tile_X4Y5_W2BEG[4] ;
 wire \Tile_X4Y5_W2BEG[5] ;
 wire \Tile_X4Y5_W2BEG[6] ;
 wire \Tile_X4Y5_W2BEG[7] ;
 wire \Tile_X4Y5_W2BEGb[0] ;
 wire \Tile_X4Y5_W2BEGb[1] ;
 wire \Tile_X4Y5_W2BEGb[2] ;
 wire \Tile_X4Y5_W2BEGb[3] ;
 wire \Tile_X4Y5_W2BEGb[4] ;
 wire \Tile_X4Y5_W2BEGb[5] ;
 wire \Tile_X4Y5_W2BEGb[6] ;
 wire \Tile_X4Y5_W2BEGb[7] ;
 wire \Tile_X4Y5_W6BEG[0] ;
 wire \Tile_X4Y5_W6BEG[10] ;
 wire \Tile_X4Y5_W6BEG[11] ;
 wire \Tile_X4Y5_W6BEG[1] ;
 wire \Tile_X4Y5_W6BEG[2] ;
 wire \Tile_X4Y5_W6BEG[3] ;
 wire \Tile_X4Y5_W6BEG[4] ;
 wire \Tile_X4Y5_W6BEG[5] ;
 wire \Tile_X4Y5_W6BEG[6] ;
 wire \Tile_X4Y5_W6BEG[7] ;
 wire \Tile_X4Y5_W6BEG[8] ;
 wire \Tile_X4Y5_W6BEG[9] ;
 wire \Tile_X4Y5_WW4BEG[0] ;
 wire \Tile_X4Y5_WW4BEG[10] ;
 wire \Tile_X4Y5_WW4BEG[11] ;
 wire \Tile_X4Y5_WW4BEG[12] ;
 wire \Tile_X4Y5_WW4BEG[13] ;
 wire \Tile_X4Y5_WW4BEG[14] ;
 wire \Tile_X4Y5_WW4BEG[15] ;
 wire \Tile_X4Y5_WW4BEG[1] ;
 wire \Tile_X4Y5_WW4BEG[2] ;
 wire \Tile_X4Y5_WW4BEG[3] ;
 wire \Tile_X4Y5_WW4BEG[4] ;
 wire \Tile_X4Y5_WW4BEG[5] ;
 wire \Tile_X4Y5_WW4BEG[6] ;
 wire \Tile_X4Y5_WW4BEG[7] ;
 wire \Tile_X4Y5_WW4BEG[8] ;
 wire \Tile_X4Y5_WW4BEG[9] ;
 wire Tile_X4Y6_Co;
 wire \Tile_X4Y6_E1BEG[0] ;
 wire \Tile_X4Y6_E1BEG[1] ;
 wire \Tile_X4Y6_E1BEG[2] ;
 wire \Tile_X4Y6_E1BEG[3] ;
 wire \Tile_X4Y6_E2BEG[0] ;
 wire \Tile_X4Y6_E2BEG[1] ;
 wire \Tile_X4Y6_E2BEG[2] ;
 wire \Tile_X4Y6_E2BEG[3] ;
 wire \Tile_X4Y6_E2BEG[4] ;
 wire \Tile_X4Y6_E2BEG[5] ;
 wire \Tile_X4Y6_E2BEG[6] ;
 wire \Tile_X4Y6_E2BEG[7] ;
 wire \Tile_X4Y6_E2BEGb[0] ;
 wire \Tile_X4Y6_E2BEGb[1] ;
 wire \Tile_X4Y6_E2BEGb[2] ;
 wire \Tile_X4Y6_E2BEGb[3] ;
 wire \Tile_X4Y6_E2BEGb[4] ;
 wire \Tile_X4Y6_E2BEGb[5] ;
 wire \Tile_X4Y6_E2BEGb[6] ;
 wire \Tile_X4Y6_E2BEGb[7] ;
 wire \Tile_X4Y6_E6BEG[0] ;
 wire \Tile_X4Y6_E6BEG[10] ;
 wire \Tile_X4Y6_E6BEG[11] ;
 wire \Tile_X4Y6_E6BEG[1] ;
 wire \Tile_X4Y6_E6BEG[2] ;
 wire \Tile_X4Y6_E6BEG[3] ;
 wire \Tile_X4Y6_E6BEG[4] ;
 wire \Tile_X4Y6_E6BEG[5] ;
 wire \Tile_X4Y6_E6BEG[6] ;
 wire \Tile_X4Y6_E6BEG[7] ;
 wire \Tile_X4Y6_E6BEG[8] ;
 wire \Tile_X4Y6_E6BEG[9] ;
 wire \Tile_X4Y6_EE4BEG[0] ;
 wire \Tile_X4Y6_EE4BEG[10] ;
 wire \Tile_X4Y6_EE4BEG[11] ;
 wire \Tile_X4Y6_EE4BEG[12] ;
 wire \Tile_X4Y6_EE4BEG[13] ;
 wire \Tile_X4Y6_EE4BEG[14] ;
 wire \Tile_X4Y6_EE4BEG[15] ;
 wire \Tile_X4Y6_EE4BEG[1] ;
 wire \Tile_X4Y6_EE4BEG[2] ;
 wire \Tile_X4Y6_EE4BEG[3] ;
 wire \Tile_X4Y6_EE4BEG[4] ;
 wire \Tile_X4Y6_EE4BEG[5] ;
 wire \Tile_X4Y6_EE4BEG[6] ;
 wire \Tile_X4Y6_EE4BEG[7] ;
 wire \Tile_X4Y6_EE4BEG[8] ;
 wire \Tile_X4Y6_EE4BEG[9] ;
 wire \Tile_X4Y6_FrameData_O[0] ;
 wire \Tile_X4Y6_FrameData_O[10] ;
 wire \Tile_X4Y6_FrameData_O[11] ;
 wire \Tile_X4Y6_FrameData_O[12] ;
 wire \Tile_X4Y6_FrameData_O[13] ;
 wire \Tile_X4Y6_FrameData_O[14] ;
 wire \Tile_X4Y6_FrameData_O[15] ;
 wire \Tile_X4Y6_FrameData_O[16] ;
 wire \Tile_X4Y6_FrameData_O[17] ;
 wire \Tile_X4Y6_FrameData_O[18] ;
 wire \Tile_X4Y6_FrameData_O[19] ;
 wire \Tile_X4Y6_FrameData_O[1] ;
 wire \Tile_X4Y6_FrameData_O[20] ;
 wire \Tile_X4Y6_FrameData_O[21] ;
 wire \Tile_X4Y6_FrameData_O[22] ;
 wire \Tile_X4Y6_FrameData_O[23] ;
 wire \Tile_X4Y6_FrameData_O[24] ;
 wire \Tile_X4Y6_FrameData_O[25] ;
 wire \Tile_X4Y6_FrameData_O[26] ;
 wire \Tile_X4Y6_FrameData_O[27] ;
 wire \Tile_X4Y6_FrameData_O[28] ;
 wire \Tile_X4Y6_FrameData_O[29] ;
 wire \Tile_X4Y6_FrameData_O[2] ;
 wire \Tile_X4Y6_FrameData_O[30] ;
 wire \Tile_X4Y6_FrameData_O[31] ;
 wire \Tile_X4Y6_FrameData_O[3] ;
 wire \Tile_X4Y6_FrameData_O[4] ;
 wire \Tile_X4Y6_FrameData_O[5] ;
 wire \Tile_X4Y6_FrameData_O[6] ;
 wire \Tile_X4Y6_FrameData_O[7] ;
 wire \Tile_X4Y6_FrameData_O[8] ;
 wire \Tile_X4Y6_FrameData_O[9] ;
 wire \Tile_X4Y6_FrameStrobe_O[0] ;
 wire \Tile_X4Y6_FrameStrobe_O[10] ;
 wire \Tile_X4Y6_FrameStrobe_O[11] ;
 wire \Tile_X4Y6_FrameStrobe_O[12] ;
 wire \Tile_X4Y6_FrameStrobe_O[13] ;
 wire \Tile_X4Y6_FrameStrobe_O[14] ;
 wire \Tile_X4Y6_FrameStrobe_O[15] ;
 wire \Tile_X4Y6_FrameStrobe_O[16] ;
 wire \Tile_X4Y6_FrameStrobe_O[17] ;
 wire \Tile_X4Y6_FrameStrobe_O[18] ;
 wire \Tile_X4Y6_FrameStrobe_O[19] ;
 wire \Tile_X4Y6_FrameStrobe_O[1] ;
 wire \Tile_X4Y6_FrameStrobe_O[2] ;
 wire \Tile_X4Y6_FrameStrobe_O[3] ;
 wire \Tile_X4Y6_FrameStrobe_O[4] ;
 wire \Tile_X4Y6_FrameStrobe_O[5] ;
 wire \Tile_X4Y6_FrameStrobe_O[6] ;
 wire \Tile_X4Y6_FrameStrobe_O[7] ;
 wire \Tile_X4Y6_FrameStrobe_O[8] ;
 wire \Tile_X4Y6_FrameStrobe_O[9] ;
 wire \Tile_X4Y6_N1BEG[0] ;
 wire \Tile_X4Y6_N1BEG[1] ;
 wire \Tile_X4Y6_N1BEG[2] ;
 wire \Tile_X4Y6_N1BEG[3] ;
 wire \Tile_X4Y6_N2BEG[0] ;
 wire \Tile_X4Y6_N2BEG[1] ;
 wire \Tile_X4Y6_N2BEG[2] ;
 wire \Tile_X4Y6_N2BEG[3] ;
 wire \Tile_X4Y6_N2BEG[4] ;
 wire \Tile_X4Y6_N2BEG[5] ;
 wire \Tile_X4Y6_N2BEG[6] ;
 wire \Tile_X4Y6_N2BEG[7] ;
 wire \Tile_X4Y6_N2BEGb[0] ;
 wire \Tile_X4Y6_N2BEGb[1] ;
 wire \Tile_X4Y6_N2BEGb[2] ;
 wire \Tile_X4Y6_N2BEGb[3] ;
 wire \Tile_X4Y6_N2BEGb[4] ;
 wire \Tile_X4Y6_N2BEGb[5] ;
 wire \Tile_X4Y6_N2BEGb[6] ;
 wire \Tile_X4Y6_N2BEGb[7] ;
 wire \Tile_X4Y6_N4BEG[0] ;
 wire \Tile_X4Y6_N4BEG[10] ;
 wire \Tile_X4Y6_N4BEG[11] ;
 wire \Tile_X4Y6_N4BEG[12] ;
 wire \Tile_X4Y6_N4BEG[13] ;
 wire \Tile_X4Y6_N4BEG[14] ;
 wire \Tile_X4Y6_N4BEG[15] ;
 wire \Tile_X4Y6_N4BEG[1] ;
 wire \Tile_X4Y6_N4BEG[2] ;
 wire \Tile_X4Y6_N4BEG[3] ;
 wire \Tile_X4Y6_N4BEG[4] ;
 wire \Tile_X4Y6_N4BEG[5] ;
 wire \Tile_X4Y6_N4BEG[6] ;
 wire \Tile_X4Y6_N4BEG[7] ;
 wire \Tile_X4Y6_N4BEG[8] ;
 wire \Tile_X4Y6_N4BEG[9] ;
 wire \Tile_X4Y6_NN4BEG[0] ;
 wire \Tile_X4Y6_NN4BEG[10] ;
 wire \Tile_X4Y6_NN4BEG[11] ;
 wire \Tile_X4Y6_NN4BEG[12] ;
 wire \Tile_X4Y6_NN4BEG[13] ;
 wire \Tile_X4Y6_NN4BEG[14] ;
 wire \Tile_X4Y6_NN4BEG[15] ;
 wire \Tile_X4Y6_NN4BEG[1] ;
 wire \Tile_X4Y6_NN4BEG[2] ;
 wire \Tile_X4Y6_NN4BEG[3] ;
 wire \Tile_X4Y6_NN4BEG[4] ;
 wire \Tile_X4Y6_NN4BEG[5] ;
 wire \Tile_X4Y6_NN4BEG[6] ;
 wire \Tile_X4Y6_NN4BEG[7] ;
 wire \Tile_X4Y6_NN4BEG[8] ;
 wire \Tile_X4Y6_NN4BEG[9] ;
 wire \Tile_X4Y6_S1BEG[0] ;
 wire \Tile_X4Y6_S1BEG[1] ;
 wire \Tile_X4Y6_S1BEG[2] ;
 wire \Tile_X4Y6_S1BEG[3] ;
 wire \Tile_X4Y6_S2BEG[0] ;
 wire \Tile_X4Y6_S2BEG[1] ;
 wire \Tile_X4Y6_S2BEG[2] ;
 wire \Tile_X4Y6_S2BEG[3] ;
 wire \Tile_X4Y6_S2BEG[4] ;
 wire \Tile_X4Y6_S2BEG[5] ;
 wire \Tile_X4Y6_S2BEG[6] ;
 wire \Tile_X4Y6_S2BEG[7] ;
 wire \Tile_X4Y6_S2BEGb[0] ;
 wire \Tile_X4Y6_S2BEGb[1] ;
 wire \Tile_X4Y6_S2BEGb[2] ;
 wire \Tile_X4Y6_S2BEGb[3] ;
 wire \Tile_X4Y6_S2BEGb[4] ;
 wire \Tile_X4Y6_S2BEGb[5] ;
 wire \Tile_X4Y6_S2BEGb[6] ;
 wire \Tile_X4Y6_S2BEGb[7] ;
 wire \Tile_X4Y6_S4BEG[0] ;
 wire \Tile_X4Y6_S4BEG[10] ;
 wire \Tile_X4Y6_S4BEG[11] ;
 wire \Tile_X4Y6_S4BEG[12] ;
 wire \Tile_X4Y6_S4BEG[13] ;
 wire \Tile_X4Y6_S4BEG[14] ;
 wire \Tile_X4Y6_S4BEG[15] ;
 wire \Tile_X4Y6_S4BEG[1] ;
 wire \Tile_X4Y6_S4BEG[2] ;
 wire \Tile_X4Y6_S4BEG[3] ;
 wire \Tile_X4Y6_S4BEG[4] ;
 wire \Tile_X4Y6_S4BEG[5] ;
 wire \Tile_X4Y6_S4BEG[6] ;
 wire \Tile_X4Y6_S4BEG[7] ;
 wire \Tile_X4Y6_S4BEG[8] ;
 wire \Tile_X4Y6_S4BEG[9] ;
 wire \Tile_X4Y6_SS4BEG[0] ;
 wire \Tile_X4Y6_SS4BEG[10] ;
 wire \Tile_X4Y6_SS4BEG[11] ;
 wire \Tile_X4Y6_SS4BEG[12] ;
 wire \Tile_X4Y6_SS4BEG[13] ;
 wire \Tile_X4Y6_SS4BEG[14] ;
 wire \Tile_X4Y6_SS4BEG[15] ;
 wire \Tile_X4Y6_SS4BEG[1] ;
 wire \Tile_X4Y6_SS4BEG[2] ;
 wire \Tile_X4Y6_SS4BEG[3] ;
 wire \Tile_X4Y6_SS4BEG[4] ;
 wire \Tile_X4Y6_SS4BEG[5] ;
 wire \Tile_X4Y6_SS4BEG[6] ;
 wire \Tile_X4Y6_SS4BEG[7] ;
 wire \Tile_X4Y6_SS4BEG[8] ;
 wire \Tile_X4Y6_SS4BEG[9] ;
 wire Tile_X4Y6_UserCLKo;
 wire \Tile_X4Y6_W1BEG[0] ;
 wire \Tile_X4Y6_W1BEG[1] ;
 wire \Tile_X4Y6_W1BEG[2] ;
 wire \Tile_X4Y6_W1BEG[3] ;
 wire \Tile_X4Y6_W2BEG[0] ;
 wire \Tile_X4Y6_W2BEG[1] ;
 wire \Tile_X4Y6_W2BEG[2] ;
 wire \Tile_X4Y6_W2BEG[3] ;
 wire \Tile_X4Y6_W2BEG[4] ;
 wire \Tile_X4Y6_W2BEG[5] ;
 wire \Tile_X4Y6_W2BEG[6] ;
 wire \Tile_X4Y6_W2BEG[7] ;
 wire \Tile_X4Y6_W2BEGb[0] ;
 wire \Tile_X4Y6_W2BEGb[1] ;
 wire \Tile_X4Y6_W2BEGb[2] ;
 wire \Tile_X4Y6_W2BEGb[3] ;
 wire \Tile_X4Y6_W2BEGb[4] ;
 wire \Tile_X4Y6_W2BEGb[5] ;
 wire \Tile_X4Y6_W2BEGb[6] ;
 wire \Tile_X4Y6_W2BEGb[7] ;
 wire \Tile_X4Y6_W6BEG[0] ;
 wire \Tile_X4Y6_W6BEG[10] ;
 wire \Tile_X4Y6_W6BEG[11] ;
 wire \Tile_X4Y6_W6BEG[1] ;
 wire \Tile_X4Y6_W6BEG[2] ;
 wire \Tile_X4Y6_W6BEG[3] ;
 wire \Tile_X4Y6_W6BEG[4] ;
 wire \Tile_X4Y6_W6BEG[5] ;
 wire \Tile_X4Y6_W6BEG[6] ;
 wire \Tile_X4Y6_W6BEG[7] ;
 wire \Tile_X4Y6_W6BEG[8] ;
 wire \Tile_X4Y6_W6BEG[9] ;
 wire \Tile_X4Y6_WW4BEG[0] ;
 wire \Tile_X4Y6_WW4BEG[10] ;
 wire \Tile_X4Y6_WW4BEG[11] ;
 wire \Tile_X4Y6_WW4BEG[12] ;
 wire \Tile_X4Y6_WW4BEG[13] ;
 wire \Tile_X4Y6_WW4BEG[14] ;
 wire \Tile_X4Y6_WW4BEG[15] ;
 wire \Tile_X4Y6_WW4BEG[1] ;
 wire \Tile_X4Y6_WW4BEG[2] ;
 wire \Tile_X4Y6_WW4BEG[3] ;
 wire \Tile_X4Y6_WW4BEG[4] ;
 wire \Tile_X4Y6_WW4BEG[5] ;
 wire \Tile_X4Y6_WW4BEG[6] ;
 wire \Tile_X4Y6_WW4BEG[7] ;
 wire \Tile_X4Y6_WW4BEG[8] ;
 wire \Tile_X4Y6_WW4BEG[9] ;
 wire Tile_X4Y7_Co;
 wire \Tile_X4Y7_E1BEG[0] ;
 wire \Tile_X4Y7_E1BEG[1] ;
 wire \Tile_X4Y7_E1BEG[2] ;
 wire \Tile_X4Y7_E1BEG[3] ;
 wire \Tile_X4Y7_E2BEG[0] ;
 wire \Tile_X4Y7_E2BEG[1] ;
 wire \Tile_X4Y7_E2BEG[2] ;
 wire \Tile_X4Y7_E2BEG[3] ;
 wire \Tile_X4Y7_E2BEG[4] ;
 wire \Tile_X4Y7_E2BEG[5] ;
 wire \Tile_X4Y7_E2BEG[6] ;
 wire \Tile_X4Y7_E2BEG[7] ;
 wire \Tile_X4Y7_E2BEGb[0] ;
 wire \Tile_X4Y7_E2BEGb[1] ;
 wire \Tile_X4Y7_E2BEGb[2] ;
 wire \Tile_X4Y7_E2BEGb[3] ;
 wire \Tile_X4Y7_E2BEGb[4] ;
 wire \Tile_X4Y7_E2BEGb[5] ;
 wire \Tile_X4Y7_E2BEGb[6] ;
 wire \Tile_X4Y7_E2BEGb[7] ;
 wire \Tile_X4Y7_E6BEG[0] ;
 wire \Tile_X4Y7_E6BEG[10] ;
 wire \Tile_X4Y7_E6BEG[11] ;
 wire \Tile_X4Y7_E6BEG[1] ;
 wire \Tile_X4Y7_E6BEG[2] ;
 wire \Tile_X4Y7_E6BEG[3] ;
 wire \Tile_X4Y7_E6BEG[4] ;
 wire \Tile_X4Y7_E6BEG[5] ;
 wire \Tile_X4Y7_E6BEG[6] ;
 wire \Tile_X4Y7_E6BEG[7] ;
 wire \Tile_X4Y7_E6BEG[8] ;
 wire \Tile_X4Y7_E6BEG[9] ;
 wire \Tile_X4Y7_EE4BEG[0] ;
 wire \Tile_X4Y7_EE4BEG[10] ;
 wire \Tile_X4Y7_EE4BEG[11] ;
 wire \Tile_X4Y7_EE4BEG[12] ;
 wire \Tile_X4Y7_EE4BEG[13] ;
 wire \Tile_X4Y7_EE4BEG[14] ;
 wire \Tile_X4Y7_EE4BEG[15] ;
 wire \Tile_X4Y7_EE4BEG[1] ;
 wire \Tile_X4Y7_EE4BEG[2] ;
 wire \Tile_X4Y7_EE4BEG[3] ;
 wire \Tile_X4Y7_EE4BEG[4] ;
 wire \Tile_X4Y7_EE4BEG[5] ;
 wire \Tile_X4Y7_EE4BEG[6] ;
 wire \Tile_X4Y7_EE4BEG[7] ;
 wire \Tile_X4Y7_EE4BEG[8] ;
 wire \Tile_X4Y7_EE4BEG[9] ;
 wire \Tile_X4Y7_FrameData_O[0] ;
 wire \Tile_X4Y7_FrameData_O[10] ;
 wire \Tile_X4Y7_FrameData_O[11] ;
 wire \Tile_X4Y7_FrameData_O[12] ;
 wire \Tile_X4Y7_FrameData_O[13] ;
 wire \Tile_X4Y7_FrameData_O[14] ;
 wire \Tile_X4Y7_FrameData_O[15] ;
 wire \Tile_X4Y7_FrameData_O[16] ;
 wire \Tile_X4Y7_FrameData_O[17] ;
 wire \Tile_X4Y7_FrameData_O[18] ;
 wire \Tile_X4Y7_FrameData_O[19] ;
 wire \Tile_X4Y7_FrameData_O[1] ;
 wire \Tile_X4Y7_FrameData_O[20] ;
 wire \Tile_X4Y7_FrameData_O[21] ;
 wire \Tile_X4Y7_FrameData_O[22] ;
 wire \Tile_X4Y7_FrameData_O[23] ;
 wire \Tile_X4Y7_FrameData_O[24] ;
 wire \Tile_X4Y7_FrameData_O[25] ;
 wire \Tile_X4Y7_FrameData_O[26] ;
 wire \Tile_X4Y7_FrameData_O[27] ;
 wire \Tile_X4Y7_FrameData_O[28] ;
 wire \Tile_X4Y7_FrameData_O[29] ;
 wire \Tile_X4Y7_FrameData_O[2] ;
 wire \Tile_X4Y7_FrameData_O[30] ;
 wire \Tile_X4Y7_FrameData_O[31] ;
 wire \Tile_X4Y7_FrameData_O[3] ;
 wire \Tile_X4Y7_FrameData_O[4] ;
 wire \Tile_X4Y7_FrameData_O[5] ;
 wire \Tile_X4Y7_FrameData_O[6] ;
 wire \Tile_X4Y7_FrameData_O[7] ;
 wire \Tile_X4Y7_FrameData_O[8] ;
 wire \Tile_X4Y7_FrameData_O[9] ;
 wire \Tile_X4Y7_FrameStrobe_O[0] ;
 wire \Tile_X4Y7_FrameStrobe_O[10] ;
 wire \Tile_X4Y7_FrameStrobe_O[11] ;
 wire \Tile_X4Y7_FrameStrobe_O[12] ;
 wire \Tile_X4Y7_FrameStrobe_O[13] ;
 wire \Tile_X4Y7_FrameStrobe_O[14] ;
 wire \Tile_X4Y7_FrameStrobe_O[15] ;
 wire \Tile_X4Y7_FrameStrobe_O[16] ;
 wire \Tile_X4Y7_FrameStrobe_O[17] ;
 wire \Tile_X4Y7_FrameStrobe_O[18] ;
 wire \Tile_X4Y7_FrameStrobe_O[19] ;
 wire \Tile_X4Y7_FrameStrobe_O[1] ;
 wire \Tile_X4Y7_FrameStrobe_O[2] ;
 wire \Tile_X4Y7_FrameStrobe_O[3] ;
 wire \Tile_X4Y7_FrameStrobe_O[4] ;
 wire \Tile_X4Y7_FrameStrobe_O[5] ;
 wire \Tile_X4Y7_FrameStrobe_O[6] ;
 wire \Tile_X4Y7_FrameStrobe_O[7] ;
 wire \Tile_X4Y7_FrameStrobe_O[8] ;
 wire \Tile_X4Y7_FrameStrobe_O[9] ;
 wire \Tile_X4Y7_N1BEG[0] ;
 wire \Tile_X4Y7_N1BEG[1] ;
 wire \Tile_X4Y7_N1BEG[2] ;
 wire \Tile_X4Y7_N1BEG[3] ;
 wire \Tile_X4Y7_N2BEG[0] ;
 wire \Tile_X4Y7_N2BEG[1] ;
 wire \Tile_X4Y7_N2BEG[2] ;
 wire \Tile_X4Y7_N2BEG[3] ;
 wire \Tile_X4Y7_N2BEG[4] ;
 wire \Tile_X4Y7_N2BEG[5] ;
 wire \Tile_X4Y7_N2BEG[6] ;
 wire \Tile_X4Y7_N2BEG[7] ;
 wire \Tile_X4Y7_N2BEGb[0] ;
 wire \Tile_X4Y7_N2BEGb[1] ;
 wire \Tile_X4Y7_N2BEGb[2] ;
 wire \Tile_X4Y7_N2BEGb[3] ;
 wire \Tile_X4Y7_N2BEGb[4] ;
 wire \Tile_X4Y7_N2BEGb[5] ;
 wire \Tile_X4Y7_N2BEGb[6] ;
 wire \Tile_X4Y7_N2BEGb[7] ;
 wire \Tile_X4Y7_N4BEG[0] ;
 wire \Tile_X4Y7_N4BEG[10] ;
 wire \Tile_X4Y7_N4BEG[11] ;
 wire \Tile_X4Y7_N4BEG[12] ;
 wire \Tile_X4Y7_N4BEG[13] ;
 wire \Tile_X4Y7_N4BEG[14] ;
 wire \Tile_X4Y7_N4BEG[15] ;
 wire \Tile_X4Y7_N4BEG[1] ;
 wire \Tile_X4Y7_N4BEG[2] ;
 wire \Tile_X4Y7_N4BEG[3] ;
 wire \Tile_X4Y7_N4BEG[4] ;
 wire \Tile_X4Y7_N4BEG[5] ;
 wire \Tile_X4Y7_N4BEG[6] ;
 wire \Tile_X4Y7_N4BEG[7] ;
 wire \Tile_X4Y7_N4BEG[8] ;
 wire \Tile_X4Y7_N4BEG[9] ;
 wire \Tile_X4Y7_NN4BEG[0] ;
 wire \Tile_X4Y7_NN4BEG[10] ;
 wire \Tile_X4Y7_NN4BEG[11] ;
 wire \Tile_X4Y7_NN4BEG[12] ;
 wire \Tile_X4Y7_NN4BEG[13] ;
 wire \Tile_X4Y7_NN4BEG[14] ;
 wire \Tile_X4Y7_NN4BEG[15] ;
 wire \Tile_X4Y7_NN4BEG[1] ;
 wire \Tile_X4Y7_NN4BEG[2] ;
 wire \Tile_X4Y7_NN4BEG[3] ;
 wire \Tile_X4Y7_NN4BEG[4] ;
 wire \Tile_X4Y7_NN4BEG[5] ;
 wire \Tile_X4Y7_NN4BEG[6] ;
 wire \Tile_X4Y7_NN4BEG[7] ;
 wire \Tile_X4Y7_NN4BEG[8] ;
 wire \Tile_X4Y7_NN4BEG[9] ;
 wire \Tile_X4Y7_S1BEG[0] ;
 wire \Tile_X4Y7_S1BEG[1] ;
 wire \Tile_X4Y7_S1BEG[2] ;
 wire \Tile_X4Y7_S1BEG[3] ;
 wire \Tile_X4Y7_S2BEG[0] ;
 wire \Tile_X4Y7_S2BEG[1] ;
 wire \Tile_X4Y7_S2BEG[2] ;
 wire \Tile_X4Y7_S2BEG[3] ;
 wire \Tile_X4Y7_S2BEG[4] ;
 wire \Tile_X4Y7_S2BEG[5] ;
 wire \Tile_X4Y7_S2BEG[6] ;
 wire \Tile_X4Y7_S2BEG[7] ;
 wire \Tile_X4Y7_S2BEGb[0] ;
 wire \Tile_X4Y7_S2BEGb[1] ;
 wire \Tile_X4Y7_S2BEGb[2] ;
 wire \Tile_X4Y7_S2BEGb[3] ;
 wire \Tile_X4Y7_S2BEGb[4] ;
 wire \Tile_X4Y7_S2BEGb[5] ;
 wire \Tile_X4Y7_S2BEGb[6] ;
 wire \Tile_X4Y7_S2BEGb[7] ;
 wire \Tile_X4Y7_S4BEG[0] ;
 wire \Tile_X4Y7_S4BEG[10] ;
 wire \Tile_X4Y7_S4BEG[11] ;
 wire \Tile_X4Y7_S4BEG[12] ;
 wire \Tile_X4Y7_S4BEG[13] ;
 wire \Tile_X4Y7_S4BEG[14] ;
 wire \Tile_X4Y7_S4BEG[15] ;
 wire \Tile_X4Y7_S4BEG[1] ;
 wire \Tile_X4Y7_S4BEG[2] ;
 wire \Tile_X4Y7_S4BEG[3] ;
 wire \Tile_X4Y7_S4BEG[4] ;
 wire \Tile_X4Y7_S4BEG[5] ;
 wire \Tile_X4Y7_S4BEG[6] ;
 wire \Tile_X4Y7_S4BEG[7] ;
 wire \Tile_X4Y7_S4BEG[8] ;
 wire \Tile_X4Y7_S4BEG[9] ;
 wire \Tile_X4Y7_SS4BEG[0] ;
 wire \Tile_X4Y7_SS4BEG[10] ;
 wire \Tile_X4Y7_SS4BEG[11] ;
 wire \Tile_X4Y7_SS4BEG[12] ;
 wire \Tile_X4Y7_SS4BEG[13] ;
 wire \Tile_X4Y7_SS4BEG[14] ;
 wire \Tile_X4Y7_SS4BEG[15] ;
 wire \Tile_X4Y7_SS4BEG[1] ;
 wire \Tile_X4Y7_SS4BEG[2] ;
 wire \Tile_X4Y7_SS4BEG[3] ;
 wire \Tile_X4Y7_SS4BEG[4] ;
 wire \Tile_X4Y7_SS4BEG[5] ;
 wire \Tile_X4Y7_SS4BEG[6] ;
 wire \Tile_X4Y7_SS4BEG[7] ;
 wire \Tile_X4Y7_SS4BEG[8] ;
 wire \Tile_X4Y7_SS4BEG[9] ;
 wire Tile_X4Y7_UserCLKo;
 wire \Tile_X4Y7_W1BEG[0] ;
 wire \Tile_X4Y7_W1BEG[1] ;
 wire \Tile_X4Y7_W1BEG[2] ;
 wire \Tile_X4Y7_W1BEG[3] ;
 wire \Tile_X4Y7_W2BEG[0] ;
 wire \Tile_X4Y7_W2BEG[1] ;
 wire \Tile_X4Y7_W2BEG[2] ;
 wire \Tile_X4Y7_W2BEG[3] ;
 wire \Tile_X4Y7_W2BEG[4] ;
 wire \Tile_X4Y7_W2BEG[5] ;
 wire \Tile_X4Y7_W2BEG[6] ;
 wire \Tile_X4Y7_W2BEG[7] ;
 wire \Tile_X4Y7_W2BEGb[0] ;
 wire \Tile_X4Y7_W2BEGb[1] ;
 wire \Tile_X4Y7_W2BEGb[2] ;
 wire \Tile_X4Y7_W2BEGb[3] ;
 wire \Tile_X4Y7_W2BEGb[4] ;
 wire \Tile_X4Y7_W2BEGb[5] ;
 wire \Tile_X4Y7_W2BEGb[6] ;
 wire \Tile_X4Y7_W2BEGb[7] ;
 wire \Tile_X4Y7_W6BEG[0] ;
 wire \Tile_X4Y7_W6BEG[10] ;
 wire \Tile_X4Y7_W6BEG[11] ;
 wire \Tile_X4Y7_W6BEG[1] ;
 wire \Tile_X4Y7_W6BEG[2] ;
 wire \Tile_X4Y7_W6BEG[3] ;
 wire \Tile_X4Y7_W6BEG[4] ;
 wire \Tile_X4Y7_W6BEG[5] ;
 wire \Tile_X4Y7_W6BEG[6] ;
 wire \Tile_X4Y7_W6BEG[7] ;
 wire \Tile_X4Y7_W6BEG[8] ;
 wire \Tile_X4Y7_W6BEG[9] ;
 wire \Tile_X4Y7_WW4BEG[0] ;
 wire \Tile_X4Y7_WW4BEG[10] ;
 wire \Tile_X4Y7_WW4BEG[11] ;
 wire \Tile_X4Y7_WW4BEG[12] ;
 wire \Tile_X4Y7_WW4BEG[13] ;
 wire \Tile_X4Y7_WW4BEG[14] ;
 wire \Tile_X4Y7_WW4BEG[15] ;
 wire \Tile_X4Y7_WW4BEG[1] ;
 wire \Tile_X4Y7_WW4BEG[2] ;
 wire \Tile_X4Y7_WW4BEG[3] ;
 wire \Tile_X4Y7_WW4BEG[4] ;
 wire \Tile_X4Y7_WW4BEG[5] ;
 wire \Tile_X4Y7_WW4BEG[6] ;
 wire \Tile_X4Y7_WW4BEG[7] ;
 wire \Tile_X4Y7_WW4BEG[8] ;
 wire \Tile_X4Y7_WW4BEG[9] ;
 wire Tile_X4Y8_Co;
 wire \Tile_X4Y8_E1BEG[0] ;
 wire \Tile_X4Y8_E1BEG[1] ;
 wire \Tile_X4Y8_E1BEG[2] ;
 wire \Tile_X4Y8_E1BEG[3] ;
 wire \Tile_X4Y8_E2BEG[0] ;
 wire \Tile_X4Y8_E2BEG[1] ;
 wire \Tile_X4Y8_E2BEG[2] ;
 wire \Tile_X4Y8_E2BEG[3] ;
 wire \Tile_X4Y8_E2BEG[4] ;
 wire \Tile_X4Y8_E2BEG[5] ;
 wire \Tile_X4Y8_E2BEG[6] ;
 wire \Tile_X4Y8_E2BEG[7] ;
 wire \Tile_X4Y8_E2BEGb[0] ;
 wire \Tile_X4Y8_E2BEGb[1] ;
 wire \Tile_X4Y8_E2BEGb[2] ;
 wire \Tile_X4Y8_E2BEGb[3] ;
 wire \Tile_X4Y8_E2BEGb[4] ;
 wire \Tile_X4Y8_E2BEGb[5] ;
 wire \Tile_X4Y8_E2BEGb[6] ;
 wire \Tile_X4Y8_E2BEGb[7] ;
 wire \Tile_X4Y8_E6BEG[0] ;
 wire \Tile_X4Y8_E6BEG[10] ;
 wire \Tile_X4Y8_E6BEG[11] ;
 wire \Tile_X4Y8_E6BEG[1] ;
 wire \Tile_X4Y8_E6BEG[2] ;
 wire \Tile_X4Y8_E6BEG[3] ;
 wire \Tile_X4Y8_E6BEG[4] ;
 wire \Tile_X4Y8_E6BEG[5] ;
 wire \Tile_X4Y8_E6BEG[6] ;
 wire \Tile_X4Y8_E6BEG[7] ;
 wire \Tile_X4Y8_E6BEG[8] ;
 wire \Tile_X4Y8_E6BEG[9] ;
 wire \Tile_X4Y8_EE4BEG[0] ;
 wire \Tile_X4Y8_EE4BEG[10] ;
 wire \Tile_X4Y8_EE4BEG[11] ;
 wire \Tile_X4Y8_EE4BEG[12] ;
 wire \Tile_X4Y8_EE4BEG[13] ;
 wire \Tile_X4Y8_EE4BEG[14] ;
 wire \Tile_X4Y8_EE4BEG[15] ;
 wire \Tile_X4Y8_EE4BEG[1] ;
 wire \Tile_X4Y8_EE4BEG[2] ;
 wire \Tile_X4Y8_EE4BEG[3] ;
 wire \Tile_X4Y8_EE4BEG[4] ;
 wire \Tile_X4Y8_EE4BEG[5] ;
 wire \Tile_X4Y8_EE4BEG[6] ;
 wire \Tile_X4Y8_EE4BEG[7] ;
 wire \Tile_X4Y8_EE4BEG[8] ;
 wire \Tile_X4Y8_EE4BEG[9] ;
 wire \Tile_X4Y8_FrameData_O[0] ;
 wire \Tile_X4Y8_FrameData_O[10] ;
 wire \Tile_X4Y8_FrameData_O[11] ;
 wire \Tile_X4Y8_FrameData_O[12] ;
 wire \Tile_X4Y8_FrameData_O[13] ;
 wire \Tile_X4Y8_FrameData_O[14] ;
 wire \Tile_X4Y8_FrameData_O[15] ;
 wire \Tile_X4Y8_FrameData_O[16] ;
 wire \Tile_X4Y8_FrameData_O[17] ;
 wire \Tile_X4Y8_FrameData_O[18] ;
 wire \Tile_X4Y8_FrameData_O[19] ;
 wire \Tile_X4Y8_FrameData_O[1] ;
 wire \Tile_X4Y8_FrameData_O[20] ;
 wire \Tile_X4Y8_FrameData_O[21] ;
 wire \Tile_X4Y8_FrameData_O[22] ;
 wire \Tile_X4Y8_FrameData_O[23] ;
 wire \Tile_X4Y8_FrameData_O[24] ;
 wire \Tile_X4Y8_FrameData_O[25] ;
 wire \Tile_X4Y8_FrameData_O[26] ;
 wire \Tile_X4Y8_FrameData_O[27] ;
 wire \Tile_X4Y8_FrameData_O[28] ;
 wire \Tile_X4Y8_FrameData_O[29] ;
 wire \Tile_X4Y8_FrameData_O[2] ;
 wire \Tile_X4Y8_FrameData_O[30] ;
 wire \Tile_X4Y8_FrameData_O[31] ;
 wire \Tile_X4Y8_FrameData_O[3] ;
 wire \Tile_X4Y8_FrameData_O[4] ;
 wire \Tile_X4Y8_FrameData_O[5] ;
 wire \Tile_X4Y8_FrameData_O[6] ;
 wire \Tile_X4Y8_FrameData_O[7] ;
 wire \Tile_X4Y8_FrameData_O[8] ;
 wire \Tile_X4Y8_FrameData_O[9] ;
 wire \Tile_X4Y8_FrameStrobe_O[0] ;
 wire \Tile_X4Y8_FrameStrobe_O[10] ;
 wire \Tile_X4Y8_FrameStrobe_O[11] ;
 wire \Tile_X4Y8_FrameStrobe_O[12] ;
 wire \Tile_X4Y8_FrameStrobe_O[13] ;
 wire \Tile_X4Y8_FrameStrobe_O[14] ;
 wire \Tile_X4Y8_FrameStrobe_O[15] ;
 wire \Tile_X4Y8_FrameStrobe_O[16] ;
 wire \Tile_X4Y8_FrameStrobe_O[17] ;
 wire \Tile_X4Y8_FrameStrobe_O[18] ;
 wire \Tile_X4Y8_FrameStrobe_O[19] ;
 wire \Tile_X4Y8_FrameStrobe_O[1] ;
 wire \Tile_X4Y8_FrameStrobe_O[2] ;
 wire \Tile_X4Y8_FrameStrobe_O[3] ;
 wire \Tile_X4Y8_FrameStrobe_O[4] ;
 wire \Tile_X4Y8_FrameStrobe_O[5] ;
 wire \Tile_X4Y8_FrameStrobe_O[6] ;
 wire \Tile_X4Y8_FrameStrobe_O[7] ;
 wire \Tile_X4Y8_FrameStrobe_O[8] ;
 wire \Tile_X4Y8_FrameStrobe_O[9] ;
 wire \Tile_X4Y8_N1BEG[0] ;
 wire \Tile_X4Y8_N1BEG[1] ;
 wire \Tile_X4Y8_N1BEG[2] ;
 wire \Tile_X4Y8_N1BEG[3] ;
 wire \Tile_X4Y8_N2BEG[0] ;
 wire \Tile_X4Y8_N2BEG[1] ;
 wire \Tile_X4Y8_N2BEG[2] ;
 wire \Tile_X4Y8_N2BEG[3] ;
 wire \Tile_X4Y8_N2BEG[4] ;
 wire \Tile_X4Y8_N2BEG[5] ;
 wire \Tile_X4Y8_N2BEG[6] ;
 wire \Tile_X4Y8_N2BEG[7] ;
 wire \Tile_X4Y8_N2BEGb[0] ;
 wire \Tile_X4Y8_N2BEGb[1] ;
 wire \Tile_X4Y8_N2BEGb[2] ;
 wire \Tile_X4Y8_N2BEGb[3] ;
 wire \Tile_X4Y8_N2BEGb[4] ;
 wire \Tile_X4Y8_N2BEGb[5] ;
 wire \Tile_X4Y8_N2BEGb[6] ;
 wire \Tile_X4Y8_N2BEGb[7] ;
 wire \Tile_X4Y8_N4BEG[0] ;
 wire \Tile_X4Y8_N4BEG[10] ;
 wire \Tile_X4Y8_N4BEG[11] ;
 wire \Tile_X4Y8_N4BEG[12] ;
 wire \Tile_X4Y8_N4BEG[13] ;
 wire \Tile_X4Y8_N4BEG[14] ;
 wire \Tile_X4Y8_N4BEG[15] ;
 wire \Tile_X4Y8_N4BEG[1] ;
 wire \Tile_X4Y8_N4BEG[2] ;
 wire \Tile_X4Y8_N4BEG[3] ;
 wire \Tile_X4Y8_N4BEG[4] ;
 wire \Tile_X4Y8_N4BEG[5] ;
 wire \Tile_X4Y8_N4BEG[6] ;
 wire \Tile_X4Y8_N4BEG[7] ;
 wire \Tile_X4Y8_N4BEG[8] ;
 wire \Tile_X4Y8_N4BEG[9] ;
 wire \Tile_X4Y8_NN4BEG[0] ;
 wire \Tile_X4Y8_NN4BEG[10] ;
 wire \Tile_X4Y8_NN4BEG[11] ;
 wire \Tile_X4Y8_NN4BEG[12] ;
 wire \Tile_X4Y8_NN4BEG[13] ;
 wire \Tile_X4Y8_NN4BEG[14] ;
 wire \Tile_X4Y8_NN4BEG[15] ;
 wire \Tile_X4Y8_NN4BEG[1] ;
 wire \Tile_X4Y8_NN4BEG[2] ;
 wire \Tile_X4Y8_NN4BEG[3] ;
 wire \Tile_X4Y8_NN4BEG[4] ;
 wire \Tile_X4Y8_NN4BEG[5] ;
 wire \Tile_X4Y8_NN4BEG[6] ;
 wire \Tile_X4Y8_NN4BEG[7] ;
 wire \Tile_X4Y8_NN4BEG[8] ;
 wire \Tile_X4Y8_NN4BEG[9] ;
 wire \Tile_X4Y8_S1BEG[0] ;
 wire \Tile_X4Y8_S1BEG[1] ;
 wire \Tile_X4Y8_S1BEG[2] ;
 wire \Tile_X4Y8_S1BEG[3] ;
 wire \Tile_X4Y8_S2BEG[0] ;
 wire \Tile_X4Y8_S2BEG[1] ;
 wire \Tile_X4Y8_S2BEG[2] ;
 wire \Tile_X4Y8_S2BEG[3] ;
 wire \Tile_X4Y8_S2BEG[4] ;
 wire \Tile_X4Y8_S2BEG[5] ;
 wire \Tile_X4Y8_S2BEG[6] ;
 wire \Tile_X4Y8_S2BEG[7] ;
 wire \Tile_X4Y8_S2BEGb[0] ;
 wire \Tile_X4Y8_S2BEGb[1] ;
 wire \Tile_X4Y8_S2BEGb[2] ;
 wire \Tile_X4Y8_S2BEGb[3] ;
 wire \Tile_X4Y8_S2BEGb[4] ;
 wire \Tile_X4Y8_S2BEGb[5] ;
 wire \Tile_X4Y8_S2BEGb[6] ;
 wire \Tile_X4Y8_S2BEGb[7] ;
 wire \Tile_X4Y8_S4BEG[0] ;
 wire \Tile_X4Y8_S4BEG[10] ;
 wire \Tile_X4Y8_S4BEG[11] ;
 wire \Tile_X4Y8_S4BEG[12] ;
 wire \Tile_X4Y8_S4BEG[13] ;
 wire \Tile_X4Y8_S4BEG[14] ;
 wire \Tile_X4Y8_S4BEG[15] ;
 wire \Tile_X4Y8_S4BEG[1] ;
 wire \Tile_X4Y8_S4BEG[2] ;
 wire \Tile_X4Y8_S4BEG[3] ;
 wire \Tile_X4Y8_S4BEG[4] ;
 wire \Tile_X4Y8_S4BEG[5] ;
 wire \Tile_X4Y8_S4BEG[6] ;
 wire \Tile_X4Y8_S4BEG[7] ;
 wire \Tile_X4Y8_S4BEG[8] ;
 wire \Tile_X4Y8_S4BEG[9] ;
 wire \Tile_X4Y8_SS4BEG[0] ;
 wire \Tile_X4Y8_SS4BEG[10] ;
 wire \Tile_X4Y8_SS4BEG[11] ;
 wire \Tile_X4Y8_SS4BEG[12] ;
 wire \Tile_X4Y8_SS4BEG[13] ;
 wire \Tile_X4Y8_SS4BEG[14] ;
 wire \Tile_X4Y8_SS4BEG[15] ;
 wire \Tile_X4Y8_SS4BEG[1] ;
 wire \Tile_X4Y8_SS4BEG[2] ;
 wire \Tile_X4Y8_SS4BEG[3] ;
 wire \Tile_X4Y8_SS4BEG[4] ;
 wire \Tile_X4Y8_SS4BEG[5] ;
 wire \Tile_X4Y8_SS4BEG[6] ;
 wire \Tile_X4Y8_SS4BEG[7] ;
 wire \Tile_X4Y8_SS4BEG[8] ;
 wire \Tile_X4Y8_SS4BEG[9] ;
 wire Tile_X4Y8_UserCLKo;
 wire \Tile_X4Y8_W1BEG[0] ;
 wire \Tile_X4Y8_W1BEG[1] ;
 wire \Tile_X4Y8_W1BEG[2] ;
 wire \Tile_X4Y8_W1BEG[3] ;
 wire \Tile_X4Y8_W2BEG[0] ;
 wire \Tile_X4Y8_W2BEG[1] ;
 wire \Tile_X4Y8_W2BEG[2] ;
 wire \Tile_X4Y8_W2BEG[3] ;
 wire \Tile_X4Y8_W2BEG[4] ;
 wire \Tile_X4Y8_W2BEG[5] ;
 wire \Tile_X4Y8_W2BEG[6] ;
 wire \Tile_X4Y8_W2BEG[7] ;
 wire \Tile_X4Y8_W2BEGb[0] ;
 wire \Tile_X4Y8_W2BEGb[1] ;
 wire \Tile_X4Y8_W2BEGb[2] ;
 wire \Tile_X4Y8_W2BEGb[3] ;
 wire \Tile_X4Y8_W2BEGb[4] ;
 wire \Tile_X4Y8_W2BEGb[5] ;
 wire \Tile_X4Y8_W2BEGb[6] ;
 wire \Tile_X4Y8_W2BEGb[7] ;
 wire \Tile_X4Y8_W6BEG[0] ;
 wire \Tile_X4Y8_W6BEG[10] ;
 wire \Tile_X4Y8_W6BEG[11] ;
 wire \Tile_X4Y8_W6BEG[1] ;
 wire \Tile_X4Y8_W6BEG[2] ;
 wire \Tile_X4Y8_W6BEG[3] ;
 wire \Tile_X4Y8_W6BEG[4] ;
 wire \Tile_X4Y8_W6BEG[5] ;
 wire \Tile_X4Y8_W6BEG[6] ;
 wire \Tile_X4Y8_W6BEG[7] ;
 wire \Tile_X4Y8_W6BEG[8] ;
 wire \Tile_X4Y8_W6BEG[9] ;
 wire \Tile_X4Y8_WW4BEG[0] ;
 wire \Tile_X4Y8_WW4BEG[10] ;
 wire \Tile_X4Y8_WW4BEG[11] ;
 wire \Tile_X4Y8_WW4BEG[12] ;
 wire \Tile_X4Y8_WW4BEG[13] ;
 wire \Tile_X4Y8_WW4BEG[14] ;
 wire \Tile_X4Y8_WW4BEG[15] ;
 wire \Tile_X4Y8_WW4BEG[1] ;
 wire \Tile_X4Y8_WW4BEG[2] ;
 wire \Tile_X4Y8_WW4BEG[3] ;
 wire \Tile_X4Y8_WW4BEG[4] ;
 wire \Tile_X4Y8_WW4BEG[5] ;
 wire \Tile_X4Y8_WW4BEG[6] ;
 wire \Tile_X4Y8_WW4BEG[7] ;
 wire \Tile_X4Y8_WW4BEG[8] ;
 wire \Tile_X4Y8_WW4BEG[9] ;
 wire Tile_X4Y9_Co;
 wire \Tile_X4Y9_FrameData_O[0] ;
 wire \Tile_X4Y9_FrameData_O[10] ;
 wire \Tile_X4Y9_FrameData_O[11] ;
 wire \Tile_X4Y9_FrameData_O[12] ;
 wire \Tile_X4Y9_FrameData_O[13] ;
 wire \Tile_X4Y9_FrameData_O[14] ;
 wire \Tile_X4Y9_FrameData_O[15] ;
 wire \Tile_X4Y9_FrameData_O[16] ;
 wire \Tile_X4Y9_FrameData_O[17] ;
 wire \Tile_X4Y9_FrameData_O[18] ;
 wire \Tile_X4Y9_FrameData_O[19] ;
 wire \Tile_X4Y9_FrameData_O[1] ;
 wire \Tile_X4Y9_FrameData_O[20] ;
 wire \Tile_X4Y9_FrameData_O[21] ;
 wire \Tile_X4Y9_FrameData_O[22] ;
 wire \Tile_X4Y9_FrameData_O[23] ;
 wire \Tile_X4Y9_FrameData_O[24] ;
 wire \Tile_X4Y9_FrameData_O[25] ;
 wire \Tile_X4Y9_FrameData_O[26] ;
 wire \Tile_X4Y9_FrameData_O[27] ;
 wire \Tile_X4Y9_FrameData_O[28] ;
 wire \Tile_X4Y9_FrameData_O[29] ;
 wire \Tile_X4Y9_FrameData_O[2] ;
 wire \Tile_X4Y9_FrameData_O[30] ;
 wire \Tile_X4Y9_FrameData_O[31] ;
 wire \Tile_X4Y9_FrameData_O[3] ;
 wire \Tile_X4Y9_FrameData_O[4] ;
 wire \Tile_X4Y9_FrameData_O[5] ;
 wire \Tile_X4Y9_FrameData_O[6] ;
 wire \Tile_X4Y9_FrameData_O[7] ;
 wire \Tile_X4Y9_FrameData_O[8] ;
 wire \Tile_X4Y9_FrameData_O[9] ;
 wire \Tile_X4Y9_FrameStrobe_O[0] ;
 wire \Tile_X4Y9_FrameStrobe_O[10] ;
 wire \Tile_X4Y9_FrameStrobe_O[11] ;
 wire \Tile_X4Y9_FrameStrobe_O[12] ;
 wire \Tile_X4Y9_FrameStrobe_O[13] ;
 wire \Tile_X4Y9_FrameStrobe_O[14] ;
 wire \Tile_X4Y9_FrameStrobe_O[15] ;
 wire \Tile_X4Y9_FrameStrobe_O[16] ;
 wire \Tile_X4Y9_FrameStrobe_O[17] ;
 wire \Tile_X4Y9_FrameStrobe_O[18] ;
 wire \Tile_X4Y9_FrameStrobe_O[19] ;
 wire \Tile_X4Y9_FrameStrobe_O[1] ;
 wire \Tile_X4Y9_FrameStrobe_O[2] ;
 wire \Tile_X4Y9_FrameStrobe_O[3] ;
 wire \Tile_X4Y9_FrameStrobe_O[4] ;
 wire \Tile_X4Y9_FrameStrobe_O[5] ;
 wire \Tile_X4Y9_FrameStrobe_O[6] ;
 wire \Tile_X4Y9_FrameStrobe_O[7] ;
 wire \Tile_X4Y9_FrameStrobe_O[8] ;
 wire \Tile_X4Y9_FrameStrobe_O[9] ;
 wire \Tile_X4Y9_N1BEG[0] ;
 wire \Tile_X4Y9_N1BEG[1] ;
 wire \Tile_X4Y9_N1BEG[2] ;
 wire \Tile_X4Y9_N1BEG[3] ;
 wire \Tile_X4Y9_N2BEG[0] ;
 wire \Tile_X4Y9_N2BEG[1] ;
 wire \Tile_X4Y9_N2BEG[2] ;
 wire \Tile_X4Y9_N2BEG[3] ;
 wire \Tile_X4Y9_N2BEG[4] ;
 wire \Tile_X4Y9_N2BEG[5] ;
 wire \Tile_X4Y9_N2BEG[6] ;
 wire \Tile_X4Y9_N2BEG[7] ;
 wire \Tile_X4Y9_N2BEGb[0] ;
 wire \Tile_X4Y9_N2BEGb[1] ;
 wire \Tile_X4Y9_N2BEGb[2] ;
 wire \Tile_X4Y9_N2BEGb[3] ;
 wire \Tile_X4Y9_N2BEGb[4] ;
 wire \Tile_X4Y9_N2BEGb[5] ;
 wire \Tile_X4Y9_N2BEGb[6] ;
 wire \Tile_X4Y9_N2BEGb[7] ;
 wire \Tile_X4Y9_N4BEG[0] ;
 wire \Tile_X4Y9_N4BEG[10] ;
 wire \Tile_X4Y9_N4BEG[11] ;
 wire \Tile_X4Y9_N4BEG[12] ;
 wire \Tile_X4Y9_N4BEG[13] ;
 wire \Tile_X4Y9_N4BEG[14] ;
 wire \Tile_X4Y9_N4BEG[15] ;
 wire \Tile_X4Y9_N4BEG[1] ;
 wire \Tile_X4Y9_N4BEG[2] ;
 wire \Tile_X4Y9_N4BEG[3] ;
 wire \Tile_X4Y9_N4BEG[4] ;
 wire \Tile_X4Y9_N4BEG[5] ;
 wire \Tile_X4Y9_N4BEG[6] ;
 wire \Tile_X4Y9_N4BEG[7] ;
 wire \Tile_X4Y9_N4BEG[8] ;
 wire \Tile_X4Y9_N4BEG[9] ;
 wire \Tile_X4Y9_NN4BEG[0] ;
 wire \Tile_X4Y9_NN4BEG[10] ;
 wire \Tile_X4Y9_NN4BEG[11] ;
 wire \Tile_X4Y9_NN4BEG[12] ;
 wire \Tile_X4Y9_NN4BEG[13] ;
 wire \Tile_X4Y9_NN4BEG[14] ;
 wire \Tile_X4Y9_NN4BEG[15] ;
 wire \Tile_X4Y9_NN4BEG[1] ;
 wire \Tile_X4Y9_NN4BEG[2] ;
 wire \Tile_X4Y9_NN4BEG[3] ;
 wire \Tile_X4Y9_NN4BEG[4] ;
 wire \Tile_X4Y9_NN4BEG[5] ;
 wire \Tile_X4Y9_NN4BEG[6] ;
 wire \Tile_X4Y9_NN4BEG[7] ;
 wire \Tile_X4Y9_NN4BEG[8] ;
 wire \Tile_X4Y9_NN4BEG[9] ;
 wire Tile_X4Y9_UserCLKo;
 wire \Tile_X5Y0_FrameData_O[0] ;
 wire \Tile_X5Y0_FrameData_O[10] ;
 wire \Tile_X5Y0_FrameData_O[11] ;
 wire \Tile_X5Y0_FrameData_O[12] ;
 wire \Tile_X5Y0_FrameData_O[13] ;
 wire \Tile_X5Y0_FrameData_O[14] ;
 wire \Tile_X5Y0_FrameData_O[15] ;
 wire \Tile_X5Y0_FrameData_O[16] ;
 wire \Tile_X5Y0_FrameData_O[17] ;
 wire \Tile_X5Y0_FrameData_O[18] ;
 wire \Tile_X5Y0_FrameData_O[19] ;
 wire \Tile_X5Y0_FrameData_O[1] ;
 wire \Tile_X5Y0_FrameData_O[20] ;
 wire \Tile_X5Y0_FrameData_O[21] ;
 wire \Tile_X5Y0_FrameData_O[22] ;
 wire \Tile_X5Y0_FrameData_O[23] ;
 wire \Tile_X5Y0_FrameData_O[24] ;
 wire \Tile_X5Y0_FrameData_O[25] ;
 wire \Tile_X5Y0_FrameData_O[26] ;
 wire \Tile_X5Y0_FrameData_O[27] ;
 wire \Tile_X5Y0_FrameData_O[28] ;
 wire \Tile_X5Y0_FrameData_O[29] ;
 wire \Tile_X5Y0_FrameData_O[2] ;
 wire \Tile_X5Y0_FrameData_O[30] ;
 wire \Tile_X5Y0_FrameData_O[31] ;
 wire \Tile_X5Y0_FrameData_O[3] ;
 wire \Tile_X5Y0_FrameData_O[4] ;
 wire \Tile_X5Y0_FrameData_O[5] ;
 wire \Tile_X5Y0_FrameData_O[6] ;
 wire \Tile_X5Y0_FrameData_O[7] ;
 wire \Tile_X5Y0_FrameData_O[8] ;
 wire \Tile_X5Y0_FrameData_O[9] ;
 wire \Tile_X5Y0_FrameStrobe_O[0] ;
 wire \Tile_X5Y0_FrameStrobe_O[10] ;
 wire \Tile_X5Y0_FrameStrobe_O[11] ;
 wire \Tile_X5Y0_FrameStrobe_O[12] ;
 wire \Tile_X5Y0_FrameStrobe_O[13] ;
 wire \Tile_X5Y0_FrameStrobe_O[14] ;
 wire \Tile_X5Y0_FrameStrobe_O[15] ;
 wire \Tile_X5Y0_FrameStrobe_O[16] ;
 wire \Tile_X5Y0_FrameStrobe_O[17] ;
 wire \Tile_X5Y0_FrameStrobe_O[18] ;
 wire \Tile_X5Y0_FrameStrobe_O[19] ;
 wire \Tile_X5Y0_FrameStrobe_O[1] ;
 wire \Tile_X5Y0_FrameStrobe_O[2] ;
 wire \Tile_X5Y0_FrameStrobe_O[3] ;
 wire \Tile_X5Y0_FrameStrobe_O[4] ;
 wire \Tile_X5Y0_FrameStrobe_O[5] ;
 wire \Tile_X5Y0_FrameStrobe_O[6] ;
 wire \Tile_X5Y0_FrameStrobe_O[7] ;
 wire \Tile_X5Y0_FrameStrobe_O[8] ;
 wire \Tile_X5Y0_FrameStrobe_O[9] ;
 wire \Tile_X5Y0_S1BEG[0] ;
 wire \Tile_X5Y0_S1BEG[1] ;
 wire \Tile_X5Y0_S1BEG[2] ;
 wire \Tile_X5Y0_S1BEG[3] ;
 wire \Tile_X5Y0_S2BEG[0] ;
 wire \Tile_X5Y0_S2BEG[1] ;
 wire \Tile_X5Y0_S2BEG[2] ;
 wire \Tile_X5Y0_S2BEG[3] ;
 wire \Tile_X5Y0_S2BEG[4] ;
 wire \Tile_X5Y0_S2BEG[5] ;
 wire \Tile_X5Y0_S2BEG[6] ;
 wire \Tile_X5Y0_S2BEG[7] ;
 wire \Tile_X5Y0_S2BEGb[0] ;
 wire \Tile_X5Y0_S2BEGb[1] ;
 wire \Tile_X5Y0_S2BEGb[2] ;
 wire \Tile_X5Y0_S2BEGb[3] ;
 wire \Tile_X5Y0_S2BEGb[4] ;
 wire \Tile_X5Y0_S2BEGb[5] ;
 wire \Tile_X5Y0_S2BEGb[6] ;
 wire \Tile_X5Y0_S2BEGb[7] ;
 wire \Tile_X5Y0_S4BEG[0] ;
 wire \Tile_X5Y0_S4BEG[10] ;
 wire \Tile_X5Y0_S4BEG[11] ;
 wire \Tile_X5Y0_S4BEG[12] ;
 wire \Tile_X5Y0_S4BEG[13] ;
 wire \Tile_X5Y0_S4BEG[14] ;
 wire \Tile_X5Y0_S4BEG[15] ;
 wire \Tile_X5Y0_S4BEG[1] ;
 wire \Tile_X5Y0_S4BEG[2] ;
 wire \Tile_X5Y0_S4BEG[3] ;
 wire \Tile_X5Y0_S4BEG[4] ;
 wire \Tile_X5Y0_S4BEG[5] ;
 wire \Tile_X5Y0_S4BEG[6] ;
 wire \Tile_X5Y0_S4BEG[7] ;
 wire \Tile_X5Y0_S4BEG[8] ;
 wire \Tile_X5Y0_S4BEG[9] ;
 wire Tile_X5Y0_UserCLKo;
 wire \Tile_X5Y1_FrameData_O[0] ;
 wire \Tile_X5Y1_FrameData_O[10] ;
 wire \Tile_X5Y1_FrameData_O[11] ;
 wire \Tile_X5Y1_FrameData_O[12] ;
 wire \Tile_X5Y1_FrameData_O[13] ;
 wire \Tile_X5Y1_FrameData_O[14] ;
 wire \Tile_X5Y1_FrameData_O[15] ;
 wire \Tile_X5Y1_FrameData_O[16] ;
 wire \Tile_X5Y1_FrameData_O[17] ;
 wire \Tile_X5Y1_FrameData_O[18] ;
 wire \Tile_X5Y1_FrameData_O[19] ;
 wire \Tile_X5Y1_FrameData_O[1] ;
 wire \Tile_X5Y1_FrameData_O[20] ;
 wire \Tile_X5Y1_FrameData_O[21] ;
 wire \Tile_X5Y1_FrameData_O[22] ;
 wire \Tile_X5Y1_FrameData_O[23] ;
 wire \Tile_X5Y1_FrameData_O[24] ;
 wire \Tile_X5Y1_FrameData_O[25] ;
 wire \Tile_X5Y1_FrameData_O[26] ;
 wire \Tile_X5Y1_FrameData_O[27] ;
 wire \Tile_X5Y1_FrameData_O[28] ;
 wire \Tile_X5Y1_FrameData_O[29] ;
 wire \Tile_X5Y1_FrameData_O[2] ;
 wire \Tile_X5Y1_FrameData_O[30] ;
 wire \Tile_X5Y1_FrameData_O[31] ;
 wire \Tile_X5Y1_FrameData_O[3] ;
 wire \Tile_X5Y1_FrameData_O[4] ;
 wire \Tile_X5Y1_FrameData_O[5] ;
 wire \Tile_X5Y1_FrameData_O[6] ;
 wire \Tile_X5Y1_FrameData_O[7] ;
 wire \Tile_X5Y1_FrameData_O[8] ;
 wire \Tile_X5Y1_FrameData_O[9] ;
 wire \Tile_X5Y1_FrameStrobe_O[0] ;
 wire \Tile_X5Y1_FrameStrobe_O[10] ;
 wire \Tile_X5Y1_FrameStrobe_O[11] ;
 wire \Tile_X5Y1_FrameStrobe_O[12] ;
 wire \Tile_X5Y1_FrameStrobe_O[13] ;
 wire \Tile_X5Y1_FrameStrobe_O[14] ;
 wire \Tile_X5Y1_FrameStrobe_O[15] ;
 wire \Tile_X5Y1_FrameStrobe_O[16] ;
 wire \Tile_X5Y1_FrameStrobe_O[17] ;
 wire \Tile_X5Y1_FrameStrobe_O[18] ;
 wire \Tile_X5Y1_FrameStrobe_O[19] ;
 wire \Tile_X5Y1_FrameStrobe_O[1] ;
 wire \Tile_X5Y1_FrameStrobe_O[2] ;
 wire \Tile_X5Y1_FrameStrobe_O[3] ;
 wire \Tile_X5Y1_FrameStrobe_O[4] ;
 wire \Tile_X5Y1_FrameStrobe_O[5] ;
 wire \Tile_X5Y1_FrameStrobe_O[6] ;
 wire \Tile_X5Y1_FrameStrobe_O[7] ;
 wire \Tile_X5Y1_FrameStrobe_O[8] ;
 wire \Tile_X5Y1_FrameStrobe_O[9] ;
 wire \Tile_X5Y1_N1BEG[0] ;
 wire \Tile_X5Y1_N1BEG[1] ;
 wire \Tile_X5Y1_N1BEG[2] ;
 wire \Tile_X5Y1_N1BEG[3] ;
 wire \Tile_X5Y1_N2BEG[0] ;
 wire \Tile_X5Y1_N2BEG[1] ;
 wire \Tile_X5Y1_N2BEG[2] ;
 wire \Tile_X5Y1_N2BEG[3] ;
 wire \Tile_X5Y1_N2BEG[4] ;
 wire \Tile_X5Y1_N2BEG[5] ;
 wire \Tile_X5Y1_N2BEG[6] ;
 wire \Tile_X5Y1_N2BEG[7] ;
 wire \Tile_X5Y1_N2BEGb[0] ;
 wire \Tile_X5Y1_N2BEGb[1] ;
 wire \Tile_X5Y1_N2BEGb[2] ;
 wire \Tile_X5Y1_N2BEGb[3] ;
 wire \Tile_X5Y1_N2BEGb[4] ;
 wire \Tile_X5Y1_N2BEGb[5] ;
 wire \Tile_X5Y1_N2BEGb[6] ;
 wire \Tile_X5Y1_N2BEGb[7] ;
 wire \Tile_X5Y1_N4BEG[0] ;
 wire \Tile_X5Y1_N4BEG[10] ;
 wire \Tile_X5Y1_N4BEG[11] ;
 wire \Tile_X5Y1_N4BEG[12] ;
 wire \Tile_X5Y1_N4BEG[13] ;
 wire \Tile_X5Y1_N4BEG[14] ;
 wire \Tile_X5Y1_N4BEG[15] ;
 wire \Tile_X5Y1_N4BEG[1] ;
 wire \Tile_X5Y1_N4BEG[2] ;
 wire \Tile_X5Y1_N4BEG[3] ;
 wire \Tile_X5Y1_N4BEG[4] ;
 wire \Tile_X5Y1_N4BEG[5] ;
 wire \Tile_X5Y1_N4BEG[6] ;
 wire \Tile_X5Y1_N4BEG[7] ;
 wire \Tile_X5Y1_N4BEG[8] ;
 wire \Tile_X5Y1_N4BEG[9] ;
 wire Tile_X5Y1_UserCLKo;
 wire \Tile_X5Y1_W1BEG[0] ;
 wire \Tile_X5Y1_W1BEG[1] ;
 wire \Tile_X5Y1_W1BEG[2] ;
 wire \Tile_X5Y1_W1BEG[3] ;
 wire \Tile_X5Y1_W2BEG[0] ;
 wire \Tile_X5Y1_W2BEG[1] ;
 wire \Tile_X5Y1_W2BEG[2] ;
 wire \Tile_X5Y1_W2BEG[3] ;
 wire \Tile_X5Y1_W2BEG[4] ;
 wire \Tile_X5Y1_W2BEG[5] ;
 wire \Tile_X5Y1_W2BEG[6] ;
 wire \Tile_X5Y1_W2BEG[7] ;
 wire \Tile_X5Y1_W2BEGb[0] ;
 wire \Tile_X5Y1_W2BEGb[1] ;
 wire \Tile_X5Y1_W2BEGb[2] ;
 wire \Tile_X5Y1_W2BEGb[3] ;
 wire \Tile_X5Y1_W2BEGb[4] ;
 wire \Tile_X5Y1_W2BEGb[5] ;
 wire \Tile_X5Y1_W2BEGb[6] ;
 wire \Tile_X5Y1_W2BEGb[7] ;
 wire \Tile_X5Y1_W6BEG[0] ;
 wire \Tile_X5Y1_W6BEG[10] ;
 wire \Tile_X5Y1_W6BEG[11] ;
 wire \Tile_X5Y1_W6BEG[1] ;
 wire \Tile_X5Y1_W6BEG[2] ;
 wire \Tile_X5Y1_W6BEG[3] ;
 wire \Tile_X5Y1_W6BEG[4] ;
 wire \Tile_X5Y1_W6BEG[5] ;
 wire \Tile_X5Y1_W6BEG[6] ;
 wire \Tile_X5Y1_W6BEG[7] ;
 wire \Tile_X5Y1_W6BEG[8] ;
 wire \Tile_X5Y1_W6BEG[9] ;
 wire \Tile_X5Y1_WW4BEG[0] ;
 wire \Tile_X5Y1_WW4BEG[10] ;
 wire \Tile_X5Y1_WW4BEG[11] ;
 wire \Tile_X5Y1_WW4BEG[12] ;
 wire \Tile_X5Y1_WW4BEG[13] ;
 wire \Tile_X5Y1_WW4BEG[14] ;
 wire \Tile_X5Y1_WW4BEG[15] ;
 wire \Tile_X5Y1_WW4BEG[1] ;
 wire \Tile_X5Y1_WW4BEG[2] ;
 wire \Tile_X5Y1_WW4BEG[3] ;
 wire \Tile_X5Y1_WW4BEG[4] ;
 wire \Tile_X5Y1_WW4BEG[5] ;
 wire \Tile_X5Y1_WW4BEG[6] ;
 wire \Tile_X5Y1_WW4BEG[7] ;
 wire \Tile_X5Y1_WW4BEG[8] ;
 wire \Tile_X5Y1_WW4BEG[9] ;
 wire \Tile_X5Y2_FrameData_O[0] ;
 wire \Tile_X5Y2_FrameData_O[10] ;
 wire \Tile_X5Y2_FrameData_O[11] ;
 wire \Tile_X5Y2_FrameData_O[12] ;
 wire \Tile_X5Y2_FrameData_O[13] ;
 wire \Tile_X5Y2_FrameData_O[14] ;
 wire \Tile_X5Y2_FrameData_O[15] ;
 wire \Tile_X5Y2_FrameData_O[16] ;
 wire \Tile_X5Y2_FrameData_O[17] ;
 wire \Tile_X5Y2_FrameData_O[18] ;
 wire \Tile_X5Y2_FrameData_O[19] ;
 wire \Tile_X5Y2_FrameData_O[1] ;
 wire \Tile_X5Y2_FrameData_O[20] ;
 wire \Tile_X5Y2_FrameData_O[21] ;
 wire \Tile_X5Y2_FrameData_O[22] ;
 wire \Tile_X5Y2_FrameData_O[23] ;
 wire \Tile_X5Y2_FrameData_O[24] ;
 wire \Tile_X5Y2_FrameData_O[25] ;
 wire \Tile_X5Y2_FrameData_O[26] ;
 wire \Tile_X5Y2_FrameData_O[27] ;
 wire \Tile_X5Y2_FrameData_O[28] ;
 wire \Tile_X5Y2_FrameData_O[29] ;
 wire \Tile_X5Y2_FrameData_O[2] ;
 wire \Tile_X5Y2_FrameData_O[30] ;
 wire \Tile_X5Y2_FrameData_O[31] ;
 wire \Tile_X5Y2_FrameData_O[3] ;
 wire \Tile_X5Y2_FrameData_O[4] ;
 wire \Tile_X5Y2_FrameData_O[5] ;
 wire \Tile_X5Y2_FrameData_O[6] ;
 wire \Tile_X5Y2_FrameData_O[7] ;
 wire \Tile_X5Y2_FrameData_O[8] ;
 wire \Tile_X5Y2_FrameData_O[9] ;
 wire \Tile_X5Y2_S1BEG[0] ;
 wire \Tile_X5Y2_S1BEG[1] ;
 wire \Tile_X5Y2_S1BEG[2] ;
 wire \Tile_X5Y2_S1BEG[3] ;
 wire \Tile_X5Y2_S2BEG[0] ;
 wire \Tile_X5Y2_S2BEG[1] ;
 wire \Tile_X5Y2_S2BEG[2] ;
 wire \Tile_X5Y2_S2BEG[3] ;
 wire \Tile_X5Y2_S2BEG[4] ;
 wire \Tile_X5Y2_S2BEG[5] ;
 wire \Tile_X5Y2_S2BEG[6] ;
 wire \Tile_X5Y2_S2BEG[7] ;
 wire \Tile_X5Y2_S2BEGb[0] ;
 wire \Tile_X5Y2_S2BEGb[1] ;
 wire \Tile_X5Y2_S2BEGb[2] ;
 wire \Tile_X5Y2_S2BEGb[3] ;
 wire \Tile_X5Y2_S2BEGb[4] ;
 wire \Tile_X5Y2_S2BEGb[5] ;
 wire \Tile_X5Y2_S2BEGb[6] ;
 wire \Tile_X5Y2_S2BEGb[7] ;
 wire \Tile_X5Y2_S4BEG[0] ;
 wire \Tile_X5Y2_S4BEG[10] ;
 wire \Tile_X5Y2_S4BEG[11] ;
 wire \Tile_X5Y2_S4BEG[12] ;
 wire \Tile_X5Y2_S4BEG[13] ;
 wire \Tile_X5Y2_S4BEG[14] ;
 wire \Tile_X5Y2_S4BEG[15] ;
 wire \Tile_X5Y2_S4BEG[1] ;
 wire \Tile_X5Y2_S4BEG[2] ;
 wire \Tile_X5Y2_S4BEG[3] ;
 wire \Tile_X5Y2_S4BEG[4] ;
 wire \Tile_X5Y2_S4BEG[5] ;
 wire \Tile_X5Y2_S4BEG[6] ;
 wire \Tile_X5Y2_S4BEG[7] ;
 wire \Tile_X5Y2_S4BEG[8] ;
 wire \Tile_X5Y2_S4BEG[9] ;
 wire \Tile_X5Y2_W1BEG[0] ;
 wire \Tile_X5Y2_W1BEG[1] ;
 wire \Tile_X5Y2_W1BEG[2] ;
 wire \Tile_X5Y2_W1BEG[3] ;
 wire \Tile_X5Y2_W2BEG[0] ;
 wire \Tile_X5Y2_W2BEG[1] ;
 wire \Tile_X5Y2_W2BEG[2] ;
 wire \Tile_X5Y2_W2BEG[3] ;
 wire \Tile_X5Y2_W2BEG[4] ;
 wire \Tile_X5Y2_W2BEG[5] ;
 wire \Tile_X5Y2_W2BEG[6] ;
 wire \Tile_X5Y2_W2BEG[7] ;
 wire \Tile_X5Y2_W2BEGb[0] ;
 wire \Tile_X5Y2_W2BEGb[1] ;
 wire \Tile_X5Y2_W2BEGb[2] ;
 wire \Tile_X5Y2_W2BEGb[3] ;
 wire \Tile_X5Y2_W2BEGb[4] ;
 wire \Tile_X5Y2_W2BEGb[5] ;
 wire \Tile_X5Y2_W2BEGb[6] ;
 wire \Tile_X5Y2_W2BEGb[7] ;
 wire \Tile_X5Y2_W6BEG[0] ;
 wire \Tile_X5Y2_W6BEG[10] ;
 wire \Tile_X5Y2_W6BEG[11] ;
 wire \Tile_X5Y2_W6BEG[1] ;
 wire \Tile_X5Y2_W6BEG[2] ;
 wire \Tile_X5Y2_W6BEG[3] ;
 wire \Tile_X5Y2_W6BEG[4] ;
 wire \Tile_X5Y2_W6BEG[5] ;
 wire \Tile_X5Y2_W6BEG[6] ;
 wire \Tile_X5Y2_W6BEG[7] ;
 wire \Tile_X5Y2_W6BEG[8] ;
 wire \Tile_X5Y2_W6BEG[9] ;
 wire \Tile_X5Y2_WW4BEG[0] ;
 wire \Tile_X5Y2_WW4BEG[10] ;
 wire \Tile_X5Y2_WW4BEG[11] ;
 wire \Tile_X5Y2_WW4BEG[12] ;
 wire \Tile_X5Y2_WW4BEG[13] ;
 wire \Tile_X5Y2_WW4BEG[14] ;
 wire \Tile_X5Y2_WW4BEG[15] ;
 wire \Tile_X5Y2_WW4BEG[1] ;
 wire \Tile_X5Y2_WW4BEG[2] ;
 wire \Tile_X5Y2_WW4BEG[3] ;
 wire \Tile_X5Y2_WW4BEG[4] ;
 wire \Tile_X5Y2_WW4BEG[5] ;
 wire \Tile_X5Y2_WW4BEG[6] ;
 wire \Tile_X5Y2_WW4BEG[7] ;
 wire \Tile_X5Y2_WW4BEG[8] ;
 wire \Tile_X5Y2_WW4BEG[9] ;
 wire \Tile_X5Y3_FrameData_O[0] ;
 wire \Tile_X5Y3_FrameData_O[10] ;
 wire \Tile_X5Y3_FrameData_O[11] ;
 wire \Tile_X5Y3_FrameData_O[12] ;
 wire \Tile_X5Y3_FrameData_O[13] ;
 wire \Tile_X5Y3_FrameData_O[14] ;
 wire \Tile_X5Y3_FrameData_O[15] ;
 wire \Tile_X5Y3_FrameData_O[16] ;
 wire \Tile_X5Y3_FrameData_O[17] ;
 wire \Tile_X5Y3_FrameData_O[18] ;
 wire \Tile_X5Y3_FrameData_O[19] ;
 wire \Tile_X5Y3_FrameData_O[1] ;
 wire \Tile_X5Y3_FrameData_O[20] ;
 wire \Tile_X5Y3_FrameData_O[21] ;
 wire \Tile_X5Y3_FrameData_O[22] ;
 wire \Tile_X5Y3_FrameData_O[23] ;
 wire \Tile_X5Y3_FrameData_O[24] ;
 wire \Tile_X5Y3_FrameData_O[25] ;
 wire \Tile_X5Y3_FrameData_O[26] ;
 wire \Tile_X5Y3_FrameData_O[27] ;
 wire \Tile_X5Y3_FrameData_O[28] ;
 wire \Tile_X5Y3_FrameData_O[29] ;
 wire \Tile_X5Y3_FrameData_O[2] ;
 wire \Tile_X5Y3_FrameData_O[30] ;
 wire \Tile_X5Y3_FrameData_O[31] ;
 wire \Tile_X5Y3_FrameData_O[3] ;
 wire \Tile_X5Y3_FrameData_O[4] ;
 wire \Tile_X5Y3_FrameData_O[5] ;
 wire \Tile_X5Y3_FrameData_O[6] ;
 wire \Tile_X5Y3_FrameData_O[7] ;
 wire \Tile_X5Y3_FrameData_O[8] ;
 wire \Tile_X5Y3_FrameData_O[9] ;
 wire \Tile_X5Y3_FrameStrobe_O[0] ;
 wire \Tile_X5Y3_FrameStrobe_O[10] ;
 wire \Tile_X5Y3_FrameStrobe_O[11] ;
 wire \Tile_X5Y3_FrameStrobe_O[12] ;
 wire \Tile_X5Y3_FrameStrobe_O[13] ;
 wire \Tile_X5Y3_FrameStrobe_O[14] ;
 wire \Tile_X5Y3_FrameStrobe_O[15] ;
 wire \Tile_X5Y3_FrameStrobe_O[16] ;
 wire \Tile_X5Y3_FrameStrobe_O[17] ;
 wire \Tile_X5Y3_FrameStrobe_O[18] ;
 wire \Tile_X5Y3_FrameStrobe_O[19] ;
 wire \Tile_X5Y3_FrameStrobe_O[1] ;
 wire \Tile_X5Y3_FrameStrobe_O[2] ;
 wire \Tile_X5Y3_FrameStrobe_O[3] ;
 wire \Tile_X5Y3_FrameStrobe_O[4] ;
 wire \Tile_X5Y3_FrameStrobe_O[5] ;
 wire \Tile_X5Y3_FrameStrobe_O[6] ;
 wire \Tile_X5Y3_FrameStrobe_O[7] ;
 wire \Tile_X5Y3_FrameStrobe_O[8] ;
 wire \Tile_X5Y3_FrameStrobe_O[9] ;
 wire \Tile_X5Y3_N1BEG[0] ;
 wire \Tile_X5Y3_N1BEG[1] ;
 wire \Tile_X5Y3_N1BEG[2] ;
 wire \Tile_X5Y3_N1BEG[3] ;
 wire \Tile_X5Y3_N2BEG[0] ;
 wire \Tile_X5Y3_N2BEG[1] ;
 wire \Tile_X5Y3_N2BEG[2] ;
 wire \Tile_X5Y3_N2BEG[3] ;
 wire \Tile_X5Y3_N2BEG[4] ;
 wire \Tile_X5Y3_N2BEG[5] ;
 wire \Tile_X5Y3_N2BEG[6] ;
 wire \Tile_X5Y3_N2BEG[7] ;
 wire \Tile_X5Y3_N2BEGb[0] ;
 wire \Tile_X5Y3_N2BEGb[1] ;
 wire \Tile_X5Y3_N2BEGb[2] ;
 wire \Tile_X5Y3_N2BEGb[3] ;
 wire \Tile_X5Y3_N2BEGb[4] ;
 wire \Tile_X5Y3_N2BEGb[5] ;
 wire \Tile_X5Y3_N2BEGb[6] ;
 wire \Tile_X5Y3_N2BEGb[7] ;
 wire \Tile_X5Y3_N4BEG[0] ;
 wire \Tile_X5Y3_N4BEG[10] ;
 wire \Tile_X5Y3_N4BEG[11] ;
 wire \Tile_X5Y3_N4BEG[12] ;
 wire \Tile_X5Y3_N4BEG[13] ;
 wire \Tile_X5Y3_N4BEG[14] ;
 wire \Tile_X5Y3_N4BEG[15] ;
 wire \Tile_X5Y3_N4BEG[1] ;
 wire \Tile_X5Y3_N4BEG[2] ;
 wire \Tile_X5Y3_N4BEG[3] ;
 wire \Tile_X5Y3_N4BEG[4] ;
 wire \Tile_X5Y3_N4BEG[5] ;
 wire \Tile_X5Y3_N4BEG[6] ;
 wire \Tile_X5Y3_N4BEG[7] ;
 wire \Tile_X5Y3_N4BEG[8] ;
 wire \Tile_X5Y3_N4BEG[9] ;
 wire Tile_X5Y3_UserCLKo;
 wire \Tile_X5Y3_W1BEG[0] ;
 wire \Tile_X5Y3_W1BEG[1] ;
 wire \Tile_X5Y3_W1BEG[2] ;
 wire \Tile_X5Y3_W1BEG[3] ;
 wire \Tile_X5Y3_W2BEG[0] ;
 wire \Tile_X5Y3_W2BEG[1] ;
 wire \Tile_X5Y3_W2BEG[2] ;
 wire \Tile_X5Y3_W2BEG[3] ;
 wire \Tile_X5Y3_W2BEG[4] ;
 wire \Tile_X5Y3_W2BEG[5] ;
 wire \Tile_X5Y3_W2BEG[6] ;
 wire \Tile_X5Y3_W2BEG[7] ;
 wire \Tile_X5Y3_W2BEGb[0] ;
 wire \Tile_X5Y3_W2BEGb[1] ;
 wire \Tile_X5Y3_W2BEGb[2] ;
 wire \Tile_X5Y3_W2BEGb[3] ;
 wire \Tile_X5Y3_W2BEGb[4] ;
 wire \Tile_X5Y3_W2BEGb[5] ;
 wire \Tile_X5Y3_W2BEGb[6] ;
 wire \Tile_X5Y3_W2BEGb[7] ;
 wire \Tile_X5Y3_W6BEG[0] ;
 wire \Tile_X5Y3_W6BEG[10] ;
 wire \Tile_X5Y3_W6BEG[11] ;
 wire \Tile_X5Y3_W6BEG[1] ;
 wire \Tile_X5Y3_W6BEG[2] ;
 wire \Tile_X5Y3_W6BEG[3] ;
 wire \Tile_X5Y3_W6BEG[4] ;
 wire \Tile_X5Y3_W6BEG[5] ;
 wire \Tile_X5Y3_W6BEG[6] ;
 wire \Tile_X5Y3_W6BEG[7] ;
 wire \Tile_X5Y3_W6BEG[8] ;
 wire \Tile_X5Y3_W6BEG[9] ;
 wire \Tile_X5Y3_WW4BEG[0] ;
 wire \Tile_X5Y3_WW4BEG[10] ;
 wire \Tile_X5Y3_WW4BEG[11] ;
 wire \Tile_X5Y3_WW4BEG[12] ;
 wire \Tile_X5Y3_WW4BEG[13] ;
 wire \Tile_X5Y3_WW4BEG[14] ;
 wire \Tile_X5Y3_WW4BEG[15] ;
 wire \Tile_X5Y3_WW4BEG[1] ;
 wire \Tile_X5Y3_WW4BEG[2] ;
 wire \Tile_X5Y3_WW4BEG[3] ;
 wire \Tile_X5Y3_WW4BEG[4] ;
 wire \Tile_X5Y3_WW4BEG[5] ;
 wire \Tile_X5Y3_WW4BEG[6] ;
 wire \Tile_X5Y3_WW4BEG[7] ;
 wire \Tile_X5Y3_WW4BEG[8] ;
 wire \Tile_X5Y3_WW4BEG[9] ;
 wire \Tile_X5Y4_FrameData_O[0] ;
 wire \Tile_X5Y4_FrameData_O[10] ;
 wire \Tile_X5Y4_FrameData_O[11] ;
 wire \Tile_X5Y4_FrameData_O[12] ;
 wire \Tile_X5Y4_FrameData_O[13] ;
 wire \Tile_X5Y4_FrameData_O[14] ;
 wire \Tile_X5Y4_FrameData_O[15] ;
 wire \Tile_X5Y4_FrameData_O[16] ;
 wire \Tile_X5Y4_FrameData_O[17] ;
 wire \Tile_X5Y4_FrameData_O[18] ;
 wire \Tile_X5Y4_FrameData_O[19] ;
 wire \Tile_X5Y4_FrameData_O[1] ;
 wire \Tile_X5Y4_FrameData_O[20] ;
 wire \Tile_X5Y4_FrameData_O[21] ;
 wire \Tile_X5Y4_FrameData_O[22] ;
 wire \Tile_X5Y4_FrameData_O[23] ;
 wire \Tile_X5Y4_FrameData_O[24] ;
 wire \Tile_X5Y4_FrameData_O[25] ;
 wire \Tile_X5Y4_FrameData_O[26] ;
 wire \Tile_X5Y4_FrameData_O[27] ;
 wire \Tile_X5Y4_FrameData_O[28] ;
 wire \Tile_X5Y4_FrameData_O[29] ;
 wire \Tile_X5Y4_FrameData_O[2] ;
 wire \Tile_X5Y4_FrameData_O[30] ;
 wire \Tile_X5Y4_FrameData_O[31] ;
 wire \Tile_X5Y4_FrameData_O[3] ;
 wire \Tile_X5Y4_FrameData_O[4] ;
 wire \Tile_X5Y4_FrameData_O[5] ;
 wire \Tile_X5Y4_FrameData_O[6] ;
 wire \Tile_X5Y4_FrameData_O[7] ;
 wire \Tile_X5Y4_FrameData_O[8] ;
 wire \Tile_X5Y4_FrameData_O[9] ;
 wire \Tile_X5Y4_S1BEG[0] ;
 wire \Tile_X5Y4_S1BEG[1] ;
 wire \Tile_X5Y4_S1BEG[2] ;
 wire \Tile_X5Y4_S1BEG[3] ;
 wire \Tile_X5Y4_S2BEG[0] ;
 wire \Tile_X5Y4_S2BEG[1] ;
 wire \Tile_X5Y4_S2BEG[2] ;
 wire \Tile_X5Y4_S2BEG[3] ;
 wire \Tile_X5Y4_S2BEG[4] ;
 wire \Tile_X5Y4_S2BEG[5] ;
 wire \Tile_X5Y4_S2BEG[6] ;
 wire \Tile_X5Y4_S2BEG[7] ;
 wire \Tile_X5Y4_S2BEGb[0] ;
 wire \Tile_X5Y4_S2BEGb[1] ;
 wire \Tile_X5Y4_S2BEGb[2] ;
 wire \Tile_X5Y4_S2BEGb[3] ;
 wire \Tile_X5Y4_S2BEGb[4] ;
 wire \Tile_X5Y4_S2BEGb[5] ;
 wire \Tile_X5Y4_S2BEGb[6] ;
 wire \Tile_X5Y4_S2BEGb[7] ;
 wire \Tile_X5Y4_S4BEG[0] ;
 wire \Tile_X5Y4_S4BEG[10] ;
 wire \Tile_X5Y4_S4BEG[11] ;
 wire \Tile_X5Y4_S4BEG[12] ;
 wire \Tile_X5Y4_S4BEG[13] ;
 wire \Tile_X5Y4_S4BEG[14] ;
 wire \Tile_X5Y4_S4BEG[15] ;
 wire \Tile_X5Y4_S4BEG[1] ;
 wire \Tile_X5Y4_S4BEG[2] ;
 wire \Tile_X5Y4_S4BEG[3] ;
 wire \Tile_X5Y4_S4BEG[4] ;
 wire \Tile_X5Y4_S4BEG[5] ;
 wire \Tile_X5Y4_S4BEG[6] ;
 wire \Tile_X5Y4_S4BEG[7] ;
 wire \Tile_X5Y4_S4BEG[8] ;
 wire \Tile_X5Y4_S4BEG[9] ;
 wire \Tile_X5Y4_W1BEG[0] ;
 wire \Tile_X5Y4_W1BEG[1] ;
 wire \Tile_X5Y4_W1BEG[2] ;
 wire \Tile_X5Y4_W1BEG[3] ;
 wire \Tile_X5Y4_W2BEG[0] ;
 wire \Tile_X5Y4_W2BEG[1] ;
 wire \Tile_X5Y4_W2BEG[2] ;
 wire \Tile_X5Y4_W2BEG[3] ;
 wire \Tile_X5Y4_W2BEG[4] ;
 wire \Tile_X5Y4_W2BEG[5] ;
 wire \Tile_X5Y4_W2BEG[6] ;
 wire \Tile_X5Y4_W2BEG[7] ;
 wire \Tile_X5Y4_W2BEGb[0] ;
 wire \Tile_X5Y4_W2BEGb[1] ;
 wire \Tile_X5Y4_W2BEGb[2] ;
 wire \Tile_X5Y4_W2BEGb[3] ;
 wire \Tile_X5Y4_W2BEGb[4] ;
 wire \Tile_X5Y4_W2BEGb[5] ;
 wire \Tile_X5Y4_W2BEGb[6] ;
 wire \Tile_X5Y4_W2BEGb[7] ;
 wire \Tile_X5Y4_W6BEG[0] ;
 wire \Tile_X5Y4_W6BEG[10] ;
 wire \Tile_X5Y4_W6BEG[11] ;
 wire \Tile_X5Y4_W6BEG[1] ;
 wire \Tile_X5Y4_W6BEG[2] ;
 wire \Tile_X5Y4_W6BEG[3] ;
 wire \Tile_X5Y4_W6BEG[4] ;
 wire \Tile_X5Y4_W6BEG[5] ;
 wire \Tile_X5Y4_W6BEG[6] ;
 wire \Tile_X5Y4_W6BEG[7] ;
 wire \Tile_X5Y4_W6BEG[8] ;
 wire \Tile_X5Y4_W6BEG[9] ;
 wire \Tile_X5Y4_WW4BEG[0] ;
 wire \Tile_X5Y4_WW4BEG[10] ;
 wire \Tile_X5Y4_WW4BEG[11] ;
 wire \Tile_X5Y4_WW4BEG[12] ;
 wire \Tile_X5Y4_WW4BEG[13] ;
 wire \Tile_X5Y4_WW4BEG[14] ;
 wire \Tile_X5Y4_WW4BEG[15] ;
 wire \Tile_X5Y4_WW4BEG[1] ;
 wire \Tile_X5Y4_WW4BEG[2] ;
 wire \Tile_X5Y4_WW4BEG[3] ;
 wire \Tile_X5Y4_WW4BEG[4] ;
 wire \Tile_X5Y4_WW4BEG[5] ;
 wire \Tile_X5Y4_WW4BEG[6] ;
 wire \Tile_X5Y4_WW4BEG[7] ;
 wire \Tile_X5Y4_WW4BEG[8] ;
 wire \Tile_X5Y4_WW4BEG[9] ;
 wire \Tile_X5Y5_FrameData_O[0] ;
 wire \Tile_X5Y5_FrameData_O[10] ;
 wire \Tile_X5Y5_FrameData_O[11] ;
 wire \Tile_X5Y5_FrameData_O[12] ;
 wire \Tile_X5Y5_FrameData_O[13] ;
 wire \Tile_X5Y5_FrameData_O[14] ;
 wire \Tile_X5Y5_FrameData_O[15] ;
 wire \Tile_X5Y5_FrameData_O[16] ;
 wire \Tile_X5Y5_FrameData_O[17] ;
 wire \Tile_X5Y5_FrameData_O[18] ;
 wire \Tile_X5Y5_FrameData_O[19] ;
 wire \Tile_X5Y5_FrameData_O[1] ;
 wire \Tile_X5Y5_FrameData_O[20] ;
 wire \Tile_X5Y5_FrameData_O[21] ;
 wire \Tile_X5Y5_FrameData_O[22] ;
 wire \Tile_X5Y5_FrameData_O[23] ;
 wire \Tile_X5Y5_FrameData_O[24] ;
 wire \Tile_X5Y5_FrameData_O[25] ;
 wire \Tile_X5Y5_FrameData_O[26] ;
 wire \Tile_X5Y5_FrameData_O[27] ;
 wire \Tile_X5Y5_FrameData_O[28] ;
 wire \Tile_X5Y5_FrameData_O[29] ;
 wire \Tile_X5Y5_FrameData_O[2] ;
 wire \Tile_X5Y5_FrameData_O[30] ;
 wire \Tile_X5Y5_FrameData_O[31] ;
 wire \Tile_X5Y5_FrameData_O[3] ;
 wire \Tile_X5Y5_FrameData_O[4] ;
 wire \Tile_X5Y5_FrameData_O[5] ;
 wire \Tile_X5Y5_FrameData_O[6] ;
 wire \Tile_X5Y5_FrameData_O[7] ;
 wire \Tile_X5Y5_FrameData_O[8] ;
 wire \Tile_X5Y5_FrameData_O[9] ;
 wire \Tile_X5Y5_FrameStrobe_O[0] ;
 wire \Tile_X5Y5_FrameStrobe_O[10] ;
 wire \Tile_X5Y5_FrameStrobe_O[11] ;
 wire \Tile_X5Y5_FrameStrobe_O[12] ;
 wire \Tile_X5Y5_FrameStrobe_O[13] ;
 wire \Tile_X5Y5_FrameStrobe_O[14] ;
 wire \Tile_X5Y5_FrameStrobe_O[15] ;
 wire \Tile_X5Y5_FrameStrobe_O[16] ;
 wire \Tile_X5Y5_FrameStrobe_O[17] ;
 wire \Tile_X5Y5_FrameStrobe_O[18] ;
 wire \Tile_X5Y5_FrameStrobe_O[19] ;
 wire \Tile_X5Y5_FrameStrobe_O[1] ;
 wire \Tile_X5Y5_FrameStrobe_O[2] ;
 wire \Tile_X5Y5_FrameStrobe_O[3] ;
 wire \Tile_X5Y5_FrameStrobe_O[4] ;
 wire \Tile_X5Y5_FrameStrobe_O[5] ;
 wire \Tile_X5Y5_FrameStrobe_O[6] ;
 wire \Tile_X5Y5_FrameStrobe_O[7] ;
 wire \Tile_X5Y5_FrameStrobe_O[8] ;
 wire \Tile_X5Y5_FrameStrobe_O[9] ;
 wire \Tile_X5Y5_N1BEG[0] ;
 wire \Tile_X5Y5_N1BEG[1] ;
 wire \Tile_X5Y5_N1BEG[2] ;
 wire \Tile_X5Y5_N1BEG[3] ;
 wire \Tile_X5Y5_N2BEG[0] ;
 wire \Tile_X5Y5_N2BEG[1] ;
 wire \Tile_X5Y5_N2BEG[2] ;
 wire \Tile_X5Y5_N2BEG[3] ;
 wire \Tile_X5Y5_N2BEG[4] ;
 wire \Tile_X5Y5_N2BEG[5] ;
 wire \Tile_X5Y5_N2BEG[6] ;
 wire \Tile_X5Y5_N2BEG[7] ;
 wire \Tile_X5Y5_N2BEGb[0] ;
 wire \Tile_X5Y5_N2BEGb[1] ;
 wire \Tile_X5Y5_N2BEGb[2] ;
 wire \Tile_X5Y5_N2BEGb[3] ;
 wire \Tile_X5Y5_N2BEGb[4] ;
 wire \Tile_X5Y5_N2BEGb[5] ;
 wire \Tile_X5Y5_N2BEGb[6] ;
 wire \Tile_X5Y5_N2BEGb[7] ;
 wire \Tile_X5Y5_N4BEG[0] ;
 wire \Tile_X5Y5_N4BEG[10] ;
 wire \Tile_X5Y5_N4BEG[11] ;
 wire \Tile_X5Y5_N4BEG[12] ;
 wire \Tile_X5Y5_N4BEG[13] ;
 wire \Tile_X5Y5_N4BEG[14] ;
 wire \Tile_X5Y5_N4BEG[15] ;
 wire \Tile_X5Y5_N4BEG[1] ;
 wire \Tile_X5Y5_N4BEG[2] ;
 wire \Tile_X5Y5_N4BEG[3] ;
 wire \Tile_X5Y5_N4BEG[4] ;
 wire \Tile_X5Y5_N4BEG[5] ;
 wire \Tile_X5Y5_N4BEG[6] ;
 wire \Tile_X5Y5_N4BEG[7] ;
 wire \Tile_X5Y5_N4BEG[8] ;
 wire \Tile_X5Y5_N4BEG[9] ;
 wire \Tile_X5Y5_S1BEG[0] ;
 wire \Tile_X5Y5_S1BEG[1] ;
 wire \Tile_X5Y5_S1BEG[2] ;
 wire \Tile_X5Y5_S1BEG[3] ;
 wire \Tile_X5Y5_S2BEG[0] ;
 wire \Tile_X5Y5_S2BEG[1] ;
 wire \Tile_X5Y5_S2BEG[2] ;
 wire \Tile_X5Y5_S2BEG[3] ;
 wire \Tile_X5Y5_S2BEG[4] ;
 wire \Tile_X5Y5_S2BEG[5] ;
 wire \Tile_X5Y5_S2BEG[6] ;
 wire \Tile_X5Y5_S2BEG[7] ;
 wire \Tile_X5Y5_S2BEGb[0] ;
 wire \Tile_X5Y5_S2BEGb[1] ;
 wire \Tile_X5Y5_S2BEGb[2] ;
 wire \Tile_X5Y5_S2BEGb[3] ;
 wire \Tile_X5Y5_S2BEGb[4] ;
 wire \Tile_X5Y5_S2BEGb[5] ;
 wire \Tile_X5Y5_S2BEGb[6] ;
 wire \Tile_X5Y5_S2BEGb[7] ;
 wire \Tile_X5Y5_S4BEG[0] ;
 wire \Tile_X5Y5_S4BEG[10] ;
 wire \Tile_X5Y5_S4BEG[11] ;
 wire \Tile_X5Y5_S4BEG[12] ;
 wire \Tile_X5Y5_S4BEG[13] ;
 wire \Tile_X5Y5_S4BEG[14] ;
 wire \Tile_X5Y5_S4BEG[15] ;
 wire \Tile_X5Y5_S4BEG[1] ;
 wire \Tile_X5Y5_S4BEG[2] ;
 wire \Tile_X5Y5_S4BEG[3] ;
 wire \Tile_X5Y5_S4BEG[4] ;
 wire \Tile_X5Y5_S4BEG[5] ;
 wire \Tile_X5Y5_S4BEG[6] ;
 wire \Tile_X5Y5_S4BEG[7] ;
 wire \Tile_X5Y5_S4BEG[8] ;
 wire \Tile_X5Y5_S4BEG[9] ;
 wire Tile_X5Y5_UserCLKo;
 wire \Tile_X5Y5_W1BEG[0] ;
 wire \Tile_X5Y5_W1BEG[1] ;
 wire \Tile_X5Y5_W1BEG[2] ;
 wire \Tile_X5Y5_W1BEG[3] ;
 wire \Tile_X5Y5_W2BEG[0] ;
 wire \Tile_X5Y5_W2BEG[1] ;
 wire \Tile_X5Y5_W2BEG[2] ;
 wire \Tile_X5Y5_W2BEG[3] ;
 wire \Tile_X5Y5_W2BEG[4] ;
 wire \Tile_X5Y5_W2BEG[5] ;
 wire \Tile_X5Y5_W2BEG[6] ;
 wire \Tile_X5Y5_W2BEG[7] ;
 wire \Tile_X5Y5_W2BEGb[0] ;
 wire \Tile_X5Y5_W2BEGb[1] ;
 wire \Tile_X5Y5_W2BEGb[2] ;
 wire \Tile_X5Y5_W2BEGb[3] ;
 wire \Tile_X5Y5_W2BEGb[4] ;
 wire \Tile_X5Y5_W2BEGb[5] ;
 wire \Tile_X5Y5_W2BEGb[6] ;
 wire \Tile_X5Y5_W2BEGb[7] ;
 wire \Tile_X5Y5_W6BEG[0] ;
 wire \Tile_X5Y5_W6BEG[10] ;
 wire \Tile_X5Y5_W6BEG[11] ;
 wire \Tile_X5Y5_W6BEG[1] ;
 wire \Tile_X5Y5_W6BEG[2] ;
 wire \Tile_X5Y5_W6BEG[3] ;
 wire \Tile_X5Y5_W6BEG[4] ;
 wire \Tile_X5Y5_W6BEG[5] ;
 wire \Tile_X5Y5_W6BEG[6] ;
 wire \Tile_X5Y5_W6BEG[7] ;
 wire \Tile_X5Y5_W6BEG[8] ;
 wire \Tile_X5Y5_W6BEG[9] ;
 wire \Tile_X5Y5_WW4BEG[0] ;
 wire \Tile_X5Y5_WW4BEG[10] ;
 wire \Tile_X5Y5_WW4BEG[11] ;
 wire \Tile_X5Y5_WW4BEG[12] ;
 wire \Tile_X5Y5_WW4BEG[13] ;
 wire \Tile_X5Y5_WW4BEG[14] ;
 wire \Tile_X5Y5_WW4BEG[15] ;
 wire \Tile_X5Y5_WW4BEG[1] ;
 wire \Tile_X5Y5_WW4BEG[2] ;
 wire \Tile_X5Y5_WW4BEG[3] ;
 wire \Tile_X5Y5_WW4BEG[4] ;
 wire \Tile_X5Y5_WW4BEG[5] ;
 wire \Tile_X5Y5_WW4BEG[6] ;
 wire \Tile_X5Y5_WW4BEG[7] ;
 wire \Tile_X5Y5_WW4BEG[8] ;
 wire \Tile_X5Y5_WW4BEG[9] ;
 wire \Tile_X5Y6_FrameData_O[0] ;
 wire \Tile_X5Y6_FrameData_O[10] ;
 wire \Tile_X5Y6_FrameData_O[11] ;
 wire \Tile_X5Y6_FrameData_O[12] ;
 wire \Tile_X5Y6_FrameData_O[13] ;
 wire \Tile_X5Y6_FrameData_O[14] ;
 wire \Tile_X5Y6_FrameData_O[15] ;
 wire \Tile_X5Y6_FrameData_O[16] ;
 wire \Tile_X5Y6_FrameData_O[17] ;
 wire \Tile_X5Y6_FrameData_O[18] ;
 wire \Tile_X5Y6_FrameData_O[19] ;
 wire \Tile_X5Y6_FrameData_O[1] ;
 wire \Tile_X5Y6_FrameData_O[20] ;
 wire \Tile_X5Y6_FrameData_O[21] ;
 wire \Tile_X5Y6_FrameData_O[22] ;
 wire \Tile_X5Y6_FrameData_O[23] ;
 wire \Tile_X5Y6_FrameData_O[24] ;
 wire \Tile_X5Y6_FrameData_O[25] ;
 wire \Tile_X5Y6_FrameData_O[26] ;
 wire \Tile_X5Y6_FrameData_O[27] ;
 wire \Tile_X5Y6_FrameData_O[28] ;
 wire \Tile_X5Y6_FrameData_O[29] ;
 wire \Tile_X5Y6_FrameData_O[2] ;
 wire \Tile_X5Y6_FrameData_O[30] ;
 wire \Tile_X5Y6_FrameData_O[31] ;
 wire \Tile_X5Y6_FrameData_O[3] ;
 wire \Tile_X5Y6_FrameData_O[4] ;
 wire \Tile_X5Y6_FrameData_O[5] ;
 wire \Tile_X5Y6_FrameData_O[6] ;
 wire \Tile_X5Y6_FrameData_O[7] ;
 wire \Tile_X5Y6_FrameData_O[8] ;
 wire \Tile_X5Y6_FrameData_O[9] ;
 wire \Tile_X5Y6_FrameStrobe_O[0] ;
 wire \Tile_X5Y6_FrameStrobe_O[10] ;
 wire \Tile_X5Y6_FrameStrobe_O[11] ;
 wire \Tile_X5Y6_FrameStrobe_O[12] ;
 wire \Tile_X5Y6_FrameStrobe_O[13] ;
 wire \Tile_X5Y6_FrameStrobe_O[14] ;
 wire \Tile_X5Y6_FrameStrobe_O[15] ;
 wire \Tile_X5Y6_FrameStrobe_O[16] ;
 wire \Tile_X5Y6_FrameStrobe_O[17] ;
 wire \Tile_X5Y6_FrameStrobe_O[18] ;
 wire \Tile_X5Y6_FrameStrobe_O[19] ;
 wire \Tile_X5Y6_FrameStrobe_O[1] ;
 wire \Tile_X5Y6_FrameStrobe_O[2] ;
 wire \Tile_X5Y6_FrameStrobe_O[3] ;
 wire \Tile_X5Y6_FrameStrobe_O[4] ;
 wire \Tile_X5Y6_FrameStrobe_O[5] ;
 wire \Tile_X5Y6_FrameStrobe_O[6] ;
 wire \Tile_X5Y6_FrameStrobe_O[7] ;
 wire \Tile_X5Y6_FrameStrobe_O[8] ;
 wire \Tile_X5Y6_FrameStrobe_O[9] ;
 wire \Tile_X5Y6_N1BEG[0] ;
 wire \Tile_X5Y6_N1BEG[1] ;
 wire \Tile_X5Y6_N1BEG[2] ;
 wire \Tile_X5Y6_N1BEG[3] ;
 wire \Tile_X5Y6_N2BEG[0] ;
 wire \Tile_X5Y6_N2BEG[1] ;
 wire \Tile_X5Y6_N2BEG[2] ;
 wire \Tile_X5Y6_N2BEG[3] ;
 wire \Tile_X5Y6_N2BEG[4] ;
 wire \Tile_X5Y6_N2BEG[5] ;
 wire \Tile_X5Y6_N2BEG[6] ;
 wire \Tile_X5Y6_N2BEG[7] ;
 wire \Tile_X5Y6_N2BEGb[0] ;
 wire \Tile_X5Y6_N2BEGb[1] ;
 wire \Tile_X5Y6_N2BEGb[2] ;
 wire \Tile_X5Y6_N2BEGb[3] ;
 wire \Tile_X5Y6_N2BEGb[4] ;
 wire \Tile_X5Y6_N2BEGb[5] ;
 wire \Tile_X5Y6_N2BEGb[6] ;
 wire \Tile_X5Y6_N2BEGb[7] ;
 wire \Tile_X5Y6_N4BEG[0] ;
 wire \Tile_X5Y6_N4BEG[10] ;
 wire \Tile_X5Y6_N4BEG[11] ;
 wire \Tile_X5Y6_N4BEG[12] ;
 wire \Tile_X5Y6_N4BEG[13] ;
 wire \Tile_X5Y6_N4BEG[14] ;
 wire \Tile_X5Y6_N4BEG[15] ;
 wire \Tile_X5Y6_N4BEG[1] ;
 wire \Tile_X5Y6_N4BEG[2] ;
 wire \Tile_X5Y6_N4BEG[3] ;
 wire \Tile_X5Y6_N4BEG[4] ;
 wire \Tile_X5Y6_N4BEG[5] ;
 wire \Tile_X5Y6_N4BEG[6] ;
 wire \Tile_X5Y6_N4BEG[7] ;
 wire \Tile_X5Y6_N4BEG[8] ;
 wire \Tile_X5Y6_N4BEG[9] ;
 wire \Tile_X5Y6_S1BEG[0] ;
 wire \Tile_X5Y6_S1BEG[1] ;
 wire \Tile_X5Y6_S1BEG[2] ;
 wire \Tile_X5Y6_S1BEG[3] ;
 wire \Tile_X5Y6_S2BEG[0] ;
 wire \Tile_X5Y6_S2BEG[1] ;
 wire \Tile_X5Y6_S2BEG[2] ;
 wire \Tile_X5Y6_S2BEG[3] ;
 wire \Tile_X5Y6_S2BEG[4] ;
 wire \Tile_X5Y6_S2BEG[5] ;
 wire \Tile_X5Y6_S2BEG[6] ;
 wire \Tile_X5Y6_S2BEG[7] ;
 wire \Tile_X5Y6_S2BEGb[0] ;
 wire \Tile_X5Y6_S2BEGb[1] ;
 wire \Tile_X5Y6_S2BEGb[2] ;
 wire \Tile_X5Y6_S2BEGb[3] ;
 wire \Tile_X5Y6_S2BEGb[4] ;
 wire \Tile_X5Y6_S2BEGb[5] ;
 wire \Tile_X5Y6_S2BEGb[6] ;
 wire \Tile_X5Y6_S2BEGb[7] ;
 wire \Tile_X5Y6_S4BEG[0] ;
 wire \Tile_X5Y6_S4BEG[10] ;
 wire \Tile_X5Y6_S4BEG[11] ;
 wire \Tile_X5Y6_S4BEG[12] ;
 wire \Tile_X5Y6_S4BEG[13] ;
 wire \Tile_X5Y6_S4BEG[14] ;
 wire \Tile_X5Y6_S4BEG[15] ;
 wire \Tile_X5Y6_S4BEG[1] ;
 wire \Tile_X5Y6_S4BEG[2] ;
 wire \Tile_X5Y6_S4BEG[3] ;
 wire \Tile_X5Y6_S4BEG[4] ;
 wire \Tile_X5Y6_S4BEG[5] ;
 wire \Tile_X5Y6_S4BEG[6] ;
 wire \Tile_X5Y6_S4BEG[7] ;
 wire \Tile_X5Y6_S4BEG[8] ;
 wire \Tile_X5Y6_S4BEG[9] ;
 wire Tile_X5Y6_UserCLKo;
 wire \Tile_X5Y6_W1BEG[0] ;
 wire \Tile_X5Y6_W1BEG[1] ;
 wire \Tile_X5Y6_W1BEG[2] ;
 wire \Tile_X5Y6_W1BEG[3] ;
 wire \Tile_X5Y6_W2BEG[0] ;
 wire \Tile_X5Y6_W2BEG[1] ;
 wire \Tile_X5Y6_W2BEG[2] ;
 wire \Tile_X5Y6_W2BEG[3] ;
 wire \Tile_X5Y6_W2BEG[4] ;
 wire \Tile_X5Y6_W2BEG[5] ;
 wire \Tile_X5Y6_W2BEG[6] ;
 wire \Tile_X5Y6_W2BEG[7] ;
 wire \Tile_X5Y6_W2BEGb[0] ;
 wire \Tile_X5Y6_W2BEGb[1] ;
 wire \Tile_X5Y6_W2BEGb[2] ;
 wire \Tile_X5Y6_W2BEGb[3] ;
 wire \Tile_X5Y6_W2BEGb[4] ;
 wire \Tile_X5Y6_W2BEGb[5] ;
 wire \Tile_X5Y6_W2BEGb[6] ;
 wire \Tile_X5Y6_W2BEGb[7] ;
 wire \Tile_X5Y6_W6BEG[0] ;
 wire \Tile_X5Y6_W6BEG[10] ;
 wire \Tile_X5Y6_W6BEG[11] ;
 wire \Tile_X5Y6_W6BEG[1] ;
 wire \Tile_X5Y6_W6BEG[2] ;
 wire \Tile_X5Y6_W6BEG[3] ;
 wire \Tile_X5Y6_W6BEG[4] ;
 wire \Tile_X5Y6_W6BEG[5] ;
 wire \Tile_X5Y6_W6BEG[6] ;
 wire \Tile_X5Y6_W6BEG[7] ;
 wire \Tile_X5Y6_W6BEG[8] ;
 wire \Tile_X5Y6_W6BEG[9] ;
 wire \Tile_X5Y6_WW4BEG[0] ;
 wire \Tile_X5Y6_WW4BEG[10] ;
 wire \Tile_X5Y6_WW4BEG[11] ;
 wire \Tile_X5Y6_WW4BEG[12] ;
 wire \Tile_X5Y6_WW4BEG[13] ;
 wire \Tile_X5Y6_WW4BEG[14] ;
 wire \Tile_X5Y6_WW4BEG[15] ;
 wire \Tile_X5Y6_WW4BEG[1] ;
 wire \Tile_X5Y6_WW4BEG[2] ;
 wire \Tile_X5Y6_WW4BEG[3] ;
 wire \Tile_X5Y6_WW4BEG[4] ;
 wire \Tile_X5Y6_WW4BEG[5] ;
 wire \Tile_X5Y6_WW4BEG[6] ;
 wire \Tile_X5Y6_WW4BEG[7] ;
 wire \Tile_X5Y6_WW4BEG[8] ;
 wire \Tile_X5Y6_WW4BEG[9] ;
 wire \Tile_X5Y7_FrameData_O[0] ;
 wire \Tile_X5Y7_FrameData_O[10] ;
 wire \Tile_X5Y7_FrameData_O[11] ;
 wire \Tile_X5Y7_FrameData_O[12] ;
 wire \Tile_X5Y7_FrameData_O[13] ;
 wire \Tile_X5Y7_FrameData_O[14] ;
 wire \Tile_X5Y7_FrameData_O[15] ;
 wire \Tile_X5Y7_FrameData_O[16] ;
 wire \Tile_X5Y7_FrameData_O[17] ;
 wire \Tile_X5Y7_FrameData_O[18] ;
 wire \Tile_X5Y7_FrameData_O[19] ;
 wire \Tile_X5Y7_FrameData_O[1] ;
 wire \Tile_X5Y7_FrameData_O[20] ;
 wire \Tile_X5Y7_FrameData_O[21] ;
 wire \Tile_X5Y7_FrameData_O[22] ;
 wire \Tile_X5Y7_FrameData_O[23] ;
 wire \Tile_X5Y7_FrameData_O[24] ;
 wire \Tile_X5Y7_FrameData_O[25] ;
 wire \Tile_X5Y7_FrameData_O[26] ;
 wire \Tile_X5Y7_FrameData_O[27] ;
 wire \Tile_X5Y7_FrameData_O[28] ;
 wire \Tile_X5Y7_FrameData_O[29] ;
 wire \Tile_X5Y7_FrameData_O[2] ;
 wire \Tile_X5Y7_FrameData_O[30] ;
 wire \Tile_X5Y7_FrameData_O[31] ;
 wire \Tile_X5Y7_FrameData_O[3] ;
 wire \Tile_X5Y7_FrameData_O[4] ;
 wire \Tile_X5Y7_FrameData_O[5] ;
 wire \Tile_X5Y7_FrameData_O[6] ;
 wire \Tile_X5Y7_FrameData_O[7] ;
 wire \Tile_X5Y7_FrameData_O[8] ;
 wire \Tile_X5Y7_FrameData_O[9] ;
 wire \Tile_X5Y7_FrameStrobe_O[0] ;
 wire \Tile_X5Y7_FrameStrobe_O[10] ;
 wire \Tile_X5Y7_FrameStrobe_O[11] ;
 wire \Tile_X5Y7_FrameStrobe_O[12] ;
 wire \Tile_X5Y7_FrameStrobe_O[13] ;
 wire \Tile_X5Y7_FrameStrobe_O[14] ;
 wire \Tile_X5Y7_FrameStrobe_O[15] ;
 wire \Tile_X5Y7_FrameStrobe_O[16] ;
 wire \Tile_X5Y7_FrameStrobe_O[17] ;
 wire \Tile_X5Y7_FrameStrobe_O[18] ;
 wire \Tile_X5Y7_FrameStrobe_O[19] ;
 wire \Tile_X5Y7_FrameStrobe_O[1] ;
 wire \Tile_X5Y7_FrameStrobe_O[2] ;
 wire \Tile_X5Y7_FrameStrobe_O[3] ;
 wire \Tile_X5Y7_FrameStrobe_O[4] ;
 wire \Tile_X5Y7_FrameStrobe_O[5] ;
 wire \Tile_X5Y7_FrameStrobe_O[6] ;
 wire \Tile_X5Y7_FrameStrobe_O[7] ;
 wire \Tile_X5Y7_FrameStrobe_O[8] ;
 wire \Tile_X5Y7_FrameStrobe_O[9] ;
 wire \Tile_X5Y7_N1BEG[0] ;
 wire \Tile_X5Y7_N1BEG[1] ;
 wire \Tile_X5Y7_N1BEG[2] ;
 wire \Tile_X5Y7_N1BEG[3] ;
 wire \Tile_X5Y7_N2BEG[0] ;
 wire \Tile_X5Y7_N2BEG[1] ;
 wire \Tile_X5Y7_N2BEG[2] ;
 wire \Tile_X5Y7_N2BEG[3] ;
 wire \Tile_X5Y7_N2BEG[4] ;
 wire \Tile_X5Y7_N2BEG[5] ;
 wire \Tile_X5Y7_N2BEG[6] ;
 wire \Tile_X5Y7_N2BEG[7] ;
 wire \Tile_X5Y7_N2BEGb[0] ;
 wire \Tile_X5Y7_N2BEGb[1] ;
 wire \Tile_X5Y7_N2BEGb[2] ;
 wire \Tile_X5Y7_N2BEGb[3] ;
 wire \Tile_X5Y7_N2BEGb[4] ;
 wire \Tile_X5Y7_N2BEGb[5] ;
 wire \Tile_X5Y7_N2BEGb[6] ;
 wire \Tile_X5Y7_N2BEGb[7] ;
 wire \Tile_X5Y7_N4BEG[0] ;
 wire \Tile_X5Y7_N4BEG[10] ;
 wire \Tile_X5Y7_N4BEG[11] ;
 wire \Tile_X5Y7_N4BEG[12] ;
 wire \Tile_X5Y7_N4BEG[13] ;
 wire \Tile_X5Y7_N4BEG[14] ;
 wire \Tile_X5Y7_N4BEG[15] ;
 wire \Tile_X5Y7_N4BEG[1] ;
 wire \Tile_X5Y7_N4BEG[2] ;
 wire \Tile_X5Y7_N4BEG[3] ;
 wire \Tile_X5Y7_N4BEG[4] ;
 wire \Tile_X5Y7_N4BEG[5] ;
 wire \Tile_X5Y7_N4BEG[6] ;
 wire \Tile_X5Y7_N4BEG[7] ;
 wire \Tile_X5Y7_N4BEG[8] ;
 wire \Tile_X5Y7_N4BEG[9] ;
 wire \Tile_X5Y7_S1BEG[0] ;
 wire \Tile_X5Y7_S1BEG[1] ;
 wire \Tile_X5Y7_S1BEG[2] ;
 wire \Tile_X5Y7_S1BEG[3] ;
 wire \Tile_X5Y7_S2BEG[0] ;
 wire \Tile_X5Y7_S2BEG[1] ;
 wire \Tile_X5Y7_S2BEG[2] ;
 wire \Tile_X5Y7_S2BEG[3] ;
 wire \Tile_X5Y7_S2BEG[4] ;
 wire \Tile_X5Y7_S2BEG[5] ;
 wire \Tile_X5Y7_S2BEG[6] ;
 wire \Tile_X5Y7_S2BEG[7] ;
 wire \Tile_X5Y7_S2BEGb[0] ;
 wire \Tile_X5Y7_S2BEGb[1] ;
 wire \Tile_X5Y7_S2BEGb[2] ;
 wire \Tile_X5Y7_S2BEGb[3] ;
 wire \Tile_X5Y7_S2BEGb[4] ;
 wire \Tile_X5Y7_S2BEGb[5] ;
 wire \Tile_X5Y7_S2BEGb[6] ;
 wire \Tile_X5Y7_S2BEGb[7] ;
 wire \Tile_X5Y7_S4BEG[0] ;
 wire \Tile_X5Y7_S4BEG[10] ;
 wire \Tile_X5Y7_S4BEG[11] ;
 wire \Tile_X5Y7_S4BEG[12] ;
 wire \Tile_X5Y7_S4BEG[13] ;
 wire \Tile_X5Y7_S4BEG[14] ;
 wire \Tile_X5Y7_S4BEG[15] ;
 wire \Tile_X5Y7_S4BEG[1] ;
 wire \Tile_X5Y7_S4BEG[2] ;
 wire \Tile_X5Y7_S4BEG[3] ;
 wire \Tile_X5Y7_S4BEG[4] ;
 wire \Tile_X5Y7_S4BEG[5] ;
 wire \Tile_X5Y7_S4BEG[6] ;
 wire \Tile_X5Y7_S4BEG[7] ;
 wire \Tile_X5Y7_S4BEG[8] ;
 wire \Tile_X5Y7_S4BEG[9] ;
 wire Tile_X5Y7_UserCLKo;
 wire \Tile_X5Y7_W1BEG[0] ;
 wire \Tile_X5Y7_W1BEG[1] ;
 wire \Tile_X5Y7_W1BEG[2] ;
 wire \Tile_X5Y7_W1BEG[3] ;
 wire \Tile_X5Y7_W2BEG[0] ;
 wire \Tile_X5Y7_W2BEG[1] ;
 wire \Tile_X5Y7_W2BEG[2] ;
 wire \Tile_X5Y7_W2BEG[3] ;
 wire \Tile_X5Y7_W2BEG[4] ;
 wire \Tile_X5Y7_W2BEG[5] ;
 wire \Tile_X5Y7_W2BEG[6] ;
 wire \Tile_X5Y7_W2BEG[7] ;
 wire \Tile_X5Y7_W2BEGb[0] ;
 wire \Tile_X5Y7_W2BEGb[1] ;
 wire \Tile_X5Y7_W2BEGb[2] ;
 wire \Tile_X5Y7_W2BEGb[3] ;
 wire \Tile_X5Y7_W2BEGb[4] ;
 wire \Tile_X5Y7_W2BEGb[5] ;
 wire \Tile_X5Y7_W2BEGb[6] ;
 wire \Tile_X5Y7_W2BEGb[7] ;
 wire \Tile_X5Y7_W6BEG[0] ;
 wire \Tile_X5Y7_W6BEG[10] ;
 wire \Tile_X5Y7_W6BEG[11] ;
 wire \Tile_X5Y7_W6BEG[1] ;
 wire \Tile_X5Y7_W6BEG[2] ;
 wire \Tile_X5Y7_W6BEG[3] ;
 wire \Tile_X5Y7_W6BEG[4] ;
 wire \Tile_X5Y7_W6BEG[5] ;
 wire \Tile_X5Y7_W6BEG[6] ;
 wire \Tile_X5Y7_W6BEG[7] ;
 wire \Tile_X5Y7_W6BEG[8] ;
 wire \Tile_X5Y7_W6BEG[9] ;
 wire \Tile_X5Y7_WW4BEG[0] ;
 wire \Tile_X5Y7_WW4BEG[10] ;
 wire \Tile_X5Y7_WW4BEG[11] ;
 wire \Tile_X5Y7_WW4BEG[12] ;
 wire \Tile_X5Y7_WW4BEG[13] ;
 wire \Tile_X5Y7_WW4BEG[14] ;
 wire \Tile_X5Y7_WW4BEG[15] ;
 wire \Tile_X5Y7_WW4BEG[1] ;
 wire \Tile_X5Y7_WW4BEG[2] ;
 wire \Tile_X5Y7_WW4BEG[3] ;
 wire \Tile_X5Y7_WW4BEG[4] ;
 wire \Tile_X5Y7_WW4BEG[5] ;
 wire \Tile_X5Y7_WW4BEG[6] ;
 wire \Tile_X5Y7_WW4BEG[7] ;
 wire \Tile_X5Y7_WW4BEG[8] ;
 wire \Tile_X5Y7_WW4BEG[9] ;
 wire \Tile_X5Y8_FrameData_O[0] ;
 wire \Tile_X5Y8_FrameData_O[10] ;
 wire \Tile_X5Y8_FrameData_O[11] ;
 wire \Tile_X5Y8_FrameData_O[12] ;
 wire \Tile_X5Y8_FrameData_O[13] ;
 wire \Tile_X5Y8_FrameData_O[14] ;
 wire \Tile_X5Y8_FrameData_O[15] ;
 wire \Tile_X5Y8_FrameData_O[16] ;
 wire \Tile_X5Y8_FrameData_O[17] ;
 wire \Tile_X5Y8_FrameData_O[18] ;
 wire \Tile_X5Y8_FrameData_O[19] ;
 wire \Tile_X5Y8_FrameData_O[1] ;
 wire \Tile_X5Y8_FrameData_O[20] ;
 wire \Tile_X5Y8_FrameData_O[21] ;
 wire \Tile_X5Y8_FrameData_O[22] ;
 wire \Tile_X5Y8_FrameData_O[23] ;
 wire \Tile_X5Y8_FrameData_O[24] ;
 wire \Tile_X5Y8_FrameData_O[25] ;
 wire \Tile_X5Y8_FrameData_O[26] ;
 wire \Tile_X5Y8_FrameData_O[27] ;
 wire \Tile_X5Y8_FrameData_O[28] ;
 wire \Tile_X5Y8_FrameData_O[29] ;
 wire \Tile_X5Y8_FrameData_O[2] ;
 wire \Tile_X5Y8_FrameData_O[30] ;
 wire \Tile_X5Y8_FrameData_O[31] ;
 wire \Tile_X5Y8_FrameData_O[3] ;
 wire \Tile_X5Y8_FrameData_O[4] ;
 wire \Tile_X5Y8_FrameData_O[5] ;
 wire \Tile_X5Y8_FrameData_O[6] ;
 wire \Tile_X5Y8_FrameData_O[7] ;
 wire \Tile_X5Y8_FrameData_O[8] ;
 wire \Tile_X5Y8_FrameData_O[9] ;
 wire \Tile_X5Y8_FrameStrobe_O[0] ;
 wire \Tile_X5Y8_FrameStrobe_O[10] ;
 wire \Tile_X5Y8_FrameStrobe_O[11] ;
 wire \Tile_X5Y8_FrameStrobe_O[12] ;
 wire \Tile_X5Y8_FrameStrobe_O[13] ;
 wire \Tile_X5Y8_FrameStrobe_O[14] ;
 wire \Tile_X5Y8_FrameStrobe_O[15] ;
 wire \Tile_X5Y8_FrameStrobe_O[16] ;
 wire \Tile_X5Y8_FrameStrobe_O[17] ;
 wire \Tile_X5Y8_FrameStrobe_O[18] ;
 wire \Tile_X5Y8_FrameStrobe_O[19] ;
 wire \Tile_X5Y8_FrameStrobe_O[1] ;
 wire \Tile_X5Y8_FrameStrobe_O[2] ;
 wire \Tile_X5Y8_FrameStrobe_O[3] ;
 wire \Tile_X5Y8_FrameStrobe_O[4] ;
 wire \Tile_X5Y8_FrameStrobe_O[5] ;
 wire \Tile_X5Y8_FrameStrobe_O[6] ;
 wire \Tile_X5Y8_FrameStrobe_O[7] ;
 wire \Tile_X5Y8_FrameStrobe_O[8] ;
 wire \Tile_X5Y8_FrameStrobe_O[9] ;
 wire \Tile_X5Y8_N1BEG[0] ;
 wire \Tile_X5Y8_N1BEG[1] ;
 wire \Tile_X5Y8_N1BEG[2] ;
 wire \Tile_X5Y8_N1BEG[3] ;
 wire \Tile_X5Y8_N2BEG[0] ;
 wire \Tile_X5Y8_N2BEG[1] ;
 wire \Tile_X5Y8_N2BEG[2] ;
 wire \Tile_X5Y8_N2BEG[3] ;
 wire \Tile_X5Y8_N2BEG[4] ;
 wire \Tile_X5Y8_N2BEG[5] ;
 wire \Tile_X5Y8_N2BEG[6] ;
 wire \Tile_X5Y8_N2BEG[7] ;
 wire \Tile_X5Y8_N2BEGb[0] ;
 wire \Tile_X5Y8_N2BEGb[1] ;
 wire \Tile_X5Y8_N2BEGb[2] ;
 wire \Tile_X5Y8_N2BEGb[3] ;
 wire \Tile_X5Y8_N2BEGb[4] ;
 wire \Tile_X5Y8_N2BEGb[5] ;
 wire \Tile_X5Y8_N2BEGb[6] ;
 wire \Tile_X5Y8_N2BEGb[7] ;
 wire \Tile_X5Y8_N4BEG[0] ;
 wire \Tile_X5Y8_N4BEG[10] ;
 wire \Tile_X5Y8_N4BEG[11] ;
 wire \Tile_X5Y8_N4BEG[12] ;
 wire \Tile_X5Y8_N4BEG[13] ;
 wire \Tile_X5Y8_N4BEG[14] ;
 wire \Tile_X5Y8_N4BEG[15] ;
 wire \Tile_X5Y8_N4BEG[1] ;
 wire \Tile_X5Y8_N4BEG[2] ;
 wire \Tile_X5Y8_N4BEG[3] ;
 wire \Tile_X5Y8_N4BEG[4] ;
 wire \Tile_X5Y8_N4BEG[5] ;
 wire \Tile_X5Y8_N4BEG[6] ;
 wire \Tile_X5Y8_N4BEG[7] ;
 wire \Tile_X5Y8_N4BEG[8] ;
 wire \Tile_X5Y8_N4BEG[9] ;
 wire \Tile_X5Y8_S1BEG[0] ;
 wire \Tile_X5Y8_S1BEG[1] ;
 wire \Tile_X5Y8_S1BEG[2] ;
 wire \Tile_X5Y8_S1BEG[3] ;
 wire \Tile_X5Y8_S2BEG[0] ;
 wire \Tile_X5Y8_S2BEG[1] ;
 wire \Tile_X5Y8_S2BEG[2] ;
 wire \Tile_X5Y8_S2BEG[3] ;
 wire \Tile_X5Y8_S2BEG[4] ;
 wire \Tile_X5Y8_S2BEG[5] ;
 wire \Tile_X5Y8_S2BEG[6] ;
 wire \Tile_X5Y8_S2BEG[7] ;
 wire \Tile_X5Y8_S2BEGb[0] ;
 wire \Tile_X5Y8_S2BEGb[1] ;
 wire \Tile_X5Y8_S2BEGb[2] ;
 wire \Tile_X5Y8_S2BEGb[3] ;
 wire \Tile_X5Y8_S2BEGb[4] ;
 wire \Tile_X5Y8_S2BEGb[5] ;
 wire \Tile_X5Y8_S2BEGb[6] ;
 wire \Tile_X5Y8_S2BEGb[7] ;
 wire \Tile_X5Y8_S4BEG[0] ;
 wire \Tile_X5Y8_S4BEG[10] ;
 wire \Tile_X5Y8_S4BEG[11] ;
 wire \Tile_X5Y8_S4BEG[12] ;
 wire \Tile_X5Y8_S4BEG[13] ;
 wire \Tile_X5Y8_S4BEG[14] ;
 wire \Tile_X5Y8_S4BEG[15] ;
 wire \Tile_X5Y8_S4BEG[1] ;
 wire \Tile_X5Y8_S4BEG[2] ;
 wire \Tile_X5Y8_S4BEG[3] ;
 wire \Tile_X5Y8_S4BEG[4] ;
 wire \Tile_X5Y8_S4BEG[5] ;
 wire \Tile_X5Y8_S4BEG[6] ;
 wire \Tile_X5Y8_S4BEG[7] ;
 wire \Tile_X5Y8_S4BEG[8] ;
 wire \Tile_X5Y8_S4BEG[9] ;
 wire Tile_X5Y8_UserCLKo;
 wire \Tile_X5Y8_W1BEG[0] ;
 wire \Tile_X5Y8_W1BEG[1] ;
 wire \Tile_X5Y8_W1BEG[2] ;
 wire \Tile_X5Y8_W1BEG[3] ;
 wire \Tile_X5Y8_W2BEG[0] ;
 wire \Tile_X5Y8_W2BEG[1] ;
 wire \Tile_X5Y8_W2BEG[2] ;
 wire \Tile_X5Y8_W2BEG[3] ;
 wire \Tile_X5Y8_W2BEG[4] ;
 wire \Tile_X5Y8_W2BEG[5] ;
 wire \Tile_X5Y8_W2BEG[6] ;
 wire \Tile_X5Y8_W2BEG[7] ;
 wire \Tile_X5Y8_W2BEGb[0] ;
 wire \Tile_X5Y8_W2BEGb[1] ;
 wire \Tile_X5Y8_W2BEGb[2] ;
 wire \Tile_X5Y8_W2BEGb[3] ;
 wire \Tile_X5Y8_W2BEGb[4] ;
 wire \Tile_X5Y8_W2BEGb[5] ;
 wire \Tile_X5Y8_W2BEGb[6] ;
 wire \Tile_X5Y8_W2BEGb[7] ;
 wire \Tile_X5Y8_W6BEG[0] ;
 wire \Tile_X5Y8_W6BEG[10] ;
 wire \Tile_X5Y8_W6BEG[11] ;
 wire \Tile_X5Y8_W6BEG[1] ;
 wire \Tile_X5Y8_W6BEG[2] ;
 wire \Tile_X5Y8_W6BEG[3] ;
 wire \Tile_X5Y8_W6BEG[4] ;
 wire \Tile_X5Y8_W6BEG[5] ;
 wire \Tile_X5Y8_W6BEG[6] ;
 wire \Tile_X5Y8_W6BEG[7] ;
 wire \Tile_X5Y8_W6BEG[8] ;
 wire \Tile_X5Y8_W6BEG[9] ;
 wire \Tile_X5Y8_WW4BEG[0] ;
 wire \Tile_X5Y8_WW4BEG[10] ;
 wire \Tile_X5Y8_WW4BEG[11] ;
 wire \Tile_X5Y8_WW4BEG[12] ;
 wire \Tile_X5Y8_WW4BEG[13] ;
 wire \Tile_X5Y8_WW4BEG[14] ;
 wire \Tile_X5Y8_WW4BEG[15] ;
 wire \Tile_X5Y8_WW4BEG[1] ;
 wire \Tile_X5Y8_WW4BEG[2] ;
 wire \Tile_X5Y8_WW4BEG[3] ;
 wire \Tile_X5Y8_WW4BEG[4] ;
 wire \Tile_X5Y8_WW4BEG[5] ;
 wire \Tile_X5Y8_WW4BEG[6] ;
 wire \Tile_X5Y8_WW4BEG[7] ;
 wire \Tile_X5Y8_WW4BEG[8] ;
 wire \Tile_X5Y8_WW4BEG[9] ;
 wire \Tile_X5Y9_FrameData_O[0] ;
 wire \Tile_X5Y9_FrameData_O[10] ;
 wire \Tile_X5Y9_FrameData_O[11] ;
 wire \Tile_X5Y9_FrameData_O[12] ;
 wire \Tile_X5Y9_FrameData_O[13] ;
 wire \Tile_X5Y9_FrameData_O[14] ;
 wire \Tile_X5Y9_FrameData_O[15] ;
 wire \Tile_X5Y9_FrameData_O[16] ;
 wire \Tile_X5Y9_FrameData_O[17] ;
 wire \Tile_X5Y9_FrameData_O[18] ;
 wire \Tile_X5Y9_FrameData_O[19] ;
 wire \Tile_X5Y9_FrameData_O[1] ;
 wire \Tile_X5Y9_FrameData_O[20] ;
 wire \Tile_X5Y9_FrameData_O[21] ;
 wire \Tile_X5Y9_FrameData_O[22] ;
 wire \Tile_X5Y9_FrameData_O[23] ;
 wire \Tile_X5Y9_FrameData_O[24] ;
 wire \Tile_X5Y9_FrameData_O[25] ;
 wire \Tile_X5Y9_FrameData_O[26] ;
 wire \Tile_X5Y9_FrameData_O[27] ;
 wire \Tile_X5Y9_FrameData_O[28] ;
 wire \Tile_X5Y9_FrameData_O[29] ;
 wire \Tile_X5Y9_FrameData_O[2] ;
 wire \Tile_X5Y9_FrameData_O[30] ;
 wire \Tile_X5Y9_FrameData_O[31] ;
 wire \Tile_X5Y9_FrameData_O[3] ;
 wire \Tile_X5Y9_FrameData_O[4] ;
 wire \Tile_X5Y9_FrameData_O[5] ;
 wire \Tile_X5Y9_FrameData_O[6] ;
 wire \Tile_X5Y9_FrameData_O[7] ;
 wire \Tile_X5Y9_FrameData_O[8] ;
 wire \Tile_X5Y9_FrameData_O[9] ;
 wire \Tile_X5Y9_FrameStrobe_O[0] ;
 wire \Tile_X5Y9_FrameStrobe_O[10] ;
 wire \Tile_X5Y9_FrameStrobe_O[11] ;
 wire \Tile_X5Y9_FrameStrobe_O[12] ;
 wire \Tile_X5Y9_FrameStrobe_O[13] ;
 wire \Tile_X5Y9_FrameStrobe_O[14] ;
 wire \Tile_X5Y9_FrameStrobe_O[15] ;
 wire \Tile_X5Y9_FrameStrobe_O[16] ;
 wire \Tile_X5Y9_FrameStrobe_O[17] ;
 wire \Tile_X5Y9_FrameStrobe_O[18] ;
 wire \Tile_X5Y9_FrameStrobe_O[19] ;
 wire \Tile_X5Y9_FrameStrobe_O[1] ;
 wire \Tile_X5Y9_FrameStrobe_O[2] ;
 wire \Tile_X5Y9_FrameStrobe_O[3] ;
 wire \Tile_X5Y9_FrameStrobe_O[4] ;
 wire \Tile_X5Y9_FrameStrobe_O[5] ;
 wire \Tile_X5Y9_FrameStrobe_O[6] ;
 wire \Tile_X5Y9_FrameStrobe_O[7] ;
 wire \Tile_X5Y9_FrameStrobe_O[8] ;
 wire \Tile_X5Y9_FrameStrobe_O[9] ;
 wire \Tile_X5Y9_N1BEG[0] ;
 wire \Tile_X5Y9_N1BEG[1] ;
 wire \Tile_X5Y9_N1BEG[2] ;
 wire \Tile_X5Y9_N1BEG[3] ;
 wire \Tile_X5Y9_N2BEG[0] ;
 wire \Tile_X5Y9_N2BEG[1] ;
 wire \Tile_X5Y9_N2BEG[2] ;
 wire \Tile_X5Y9_N2BEG[3] ;
 wire \Tile_X5Y9_N2BEG[4] ;
 wire \Tile_X5Y9_N2BEG[5] ;
 wire \Tile_X5Y9_N2BEG[6] ;
 wire \Tile_X5Y9_N2BEG[7] ;
 wire \Tile_X5Y9_N2BEGb[0] ;
 wire \Tile_X5Y9_N2BEGb[1] ;
 wire \Tile_X5Y9_N2BEGb[2] ;
 wire \Tile_X5Y9_N2BEGb[3] ;
 wire \Tile_X5Y9_N2BEGb[4] ;
 wire \Tile_X5Y9_N2BEGb[5] ;
 wire \Tile_X5Y9_N2BEGb[6] ;
 wire \Tile_X5Y9_N2BEGb[7] ;
 wire \Tile_X5Y9_N4BEG[0] ;
 wire \Tile_X5Y9_N4BEG[10] ;
 wire \Tile_X5Y9_N4BEG[11] ;
 wire \Tile_X5Y9_N4BEG[12] ;
 wire \Tile_X5Y9_N4BEG[13] ;
 wire \Tile_X5Y9_N4BEG[14] ;
 wire \Tile_X5Y9_N4BEG[15] ;
 wire \Tile_X5Y9_N4BEG[1] ;
 wire \Tile_X5Y9_N4BEG[2] ;
 wire \Tile_X5Y9_N4BEG[3] ;
 wire \Tile_X5Y9_N4BEG[4] ;
 wire \Tile_X5Y9_N4BEG[5] ;
 wire \Tile_X5Y9_N4BEG[6] ;
 wire \Tile_X5Y9_N4BEG[7] ;
 wire \Tile_X5Y9_N4BEG[8] ;
 wire \Tile_X5Y9_N4BEG[9] ;
 wire Tile_X5Y9_UserCLKo;

 NW_term Tile_X0Y0_NW_term (.UserCLK(Tile_X0Y1_UserCLKo),
    .UserCLKo(Tile_X0Y0_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .FrameData({FrameData[31],
    FrameData[30],
    FrameData[29],
    FrameData[28],
    FrameData[27],
    FrameData[26],
    FrameData[25],
    FrameData[24],
    FrameData[23],
    FrameData[22],
    FrameData[21],
    FrameData[20],
    FrameData[19],
    FrameData[18],
    FrameData[17],
    FrameData[16],
    FrameData[15],
    FrameData[14],
    FrameData[13],
    FrameData[12],
    FrameData[11],
    FrameData[10],
    FrameData[9],
    FrameData[8],
    FrameData[7],
    FrameData[6],
    FrameData[5],
    FrameData[4],
    FrameData[3],
    FrameData[2],
    FrameData[1],
    FrameData[0]}),
    .FrameData_O({\Tile_X0Y0_FrameData_O[31] ,
    \Tile_X0Y0_FrameData_O[30] ,
    \Tile_X0Y0_FrameData_O[29] ,
    \Tile_X0Y0_FrameData_O[28] ,
    \Tile_X0Y0_FrameData_O[27] ,
    \Tile_X0Y0_FrameData_O[26] ,
    \Tile_X0Y0_FrameData_O[25] ,
    \Tile_X0Y0_FrameData_O[24] ,
    \Tile_X0Y0_FrameData_O[23] ,
    \Tile_X0Y0_FrameData_O[22] ,
    \Tile_X0Y0_FrameData_O[21] ,
    \Tile_X0Y0_FrameData_O[20] ,
    \Tile_X0Y0_FrameData_O[19] ,
    \Tile_X0Y0_FrameData_O[18] ,
    \Tile_X0Y0_FrameData_O[17] ,
    \Tile_X0Y0_FrameData_O[16] ,
    \Tile_X0Y0_FrameData_O[15] ,
    \Tile_X0Y0_FrameData_O[14] ,
    \Tile_X0Y0_FrameData_O[13] ,
    \Tile_X0Y0_FrameData_O[12] ,
    \Tile_X0Y0_FrameData_O[11] ,
    \Tile_X0Y0_FrameData_O[10] ,
    \Tile_X0Y0_FrameData_O[9] ,
    \Tile_X0Y0_FrameData_O[8] ,
    \Tile_X0Y0_FrameData_O[7] ,
    \Tile_X0Y0_FrameData_O[6] ,
    \Tile_X0Y0_FrameData_O[5] ,
    \Tile_X0Y0_FrameData_O[4] ,
    \Tile_X0Y0_FrameData_O[3] ,
    \Tile_X0Y0_FrameData_O[2] ,
    \Tile_X0Y0_FrameData_O[1] ,
    \Tile_X0Y0_FrameData_O[0] }),
    .FrameStrobe({\Tile_X0Y1_FrameStrobe_O[19] ,
    \Tile_X0Y1_FrameStrobe_O[18] ,
    \Tile_X0Y1_FrameStrobe_O[17] ,
    \Tile_X0Y1_FrameStrobe_O[16] ,
    \Tile_X0Y1_FrameStrobe_O[15] ,
    \Tile_X0Y1_FrameStrobe_O[14] ,
    \Tile_X0Y1_FrameStrobe_O[13] ,
    \Tile_X0Y1_FrameStrobe_O[12] ,
    \Tile_X0Y1_FrameStrobe_O[11] ,
    \Tile_X0Y1_FrameStrobe_O[10] ,
    \Tile_X0Y1_FrameStrobe_O[9] ,
    \Tile_X0Y1_FrameStrobe_O[8] ,
    \Tile_X0Y1_FrameStrobe_O[7] ,
    \Tile_X0Y1_FrameStrobe_O[6] ,
    \Tile_X0Y1_FrameStrobe_O[5] ,
    \Tile_X0Y1_FrameStrobe_O[4] ,
    \Tile_X0Y1_FrameStrobe_O[3] ,
    \Tile_X0Y1_FrameStrobe_O[2] ,
    \Tile_X0Y1_FrameStrobe_O[1] ,
    \Tile_X0Y1_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X0Y0_FrameStrobe_O[19] ,
    \Tile_X0Y0_FrameStrobe_O[18] ,
    \Tile_X0Y0_FrameStrobe_O[17] ,
    \Tile_X0Y0_FrameStrobe_O[16] ,
    \Tile_X0Y0_FrameStrobe_O[15] ,
    \Tile_X0Y0_FrameStrobe_O[14] ,
    \Tile_X0Y0_FrameStrobe_O[13] ,
    \Tile_X0Y0_FrameStrobe_O[12] ,
    \Tile_X0Y0_FrameStrobe_O[11] ,
    \Tile_X0Y0_FrameStrobe_O[10] ,
    \Tile_X0Y0_FrameStrobe_O[9] ,
    \Tile_X0Y0_FrameStrobe_O[8] ,
    \Tile_X0Y0_FrameStrobe_O[7] ,
    \Tile_X0Y0_FrameStrobe_O[6] ,
    \Tile_X0Y0_FrameStrobe_O[5] ,
    \Tile_X0Y0_FrameStrobe_O[4] ,
    \Tile_X0Y0_FrameStrobe_O[3] ,
    \Tile_X0Y0_FrameStrobe_O[2] ,
    \Tile_X0Y0_FrameStrobe_O[1] ,
    \Tile_X0Y0_FrameStrobe_O[0] }),
    .N1END({\Tile_X0Y1_N1BEG[3] ,
    \Tile_X0Y1_N1BEG[2] ,
    \Tile_X0Y1_N1BEG[1] ,
    \Tile_X0Y1_N1BEG[0] }),
    .N2END({\Tile_X0Y1_N2BEGb[7] ,
    \Tile_X0Y1_N2BEGb[6] ,
    \Tile_X0Y1_N2BEGb[5] ,
    \Tile_X0Y1_N2BEGb[4] ,
    \Tile_X0Y1_N2BEGb[3] ,
    \Tile_X0Y1_N2BEGb[2] ,
    \Tile_X0Y1_N2BEGb[1] ,
    \Tile_X0Y1_N2BEGb[0] }),
    .N2MID({\Tile_X0Y1_N2BEG[7] ,
    \Tile_X0Y1_N2BEG[6] ,
    \Tile_X0Y1_N2BEG[5] ,
    \Tile_X0Y1_N2BEG[4] ,
    \Tile_X0Y1_N2BEG[3] ,
    \Tile_X0Y1_N2BEG[2] ,
    \Tile_X0Y1_N2BEG[1] ,
    \Tile_X0Y1_N2BEG[0] }),
    .N4END({\Tile_X0Y1_N4BEG[15] ,
    \Tile_X0Y1_N4BEG[14] ,
    \Tile_X0Y1_N4BEG[13] ,
    \Tile_X0Y1_N4BEG[12] ,
    \Tile_X0Y1_N4BEG[11] ,
    \Tile_X0Y1_N4BEG[10] ,
    \Tile_X0Y1_N4BEG[9] ,
    \Tile_X0Y1_N4BEG[8] ,
    \Tile_X0Y1_N4BEG[7] ,
    \Tile_X0Y1_N4BEG[6] ,
    \Tile_X0Y1_N4BEG[5] ,
    \Tile_X0Y1_N4BEG[4] ,
    \Tile_X0Y1_N4BEG[3] ,
    \Tile_X0Y1_N4BEG[2] ,
    \Tile_X0Y1_N4BEG[1] ,
    \Tile_X0Y1_N4BEG[0] }),
    .S1BEG({\Tile_X0Y0_S1BEG[3] ,
    \Tile_X0Y0_S1BEG[2] ,
    \Tile_X0Y0_S1BEG[1] ,
    \Tile_X0Y0_S1BEG[0] }),
    .S2BEG({\Tile_X0Y0_S2BEG[7] ,
    \Tile_X0Y0_S2BEG[6] ,
    \Tile_X0Y0_S2BEG[5] ,
    \Tile_X0Y0_S2BEG[4] ,
    \Tile_X0Y0_S2BEG[3] ,
    \Tile_X0Y0_S2BEG[2] ,
    \Tile_X0Y0_S2BEG[1] ,
    \Tile_X0Y0_S2BEG[0] }),
    .S2BEGb({\Tile_X0Y0_S2BEGb[7] ,
    \Tile_X0Y0_S2BEGb[6] ,
    \Tile_X0Y0_S2BEGb[5] ,
    \Tile_X0Y0_S2BEGb[4] ,
    \Tile_X0Y0_S2BEGb[3] ,
    \Tile_X0Y0_S2BEGb[2] ,
    \Tile_X0Y0_S2BEGb[1] ,
    \Tile_X0Y0_S2BEGb[0] }),
    .S4BEG({\Tile_X0Y0_S4BEG[15] ,
    \Tile_X0Y0_S4BEG[14] ,
    \Tile_X0Y0_S4BEG[13] ,
    \Tile_X0Y0_S4BEG[12] ,
    \Tile_X0Y0_S4BEG[11] ,
    \Tile_X0Y0_S4BEG[10] ,
    \Tile_X0Y0_S4BEG[9] ,
    \Tile_X0Y0_S4BEG[8] ,
    \Tile_X0Y0_S4BEG[7] ,
    \Tile_X0Y0_S4BEG[6] ,
    \Tile_X0Y0_S4BEG[5] ,
    \Tile_X0Y0_S4BEG[4] ,
    \Tile_X0Y0_S4BEG[3] ,
    \Tile_X0Y0_S4BEG[2] ,
    \Tile_X0Y0_S4BEG[1] ,
    \Tile_X0Y0_S4BEG[0] }));
 W_TT_IF2 Tile_X0Y1_W_TT_IF2 (.CLK_TT_PROJECT(Tile_X0Y2_CLK_TT_PROJECT),
    .ENA_TT_PROJECT(Tile_X0Y2_ENA_TT_PROJECT),
    .RST_N_TT_PROJECT(Tile_X0Y2_RST_N_TT_PROJECT),
    .Tile_X0Y0_UserCLKo(Tile_X0Y1_UserCLKo),
    .Tile_X0Y1_UserCLK(Tile_X0Y3_UserCLKo),
    .UIO_IN_TT_PROJECT0(Tile_X0Y2_UIO_IN_TT_PROJECT0),
    .UIO_IN_TT_PROJECT1(Tile_X0Y2_UIO_IN_TT_PROJECT1),
    .UIO_IN_TT_PROJECT2(Tile_X0Y2_UIO_IN_TT_PROJECT2),
    .UIO_IN_TT_PROJECT3(Tile_X0Y2_UIO_IN_TT_PROJECT3),
    .UIO_IN_TT_PROJECT4(Tile_X0Y2_UIO_IN_TT_PROJECT4),
    .UIO_IN_TT_PROJECT5(Tile_X0Y2_UIO_IN_TT_PROJECT5),
    .UIO_IN_TT_PROJECT6(Tile_X0Y2_UIO_IN_TT_PROJECT6),
    .UIO_IN_TT_PROJECT7(Tile_X0Y2_UIO_IN_TT_PROJECT7),
    .UIO_OE_TT_PROJECT0(Tile_X0Y2_UIO_OE_TT_PROJECT0),
    .UIO_OE_TT_PROJECT1(Tile_X0Y2_UIO_OE_TT_PROJECT1),
    .UIO_OE_TT_PROJECT2(Tile_X0Y2_UIO_OE_TT_PROJECT2),
    .UIO_OE_TT_PROJECT3(Tile_X0Y2_UIO_OE_TT_PROJECT3),
    .UIO_OE_TT_PROJECT4(Tile_X0Y2_UIO_OE_TT_PROJECT4),
    .UIO_OE_TT_PROJECT5(Tile_X0Y2_UIO_OE_TT_PROJECT5),
    .UIO_OE_TT_PROJECT6(Tile_X0Y2_UIO_OE_TT_PROJECT6),
    .UIO_OE_TT_PROJECT7(Tile_X0Y2_UIO_OE_TT_PROJECT7),
    .UIO_OUT_TT_PROJECT0(Tile_X0Y2_UIO_OUT_TT_PROJECT0),
    .UIO_OUT_TT_PROJECT1(Tile_X0Y2_UIO_OUT_TT_PROJECT1),
    .UIO_OUT_TT_PROJECT2(Tile_X0Y2_UIO_OUT_TT_PROJECT2),
    .UIO_OUT_TT_PROJECT3(Tile_X0Y2_UIO_OUT_TT_PROJECT3),
    .UIO_OUT_TT_PROJECT4(Tile_X0Y2_UIO_OUT_TT_PROJECT4),
    .UIO_OUT_TT_PROJECT5(Tile_X0Y2_UIO_OUT_TT_PROJECT5),
    .UIO_OUT_TT_PROJECT6(Tile_X0Y2_UIO_OUT_TT_PROJECT6),
    .UIO_OUT_TT_PROJECT7(Tile_X0Y2_UIO_OUT_TT_PROJECT7),
    .UI_IN_TT_PROJECT0(Tile_X0Y2_UI_IN_TT_PROJECT0),
    .UI_IN_TT_PROJECT1(Tile_X0Y2_UI_IN_TT_PROJECT1),
    .UI_IN_TT_PROJECT2(Tile_X0Y2_UI_IN_TT_PROJECT2),
    .UI_IN_TT_PROJECT3(Tile_X0Y2_UI_IN_TT_PROJECT3),
    .UI_IN_TT_PROJECT4(Tile_X0Y2_UI_IN_TT_PROJECT4),
    .UI_IN_TT_PROJECT5(Tile_X0Y2_UI_IN_TT_PROJECT5),
    .UI_IN_TT_PROJECT6(Tile_X0Y2_UI_IN_TT_PROJECT6),
    .UI_IN_TT_PROJECT7(Tile_X0Y2_UI_IN_TT_PROJECT7),
    .UO_OUT_TT_PROJECT0(Tile_X0Y2_UO_OUT_TT_PROJECT0),
    .UO_OUT_TT_PROJECT1(Tile_X0Y2_UO_OUT_TT_PROJECT1),
    .UO_OUT_TT_PROJECT2(Tile_X0Y2_UO_OUT_TT_PROJECT2),
    .UO_OUT_TT_PROJECT3(Tile_X0Y2_UO_OUT_TT_PROJECT3),
    .UO_OUT_TT_PROJECT4(Tile_X0Y2_UO_OUT_TT_PROJECT4),
    .UO_OUT_TT_PROJECT5(Tile_X0Y2_UO_OUT_TT_PROJECT5),
    .UO_OUT_TT_PROJECT6(Tile_X0Y2_UO_OUT_TT_PROJECT6),
    .UO_OUT_TT_PROJECT7(Tile_X0Y2_UO_OUT_TT_PROJECT7),
    .VGND(VGND),
    .VPWR(VPWR),
    .Tile_X0Y0_E1BEG({\Tile_X0Y1_E1BEG[3] ,
    \Tile_X0Y1_E1BEG[2] ,
    \Tile_X0Y1_E1BEG[1] ,
    \Tile_X0Y1_E1BEG[0] }),
    .Tile_X0Y0_E2BEG({\Tile_X0Y1_E2BEG[7] ,
    \Tile_X0Y1_E2BEG[6] ,
    \Tile_X0Y1_E2BEG[5] ,
    \Tile_X0Y1_E2BEG[4] ,
    \Tile_X0Y1_E2BEG[3] ,
    \Tile_X0Y1_E2BEG[2] ,
    \Tile_X0Y1_E2BEG[1] ,
    \Tile_X0Y1_E2BEG[0] }),
    .Tile_X0Y0_E2BEGb({\Tile_X0Y1_E2BEGb[7] ,
    \Tile_X0Y1_E2BEGb[6] ,
    \Tile_X0Y1_E2BEGb[5] ,
    \Tile_X0Y1_E2BEGb[4] ,
    \Tile_X0Y1_E2BEGb[3] ,
    \Tile_X0Y1_E2BEGb[2] ,
    \Tile_X0Y1_E2BEGb[1] ,
    \Tile_X0Y1_E2BEGb[0] }),
    .Tile_X0Y0_E6BEG({\Tile_X0Y1_E6BEG[11] ,
    \Tile_X0Y1_E6BEG[10] ,
    \Tile_X0Y1_E6BEG[9] ,
    \Tile_X0Y1_E6BEG[8] ,
    \Tile_X0Y1_E6BEG[7] ,
    \Tile_X0Y1_E6BEG[6] ,
    \Tile_X0Y1_E6BEG[5] ,
    \Tile_X0Y1_E6BEG[4] ,
    \Tile_X0Y1_E6BEG[3] ,
    \Tile_X0Y1_E6BEG[2] ,
    \Tile_X0Y1_E6BEG[1] ,
    \Tile_X0Y1_E6BEG[0] }),
    .Tile_X0Y0_EE4BEG({\Tile_X0Y1_EE4BEG[15] ,
    \Tile_X0Y1_EE4BEG[14] ,
    \Tile_X0Y1_EE4BEG[13] ,
    \Tile_X0Y1_EE4BEG[12] ,
    \Tile_X0Y1_EE4BEG[11] ,
    \Tile_X0Y1_EE4BEG[10] ,
    \Tile_X0Y1_EE4BEG[9] ,
    \Tile_X0Y1_EE4BEG[8] ,
    \Tile_X0Y1_EE4BEG[7] ,
    \Tile_X0Y1_EE4BEG[6] ,
    \Tile_X0Y1_EE4BEG[5] ,
    \Tile_X0Y1_EE4BEG[4] ,
    \Tile_X0Y1_EE4BEG[3] ,
    \Tile_X0Y1_EE4BEG[2] ,
    \Tile_X0Y1_EE4BEG[1] ,
    \Tile_X0Y1_EE4BEG[0] }),
    .Tile_X0Y0_FrameData({FrameData[63],
    FrameData[62],
    FrameData[61],
    FrameData[60],
    FrameData[59],
    FrameData[58],
    FrameData[57],
    FrameData[56],
    FrameData[55],
    FrameData[54],
    FrameData[53],
    FrameData[52],
    FrameData[51],
    FrameData[50],
    FrameData[49],
    FrameData[48],
    FrameData[47],
    FrameData[46],
    FrameData[45],
    FrameData[44],
    FrameData[43],
    FrameData[42],
    FrameData[41],
    FrameData[40],
    FrameData[39],
    FrameData[38],
    FrameData[37],
    FrameData[36],
    FrameData[35],
    FrameData[34],
    FrameData[33],
    FrameData[32]}),
    .Tile_X0Y0_FrameData_O({\Tile_X0Y1_FrameData_O[31] ,
    \Tile_X0Y1_FrameData_O[30] ,
    \Tile_X0Y1_FrameData_O[29] ,
    \Tile_X0Y1_FrameData_O[28] ,
    \Tile_X0Y1_FrameData_O[27] ,
    \Tile_X0Y1_FrameData_O[26] ,
    \Tile_X0Y1_FrameData_O[25] ,
    \Tile_X0Y1_FrameData_O[24] ,
    \Tile_X0Y1_FrameData_O[23] ,
    \Tile_X0Y1_FrameData_O[22] ,
    \Tile_X0Y1_FrameData_O[21] ,
    \Tile_X0Y1_FrameData_O[20] ,
    \Tile_X0Y1_FrameData_O[19] ,
    \Tile_X0Y1_FrameData_O[18] ,
    \Tile_X0Y1_FrameData_O[17] ,
    \Tile_X0Y1_FrameData_O[16] ,
    \Tile_X0Y1_FrameData_O[15] ,
    \Tile_X0Y1_FrameData_O[14] ,
    \Tile_X0Y1_FrameData_O[13] ,
    \Tile_X0Y1_FrameData_O[12] ,
    \Tile_X0Y1_FrameData_O[11] ,
    \Tile_X0Y1_FrameData_O[10] ,
    \Tile_X0Y1_FrameData_O[9] ,
    \Tile_X0Y1_FrameData_O[8] ,
    \Tile_X0Y1_FrameData_O[7] ,
    \Tile_X0Y1_FrameData_O[6] ,
    \Tile_X0Y1_FrameData_O[5] ,
    \Tile_X0Y1_FrameData_O[4] ,
    \Tile_X0Y1_FrameData_O[3] ,
    \Tile_X0Y1_FrameData_O[2] ,
    \Tile_X0Y1_FrameData_O[1] ,
    \Tile_X0Y1_FrameData_O[0] }),
    .Tile_X0Y0_FrameStrobe_O({\Tile_X0Y1_FrameStrobe_O[19] ,
    \Tile_X0Y1_FrameStrobe_O[18] ,
    \Tile_X0Y1_FrameStrobe_O[17] ,
    \Tile_X0Y1_FrameStrobe_O[16] ,
    \Tile_X0Y1_FrameStrobe_O[15] ,
    \Tile_X0Y1_FrameStrobe_O[14] ,
    \Tile_X0Y1_FrameStrobe_O[13] ,
    \Tile_X0Y1_FrameStrobe_O[12] ,
    \Tile_X0Y1_FrameStrobe_O[11] ,
    \Tile_X0Y1_FrameStrobe_O[10] ,
    \Tile_X0Y1_FrameStrobe_O[9] ,
    \Tile_X0Y1_FrameStrobe_O[8] ,
    \Tile_X0Y1_FrameStrobe_O[7] ,
    \Tile_X0Y1_FrameStrobe_O[6] ,
    \Tile_X0Y1_FrameStrobe_O[5] ,
    \Tile_X0Y1_FrameStrobe_O[4] ,
    \Tile_X0Y1_FrameStrobe_O[3] ,
    \Tile_X0Y1_FrameStrobe_O[2] ,
    \Tile_X0Y1_FrameStrobe_O[1] ,
    \Tile_X0Y1_FrameStrobe_O[0] }),
    .Tile_X0Y0_N1BEG({\Tile_X0Y1_N1BEG[3] ,
    \Tile_X0Y1_N1BEG[2] ,
    \Tile_X0Y1_N1BEG[1] ,
    \Tile_X0Y1_N1BEG[0] }),
    .Tile_X0Y0_N2BEG({\Tile_X0Y1_N2BEG[7] ,
    \Tile_X0Y1_N2BEG[6] ,
    \Tile_X0Y1_N2BEG[5] ,
    \Tile_X0Y1_N2BEG[4] ,
    \Tile_X0Y1_N2BEG[3] ,
    \Tile_X0Y1_N2BEG[2] ,
    \Tile_X0Y1_N2BEG[1] ,
    \Tile_X0Y1_N2BEG[0] }),
    .Tile_X0Y0_N2BEGb({\Tile_X0Y1_N2BEGb[7] ,
    \Tile_X0Y1_N2BEGb[6] ,
    \Tile_X0Y1_N2BEGb[5] ,
    \Tile_X0Y1_N2BEGb[4] ,
    \Tile_X0Y1_N2BEGb[3] ,
    \Tile_X0Y1_N2BEGb[2] ,
    \Tile_X0Y1_N2BEGb[1] ,
    \Tile_X0Y1_N2BEGb[0] }),
    .Tile_X0Y0_N4BEG({\Tile_X0Y1_N4BEG[15] ,
    \Tile_X0Y1_N4BEG[14] ,
    \Tile_X0Y1_N4BEG[13] ,
    \Tile_X0Y1_N4BEG[12] ,
    \Tile_X0Y1_N4BEG[11] ,
    \Tile_X0Y1_N4BEG[10] ,
    \Tile_X0Y1_N4BEG[9] ,
    \Tile_X0Y1_N4BEG[8] ,
    \Tile_X0Y1_N4BEG[7] ,
    \Tile_X0Y1_N4BEG[6] ,
    \Tile_X0Y1_N4BEG[5] ,
    \Tile_X0Y1_N4BEG[4] ,
    \Tile_X0Y1_N4BEG[3] ,
    \Tile_X0Y1_N4BEG[2] ,
    \Tile_X0Y1_N4BEG[1] ,
    \Tile_X0Y1_N4BEG[0] }),
    .Tile_X0Y0_S1END({\Tile_X0Y0_S1BEG[3] ,
    \Tile_X0Y0_S1BEG[2] ,
    \Tile_X0Y0_S1BEG[1] ,
    \Tile_X0Y0_S1BEG[0] }),
    .Tile_X0Y0_S2END({\Tile_X0Y0_S2BEGb[7] ,
    \Tile_X0Y0_S2BEGb[6] ,
    \Tile_X0Y0_S2BEGb[5] ,
    \Tile_X0Y0_S2BEGb[4] ,
    \Tile_X0Y0_S2BEGb[3] ,
    \Tile_X0Y0_S2BEGb[2] ,
    \Tile_X0Y0_S2BEGb[1] ,
    \Tile_X0Y0_S2BEGb[0] }),
    .Tile_X0Y0_S2MID({\Tile_X0Y0_S2BEG[7] ,
    \Tile_X0Y0_S2BEG[6] ,
    \Tile_X0Y0_S2BEG[5] ,
    \Tile_X0Y0_S2BEG[4] ,
    \Tile_X0Y0_S2BEG[3] ,
    \Tile_X0Y0_S2BEG[2] ,
    \Tile_X0Y0_S2BEG[1] ,
    \Tile_X0Y0_S2BEG[0] }),
    .Tile_X0Y0_S4END({\Tile_X0Y0_S4BEG[15] ,
    \Tile_X0Y0_S4BEG[14] ,
    \Tile_X0Y0_S4BEG[13] ,
    \Tile_X0Y0_S4BEG[12] ,
    \Tile_X0Y0_S4BEG[11] ,
    \Tile_X0Y0_S4BEG[10] ,
    \Tile_X0Y0_S4BEG[9] ,
    \Tile_X0Y0_S4BEG[8] ,
    \Tile_X0Y0_S4BEG[7] ,
    \Tile_X0Y0_S4BEG[6] ,
    \Tile_X0Y0_S4BEG[5] ,
    \Tile_X0Y0_S4BEG[4] ,
    \Tile_X0Y0_S4BEG[3] ,
    \Tile_X0Y0_S4BEG[2] ,
    \Tile_X0Y0_S4BEG[1] ,
    \Tile_X0Y0_S4BEG[0] }),
    .Tile_X0Y0_W1END({\Tile_X1Y1_W1BEG[3] ,
    \Tile_X1Y1_W1BEG[2] ,
    \Tile_X1Y1_W1BEG[1] ,
    \Tile_X1Y1_W1BEG[0] }),
    .Tile_X0Y0_W2END({\Tile_X1Y1_W2BEGb[7] ,
    \Tile_X1Y1_W2BEGb[6] ,
    \Tile_X1Y1_W2BEGb[5] ,
    \Tile_X1Y1_W2BEGb[4] ,
    \Tile_X1Y1_W2BEGb[3] ,
    \Tile_X1Y1_W2BEGb[2] ,
    \Tile_X1Y1_W2BEGb[1] ,
    \Tile_X1Y1_W2BEGb[0] }),
    .Tile_X0Y0_W2MID({\Tile_X1Y1_W2BEG[7] ,
    \Tile_X1Y1_W2BEG[6] ,
    \Tile_X1Y1_W2BEG[5] ,
    \Tile_X1Y1_W2BEG[4] ,
    \Tile_X1Y1_W2BEG[3] ,
    \Tile_X1Y1_W2BEG[2] ,
    \Tile_X1Y1_W2BEG[1] ,
    \Tile_X1Y1_W2BEG[0] }),
    .Tile_X0Y0_W6END({\Tile_X1Y1_W6BEG[11] ,
    \Tile_X1Y1_W6BEG[10] ,
    \Tile_X1Y1_W6BEG[9] ,
    \Tile_X1Y1_W6BEG[8] ,
    \Tile_X1Y1_W6BEG[7] ,
    \Tile_X1Y1_W6BEG[6] ,
    \Tile_X1Y1_W6BEG[5] ,
    \Tile_X1Y1_W6BEG[4] ,
    \Tile_X1Y1_W6BEG[3] ,
    \Tile_X1Y1_W6BEG[2] ,
    \Tile_X1Y1_W6BEG[1] ,
    \Tile_X1Y1_W6BEG[0] }),
    .Tile_X0Y0_WW4END({\Tile_X1Y1_WW4BEG[15] ,
    \Tile_X1Y1_WW4BEG[14] ,
    \Tile_X1Y1_WW4BEG[13] ,
    \Tile_X1Y1_WW4BEG[12] ,
    \Tile_X1Y1_WW4BEG[11] ,
    \Tile_X1Y1_WW4BEG[10] ,
    \Tile_X1Y1_WW4BEG[9] ,
    \Tile_X1Y1_WW4BEG[8] ,
    \Tile_X1Y1_WW4BEG[7] ,
    \Tile_X1Y1_WW4BEG[6] ,
    \Tile_X1Y1_WW4BEG[5] ,
    \Tile_X1Y1_WW4BEG[4] ,
    \Tile_X1Y1_WW4BEG[3] ,
    \Tile_X1Y1_WW4BEG[2] ,
    \Tile_X1Y1_WW4BEG[1] ,
    \Tile_X1Y1_WW4BEG[0] }),
    .Tile_X0Y1_E1BEG({\Tile_X0Y2_E1BEG[3] ,
    \Tile_X0Y2_E1BEG[2] ,
    \Tile_X0Y2_E1BEG[1] ,
    \Tile_X0Y2_E1BEG[0] }),
    .Tile_X0Y1_E2BEG({\Tile_X0Y2_E2BEG[7] ,
    \Tile_X0Y2_E2BEG[6] ,
    \Tile_X0Y2_E2BEG[5] ,
    \Tile_X0Y2_E2BEG[4] ,
    \Tile_X0Y2_E2BEG[3] ,
    \Tile_X0Y2_E2BEG[2] ,
    \Tile_X0Y2_E2BEG[1] ,
    \Tile_X0Y2_E2BEG[0] }),
    .Tile_X0Y1_E2BEGb({\Tile_X0Y2_E2BEGb[7] ,
    \Tile_X0Y2_E2BEGb[6] ,
    \Tile_X0Y2_E2BEGb[5] ,
    \Tile_X0Y2_E2BEGb[4] ,
    \Tile_X0Y2_E2BEGb[3] ,
    \Tile_X0Y2_E2BEGb[2] ,
    \Tile_X0Y2_E2BEGb[1] ,
    \Tile_X0Y2_E2BEGb[0] }),
    .Tile_X0Y1_E6BEG({\Tile_X0Y2_E6BEG[11] ,
    \Tile_X0Y2_E6BEG[10] ,
    \Tile_X0Y2_E6BEG[9] ,
    \Tile_X0Y2_E6BEG[8] ,
    \Tile_X0Y2_E6BEG[7] ,
    \Tile_X0Y2_E6BEG[6] ,
    \Tile_X0Y2_E6BEG[5] ,
    \Tile_X0Y2_E6BEG[4] ,
    \Tile_X0Y2_E6BEG[3] ,
    \Tile_X0Y2_E6BEG[2] ,
    \Tile_X0Y2_E6BEG[1] ,
    \Tile_X0Y2_E6BEG[0] }),
    .Tile_X0Y1_EE4BEG({\Tile_X0Y2_EE4BEG[15] ,
    \Tile_X0Y2_EE4BEG[14] ,
    \Tile_X0Y2_EE4BEG[13] ,
    \Tile_X0Y2_EE4BEG[12] ,
    \Tile_X0Y2_EE4BEG[11] ,
    \Tile_X0Y2_EE4BEG[10] ,
    \Tile_X0Y2_EE4BEG[9] ,
    \Tile_X0Y2_EE4BEG[8] ,
    \Tile_X0Y2_EE4BEG[7] ,
    \Tile_X0Y2_EE4BEG[6] ,
    \Tile_X0Y2_EE4BEG[5] ,
    \Tile_X0Y2_EE4BEG[4] ,
    \Tile_X0Y2_EE4BEG[3] ,
    \Tile_X0Y2_EE4BEG[2] ,
    \Tile_X0Y2_EE4BEG[1] ,
    \Tile_X0Y2_EE4BEG[0] }),
    .Tile_X0Y1_FrameData({FrameData[95],
    FrameData[94],
    FrameData[93],
    FrameData[92],
    FrameData[91],
    FrameData[90],
    FrameData[89],
    FrameData[88],
    FrameData[87],
    FrameData[86],
    FrameData[85],
    FrameData[84],
    FrameData[83],
    FrameData[82],
    FrameData[81],
    FrameData[80],
    FrameData[79],
    FrameData[78],
    FrameData[77],
    FrameData[76],
    FrameData[75],
    FrameData[74],
    FrameData[73],
    FrameData[72],
    FrameData[71],
    FrameData[70],
    FrameData[69],
    FrameData[68],
    FrameData[67],
    FrameData[66],
    FrameData[65],
    FrameData[64]}),
    .Tile_X0Y1_FrameData_O({\Tile_X0Y2_FrameData_O[31] ,
    \Tile_X0Y2_FrameData_O[30] ,
    \Tile_X0Y2_FrameData_O[29] ,
    \Tile_X0Y2_FrameData_O[28] ,
    \Tile_X0Y2_FrameData_O[27] ,
    \Tile_X0Y2_FrameData_O[26] ,
    \Tile_X0Y2_FrameData_O[25] ,
    \Tile_X0Y2_FrameData_O[24] ,
    \Tile_X0Y2_FrameData_O[23] ,
    \Tile_X0Y2_FrameData_O[22] ,
    \Tile_X0Y2_FrameData_O[21] ,
    \Tile_X0Y2_FrameData_O[20] ,
    \Tile_X0Y2_FrameData_O[19] ,
    \Tile_X0Y2_FrameData_O[18] ,
    \Tile_X0Y2_FrameData_O[17] ,
    \Tile_X0Y2_FrameData_O[16] ,
    \Tile_X0Y2_FrameData_O[15] ,
    \Tile_X0Y2_FrameData_O[14] ,
    \Tile_X0Y2_FrameData_O[13] ,
    \Tile_X0Y2_FrameData_O[12] ,
    \Tile_X0Y2_FrameData_O[11] ,
    \Tile_X0Y2_FrameData_O[10] ,
    \Tile_X0Y2_FrameData_O[9] ,
    \Tile_X0Y2_FrameData_O[8] ,
    \Tile_X0Y2_FrameData_O[7] ,
    \Tile_X0Y2_FrameData_O[6] ,
    \Tile_X0Y2_FrameData_O[5] ,
    \Tile_X0Y2_FrameData_O[4] ,
    \Tile_X0Y2_FrameData_O[3] ,
    \Tile_X0Y2_FrameData_O[2] ,
    \Tile_X0Y2_FrameData_O[1] ,
    \Tile_X0Y2_FrameData_O[0] }),
    .Tile_X0Y1_FrameStrobe({\Tile_X0Y3_FrameStrobe_O[19] ,
    \Tile_X0Y3_FrameStrobe_O[18] ,
    \Tile_X0Y3_FrameStrobe_O[17] ,
    \Tile_X0Y3_FrameStrobe_O[16] ,
    \Tile_X0Y3_FrameStrobe_O[15] ,
    \Tile_X0Y3_FrameStrobe_O[14] ,
    \Tile_X0Y3_FrameStrobe_O[13] ,
    \Tile_X0Y3_FrameStrobe_O[12] ,
    \Tile_X0Y3_FrameStrobe_O[11] ,
    \Tile_X0Y3_FrameStrobe_O[10] ,
    \Tile_X0Y3_FrameStrobe_O[9] ,
    \Tile_X0Y3_FrameStrobe_O[8] ,
    \Tile_X0Y3_FrameStrobe_O[7] ,
    \Tile_X0Y3_FrameStrobe_O[6] ,
    \Tile_X0Y3_FrameStrobe_O[5] ,
    \Tile_X0Y3_FrameStrobe_O[4] ,
    \Tile_X0Y3_FrameStrobe_O[3] ,
    \Tile_X0Y3_FrameStrobe_O[2] ,
    \Tile_X0Y3_FrameStrobe_O[1] ,
    \Tile_X0Y3_FrameStrobe_O[0] }),
    .Tile_X0Y1_N1END({\Tile_X0Y3_N1BEG[3] ,
    \Tile_X0Y3_N1BEG[2] ,
    \Tile_X0Y3_N1BEG[1] ,
    \Tile_X0Y3_N1BEG[0] }),
    .Tile_X0Y1_N2END({\Tile_X0Y3_N2BEGb[7] ,
    \Tile_X0Y3_N2BEGb[6] ,
    \Tile_X0Y3_N2BEGb[5] ,
    \Tile_X0Y3_N2BEGb[4] ,
    \Tile_X0Y3_N2BEGb[3] ,
    \Tile_X0Y3_N2BEGb[2] ,
    \Tile_X0Y3_N2BEGb[1] ,
    \Tile_X0Y3_N2BEGb[0] }),
    .Tile_X0Y1_N2MID({\Tile_X0Y3_N2BEG[7] ,
    \Tile_X0Y3_N2BEG[6] ,
    \Tile_X0Y3_N2BEG[5] ,
    \Tile_X0Y3_N2BEG[4] ,
    \Tile_X0Y3_N2BEG[3] ,
    \Tile_X0Y3_N2BEG[2] ,
    \Tile_X0Y3_N2BEG[1] ,
    \Tile_X0Y3_N2BEG[0] }),
    .Tile_X0Y1_N4END({\Tile_X0Y3_N4BEG[15] ,
    \Tile_X0Y3_N4BEG[14] ,
    \Tile_X0Y3_N4BEG[13] ,
    \Tile_X0Y3_N4BEG[12] ,
    \Tile_X0Y3_N4BEG[11] ,
    \Tile_X0Y3_N4BEG[10] ,
    \Tile_X0Y3_N4BEG[9] ,
    \Tile_X0Y3_N4BEG[8] ,
    \Tile_X0Y3_N4BEG[7] ,
    \Tile_X0Y3_N4BEG[6] ,
    \Tile_X0Y3_N4BEG[5] ,
    \Tile_X0Y3_N4BEG[4] ,
    \Tile_X0Y3_N4BEG[3] ,
    \Tile_X0Y3_N4BEG[2] ,
    \Tile_X0Y3_N4BEG[1] ,
    \Tile_X0Y3_N4BEG[0] }),
    .Tile_X0Y1_S1BEG({\Tile_X0Y2_S1BEG[3] ,
    \Tile_X0Y2_S1BEG[2] ,
    \Tile_X0Y2_S1BEG[1] ,
    \Tile_X0Y2_S1BEG[0] }),
    .Tile_X0Y1_S2BEG({\Tile_X0Y2_S2BEG[7] ,
    \Tile_X0Y2_S2BEG[6] ,
    \Tile_X0Y2_S2BEG[5] ,
    \Tile_X0Y2_S2BEG[4] ,
    \Tile_X0Y2_S2BEG[3] ,
    \Tile_X0Y2_S2BEG[2] ,
    \Tile_X0Y2_S2BEG[1] ,
    \Tile_X0Y2_S2BEG[0] }),
    .Tile_X0Y1_S2BEGb({\Tile_X0Y2_S2BEGb[7] ,
    \Tile_X0Y2_S2BEGb[6] ,
    \Tile_X0Y2_S2BEGb[5] ,
    \Tile_X0Y2_S2BEGb[4] ,
    \Tile_X0Y2_S2BEGb[3] ,
    \Tile_X0Y2_S2BEGb[2] ,
    \Tile_X0Y2_S2BEGb[1] ,
    \Tile_X0Y2_S2BEGb[0] }),
    .Tile_X0Y1_S4BEG({\Tile_X0Y2_S4BEG[15] ,
    \Tile_X0Y2_S4BEG[14] ,
    \Tile_X0Y2_S4BEG[13] ,
    \Tile_X0Y2_S4BEG[12] ,
    \Tile_X0Y2_S4BEG[11] ,
    \Tile_X0Y2_S4BEG[10] ,
    \Tile_X0Y2_S4BEG[9] ,
    \Tile_X0Y2_S4BEG[8] ,
    \Tile_X0Y2_S4BEG[7] ,
    \Tile_X0Y2_S4BEG[6] ,
    \Tile_X0Y2_S4BEG[5] ,
    \Tile_X0Y2_S4BEG[4] ,
    \Tile_X0Y2_S4BEG[3] ,
    \Tile_X0Y2_S4BEG[2] ,
    \Tile_X0Y2_S4BEG[1] ,
    \Tile_X0Y2_S4BEG[0] }),
    .Tile_X0Y1_W1END({\Tile_X1Y2_W1BEG[3] ,
    \Tile_X1Y2_W1BEG[2] ,
    \Tile_X1Y2_W1BEG[1] ,
    \Tile_X1Y2_W1BEG[0] }),
    .Tile_X0Y1_W2END({\Tile_X1Y2_W2BEGb[7] ,
    \Tile_X1Y2_W2BEGb[6] ,
    \Tile_X1Y2_W2BEGb[5] ,
    \Tile_X1Y2_W2BEGb[4] ,
    \Tile_X1Y2_W2BEGb[3] ,
    \Tile_X1Y2_W2BEGb[2] ,
    \Tile_X1Y2_W2BEGb[1] ,
    \Tile_X1Y2_W2BEGb[0] }),
    .Tile_X0Y1_W2MID({\Tile_X1Y2_W2BEG[7] ,
    \Tile_X1Y2_W2BEG[6] ,
    \Tile_X1Y2_W2BEG[5] ,
    \Tile_X1Y2_W2BEG[4] ,
    \Tile_X1Y2_W2BEG[3] ,
    \Tile_X1Y2_W2BEG[2] ,
    \Tile_X1Y2_W2BEG[1] ,
    \Tile_X1Y2_W2BEG[0] }),
    .Tile_X0Y1_W6END({\Tile_X1Y2_W6BEG[11] ,
    \Tile_X1Y2_W6BEG[10] ,
    \Tile_X1Y2_W6BEG[9] ,
    \Tile_X1Y2_W6BEG[8] ,
    \Tile_X1Y2_W6BEG[7] ,
    \Tile_X1Y2_W6BEG[6] ,
    \Tile_X1Y2_W6BEG[5] ,
    \Tile_X1Y2_W6BEG[4] ,
    \Tile_X1Y2_W6BEG[3] ,
    \Tile_X1Y2_W6BEG[2] ,
    \Tile_X1Y2_W6BEG[1] ,
    \Tile_X1Y2_W6BEG[0] }),
    .Tile_X0Y1_WW4END({\Tile_X1Y2_WW4BEG[15] ,
    \Tile_X1Y2_WW4BEG[14] ,
    \Tile_X1Y2_WW4BEG[13] ,
    \Tile_X1Y2_WW4BEG[12] ,
    \Tile_X1Y2_WW4BEG[11] ,
    \Tile_X1Y2_WW4BEG[10] ,
    \Tile_X1Y2_WW4BEG[9] ,
    \Tile_X1Y2_WW4BEG[8] ,
    \Tile_X1Y2_WW4BEG[7] ,
    \Tile_X1Y2_WW4BEG[6] ,
    \Tile_X1Y2_WW4BEG[5] ,
    \Tile_X1Y2_WW4BEG[4] ,
    \Tile_X1Y2_WW4BEG[3] ,
    \Tile_X1Y2_WW4BEG[2] ,
    \Tile_X1Y2_WW4BEG[1] ,
    \Tile_X1Y2_WW4BEG[0] }));
 W_TT_IF Tile_X0Y3_W_TT_IF (.CLK_TT_PROJECT(Tile_X0Y3_CLK_TT_PROJECT),
    .ENA_TT_PROJECT(Tile_X0Y3_ENA_TT_PROJECT),
    .RST_N_TT_PROJECT(Tile_X0Y3_RST_N_TT_PROJECT),
    .UIO_IN_TT_PROJECT0(Tile_X0Y3_UIO_IN_TT_PROJECT0),
    .UIO_IN_TT_PROJECT1(Tile_X0Y3_UIO_IN_TT_PROJECT1),
    .UIO_IN_TT_PROJECT2(Tile_X0Y3_UIO_IN_TT_PROJECT2),
    .UIO_IN_TT_PROJECT3(Tile_X0Y3_UIO_IN_TT_PROJECT3),
    .UIO_IN_TT_PROJECT4(Tile_X0Y3_UIO_IN_TT_PROJECT4),
    .UIO_IN_TT_PROJECT5(Tile_X0Y3_UIO_IN_TT_PROJECT5),
    .UIO_IN_TT_PROJECT6(Tile_X0Y3_UIO_IN_TT_PROJECT6),
    .UIO_IN_TT_PROJECT7(Tile_X0Y3_UIO_IN_TT_PROJECT7),
    .UIO_OE_TT_PROJECT0(Tile_X0Y3_UIO_OE_TT_PROJECT0),
    .UIO_OE_TT_PROJECT1(Tile_X0Y3_UIO_OE_TT_PROJECT1),
    .UIO_OE_TT_PROJECT2(Tile_X0Y3_UIO_OE_TT_PROJECT2),
    .UIO_OE_TT_PROJECT3(Tile_X0Y3_UIO_OE_TT_PROJECT3),
    .UIO_OE_TT_PROJECT4(Tile_X0Y3_UIO_OE_TT_PROJECT4),
    .UIO_OE_TT_PROJECT5(Tile_X0Y3_UIO_OE_TT_PROJECT5),
    .UIO_OE_TT_PROJECT6(Tile_X0Y3_UIO_OE_TT_PROJECT6),
    .UIO_OE_TT_PROJECT7(Tile_X0Y3_UIO_OE_TT_PROJECT7),
    .UIO_OUT_TT_PROJECT0(Tile_X0Y3_UIO_OUT_TT_PROJECT0),
    .UIO_OUT_TT_PROJECT1(Tile_X0Y3_UIO_OUT_TT_PROJECT1),
    .UIO_OUT_TT_PROJECT2(Tile_X0Y3_UIO_OUT_TT_PROJECT2),
    .UIO_OUT_TT_PROJECT3(Tile_X0Y3_UIO_OUT_TT_PROJECT3),
    .UIO_OUT_TT_PROJECT4(Tile_X0Y3_UIO_OUT_TT_PROJECT4),
    .UIO_OUT_TT_PROJECT5(Tile_X0Y3_UIO_OUT_TT_PROJECT5),
    .UIO_OUT_TT_PROJECT6(Tile_X0Y3_UIO_OUT_TT_PROJECT6),
    .UIO_OUT_TT_PROJECT7(Tile_X0Y3_UIO_OUT_TT_PROJECT7),
    .UI_IN_TT_PROJECT0(Tile_X0Y3_UI_IN_TT_PROJECT0),
    .UI_IN_TT_PROJECT1(Tile_X0Y3_UI_IN_TT_PROJECT1),
    .UI_IN_TT_PROJECT2(Tile_X0Y3_UI_IN_TT_PROJECT2),
    .UI_IN_TT_PROJECT3(Tile_X0Y3_UI_IN_TT_PROJECT3),
    .UI_IN_TT_PROJECT4(Tile_X0Y3_UI_IN_TT_PROJECT4),
    .UI_IN_TT_PROJECT5(Tile_X0Y3_UI_IN_TT_PROJECT5),
    .UI_IN_TT_PROJECT6(Tile_X0Y3_UI_IN_TT_PROJECT6),
    .UI_IN_TT_PROJECT7(Tile_X0Y3_UI_IN_TT_PROJECT7),
    .UO_OUT_TT_PROJECT0(Tile_X0Y3_UO_OUT_TT_PROJECT0),
    .UO_OUT_TT_PROJECT1(Tile_X0Y3_UO_OUT_TT_PROJECT1),
    .UO_OUT_TT_PROJECT2(Tile_X0Y3_UO_OUT_TT_PROJECT2),
    .UO_OUT_TT_PROJECT3(Tile_X0Y3_UO_OUT_TT_PROJECT3),
    .UO_OUT_TT_PROJECT4(Tile_X0Y3_UO_OUT_TT_PROJECT4),
    .UO_OUT_TT_PROJECT5(Tile_X0Y3_UO_OUT_TT_PROJECT5),
    .UO_OUT_TT_PROJECT6(Tile_X0Y3_UO_OUT_TT_PROJECT6),
    .UO_OUT_TT_PROJECT7(Tile_X0Y3_UO_OUT_TT_PROJECT7),
    .UserCLK(Tile_X0Y4_UserCLKo),
    .UserCLKo(Tile_X0Y3_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X0Y3_E1BEG[3] ,
    \Tile_X0Y3_E1BEG[2] ,
    \Tile_X0Y3_E1BEG[1] ,
    \Tile_X0Y3_E1BEG[0] }),
    .E2BEG({\Tile_X0Y3_E2BEG[7] ,
    \Tile_X0Y3_E2BEG[6] ,
    \Tile_X0Y3_E2BEG[5] ,
    \Tile_X0Y3_E2BEG[4] ,
    \Tile_X0Y3_E2BEG[3] ,
    \Tile_X0Y3_E2BEG[2] ,
    \Tile_X0Y3_E2BEG[1] ,
    \Tile_X0Y3_E2BEG[0] }),
    .E2BEGb({\Tile_X0Y3_E2BEGb[7] ,
    \Tile_X0Y3_E2BEGb[6] ,
    \Tile_X0Y3_E2BEGb[5] ,
    \Tile_X0Y3_E2BEGb[4] ,
    \Tile_X0Y3_E2BEGb[3] ,
    \Tile_X0Y3_E2BEGb[2] ,
    \Tile_X0Y3_E2BEGb[1] ,
    \Tile_X0Y3_E2BEGb[0] }),
    .E6BEG({\Tile_X0Y3_E6BEG[11] ,
    \Tile_X0Y3_E6BEG[10] ,
    \Tile_X0Y3_E6BEG[9] ,
    \Tile_X0Y3_E6BEG[8] ,
    \Tile_X0Y3_E6BEG[7] ,
    \Tile_X0Y3_E6BEG[6] ,
    \Tile_X0Y3_E6BEG[5] ,
    \Tile_X0Y3_E6BEG[4] ,
    \Tile_X0Y3_E6BEG[3] ,
    \Tile_X0Y3_E6BEG[2] ,
    \Tile_X0Y3_E6BEG[1] ,
    \Tile_X0Y3_E6BEG[0] }),
    .EE4BEG({\Tile_X0Y3_EE4BEG[15] ,
    \Tile_X0Y3_EE4BEG[14] ,
    \Tile_X0Y3_EE4BEG[13] ,
    \Tile_X0Y3_EE4BEG[12] ,
    \Tile_X0Y3_EE4BEG[11] ,
    \Tile_X0Y3_EE4BEG[10] ,
    \Tile_X0Y3_EE4BEG[9] ,
    \Tile_X0Y3_EE4BEG[8] ,
    \Tile_X0Y3_EE4BEG[7] ,
    \Tile_X0Y3_EE4BEG[6] ,
    \Tile_X0Y3_EE4BEG[5] ,
    \Tile_X0Y3_EE4BEG[4] ,
    \Tile_X0Y3_EE4BEG[3] ,
    \Tile_X0Y3_EE4BEG[2] ,
    \Tile_X0Y3_EE4BEG[1] ,
    \Tile_X0Y3_EE4BEG[0] }),
    .FrameData({FrameData[127],
    FrameData[126],
    FrameData[125],
    FrameData[124],
    FrameData[123],
    FrameData[122],
    FrameData[121],
    FrameData[120],
    FrameData[119],
    FrameData[118],
    FrameData[117],
    FrameData[116],
    FrameData[115],
    FrameData[114],
    FrameData[113],
    FrameData[112],
    FrameData[111],
    FrameData[110],
    FrameData[109],
    FrameData[108],
    FrameData[107],
    FrameData[106],
    FrameData[105],
    FrameData[104],
    FrameData[103],
    FrameData[102],
    FrameData[101],
    FrameData[100],
    FrameData[99],
    FrameData[98],
    FrameData[97],
    FrameData[96]}),
    .FrameData_O({\Tile_X0Y3_FrameData_O[31] ,
    \Tile_X0Y3_FrameData_O[30] ,
    \Tile_X0Y3_FrameData_O[29] ,
    \Tile_X0Y3_FrameData_O[28] ,
    \Tile_X0Y3_FrameData_O[27] ,
    \Tile_X0Y3_FrameData_O[26] ,
    \Tile_X0Y3_FrameData_O[25] ,
    \Tile_X0Y3_FrameData_O[24] ,
    \Tile_X0Y3_FrameData_O[23] ,
    \Tile_X0Y3_FrameData_O[22] ,
    \Tile_X0Y3_FrameData_O[21] ,
    \Tile_X0Y3_FrameData_O[20] ,
    \Tile_X0Y3_FrameData_O[19] ,
    \Tile_X0Y3_FrameData_O[18] ,
    \Tile_X0Y3_FrameData_O[17] ,
    \Tile_X0Y3_FrameData_O[16] ,
    \Tile_X0Y3_FrameData_O[15] ,
    \Tile_X0Y3_FrameData_O[14] ,
    \Tile_X0Y3_FrameData_O[13] ,
    \Tile_X0Y3_FrameData_O[12] ,
    \Tile_X0Y3_FrameData_O[11] ,
    \Tile_X0Y3_FrameData_O[10] ,
    \Tile_X0Y3_FrameData_O[9] ,
    \Tile_X0Y3_FrameData_O[8] ,
    \Tile_X0Y3_FrameData_O[7] ,
    \Tile_X0Y3_FrameData_O[6] ,
    \Tile_X0Y3_FrameData_O[5] ,
    \Tile_X0Y3_FrameData_O[4] ,
    \Tile_X0Y3_FrameData_O[3] ,
    \Tile_X0Y3_FrameData_O[2] ,
    \Tile_X0Y3_FrameData_O[1] ,
    \Tile_X0Y3_FrameData_O[0] }),
    .FrameStrobe({\Tile_X0Y4_FrameStrobe_O[19] ,
    \Tile_X0Y4_FrameStrobe_O[18] ,
    \Tile_X0Y4_FrameStrobe_O[17] ,
    \Tile_X0Y4_FrameStrobe_O[16] ,
    \Tile_X0Y4_FrameStrobe_O[15] ,
    \Tile_X0Y4_FrameStrobe_O[14] ,
    \Tile_X0Y4_FrameStrobe_O[13] ,
    \Tile_X0Y4_FrameStrobe_O[12] ,
    \Tile_X0Y4_FrameStrobe_O[11] ,
    \Tile_X0Y4_FrameStrobe_O[10] ,
    \Tile_X0Y4_FrameStrobe_O[9] ,
    \Tile_X0Y4_FrameStrobe_O[8] ,
    \Tile_X0Y4_FrameStrobe_O[7] ,
    \Tile_X0Y4_FrameStrobe_O[6] ,
    \Tile_X0Y4_FrameStrobe_O[5] ,
    \Tile_X0Y4_FrameStrobe_O[4] ,
    \Tile_X0Y4_FrameStrobe_O[3] ,
    \Tile_X0Y4_FrameStrobe_O[2] ,
    \Tile_X0Y4_FrameStrobe_O[1] ,
    \Tile_X0Y4_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X0Y3_FrameStrobe_O[19] ,
    \Tile_X0Y3_FrameStrobe_O[18] ,
    \Tile_X0Y3_FrameStrobe_O[17] ,
    \Tile_X0Y3_FrameStrobe_O[16] ,
    \Tile_X0Y3_FrameStrobe_O[15] ,
    \Tile_X0Y3_FrameStrobe_O[14] ,
    \Tile_X0Y3_FrameStrobe_O[13] ,
    \Tile_X0Y3_FrameStrobe_O[12] ,
    \Tile_X0Y3_FrameStrobe_O[11] ,
    \Tile_X0Y3_FrameStrobe_O[10] ,
    \Tile_X0Y3_FrameStrobe_O[9] ,
    \Tile_X0Y3_FrameStrobe_O[8] ,
    \Tile_X0Y3_FrameStrobe_O[7] ,
    \Tile_X0Y3_FrameStrobe_O[6] ,
    \Tile_X0Y3_FrameStrobe_O[5] ,
    \Tile_X0Y3_FrameStrobe_O[4] ,
    \Tile_X0Y3_FrameStrobe_O[3] ,
    \Tile_X0Y3_FrameStrobe_O[2] ,
    \Tile_X0Y3_FrameStrobe_O[1] ,
    \Tile_X0Y3_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X0Y3_N1BEG[3] ,
    \Tile_X0Y3_N1BEG[2] ,
    \Tile_X0Y3_N1BEG[1] ,
    \Tile_X0Y3_N1BEG[0] }),
    .N1END({\Tile_X0Y4_N1BEG[3] ,
    \Tile_X0Y4_N1BEG[2] ,
    \Tile_X0Y4_N1BEG[1] ,
    \Tile_X0Y4_N1BEG[0] }),
    .N2BEG({\Tile_X0Y3_N2BEG[7] ,
    \Tile_X0Y3_N2BEG[6] ,
    \Tile_X0Y3_N2BEG[5] ,
    \Tile_X0Y3_N2BEG[4] ,
    \Tile_X0Y3_N2BEG[3] ,
    \Tile_X0Y3_N2BEG[2] ,
    \Tile_X0Y3_N2BEG[1] ,
    \Tile_X0Y3_N2BEG[0] }),
    .N2BEGb({\Tile_X0Y3_N2BEGb[7] ,
    \Tile_X0Y3_N2BEGb[6] ,
    \Tile_X0Y3_N2BEGb[5] ,
    \Tile_X0Y3_N2BEGb[4] ,
    \Tile_X0Y3_N2BEGb[3] ,
    \Tile_X0Y3_N2BEGb[2] ,
    \Tile_X0Y3_N2BEGb[1] ,
    \Tile_X0Y3_N2BEGb[0] }),
    .N2END({\Tile_X0Y4_N2BEGb[7] ,
    \Tile_X0Y4_N2BEGb[6] ,
    \Tile_X0Y4_N2BEGb[5] ,
    \Tile_X0Y4_N2BEGb[4] ,
    \Tile_X0Y4_N2BEGb[3] ,
    \Tile_X0Y4_N2BEGb[2] ,
    \Tile_X0Y4_N2BEGb[1] ,
    \Tile_X0Y4_N2BEGb[0] }),
    .N2MID({\Tile_X0Y4_N2BEG[7] ,
    \Tile_X0Y4_N2BEG[6] ,
    \Tile_X0Y4_N2BEG[5] ,
    \Tile_X0Y4_N2BEG[4] ,
    \Tile_X0Y4_N2BEG[3] ,
    \Tile_X0Y4_N2BEG[2] ,
    \Tile_X0Y4_N2BEG[1] ,
    \Tile_X0Y4_N2BEG[0] }),
    .N4BEG({\Tile_X0Y3_N4BEG[15] ,
    \Tile_X0Y3_N4BEG[14] ,
    \Tile_X0Y3_N4BEG[13] ,
    \Tile_X0Y3_N4BEG[12] ,
    \Tile_X0Y3_N4BEG[11] ,
    \Tile_X0Y3_N4BEG[10] ,
    \Tile_X0Y3_N4BEG[9] ,
    \Tile_X0Y3_N4BEG[8] ,
    \Tile_X0Y3_N4BEG[7] ,
    \Tile_X0Y3_N4BEG[6] ,
    \Tile_X0Y3_N4BEG[5] ,
    \Tile_X0Y3_N4BEG[4] ,
    \Tile_X0Y3_N4BEG[3] ,
    \Tile_X0Y3_N4BEG[2] ,
    \Tile_X0Y3_N4BEG[1] ,
    \Tile_X0Y3_N4BEG[0] }),
    .N4END({\Tile_X0Y4_N4BEG[15] ,
    \Tile_X0Y4_N4BEG[14] ,
    \Tile_X0Y4_N4BEG[13] ,
    \Tile_X0Y4_N4BEG[12] ,
    \Tile_X0Y4_N4BEG[11] ,
    \Tile_X0Y4_N4BEG[10] ,
    \Tile_X0Y4_N4BEG[9] ,
    \Tile_X0Y4_N4BEG[8] ,
    \Tile_X0Y4_N4BEG[7] ,
    \Tile_X0Y4_N4BEG[6] ,
    \Tile_X0Y4_N4BEG[5] ,
    \Tile_X0Y4_N4BEG[4] ,
    \Tile_X0Y4_N4BEG[3] ,
    \Tile_X0Y4_N4BEG[2] ,
    \Tile_X0Y4_N4BEG[1] ,
    \Tile_X0Y4_N4BEG[0] }),
    .S1BEG({\Tile_X0Y3_S1BEG[3] ,
    \Tile_X0Y3_S1BEG[2] ,
    \Tile_X0Y3_S1BEG[1] ,
    \Tile_X0Y3_S1BEG[0] }),
    .S1END({\Tile_X0Y2_S1BEG[3] ,
    \Tile_X0Y2_S1BEG[2] ,
    \Tile_X0Y2_S1BEG[1] ,
    \Tile_X0Y2_S1BEG[0] }),
    .S2BEG({\Tile_X0Y3_S2BEG[7] ,
    \Tile_X0Y3_S2BEG[6] ,
    \Tile_X0Y3_S2BEG[5] ,
    \Tile_X0Y3_S2BEG[4] ,
    \Tile_X0Y3_S2BEG[3] ,
    \Tile_X0Y3_S2BEG[2] ,
    \Tile_X0Y3_S2BEG[1] ,
    \Tile_X0Y3_S2BEG[0] }),
    .S2BEGb({\Tile_X0Y3_S2BEGb[7] ,
    \Tile_X0Y3_S2BEGb[6] ,
    \Tile_X0Y3_S2BEGb[5] ,
    \Tile_X0Y3_S2BEGb[4] ,
    \Tile_X0Y3_S2BEGb[3] ,
    \Tile_X0Y3_S2BEGb[2] ,
    \Tile_X0Y3_S2BEGb[1] ,
    \Tile_X0Y3_S2BEGb[0] }),
    .S2END({\Tile_X0Y2_S2BEGb[7] ,
    \Tile_X0Y2_S2BEGb[6] ,
    \Tile_X0Y2_S2BEGb[5] ,
    \Tile_X0Y2_S2BEGb[4] ,
    \Tile_X0Y2_S2BEGb[3] ,
    \Tile_X0Y2_S2BEGb[2] ,
    \Tile_X0Y2_S2BEGb[1] ,
    \Tile_X0Y2_S2BEGb[0] }),
    .S2MID({\Tile_X0Y2_S2BEG[7] ,
    \Tile_X0Y2_S2BEG[6] ,
    \Tile_X0Y2_S2BEG[5] ,
    \Tile_X0Y2_S2BEG[4] ,
    \Tile_X0Y2_S2BEG[3] ,
    \Tile_X0Y2_S2BEG[2] ,
    \Tile_X0Y2_S2BEG[1] ,
    \Tile_X0Y2_S2BEG[0] }),
    .S4BEG({\Tile_X0Y3_S4BEG[15] ,
    \Tile_X0Y3_S4BEG[14] ,
    \Tile_X0Y3_S4BEG[13] ,
    \Tile_X0Y3_S4BEG[12] ,
    \Tile_X0Y3_S4BEG[11] ,
    \Tile_X0Y3_S4BEG[10] ,
    \Tile_X0Y3_S4BEG[9] ,
    \Tile_X0Y3_S4BEG[8] ,
    \Tile_X0Y3_S4BEG[7] ,
    \Tile_X0Y3_S4BEG[6] ,
    \Tile_X0Y3_S4BEG[5] ,
    \Tile_X0Y3_S4BEG[4] ,
    \Tile_X0Y3_S4BEG[3] ,
    \Tile_X0Y3_S4BEG[2] ,
    \Tile_X0Y3_S4BEG[1] ,
    \Tile_X0Y3_S4BEG[0] }),
    .S4END({\Tile_X0Y2_S4BEG[15] ,
    \Tile_X0Y2_S4BEG[14] ,
    \Tile_X0Y2_S4BEG[13] ,
    \Tile_X0Y2_S4BEG[12] ,
    \Tile_X0Y2_S4BEG[11] ,
    \Tile_X0Y2_S4BEG[10] ,
    \Tile_X0Y2_S4BEG[9] ,
    \Tile_X0Y2_S4BEG[8] ,
    \Tile_X0Y2_S4BEG[7] ,
    \Tile_X0Y2_S4BEG[6] ,
    \Tile_X0Y2_S4BEG[5] ,
    \Tile_X0Y2_S4BEG[4] ,
    \Tile_X0Y2_S4BEG[3] ,
    \Tile_X0Y2_S4BEG[2] ,
    \Tile_X0Y2_S4BEG[1] ,
    \Tile_X0Y2_S4BEG[0] }),
    .W1END({\Tile_X1Y3_W1BEG[3] ,
    \Tile_X1Y3_W1BEG[2] ,
    \Tile_X1Y3_W1BEG[1] ,
    \Tile_X1Y3_W1BEG[0] }),
    .W2END({\Tile_X1Y3_W2BEGb[7] ,
    \Tile_X1Y3_W2BEGb[6] ,
    \Tile_X1Y3_W2BEGb[5] ,
    \Tile_X1Y3_W2BEGb[4] ,
    \Tile_X1Y3_W2BEGb[3] ,
    \Tile_X1Y3_W2BEGb[2] ,
    \Tile_X1Y3_W2BEGb[1] ,
    \Tile_X1Y3_W2BEGb[0] }),
    .W2MID({\Tile_X1Y3_W2BEG[7] ,
    \Tile_X1Y3_W2BEG[6] ,
    \Tile_X1Y3_W2BEG[5] ,
    \Tile_X1Y3_W2BEG[4] ,
    \Tile_X1Y3_W2BEG[3] ,
    \Tile_X1Y3_W2BEG[2] ,
    \Tile_X1Y3_W2BEG[1] ,
    \Tile_X1Y3_W2BEG[0] }),
    .W6END({\Tile_X1Y3_W6BEG[11] ,
    \Tile_X1Y3_W6BEG[10] ,
    \Tile_X1Y3_W6BEG[9] ,
    \Tile_X1Y3_W6BEG[8] ,
    \Tile_X1Y3_W6BEG[7] ,
    \Tile_X1Y3_W6BEG[6] ,
    \Tile_X1Y3_W6BEG[5] ,
    \Tile_X1Y3_W6BEG[4] ,
    \Tile_X1Y3_W6BEG[3] ,
    \Tile_X1Y3_W6BEG[2] ,
    \Tile_X1Y3_W6BEG[1] ,
    \Tile_X1Y3_W6BEG[0] }),
    .WW4END({\Tile_X1Y3_WW4BEG[15] ,
    \Tile_X1Y3_WW4BEG[14] ,
    \Tile_X1Y3_WW4BEG[13] ,
    \Tile_X1Y3_WW4BEG[12] ,
    \Tile_X1Y3_WW4BEG[11] ,
    \Tile_X1Y3_WW4BEG[10] ,
    \Tile_X1Y3_WW4BEG[9] ,
    \Tile_X1Y3_WW4BEG[8] ,
    \Tile_X1Y3_WW4BEG[7] ,
    \Tile_X1Y3_WW4BEG[6] ,
    \Tile_X1Y3_WW4BEG[5] ,
    \Tile_X1Y3_WW4BEG[4] ,
    \Tile_X1Y3_WW4BEG[3] ,
    \Tile_X1Y3_WW4BEG[2] ,
    \Tile_X1Y3_WW4BEG[1] ,
    \Tile_X1Y3_WW4BEG[0] }));
 W_TT_IF Tile_X0Y4_W_TT_IF (.CLK_TT_PROJECT(Tile_X0Y4_CLK_TT_PROJECT),
    .ENA_TT_PROJECT(Tile_X0Y4_ENA_TT_PROJECT),
    .RST_N_TT_PROJECT(Tile_X0Y4_RST_N_TT_PROJECT),
    .UIO_IN_TT_PROJECT0(Tile_X0Y4_UIO_IN_TT_PROJECT0),
    .UIO_IN_TT_PROJECT1(Tile_X0Y4_UIO_IN_TT_PROJECT1),
    .UIO_IN_TT_PROJECT2(Tile_X0Y4_UIO_IN_TT_PROJECT2),
    .UIO_IN_TT_PROJECT3(Tile_X0Y4_UIO_IN_TT_PROJECT3),
    .UIO_IN_TT_PROJECT4(Tile_X0Y4_UIO_IN_TT_PROJECT4),
    .UIO_IN_TT_PROJECT5(Tile_X0Y4_UIO_IN_TT_PROJECT5),
    .UIO_IN_TT_PROJECT6(Tile_X0Y4_UIO_IN_TT_PROJECT6),
    .UIO_IN_TT_PROJECT7(Tile_X0Y4_UIO_IN_TT_PROJECT7),
    .UIO_OE_TT_PROJECT0(Tile_X0Y4_UIO_OE_TT_PROJECT0),
    .UIO_OE_TT_PROJECT1(Tile_X0Y4_UIO_OE_TT_PROJECT1),
    .UIO_OE_TT_PROJECT2(Tile_X0Y4_UIO_OE_TT_PROJECT2),
    .UIO_OE_TT_PROJECT3(Tile_X0Y4_UIO_OE_TT_PROJECT3),
    .UIO_OE_TT_PROJECT4(Tile_X0Y4_UIO_OE_TT_PROJECT4),
    .UIO_OE_TT_PROJECT5(Tile_X0Y4_UIO_OE_TT_PROJECT5),
    .UIO_OE_TT_PROJECT6(Tile_X0Y4_UIO_OE_TT_PROJECT6),
    .UIO_OE_TT_PROJECT7(Tile_X0Y4_UIO_OE_TT_PROJECT7),
    .UIO_OUT_TT_PROJECT0(Tile_X0Y4_UIO_OUT_TT_PROJECT0),
    .UIO_OUT_TT_PROJECT1(Tile_X0Y4_UIO_OUT_TT_PROJECT1),
    .UIO_OUT_TT_PROJECT2(Tile_X0Y4_UIO_OUT_TT_PROJECT2),
    .UIO_OUT_TT_PROJECT3(Tile_X0Y4_UIO_OUT_TT_PROJECT3),
    .UIO_OUT_TT_PROJECT4(Tile_X0Y4_UIO_OUT_TT_PROJECT4),
    .UIO_OUT_TT_PROJECT5(Tile_X0Y4_UIO_OUT_TT_PROJECT5),
    .UIO_OUT_TT_PROJECT6(Tile_X0Y4_UIO_OUT_TT_PROJECT6),
    .UIO_OUT_TT_PROJECT7(Tile_X0Y4_UIO_OUT_TT_PROJECT7),
    .UI_IN_TT_PROJECT0(Tile_X0Y4_UI_IN_TT_PROJECT0),
    .UI_IN_TT_PROJECT1(Tile_X0Y4_UI_IN_TT_PROJECT1),
    .UI_IN_TT_PROJECT2(Tile_X0Y4_UI_IN_TT_PROJECT2),
    .UI_IN_TT_PROJECT3(Tile_X0Y4_UI_IN_TT_PROJECT3),
    .UI_IN_TT_PROJECT4(Tile_X0Y4_UI_IN_TT_PROJECT4),
    .UI_IN_TT_PROJECT5(Tile_X0Y4_UI_IN_TT_PROJECT5),
    .UI_IN_TT_PROJECT6(Tile_X0Y4_UI_IN_TT_PROJECT6),
    .UI_IN_TT_PROJECT7(Tile_X0Y4_UI_IN_TT_PROJECT7),
    .UO_OUT_TT_PROJECT0(Tile_X0Y4_UO_OUT_TT_PROJECT0),
    .UO_OUT_TT_PROJECT1(Tile_X0Y4_UO_OUT_TT_PROJECT1),
    .UO_OUT_TT_PROJECT2(Tile_X0Y4_UO_OUT_TT_PROJECT2),
    .UO_OUT_TT_PROJECT3(Tile_X0Y4_UO_OUT_TT_PROJECT3),
    .UO_OUT_TT_PROJECT4(Tile_X0Y4_UO_OUT_TT_PROJECT4),
    .UO_OUT_TT_PROJECT5(Tile_X0Y4_UO_OUT_TT_PROJECT5),
    .UO_OUT_TT_PROJECT6(Tile_X0Y4_UO_OUT_TT_PROJECT6),
    .UO_OUT_TT_PROJECT7(Tile_X0Y4_UO_OUT_TT_PROJECT7),
    .UserCLK(Tile_X0Y5_UserCLKo),
    .UserCLKo(Tile_X0Y4_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X0Y4_E1BEG[3] ,
    \Tile_X0Y4_E1BEG[2] ,
    \Tile_X0Y4_E1BEG[1] ,
    \Tile_X0Y4_E1BEG[0] }),
    .E2BEG({\Tile_X0Y4_E2BEG[7] ,
    \Tile_X0Y4_E2BEG[6] ,
    \Tile_X0Y4_E2BEG[5] ,
    \Tile_X0Y4_E2BEG[4] ,
    \Tile_X0Y4_E2BEG[3] ,
    \Tile_X0Y4_E2BEG[2] ,
    \Tile_X0Y4_E2BEG[1] ,
    \Tile_X0Y4_E2BEG[0] }),
    .E2BEGb({\Tile_X0Y4_E2BEGb[7] ,
    \Tile_X0Y4_E2BEGb[6] ,
    \Tile_X0Y4_E2BEGb[5] ,
    \Tile_X0Y4_E2BEGb[4] ,
    \Tile_X0Y4_E2BEGb[3] ,
    \Tile_X0Y4_E2BEGb[2] ,
    \Tile_X0Y4_E2BEGb[1] ,
    \Tile_X0Y4_E2BEGb[0] }),
    .E6BEG({\Tile_X0Y4_E6BEG[11] ,
    \Tile_X0Y4_E6BEG[10] ,
    \Tile_X0Y4_E6BEG[9] ,
    \Tile_X0Y4_E6BEG[8] ,
    \Tile_X0Y4_E6BEG[7] ,
    \Tile_X0Y4_E6BEG[6] ,
    \Tile_X0Y4_E6BEG[5] ,
    \Tile_X0Y4_E6BEG[4] ,
    \Tile_X0Y4_E6BEG[3] ,
    \Tile_X0Y4_E6BEG[2] ,
    \Tile_X0Y4_E6BEG[1] ,
    \Tile_X0Y4_E6BEG[0] }),
    .EE4BEG({\Tile_X0Y4_EE4BEG[15] ,
    \Tile_X0Y4_EE4BEG[14] ,
    \Tile_X0Y4_EE4BEG[13] ,
    \Tile_X0Y4_EE4BEG[12] ,
    \Tile_X0Y4_EE4BEG[11] ,
    \Tile_X0Y4_EE4BEG[10] ,
    \Tile_X0Y4_EE4BEG[9] ,
    \Tile_X0Y4_EE4BEG[8] ,
    \Tile_X0Y4_EE4BEG[7] ,
    \Tile_X0Y4_EE4BEG[6] ,
    \Tile_X0Y4_EE4BEG[5] ,
    \Tile_X0Y4_EE4BEG[4] ,
    \Tile_X0Y4_EE4BEG[3] ,
    \Tile_X0Y4_EE4BEG[2] ,
    \Tile_X0Y4_EE4BEG[1] ,
    \Tile_X0Y4_EE4BEG[0] }),
    .FrameData({FrameData[159],
    FrameData[158],
    FrameData[157],
    FrameData[156],
    FrameData[155],
    FrameData[154],
    FrameData[153],
    FrameData[152],
    FrameData[151],
    FrameData[150],
    FrameData[149],
    FrameData[148],
    FrameData[147],
    FrameData[146],
    FrameData[145],
    FrameData[144],
    FrameData[143],
    FrameData[142],
    FrameData[141],
    FrameData[140],
    FrameData[139],
    FrameData[138],
    FrameData[137],
    FrameData[136],
    FrameData[135],
    FrameData[134],
    FrameData[133],
    FrameData[132],
    FrameData[131],
    FrameData[130],
    FrameData[129],
    FrameData[128]}),
    .FrameData_O({\Tile_X0Y4_FrameData_O[31] ,
    \Tile_X0Y4_FrameData_O[30] ,
    \Tile_X0Y4_FrameData_O[29] ,
    \Tile_X0Y4_FrameData_O[28] ,
    \Tile_X0Y4_FrameData_O[27] ,
    \Tile_X0Y4_FrameData_O[26] ,
    \Tile_X0Y4_FrameData_O[25] ,
    \Tile_X0Y4_FrameData_O[24] ,
    \Tile_X0Y4_FrameData_O[23] ,
    \Tile_X0Y4_FrameData_O[22] ,
    \Tile_X0Y4_FrameData_O[21] ,
    \Tile_X0Y4_FrameData_O[20] ,
    \Tile_X0Y4_FrameData_O[19] ,
    \Tile_X0Y4_FrameData_O[18] ,
    \Tile_X0Y4_FrameData_O[17] ,
    \Tile_X0Y4_FrameData_O[16] ,
    \Tile_X0Y4_FrameData_O[15] ,
    \Tile_X0Y4_FrameData_O[14] ,
    \Tile_X0Y4_FrameData_O[13] ,
    \Tile_X0Y4_FrameData_O[12] ,
    \Tile_X0Y4_FrameData_O[11] ,
    \Tile_X0Y4_FrameData_O[10] ,
    \Tile_X0Y4_FrameData_O[9] ,
    \Tile_X0Y4_FrameData_O[8] ,
    \Tile_X0Y4_FrameData_O[7] ,
    \Tile_X0Y4_FrameData_O[6] ,
    \Tile_X0Y4_FrameData_O[5] ,
    \Tile_X0Y4_FrameData_O[4] ,
    \Tile_X0Y4_FrameData_O[3] ,
    \Tile_X0Y4_FrameData_O[2] ,
    \Tile_X0Y4_FrameData_O[1] ,
    \Tile_X0Y4_FrameData_O[0] }),
    .FrameStrobe({\Tile_X0Y5_FrameStrobe_O[19] ,
    \Tile_X0Y5_FrameStrobe_O[18] ,
    \Tile_X0Y5_FrameStrobe_O[17] ,
    \Tile_X0Y5_FrameStrobe_O[16] ,
    \Tile_X0Y5_FrameStrobe_O[15] ,
    \Tile_X0Y5_FrameStrobe_O[14] ,
    \Tile_X0Y5_FrameStrobe_O[13] ,
    \Tile_X0Y5_FrameStrobe_O[12] ,
    \Tile_X0Y5_FrameStrobe_O[11] ,
    \Tile_X0Y5_FrameStrobe_O[10] ,
    \Tile_X0Y5_FrameStrobe_O[9] ,
    \Tile_X0Y5_FrameStrobe_O[8] ,
    \Tile_X0Y5_FrameStrobe_O[7] ,
    \Tile_X0Y5_FrameStrobe_O[6] ,
    \Tile_X0Y5_FrameStrobe_O[5] ,
    \Tile_X0Y5_FrameStrobe_O[4] ,
    \Tile_X0Y5_FrameStrobe_O[3] ,
    \Tile_X0Y5_FrameStrobe_O[2] ,
    \Tile_X0Y5_FrameStrobe_O[1] ,
    \Tile_X0Y5_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X0Y4_FrameStrobe_O[19] ,
    \Tile_X0Y4_FrameStrobe_O[18] ,
    \Tile_X0Y4_FrameStrobe_O[17] ,
    \Tile_X0Y4_FrameStrobe_O[16] ,
    \Tile_X0Y4_FrameStrobe_O[15] ,
    \Tile_X0Y4_FrameStrobe_O[14] ,
    \Tile_X0Y4_FrameStrobe_O[13] ,
    \Tile_X0Y4_FrameStrobe_O[12] ,
    \Tile_X0Y4_FrameStrobe_O[11] ,
    \Tile_X0Y4_FrameStrobe_O[10] ,
    \Tile_X0Y4_FrameStrobe_O[9] ,
    \Tile_X0Y4_FrameStrobe_O[8] ,
    \Tile_X0Y4_FrameStrobe_O[7] ,
    \Tile_X0Y4_FrameStrobe_O[6] ,
    \Tile_X0Y4_FrameStrobe_O[5] ,
    \Tile_X0Y4_FrameStrobe_O[4] ,
    \Tile_X0Y4_FrameStrobe_O[3] ,
    \Tile_X0Y4_FrameStrobe_O[2] ,
    \Tile_X0Y4_FrameStrobe_O[1] ,
    \Tile_X0Y4_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X0Y4_N1BEG[3] ,
    \Tile_X0Y4_N1BEG[2] ,
    \Tile_X0Y4_N1BEG[1] ,
    \Tile_X0Y4_N1BEG[0] }),
    .N1END({\Tile_X0Y5_N1BEG[3] ,
    \Tile_X0Y5_N1BEG[2] ,
    \Tile_X0Y5_N1BEG[1] ,
    \Tile_X0Y5_N1BEG[0] }),
    .N2BEG({\Tile_X0Y4_N2BEG[7] ,
    \Tile_X0Y4_N2BEG[6] ,
    \Tile_X0Y4_N2BEG[5] ,
    \Tile_X0Y4_N2BEG[4] ,
    \Tile_X0Y4_N2BEG[3] ,
    \Tile_X0Y4_N2BEG[2] ,
    \Tile_X0Y4_N2BEG[1] ,
    \Tile_X0Y4_N2BEG[0] }),
    .N2BEGb({\Tile_X0Y4_N2BEGb[7] ,
    \Tile_X0Y4_N2BEGb[6] ,
    \Tile_X0Y4_N2BEGb[5] ,
    \Tile_X0Y4_N2BEGb[4] ,
    \Tile_X0Y4_N2BEGb[3] ,
    \Tile_X0Y4_N2BEGb[2] ,
    \Tile_X0Y4_N2BEGb[1] ,
    \Tile_X0Y4_N2BEGb[0] }),
    .N2END({\Tile_X0Y5_N2BEGb[7] ,
    \Tile_X0Y5_N2BEGb[6] ,
    \Tile_X0Y5_N2BEGb[5] ,
    \Tile_X0Y5_N2BEGb[4] ,
    \Tile_X0Y5_N2BEGb[3] ,
    \Tile_X0Y5_N2BEGb[2] ,
    \Tile_X0Y5_N2BEGb[1] ,
    \Tile_X0Y5_N2BEGb[0] }),
    .N2MID({\Tile_X0Y5_N2BEG[7] ,
    \Tile_X0Y5_N2BEG[6] ,
    \Tile_X0Y5_N2BEG[5] ,
    \Tile_X0Y5_N2BEG[4] ,
    \Tile_X0Y5_N2BEG[3] ,
    \Tile_X0Y5_N2BEG[2] ,
    \Tile_X0Y5_N2BEG[1] ,
    \Tile_X0Y5_N2BEG[0] }),
    .N4BEG({\Tile_X0Y4_N4BEG[15] ,
    \Tile_X0Y4_N4BEG[14] ,
    \Tile_X0Y4_N4BEG[13] ,
    \Tile_X0Y4_N4BEG[12] ,
    \Tile_X0Y4_N4BEG[11] ,
    \Tile_X0Y4_N4BEG[10] ,
    \Tile_X0Y4_N4BEG[9] ,
    \Tile_X0Y4_N4BEG[8] ,
    \Tile_X0Y4_N4BEG[7] ,
    \Tile_X0Y4_N4BEG[6] ,
    \Tile_X0Y4_N4BEG[5] ,
    \Tile_X0Y4_N4BEG[4] ,
    \Tile_X0Y4_N4BEG[3] ,
    \Tile_X0Y4_N4BEG[2] ,
    \Tile_X0Y4_N4BEG[1] ,
    \Tile_X0Y4_N4BEG[0] }),
    .N4END({\Tile_X0Y5_N4BEG[15] ,
    \Tile_X0Y5_N4BEG[14] ,
    \Tile_X0Y5_N4BEG[13] ,
    \Tile_X0Y5_N4BEG[12] ,
    \Tile_X0Y5_N4BEG[11] ,
    \Tile_X0Y5_N4BEG[10] ,
    \Tile_X0Y5_N4BEG[9] ,
    \Tile_X0Y5_N4BEG[8] ,
    \Tile_X0Y5_N4BEG[7] ,
    \Tile_X0Y5_N4BEG[6] ,
    \Tile_X0Y5_N4BEG[5] ,
    \Tile_X0Y5_N4BEG[4] ,
    \Tile_X0Y5_N4BEG[3] ,
    \Tile_X0Y5_N4BEG[2] ,
    \Tile_X0Y5_N4BEG[1] ,
    \Tile_X0Y5_N4BEG[0] }),
    .S1BEG({\Tile_X0Y4_S1BEG[3] ,
    \Tile_X0Y4_S1BEG[2] ,
    \Tile_X0Y4_S1BEG[1] ,
    \Tile_X0Y4_S1BEG[0] }),
    .S1END({\Tile_X0Y3_S1BEG[3] ,
    \Tile_X0Y3_S1BEG[2] ,
    \Tile_X0Y3_S1BEG[1] ,
    \Tile_X0Y3_S1BEG[0] }),
    .S2BEG({\Tile_X0Y4_S2BEG[7] ,
    \Tile_X0Y4_S2BEG[6] ,
    \Tile_X0Y4_S2BEG[5] ,
    \Tile_X0Y4_S2BEG[4] ,
    \Tile_X0Y4_S2BEG[3] ,
    \Tile_X0Y4_S2BEG[2] ,
    \Tile_X0Y4_S2BEG[1] ,
    \Tile_X0Y4_S2BEG[0] }),
    .S2BEGb({\Tile_X0Y4_S2BEGb[7] ,
    \Tile_X0Y4_S2BEGb[6] ,
    \Tile_X0Y4_S2BEGb[5] ,
    \Tile_X0Y4_S2BEGb[4] ,
    \Tile_X0Y4_S2BEGb[3] ,
    \Tile_X0Y4_S2BEGb[2] ,
    \Tile_X0Y4_S2BEGb[1] ,
    \Tile_X0Y4_S2BEGb[0] }),
    .S2END({\Tile_X0Y3_S2BEGb[7] ,
    \Tile_X0Y3_S2BEGb[6] ,
    \Tile_X0Y3_S2BEGb[5] ,
    \Tile_X0Y3_S2BEGb[4] ,
    \Tile_X0Y3_S2BEGb[3] ,
    \Tile_X0Y3_S2BEGb[2] ,
    \Tile_X0Y3_S2BEGb[1] ,
    \Tile_X0Y3_S2BEGb[0] }),
    .S2MID({\Tile_X0Y3_S2BEG[7] ,
    \Tile_X0Y3_S2BEG[6] ,
    \Tile_X0Y3_S2BEG[5] ,
    \Tile_X0Y3_S2BEG[4] ,
    \Tile_X0Y3_S2BEG[3] ,
    \Tile_X0Y3_S2BEG[2] ,
    \Tile_X0Y3_S2BEG[1] ,
    \Tile_X0Y3_S2BEG[0] }),
    .S4BEG({\Tile_X0Y4_S4BEG[15] ,
    \Tile_X0Y4_S4BEG[14] ,
    \Tile_X0Y4_S4BEG[13] ,
    \Tile_X0Y4_S4BEG[12] ,
    \Tile_X0Y4_S4BEG[11] ,
    \Tile_X0Y4_S4BEG[10] ,
    \Tile_X0Y4_S4BEG[9] ,
    \Tile_X0Y4_S4BEG[8] ,
    \Tile_X0Y4_S4BEG[7] ,
    \Tile_X0Y4_S4BEG[6] ,
    \Tile_X0Y4_S4BEG[5] ,
    \Tile_X0Y4_S4BEG[4] ,
    \Tile_X0Y4_S4BEG[3] ,
    \Tile_X0Y4_S4BEG[2] ,
    \Tile_X0Y4_S4BEG[1] ,
    \Tile_X0Y4_S4BEG[0] }),
    .S4END({\Tile_X0Y3_S4BEG[15] ,
    \Tile_X0Y3_S4BEG[14] ,
    \Tile_X0Y3_S4BEG[13] ,
    \Tile_X0Y3_S4BEG[12] ,
    \Tile_X0Y3_S4BEG[11] ,
    \Tile_X0Y3_S4BEG[10] ,
    \Tile_X0Y3_S4BEG[9] ,
    \Tile_X0Y3_S4BEG[8] ,
    \Tile_X0Y3_S4BEG[7] ,
    \Tile_X0Y3_S4BEG[6] ,
    \Tile_X0Y3_S4BEG[5] ,
    \Tile_X0Y3_S4BEG[4] ,
    \Tile_X0Y3_S4BEG[3] ,
    \Tile_X0Y3_S4BEG[2] ,
    \Tile_X0Y3_S4BEG[1] ,
    \Tile_X0Y3_S4BEG[0] }),
    .W1END({\Tile_X1Y4_W1BEG[3] ,
    \Tile_X1Y4_W1BEG[2] ,
    \Tile_X1Y4_W1BEG[1] ,
    \Tile_X1Y4_W1BEG[0] }),
    .W2END({\Tile_X1Y4_W2BEGb[7] ,
    \Tile_X1Y4_W2BEGb[6] ,
    \Tile_X1Y4_W2BEGb[5] ,
    \Tile_X1Y4_W2BEGb[4] ,
    \Tile_X1Y4_W2BEGb[3] ,
    \Tile_X1Y4_W2BEGb[2] ,
    \Tile_X1Y4_W2BEGb[1] ,
    \Tile_X1Y4_W2BEGb[0] }),
    .W2MID({\Tile_X1Y4_W2BEG[7] ,
    \Tile_X1Y4_W2BEG[6] ,
    \Tile_X1Y4_W2BEG[5] ,
    \Tile_X1Y4_W2BEG[4] ,
    \Tile_X1Y4_W2BEG[3] ,
    \Tile_X1Y4_W2BEG[2] ,
    \Tile_X1Y4_W2BEG[1] ,
    \Tile_X1Y4_W2BEG[0] }),
    .W6END({\Tile_X1Y4_W6BEG[11] ,
    \Tile_X1Y4_W6BEG[10] ,
    \Tile_X1Y4_W6BEG[9] ,
    \Tile_X1Y4_W6BEG[8] ,
    \Tile_X1Y4_W6BEG[7] ,
    \Tile_X1Y4_W6BEG[6] ,
    \Tile_X1Y4_W6BEG[5] ,
    \Tile_X1Y4_W6BEG[4] ,
    \Tile_X1Y4_W6BEG[3] ,
    \Tile_X1Y4_W6BEG[2] ,
    \Tile_X1Y4_W6BEG[1] ,
    \Tile_X1Y4_W6BEG[0] }),
    .WW4END({\Tile_X1Y4_WW4BEG[15] ,
    \Tile_X1Y4_WW4BEG[14] ,
    \Tile_X1Y4_WW4BEG[13] ,
    \Tile_X1Y4_WW4BEG[12] ,
    \Tile_X1Y4_WW4BEG[11] ,
    \Tile_X1Y4_WW4BEG[10] ,
    \Tile_X1Y4_WW4BEG[9] ,
    \Tile_X1Y4_WW4BEG[8] ,
    \Tile_X1Y4_WW4BEG[7] ,
    \Tile_X1Y4_WW4BEG[6] ,
    \Tile_X1Y4_WW4BEG[5] ,
    \Tile_X1Y4_WW4BEG[4] ,
    \Tile_X1Y4_WW4BEG[3] ,
    \Tile_X1Y4_WW4BEG[2] ,
    \Tile_X1Y4_WW4BEG[1] ,
    \Tile_X1Y4_WW4BEG[0] }));
 W_TT_IF Tile_X0Y5_W_TT_IF (.CLK_TT_PROJECT(Tile_X0Y5_CLK_TT_PROJECT),
    .ENA_TT_PROJECT(Tile_X0Y5_ENA_TT_PROJECT),
    .RST_N_TT_PROJECT(Tile_X0Y5_RST_N_TT_PROJECT),
    .UIO_IN_TT_PROJECT0(Tile_X0Y5_UIO_IN_TT_PROJECT0),
    .UIO_IN_TT_PROJECT1(Tile_X0Y5_UIO_IN_TT_PROJECT1),
    .UIO_IN_TT_PROJECT2(Tile_X0Y5_UIO_IN_TT_PROJECT2),
    .UIO_IN_TT_PROJECT3(Tile_X0Y5_UIO_IN_TT_PROJECT3),
    .UIO_IN_TT_PROJECT4(Tile_X0Y5_UIO_IN_TT_PROJECT4),
    .UIO_IN_TT_PROJECT5(Tile_X0Y5_UIO_IN_TT_PROJECT5),
    .UIO_IN_TT_PROJECT6(Tile_X0Y5_UIO_IN_TT_PROJECT6),
    .UIO_IN_TT_PROJECT7(Tile_X0Y5_UIO_IN_TT_PROJECT7),
    .UIO_OE_TT_PROJECT0(Tile_X0Y5_UIO_OE_TT_PROJECT0),
    .UIO_OE_TT_PROJECT1(Tile_X0Y5_UIO_OE_TT_PROJECT1),
    .UIO_OE_TT_PROJECT2(Tile_X0Y5_UIO_OE_TT_PROJECT2),
    .UIO_OE_TT_PROJECT3(Tile_X0Y5_UIO_OE_TT_PROJECT3),
    .UIO_OE_TT_PROJECT4(Tile_X0Y5_UIO_OE_TT_PROJECT4),
    .UIO_OE_TT_PROJECT5(Tile_X0Y5_UIO_OE_TT_PROJECT5),
    .UIO_OE_TT_PROJECT6(Tile_X0Y5_UIO_OE_TT_PROJECT6),
    .UIO_OE_TT_PROJECT7(Tile_X0Y5_UIO_OE_TT_PROJECT7),
    .UIO_OUT_TT_PROJECT0(Tile_X0Y5_UIO_OUT_TT_PROJECT0),
    .UIO_OUT_TT_PROJECT1(Tile_X0Y5_UIO_OUT_TT_PROJECT1),
    .UIO_OUT_TT_PROJECT2(Tile_X0Y5_UIO_OUT_TT_PROJECT2),
    .UIO_OUT_TT_PROJECT3(Tile_X0Y5_UIO_OUT_TT_PROJECT3),
    .UIO_OUT_TT_PROJECT4(Tile_X0Y5_UIO_OUT_TT_PROJECT4),
    .UIO_OUT_TT_PROJECT5(Tile_X0Y5_UIO_OUT_TT_PROJECT5),
    .UIO_OUT_TT_PROJECT6(Tile_X0Y5_UIO_OUT_TT_PROJECT6),
    .UIO_OUT_TT_PROJECT7(Tile_X0Y5_UIO_OUT_TT_PROJECT7),
    .UI_IN_TT_PROJECT0(Tile_X0Y5_UI_IN_TT_PROJECT0),
    .UI_IN_TT_PROJECT1(Tile_X0Y5_UI_IN_TT_PROJECT1),
    .UI_IN_TT_PROJECT2(Tile_X0Y5_UI_IN_TT_PROJECT2),
    .UI_IN_TT_PROJECT3(Tile_X0Y5_UI_IN_TT_PROJECT3),
    .UI_IN_TT_PROJECT4(Tile_X0Y5_UI_IN_TT_PROJECT4),
    .UI_IN_TT_PROJECT5(Tile_X0Y5_UI_IN_TT_PROJECT5),
    .UI_IN_TT_PROJECT6(Tile_X0Y5_UI_IN_TT_PROJECT6),
    .UI_IN_TT_PROJECT7(Tile_X0Y5_UI_IN_TT_PROJECT7),
    .UO_OUT_TT_PROJECT0(Tile_X0Y5_UO_OUT_TT_PROJECT0),
    .UO_OUT_TT_PROJECT1(Tile_X0Y5_UO_OUT_TT_PROJECT1),
    .UO_OUT_TT_PROJECT2(Tile_X0Y5_UO_OUT_TT_PROJECT2),
    .UO_OUT_TT_PROJECT3(Tile_X0Y5_UO_OUT_TT_PROJECT3),
    .UO_OUT_TT_PROJECT4(Tile_X0Y5_UO_OUT_TT_PROJECT4),
    .UO_OUT_TT_PROJECT5(Tile_X0Y5_UO_OUT_TT_PROJECT5),
    .UO_OUT_TT_PROJECT6(Tile_X0Y5_UO_OUT_TT_PROJECT6),
    .UO_OUT_TT_PROJECT7(Tile_X0Y5_UO_OUT_TT_PROJECT7),
    .UserCLK(Tile_X0Y6_UserCLKo),
    .UserCLKo(Tile_X0Y5_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X0Y5_E1BEG[3] ,
    \Tile_X0Y5_E1BEG[2] ,
    \Tile_X0Y5_E1BEG[1] ,
    \Tile_X0Y5_E1BEG[0] }),
    .E2BEG({\Tile_X0Y5_E2BEG[7] ,
    \Tile_X0Y5_E2BEG[6] ,
    \Tile_X0Y5_E2BEG[5] ,
    \Tile_X0Y5_E2BEG[4] ,
    \Tile_X0Y5_E2BEG[3] ,
    \Tile_X0Y5_E2BEG[2] ,
    \Tile_X0Y5_E2BEG[1] ,
    \Tile_X0Y5_E2BEG[0] }),
    .E2BEGb({\Tile_X0Y5_E2BEGb[7] ,
    \Tile_X0Y5_E2BEGb[6] ,
    \Tile_X0Y5_E2BEGb[5] ,
    \Tile_X0Y5_E2BEGb[4] ,
    \Tile_X0Y5_E2BEGb[3] ,
    \Tile_X0Y5_E2BEGb[2] ,
    \Tile_X0Y5_E2BEGb[1] ,
    \Tile_X0Y5_E2BEGb[0] }),
    .E6BEG({\Tile_X0Y5_E6BEG[11] ,
    \Tile_X0Y5_E6BEG[10] ,
    \Tile_X0Y5_E6BEG[9] ,
    \Tile_X0Y5_E6BEG[8] ,
    \Tile_X0Y5_E6BEG[7] ,
    \Tile_X0Y5_E6BEG[6] ,
    \Tile_X0Y5_E6BEG[5] ,
    \Tile_X0Y5_E6BEG[4] ,
    \Tile_X0Y5_E6BEG[3] ,
    \Tile_X0Y5_E6BEG[2] ,
    \Tile_X0Y5_E6BEG[1] ,
    \Tile_X0Y5_E6BEG[0] }),
    .EE4BEG({\Tile_X0Y5_EE4BEG[15] ,
    \Tile_X0Y5_EE4BEG[14] ,
    \Tile_X0Y5_EE4BEG[13] ,
    \Tile_X0Y5_EE4BEG[12] ,
    \Tile_X0Y5_EE4BEG[11] ,
    \Tile_X0Y5_EE4BEG[10] ,
    \Tile_X0Y5_EE4BEG[9] ,
    \Tile_X0Y5_EE4BEG[8] ,
    \Tile_X0Y5_EE4BEG[7] ,
    \Tile_X0Y5_EE4BEG[6] ,
    \Tile_X0Y5_EE4BEG[5] ,
    \Tile_X0Y5_EE4BEG[4] ,
    \Tile_X0Y5_EE4BEG[3] ,
    \Tile_X0Y5_EE4BEG[2] ,
    \Tile_X0Y5_EE4BEG[1] ,
    \Tile_X0Y5_EE4BEG[0] }),
    .FrameData({FrameData[191],
    FrameData[190],
    FrameData[189],
    FrameData[188],
    FrameData[187],
    FrameData[186],
    FrameData[185],
    FrameData[184],
    FrameData[183],
    FrameData[182],
    FrameData[181],
    FrameData[180],
    FrameData[179],
    FrameData[178],
    FrameData[177],
    FrameData[176],
    FrameData[175],
    FrameData[174],
    FrameData[173],
    FrameData[172],
    FrameData[171],
    FrameData[170],
    FrameData[169],
    FrameData[168],
    FrameData[167],
    FrameData[166],
    FrameData[165],
    FrameData[164],
    FrameData[163],
    FrameData[162],
    FrameData[161],
    FrameData[160]}),
    .FrameData_O({\Tile_X0Y5_FrameData_O[31] ,
    \Tile_X0Y5_FrameData_O[30] ,
    \Tile_X0Y5_FrameData_O[29] ,
    \Tile_X0Y5_FrameData_O[28] ,
    \Tile_X0Y5_FrameData_O[27] ,
    \Tile_X0Y5_FrameData_O[26] ,
    \Tile_X0Y5_FrameData_O[25] ,
    \Tile_X0Y5_FrameData_O[24] ,
    \Tile_X0Y5_FrameData_O[23] ,
    \Tile_X0Y5_FrameData_O[22] ,
    \Tile_X0Y5_FrameData_O[21] ,
    \Tile_X0Y5_FrameData_O[20] ,
    \Tile_X0Y5_FrameData_O[19] ,
    \Tile_X0Y5_FrameData_O[18] ,
    \Tile_X0Y5_FrameData_O[17] ,
    \Tile_X0Y5_FrameData_O[16] ,
    \Tile_X0Y5_FrameData_O[15] ,
    \Tile_X0Y5_FrameData_O[14] ,
    \Tile_X0Y5_FrameData_O[13] ,
    \Tile_X0Y5_FrameData_O[12] ,
    \Tile_X0Y5_FrameData_O[11] ,
    \Tile_X0Y5_FrameData_O[10] ,
    \Tile_X0Y5_FrameData_O[9] ,
    \Tile_X0Y5_FrameData_O[8] ,
    \Tile_X0Y5_FrameData_O[7] ,
    \Tile_X0Y5_FrameData_O[6] ,
    \Tile_X0Y5_FrameData_O[5] ,
    \Tile_X0Y5_FrameData_O[4] ,
    \Tile_X0Y5_FrameData_O[3] ,
    \Tile_X0Y5_FrameData_O[2] ,
    \Tile_X0Y5_FrameData_O[1] ,
    \Tile_X0Y5_FrameData_O[0] }),
    .FrameStrobe({\Tile_X0Y6_FrameStrobe_O[19] ,
    \Tile_X0Y6_FrameStrobe_O[18] ,
    \Tile_X0Y6_FrameStrobe_O[17] ,
    \Tile_X0Y6_FrameStrobe_O[16] ,
    \Tile_X0Y6_FrameStrobe_O[15] ,
    \Tile_X0Y6_FrameStrobe_O[14] ,
    \Tile_X0Y6_FrameStrobe_O[13] ,
    \Tile_X0Y6_FrameStrobe_O[12] ,
    \Tile_X0Y6_FrameStrobe_O[11] ,
    \Tile_X0Y6_FrameStrobe_O[10] ,
    \Tile_X0Y6_FrameStrobe_O[9] ,
    \Tile_X0Y6_FrameStrobe_O[8] ,
    \Tile_X0Y6_FrameStrobe_O[7] ,
    \Tile_X0Y6_FrameStrobe_O[6] ,
    \Tile_X0Y6_FrameStrobe_O[5] ,
    \Tile_X0Y6_FrameStrobe_O[4] ,
    \Tile_X0Y6_FrameStrobe_O[3] ,
    \Tile_X0Y6_FrameStrobe_O[2] ,
    \Tile_X0Y6_FrameStrobe_O[1] ,
    \Tile_X0Y6_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X0Y5_FrameStrobe_O[19] ,
    \Tile_X0Y5_FrameStrobe_O[18] ,
    \Tile_X0Y5_FrameStrobe_O[17] ,
    \Tile_X0Y5_FrameStrobe_O[16] ,
    \Tile_X0Y5_FrameStrobe_O[15] ,
    \Tile_X0Y5_FrameStrobe_O[14] ,
    \Tile_X0Y5_FrameStrobe_O[13] ,
    \Tile_X0Y5_FrameStrobe_O[12] ,
    \Tile_X0Y5_FrameStrobe_O[11] ,
    \Tile_X0Y5_FrameStrobe_O[10] ,
    \Tile_X0Y5_FrameStrobe_O[9] ,
    \Tile_X0Y5_FrameStrobe_O[8] ,
    \Tile_X0Y5_FrameStrobe_O[7] ,
    \Tile_X0Y5_FrameStrobe_O[6] ,
    \Tile_X0Y5_FrameStrobe_O[5] ,
    \Tile_X0Y5_FrameStrobe_O[4] ,
    \Tile_X0Y5_FrameStrobe_O[3] ,
    \Tile_X0Y5_FrameStrobe_O[2] ,
    \Tile_X0Y5_FrameStrobe_O[1] ,
    \Tile_X0Y5_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X0Y5_N1BEG[3] ,
    \Tile_X0Y5_N1BEG[2] ,
    \Tile_X0Y5_N1BEG[1] ,
    \Tile_X0Y5_N1BEG[0] }),
    .N1END({\Tile_X0Y6_N1BEG[3] ,
    \Tile_X0Y6_N1BEG[2] ,
    \Tile_X0Y6_N1BEG[1] ,
    \Tile_X0Y6_N1BEG[0] }),
    .N2BEG({\Tile_X0Y5_N2BEG[7] ,
    \Tile_X0Y5_N2BEG[6] ,
    \Tile_X0Y5_N2BEG[5] ,
    \Tile_X0Y5_N2BEG[4] ,
    \Tile_X0Y5_N2BEG[3] ,
    \Tile_X0Y5_N2BEG[2] ,
    \Tile_X0Y5_N2BEG[1] ,
    \Tile_X0Y5_N2BEG[0] }),
    .N2BEGb({\Tile_X0Y5_N2BEGb[7] ,
    \Tile_X0Y5_N2BEGb[6] ,
    \Tile_X0Y5_N2BEGb[5] ,
    \Tile_X0Y5_N2BEGb[4] ,
    \Tile_X0Y5_N2BEGb[3] ,
    \Tile_X0Y5_N2BEGb[2] ,
    \Tile_X0Y5_N2BEGb[1] ,
    \Tile_X0Y5_N2BEGb[0] }),
    .N2END({\Tile_X0Y6_N2BEGb[7] ,
    \Tile_X0Y6_N2BEGb[6] ,
    \Tile_X0Y6_N2BEGb[5] ,
    \Tile_X0Y6_N2BEGb[4] ,
    \Tile_X0Y6_N2BEGb[3] ,
    \Tile_X0Y6_N2BEGb[2] ,
    \Tile_X0Y6_N2BEGb[1] ,
    \Tile_X0Y6_N2BEGb[0] }),
    .N2MID({\Tile_X0Y6_N2BEG[7] ,
    \Tile_X0Y6_N2BEG[6] ,
    \Tile_X0Y6_N2BEG[5] ,
    \Tile_X0Y6_N2BEG[4] ,
    \Tile_X0Y6_N2BEG[3] ,
    \Tile_X0Y6_N2BEG[2] ,
    \Tile_X0Y6_N2BEG[1] ,
    \Tile_X0Y6_N2BEG[0] }),
    .N4BEG({\Tile_X0Y5_N4BEG[15] ,
    \Tile_X0Y5_N4BEG[14] ,
    \Tile_X0Y5_N4BEG[13] ,
    \Tile_X0Y5_N4BEG[12] ,
    \Tile_X0Y5_N4BEG[11] ,
    \Tile_X0Y5_N4BEG[10] ,
    \Tile_X0Y5_N4BEG[9] ,
    \Tile_X0Y5_N4BEG[8] ,
    \Tile_X0Y5_N4BEG[7] ,
    \Tile_X0Y5_N4BEG[6] ,
    \Tile_X0Y5_N4BEG[5] ,
    \Tile_X0Y5_N4BEG[4] ,
    \Tile_X0Y5_N4BEG[3] ,
    \Tile_X0Y5_N4BEG[2] ,
    \Tile_X0Y5_N4BEG[1] ,
    \Tile_X0Y5_N4BEG[0] }),
    .N4END({\Tile_X0Y6_N4BEG[15] ,
    \Tile_X0Y6_N4BEG[14] ,
    \Tile_X0Y6_N4BEG[13] ,
    \Tile_X0Y6_N4BEG[12] ,
    \Tile_X0Y6_N4BEG[11] ,
    \Tile_X0Y6_N4BEG[10] ,
    \Tile_X0Y6_N4BEG[9] ,
    \Tile_X0Y6_N4BEG[8] ,
    \Tile_X0Y6_N4BEG[7] ,
    \Tile_X0Y6_N4BEG[6] ,
    \Tile_X0Y6_N4BEG[5] ,
    \Tile_X0Y6_N4BEG[4] ,
    \Tile_X0Y6_N4BEG[3] ,
    \Tile_X0Y6_N4BEG[2] ,
    \Tile_X0Y6_N4BEG[1] ,
    \Tile_X0Y6_N4BEG[0] }),
    .S1BEG({\Tile_X0Y5_S1BEG[3] ,
    \Tile_X0Y5_S1BEG[2] ,
    \Tile_X0Y5_S1BEG[1] ,
    \Tile_X0Y5_S1BEG[0] }),
    .S1END({\Tile_X0Y4_S1BEG[3] ,
    \Tile_X0Y4_S1BEG[2] ,
    \Tile_X0Y4_S1BEG[1] ,
    \Tile_X0Y4_S1BEG[0] }),
    .S2BEG({\Tile_X0Y5_S2BEG[7] ,
    \Tile_X0Y5_S2BEG[6] ,
    \Tile_X0Y5_S2BEG[5] ,
    \Tile_X0Y5_S2BEG[4] ,
    \Tile_X0Y5_S2BEG[3] ,
    \Tile_X0Y5_S2BEG[2] ,
    \Tile_X0Y5_S2BEG[1] ,
    \Tile_X0Y5_S2BEG[0] }),
    .S2BEGb({\Tile_X0Y5_S2BEGb[7] ,
    \Tile_X0Y5_S2BEGb[6] ,
    \Tile_X0Y5_S2BEGb[5] ,
    \Tile_X0Y5_S2BEGb[4] ,
    \Tile_X0Y5_S2BEGb[3] ,
    \Tile_X0Y5_S2BEGb[2] ,
    \Tile_X0Y5_S2BEGb[1] ,
    \Tile_X0Y5_S2BEGb[0] }),
    .S2END({\Tile_X0Y4_S2BEGb[7] ,
    \Tile_X0Y4_S2BEGb[6] ,
    \Tile_X0Y4_S2BEGb[5] ,
    \Tile_X0Y4_S2BEGb[4] ,
    \Tile_X0Y4_S2BEGb[3] ,
    \Tile_X0Y4_S2BEGb[2] ,
    \Tile_X0Y4_S2BEGb[1] ,
    \Tile_X0Y4_S2BEGb[0] }),
    .S2MID({\Tile_X0Y4_S2BEG[7] ,
    \Tile_X0Y4_S2BEG[6] ,
    \Tile_X0Y4_S2BEG[5] ,
    \Tile_X0Y4_S2BEG[4] ,
    \Tile_X0Y4_S2BEG[3] ,
    \Tile_X0Y4_S2BEG[2] ,
    \Tile_X0Y4_S2BEG[1] ,
    \Tile_X0Y4_S2BEG[0] }),
    .S4BEG({\Tile_X0Y5_S4BEG[15] ,
    \Tile_X0Y5_S4BEG[14] ,
    \Tile_X0Y5_S4BEG[13] ,
    \Tile_X0Y5_S4BEG[12] ,
    \Tile_X0Y5_S4BEG[11] ,
    \Tile_X0Y5_S4BEG[10] ,
    \Tile_X0Y5_S4BEG[9] ,
    \Tile_X0Y5_S4BEG[8] ,
    \Tile_X0Y5_S4BEG[7] ,
    \Tile_X0Y5_S4BEG[6] ,
    \Tile_X0Y5_S4BEG[5] ,
    \Tile_X0Y5_S4BEG[4] ,
    \Tile_X0Y5_S4BEG[3] ,
    \Tile_X0Y5_S4BEG[2] ,
    \Tile_X0Y5_S4BEG[1] ,
    \Tile_X0Y5_S4BEG[0] }),
    .S4END({\Tile_X0Y4_S4BEG[15] ,
    \Tile_X0Y4_S4BEG[14] ,
    \Tile_X0Y4_S4BEG[13] ,
    \Tile_X0Y4_S4BEG[12] ,
    \Tile_X0Y4_S4BEG[11] ,
    \Tile_X0Y4_S4BEG[10] ,
    \Tile_X0Y4_S4BEG[9] ,
    \Tile_X0Y4_S4BEG[8] ,
    \Tile_X0Y4_S4BEG[7] ,
    \Tile_X0Y4_S4BEG[6] ,
    \Tile_X0Y4_S4BEG[5] ,
    \Tile_X0Y4_S4BEG[4] ,
    \Tile_X0Y4_S4BEG[3] ,
    \Tile_X0Y4_S4BEG[2] ,
    \Tile_X0Y4_S4BEG[1] ,
    \Tile_X0Y4_S4BEG[0] }),
    .W1END({\Tile_X1Y5_W1BEG[3] ,
    \Tile_X1Y5_W1BEG[2] ,
    \Tile_X1Y5_W1BEG[1] ,
    \Tile_X1Y5_W1BEG[0] }),
    .W2END({\Tile_X1Y5_W2BEGb[7] ,
    \Tile_X1Y5_W2BEGb[6] ,
    \Tile_X1Y5_W2BEGb[5] ,
    \Tile_X1Y5_W2BEGb[4] ,
    \Tile_X1Y5_W2BEGb[3] ,
    \Tile_X1Y5_W2BEGb[2] ,
    \Tile_X1Y5_W2BEGb[1] ,
    \Tile_X1Y5_W2BEGb[0] }),
    .W2MID({\Tile_X1Y5_W2BEG[7] ,
    \Tile_X1Y5_W2BEG[6] ,
    \Tile_X1Y5_W2BEG[5] ,
    \Tile_X1Y5_W2BEG[4] ,
    \Tile_X1Y5_W2BEG[3] ,
    \Tile_X1Y5_W2BEG[2] ,
    \Tile_X1Y5_W2BEG[1] ,
    \Tile_X1Y5_W2BEG[0] }),
    .W6END({\Tile_X1Y5_W6BEG[11] ,
    \Tile_X1Y5_W6BEG[10] ,
    \Tile_X1Y5_W6BEG[9] ,
    \Tile_X1Y5_W6BEG[8] ,
    \Tile_X1Y5_W6BEG[7] ,
    \Tile_X1Y5_W6BEG[6] ,
    \Tile_X1Y5_W6BEG[5] ,
    \Tile_X1Y5_W6BEG[4] ,
    \Tile_X1Y5_W6BEG[3] ,
    \Tile_X1Y5_W6BEG[2] ,
    \Tile_X1Y5_W6BEG[1] ,
    \Tile_X1Y5_W6BEG[0] }),
    .WW4END({\Tile_X1Y5_WW4BEG[15] ,
    \Tile_X1Y5_WW4BEG[14] ,
    \Tile_X1Y5_WW4BEG[13] ,
    \Tile_X1Y5_WW4BEG[12] ,
    \Tile_X1Y5_WW4BEG[11] ,
    \Tile_X1Y5_WW4BEG[10] ,
    \Tile_X1Y5_WW4BEG[9] ,
    \Tile_X1Y5_WW4BEG[8] ,
    \Tile_X1Y5_WW4BEG[7] ,
    \Tile_X1Y5_WW4BEG[6] ,
    \Tile_X1Y5_WW4BEG[5] ,
    \Tile_X1Y5_WW4BEG[4] ,
    \Tile_X1Y5_WW4BEG[3] ,
    \Tile_X1Y5_WW4BEG[2] ,
    \Tile_X1Y5_WW4BEG[1] ,
    \Tile_X1Y5_WW4BEG[0] }));
 W_TT_IF Tile_X0Y6_W_TT_IF (.CLK_TT_PROJECT(Tile_X0Y6_CLK_TT_PROJECT),
    .ENA_TT_PROJECT(Tile_X0Y6_ENA_TT_PROJECT),
    .RST_N_TT_PROJECT(Tile_X0Y6_RST_N_TT_PROJECT),
    .UIO_IN_TT_PROJECT0(Tile_X0Y6_UIO_IN_TT_PROJECT0),
    .UIO_IN_TT_PROJECT1(Tile_X0Y6_UIO_IN_TT_PROJECT1),
    .UIO_IN_TT_PROJECT2(Tile_X0Y6_UIO_IN_TT_PROJECT2),
    .UIO_IN_TT_PROJECT3(Tile_X0Y6_UIO_IN_TT_PROJECT3),
    .UIO_IN_TT_PROJECT4(Tile_X0Y6_UIO_IN_TT_PROJECT4),
    .UIO_IN_TT_PROJECT5(Tile_X0Y6_UIO_IN_TT_PROJECT5),
    .UIO_IN_TT_PROJECT6(Tile_X0Y6_UIO_IN_TT_PROJECT6),
    .UIO_IN_TT_PROJECT7(Tile_X0Y6_UIO_IN_TT_PROJECT7),
    .UIO_OE_TT_PROJECT0(Tile_X0Y6_UIO_OE_TT_PROJECT0),
    .UIO_OE_TT_PROJECT1(Tile_X0Y6_UIO_OE_TT_PROJECT1),
    .UIO_OE_TT_PROJECT2(Tile_X0Y6_UIO_OE_TT_PROJECT2),
    .UIO_OE_TT_PROJECT3(Tile_X0Y6_UIO_OE_TT_PROJECT3),
    .UIO_OE_TT_PROJECT4(Tile_X0Y6_UIO_OE_TT_PROJECT4),
    .UIO_OE_TT_PROJECT5(Tile_X0Y6_UIO_OE_TT_PROJECT5),
    .UIO_OE_TT_PROJECT6(Tile_X0Y6_UIO_OE_TT_PROJECT6),
    .UIO_OE_TT_PROJECT7(Tile_X0Y6_UIO_OE_TT_PROJECT7),
    .UIO_OUT_TT_PROJECT0(Tile_X0Y6_UIO_OUT_TT_PROJECT0),
    .UIO_OUT_TT_PROJECT1(Tile_X0Y6_UIO_OUT_TT_PROJECT1),
    .UIO_OUT_TT_PROJECT2(Tile_X0Y6_UIO_OUT_TT_PROJECT2),
    .UIO_OUT_TT_PROJECT3(Tile_X0Y6_UIO_OUT_TT_PROJECT3),
    .UIO_OUT_TT_PROJECT4(Tile_X0Y6_UIO_OUT_TT_PROJECT4),
    .UIO_OUT_TT_PROJECT5(Tile_X0Y6_UIO_OUT_TT_PROJECT5),
    .UIO_OUT_TT_PROJECT6(Tile_X0Y6_UIO_OUT_TT_PROJECT6),
    .UIO_OUT_TT_PROJECT7(Tile_X0Y6_UIO_OUT_TT_PROJECT7),
    .UI_IN_TT_PROJECT0(Tile_X0Y6_UI_IN_TT_PROJECT0),
    .UI_IN_TT_PROJECT1(Tile_X0Y6_UI_IN_TT_PROJECT1),
    .UI_IN_TT_PROJECT2(Tile_X0Y6_UI_IN_TT_PROJECT2),
    .UI_IN_TT_PROJECT3(Tile_X0Y6_UI_IN_TT_PROJECT3),
    .UI_IN_TT_PROJECT4(Tile_X0Y6_UI_IN_TT_PROJECT4),
    .UI_IN_TT_PROJECT5(Tile_X0Y6_UI_IN_TT_PROJECT5),
    .UI_IN_TT_PROJECT6(Tile_X0Y6_UI_IN_TT_PROJECT6),
    .UI_IN_TT_PROJECT7(Tile_X0Y6_UI_IN_TT_PROJECT7),
    .UO_OUT_TT_PROJECT0(Tile_X0Y6_UO_OUT_TT_PROJECT0),
    .UO_OUT_TT_PROJECT1(Tile_X0Y6_UO_OUT_TT_PROJECT1),
    .UO_OUT_TT_PROJECT2(Tile_X0Y6_UO_OUT_TT_PROJECT2),
    .UO_OUT_TT_PROJECT3(Tile_X0Y6_UO_OUT_TT_PROJECT3),
    .UO_OUT_TT_PROJECT4(Tile_X0Y6_UO_OUT_TT_PROJECT4),
    .UO_OUT_TT_PROJECT5(Tile_X0Y6_UO_OUT_TT_PROJECT5),
    .UO_OUT_TT_PROJECT6(Tile_X0Y6_UO_OUT_TT_PROJECT6),
    .UO_OUT_TT_PROJECT7(Tile_X0Y6_UO_OUT_TT_PROJECT7),
    .UserCLK(Tile_X0Y7_UserCLKo),
    .UserCLKo(Tile_X0Y6_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X0Y6_E1BEG[3] ,
    \Tile_X0Y6_E1BEG[2] ,
    \Tile_X0Y6_E1BEG[1] ,
    \Tile_X0Y6_E1BEG[0] }),
    .E2BEG({\Tile_X0Y6_E2BEG[7] ,
    \Tile_X0Y6_E2BEG[6] ,
    \Tile_X0Y6_E2BEG[5] ,
    \Tile_X0Y6_E2BEG[4] ,
    \Tile_X0Y6_E2BEG[3] ,
    \Tile_X0Y6_E2BEG[2] ,
    \Tile_X0Y6_E2BEG[1] ,
    \Tile_X0Y6_E2BEG[0] }),
    .E2BEGb({\Tile_X0Y6_E2BEGb[7] ,
    \Tile_X0Y6_E2BEGb[6] ,
    \Tile_X0Y6_E2BEGb[5] ,
    \Tile_X0Y6_E2BEGb[4] ,
    \Tile_X0Y6_E2BEGb[3] ,
    \Tile_X0Y6_E2BEGb[2] ,
    \Tile_X0Y6_E2BEGb[1] ,
    \Tile_X0Y6_E2BEGb[0] }),
    .E6BEG({\Tile_X0Y6_E6BEG[11] ,
    \Tile_X0Y6_E6BEG[10] ,
    \Tile_X0Y6_E6BEG[9] ,
    \Tile_X0Y6_E6BEG[8] ,
    \Tile_X0Y6_E6BEG[7] ,
    \Tile_X0Y6_E6BEG[6] ,
    \Tile_X0Y6_E6BEG[5] ,
    \Tile_X0Y6_E6BEG[4] ,
    \Tile_X0Y6_E6BEG[3] ,
    \Tile_X0Y6_E6BEG[2] ,
    \Tile_X0Y6_E6BEG[1] ,
    \Tile_X0Y6_E6BEG[0] }),
    .EE4BEG({\Tile_X0Y6_EE4BEG[15] ,
    \Tile_X0Y6_EE4BEG[14] ,
    \Tile_X0Y6_EE4BEG[13] ,
    \Tile_X0Y6_EE4BEG[12] ,
    \Tile_X0Y6_EE4BEG[11] ,
    \Tile_X0Y6_EE4BEG[10] ,
    \Tile_X0Y6_EE4BEG[9] ,
    \Tile_X0Y6_EE4BEG[8] ,
    \Tile_X0Y6_EE4BEG[7] ,
    \Tile_X0Y6_EE4BEG[6] ,
    \Tile_X0Y6_EE4BEG[5] ,
    \Tile_X0Y6_EE4BEG[4] ,
    \Tile_X0Y6_EE4BEG[3] ,
    \Tile_X0Y6_EE4BEG[2] ,
    \Tile_X0Y6_EE4BEG[1] ,
    \Tile_X0Y6_EE4BEG[0] }),
    .FrameData({FrameData[223],
    FrameData[222],
    FrameData[221],
    FrameData[220],
    FrameData[219],
    FrameData[218],
    FrameData[217],
    FrameData[216],
    FrameData[215],
    FrameData[214],
    FrameData[213],
    FrameData[212],
    FrameData[211],
    FrameData[210],
    FrameData[209],
    FrameData[208],
    FrameData[207],
    FrameData[206],
    FrameData[205],
    FrameData[204],
    FrameData[203],
    FrameData[202],
    FrameData[201],
    FrameData[200],
    FrameData[199],
    FrameData[198],
    FrameData[197],
    FrameData[196],
    FrameData[195],
    FrameData[194],
    FrameData[193],
    FrameData[192]}),
    .FrameData_O({\Tile_X0Y6_FrameData_O[31] ,
    \Tile_X0Y6_FrameData_O[30] ,
    \Tile_X0Y6_FrameData_O[29] ,
    \Tile_X0Y6_FrameData_O[28] ,
    \Tile_X0Y6_FrameData_O[27] ,
    \Tile_X0Y6_FrameData_O[26] ,
    \Tile_X0Y6_FrameData_O[25] ,
    \Tile_X0Y6_FrameData_O[24] ,
    \Tile_X0Y6_FrameData_O[23] ,
    \Tile_X0Y6_FrameData_O[22] ,
    \Tile_X0Y6_FrameData_O[21] ,
    \Tile_X0Y6_FrameData_O[20] ,
    \Tile_X0Y6_FrameData_O[19] ,
    \Tile_X0Y6_FrameData_O[18] ,
    \Tile_X0Y6_FrameData_O[17] ,
    \Tile_X0Y6_FrameData_O[16] ,
    \Tile_X0Y6_FrameData_O[15] ,
    \Tile_X0Y6_FrameData_O[14] ,
    \Tile_X0Y6_FrameData_O[13] ,
    \Tile_X0Y6_FrameData_O[12] ,
    \Tile_X0Y6_FrameData_O[11] ,
    \Tile_X0Y6_FrameData_O[10] ,
    \Tile_X0Y6_FrameData_O[9] ,
    \Tile_X0Y6_FrameData_O[8] ,
    \Tile_X0Y6_FrameData_O[7] ,
    \Tile_X0Y6_FrameData_O[6] ,
    \Tile_X0Y6_FrameData_O[5] ,
    \Tile_X0Y6_FrameData_O[4] ,
    \Tile_X0Y6_FrameData_O[3] ,
    \Tile_X0Y6_FrameData_O[2] ,
    \Tile_X0Y6_FrameData_O[1] ,
    \Tile_X0Y6_FrameData_O[0] }),
    .FrameStrobe({\Tile_X0Y7_FrameStrobe_O[19] ,
    \Tile_X0Y7_FrameStrobe_O[18] ,
    \Tile_X0Y7_FrameStrobe_O[17] ,
    \Tile_X0Y7_FrameStrobe_O[16] ,
    \Tile_X0Y7_FrameStrobe_O[15] ,
    \Tile_X0Y7_FrameStrobe_O[14] ,
    \Tile_X0Y7_FrameStrobe_O[13] ,
    \Tile_X0Y7_FrameStrobe_O[12] ,
    \Tile_X0Y7_FrameStrobe_O[11] ,
    \Tile_X0Y7_FrameStrobe_O[10] ,
    \Tile_X0Y7_FrameStrobe_O[9] ,
    \Tile_X0Y7_FrameStrobe_O[8] ,
    \Tile_X0Y7_FrameStrobe_O[7] ,
    \Tile_X0Y7_FrameStrobe_O[6] ,
    \Tile_X0Y7_FrameStrobe_O[5] ,
    \Tile_X0Y7_FrameStrobe_O[4] ,
    \Tile_X0Y7_FrameStrobe_O[3] ,
    \Tile_X0Y7_FrameStrobe_O[2] ,
    \Tile_X0Y7_FrameStrobe_O[1] ,
    \Tile_X0Y7_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X0Y6_FrameStrobe_O[19] ,
    \Tile_X0Y6_FrameStrobe_O[18] ,
    \Tile_X0Y6_FrameStrobe_O[17] ,
    \Tile_X0Y6_FrameStrobe_O[16] ,
    \Tile_X0Y6_FrameStrobe_O[15] ,
    \Tile_X0Y6_FrameStrobe_O[14] ,
    \Tile_X0Y6_FrameStrobe_O[13] ,
    \Tile_X0Y6_FrameStrobe_O[12] ,
    \Tile_X0Y6_FrameStrobe_O[11] ,
    \Tile_X0Y6_FrameStrobe_O[10] ,
    \Tile_X0Y6_FrameStrobe_O[9] ,
    \Tile_X0Y6_FrameStrobe_O[8] ,
    \Tile_X0Y6_FrameStrobe_O[7] ,
    \Tile_X0Y6_FrameStrobe_O[6] ,
    \Tile_X0Y6_FrameStrobe_O[5] ,
    \Tile_X0Y6_FrameStrobe_O[4] ,
    \Tile_X0Y6_FrameStrobe_O[3] ,
    \Tile_X0Y6_FrameStrobe_O[2] ,
    \Tile_X0Y6_FrameStrobe_O[1] ,
    \Tile_X0Y6_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X0Y6_N1BEG[3] ,
    \Tile_X0Y6_N1BEG[2] ,
    \Tile_X0Y6_N1BEG[1] ,
    \Tile_X0Y6_N1BEG[0] }),
    .N1END({\Tile_X0Y7_N1BEG[3] ,
    \Tile_X0Y7_N1BEG[2] ,
    \Tile_X0Y7_N1BEG[1] ,
    \Tile_X0Y7_N1BEG[0] }),
    .N2BEG({\Tile_X0Y6_N2BEG[7] ,
    \Tile_X0Y6_N2BEG[6] ,
    \Tile_X0Y6_N2BEG[5] ,
    \Tile_X0Y6_N2BEG[4] ,
    \Tile_X0Y6_N2BEG[3] ,
    \Tile_X0Y6_N2BEG[2] ,
    \Tile_X0Y6_N2BEG[1] ,
    \Tile_X0Y6_N2BEG[0] }),
    .N2BEGb({\Tile_X0Y6_N2BEGb[7] ,
    \Tile_X0Y6_N2BEGb[6] ,
    \Tile_X0Y6_N2BEGb[5] ,
    \Tile_X0Y6_N2BEGb[4] ,
    \Tile_X0Y6_N2BEGb[3] ,
    \Tile_X0Y6_N2BEGb[2] ,
    \Tile_X0Y6_N2BEGb[1] ,
    \Tile_X0Y6_N2BEGb[0] }),
    .N2END({\Tile_X0Y7_N2BEGb[7] ,
    \Tile_X0Y7_N2BEGb[6] ,
    \Tile_X0Y7_N2BEGb[5] ,
    \Tile_X0Y7_N2BEGb[4] ,
    \Tile_X0Y7_N2BEGb[3] ,
    \Tile_X0Y7_N2BEGb[2] ,
    \Tile_X0Y7_N2BEGb[1] ,
    \Tile_X0Y7_N2BEGb[0] }),
    .N2MID({\Tile_X0Y7_N2BEG[7] ,
    \Tile_X0Y7_N2BEG[6] ,
    \Tile_X0Y7_N2BEG[5] ,
    \Tile_X0Y7_N2BEG[4] ,
    \Tile_X0Y7_N2BEG[3] ,
    \Tile_X0Y7_N2BEG[2] ,
    \Tile_X0Y7_N2BEG[1] ,
    \Tile_X0Y7_N2BEG[0] }),
    .N4BEG({\Tile_X0Y6_N4BEG[15] ,
    \Tile_X0Y6_N4BEG[14] ,
    \Tile_X0Y6_N4BEG[13] ,
    \Tile_X0Y6_N4BEG[12] ,
    \Tile_X0Y6_N4BEG[11] ,
    \Tile_X0Y6_N4BEG[10] ,
    \Tile_X0Y6_N4BEG[9] ,
    \Tile_X0Y6_N4BEG[8] ,
    \Tile_X0Y6_N4BEG[7] ,
    \Tile_X0Y6_N4BEG[6] ,
    \Tile_X0Y6_N4BEG[5] ,
    \Tile_X0Y6_N4BEG[4] ,
    \Tile_X0Y6_N4BEG[3] ,
    \Tile_X0Y6_N4BEG[2] ,
    \Tile_X0Y6_N4BEG[1] ,
    \Tile_X0Y6_N4BEG[0] }),
    .N4END({\Tile_X0Y7_N4BEG[15] ,
    \Tile_X0Y7_N4BEG[14] ,
    \Tile_X0Y7_N4BEG[13] ,
    \Tile_X0Y7_N4BEG[12] ,
    \Tile_X0Y7_N4BEG[11] ,
    \Tile_X0Y7_N4BEG[10] ,
    \Tile_X0Y7_N4BEG[9] ,
    \Tile_X0Y7_N4BEG[8] ,
    \Tile_X0Y7_N4BEG[7] ,
    \Tile_X0Y7_N4BEG[6] ,
    \Tile_X0Y7_N4BEG[5] ,
    \Tile_X0Y7_N4BEG[4] ,
    \Tile_X0Y7_N4BEG[3] ,
    \Tile_X0Y7_N4BEG[2] ,
    \Tile_X0Y7_N4BEG[1] ,
    \Tile_X0Y7_N4BEG[0] }),
    .S1BEG({\Tile_X0Y6_S1BEG[3] ,
    \Tile_X0Y6_S1BEG[2] ,
    \Tile_X0Y6_S1BEG[1] ,
    \Tile_X0Y6_S1BEG[0] }),
    .S1END({\Tile_X0Y5_S1BEG[3] ,
    \Tile_X0Y5_S1BEG[2] ,
    \Tile_X0Y5_S1BEG[1] ,
    \Tile_X0Y5_S1BEG[0] }),
    .S2BEG({\Tile_X0Y6_S2BEG[7] ,
    \Tile_X0Y6_S2BEG[6] ,
    \Tile_X0Y6_S2BEG[5] ,
    \Tile_X0Y6_S2BEG[4] ,
    \Tile_X0Y6_S2BEG[3] ,
    \Tile_X0Y6_S2BEG[2] ,
    \Tile_X0Y6_S2BEG[1] ,
    \Tile_X0Y6_S2BEG[0] }),
    .S2BEGb({\Tile_X0Y6_S2BEGb[7] ,
    \Tile_X0Y6_S2BEGb[6] ,
    \Tile_X0Y6_S2BEGb[5] ,
    \Tile_X0Y6_S2BEGb[4] ,
    \Tile_X0Y6_S2BEGb[3] ,
    \Tile_X0Y6_S2BEGb[2] ,
    \Tile_X0Y6_S2BEGb[1] ,
    \Tile_X0Y6_S2BEGb[0] }),
    .S2END({\Tile_X0Y5_S2BEGb[7] ,
    \Tile_X0Y5_S2BEGb[6] ,
    \Tile_X0Y5_S2BEGb[5] ,
    \Tile_X0Y5_S2BEGb[4] ,
    \Tile_X0Y5_S2BEGb[3] ,
    \Tile_X0Y5_S2BEGb[2] ,
    \Tile_X0Y5_S2BEGb[1] ,
    \Tile_X0Y5_S2BEGb[0] }),
    .S2MID({\Tile_X0Y5_S2BEG[7] ,
    \Tile_X0Y5_S2BEG[6] ,
    \Tile_X0Y5_S2BEG[5] ,
    \Tile_X0Y5_S2BEG[4] ,
    \Tile_X0Y5_S2BEG[3] ,
    \Tile_X0Y5_S2BEG[2] ,
    \Tile_X0Y5_S2BEG[1] ,
    \Tile_X0Y5_S2BEG[0] }),
    .S4BEG({\Tile_X0Y6_S4BEG[15] ,
    \Tile_X0Y6_S4BEG[14] ,
    \Tile_X0Y6_S4BEG[13] ,
    \Tile_X0Y6_S4BEG[12] ,
    \Tile_X0Y6_S4BEG[11] ,
    \Tile_X0Y6_S4BEG[10] ,
    \Tile_X0Y6_S4BEG[9] ,
    \Tile_X0Y6_S4BEG[8] ,
    \Tile_X0Y6_S4BEG[7] ,
    \Tile_X0Y6_S4BEG[6] ,
    \Tile_X0Y6_S4BEG[5] ,
    \Tile_X0Y6_S4BEG[4] ,
    \Tile_X0Y6_S4BEG[3] ,
    \Tile_X0Y6_S4BEG[2] ,
    \Tile_X0Y6_S4BEG[1] ,
    \Tile_X0Y6_S4BEG[0] }),
    .S4END({\Tile_X0Y5_S4BEG[15] ,
    \Tile_X0Y5_S4BEG[14] ,
    \Tile_X0Y5_S4BEG[13] ,
    \Tile_X0Y5_S4BEG[12] ,
    \Tile_X0Y5_S4BEG[11] ,
    \Tile_X0Y5_S4BEG[10] ,
    \Tile_X0Y5_S4BEG[9] ,
    \Tile_X0Y5_S4BEG[8] ,
    \Tile_X0Y5_S4BEG[7] ,
    \Tile_X0Y5_S4BEG[6] ,
    \Tile_X0Y5_S4BEG[5] ,
    \Tile_X0Y5_S4BEG[4] ,
    \Tile_X0Y5_S4BEG[3] ,
    \Tile_X0Y5_S4BEG[2] ,
    \Tile_X0Y5_S4BEG[1] ,
    \Tile_X0Y5_S4BEG[0] }),
    .W1END({\Tile_X1Y6_W1BEG[3] ,
    \Tile_X1Y6_W1BEG[2] ,
    \Tile_X1Y6_W1BEG[1] ,
    \Tile_X1Y6_W1BEG[0] }),
    .W2END({\Tile_X1Y6_W2BEGb[7] ,
    \Tile_X1Y6_W2BEGb[6] ,
    \Tile_X1Y6_W2BEGb[5] ,
    \Tile_X1Y6_W2BEGb[4] ,
    \Tile_X1Y6_W2BEGb[3] ,
    \Tile_X1Y6_W2BEGb[2] ,
    \Tile_X1Y6_W2BEGb[1] ,
    \Tile_X1Y6_W2BEGb[0] }),
    .W2MID({\Tile_X1Y6_W2BEG[7] ,
    \Tile_X1Y6_W2BEG[6] ,
    \Tile_X1Y6_W2BEG[5] ,
    \Tile_X1Y6_W2BEG[4] ,
    \Tile_X1Y6_W2BEG[3] ,
    \Tile_X1Y6_W2BEG[2] ,
    \Tile_X1Y6_W2BEG[1] ,
    \Tile_X1Y6_W2BEG[0] }),
    .W6END({\Tile_X1Y6_W6BEG[11] ,
    \Tile_X1Y6_W6BEG[10] ,
    \Tile_X1Y6_W6BEG[9] ,
    \Tile_X1Y6_W6BEG[8] ,
    \Tile_X1Y6_W6BEG[7] ,
    \Tile_X1Y6_W6BEG[6] ,
    \Tile_X1Y6_W6BEG[5] ,
    \Tile_X1Y6_W6BEG[4] ,
    \Tile_X1Y6_W6BEG[3] ,
    \Tile_X1Y6_W6BEG[2] ,
    \Tile_X1Y6_W6BEG[1] ,
    \Tile_X1Y6_W6BEG[0] }),
    .WW4END({\Tile_X1Y6_WW4BEG[15] ,
    \Tile_X1Y6_WW4BEG[14] ,
    \Tile_X1Y6_WW4BEG[13] ,
    \Tile_X1Y6_WW4BEG[12] ,
    \Tile_X1Y6_WW4BEG[11] ,
    \Tile_X1Y6_WW4BEG[10] ,
    \Tile_X1Y6_WW4BEG[9] ,
    \Tile_X1Y6_WW4BEG[8] ,
    \Tile_X1Y6_WW4BEG[7] ,
    \Tile_X1Y6_WW4BEG[6] ,
    \Tile_X1Y6_WW4BEG[5] ,
    \Tile_X1Y6_WW4BEG[4] ,
    \Tile_X1Y6_WW4BEG[3] ,
    \Tile_X1Y6_WW4BEG[2] ,
    \Tile_X1Y6_WW4BEG[1] ,
    \Tile_X1Y6_WW4BEG[0] }));
 W_TT_IF Tile_X0Y7_W_TT_IF (.CLK_TT_PROJECT(Tile_X0Y7_CLK_TT_PROJECT),
    .ENA_TT_PROJECT(Tile_X0Y7_ENA_TT_PROJECT),
    .RST_N_TT_PROJECT(Tile_X0Y7_RST_N_TT_PROJECT),
    .UIO_IN_TT_PROJECT0(Tile_X0Y7_UIO_IN_TT_PROJECT0),
    .UIO_IN_TT_PROJECT1(Tile_X0Y7_UIO_IN_TT_PROJECT1),
    .UIO_IN_TT_PROJECT2(Tile_X0Y7_UIO_IN_TT_PROJECT2),
    .UIO_IN_TT_PROJECT3(Tile_X0Y7_UIO_IN_TT_PROJECT3),
    .UIO_IN_TT_PROJECT4(Tile_X0Y7_UIO_IN_TT_PROJECT4),
    .UIO_IN_TT_PROJECT5(Tile_X0Y7_UIO_IN_TT_PROJECT5),
    .UIO_IN_TT_PROJECT6(Tile_X0Y7_UIO_IN_TT_PROJECT6),
    .UIO_IN_TT_PROJECT7(Tile_X0Y7_UIO_IN_TT_PROJECT7),
    .UIO_OE_TT_PROJECT0(Tile_X0Y7_UIO_OE_TT_PROJECT0),
    .UIO_OE_TT_PROJECT1(Tile_X0Y7_UIO_OE_TT_PROJECT1),
    .UIO_OE_TT_PROJECT2(Tile_X0Y7_UIO_OE_TT_PROJECT2),
    .UIO_OE_TT_PROJECT3(Tile_X0Y7_UIO_OE_TT_PROJECT3),
    .UIO_OE_TT_PROJECT4(Tile_X0Y7_UIO_OE_TT_PROJECT4),
    .UIO_OE_TT_PROJECT5(Tile_X0Y7_UIO_OE_TT_PROJECT5),
    .UIO_OE_TT_PROJECT6(Tile_X0Y7_UIO_OE_TT_PROJECT6),
    .UIO_OE_TT_PROJECT7(Tile_X0Y7_UIO_OE_TT_PROJECT7),
    .UIO_OUT_TT_PROJECT0(Tile_X0Y7_UIO_OUT_TT_PROJECT0),
    .UIO_OUT_TT_PROJECT1(Tile_X0Y7_UIO_OUT_TT_PROJECT1),
    .UIO_OUT_TT_PROJECT2(Tile_X0Y7_UIO_OUT_TT_PROJECT2),
    .UIO_OUT_TT_PROJECT3(Tile_X0Y7_UIO_OUT_TT_PROJECT3),
    .UIO_OUT_TT_PROJECT4(Tile_X0Y7_UIO_OUT_TT_PROJECT4),
    .UIO_OUT_TT_PROJECT5(Tile_X0Y7_UIO_OUT_TT_PROJECT5),
    .UIO_OUT_TT_PROJECT6(Tile_X0Y7_UIO_OUT_TT_PROJECT6),
    .UIO_OUT_TT_PROJECT7(Tile_X0Y7_UIO_OUT_TT_PROJECT7),
    .UI_IN_TT_PROJECT0(Tile_X0Y7_UI_IN_TT_PROJECT0),
    .UI_IN_TT_PROJECT1(Tile_X0Y7_UI_IN_TT_PROJECT1),
    .UI_IN_TT_PROJECT2(Tile_X0Y7_UI_IN_TT_PROJECT2),
    .UI_IN_TT_PROJECT3(Tile_X0Y7_UI_IN_TT_PROJECT3),
    .UI_IN_TT_PROJECT4(Tile_X0Y7_UI_IN_TT_PROJECT4),
    .UI_IN_TT_PROJECT5(Tile_X0Y7_UI_IN_TT_PROJECT5),
    .UI_IN_TT_PROJECT6(Tile_X0Y7_UI_IN_TT_PROJECT6),
    .UI_IN_TT_PROJECT7(Tile_X0Y7_UI_IN_TT_PROJECT7),
    .UO_OUT_TT_PROJECT0(Tile_X0Y7_UO_OUT_TT_PROJECT0),
    .UO_OUT_TT_PROJECT1(Tile_X0Y7_UO_OUT_TT_PROJECT1),
    .UO_OUT_TT_PROJECT2(Tile_X0Y7_UO_OUT_TT_PROJECT2),
    .UO_OUT_TT_PROJECT3(Tile_X0Y7_UO_OUT_TT_PROJECT3),
    .UO_OUT_TT_PROJECT4(Tile_X0Y7_UO_OUT_TT_PROJECT4),
    .UO_OUT_TT_PROJECT5(Tile_X0Y7_UO_OUT_TT_PROJECT5),
    .UO_OUT_TT_PROJECT6(Tile_X0Y7_UO_OUT_TT_PROJECT6),
    .UO_OUT_TT_PROJECT7(Tile_X0Y7_UO_OUT_TT_PROJECT7),
    .UserCLK(Tile_X0Y8_UserCLKo),
    .UserCLKo(Tile_X0Y7_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X0Y7_E1BEG[3] ,
    \Tile_X0Y7_E1BEG[2] ,
    \Tile_X0Y7_E1BEG[1] ,
    \Tile_X0Y7_E1BEG[0] }),
    .E2BEG({\Tile_X0Y7_E2BEG[7] ,
    \Tile_X0Y7_E2BEG[6] ,
    \Tile_X0Y7_E2BEG[5] ,
    \Tile_X0Y7_E2BEG[4] ,
    \Tile_X0Y7_E2BEG[3] ,
    \Tile_X0Y7_E2BEG[2] ,
    \Tile_X0Y7_E2BEG[1] ,
    \Tile_X0Y7_E2BEG[0] }),
    .E2BEGb({\Tile_X0Y7_E2BEGb[7] ,
    \Tile_X0Y7_E2BEGb[6] ,
    \Tile_X0Y7_E2BEGb[5] ,
    \Tile_X0Y7_E2BEGb[4] ,
    \Tile_X0Y7_E2BEGb[3] ,
    \Tile_X0Y7_E2BEGb[2] ,
    \Tile_X0Y7_E2BEGb[1] ,
    \Tile_X0Y7_E2BEGb[0] }),
    .E6BEG({\Tile_X0Y7_E6BEG[11] ,
    \Tile_X0Y7_E6BEG[10] ,
    \Tile_X0Y7_E6BEG[9] ,
    \Tile_X0Y7_E6BEG[8] ,
    \Tile_X0Y7_E6BEG[7] ,
    \Tile_X0Y7_E6BEG[6] ,
    \Tile_X0Y7_E6BEG[5] ,
    \Tile_X0Y7_E6BEG[4] ,
    \Tile_X0Y7_E6BEG[3] ,
    \Tile_X0Y7_E6BEG[2] ,
    \Tile_X0Y7_E6BEG[1] ,
    \Tile_X0Y7_E6BEG[0] }),
    .EE4BEG({\Tile_X0Y7_EE4BEG[15] ,
    \Tile_X0Y7_EE4BEG[14] ,
    \Tile_X0Y7_EE4BEG[13] ,
    \Tile_X0Y7_EE4BEG[12] ,
    \Tile_X0Y7_EE4BEG[11] ,
    \Tile_X0Y7_EE4BEG[10] ,
    \Tile_X0Y7_EE4BEG[9] ,
    \Tile_X0Y7_EE4BEG[8] ,
    \Tile_X0Y7_EE4BEG[7] ,
    \Tile_X0Y7_EE4BEG[6] ,
    \Tile_X0Y7_EE4BEG[5] ,
    \Tile_X0Y7_EE4BEG[4] ,
    \Tile_X0Y7_EE4BEG[3] ,
    \Tile_X0Y7_EE4BEG[2] ,
    \Tile_X0Y7_EE4BEG[1] ,
    \Tile_X0Y7_EE4BEG[0] }),
    .FrameData({FrameData[255],
    FrameData[254],
    FrameData[253],
    FrameData[252],
    FrameData[251],
    FrameData[250],
    FrameData[249],
    FrameData[248],
    FrameData[247],
    FrameData[246],
    FrameData[245],
    FrameData[244],
    FrameData[243],
    FrameData[242],
    FrameData[241],
    FrameData[240],
    FrameData[239],
    FrameData[238],
    FrameData[237],
    FrameData[236],
    FrameData[235],
    FrameData[234],
    FrameData[233],
    FrameData[232],
    FrameData[231],
    FrameData[230],
    FrameData[229],
    FrameData[228],
    FrameData[227],
    FrameData[226],
    FrameData[225],
    FrameData[224]}),
    .FrameData_O({\Tile_X0Y7_FrameData_O[31] ,
    \Tile_X0Y7_FrameData_O[30] ,
    \Tile_X0Y7_FrameData_O[29] ,
    \Tile_X0Y7_FrameData_O[28] ,
    \Tile_X0Y7_FrameData_O[27] ,
    \Tile_X0Y7_FrameData_O[26] ,
    \Tile_X0Y7_FrameData_O[25] ,
    \Tile_X0Y7_FrameData_O[24] ,
    \Tile_X0Y7_FrameData_O[23] ,
    \Tile_X0Y7_FrameData_O[22] ,
    \Tile_X0Y7_FrameData_O[21] ,
    \Tile_X0Y7_FrameData_O[20] ,
    \Tile_X0Y7_FrameData_O[19] ,
    \Tile_X0Y7_FrameData_O[18] ,
    \Tile_X0Y7_FrameData_O[17] ,
    \Tile_X0Y7_FrameData_O[16] ,
    \Tile_X0Y7_FrameData_O[15] ,
    \Tile_X0Y7_FrameData_O[14] ,
    \Tile_X0Y7_FrameData_O[13] ,
    \Tile_X0Y7_FrameData_O[12] ,
    \Tile_X0Y7_FrameData_O[11] ,
    \Tile_X0Y7_FrameData_O[10] ,
    \Tile_X0Y7_FrameData_O[9] ,
    \Tile_X0Y7_FrameData_O[8] ,
    \Tile_X0Y7_FrameData_O[7] ,
    \Tile_X0Y7_FrameData_O[6] ,
    \Tile_X0Y7_FrameData_O[5] ,
    \Tile_X0Y7_FrameData_O[4] ,
    \Tile_X0Y7_FrameData_O[3] ,
    \Tile_X0Y7_FrameData_O[2] ,
    \Tile_X0Y7_FrameData_O[1] ,
    \Tile_X0Y7_FrameData_O[0] }),
    .FrameStrobe({\Tile_X0Y8_FrameStrobe_O[19] ,
    \Tile_X0Y8_FrameStrobe_O[18] ,
    \Tile_X0Y8_FrameStrobe_O[17] ,
    \Tile_X0Y8_FrameStrobe_O[16] ,
    \Tile_X0Y8_FrameStrobe_O[15] ,
    \Tile_X0Y8_FrameStrobe_O[14] ,
    \Tile_X0Y8_FrameStrobe_O[13] ,
    \Tile_X0Y8_FrameStrobe_O[12] ,
    \Tile_X0Y8_FrameStrobe_O[11] ,
    \Tile_X0Y8_FrameStrobe_O[10] ,
    \Tile_X0Y8_FrameStrobe_O[9] ,
    \Tile_X0Y8_FrameStrobe_O[8] ,
    \Tile_X0Y8_FrameStrobe_O[7] ,
    \Tile_X0Y8_FrameStrobe_O[6] ,
    \Tile_X0Y8_FrameStrobe_O[5] ,
    \Tile_X0Y8_FrameStrobe_O[4] ,
    \Tile_X0Y8_FrameStrobe_O[3] ,
    \Tile_X0Y8_FrameStrobe_O[2] ,
    \Tile_X0Y8_FrameStrobe_O[1] ,
    \Tile_X0Y8_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X0Y7_FrameStrobe_O[19] ,
    \Tile_X0Y7_FrameStrobe_O[18] ,
    \Tile_X0Y7_FrameStrobe_O[17] ,
    \Tile_X0Y7_FrameStrobe_O[16] ,
    \Tile_X0Y7_FrameStrobe_O[15] ,
    \Tile_X0Y7_FrameStrobe_O[14] ,
    \Tile_X0Y7_FrameStrobe_O[13] ,
    \Tile_X0Y7_FrameStrobe_O[12] ,
    \Tile_X0Y7_FrameStrobe_O[11] ,
    \Tile_X0Y7_FrameStrobe_O[10] ,
    \Tile_X0Y7_FrameStrobe_O[9] ,
    \Tile_X0Y7_FrameStrobe_O[8] ,
    \Tile_X0Y7_FrameStrobe_O[7] ,
    \Tile_X0Y7_FrameStrobe_O[6] ,
    \Tile_X0Y7_FrameStrobe_O[5] ,
    \Tile_X0Y7_FrameStrobe_O[4] ,
    \Tile_X0Y7_FrameStrobe_O[3] ,
    \Tile_X0Y7_FrameStrobe_O[2] ,
    \Tile_X0Y7_FrameStrobe_O[1] ,
    \Tile_X0Y7_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X0Y7_N1BEG[3] ,
    \Tile_X0Y7_N1BEG[2] ,
    \Tile_X0Y7_N1BEG[1] ,
    \Tile_X0Y7_N1BEG[0] }),
    .N1END({\Tile_X0Y8_N1BEG[3] ,
    \Tile_X0Y8_N1BEG[2] ,
    \Tile_X0Y8_N1BEG[1] ,
    \Tile_X0Y8_N1BEG[0] }),
    .N2BEG({\Tile_X0Y7_N2BEG[7] ,
    \Tile_X0Y7_N2BEG[6] ,
    \Tile_X0Y7_N2BEG[5] ,
    \Tile_X0Y7_N2BEG[4] ,
    \Tile_X0Y7_N2BEG[3] ,
    \Tile_X0Y7_N2BEG[2] ,
    \Tile_X0Y7_N2BEG[1] ,
    \Tile_X0Y7_N2BEG[0] }),
    .N2BEGb({\Tile_X0Y7_N2BEGb[7] ,
    \Tile_X0Y7_N2BEGb[6] ,
    \Tile_X0Y7_N2BEGb[5] ,
    \Tile_X0Y7_N2BEGb[4] ,
    \Tile_X0Y7_N2BEGb[3] ,
    \Tile_X0Y7_N2BEGb[2] ,
    \Tile_X0Y7_N2BEGb[1] ,
    \Tile_X0Y7_N2BEGb[0] }),
    .N2END({\Tile_X0Y8_N2BEGb[7] ,
    \Tile_X0Y8_N2BEGb[6] ,
    \Tile_X0Y8_N2BEGb[5] ,
    \Tile_X0Y8_N2BEGb[4] ,
    \Tile_X0Y8_N2BEGb[3] ,
    \Tile_X0Y8_N2BEGb[2] ,
    \Tile_X0Y8_N2BEGb[1] ,
    \Tile_X0Y8_N2BEGb[0] }),
    .N2MID({\Tile_X0Y8_N2BEG[7] ,
    \Tile_X0Y8_N2BEG[6] ,
    \Tile_X0Y8_N2BEG[5] ,
    \Tile_X0Y8_N2BEG[4] ,
    \Tile_X0Y8_N2BEG[3] ,
    \Tile_X0Y8_N2BEG[2] ,
    \Tile_X0Y8_N2BEG[1] ,
    \Tile_X0Y8_N2BEG[0] }),
    .N4BEG({\Tile_X0Y7_N4BEG[15] ,
    \Tile_X0Y7_N4BEG[14] ,
    \Tile_X0Y7_N4BEG[13] ,
    \Tile_X0Y7_N4BEG[12] ,
    \Tile_X0Y7_N4BEG[11] ,
    \Tile_X0Y7_N4BEG[10] ,
    \Tile_X0Y7_N4BEG[9] ,
    \Tile_X0Y7_N4BEG[8] ,
    \Tile_X0Y7_N4BEG[7] ,
    \Tile_X0Y7_N4BEG[6] ,
    \Tile_X0Y7_N4BEG[5] ,
    \Tile_X0Y7_N4BEG[4] ,
    \Tile_X0Y7_N4BEG[3] ,
    \Tile_X0Y7_N4BEG[2] ,
    \Tile_X0Y7_N4BEG[1] ,
    \Tile_X0Y7_N4BEG[0] }),
    .N4END({\Tile_X0Y8_N4BEG[15] ,
    \Tile_X0Y8_N4BEG[14] ,
    \Tile_X0Y8_N4BEG[13] ,
    \Tile_X0Y8_N4BEG[12] ,
    \Tile_X0Y8_N4BEG[11] ,
    \Tile_X0Y8_N4BEG[10] ,
    \Tile_X0Y8_N4BEG[9] ,
    \Tile_X0Y8_N4BEG[8] ,
    \Tile_X0Y8_N4BEG[7] ,
    \Tile_X0Y8_N4BEG[6] ,
    \Tile_X0Y8_N4BEG[5] ,
    \Tile_X0Y8_N4BEG[4] ,
    \Tile_X0Y8_N4BEG[3] ,
    \Tile_X0Y8_N4BEG[2] ,
    \Tile_X0Y8_N4BEG[1] ,
    \Tile_X0Y8_N4BEG[0] }),
    .S1BEG({\Tile_X0Y7_S1BEG[3] ,
    \Tile_X0Y7_S1BEG[2] ,
    \Tile_X0Y7_S1BEG[1] ,
    \Tile_X0Y7_S1BEG[0] }),
    .S1END({\Tile_X0Y6_S1BEG[3] ,
    \Tile_X0Y6_S1BEG[2] ,
    \Tile_X0Y6_S1BEG[1] ,
    \Tile_X0Y6_S1BEG[0] }),
    .S2BEG({\Tile_X0Y7_S2BEG[7] ,
    \Tile_X0Y7_S2BEG[6] ,
    \Tile_X0Y7_S2BEG[5] ,
    \Tile_X0Y7_S2BEG[4] ,
    \Tile_X0Y7_S2BEG[3] ,
    \Tile_X0Y7_S2BEG[2] ,
    \Tile_X0Y7_S2BEG[1] ,
    \Tile_X0Y7_S2BEG[0] }),
    .S2BEGb({\Tile_X0Y7_S2BEGb[7] ,
    \Tile_X0Y7_S2BEGb[6] ,
    \Tile_X0Y7_S2BEGb[5] ,
    \Tile_X0Y7_S2BEGb[4] ,
    \Tile_X0Y7_S2BEGb[3] ,
    \Tile_X0Y7_S2BEGb[2] ,
    \Tile_X0Y7_S2BEGb[1] ,
    \Tile_X0Y7_S2BEGb[0] }),
    .S2END({\Tile_X0Y6_S2BEGb[7] ,
    \Tile_X0Y6_S2BEGb[6] ,
    \Tile_X0Y6_S2BEGb[5] ,
    \Tile_X0Y6_S2BEGb[4] ,
    \Tile_X0Y6_S2BEGb[3] ,
    \Tile_X0Y6_S2BEGb[2] ,
    \Tile_X0Y6_S2BEGb[1] ,
    \Tile_X0Y6_S2BEGb[0] }),
    .S2MID({\Tile_X0Y6_S2BEG[7] ,
    \Tile_X0Y6_S2BEG[6] ,
    \Tile_X0Y6_S2BEG[5] ,
    \Tile_X0Y6_S2BEG[4] ,
    \Tile_X0Y6_S2BEG[3] ,
    \Tile_X0Y6_S2BEG[2] ,
    \Tile_X0Y6_S2BEG[1] ,
    \Tile_X0Y6_S2BEG[0] }),
    .S4BEG({\Tile_X0Y7_S4BEG[15] ,
    \Tile_X0Y7_S4BEG[14] ,
    \Tile_X0Y7_S4BEG[13] ,
    \Tile_X0Y7_S4BEG[12] ,
    \Tile_X0Y7_S4BEG[11] ,
    \Tile_X0Y7_S4BEG[10] ,
    \Tile_X0Y7_S4BEG[9] ,
    \Tile_X0Y7_S4BEG[8] ,
    \Tile_X0Y7_S4BEG[7] ,
    \Tile_X0Y7_S4BEG[6] ,
    \Tile_X0Y7_S4BEG[5] ,
    \Tile_X0Y7_S4BEG[4] ,
    \Tile_X0Y7_S4BEG[3] ,
    \Tile_X0Y7_S4BEG[2] ,
    \Tile_X0Y7_S4BEG[1] ,
    \Tile_X0Y7_S4BEG[0] }),
    .S4END({\Tile_X0Y6_S4BEG[15] ,
    \Tile_X0Y6_S4BEG[14] ,
    \Tile_X0Y6_S4BEG[13] ,
    \Tile_X0Y6_S4BEG[12] ,
    \Tile_X0Y6_S4BEG[11] ,
    \Tile_X0Y6_S4BEG[10] ,
    \Tile_X0Y6_S4BEG[9] ,
    \Tile_X0Y6_S4BEG[8] ,
    \Tile_X0Y6_S4BEG[7] ,
    \Tile_X0Y6_S4BEG[6] ,
    \Tile_X0Y6_S4BEG[5] ,
    \Tile_X0Y6_S4BEG[4] ,
    \Tile_X0Y6_S4BEG[3] ,
    \Tile_X0Y6_S4BEG[2] ,
    \Tile_X0Y6_S4BEG[1] ,
    \Tile_X0Y6_S4BEG[0] }),
    .W1END({\Tile_X1Y7_W1BEG[3] ,
    \Tile_X1Y7_W1BEG[2] ,
    \Tile_X1Y7_W1BEG[1] ,
    \Tile_X1Y7_W1BEG[0] }),
    .W2END({\Tile_X1Y7_W2BEGb[7] ,
    \Tile_X1Y7_W2BEGb[6] ,
    \Tile_X1Y7_W2BEGb[5] ,
    \Tile_X1Y7_W2BEGb[4] ,
    \Tile_X1Y7_W2BEGb[3] ,
    \Tile_X1Y7_W2BEGb[2] ,
    \Tile_X1Y7_W2BEGb[1] ,
    \Tile_X1Y7_W2BEGb[0] }),
    .W2MID({\Tile_X1Y7_W2BEG[7] ,
    \Tile_X1Y7_W2BEG[6] ,
    \Tile_X1Y7_W2BEG[5] ,
    \Tile_X1Y7_W2BEG[4] ,
    \Tile_X1Y7_W2BEG[3] ,
    \Tile_X1Y7_W2BEG[2] ,
    \Tile_X1Y7_W2BEG[1] ,
    \Tile_X1Y7_W2BEG[0] }),
    .W6END({\Tile_X1Y7_W6BEG[11] ,
    \Tile_X1Y7_W6BEG[10] ,
    \Tile_X1Y7_W6BEG[9] ,
    \Tile_X1Y7_W6BEG[8] ,
    \Tile_X1Y7_W6BEG[7] ,
    \Tile_X1Y7_W6BEG[6] ,
    \Tile_X1Y7_W6BEG[5] ,
    \Tile_X1Y7_W6BEG[4] ,
    \Tile_X1Y7_W6BEG[3] ,
    \Tile_X1Y7_W6BEG[2] ,
    \Tile_X1Y7_W6BEG[1] ,
    \Tile_X1Y7_W6BEG[0] }),
    .WW4END({\Tile_X1Y7_WW4BEG[15] ,
    \Tile_X1Y7_WW4BEG[14] ,
    \Tile_X1Y7_WW4BEG[13] ,
    \Tile_X1Y7_WW4BEG[12] ,
    \Tile_X1Y7_WW4BEG[11] ,
    \Tile_X1Y7_WW4BEG[10] ,
    \Tile_X1Y7_WW4BEG[9] ,
    \Tile_X1Y7_WW4BEG[8] ,
    \Tile_X1Y7_WW4BEG[7] ,
    \Tile_X1Y7_WW4BEG[6] ,
    \Tile_X1Y7_WW4BEG[5] ,
    \Tile_X1Y7_WW4BEG[4] ,
    \Tile_X1Y7_WW4BEG[3] ,
    \Tile_X1Y7_WW4BEG[2] ,
    \Tile_X1Y7_WW4BEG[1] ,
    \Tile_X1Y7_WW4BEG[0] }));
 W_TT_IF Tile_X0Y8_W_TT_IF (.CLK_TT_PROJECT(Tile_X0Y8_CLK_TT_PROJECT),
    .ENA_TT_PROJECT(Tile_X0Y8_ENA_TT_PROJECT),
    .RST_N_TT_PROJECT(Tile_X0Y8_RST_N_TT_PROJECT),
    .UIO_IN_TT_PROJECT0(Tile_X0Y8_UIO_IN_TT_PROJECT0),
    .UIO_IN_TT_PROJECT1(Tile_X0Y8_UIO_IN_TT_PROJECT1),
    .UIO_IN_TT_PROJECT2(Tile_X0Y8_UIO_IN_TT_PROJECT2),
    .UIO_IN_TT_PROJECT3(Tile_X0Y8_UIO_IN_TT_PROJECT3),
    .UIO_IN_TT_PROJECT4(Tile_X0Y8_UIO_IN_TT_PROJECT4),
    .UIO_IN_TT_PROJECT5(Tile_X0Y8_UIO_IN_TT_PROJECT5),
    .UIO_IN_TT_PROJECT6(Tile_X0Y8_UIO_IN_TT_PROJECT6),
    .UIO_IN_TT_PROJECT7(Tile_X0Y8_UIO_IN_TT_PROJECT7),
    .UIO_OE_TT_PROJECT0(Tile_X0Y8_UIO_OE_TT_PROJECT0),
    .UIO_OE_TT_PROJECT1(Tile_X0Y8_UIO_OE_TT_PROJECT1),
    .UIO_OE_TT_PROJECT2(Tile_X0Y8_UIO_OE_TT_PROJECT2),
    .UIO_OE_TT_PROJECT3(Tile_X0Y8_UIO_OE_TT_PROJECT3),
    .UIO_OE_TT_PROJECT4(Tile_X0Y8_UIO_OE_TT_PROJECT4),
    .UIO_OE_TT_PROJECT5(Tile_X0Y8_UIO_OE_TT_PROJECT5),
    .UIO_OE_TT_PROJECT6(Tile_X0Y8_UIO_OE_TT_PROJECT6),
    .UIO_OE_TT_PROJECT7(Tile_X0Y8_UIO_OE_TT_PROJECT7),
    .UIO_OUT_TT_PROJECT0(Tile_X0Y8_UIO_OUT_TT_PROJECT0),
    .UIO_OUT_TT_PROJECT1(Tile_X0Y8_UIO_OUT_TT_PROJECT1),
    .UIO_OUT_TT_PROJECT2(Tile_X0Y8_UIO_OUT_TT_PROJECT2),
    .UIO_OUT_TT_PROJECT3(Tile_X0Y8_UIO_OUT_TT_PROJECT3),
    .UIO_OUT_TT_PROJECT4(Tile_X0Y8_UIO_OUT_TT_PROJECT4),
    .UIO_OUT_TT_PROJECT5(Tile_X0Y8_UIO_OUT_TT_PROJECT5),
    .UIO_OUT_TT_PROJECT6(Tile_X0Y8_UIO_OUT_TT_PROJECT6),
    .UIO_OUT_TT_PROJECT7(Tile_X0Y8_UIO_OUT_TT_PROJECT7),
    .UI_IN_TT_PROJECT0(Tile_X0Y8_UI_IN_TT_PROJECT0),
    .UI_IN_TT_PROJECT1(Tile_X0Y8_UI_IN_TT_PROJECT1),
    .UI_IN_TT_PROJECT2(Tile_X0Y8_UI_IN_TT_PROJECT2),
    .UI_IN_TT_PROJECT3(Tile_X0Y8_UI_IN_TT_PROJECT3),
    .UI_IN_TT_PROJECT4(Tile_X0Y8_UI_IN_TT_PROJECT4),
    .UI_IN_TT_PROJECT5(Tile_X0Y8_UI_IN_TT_PROJECT5),
    .UI_IN_TT_PROJECT6(Tile_X0Y8_UI_IN_TT_PROJECT6),
    .UI_IN_TT_PROJECT7(Tile_X0Y8_UI_IN_TT_PROJECT7),
    .UO_OUT_TT_PROJECT0(Tile_X0Y8_UO_OUT_TT_PROJECT0),
    .UO_OUT_TT_PROJECT1(Tile_X0Y8_UO_OUT_TT_PROJECT1),
    .UO_OUT_TT_PROJECT2(Tile_X0Y8_UO_OUT_TT_PROJECT2),
    .UO_OUT_TT_PROJECT3(Tile_X0Y8_UO_OUT_TT_PROJECT3),
    .UO_OUT_TT_PROJECT4(Tile_X0Y8_UO_OUT_TT_PROJECT4),
    .UO_OUT_TT_PROJECT5(Tile_X0Y8_UO_OUT_TT_PROJECT5),
    .UO_OUT_TT_PROJECT6(Tile_X0Y8_UO_OUT_TT_PROJECT6),
    .UO_OUT_TT_PROJECT7(Tile_X0Y8_UO_OUT_TT_PROJECT7),
    .UserCLK(Tile_X0Y9_UserCLKo),
    .UserCLKo(Tile_X0Y8_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X0Y8_E1BEG[3] ,
    \Tile_X0Y8_E1BEG[2] ,
    \Tile_X0Y8_E1BEG[1] ,
    \Tile_X0Y8_E1BEG[0] }),
    .E2BEG({\Tile_X0Y8_E2BEG[7] ,
    \Tile_X0Y8_E2BEG[6] ,
    \Tile_X0Y8_E2BEG[5] ,
    \Tile_X0Y8_E2BEG[4] ,
    \Tile_X0Y8_E2BEG[3] ,
    \Tile_X0Y8_E2BEG[2] ,
    \Tile_X0Y8_E2BEG[1] ,
    \Tile_X0Y8_E2BEG[0] }),
    .E2BEGb({\Tile_X0Y8_E2BEGb[7] ,
    \Tile_X0Y8_E2BEGb[6] ,
    \Tile_X0Y8_E2BEGb[5] ,
    \Tile_X0Y8_E2BEGb[4] ,
    \Tile_X0Y8_E2BEGb[3] ,
    \Tile_X0Y8_E2BEGb[2] ,
    \Tile_X0Y8_E2BEGb[1] ,
    \Tile_X0Y8_E2BEGb[0] }),
    .E6BEG({\Tile_X0Y8_E6BEG[11] ,
    \Tile_X0Y8_E6BEG[10] ,
    \Tile_X0Y8_E6BEG[9] ,
    \Tile_X0Y8_E6BEG[8] ,
    \Tile_X0Y8_E6BEG[7] ,
    \Tile_X0Y8_E6BEG[6] ,
    \Tile_X0Y8_E6BEG[5] ,
    \Tile_X0Y8_E6BEG[4] ,
    \Tile_X0Y8_E6BEG[3] ,
    \Tile_X0Y8_E6BEG[2] ,
    \Tile_X0Y8_E6BEG[1] ,
    \Tile_X0Y8_E6BEG[0] }),
    .EE4BEG({\Tile_X0Y8_EE4BEG[15] ,
    \Tile_X0Y8_EE4BEG[14] ,
    \Tile_X0Y8_EE4BEG[13] ,
    \Tile_X0Y8_EE4BEG[12] ,
    \Tile_X0Y8_EE4BEG[11] ,
    \Tile_X0Y8_EE4BEG[10] ,
    \Tile_X0Y8_EE4BEG[9] ,
    \Tile_X0Y8_EE4BEG[8] ,
    \Tile_X0Y8_EE4BEG[7] ,
    \Tile_X0Y8_EE4BEG[6] ,
    \Tile_X0Y8_EE4BEG[5] ,
    \Tile_X0Y8_EE4BEG[4] ,
    \Tile_X0Y8_EE4BEG[3] ,
    \Tile_X0Y8_EE4BEG[2] ,
    \Tile_X0Y8_EE4BEG[1] ,
    \Tile_X0Y8_EE4BEG[0] }),
    .FrameData({FrameData[287],
    FrameData[286],
    FrameData[285],
    FrameData[284],
    FrameData[283],
    FrameData[282],
    FrameData[281],
    FrameData[280],
    FrameData[279],
    FrameData[278],
    FrameData[277],
    FrameData[276],
    FrameData[275],
    FrameData[274],
    FrameData[273],
    FrameData[272],
    FrameData[271],
    FrameData[270],
    FrameData[269],
    FrameData[268],
    FrameData[267],
    FrameData[266],
    FrameData[265],
    FrameData[264],
    FrameData[263],
    FrameData[262],
    FrameData[261],
    FrameData[260],
    FrameData[259],
    FrameData[258],
    FrameData[257],
    FrameData[256]}),
    .FrameData_O({\Tile_X0Y8_FrameData_O[31] ,
    \Tile_X0Y8_FrameData_O[30] ,
    \Tile_X0Y8_FrameData_O[29] ,
    \Tile_X0Y8_FrameData_O[28] ,
    \Tile_X0Y8_FrameData_O[27] ,
    \Tile_X0Y8_FrameData_O[26] ,
    \Tile_X0Y8_FrameData_O[25] ,
    \Tile_X0Y8_FrameData_O[24] ,
    \Tile_X0Y8_FrameData_O[23] ,
    \Tile_X0Y8_FrameData_O[22] ,
    \Tile_X0Y8_FrameData_O[21] ,
    \Tile_X0Y8_FrameData_O[20] ,
    \Tile_X0Y8_FrameData_O[19] ,
    \Tile_X0Y8_FrameData_O[18] ,
    \Tile_X0Y8_FrameData_O[17] ,
    \Tile_X0Y8_FrameData_O[16] ,
    \Tile_X0Y8_FrameData_O[15] ,
    \Tile_X0Y8_FrameData_O[14] ,
    \Tile_X0Y8_FrameData_O[13] ,
    \Tile_X0Y8_FrameData_O[12] ,
    \Tile_X0Y8_FrameData_O[11] ,
    \Tile_X0Y8_FrameData_O[10] ,
    \Tile_X0Y8_FrameData_O[9] ,
    \Tile_X0Y8_FrameData_O[8] ,
    \Tile_X0Y8_FrameData_O[7] ,
    \Tile_X0Y8_FrameData_O[6] ,
    \Tile_X0Y8_FrameData_O[5] ,
    \Tile_X0Y8_FrameData_O[4] ,
    \Tile_X0Y8_FrameData_O[3] ,
    \Tile_X0Y8_FrameData_O[2] ,
    \Tile_X0Y8_FrameData_O[1] ,
    \Tile_X0Y8_FrameData_O[0] }),
    .FrameStrobe({\Tile_X0Y9_FrameStrobe_O[19] ,
    \Tile_X0Y9_FrameStrobe_O[18] ,
    \Tile_X0Y9_FrameStrobe_O[17] ,
    \Tile_X0Y9_FrameStrobe_O[16] ,
    \Tile_X0Y9_FrameStrobe_O[15] ,
    \Tile_X0Y9_FrameStrobe_O[14] ,
    \Tile_X0Y9_FrameStrobe_O[13] ,
    \Tile_X0Y9_FrameStrobe_O[12] ,
    \Tile_X0Y9_FrameStrobe_O[11] ,
    \Tile_X0Y9_FrameStrobe_O[10] ,
    \Tile_X0Y9_FrameStrobe_O[9] ,
    \Tile_X0Y9_FrameStrobe_O[8] ,
    \Tile_X0Y9_FrameStrobe_O[7] ,
    \Tile_X0Y9_FrameStrobe_O[6] ,
    \Tile_X0Y9_FrameStrobe_O[5] ,
    \Tile_X0Y9_FrameStrobe_O[4] ,
    \Tile_X0Y9_FrameStrobe_O[3] ,
    \Tile_X0Y9_FrameStrobe_O[2] ,
    \Tile_X0Y9_FrameStrobe_O[1] ,
    \Tile_X0Y9_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X0Y8_FrameStrobe_O[19] ,
    \Tile_X0Y8_FrameStrobe_O[18] ,
    \Tile_X0Y8_FrameStrobe_O[17] ,
    \Tile_X0Y8_FrameStrobe_O[16] ,
    \Tile_X0Y8_FrameStrobe_O[15] ,
    \Tile_X0Y8_FrameStrobe_O[14] ,
    \Tile_X0Y8_FrameStrobe_O[13] ,
    \Tile_X0Y8_FrameStrobe_O[12] ,
    \Tile_X0Y8_FrameStrobe_O[11] ,
    \Tile_X0Y8_FrameStrobe_O[10] ,
    \Tile_X0Y8_FrameStrobe_O[9] ,
    \Tile_X0Y8_FrameStrobe_O[8] ,
    \Tile_X0Y8_FrameStrobe_O[7] ,
    \Tile_X0Y8_FrameStrobe_O[6] ,
    \Tile_X0Y8_FrameStrobe_O[5] ,
    \Tile_X0Y8_FrameStrobe_O[4] ,
    \Tile_X0Y8_FrameStrobe_O[3] ,
    \Tile_X0Y8_FrameStrobe_O[2] ,
    \Tile_X0Y8_FrameStrobe_O[1] ,
    \Tile_X0Y8_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X0Y8_N1BEG[3] ,
    \Tile_X0Y8_N1BEG[2] ,
    \Tile_X0Y8_N1BEG[1] ,
    \Tile_X0Y8_N1BEG[0] }),
    .N1END({\Tile_X0Y9_N1BEG[3] ,
    \Tile_X0Y9_N1BEG[2] ,
    \Tile_X0Y9_N1BEG[1] ,
    \Tile_X0Y9_N1BEG[0] }),
    .N2BEG({\Tile_X0Y8_N2BEG[7] ,
    \Tile_X0Y8_N2BEG[6] ,
    \Tile_X0Y8_N2BEG[5] ,
    \Tile_X0Y8_N2BEG[4] ,
    \Tile_X0Y8_N2BEG[3] ,
    \Tile_X0Y8_N2BEG[2] ,
    \Tile_X0Y8_N2BEG[1] ,
    \Tile_X0Y8_N2BEG[0] }),
    .N2BEGb({\Tile_X0Y8_N2BEGb[7] ,
    \Tile_X0Y8_N2BEGb[6] ,
    \Tile_X0Y8_N2BEGb[5] ,
    \Tile_X0Y8_N2BEGb[4] ,
    \Tile_X0Y8_N2BEGb[3] ,
    \Tile_X0Y8_N2BEGb[2] ,
    \Tile_X0Y8_N2BEGb[1] ,
    \Tile_X0Y8_N2BEGb[0] }),
    .N2END({\Tile_X0Y9_N2BEGb[7] ,
    \Tile_X0Y9_N2BEGb[6] ,
    \Tile_X0Y9_N2BEGb[5] ,
    \Tile_X0Y9_N2BEGb[4] ,
    \Tile_X0Y9_N2BEGb[3] ,
    \Tile_X0Y9_N2BEGb[2] ,
    \Tile_X0Y9_N2BEGb[1] ,
    \Tile_X0Y9_N2BEGb[0] }),
    .N2MID({\Tile_X0Y9_N2BEG[7] ,
    \Tile_X0Y9_N2BEG[6] ,
    \Tile_X0Y9_N2BEG[5] ,
    \Tile_X0Y9_N2BEG[4] ,
    \Tile_X0Y9_N2BEG[3] ,
    \Tile_X0Y9_N2BEG[2] ,
    \Tile_X0Y9_N2BEG[1] ,
    \Tile_X0Y9_N2BEG[0] }),
    .N4BEG({\Tile_X0Y8_N4BEG[15] ,
    \Tile_X0Y8_N4BEG[14] ,
    \Tile_X0Y8_N4BEG[13] ,
    \Tile_X0Y8_N4BEG[12] ,
    \Tile_X0Y8_N4BEG[11] ,
    \Tile_X0Y8_N4BEG[10] ,
    \Tile_X0Y8_N4BEG[9] ,
    \Tile_X0Y8_N4BEG[8] ,
    \Tile_X0Y8_N4BEG[7] ,
    \Tile_X0Y8_N4BEG[6] ,
    \Tile_X0Y8_N4BEG[5] ,
    \Tile_X0Y8_N4BEG[4] ,
    \Tile_X0Y8_N4BEG[3] ,
    \Tile_X0Y8_N4BEG[2] ,
    \Tile_X0Y8_N4BEG[1] ,
    \Tile_X0Y8_N4BEG[0] }),
    .N4END({\Tile_X0Y9_N4BEG[15] ,
    \Tile_X0Y9_N4BEG[14] ,
    \Tile_X0Y9_N4BEG[13] ,
    \Tile_X0Y9_N4BEG[12] ,
    \Tile_X0Y9_N4BEG[11] ,
    \Tile_X0Y9_N4BEG[10] ,
    \Tile_X0Y9_N4BEG[9] ,
    \Tile_X0Y9_N4BEG[8] ,
    \Tile_X0Y9_N4BEG[7] ,
    \Tile_X0Y9_N4BEG[6] ,
    \Tile_X0Y9_N4BEG[5] ,
    \Tile_X0Y9_N4BEG[4] ,
    \Tile_X0Y9_N4BEG[3] ,
    \Tile_X0Y9_N4BEG[2] ,
    \Tile_X0Y9_N4BEG[1] ,
    \Tile_X0Y9_N4BEG[0] }),
    .S1BEG({\Tile_X0Y8_S1BEG[3] ,
    \Tile_X0Y8_S1BEG[2] ,
    \Tile_X0Y8_S1BEG[1] ,
    \Tile_X0Y8_S1BEG[0] }),
    .S1END({\Tile_X0Y7_S1BEG[3] ,
    \Tile_X0Y7_S1BEG[2] ,
    \Tile_X0Y7_S1BEG[1] ,
    \Tile_X0Y7_S1BEG[0] }),
    .S2BEG({\Tile_X0Y8_S2BEG[7] ,
    \Tile_X0Y8_S2BEG[6] ,
    \Tile_X0Y8_S2BEG[5] ,
    \Tile_X0Y8_S2BEG[4] ,
    \Tile_X0Y8_S2BEG[3] ,
    \Tile_X0Y8_S2BEG[2] ,
    \Tile_X0Y8_S2BEG[1] ,
    \Tile_X0Y8_S2BEG[0] }),
    .S2BEGb({\Tile_X0Y8_S2BEGb[7] ,
    \Tile_X0Y8_S2BEGb[6] ,
    \Tile_X0Y8_S2BEGb[5] ,
    \Tile_X0Y8_S2BEGb[4] ,
    \Tile_X0Y8_S2BEGb[3] ,
    \Tile_X0Y8_S2BEGb[2] ,
    \Tile_X0Y8_S2BEGb[1] ,
    \Tile_X0Y8_S2BEGb[0] }),
    .S2END({\Tile_X0Y7_S2BEGb[7] ,
    \Tile_X0Y7_S2BEGb[6] ,
    \Tile_X0Y7_S2BEGb[5] ,
    \Tile_X0Y7_S2BEGb[4] ,
    \Tile_X0Y7_S2BEGb[3] ,
    \Tile_X0Y7_S2BEGb[2] ,
    \Tile_X0Y7_S2BEGb[1] ,
    \Tile_X0Y7_S2BEGb[0] }),
    .S2MID({\Tile_X0Y7_S2BEG[7] ,
    \Tile_X0Y7_S2BEG[6] ,
    \Tile_X0Y7_S2BEG[5] ,
    \Tile_X0Y7_S2BEG[4] ,
    \Tile_X0Y7_S2BEG[3] ,
    \Tile_X0Y7_S2BEG[2] ,
    \Tile_X0Y7_S2BEG[1] ,
    \Tile_X0Y7_S2BEG[0] }),
    .S4BEG({\Tile_X0Y8_S4BEG[15] ,
    \Tile_X0Y8_S4BEG[14] ,
    \Tile_X0Y8_S4BEG[13] ,
    \Tile_X0Y8_S4BEG[12] ,
    \Tile_X0Y8_S4BEG[11] ,
    \Tile_X0Y8_S4BEG[10] ,
    \Tile_X0Y8_S4BEG[9] ,
    \Tile_X0Y8_S4BEG[8] ,
    \Tile_X0Y8_S4BEG[7] ,
    \Tile_X0Y8_S4BEG[6] ,
    \Tile_X0Y8_S4BEG[5] ,
    \Tile_X0Y8_S4BEG[4] ,
    \Tile_X0Y8_S4BEG[3] ,
    \Tile_X0Y8_S4BEG[2] ,
    \Tile_X0Y8_S4BEG[1] ,
    \Tile_X0Y8_S4BEG[0] }),
    .S4END({\Tile_X0Y7_S4BEG[15] ,
    \Tile_X0Y7_S4BEG[14] ,
    \Tile_X0Y7_S4BEG[13] ,
    \Tile_X0Y7_S4BEG[12] ,
    \Tile_X0Y7_S4BEG[11] ,
    \Tile_X0Y7_S4BEG[10] ,
    \Tile_X0Y7_S4BEG[9] ,
    \Tile_X0Y7_S4BEG[8] ,
    \Tile_X0Y7_S4BEG[7] ,
    \Tile_X0Y7_S4BEG[6] ,
    \Tile_X0Y7_S4BEG[5] ,
    \Tile_X0Y7_S4BEG[4] ,
    \Tile_X0Y7_S4BEG[3] ,
    \Tile_X0Y7_S4BEG[2] ,
    \Tile_X0Y7_S4BEG[1] ,
    \Tile_X0Y7_S4BEG[0] }),
    .W1END({\Tile_X1Y8_W1BEG[3] ,
    \Tile_X1Y8_W1BEG[2] ,
    \Tile_X1Y8_W1BEG[1] ,
    \Tile_X1Y8_W1BEG[0] }),
    .W2END({\Tile_X1Y8_W2BEGb[7] ,
    \Tile_X1Y8_W2BEGb[6] ,
    \Tile_X1Y8_W2BEGb[5] ,
    \Tile_X1Y8_W2BEGb[4] ,
    \Tile_X1Y8_W2BEGb[3] ,
    \Tile_X1Y8_W2BEGb[2] ,
    \Tile_X1Y8_W2BEGb[1] ,
    \Tile_X1Y8_W2BEGb[0] }),
    .W2MID({\Tile_X1Y8_W2BEG[7] ,
    \Tile_X1Y8_W2BEG[6] ,
    \Tile_X1Y8_W2BEG[5] ,
    \Tile_X1Y8_W2BEG[4] ,
    \Tile_X1Y8_W2BEG[3] ,
    \Tile_X1Y8_W2BEG[2] ,
    \Tile_X1Y8_W2BEG[1] ,
    \Tile_X1Y8_W2BEG[0] }),
    .W6END({\Tile_X1Y8_W6BEG[11] ,
    \Tile_X1Y8_W6BEG[10] ,
    \Tile_X1Y8_W6BEG[9] ,
    \Tile_X1Y8_W6BEG[8] ,
    \Tile_X1Y8_W6BEG[7] ,
    \Tile_X1Y8_W6BEG[6] ,
    \Tile_X1Y8_W6BEG[5] ,
    \Tile_X1Y8_W6BEG[4] ,
    \Tile_X1Y8_W6BEG[3] ,
    \Tile_X1Y8_W6BEG[2] ,
    \Tile_X1Y8_W6BEG[1] ,
    \Tile_X1Y8_W6BEG[0] }),
    .WW4END({\Tile_X1Y8_WW4BEG[15] ,
    \Tile_X1Y8_WW4BEG[14] ,
    \Tile_X1Y8_WW4BEG[13] ,
    \Tile_X1Y8_WW4BEG[12] ,
    \Tile_X1Y8_WW4BEG[11] ,
    \Tile_X1Y8_WW4BEG[10] ,
    \Tile_X1Y8_WW4BEG[9] ,
    \Tile_X1Y8_WW4BEG[8] ,
    \Tile_X1Y8_WW4BEG[7] ,
    \Tile_X1Y8_WW4BEG[6] ,
    \Tile_X1Y8_WW4BEG[5] ,
    \Tile_X1Y8_WW4BEG[4] ,
    \Tile_X1Y8_WW4BEG[3] ,
    \Tile_X1Y8_WW4BEG[2] ,
    \Tile_X1Y8_WW4BEG[1] ,
    \Tile_X1Y8_WW4BEG[0] }));
 SW_term Tile_X0Y9_SW_term (.UserCLK(UserCLK),
    .UserCLKo(Tile_X0Y9_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .FrameData({FrameData[319],
    FrameData[318],
    FrameData[317],
    FrameData[316],
    FrameData[315],
    FrameData[314],
    FrameData[313],
    FrameData[312],
    FrameData[311],
    FrameData[310],
    FrameData[309],
    FrameData[308],
    FrameData[307],
    FrameData[306],
    FrameData[305],
    FrameData[304],
    FrameData[303],
    FrameData[302],
    FrameData[301],
    FrameData[300],
    FrameData[299],
    FrameData[298],
    FrameData[297],
    FrameData[296],
    FrameData[295],
    FrameData[294],
    FrameData[293],
    FrameData[292],
    FrameData[291],
    FrameData[290],
    FrameData[289],
    FrameData[288]}),
    .FrameData_O({\Tile_X0Y9_FrameData_O[31] ,
    \Tile_X0Y9_FrameData_O[30] ,
    \Tile_X0Y9_FrameData_O[29] ,
    \Tile_X0Y9_FrameData_O[28] ,
    \Tile_X0Y9_FrameData_O[27] ,
    \Tile_X0Y9_FrameData_O[26] ,
    \Tile_X0Y9_FrameData_O[25] ,
    \Tile_X0Y9_FrameData_O[24] ,
    \Tile_X0Y9_FrameData_O[23] ,
    \Tile_X0Y9_FrameData_O[22] ,
    \Tile_X0Y9_FrameData_O[21] ,
    \Tile_X0Y9_FrameData_O[20] ,
    \Tile_X0Y9_FrameData_O[19] ,
    \Tile_X0Y9_FrameData_O[18] ,
    \Tile_X0Y9_FrameData_O[17] ,
    \Tile_X0Y9_FrameData_O[16] ,
    \Tile_X0Y9_FrameData_O[15] ,
    \Tile_X0Y9_FrameData_O[14] ,
    \Tile_X0Y9_FrameData_O[13] ,
    \Tile_X0Y9_FrameData_O[12] ,
    \Tile_X0Y9_FrameData_O[11] ,
    \Tile_X0Y9_FrameData_O[10] ,
    \Tile_X0Y9_FrameData_O[9] ,
    \Tile_X0Y9_FrameData_O[8] ,
    \Tile_X0Y9_FrameData_O[7] ,
    \Tile_X0Y9_FrameData_O[6] ,
    \Tile_X0Y9_FrameData_O[5] ,
    \Tile_X0Y9_FrameData_O[4] ,
    \Tile_X0Y9_FrameData_O[3] ,
    \Tile_X0Y9_FrameData_O[2] ,
    \Tile_X0Y9_FrameData_O[1] ,
    \Tile_X0Y9_FrameData_O[0] }),
    .FrameStrobe({FrameStrobe[19],
    FrameStrobe[18],
    FrameStrobe[17],
    FrameStrobe[16],
    FrameStrobe[15],
    FrameStrobe[14],
    FrameStrobe[13],
    FrameStrobe[12],
    FrameStrobe[11],
    FrameStrobe[10],
    FrameStrobe[9],
    FrameStrobe[8],
    FrameStrobe[7],
    FrameStrobe[6],
    FrameStrobe[5],
    FrameStrobe[4],
    FrameStrobe[3],
    FrameStrobe[2],
    FrameStrobe[1],
    FrameStrobe[0]}),
    .FrameStrobe_O({\Tile_X0Y9_FrameStrobe_O[19] ,
    \Tile_X0Y9_FrameStrobe_O[18] ,
    \Tile_X0Y9_FrameStrobe_O[17] ,
    \Tile_X0Y9_FrameStrobe_O[16] ,
    \Tile_X0Y9_FrameStrobe_O[15] ,
    \Tile_X0Y9_FrameStrobe_O[14] ,
    \Tile_X0Y9_FrameStrobe_O[13] ,
    \Tile_X0Y9_FrameStrobe_O[12] ,
    \Tile_X0Y9_FrameStrobe_O[11] ,
    \Tile_X0Y9_FrameStrobe_O[10] ,
    \Tile_X0Y9_FrameStrobe_O[9] ,
    \Tile_X0Y9_FrameStrobe_O[8] ,
    \Tile_X0Y9_FrameStrobe_O[7] ,
    \Tile_X0Y9_FrameStrobe_O[6] ,
    \Tile_X0Y9_FrameStrobe_O[5] ,
    \Tile_X0Y9_FrameStrobe_O[4] ,
    \Tile_X0Y9_FrameStrobe_O[3] ,
    \Tile_X0Y9_FrameStrobe_O[2] ,
    \Tile_X0Y9_FrameStrobe_O[1] ,
    \Tile_X0Y9_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X0Y9_N1BEG[3] ,
    \Tile_X0Y9_N1BEG[2] ,
    \Tile_X0Y9_N1BEG[1] ,
    \Tile_X0Y9_N1BEG[0] }),
    .N2BEG({\Tile_X0Y9_N2BEG[7] ,
    \Tile_X0Y9_N2BEG[6] ,
    \Tile_X0Y9_N2BEG[5] ,
    \Tile_X0Y9_N2BEG[4] ,
    \Tile_X0Y9_N2BEG[3] ,
    \Tile_X0Y9_N2BEG[2] ,
    \Tile_X0Y9_N2BEG[1] ,
    \Tile_X0Y9_N2BEG[0] }),
    .N2BEGb({\Tile_X0Y9_N2BEGb[7] ,
    \Tile_X0Y9_N2BEGb[6] ,
    \Tile_X0Y9_N2BEGb[5] ,
    \Tile_X0Y9_N2BEGb[4] ,
    \Tile_X0Y9_N2BEGb[3] ,
    \Tile_X0Y9_N2BEGb[2] ,
    \Tile_X0Y9_N2BEGb[1] ,
    \Tile_X0Y9_N2BEGb[0] }),
    .N4BEG({\Tile_X0Y9_N4BEG[15] ,
    \Tile_X0Y9_N4BEG[14] ,
    \Tile_X0Y9_N4BEG[13] ,
    \Tile_X0Y9_N4BEG[12] ,
    \Tile_X0Y9_N4BEG[11] ,
    \Tile_X0Y9_N4BEG[10] ,
    \Tile_X0Y9_N4BEG[9] ,
    \Tile_X0Y9_N4BEG[8] ,
    \Tile_X0Y9_N4BEG[7] ,
    \Tile_X0Y9_N4BEG[6] ,
    \Tile_X0Y9_N4BEG[5] ,
    \Tile_X0Y9_N4BEG[4] ,
    \Tile_X0Y9_N4BEG[3] ,
    \Tile_X0Y9_N4BEG[2] ,
    \Tile_X0Y9_N4BEG[1] ,
    \Tile_X0Y9_N4BEG[0] }),
    .S1END({\Tile_X0Y8_S1BEG[3] ,
    \Tile_X0Y8_S1BEG[2] ,
    \Tile_X0Y8_S1BEG[1] ,
    \Tile_X0Y8_S1BEG[0] }),
    .S2END({\Tile_X0Y8_S2BEGb[7] ,
    \Tile_X0Y8_S2BEGb[6] ,
    \Tile_X0Y8_S2BEGb[5] ,
    \Tile_X0Y8_S2BEGb[4] ,
    \Tile_X0Y8_S2BEGb[3] ,
    \Tile_X0Y8_S2BEGb[2] ,
    \Tile_X0Y8_S2BEGb[1] ,
    \Tile_X0Y8_S2BEGb[0] }),
    .S2MID({\Tile_X0Y8_S2BEG[7] ,
    \Tile_X0Y8_S2BEG[6] ,
    \Tile_X0Y8_S2BEG[5] ,
    \Tile_X0Y8_S2BEG[4] ,
    \Tile_X0Y8_S2BEG[3] ,
    \Tile_X0Y8_S2BEG[2] ,
    \Tile_X0Y8_S2BEG[1] ,
    \Tile_X0Y8_S2BEG[0] }),
    .S4END({\Tile_X0Y8_S4BEG[15] ,
    \Tile_X0Y8_S4BEG[14] ,
    \Tile_X0Y8_S4BEG[13] ,
    \Tile_X0Y8_S4BEG[12] ,
    \Tile_X0Y8_S4BEG[11] ,
    \Tile_X0Y8_S4BEG[10] ,
    \Tile_X0Y8_S4BEG[9] ,
    \Tile_X0Y8_S4BEG[8] ,
    \Tile_X0Y8_S4BEG[7] ,
    \Tile_X0Y8_S4BEG[6] ,
    \Tile_X0Y8_S4BEG[5] ,
    \Tile_X0Y8_S4BEG[4] ,
    \Tile_X0Y8_S4BEG[3] ,
    \Tile_X0Y8_S4BEG[2] ,
    \Tile_X0Y8_S4BEG[1] ,
    \Tile_X0Y8_S4BEG[0] }));
 N_IO4 Tile_X1Y0_N_IO4 (.A_I_top(Tile_X1Y0_A_I_top),
    .A_O_top(Tile_X1Y0_A_O_top),
    .A_T_top(Tile_X1Y0_A_T_top),
    .B_I_top(Tile_X1Y0_B_I_top),
    .B_O_top(Tile_X1Y0_B_O_top),
    .B_T_top(Tile_X1Y0_B_T_top),
    .C_I_top(Tile_X1Y0_C_I_top),
    .C_O_top(Tile_X1Y0_C_O_top),
    .C_T_top(Tile_X1Y0_C_T_top),
    .Ci(Tile_X1Y1_Co),
    .D_I_top(Tile_X1Y0_D_I_top),
    .D_O_top(Tile_X1Y0_D_O_top),
    .D_T_top(Tile_X1Y0_D_T_top),
    .UserCLK(Tile_X1Y1_UserCLKo),
    .UserCLKo(Tile_X1Y0_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .FrameData({\Tile_X0Y0_FrameData_O[31] ,
    \Tile_X0Y0_FrameData_O[30] ,
    \Tile_X0Y0_FrameData_O[29] ,
    \Tile_X0Y0_FrameData_O[28] ,
    \Tile_X0Y0_FrameData_O[27] ,
    \Tile_X0Y0_FrameData_O[26] ,
    \Tile_X0Y0_FrameData_O[25] ,
    \Tile_X0Y0_FrameData_O[24] ,
    \Tile_X0Y0_FrameData_O[23] ,
    \Tile_X0Y0_FrameData_O[22] ,
    \Tile_X0Y0_FrameData_O[21] ,
    \Tile_X0Y0_FrameData_O[20] ,
    \Tile_X0Y0_FrameData_O[19] ,
    \Tile_X0Y0_FrameData_O[18] ,
    \Tile_X0Y0_FrameData_O[17] ,
    \Tile_X0Y0_FrameData_O[16] ,
    \Tile_X0Y0_FrameData_O[15] ,
    \Tile_X0Y0_FrameData_O[14] ,
    \Tile_X0Y0_FrameData_O[13] ,
    \Tile_X0Y0_FrameData_O[12] ,
    \Tile_X0Y0_FrameData_O[11] ,
    \Tile_X0Y0_FrameData_O[10] ,
    \Tile_X0Y0_FrameData_O[9] ,
    \Tile_X0Y0_FrameData_O[8] ,
    \Tile_X0Y0_FrameData_O[7] ,
    \Tile_X0Y0_FrameData_O[6] ,
    \Tile_X0Y0_FrameData_O[5] ,
    \Tile_X0Y0_FrameData_O[4] ,
    \Tile_X0Y0_FrameData_O[3] ,
    \Tile_X0Y0_FrameData_O[2] ,
    \Tile_X0Y0_FrameData_O[1] ,
    \Tile_X0Y0_FrameData_O[0] }),
    .FrameData_O({\Tile_X1Y0_FrameData_O[31] ,
    \Tile_X1Y0_FrameData_O[30] ,
    \Tile_X1Y0_FrameData_O[29] ,
    \Tile_X1Y0_FrameData_O[28] ,
    \Tile_X1Y0_FrameData_O[27] ,
    \Tile_X1Y0_FrameData_O[26] ,
    \Tile_X1Y0_FrameData_O[25] ,
    \Tile_X1Y0_FrameData_O[24] ,
    \Tile_X1Y0_FrameData_O[23] ,
    \Tile_X1Y0_FrameData_O[22] ,
    \Tile_X1Y0_FrameData_O[21] ,
    \Tile_X1Y0_FrameData_O[20] ,
    \Tile_X1Y0_FrameData_O[19] ,
    \Tile_X1Y0_FrameData_O[18] ,
    \Tile_X1Y0_FrameData_O[17] ,
    \Tile_X1Y0_FrameData_O[16] ,
    \Tile_X1Y0_FrameData_O[15] ,
    \Tile_X1Y0_FrameData_O[14] ,
    \Tile_X1Y0_FrameData_O[13] ,
    \Tile_X1Y0_FrameData_O[12] ,
    \Tile_X1Y0_FrameData_O[11] ,
    \Tile_X1Y0_FrameData_O[10] ,
    \Tile_X1Y0_FrameData_O[9] ,
    \Tile_X1Y0_FrameData_O[8] ,
    \Tile_X1Y0_FrameData_O[7] ,
    \Tile_X1Y0_FrameData_O[6] ,
    \Tile_X1Y0_FrameData_O[5] ,
    \Tile_X1Y0_FrameData_O[4] ,
    \Tile_X1Y0_FrameData_O[3] ,
    \Tile_X1Y0_FrameData_O[2] ,
    \Tile_X1Y0_FrameData_O[1] ,
    \Tile_X1Y0_FrameData_O[0] }),
    .FrameStrobe({\Tile_X1Y1_FrameStrobe_O[19] ,
    \Tile_X1Y1_FrameStrobe_O[18] ,
    \Tile_X1Y1_FrameStrobe_O[17] ,
    \Tile_X1Y1_FrameStrobe_O[16] ,
    \Tile_X1Y1_FrameStrobe_O[15] ,
    \Tile_X1Y1_FrameStrobe_O[14] ,
    \Tile_X1Y1_FrameStrobe_O[13] ,
    \Tile_X1Y1_FrameStrobe_O[12] ,
    \Tile_X1Y1_FrameStrobe_O[11] ,
    \Tile_X1Y1_FrameStrobe_O[10] ,
    \Tile_X1Y1_FrameStrobe_O[9] ,
    \Tile_X1Y1_FrameStrobe_O[8] ,
    \Tile_X1Y1_FrameStrobe_O[7] ,
    \Tile_X1Y1_FrameStrobe_O[6] ,
    \Tile_X1Y1_FrameStrobe_O[5] ,
    \Tile_X1Y1_FrameStrobe_O[4] ,
    \Tile_X1Y1_FrameStrobe_O[3] ,
    \Tile_X1Y1_FrameStrobe_O[2] ,
    \Tile_X1Y1_FrameStrobe_O[1] ,
    \Tile_X1Y1_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X1Y0_FrameStrobe_O[19] ,
    \Tile_X1Y0_FrameStrobe_O[18] ,
    \Tile_X1Y0_FrameStrobe_O[17] ,
    \Tile_X1Y0_FrameStrobe_O[16] ,
    \Tile_X1Y0_FrameStrobe_O[15] ,
    \Tile_X1Y0_FrameStrobe_O[14] ,
    \Tile_X1Y0_FrameStrobe_O[13] ,
    \Tile_X1Y0_FrameStrobe_O[12] ,
    \Tile_X1Y0_FrameStrobe_O[11] ,
    \Tile_X1Y0_FrameStrobe_O[10] ,
    \Tile_X1Y0_FrameStrobe_O[9] ,
    \Tile_X1Y0_FrameStrobe_O[8] ,
    \Tile_X1Y0_FrameStrobe_O[7] ,
    \Tile_X1Y0_FrameStrobe_O[6] ,
    \Tile_X1Y0_FrameStrobe_O[5] ,
    \Tile_X1Y0_FrameStrobe_O[4] ,
    \Tile_X1Y0_FrameStrobe_O[3] ,
    \Tile_X1Y0_FrameStrobe_O[2] ,
    \Tile_X1Y0_FrameStrobe_O[1] ,
    \Tile_X1Y0_FrameStrobe_O[0] }),
    .N1END({\Tile_X1Y1_N1BEG[3] ,
    \Tile_X1Y1_N1BEG[2] ,
    \Tile_X1Y1_N1BEG[1] ,
    \Tile_X1Y1_N1BEG[0] }),
    .N2END({\Tile_X1Y1_N2BEGb[7] ,
    \Tile_X1Y1_N2BEGb[6] ,
    \Tile_X1Y1_N2BEGb[5] ,
    \Tile_X1Y1_N2BEGb[4] ,
    \Tile_X1Y1_N2BEGb[3] ,
    \Tile_X1Y1_N2BEGb[2] ,
    \Tile_X1Y1_N2BEGb[1] ,
    \Tile_X1Y1_N2BEGb[0] }),
    .N2MID({\Tile_X1Y1_N2BEG[7] ,
    \Tile_X1Y1_N2BEG[6] ,
    \Tile_X1Y1_N2BEG[5] ,
    \Tile_X1Y1_N2BEG[4] ,
    \Tile_X1Y1_N2BEG[3] ,
    \Tile_X1Y1_N2BEG[2] ,
    \Tile_X1Y1_N2BEG[1] ,
    \Tile_X1Y1_N2BEG[0] }),
    .N4END({\Tile_X1Y1_N4BEG[15] ,
    \Tile_X1Y1_N4BEG[14] ,
    \Tile_X1Y1_N4BEG[13] ,
    \Tile_X1Y1_N4BEG[12] ,
    \Tile_X1Y1_N4BEG[11] ,
    \Tile_X1Y1_N4BEG[10] ,
    \Tile_X1Y1_N4BEG[9] ,
    \Tile_X1Y1_N4BEG[8] ,
    \Tile_X1Y1_N4BEG[7] ,
    \Tile_X1Y1_N4BEG[6] ,
    \Tile_X1Y1_N4BEG[5] ,
    \Tile_X1Y1_N4BEG[4] ,
    \Tile_X1Y1_N4BEG[3] ,
    \Tile_X1Y1_N4BEG[2] ,
    \Tile_X1Y1_N4BEG[1] ,
    \Tile_X1Y1_N4BEG[0] }),
    .NN4END({\Tile_X1Y1_NN4BEG[15] ,
    \Tile_X1Y1_NN4BEG[14] ,
    \Tile_X1Y1_NN4BEG[13] ,
    \Tile_X1Y1_NN4BEG[12] ,
    \Tile_X1Y1_NN4BEG[11] ,
    \Tile_X1Y1_NN4BEG[10] ,
    \Tile_X1Y1_NN4BEG[9] ,
    \Tile_X1Y1_NN4BEG[8] ,
    \Tile_X1Y1_NN4BEG[7] ,
    \Tile_X1Y1_NN4BEG[6] ,
    \Tile_X1Y1_NN4BEG[5] ,
    \Tile_X1Y1_NN4BEG[4] ,
    \Tile_X1Y1_NN4BEG[3] ,
    \Tile_X1Y1_NN4BEG[2] ,
    \Tile_X1Y1_NN4BEG[1] ,
    \Tile_X1Y1_NN4BEG[0] }),
    .S1BEG({\Tile_X1Y0_S1BEG[3] ,
    \Tile_X1Y0_S1BEG[2] ,
    \Tile_X1Y0_S1BEG[1] ,
    \Tile_X1Y0_S1BEG[0] }),
    .S2BEG({\Tile_X1Y0_S2BEG[7] ,
    \Tile_X1Y0_S2BEG[6] ,
    \Tile_X1Y0_S2BEG[5] ,
    \Tile_X1Y0_S2BEG[4] ,
    \Tile_X1Y0_S2BEG[3] ,
    \Tile_X1Y0_S2BEG[2] ,
    \Tile_X1Y0_S2BEG[1] ,
    \Tile_X1Y0_S2BEG[0] }),
    .S2BEGb({\Tile_X1Y0_S2BEGb[7] ,
    \Tile_X1Y0_S2BEGb[6] ,
    \Tile_X1Y0_S2BEGb[5] ,
    \Tile_X1Y0_S2BEGb[4] ,
    \Tile_X1Y0_S2BEGb[3] ,
    \Tile_X1Y0_S2BEGb[2] ,
    \Tile_X1Y0_S2BEGb[1] ,
    \Tile_X1Y0_S2BEGb[0] }),
    .S4BEG({\Tile_X1Y0_S4BEG[15] ,
    \Tile_X1Y0_S4BEG[14] ,
    \Tile_X1Y0_S4BEG[13] ,
    \Tile_X1Y0_S4BEG[12] ,
    \Tile_X1Y0_S4BEG[11] ,
    \Tile_X1Y0_S4BEG[10] ,
    \Tile_X1Y0_S4BEG[9] ,
    \Tile_X1Y0_S4BEG[8] ,
    \Tile_X1Y0_S4BEG[7] ,
    \Tile_X1Y0_S4BEG[6] ,
    \Tile_X1Y0_S4BEG[5] ,
    \Tile_X1Y0_S4BEG[4] ,
    \Tile_X1Y0_S4BEG[3] ,
    \Tile_X1Y0_S4BEG[2] ,
    \Tile_X1Y0_S4BEG[1] ,
    \Tile_X1Y0_S4BEG[0] }),
    .SS4BEG({\Tile_X1Y0_SS4BEG[15] ,
    \Tile_X1Y0_SS4BEG[14] ,
    \Tile_X1Y0_SS4BEG[13] ,
    \Tile_X1Y0_SS4BEG[12] ,
    \Tile_X1Y0_SS4BEG[11] ,
    \Tile_X1Y0_SS4BEG[10] ,
    \Tile_X1Y0_SS4BEG[9] ,
    \Tile_X1Y0_SS4BEG[8] ,
    \Tile_X1Y0_SS4BEG[7] ,
    \Tile_X1Y0_SS4BEG[6] ,
    \Tile_X1Y0_SS4BEG[5] ,
    \Tile_X1Y0_SS4BEG[4] ,
    \Tile_X1Y0_SS4BEG[3] ,
    \Tile_X1Y0_SS4BEG[2] ,
    \Tile_X1Y0_SS4BEG[1] ,
    \Tile_X1Y0_SS4BEG[0] }));
 LUT4AB Tile_X1Y1_LUT4AB (.Ci(Tile_X1Y2_Co),
    .Co(Tile_X1Y1_Co),
    .UserCLK(Tile_X1Y2_UserCLKo),
    .UserCLKo(Tile_X1Y1_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X1Y1_E1BEG[3] ,
    \Tile_X1Y1_E1BEG[2] ,
    \Tile_X1Y1_E1BEG[1] ,
    \Tile_X1Y1_E1BEG[0] }),
    .E1END({\Tile_X0Y1_E1BEG[3] ,
    \Tile_X0Y1_E1BEG[2] ,
    \Tile_X0Y1_E1BEG[1] ,
    \Tile_X0Y1_E1BEG[0] }),
    .E2BEG({\Tile_X1Y1_E2BEG[7] ,
    \Tile_X1Y1_E2BEG[6] ,
    \Tile_X1Y1_E2BEG[5] ,
    \Tile_X1Y1_E2BEG[4] ,
    \Tile_X1Y1_E2BEG[3] ,
    \Tile_X1Y1_E2BEG[2] ,
    \Tile_X1Y1_E2BEG[1] ,
    \Tile_X1Y1_E2BEG[0] }),
    .E2BEGb({\Tile_X1Y1_E2BEGb[7] ,
    \Tile_X1Y1_E2BEGb[6] ,
    \Tile_X1Y1_E2BEGb[5] ,
    \Tile_X1Y1_E2BEGb[4] ,
    \Tile_X1Y1_E2BEGb[3] ,
    \Tile_X1Y1_E2BEGb[2] ,
    \Tile_X1Y1_E2BEGb[1] ,
    \Tile_X1Y1_E2BEGb[0] }),
    .E2END({\Tile_X0Y1_E2BEGb[7] ,
    \Tile_X0Y1_E2BEGb[6] ,
    \Tile_X0Y1_E2BEGb[5] ,
    \Tile_X0Y1_E2BEGb[4] ,
    \Tile_X0Y1_E2BEGb[3] ,
    \Tile_X0Y1_E2BEGb[2] ,
    \Tile_X0Y1_E2BEGb[1] ,
    \Tile_X0Y1_E2BEGb[0] }),
    .E2MID({\Tile_X0Y1_E2BEG[7] ,
    \Tile_X0Y1_E2BEG[6] ,
    \Tile_X0Y1_E2BEG[5] ,
    \Tile_X0Y1_E2BEG[4] ,
    \Tile_X0Y1_E2BEG[3] ,
    \Tile_X0Y1_E2BEG[2] ,
    \Tile_X0Y1_E2BEG[1] ,
    \Tile_X0Y1_E2BEG[0] }),
    .E6BEG({\Tile_X1Y1_E6BEG[11] ,
    \Tile_X1Y1_E6BEG[10] ,
    \Tile_X1Y1_E6BEG[9] ,
    \Tile_X1Y1_E6BEG[8] ,
    \Tile_X1Y1_E6BEG[7] ,
    \Tile_X1Y1_E6BEG[6] ,
    \Tile_X1Y1_E6BEG[5] ,
    \Tile_X1Y1_E6BEG[4] ,
    \Tile_X1Y1_E6BEG[3] ,
    \Tile_X1Y1_E6BEG[2] ,
    \Tile_X1Y1_E6BEG[1] ,
    \Tile_X1Y1_E6BEG[0] }),
    .E6END({\Tile_X0Y1_E6BEG[11] ,
    \Tile_X0Y1_E6BEG[10] ,
    \Tile_X0Y1_E6BEG[9] ,
    \Tile_X0Y1_E6BEG[8] ,
    \Tile_X0Y1_E6BEG[7] ,
    \Tile_X0Y1_E6BEG[6] ,
    \Tile_X0Y1_E6BEG[5] ,
    \Tile_X0Y1_E6BEG[4] ,
    \Tile_X0Y1_E6BEG[3] ,
    \Tile_X0Y1_E6BEG[2] ,
    \Tile_X0Y1_E6BEG[1] ,
    \Tile_X0Y1_E6BEG[0] }),
    .EE4BEG({\Tile_X1Y1_EE4BEG[15] ,
    \Tile_X1Y1_EE4BEG[14] ,
    \Tile_X1Y1_EE4BEG[13] ,
    \Tile_X1Y1_EE4BEG[12] ,
    \Tile_X1Y1_EE4BEG[11] ,
    \Tile_X1Y1_EE4BEG[10] ,
    \Tile_X1Y1_EE4BEG[9] ,
    \Tile_X1Y1_EE4BEG[8] ,
    \Tile_X1Y1_EE4BEG[7] ,
    \Tile_X1Y1_EE4BEG[6] ,
    \Tile_X1Y1_EE4BEG[5] ,
    \Tile_X1Y1_EE4BEG[4] ,
    \Tile_X1Y1_EE4BEG[3] ,
    \Tile_X1Y1_EE4BEG[2] ,
    \Tile_X1Y1_EE4BEG[1] ,
    \Tile_X1Y1_EE4BEG[0] }),
    .EE4END({\Tile_X0Y1_EE4BEG[15] ,
    \Tile_X0Y1_EE4BEG[14] ,
    \Tile_X0Y1_EE4BEG[13] ,
    \Tile_X0Y1_EE4BEG[12] ,
    \Tile_X0Y1_EE4BEG[11] ,
    \Tile_X0Y1_EE4BEG[10] ,
    \Tile_X0Y1_EE4BEG[9] ,
    \Tile_X0Y1_EE4BEG[8] ,
    \Tile_X0Y1_EE4BEG[7] ,
    \Tile_X0Y1_EE4BEG[6] ,
    \Tile_X0Y1_EE4BEG[5] ,
    \Tile_X0Y1_EE4BEG[4] ,
    \Tile_X0Y1_EE4BEG[3] ,
    \Tile_X0Y1_EE4BEG[2] ,
    \Tile_X0Y1_EE4BEG[1] ,
    \Tile_X0Y1_EE4BEG[0] }),
    .FrameData({\Tile_X0Y1_FrameData_O[31] ,
    \Tile_X0Y1_FrameData_O[30] ,
    \Tile_X0Y1_FrameData_O[29] ,
    \Tile_X0Y1_FrameData_O[28] ,
    \Tile_X0Y1_FrameData_O[27] ,
    \Tile_X0Y1_FrameData_O[26] ,
    \Tile_X0Y1_FrameData_O[25] ,
    \Tile_X0Y1_FrameData_O[24] ,
    \Tile_X0Y1_FrameData_O[23] ,
    \Tile_X0Y1_FrameData_O[22] ,
    \Tile_X0Y1_FrameData_O[21] ,
    \Tile_X0Y1_FrameData_O[20] ,
    \Tile_X0Y1_FrameData_O[19] ,
    \Tile_X0Y1_FrameData_O[18] ,
    \Tile_X0Y1_FrameData_O[17] ,
    \Tile_X0Y1_FrameData_O[16] ,
    \Tile_X0Y1_FrameData_O[15] ,
    \Tile_X0Y1_FrameData_O[14] ,
    \Tile_X0Y1_FrameData_O[13] ,
    \Tile_X0Y1_FrameData_O[12] ,
    \Tile_X0Y1_FrameData_O[11] ,
    \Tile_X0Y1_FrameData_O[10] ,
    \Tile_X0Y1_FrameData_O[9] ,
    \Tile_X0Y1_FrameData_O[8] ,
    \Tile_X0Y1_FrameData_O[7] ,
    \Tile_X0Y1_FrameData_O[6] ,
    \Tile_X0Y1_FrameData_O[5] ,
    \Tile_X0Y1_FrameData_O[4] ,
    \Tile_X0Y1_FrameData_O[3] ,
    \Tile_X0Y1_FrameData_O[2] ,
    \Tile_X0Y1_FrameData_O[1] ,
    \Tile_X0Y1_FrameData_O[0] }),
    .FrameData_O({\Tile_X1Y1_FrameData_O[31] ,
    \Tile_X1Y1_FrameData_O[30] ,
    \Tile_X1Y1_FrameData_O[29] ,
    \Tile_X1Y1_FrameData_O[28] ,
    \Tile_X1Y1_FrameData_O[27] ,
    \Tile_X1Y1_FrameData_O[26] ,
    \Tile_X1Y1_FrameData_O[25] ,
    \Tile_X1Y1_FrameData_O[24] ,
    \Tile_X1Y1_FrameData_O[23] ,
    \Tile_X1Y1_FrameData_O[22] ,
    \Tile_X1Y1_FrameData_O[21] ,
    \Tile_X1Y1_FrameData_O[20] ,
    \Tile_X1Y1_FrameData_O[19] ,
    \Tile_X1Y1_FrameData_O[18] ,
    \Tile_X1Y1_FrameData_O[17] ,
    \Tile_X1Y1_FrameData_O[16] ,
    \Tile_X1Y1_FrameData_O[15] ,
    \Tile_X1Y1_FrameData_O[14] ,
    \Tile_X1Y1_FrameData_O[13] ,
    \Tile_X1Y1_FrameData_O[12] ,
    \Tile_X1Y1_FrameData_O[11] ,
    \Tile_X1Y1_FrameData_O[10] ,
    \Tile_X1Y1_FrameData_O[9] ,
    \Tile_X1Y1_FrameData_O[8] ,
    \Tile_X1Y1_FrameData_O[7] ,
    \Tile_X1Y1_FrameData_O[6] ,
    \Tile_X1Y1_FrameData_O[5] ,
    \Tile_X1Y1_FrameData_O[4] ,
    \Tile_X1Y1_FrameData_O[3] ,
    \Tile_X1Y1_FrameData_O[2] ,
    \Tile_X1Y1_FrameData_O[1] ,
    \Tile_X1Y1_FrameData_O[0] }),
    .FrameStrobe({\Tile_X1Y2_FrameStrobe_O[19] ,
    \Tile_X1Y2_FrameStrobe_O[18] ,
    \Tile_X1Y2_FrameStrobe_O[17] ,
    \Tile_X1Y2_FrameStrobe_O[16] ,
    \Tile_X1Y2_FrameStrobe_O[15] ,
    \Tile_X1Y2_FrameStrobe_O[14] ,
    \Tile_X1Y2_FrameStrobe_O[13] ,
    \Tile_X1Y2_FrameStrobe_O[12] ,
    \Tile_X1Y2_FrameStrobe_O[11] ,
    \Tile_X1Y2_FrameStrobe_O[10] ,
    \Tile_X1Y2_FrameStrobe_O[9] ,
    \Tile_X1Y2_FrameStrobe_O[8] ,
    \Tile_X1Y2_FrameStrobe_O[7] ,
    \Tile_X1Y2_FrameStrobe_O[6] ,
    \Tile_X1Y2_FrameStrobe_O[5] ,
    \Tile_X1Y2_FrameStrobe_O[4] ,
    \Tile_X1Y2_FrameStrobe_O[3] ,
    \Tile_X1Y2_FrameStrobe_O[2] ,
    \Tile_X1Y2_FrameStrobe_O[1] ,
    \Tile_X1Y2_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X1Y1_FrameStrobe_O[19] ,
    \Tile_X1Y1_FrameStrobe_O[18] ,
    \Tile_X1Y1_FrameStrobe_O[17] ,
    \Tile_X1Y1_FrameStrobe_O[16] ,
    \Tile_X1Y1_FrameStrobe_O[15] ,
    \Tile_X1Y1_FrameStrobe_O[14] ,
    \Tile_X1Y1_FrameStrobe_O[13] ,
    \Tile_X1Y1_FrameStrobe_O[12] ,
    \Tile_X1Y1_FrameStrobe_O[11] ,
    \Tile_X1Y1_FrameStrobe_O[10] ,
    \Tile_X1Y1_FrameStrobe_O[9] ,
    \Tile_X1Y1_FrameStrobe_O[8] ,
    \Tile_X1Y1_FrameStrobe_O[7] ,
    \Tile_X1Y1_FrameStrobe_O[6] ,
    \Tile_X1Y1_FrameStrobe_O[5] ,
    \Tile_X1Y1_FrameStrobe_O[4] ,
    \Tile_X1Y1_FrameStrobe_O[3] ,
    \Tile_X1Y1_FrameStrobe_O[2] ,
    \Tile_X1Y1_FrameStrobe_O[1] ,
    \Tile_X1Y1_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X1Y1_N1BEG[3] ,
    \Tile_X1Y1_N1BEG[2] ,
    \Tile_X1Y1_N1BEG[1] ,
    \Tile_X1Y1_N1BEG[0] }),
    .N1END({\Tile_X1Y2_N1BEG[3] ,
    \Tile_X1Y2_N1BEG[2] ,
    \Tile_X1Y2_N1BEG[1] ,
    \Tile_X1Y2_N1BEG[0] }),
    .N2BEG({\Tile_X1Y1_N2BEG[7] ,
    \Tile_X1Y1_N2BEG[6] ,
    \Tile_X1Y1_N2BEG[5] ,
    \Tile_X1Y1_N2BEG[4] ,
    \Tile_X1Y1_N2BEG[3] ,
    \Tile_X1Y1_N2BEG[2] ,
    \Tile_X1Y1_N2BEG[1] ,
    \Tile_X1Y1_N2BEG[0] }),
    .N2BEGb({\Tile_X1Y1_N2BEGb[7] ,
    \Tile_X1Y1_N2BEGb[6] ,
    \Tile_X1Y1_N2BEGb[5] ,
    \Tile_X1Y1_N2BEGb[4] ,
    \Tile_X1Y1_N2BEGb[3] ,
    \Tile_X1Y1_N2BEGb[2] ,
    \Tile_X1Y1_N2BEGb[1] ,
    \Tile_X1Y1_N2BEGb[0] }),
    .N2END({\Tile_X1Y2_N2BEGb[7] ,
    \Tile_X1Y2_N2BEGb[6] ,
    \Tile_X1Y2_N2BEGb[5] ,
    \Tile_X1Y2_N2BEGb[4] ,
    \Tile_X1Y2_N2BEGb[3] ,
    \Tile_X1Y2_N2BEGb[2] ,
    \Tile_X1Y2_N2BEGb[1] ,
    \Tile_X1Y2_N2BEGb[0] }),
    .N2MID({\Tile_X1Y2_N2BEG[7] ,
    \Tile_X1Y2_N2BEG[6] ,
    \Tile_X1Y2_N2BEG[5] ,
    \Tile_X1Y2_N2BEG[4] ,
    \Tile_X1Y2_N2BEG[3] ,
    \Tile_X1Y2_N2BEG[2] ,
    \Tile_X1Y2_N2BEG[1] ,
    \Tile_X1Y2_N2BEG[0] }),
    .N4BEG({\Tile_X1Y1_N4BEG[15] ,
    \Tile_X1Y1_N4BEG[14] ,
    \Tile_X1Y1_N4BEG[13] ,
    \Tile_X1Y1_N4BEG[12] ,
    \Tile_X1Y1_N4BEG[11] ,
    \Tile_X1Y1_N4BEG[10] ,
    \Tile_X1Y1_N4BEG[9] ,
    \Tile_X1Y1_N4BEG[8] ,
    \Tile_X1Y1_N4BEG[7] ,
    \Tile_X1Y1_N4BEG[6] ,
    \Tile_X1Y1_N4BEG[5] ,
    \Tile_X1Y1_N4BEG[4] ,
    \Tile_X1Y1_N4BEG[3] ,
    \Tile_X1Y1_N4BEG[2] ,
    \Tile_X1Y1_N4BEG[1] ,
    \Tile_X1Y1_N4BEG[0] }),
    .N4END({\Tile_X1Y2_N4BEG[15] ,
    \Tile_X1Y2_N4BEG[14] ,
    \Tile_X1Y2_N4BEG[13] ,
    \Tile_X1Y2_N4BEG[12] ,
    \Tile_X1Y2_N4BEG[11] ,
    \Tile_X1Y2_N4BEG[10] ,
    \Tile_X1Y2_N4BEG[9] ,
    \Tile_X1Y2_N4BEG[8] ,
    \Tile_X1Y2_N4BEG[7] ,
    \Tile_X1Y2_N4BEG[6] ,
    \Tile_X1Y2_N4BEG[5] ,
    \Tile_X1Y2_N4BEG[4] ,
    \Tile_X1Y2_N4BEG[3] ,
    \Tile_X1Y2_N4BEG[2] ,
    \Tile_X1Y2_N4BEG[1] ,
    \Tile_X1Y2_N4BEG[0] }),
    .NN4BEG({\Tile_X1Y1_NN4BEG[15] ,
    \Tile_X1Y1_NN4BEG[14] ,
    \Tile_X1Y1_NN4BEG[13] ,
    \Tile_X1Y1_NN4BEG[12] ,
    \Tile_X1Y1_NN4BEG[11] ,
    \Tile_X1Y1_NN4BEG[10] ,
    \Tile_X1Y1_NN4BEG[9] ,
    \Tile_X1Y1_NN4BEG[8] ,
    \Tile_X1Y1_NN4BEG[7] ,
    \Tile_X1Y1_NN4BEG[6] ,
    \Tile_X1Y1_NN4BEG[5] ,
    \Tile_X1Y1_NN4BEG[4] ,
    \Tile_X1Y1_NN4BEG[3] ,
    \Tile_X1Y1_NN4BEG[2] ,
    \Tile_X1Y1_NN4BEG[1] ,
    \Tile_X1Y1_NN4BEG[0] }),
    .NN4END({\Tile_X1Y2_NN4BEG[15] ,
    \Tile_X1Y2_NN4BEG[14] ,
    \Tile_X1Y2_NN4BEG[13] ,
    \Tile_X1Y2_NN4BEG[12] ,
    \Tile_X1Y2_NN4BEG[11] ,
    \Tile_X1Y2_NN4BEG[10] ,
    \Tile_X1Y2_NN4BEG[9] ,
    \Tile_X1Y2_NN4BEG[8] ,
    \Tile_X1Y2_NN4BEG[7] ,
    \Tile_X1Y2_NN4BEG[6] ,
    \Tile_X1Y2_NN4BEG[5] ,
    \Tile_X1Y2_NN4BEG[4] ,
    \Tile_X1Y2_NN4BEG[3] ,
    \Tile_X1Y2_NN4BEG[2] ,
    \Tile_X1Y2_NN4BEG[1] ,
    \Tile_X1Y2_NN4BEG[0] }),
    .S1BEG({\Tile_X1Y1_S1BEG[3] ,
    \Tile_X1Y1_S1BEG[2] ,
    \Tile_X1Y1_S1BEG[1] ,
    \Tile_X1Y1_S1BEG[0] }),
    .S1END({\Tile_X1Y0_S1BEG[3] ,
    \Tile_X1Y0_S1BEG[2] ,
    \Tile_X1Y0_S1BEG[1] ,
    \Tile_X1Y0_S1BEG[0] }),
    .S2BEG({\Tile_X1Y1_S2BEG[7] ,
    \Tile_X1Y1_S2BEG[6] ,
    \Tile_X1Y1_S2BEG[5] ,
    \Tile_X1Y1_S2BEG[4] ,
    \Tile_X1Y1_S2BEG[3] ,
    \Tile_X1Y1_S2BEG[2] ,
    \Tile_X1Y1_S2BEG[1] ,
    \Tile_X1Y1_S2BEG[0] }),
    .S2BEGb({\Tile_X1Y1_S2BEGb[7] ,
    \Tile_X1Y1_S2BEGb[6] ,
    \Tile_X1Y1_S2BEGb[5] ,
    \Tile_X1Y1_S2BEGb[4] ,
    \Tile_X1Y1_S2BEGb[3] ,
    \Tile_X1Y1_S2BEGb[2] ,
    \Tile_X1Y1_S2BEGb[1] ,
    \Tile_X1Y1_S2BEGb[0] }),
    .S2END({\Tile_X1Y0_S2BEGb[7] ,
    \Tile_X1Y0_S2BEGb[6] ,
    \Tile_X1Y0_S2BEGb[5] ,
    \Tile_X1Y0_S2BEGb[4] ,
    \Tile_X1Y0_S2BEGb[3] ,
    \Tile_X1Y0_S2BEGb[2] ,
    \Tile_X1Y0_S2BEGb[1] ,
    \Tile_X1Y0_S2BEGb[0] }),
    .S2MID({\Tile_X1Y0_S2BEG[7] ,
    \Tile_X1Y0_S2BEG[6] ,
    \Tile_X1Y0_S2BEG[5] ,
    \Tile_X1Y0_S2BEG[4] ,
    \Tile_X1Y0_S2BEG[3] ,
    \Tile_X1Y0_S2BEG[2] ,
    \Tile_X1Y0_S2BEG[1] ,
    \Tile_X1Y0_S2BEG[0] }),
    .S4BEG({\Tile_X1Y1_S4BEG[15] ,
    \Tile_X1Y1_S4BEG[14] ,
    \Tile_X1Y1_S4BEG[13] ,
    \Tile_X1Y1_S4BEG[12] ,
    \Tile_X1Y1_S4BEG[11] ,
    \Tile_X1Y1_S4BEG[10] ,
    \Tile_X1Y1_S4BEG[9] ,
    \Tile_X1Y1_S4BEG[8] ,
    \Tile_X1Y1_S4BEG[7] ,
    \Tile_X1Y1_S4BEG[6] ,
    \Tile_X1Y1_S4BEG[5] ,
    \Tile_X1Y1_S4BEG[4] ,
    \Tile_X1Y1_S4BEG[3] ,
    \Tile_X1Y1_S4BEG[2] ,
    \Tile_X1Y1_S4BEG[1] ,
    \Tile_X1Y1_S4BEG[0] }),
    .S4END({\Tile_X1Y0_S4BEG[15] ,
    \Tile_X1Y0_S4BEG[14] ,
    \Tile_X1Y0_S4BEG[13] ,
    \Tile_X1Y0_S4BEG[12] ,
    \Tile_X1Y0_S4BEG[11] ,
    \Tile_X1Y0_S4BEG[10] ,
    \Tile_X1Y0_S4BEG[9] ,
    \Tile_X1Y0_S4BEG[8] ,
    \Tile_X1Y0_S4BEG[7] ,
    \Tile_X1Y0_S4BEG[6] ,
    \Tile_X1Y0_S4BEG[5] ,
    \Tile_X1Y0_S4BEG[4] ,
    \Tile_X1Y0_S4BEG[3] ,
    \Tile_X1Y0_S4BEG[2] ,
    \Tile_X1Y0_S4BEG[1] ,
    \Tile_X1Y0_S4BEG[0] }),
    .SS4BEG({\Tile_X1Y1_SS4BEG[15] ,
    \Tile_X1Y1_SS4BEG[14] ,
    \Tile_X1Y1_SS4BEG[13] ,
    \Tile_X1Y1_SS4BEG[12] ,
    \Tile_X1Y1_SS4BEG[11] ,
    \Tile_X1Y1_SS4BEG[10] ,
    \Tile_X1Y1_SS4BEG[9] ,
    \Tile_X1Y1_SS4BEG[8] ,
    \Tile_X1Y1_SS4BEG[7] ,
    \Tile_X1Y1_SS4BEG[6] ,
    \Tile_X1Y1_SS4BEG[5] ,
    \Tile_X1Y1_SS4BEG[4] ,
    \Tile_X1Y1_SS4BEG[3] ,
    \Tile_X1Y1_SS4BEG[2] ,
    \Tile_X1Y1_SS4BEG[1] ,
    \Tile_X1Y1_SS4BEG[0] }),
    .SS4END({\Tile_X1Y0_SS4BEG[15] ,
    \Tile_X1Y0_SS4BEG[14] ,
    \Tile_X1Y0_SS4BEG[13] ,
    \Tile_X1Y0_SS4BEG[12] ,
    \Tile_X1Y0_SS4BEG[11] ,
    \Tile_X1Y0_SS4BEG[10] ,
    \Tile_X1Y0_SS4BEG[9] ,
    \Tile_X1Y0_SS4BEG[8] ,
    \Tile_X1Y0_SS4BEG[7] ,
    \Tile_X1Y0_SS4BEG[6] ,
    \Tile_X1Y0_SS4BEG[5] ,
    \Tile_X1Y0_SS4BEG[4] ,
    \Tile_X1Y0_SS4BEG[3] ,
    \Tile_X1Y0_SS4BEG[2] ,
    \Tile_X1Y0_SS4BEG[1] ,
    \Tile_X1Y0_SS4BEG[0] }),
    .W1BEG({\Tile_X1Y1_W1BEG[3] ,
    \Tile_X1Y1_W1BEG[2] ,
    \Tile_X1Y1_W1BEG[1] ,
    \Tile_X1Y1_W1BEG[0] }),
    .W1END({\Tile_X2Y1_W1BEG[3] ,
    \Tile_X2Y1_W1BEG[2] ,
    \Tile_X2Y1_W1BEG[1] ,
    \Tile_X2Y1_W1BEG[0] }),
    .W2BEG({\Tile_X1Y1_W2BEG[7] ,
    \Tile_X1Y1_W2BEG[6] ,
    \Tile_X1Y1_W2BEG[5] ,
    \Tile_X1Y1_W2BEG[4] ,
    \Tile_X1Y1_W2BEG[3] ,
    \Tile_X1Y1_W2BEG[2] ,
    \Tile_X1Y1_W2BEG[1] ,
    \Tile_X1Y1_W2BEG[0] }),
    .W2BEGb({\Tile_X1Y1_W2BEGb[7] ,
    \Tile_X1Y1_W2BEGb[6] ,
    \Tile_X1Y1_W2BEGb[5] ,
    \Tile_X1Y1_W2BEGb[4] ,
    \Tile_X1Y1_W2BEGb[3] ,
    \Tile_X1Y1_W2BEGb[2] ,
    \Tile_X1Y1_W2BEGb[1] ,
    \Tile_X1Y1_W2BEGb[0] }),
    .W2END({\Tile_X2Y1_W2BEGb[7] ,
    \Tile_X2Y1_W2BEGb[6] ,
    \Tile_X2Y1_W2BEGb[5] ,
    \Tile_X2Y1_W2BEGb[4] ,
    \Tile_X2Y1_W2BEGb[3] ,
    \Tile_X2Y1_W2BEGb[2] ,
    \Tile_X2Y1_W2BEGb[1] ,
    \Tile_X2Y1_W2BEGb[0] }),
    .W2MID({\Tile_X2Y1_W2BEG[7] ,
    \Tile_X2Y1_W2BEG[6] ,
    \Tile_X2Y1_W2BEG[5] ,
    \Tile_X2Y1_W2BEG[4] ,
    \Tile_X2Y1_W2BEG[3] ,
    \Tile_X2Y1_W2BEG[2] ,
    \Tile_X2Y1_W2BEG[1] ,
    \Tile_X2Y1_W2BEG[0] }),
    .W6BEG({\Tile_X1Y1_W6BEG[11] ,
    \Tile_X1Y1_W6BEG[10] ,
    \Tile_X1Y1_W6BEG[9] ,
    \Tile_X1Y1_W6BEG[8] ,
    \Tile_X1Y1_W6BEG[7] ,
    \Tile_X1Y1_W6BEG[6] ,
    \Tile_X1Y1_W6BEG[5] ,
    \Tile_X1Y1_W6BEG[4] ,
    \Tile_X1Y1_W6BEG[3] ,
    \Tile_X1Y1_W6BEG[2] ,
    \Tile_X1Y1_W6BEG[1] ,
    \Tile_X1Y1_W6BEG[0] }),
    .W6END({\Tile_X2Y1_W6BEG[11] ,
    \Tile_X2Y1_W6BEG[10] ,
    \Tile_X2Y1_W6BEG[9] ,
    \Tile_X2Y1_W6BEG[8] ,
    \Tile_X2Y1_W6BEG[7] ,
    \Tile_X2Y1_W6BEG[6] ,
    \Tile_X2Y1_W6BEG[5] ,
    \Tile_X2Y1_W6BEG[4] ,
    \Tile_X2Y1_W6BEG[3] ,
    \Tile_X2Y1_W6BEG[2] ,
    \Tile_X2Y1_W6BEG[1] ,
    \Tile_X2Y1_W6BEG[0] }),
    .WW4BEG({\Tile_X1Y1_WW4BEG[15] ,
    \Tile_X1Y1_WW4BEG[14] ,
    \Tile_X1Y1_WW4BEG[13] ,
    \Tile_X1Y1_WW4BEG[12] ,
    \Tile_X1Y1_WW4BEG[11] ,
    \Tile_X1Y1_WW4BEG[10] ,
    \Tile_X1Y1_WW4BEG[9] ,
    \Tile_X1Y1_WW4BEG[8] ,
    \Tile_X1Y1_WW4BEG[7] ,
    \Tile_X1Y1_WW4BEG[6] ,
    \Tile_X1Y1_WW4BEG[5] ,
    \Tile_X1Y1_WW4BEG[4] ,
    \Tile_X1Y1_WW4BEG[3] ,
    \Tile_X1Y1_WW4BEG[2] ,
    \Tile_X1Y1_WW4BEG[1] ,
    \Tile_X1Y1_WW4BEG[0] }),
    .WW4END({\Tile_X2Y1_WW4BEG[15] ,
    \Tile_X2Y1_WW4BEG[14] ,
    \Tile_X2Y1_WW4BEG[13] ,
    \Tile_X2Y1_WW4BEG[12] ,
    \Tile_X2Y1_WW4BEG[11] ,
    \Tile_X2Y1_WW4BEG[10] ,
    \Tile_X2Y1_WW4BEG[9] ,
    \Tile_X2Y1_WW4BEG[8] ,
    \Tile_X2Y1_WW4BEG[7] ,
    \Tile_X2Y1_WW4BEG[6] ,
    \Tile_X2Y1_WW4BEG[5] ,
    \Tile_X2Y1_WW4BEG[4] ,
    \Tile_X2Y1_WW4BEG[3] ,
    \Tile_X2Y1_WW4BEG[2] ,
    \Tile_X2Y1_WW4BEG[1] ,
    \Tile_X2Y1_WW4BEG[0] }));
 LUT4AB Tile_X1Y2_LUT4AB (.Ci(Tile_X1Y3_Co),
    .Co(Tile_X1Y2_Co),
    .UserCLK(Tile_X1Y3_UserCLKo),
    .UserCLKo(Tile_X1Y2_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X1Y2_E1BEG[3] ,
    \Tile_X1Y2_E1BEG[2] ,
    \Tile_X1Y2_E1BEG[1] ,
    \Tile_X1Y2_E1BEG[0] }),
    .E1END({\Tile_X0Y2_E1BEG[3] ,
    \Tile_X0Y2_E1BEG[2] ,
    \Tile_X0Y2_E1BEG[1] ,
    \Tile_X0Y2_E1BEG[0] }),
    .E2BEG({\Tile_X1Y2_E2BEG[7] ,
    \Tile_X1Y2_E2BEG[6] ,
    \Tile_X1Y2_E2BEG[5] ,
    \Tile_X1Y2_E2BEG[4] ,
    \Tile_X1Y2_E2BEG[3] ,
    \Tile_X1Y2_E2BEG[2] ,
    \Tile_X1Y2_E2BEG[1] ,
    \Tile_X1Y2_E2BEG[0] }),
    .E2BEGb({\Tile_X1Y2_E2BEGb[7] ,
    \Tile_X1Y2_E2BEGb[6] ,
    \Tile_X1Y2_E2BEGb[5] ,
    \Tile_X1Y2_E2BEGb[4] ,
    \Tile_X1Y2_E2BEGb[3] ,
    \Tile_X1Y2_E2BEGb[2] ,
    \Tile_X1Y2_E2BEGb[1] ,
    \Tile_X1Y2_E2BEGb[0] }),
    .E2END({\Tile_X0Y2_E2BEGb[7] ,
    \Tile_X0Y2_E2BEGb[6] ,
    \Tile_X0Y2_E2BEGb[5] ,
    \Tile_X0Y2_E2BEGb[4] ,
    \Tile_X0Y2_E2BEGb[3] ,
    \Tile_X0Y2_E2BEGb[2] ,
    \Tile_X0Y2_E2BEGb[1] ,
    \Tile_X0Y2_E2BEGb[0] }),
    .E2MID({\Tile_X0Y2_E2BEG[7] ,
    \Tile_X0Y2_E2BEG[6] ,
    \Tile_X0Y2_E2BEG[5] ,
    \Tile_X0Y2_E2BEG[4] ,
    \Tile_X0Y2_E2BEG[3] ,
    \Tile_X0Y2_E2BEG[2] ,
    \Tile_X0Y2_E2BEG[1] ,
    \Tile_X0Y2_E2BEG[0] }),
    .E6BEG({\Tile_X1Y2_E6BEG[11] ,
    \Tile_X1Y2_E6BEG[10] ,
    \Tile_X1Y2_E6BEG[9] ,
    \Tile_X1Y2_E6BEG[8] ,
    \Tile_X1Y2_E6BEG[7] ,
    \Tile_X1Y2_E6BEG[6] ,
    \Tile_X1Y2_E6BEG[5] ,
    \Tile_X1Y2_E6BEG[4] ,
    \Tile_X1Y2_E6BEG[3] ,
    \Tile_X1Y2_E6BEG[2] ,
    \Tile_X1Y2_E6BEG[1] ,
    \Tile_X1Y2_E6BEG[0] }),
    .E6END({\Tile_X0Y2_E6BEG[11] ,
    \Tile_X0Y2_E6BEG[10] ,
    \Tile_X0Y2_E6BEG[9] ,
    \Tile_X0Y2_E6BEG[8] ,
    \Tile_X0Y2_E6BEG[7] ,
    \Tile_X0Y2_E6BEG[6] ,
    \Tile_X0Y2_E6BEG[5] ,
    \Tile_X0Y2_E6BEG[4] ,
    \Tile_X0Y2_E6BEG[3] ,
    \Tile_X0Y2_E6BEG[2] ,
    \Tile_X0Y2_E6BEG[1] ,
    \Tile_X0Y2_E6BEG[0] }),
    .EE4BEG({\Tile_X1Y2_EE4BEG[15] ,
    \Tile_X1Y2_EE4BEG[14] ,
    \Tile_X1Y2_EE4BEG[13] ,
    \Tile_X1Y2_EE4BEG[12] ,
    \Tile_X1Y2_EE4BEG[11] ,
    \Tile_X1Y2_EE4BEG[10] ,
    \Tile_X1Y2_EE4BEG[9] ,
    \Tile_X1Y2_EE4BEG[8] ,
    \Tile_X1Y2_EE4BEG[7] ,
    \Tile_X1Y2_EE4BEG[6] ,
    \Tile_X1Y2_EE4BEG[5] ,
    \Tile_X1Y2_EE4BEG[4] ,
    \Tile_X1Y2_EE4BEG[3] ,
    \Tile_X1Y2_EE4BEG[2] ,
    \Tile_X1Y2_EE4BEG[1] ,
    \Tile_X1Y2_EE4BEG[0] }),
    .EE4END({\Tile_X0Y2_EE4BEG[15] ,
    \Tile_X0Y2_EE4BEG[14] ,
    \Tile_X0Y2_EE4BEG[13] ,
    \Tile_X0Y2_EE4BEG[12] ,
    \Tile_X0Y2_EE4BEG[11] ,
    \Tile_X0Y2_EE4BEG[10] ,
    \Tile_X0Y2_EE4BEG[9] ,
    \Tile_X0Y2_EE4BEG[8] ,
    \Tile_X0Y2_EE4BEG[7] ,
    \Tile_X0Y2_EE4BEG[6] ,
    \Tile_X0Y2_EE4BEG[5] ,
    \Tile_X0Y2_EE4BEG[4] ,
    \Tile_X0Y2_EE4BEG[3] ,
    \Tile_X0Y2_EE4BEG[2] ,
    \Tile_X0Y2_EE4BEG[1] ,
    \Tile_X0Y2_EE4BEG[0] }),
    .FrameData({\Tile_X0Y2_FrameData_O[31] ,
    \Tile_X0Y2_FrameData_O[30] ,
    \Tile_X0Y2_FrameData_O[29] ,
    \Tile_X0Y2_FrameData_O[28] ,
    \Tile_X0Y2_FrameData_O[27] ,
    \Tile_X0Y2_FrameData_O[26] ,
    \Tile_X0Y2_FrameData_O[25] ,
    \Tile_X0Y2_FrameData_O[24] ,
    \Tile_X0Y2_FrameData_O[23] ,
    \Tile_X0Y2_FrameData_O[22] ,
    \Tile_X0Y2_FrameData_O[21] ,
    \Tile_X0Y2_FrameData_O[20] ,
    \Tile_X0Y2_FrameData_O[19] ,
    \Tile_X0Y2_FrameData_O[18] ,
    \Tile_X0Y2_FrameData_O[17] ,
    \Tile_X0Y2_FrameData_O[16] ,
    \Tile_X0Y2_FrameData_O[15] ,
    \Tile_X0Y2_FrameData_O[14] ,
    \Tile_X0Y2_FrameData_O[13] ,
    \Tile_X0Y2_FrameData_O[12] ,
    \Tile_X0Y2_FrameData_O[11] ,
    \Tile_X0Y2_FrameData_O[10] ,
    \Tile_X0Y2_FrameData_O[9] ,
    \Tile_X0Y2_FrameData_O[8] ,
    \Tile_X0Y2_FrameData_O[7] ,
    \Tile_X0Y2_FrameData_O[6] ,
    \Tile_X0Y2_FrameData_O[5] ,
    \Tile_X0Y2_FrameData_O[4] ,
    \Tile_X0Y2_FrameData_O[3] ,
    \Tile_X0Y2_FrameData_O[2] ,
    \Tile_X0Y2_FrameData_O[1] ,
    \Tile_X0Y2_FrameData_O[0] }),
    .FrameData_O({\Tile_X1Y2_FrameData_O[31] ,
    \Tile_X1Y2_FrameData_O[30] ,
    \Tile_X1Y2_FrameData_O[29] ,
    \Tile_X1Y2_FrameData_O[28] ,
    \Tile_X1Y2_FrameData_O[27] ,
    \Tile_X1Y2_FrameData_O[26] ,
    \Tile_X1Y2_FrameData_O[25] ,
    \Tile_X1Y2_FrameData_O[24] ,
    \Tile_X1Y2_FrameData_O[23] ,
    \Tile_X1Y2_FrameData_O[22] ,
    \Tile_X1Y2_FrameData_O[21] ,
    \Tile_X1Y2_FrameData_O[20] ,
    \Tile_X1Y2_FrameData_O[19] ,
    \Tile_X1Y2_FrameData_O[18] ,
    \Tile_X1Y2_FrameData_O[17] ,
    \Tile_X1Y2_FrameData_O[16] ,
    \Tile_X1Y2_FrameData_O[15] ,
    \Tile_X1Y2_FrameData_O[14] ,
    \Tile_X1Y2_FrameData_O[13] ,
    \Tile_X1Y2_FrameData_O[12] ,
    \Tile_X1Y2_FrameData_O[11] ,
    \Tile_X1Y2_FrameData_O[10] ,
    \Tile_X1Y2_FrameData_O[9] ,
    \Tile_X1Y2_FrameData_O[8] ,
    \Tile_X1Y2_FrameData_O[7] ,
    \Tile_X1Y2_FrameData_O[6] ,
    \Tile_X1Y2_FrameData_O[5] ,
    \Tile_X1Y2_FrameData_O[4] ,
    \Tile_X1Y2_FrameData_O[3] ,
    \Tile_X1Y2_FrameData_O[2] ,
    \Tile_X1Y2_FrameData_O[1] ,
    \Tile_X1Y2_FrameData_O[0] }),
    .FrameStrobe({\Tile_X1Y3_FrameStrobe_O[19] ,
    \Tile_X1Y3_FrameStrobe_O[18] ,
    \Tile_X1Y3_FrameStrobe_O[17] ,
    \Tile_X1Y3_FrameStrobe_O[16] ,
    \Tile_X1Y3_FrameStrobe_O[15] ,
    \Tile_X1Y3_FrameStrobe_O[14] ,
    \Tile_X1Y3_FrameStrobe_O[13] ,
    \Tile_X1Y3_FrameStrobe_O[12] ,
    \Tile_X1Y3_FrameStrobe_O[11] ,
    \Tile_X1Y3_FrameStrobe_O[10] ,
    \Tile_X1Y3_FrameStrobe_O[9] ,
    \Tile_X1Y3_FrameStrobe_O[8] ,
    \Tile_X1Y3_FrameStrobe_O[7] ,
    \Tile_X1Y3_FrameStrobe_O[6] ,
    \Tile_X1Y3_FrameStrobe_O[5] ,
    \Tile_X1Y3_FrameStrobe_O[4] ,
    \Tile_X1Y3_FrameStrobe_O[3] ,
    \Tile_X1Y3_FrameStrobe_O[2] ,
    \Tile_X1Y3_FrameStrobe_O[1] ,
    \Tile_X1Y3_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X1Y2_FrameStrobe_O[19] ,
    \Tile_X1Y2_FrameStrobe_O[18] ,
    \Tile_X1Y2_FrameStrobe_O[17] ,
    \Tile_X1Y2_FrameStrobe_O[16] ,
    \Tile_X1Y2_FrameStrobe_O[15] ,
    \Tile_X1Y2_FrameStrobe_O[14] ,
    \Tile_X1Y2_FrameStrobe_O[13] ,
    \Tile_X1Y2_FrameStrobe_O[12] ,
    \Tile_X1Y2_FrameStrobe_O[11] ,
    \Tile_X1Y2_FrameStrobe_O[10] ,
    \Tile_X1Y2_FrameStrobe_O[9] ,
    \Tile_X1Y2_FrameStrobe_O[8] ,
    \Tile_X1Y2_FrameStrobe_O[7] ,
    \Tile_X1Y2_FrameStrobe_O[6] ,
    \Tile_X1Y2_FrameStrobe_O[5] ,
    \Tile_X1Y2_FrameStrobe_O[4] ,
    \Tile_X1Y2_FrameStrobe_O[3] ,
    \Tile_X1Y2_FrameStrobe_O[2] ,
    \Tile_X1Y2_FrameStrobe_O[1] ,
    \Tile_X1Y2_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X1Y2_N1BEG[3] ,
    \Tile_X1Y2_N1BEG[2] ,
    \Tile_X1Y2_N1BEG[1] ,
    \Tile_X1Y2_N1BEG[0] }),
    .N1END({\Tile_X1Y3_N1BEG[3] ,
    \Tile_X1Y3_N1BEG[2] ,
    \Tile_X1Y3_N1BEG[1] ,
    \Tile_X1Y3_N1BEG[0] }),
    .N2BEG({\Tile_X1Y2_N2BEG[7] ,
    \Tile_X1Y2_N2BEG[6] ,
    \Tile_X1Y2_N2BEG[5] ,
    \Tile_X1Y2_N2BEG[4] ,
    \Tile_X1Y2_N2BEG[3] ,
    \Tile_X1Y2_N2BEG[2] ,
    \Tile_X1Y2_N2BEG[1] ,
    \Tile_X1Y2_N2BEG[0] }),
    .N2BEGb({\Tile_X1Y2_N2BEGb[7] ,
    \Tile_X1Y2_N2BEGb[6] ,
    \Tile_X1Y2_N2BEGb[5] ,
    \Tile_X1Y2_N2BEGb[4] ,
    \Tile_X1Y2_N2BEGb[3] ,
    \Tile_X1Y2_N2BEGb[2] ,
    \Tile_X1Y2_N2BEGb[1] ,
    \Tile_X1Y2_N2BEGb[0] }),
    .N2END({\Tile_X1Y3_N2BEGb[7] ,
    \Tile_X1Y3_N2BEGb[6] ,
    \Tile_X1Y3_N2BEGb[5] ,
    \Tile_X1Y3_N2BEGb[4] ,
    \Tile_X1Y3_N2BEGb[3] ,
    \Tile_X1Y3_N2BEGb[2] ,
    \Tile_X1Y3_N2BEGb[1] ,
    \Tile_X1Y3_N2BEGb[0] }),
    .N2MID({\Tile_X1Y3_N2BEG[7] ,
    \Tile_X1Y3_N2BEG[6] ,
    \Tile_X1Y3_N2BEG[5] ,
    \Tile_X1Y3_N2BEG[4] ,
    \Tile_X1Y3_N2BEG[3] ,
    \Tile_X1Y3_N2BEG[2] ,
    \Tile_X1Y3_N2BEG[1] ,
    \Tile_X1Y3_N2BEG[0] }),
    .N4BEG({\Tile_X1Y2_N4BEG[15] ,
    \Tile_X1Y2_N4BEG[14] ,
    \Tile_X1Y2_N4BEG[13] ,
    \Tile_X1Y2_N4BEG[12] ,
    \Tile_X1Y2_N4BEG[11] ,
    \Tile_X1Y2_N4BEG[10] ,
    \Tile_X1Y2_N4BEG[9] ,
    \Tile_X1Y2_N4BEG[8] ,
    \Tile_X1Y2_N4BEG[7] ,
    \Tile_X1Y2_N4BEG[6] ,
    \Tile_X1Y2_N4BEG[5] ,
    \Tile_X1Y2_N4BEG[4] ,
    \Tile_X1Y2_N4BEG[3] ,
    \Tile_X1Y2_N4BEG[2] ,
    \Tile_X1Y2_N4BEG[1] ,
    \Tile_X1Y2_N4BEG[0] }),
    .N4END({\Tile_X1Y3_N4BEG[15] ,
    \Tile_X1Y3_N4BEG[14] ,
    \Tile_X1Y3_N4BEG[13] ,
    \Tile_X1Y3_N4BEG[12] ,
    \Tile_X1Y3_N4BEG[11] ,
    \Tile_X1Y3_N4BEG[10] ,
    \Tile_X1Y3_N4BEG[9] ,
    \Tile_X1Y3_N4BEG[8] ,
    \Tile_X1Y3_N4BEG[7] ,
    \Tile_X1Y3_N4BEG[6] ,
    \Tile_X1Y3_N4BEG[5] ,
    \Tile_X1Y3_N4BEG[4] ,
    \Tile_X1Y3_N4BEG[3] ,
    \Tile_X1Y3_N4BEG[2] ,
    \Tile_X1Y3_N4BEG[1] ,
    \Tile_X1Y3_N4BEG[0] }),
    .NN4BEG({\Tile_X1Y2_NN4BEG[15] ,
    \Tile_X1Y2_NN4BEG[14] ,
    \Tile_X1Y2_NN4BEG[13] ,
    \Tile_X1Y2_NN4BEG[12] ,
    \Tile_X1Y2_NN4BEG[11] ,
    \Tile_X1Y2_NN4BEG[10] ,
    \Tile_X1Y2_NN4BEG[9] ,
    \Tile_X1Y2_NN4BEG[8] ,
    \Tile_X1Y2_NN4BEG[7] ,
    \Tile_X1Y2_NN4BEG[6] ,
    \Tile_X1Y2_NN4BEG[5] ,
    \Tile_X1Y2_NN4BEG[4] ,
    \Tile_X1Y2_NN4BEG[3] ,
    \Tile_X1Y2_NN4BEG[2] ,
    \Tile_X1Y2_NN4BEG[1] ,
    \Tile_X1Y2_NN4BEG[0] }),
    .NN4END({\Tile_X1Y3_NN4BEG[15] ,
    \Tile_X1Y3_NN4BEG[14] ,
    \Tile_X1Y3_NN4BEG[13] ,
    \Tile_X1Y3_NN4BEG[12] ,
    \Tile_X1Y3_NN4BEG[11] ,
    \Tile_X1Y3_NN4BEG[10] ,
    \Tile_X1Y3_NN4BEG[9] ,
    \Tile_X1Y3_NN4BEG[8] ,
    \Tile_X1Y3_NN4BEG[7] ,
    \Tile_X1Y3_NN4BEG[6] ,
    \Tile_X1Y3_NN4BEG[5] ,
    \Tile_X1Y3_NN4BEG[4] ,
    \Tile_X1Y3_NN4BEG[3] ,
    \Tile_X1Y3_NN4BEG[2] ,
    \Tile_X1Y3_NN4BEG[1] ,
    \Tile_X1Y3_NN4BEG[0] }),
    .S1BEG({\Tile_X1Y2_S1BEG[3] ,
    \Tile_X1Y2_S1BEG[2] ,
    \Tile_X1Y2_S1BEG[1] ,
    \Tile_X1Y2_S1BEG[0] }),
    .S1END({\Tile_X1Y1_S1BEG[3] ,
    \Tile_X1Y1_S1BEG[2] ,
    \Tile_X1Y1_S1BEG[1] ,
    \Tile_X1Y1_S1BEG[0] }),
    .S2BEG({\Tile_X1Y2_S2BEG[7] ,
    \Tile_X1Y2_S2BEG[6] ,
    \Tile_X1Y2_S2BEG[5] ,
    \Tile_X1Y2_S2BEG[4] ,
    \Tile_X1Y2_S2BEG[3] ,
    \Tile_X1Y2_S2BEG[2] ,
    \Tile_X1Y2_S2BEG[1] ,
    \Tile_X1Y2_S2BEG[0] }),
    .S2BEGb({\Tile_X1Y2_S2BEGb[7] ,
    \Tile_X1Y2_S2BEGb[6] ,
    \Tile_X1Y2_S2BEGb[5] ,
    \Tile_X1Y2_S2BEGb[4] ,
    \Tile_X1Y2_S2BEGb[3] ,
    \Tile_X1Y2_S2BEGb[2] ,
    \Tile_X1Y2_S2BEGb[1] ,
    \Tile_X1Y2_S2BEGb[0] }),
    .S2END({\Tile_X1Y1_S2BEGb[7] ,
    \Tile_X1Y1_S2BEGb[6] ,
    \Tile_X1Y1_S2BEGb[5] ,
    \Tile_X1Y1_S2BEGb[4] ,
    \Tile_X1Y1_S2BEGb[3] ,
    \Tile_X1Y1_S2BEGb[2] ,
    \Tile_X1Y1_S2BEGb[1] ,
    \Tile_X1Y1_S2BEGb[0] }),
    .S2MID({\Tile_X1Y1_S2BEG[7] ,
    \Tile_X1Y1_S2BEG[6] ,
    \Tile_X1Y1_S2BEG[5] ,
    \Tile_X1Y1_S2BEG[4] ,
    \Tile_X1Y1_S2BEG[3] ,
    \Tile_X1Y1_S2BEG[2] ,
    \Tile_X1Y1_S2BEG[1] ,
    \Tile_X1Y1_S2BEG[0] }),
    .S4BEG({\Tile_X1Y2_S4BEG[15] ,
    \Tile_X1Y2_S4BEG[14] ,
    \Tile_X1Y2_S4BEG[13] ,
    \Tile_X1Y2_S4BEG[12] ,
    \Tile_X1Y2_S4BEG[11] ,
    \Tile_X1Y2_S4BEG[10] ,
    \Tile_X1Y2_S4BEG[9] ,
    \Tile_X1Y2_S4BEG[8] ,
    \Tile_X1Y2_S4BEG[7] ,
    \Tile_X1Y2_S4BEG[6] ,
    \Tile_X1Y2_S4BEG[5] ,
    \Tile_X1Y2_S4BEG[4] ,
    \Tile_X1Y2_S4BEG[3] ,
    \Tile_X1Y2_S4BEG[2] ,
    \Tile_X1Y2_S4BEG[1] ,
    \Tile_X1Y2_S4BEG[0] }),
    .S4END({\Tile_X1Y1_S4BEG[15] ,
    \Tile_X1Y1_S4BEG[14] ,
    \Tile_X1Y1_S4BEG[13] ,
    \Tile_X1Y1_S4BEG[12] ,
    \Tile_X1Y1_S4BEG[11] ,
    \Tile_X1Y1_S4BEG[10] ,
    \Tile_X1Y1_S4BEG[9] ,
    \Tile_X1Y1_S4BEG[8] ,
    \Tile_X1Y1_S4BEG[7] ,
    \Tile_X1Y1_S4BEG[6] ,
    \Tile_X1Y1_S4BEG[5] ,
    \Tile_X1Y1_S4BEG[4] ,
    \Tile_X1Y1_S4BEG[3] ,
    \Tile_X1Y1_S4BEG[2] ,
    \Tile_X1Y1_S4BEG[1] ,
    \Tile_X1Y1_S4BEG[0] }),
    .SS4BEG({\Tile_X1Y2_SS4BEG[15] ,
    \Tile_X1Y2_SS4BEG[14] ,
    \Tile_X1Y2_SS4BEG[13] ,
    \Tile_X1Y2_SS4BEG[12] ,
    \Tile_X1Y2_SS4BEG[11] ,
    \Tile_X1Y2_SS4BEG[10] ,
    \Tile_X1Y2_SS4BEG[9] ,
    \Tile_X1Y2_SS4BEG[8] ,
    \Tile_X1Y2_SS4BEG[7] ,
    \Tile_X1Y2_SS4BEG[6] ,
    \Tile_X1Y2_SS4BEG[5] ,
    \Tile_X1Y2_SS4BEG[4] ,
    \Tile_X1Y2_SS4BEG[3] ,
    \Tile_X1Y2_SS4BEG[2] ,
    \Tile_X1Y2_SS4BEG[1] ,
    \Tile_X1Y2_SS4BEG[0] }),
    .SS4END({\Tile_X1Y1_SS4BEG[15] ,
    \Tile_X1Y1_SS4BEG[14] ,
    \Tile_X1Y1_SS4BEG[13] ,
    \Tile_X1Y1_SS4BEG[12] ,
    \Tile_X1Y1_SS4BEG[11] ,
    \Tile_X1Y1_SS4BEG[10] ,
    \Tile_X1Y1_SS4BEG[9] ,
    \Tile_X1Y1_SS4BEG[8] ,
    \Tile_X1Y1_SS4BEG[7] ,
    \Tile_X1Y1_SS4BEG[6] ,
    \Tile_X1Y1_SS4BEG[5] ,
    \Tile_X1Y1_SS4BEG[4] ,
    \Tile_X1Y1_SS4BEG[3] ,
    \Tile_X1Y1_SS4BEG[2] ,
    \Tile_X1Y1_SS4BEG[1] ,
    \Tile_X1Y1_SS4BEG[0] }),
    .W1BEG({\Tile_X1Y2_W1BEG[3] ,
    \Tile_X1Y2_W1BEG[2] ,
    \Tile_X1Y2_W1BEG[1] ,
    \Tile_X1Y2_W1BEG[0] }),
    .W1END({\Tile_X2Y2_W1BEG[3] ,
    \Tile_X2Y2_W1BEG[2] ,
    \Tile_X2Y2_W1BEG[1] ,
    \Tile_X2Y2_W1BEG[0] }),
    .W2BEG({\Tile_X1Y2_W2BEG[7] ,
    \Tile_X1Y2_W2BEG[6] ,
    \Tile_X1Y2_W2BEG[5] ,
    \Tile_X1Y2_W2BEG[4] ,
    \Tile_X1Y2_W2BEG[3] ,
    \Tile_X1Y2_W2BEG[2] ,
    \Tile_X1Y2_W2BEG[1] ,
    \Tile_X1Y2_W2BEG[0] }),
    .W2BEGb({\Tile_X1Y2_W2BEGb[7] ,
    \Tile_X1Y2_W2BEGb[6] ,
    \Tile_X1Y2_W2BEGb[5] ,
    \Tile_X1Y2_W2BEGb[4] ,
    \Tile_X1Y2_W2BEGb[3] ,
    \Tile_X1Y2_W2BEGb[2] ,
    \Tile_X1Y2_W2BEGb[1] ,
    \Tile_X1Y2_W2BEGb[0] }),
    .W2END({\Tile_X2Y2_W2BEGb[7] ,
    \Tile_X2Y2_W2BEGb[6] ,
    \Tile_X2Y2_W2BEGb[5] ,
    \Tile_X2Y2_W2BEGb[4] ,
    \Tile_X2Y2_W2BEGb[3] ,
    \Tile_X2Y2_W2BEGb[2] ,
    \Tile_X2Y2_W2BEGb[1] ,
    \Tile_X2Y2_W2BEGb[0] }),
    .W2MID({\Tile_X2Y2_W2BEG[7] ,
    \Tile_X2Y2_W2BEG[6] ,
    \Tile_X2Y2_W2BEG[5] ,
    \Tile_X2Y2_W2BEG[4] ,
    \Tile_X2Y2_W2BEG[3] ,
    \Tile_X2Y2_W2BEG[2] ,
    \Tile_X2Y2_W2BEG[1] ,
    \Tile_X2Y2_W2BEG[0] }),
    .W6BEG({\Tile_X1Y2_W6BEG[11] ,
    \Tile_X1Y2_W6BEG[10] ,
    \Tile_X1Y2_W6BEG[9] ,
    \Tile_X1Y2_W6BEG[8] ,
    \Tile_X1Y2_W6BEG[7] ,
    \Tile_X1Y2_W6BEG[6] ,
    \Tile_X1Y2_W6BEG[5] ,
    \Tile_X1Y2_W6BEG[4] ,
    \Tile_X1Y2_W6BEG[3] ,
    \Tile_X1Y2_W6BEG[2] ,
    \Tile_X1Y2_W6BEG[1] ,
    \Tile_X1Y2_W6BEG[0] }),
    .W6END({\Tile_X2Y2_W6BEG[11] ,
    \Tile_X2Y2_W6BEG[10] ,
    \Tile_X2Y2_W6BEG[9] ,
    \Tile_X2Y2_W6BEG[8] ,
    \Tile_X2Y2_W6BEG[7] ,
    \Tile_X2Y2_W6BEG[6] ,
    \Tile_X2Y2_W6BEG[5] ,
    \Tile_X2Y2_W6BEG[4] ,
    \Tile_X2Y2_W6BEG[3] ,
    \Tile_X2Y2_W6BEG[2] ,
    \Tile_X2Y2_W6BEG[1] ,
    \Tile_X2Y2_W6BEG[0] }),
    .WW4BEG({\Tile_X1Y2_WW4BEG[15] ,
    \Tile_X1Y2_WW4BEG[14] ,
    \Tile_X1Y2_WW4BEG[13] ,
    \Tile_X1Y2_WW4BEG[12] ,
    \Tile_X1Y2_WW4BEG[11] ,
    \Tile_X1Y2_WW4BEG[10] ,
    \Tile_X1Y2_WW4BEG[9] ,
    \Tile_X1Y2_WW4BEG[8] ,
    \Tile_X1Y2_WW4BEG[7] ,
    \Tile_X1Y2_WW4BEG[6] ,
    \Tile_X1Y2_WW4BEG[5] ,
    \Tile_X1Y2_WW4BEG[4] ,
    \Tile_X1Y2_WW4BEG[3] ,
    \Tile_X1Y2_WW4BEG[2] ,
    \Tile_X1Y2_WW4BEG[1] ,
    \Tile_X1Y2_WW4BEG[0] }),
    .WW4END({\Tile_X2Y2_WW4BEG[15] ,
    \Tile_X2Y2_WW4BEG[14] ,
    \Tile_X2Y2_WW4BEG[13] ,
    \Tile_X2Y2_WW4BEG[12] ,
    \Tile_X2Y2_WW4BEG[11] ,
    \Tile_X2Y2_WW4BEG[10] ,
    \Tile_X2Y2_WW4BEG[9] ,
    \Tile_X2Y2_WW4BEG[8] ,
    \Tile_X2Y2_WW4BEG[7] ,
    \Tile_X2Y2_WW4BEG[6] ,
    \Tile_X2Y2_WW4BEG[5] ,
    \Tile_X2Y2_WW4BEG[4] ,
    \Tile_X2Y2_WW4BEG[3] ,
    \Tile_X2Y2_WW4BEG[2] ,
    \Tile_X2Y2_WW4BEG[1] ,
    \Tile_X2Y2_WW4BEG[0] }));
 LUT4AB Tile_X1Y3_LUT4AB (.Ci(Tile_X1Y4_Co),
    .Co(Tile_X1Y3_Co),
    .UserCLK(Tile_X1Y4_UserCLKo),
    .UserCLKo(Tile_X1Y3_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X1Y3_E1BEG[3] ,
    \Tile_X1Y3_E1BEG[2] ,
    \Tile_X1Y3_E1BEG[1] ,
    \Tile_X1Y3_E1BEG[0] }),
    .E1END({\Tile_X0Y3_E1BEG[3] ,
    \Tile_X0Y3_E1BEG[2] ,
    \Tile_X0Y3_E1BEG[1] ,
    \Tile_X0Y3_E1BEG[0] }),
    .E2BEG({\Tile_X1Y3_E2BEG[7] ,
    \Tile_X1Y3_E2BEG[6] ,
    \Tile_X1Y3_E2BEG[5] ,
    \Tile_X1Y3_E2BEG[4] ,
    \Tile_X1Y3_E2BEG[3] ,
    \Tile_X1Y3_E2BEG[2] ,
    \Tile_X1Y3_E2BEG[1] ,
    \Tile_X1Y3_E2BEG[0] }),
    .E2BEGb({\Tile_X1Y3_E2BEGb[7] ,
    \Tile_X1Y3_E2BEGb[6] ,
    \Tile_X1Y3_E2BEGb[5] ,
    \Tile_X1Y3_E2BEGb[4] ,
    \Tile_X1Y3_E2BEGb[3] ,
    \Tile_X1Y3_E2BEGb[2] ,
    \Tile_X1Y3_E2BEGb[1] ,
    \Tile_X1Y3_E2BEGb[0] }),
    .E2END({\Tile_X0Y3_E2BEGb[7] ,
    \Tile_X0Y3_E2BEGb[6] ,
    \Tile_X0Y3_E2BEGb[5] ,
    \Tile_X0Y3_E2BEGb[4] ,
    \Tile_X0Y3_E2BEGb[3] ,
    \Tile_X0Y3_E2BEGb[2] ,
    \Tile_X0Y3_E2BEGb[1] ,
    \Tile_X0Y3_E2BEGb[0] }),
    .E2MID({\Tile_X0Y3_E2BEG[7] ,
    \Tile_X0Y3_E2BEG[6] ,
    \Tile_X0Y3_E2BEG[5] ,
    \Tile_X0Y3_E2BEG[4] ,
    \Tile_X0Y3_E2BEG[3] ,
    \Tile_X0Y3_E2BEG[2] ,
    \Tile_X0Y3_E2BEG[1] ,
    \Tile_X0Y3_E2BEG[0] }),
    .E6BEG({\Tile_X1Y3_E6BEG[11] ,
    \Tile_X1Y3_E6BEG[10] ,
    \Tile_X1Y3_E6BEG[9] ,
    \Tile_X1Y3_E6BEG[8] ,
    \Tile_X1Y3_E6BEG[7] ,
    \Tile_X1Y3_E6BEG[6] ,
    \Tile_X1Y3_E6BEG[5] ,
    \Tile_X1Y3_E6BEG[4] ,
    \Tile_X1Y3_E6BEG[3] ,
    \Tile_X1Y3_E6BEG[2] ,
    \Tile_X1Y3_E6BEG[1] ,
    \Tile_X1Y3_E6BEG[0] }),
    .E6END({\Tile_X0Y3_E6BEG[11] ,
    \Tile_X0Y3_E6BEG[10] ,
    \Tile_X0Y3_E6BEG[9] ,
    \Tile_X0Y3_E6BEG[8] ,
    \Tile_X0Y3_E6BEG[7] ,
    \Tile_X0Y3_E6BEG[6] ,
    \Tile_X0Y3_E6BEG[5] ,
    \Tile_X0Y3_E6BEG[4] ,
    \Tile_X0Y3_E6BEG[3] ,
    \Tile_X0Y3_E6BEG[2] ,
    \Tile_X0Y3_E6BEG[1] ,
    \Tile_X0Y3_E6BEG[0] }),
    .EE4BEG({\Tile_X1Y3_EE4BEG[15] ,
    \Tile_X1Y3_EE4BEG[14] ,
    \Tile_X1Y3_EE4BEG[13] ,
    \Tile_X1Y3_EE4BEG[12] ,
    \Tile_X1Y3_EE4BEG[11] ,
    \Tile_X1Y3_EE4BEG[10] ,
    \Tile_X1Y3_EE4BEG[9] ,
    \Tile_X1Y3_EE4BEG[8] ,
    \Tile_X1Y3_EE4BEG[7] ,
    \Tile_X1Y3_EE4BEG[6] ,
    \Tile_X1Y3_EE4BEG[5] ,
    \Tile_X1Y3_EE4BEG[4] ,
    \Tile_X1Y3_EE4BEG[3] ,
    \Tile_X1Y3_EE4BEG[2] ,
    \Tile_X1Y3_EE4BEG[1] ,
    \Tile_X1Y3_EE4BEG[0] }),
    .EE4END({\Tile_X0Y3_EE4BEG[15] ,
    \Tile_X0Y3_EE4BEG[14] ,
    \Tile_X0Y3_EE4BEG[13] ,
    \Tile_X0Y3_EE4BEG[12] ,
    \Tile_X0Y3_EE4BEG[11] ,
    \Tile_X0Y3_EE4BEG[10] ,
    \Tile_X0Y3_EE4BEG[9] ,
    \Tile_X0Y3_EE4BEG[8] ,
    \Tile_X0Y3_EE4BEG[7] ,
    \Tile_X0Y3_EE4BEG[6] ,
    \Tile_X0Y3_EE4BEG[5] ,
    \Tile_X0Y3_EE4BEG[4] ,
    \Tile_X0Y3_EE4BEG[3] ,
    \Tile_X0Y3_EE4BEG[2] ,
    \Tile_X0Y3_EE4BEG[1] ,
    \Tile_X0Y3_EE4BEG[0] }),
    .FrameData({\Tile_X0Y3_FrameData_O[31] ,
    \Tile_X0Y3_FrameData_O[30] ,
    \Tile_X0Y3_FrameData_O[29] ,
    \Tile_X0Y3_FrameData_O[28] ,
    \Tile_X0Y3_FrameData_O[27] ,
    \Tile_X0Y3_FrameData_O[26] ,
    \Tile_X0Y3_FrameData_O[25] ,
    \Tile_X0Y3_FrameData_O[24] ,
    \Tile_X0Y3_FrameData_O[23] ,
    \Tile_X0Y3_FrameData_O[22] ,
    \Tile_X0Y3_FrameData_O[21] ,
    \Tile_X0Y3_FrameData_O[20] ,
    \Tile_X0Y3_FrameData_O[19] ,
    \Tile_X0Y3_FrameData_O[18] ,
    \Tile_X0Y3_FrameData_O[17] ,
    \Tile_X0Y3_FrameData_O[16] ,
    \Tile_X0Y3_FrameData_O[15] ,
    \Tile_X0Y3_FrameData_O[14] ,
    \Tile_X0Y3_FrameData_O[13] ,
    \Tile_X0Y3_FrameData_O[12] ,
    \Tile_X0Y3_FrameData_O[11] ,
    \Tile_X0Y3_FrameData_O[10] ,
    \Tile_X0Y3_FrameData_O[9] ,
    \Tile_X0Y3_FrameData_O[8] ,
    \Tile_X0Y3_FrameData_O[7] ,
    \Tile_X0Y3_FrameData_O[6] ,
    \Tile_X0Y3_FrameData_O[5] ,
    \Tile_X0Y3_FrameData_O[4] ,
    \Tile_X0Y3_FrameData_O[3] ,
    \Tile_X0Y3_FrameData_O[2] ,
    \Tile_X0Y3_FrameData_O[1] ,
    \Tile_X0Y3_FrameData_O[0] }),
    .FrameData_O({\Tile_X1Y3_FrameData_O[31] ,
    \Tile_X1Y3_FrameData_O[30] ,
    \Tile_X1Y3_FrameData_O[29] ,
    \Tile_X1Y3_FrameData_O[28] ,
    \Tile_X1Y3_FrameData_O[27] ,
    \Tile_X1Y3_FrameData_O[26] ,
    \Tile_X1Y3_FrameData_O[25] ,
    \Tile_X1Y3_FrameData_O[24] ,
    \Tile_X1Y3_FrameData_O[23] ,
    \Tile_X1Y3_FrameData_O[22] ,
    \Tile_X1Y3_FrameData_O[21] ,
    \Tile_X1Y3_FrameData_O[20] ,
    \Tile_X1Y3_FrameData_O[19] ,
    \Tile_X1Y3_FrameData_O[18] ,
    \Tile_X1Y3_FrameData_O[17] ,
    \Tile_X1Y3_FrameData_O[16] ,
    \Tile_X1Y3_FrameData_O[15] ,
    \Tile_X1Y3_FrameData_O[14] ,
    \Tile_X1Y3_FrameData_O[13] ,
    \Tile_X1Y3_FrameData_O[12] ,
    \Tile_X1Y3_FrameData_O[11] ,
    \Tile_X1Y3_FrameData_O[10] ,
    \Tile_X1Y3_FrameData_O[9] ,
    \Tile_X1Y3_FrameData_O[8] ,
    \Tile_X1Y3_FrameData_O[7] ,
    \Tile_X1Y3_FrameData_O[6] ,
    \Tile_X1Y3_FrameData_O[5] ,
    \Tile_X1Y3_FrameData_O[4] ,
    \Tile_X1Y3_FrameData_O[3] ,
    \Tile_X1Y3_FrameData_O[2] ,
    \Tile_X1Y3_FrameData_O[1] ,
    \Tile_X1Y3_FrameData_O[0] }),
    .FrameStrobe({\Tile_X1Y4_FrameStrobe_O[19] ,
    \Tile_X1Y4_FrameStrobe_O[18] ,
    \Tile_X1Y4_FrameStrobe_O[17] ,
    \Tile_X1Y4_FrameStrobe_O[16] ,
    \Tile_X1Y4_FrameStrobe_O[15] ,
    \Tile_X1Y4_FrameStrobe_O[14] ,
    \Tile_X1Y4_FrameStrobe_O[13] ,
    \Tile_X1Y4_FrameStrobe_O[12] ,
    \Tile_X1Y4_FrameStrobe_O[11] ,
    \Tile_X1Y4_FrameStrobe_O[10] ,
    \Tile_X1Y4_FrameStrobe_O[9] ,
    \Tile_X1Y4_FrameStrobe_O[8] ,
    \Tile_X1Y4_FrameStrobe_O[7] ,
    \Tile_X1Y4_FrameStrobe_O[6] ,
    \Tile_X1Y4_FrameStrobe_O[5] ,
    \Tile_X1Y4_FrameStrobe_O[4] ,
    \Tile_X1Y4_FrameStrobe_O[3] ,
    \Tile_X1Y4_FrameStrobe_O[2] ,
    \Tile_X1Y4_FrameStrobe_O[1] ,
    \Tile_X1Y4_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X1Y3_FrameStrobe_O[19] ,
    \Tile_X1Y3_FrameStrobe_O[18] ,
    \Tile_X1Y3_FrameStrobe_O[17] ,
    \Tile_X1Y3_FrameStrobe_O[16] ,
    \Tile_X1Y3_FrameStrobe_O[15] ,
    \Tile_X1Y3_FrameStrobe_O[14] ,
    \Tile_X1Y3_FrameStrobe_O[13] ,
    \Tile_X1Y3_FrameStrobe_O[12] ,
    \Tile_X1Y3_FrameStrobe_O[11] ,
    \Tile_X1Y3_FrameStrobe_O[10] ,
    \Tile_X1Y3_FrameStrobe_O[9] ,
    \Tile_X1Y3_FrameStrobe_O[8] ,
    \Tile_X1Y3_FrameStrobe_O[7] ,
    \Tile_X1Y3_FrameStrobe_O[6] ,
    \Tile_X1Y3_FrameStrobe_O[5] ,
    \Tile_X1Y3_FrameStrobe_O[4] ,
    \Tile_X1Y3_FrameStrobe_O[3] ,
    \Tile_X1Y3_FrameStrobe_O[2] ,
    \Tile_X1Y3_FrameStrobe_O[1] ,
    \Tile_X1Y3_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X1Y3_N1BEG[3] ,
    \Tile_X1Y3_N1BEG[2] ,
    \Tile_X1Y3_N1BEG[1] ,
    \Tile_X1Y3_N1BEG[0] }),
    .N1END({\Tile_X1Y4_N1BEG[3] ,
    \Tile_X1Y4_N1BEG[2] ,
    \Tile_X1Y4_N1BEG[1] ,
    \Tile_X1Y4_N1BEG[0] }),
    .N2BEG({\Tile_X1Y3_N2BEG[7] ,
    \Tile_X1Y3_N2BEG[6] ,
    \Tile_X1Y3_N2BEG[5] ,
    \Tile_X1Y3_N2BEG[4] ,
    \Tile_X1Y3_N2BEG[3] ,
    \Tile_X1Y3_N2BEG[2] ,
    \Tile_X1Y3_N2BEG[1] ,
    \Tile_X1Y3_N2BEG[0] }),
    .N2BEGb({\Tile_X1Y3_N2BEGb[7] ,
    \Tile_X1Y3_N2BEGb[6] ,
    \Tile_X1Y3_N2BEGb[5] ,
    \Tile_X1Y3_N2BEGb[4] ,
    \Tile_X1Y3_N2BEGb[3] ,
    \Tile_X1Y3_N2BEGb[2] ,
    \Tile_X1Y3_N2BEGb[1] ,
    \Tile_X1Y3_N2BEGb[0] }),
    .N2END({\Tile_X1Y4_N2BEGb[7] ,
    \Tile_X1Y4_N2BEGb[6] ,
    \Tile_X1Y4_N2BEGb[5] ,
    \Tile_X1Y4_N2BEGb[4] ,
    \Tile_X1Y4_N2BEGb[3] ,
    \Tile_X1Y4_N2BEGb[2] ,
    \Tile_X1Y4_N2BEGb[1] ,
    \Tile_X1Y4_N2BEGb[0] }),
    .N2MID({\Tile_X1Y4_N2BEG[7] ,
    \Tile_X1Y4_N2BEG[6] ,
    \Tile_X1Y4_N2BEG[5] ,
    \Tile_X1Y4_N2BEG[4] ,
    \Tile_X1Y4_N2BEG[3] ,
    \Tile_X1Y4_N2BEG[2] ,
    \Tile_X1Y4_N2BEG[1] ,
    \Tile_X1Y4_N2BEG[0] }),
    .N4BEG({\Tile_X1Y3_N4BEG[15] ,
    \Tile_X1Y3_N4BEG[14] ,
    \Tile_X1Y3_N4BEG[13] ,
    \Tile_X1Y3_N4BEG[12] ,
    \Tile_X1Y3_N4BEG[11] ,
    \Tile_X1Y3_N4BEG[10] ,
    \Tile_X1Y3_N4BEG[9] ,
    \Tile_X1Y3_N4BEG[8] ,
    \Tile_X1Y3_N4BEG[7] ,
    \Tile_X1Y3_N4BEG[6] ,
    \Tile_X1Y3_N4BEG[5] ,
    \Tile_X1Y3_N4BEG[4] ,
    \Tile_X1Y3_N4BEG[3] ,
    \Tile_X1Y3_N4BEG[2] ,
    \Tile_X1Y3_N4BEG[1] ,
    \Tile_X1Y3_N4BEG[0] }),
    .N4END({\Tile_X1Y4_N4BEG[15] ,
    \Tile_X1Y4_N4BEG[14] ,
    \Tile_X1Y4_N4BEG[13] ,
    \Tile_X1Y4_N4BEG[12] ,
    \Tile_X1Y4_N4BEG[11] ,
    \Tile_X1Y4_N4BEG[10] ,
    \Tile_X1Y4_N4BEG[9] ,
    \Tile_X1Y4_N4BEG[8] ,
    \Tile_X1Y4_N4BEG[7] ,
    \Tile_X1Y4_N4BEG[6] ,
    \Tile_X1Y4_N4BEG[5] ,
    \Tile_X1Y4_N4BEG[4] ,
    \Tile_X1Y4_N4BEG[3] ,
    \Tile_X1Y4_N4BEG[2] ,
    \Tile_X1Y4_N4BEG[1] ,
    \Tile_X1Y4_N4BEG[0] }),
    .NN4BEG({\Tile_X1Y3_NN4BEG[15] ,
    \Tile_X1Y3_NN4BEG[14] ,
    \Tile_X1Y3_NN4BEG[13] ,
    \Tile_X1Y3_NN4BEG[12] ,
    \Tile_X1Y3_NN4BEG[11] ,
    \Tile_X1Y3_NN4BEG[10] ,
    \Tile_X1Y3_NN4BEG[9] ,
    \Tile_X1Y3_NN4BEG[8] ,
    \Tile_X1Y3_NN4BEG[7] ,
    \Tile_X1Y3_NN4BEG[6] ,
    \Tile_X1Y3_NN4BEG[5] ,
    \Tile_X1Y3_NN4BEG[4] ,
    \Tile_X1Y3_NN4BEG[3] ,
    \Tile_X1Y3_NN4BEG[2] ,
    \Tile_X1Y3_NN4BEG[1] ,
    \Tile_X1Y3_NN4BEG[0] }),
    .NN4END({\Tile_X1Y4_NN4BEG[15] ,
    \Tile_X1Y4_NN4BEG[14] ,
    \Tile_X1Y4_NN4BEG[13] ,
    \Tile_X1Y4_NN4BEG[12] ,
    \Tile_X1Y4_NN4BEG[11] ,
    \Tile_X1Y4_NN4BEG[10] ,
    \Tile_X1Y4_NN4BEG[9] ,
    \Tile_X1Y4_NN4BEG[8] ,
    \Tile_X1Y4_NN4BEG[7] ,
    \Tile_X1Y4_NN4BEG[6] ,
    \Tile_X1Y4_NN4BEG[5] ,
    \Tile_X1Y4_NN4BEG[4] ,
    \Tile_X1Y4_NN4BEG[3] ,
    \Tile_X1Y4_NN4BEG[2] ,
    \Tile_X1Y4_NN4BEG[1] ,
    \Tile_X1Y4_NN4BEG[0] }),
    .S1BEG({\Tile_X1Y3_S1BEG[3] ,
    \Tile_X1Y3_S1BEG[2] ,
    \Tile_X1Y3_S1BEG[1] ,
    \Tile_X1Y3_S1BEG[0] }),
    .S1END({\Tile_X1Y2_S1BEG[3] ,
    \Tile_X1Y2_S1BEG[2] ,
    \Tile_X1Y2_S1BEG[1] ,
    \Tile_X1Y2_S1BEG[0] }),
    .S2BEG({\Tile_X1Y3_S2BEG[7] ,
    \Tile_X1Y3_S2BEG[6] ,
    \Tile_X1Y3_S2BEG[5] ,
    \Tile_X1Y3_S2BEG[4] ,
    \Tile_X1Y3_S2BEG[3] ,
    \Tile_X1Y3_S2BEG[2] ,
    \Tile_X1Y3_S2BEG[1] ,
    \Tile_X1Y3_S2BEG[0] }),
    .S2BEGb({\Tile_X1Y3_S2BEGb[7] ,
    \Tile_X1Y3_S2BEGb[6] ,
    \Tile_X1Y3_S2BEGb[5] ,
    \Tile_X1Y3_S2BEGb[4] ,
    \Tile_X1Y3_S2BEGb[3] ,
    \Tile_X1Y3_S2BEGb[2] ,
    \Tile_X1Y3_S2BEGb[1] ,
    \Tile_X1Y3_S2BEGb[0] }),
    .S2END({\Tile_X1Y2_S2BEGb[7] ,
    \Tile_X1Y2_S2BEGb[6] ,
    \Tile_X1Y2_S2BEGb[5] ,
    \Tile_X1Y2_S2BEGb[4] ,
    \Tile_X1Y2_S2BEGb[3] ,
    \Tile_X1Y2_S2BEGb[2] ,
    \Tile_X1Y2_S2BEGb[1] ,
    \Tile_X1Y2_S2BEGb[0] }),
    .S2MID({\Tile_X1Y2_S2BEG[7] ,
    \Tile_X1Y2_S2BEG[6] ,
    \Tile_X1Y2_S2BEG[5] ,
    \Tile_X1Y2_S2BEG[4] ,
    \Tile_X1Y2_S2BEG[3] ,
    \Tile_X1Y2_S2BEG[2] ,
    \Tile_X1Y2_S2BEG[1] ,
    \Tile_X1Y2_S2BEG[0] }),
    .S4BEG({\Tile_X1Y3_S4BEG[15] ,
    \Tile_X1Y3_S4BEG[14] ,
    \Tile_X1Y3_S4BEG[13] ,
    \Tile_X1Y3_S4BEG[12] ,
    \Tile_X1Y3_S4BEG[11] ,
    \Tile_X1Y3_S4BEG[10] ,
    \Tile_X1Y3_S4BEG[9] ,
    \Tile_X1Y3_S4BEG[8] ,
    \Tile_X1Y3_S4BEG[7] ,
    \Tile_X1Y3_S4BEG[6] ,
    \Tile_X1Y3_S4BEG[5] ,
    \Tile_X1Y3_S4BEG[4] ,
    \Tile_X1Y3_S4BEG[3] ,
    \Tile_X1Y3_S4BEG[2] ,
    \Tile_X1Y3_S4BEG[1] ,
    \Tile_X1Y3_S4BEG[0] }),
    .S4END({\Tile_X1Y2_S4BEG[15] ,
    \Tile_X1Y2_S4BEG[14] ,
    \Tile_X1Y2_S4BEG[13] ,
    \Tile_X1Y2_S4BEG[12] ,
    \Tile_X1Y2_S4BEG[11] ,
    \Tile_X1Y2_S4BEG[10] ,
    \Tile_X1Y2_S4BEG[9] ,
    \Tile_X1Y2_S4BEG[8] ,
    \Tile_X1Y2_S4BEG[7] ,
    \Tile_X1Y2_S4BEG[6] ,
    \Tile_X1Y2_S4BEG[5] ,
    \Tile_X1Y2_S4BEG[4] ,
    \Tile_X1Y2_S4BEG[3] ,
    \Tile_X1Y2_S4BEG[2] ,
    \Tile_X1Y2_S4BEG[1] ,
    \Tile_X1Y2_S4BEG[0] }),
    .SS4BEG({\Tile_X1Y3_SS4BEG[15] ,
    \Tile_X1Y3_SS4BEG[14] ,
    \Tile_X1Y3_SS4BEG[13] ,
    \Tile_X1Y3_SS4BEG[12] ,
    \Tile_X1Y3_SS4BEG[11] ,
    \Tile_X1Y3_SS4BEG[10] ,
    \Tile_X1Y3_SS4BEG[9] ,
    \Tile_X1Y3_SS4BEG[8] ,
    \Tile_X1Y3_SS4BEG[7] ,
    \Tile_X1Y3_SS4BEG[6] ,
    \Tile_X1Y3_SS4BEG[5] ,
    \Tile_X1Y3_SS4BEG[4] ,
    \Tile_X1Y3_SS4BEG[3] ,
    \Tile_X1Y3_SS4BEG[2] ,
    \Tile_X1Y3_SS4BEG[1] ,
    \Tile_X1Y3_SS4BEG[0] }),
    .SS4END({\Tile_X1Y2_SS4BEG[15] ,
    \Tile_X1Y2_SS4BEG[14] ,
    \Tile_X1Y2_SS4BEG[13] ,
    \Tile_X1Y2_SS4BEG[12] ,
    \Tile_X1Y2_SS4BEG[11] ,
    \Tile_X1Y2_SS4BEG[10] ,
    \Tile_X1Y2_SS4BEG[9] ,
    \Tile_X1Y2_SS4BEG[8] ,
    \Tile_X1Y2_SS4BEG[7] ,
    \Tile_X1Y2_SS4BEG[6] ,
    \Tile_X1Y2_SS4BEG[5] ,
    \Tile_X1Y2_SS4BEG[4] ,
    \Tile_X1Y2_SS4BEG[3] ,
    \Tile_X1Y2_SS4BEG[2] ,
    \Tile_X1Y2_SS4BEG[1] ,
    \Tile_X1Y2_SS4BEG[0] }),
    .W1BEG({\Tile_X1Y3_W1BEG[3] ,
    \Tile_X1Y3_W1BEG[2] ,
    \Tile_X1Y3_W1BEG[1] ,
    \Tile_X1Y3_W1BEG[0] }),
    .W1END({\Tile_X2Y3_W1BEG[3] ,
    \Tile_X2Y3_W1BEG[2] ,
    \Tile_X2Y3_W1BEG[1] ,
    \Tile_X2Y3_W1BEG[0] }),
    .W2BEG({\Tile_X1Y3_W2BEG[7] ,
    \Tile_X1Y3_W2BEG[6] ,
    \Tile_X1Y3_W2BEG[5] ,
    \Tile_X1Y3_W2BEG[4] ,
    \Tile_X1Y3_W2BEG[3] ,
    \Tile_X1Y3_W2BEG[2] ,
    \Tile_X1Y3_W2BEG[1] ,
    \Tile_X1Y3_W2BEG[0] }),
    .W2BEGb({\Tile_X1Y3_W2BEGb[7] ,
    \Tile_X1Y3_W2BEGb[6] ,
    \Tile_X1Y3_W2BEGb[5] ,
    \Tile_X1Y3_W2BEGb[4] ,
    \Tile_X1Y3_W2BEGb[3] ,
    \Tile_X1Y3_W2BEGb[2] ,
    \Tile_X1Y3_W2BEGb[1] ,
    \Tile_X1Y3_W2BEGb[0] }),
    .W2END({\Tile_X2Y3_W2BEGb[7] ,
    \Tile_X2Y3_W2BEGb[6] ,
    \Tile_X2Y3_W2BEGb[5] ,
    \Tile_X2Y3_W2BEGb[4] ,
    \Tile_X2Y3_W2BEGb[3] ,
    \Tile_X2Y3_W2BEGb[2] ,
    \Tile_X2Y3_W2BEGb[1] ,
    \Tile_X2Y3_W2BEGb[0] }),
    .W2MID({\Tile_X2Y3_W2BEG[7] ,
    \Tile_X2Y3_W2BEG[6] ,
    \Tile_X2Y3_W2BEG[5] ,
    \Tile_X2Y3_W2BEG[4] ,
    \Tile_X2Y3_W2BEG[3] ,
    \Tile_X2Y3_W2BEG[2] ,
    \Tile_X2Y3_W2BEG[1] ,
    \Tile_X2Y3_W2BEG[0] }),
    .W6BEG({\Tile_X1Y3_W6BEG[11] ,
    \Tile_X1Y3_W6BEG[10] ,
    \Tile_X1Y3_W6BEG[9] ,
    \Tile_X1Y3_W6BEG[8] ,
    \Tile_X1Y3_W6BEG[7] ,
    \Tile_X1Y3_W6BEG[6] ,
    \Tile_X1Y3_W6BEG[5] ,
    \Tile_X1Y3_W6BEG[4] ,
    \Tile_X1Y3_W6BEG[3] ,
    \Tile_X1Y3_W6BEG[2] ,
    \Tile_X1Y3_W6BEG[1] ,
    \Tile_X1Y3_W6BEG[0] }),
    .W6END({\Tile_X2Y3_W6BEG[11] ,
    \Tile_X2Y3_W6BEG[10] ,
    \Tile_X2Y3_W6BEG[9] ,
    \Tile_X2Y3_W6BEG[8] ,
    \Tile_X2Y3_W6BEG[7] ,
    \Tile_X2Y3_W6BEG[6] ,
    \Tile_X2Y3_W6BEG[5] ,
    \Tile_X2Y3_W6BEG[4] ,
    \Tile_X2Y3_W6BEG[3] ,
    \Tile_X2Y3_W6BEG[2] ,
    \Tile_X2Y3_W6BEG[1] ,
    \Tile_X2Y3_W6BEG[0] }),
    .WW4BEG({\Tile_X1Y3_WW4BEG[15] ,
    \Tile_X1Y3_WW4BEG[14] ,
    \Tile_X1Y3_WW4BEG[13] ,
    \Tile_X1Y3_WW4BEG[12] ,
    \Tile_X1Y3_WW4BEG[11] ,
    \Tile_X1Y3_WW4BEG[10] ,
    \Tile_X1Y3_WW4BEG[9] ,
    \Tile_X1Y3_WW4BEG[8] ,
    \Tile_X1Y3_WW4BEG[7] ,
    \Tile_X1Y3_WW4BEG[6] ,
    \Tile_X1Y3_WW4BEG[5] ,
    \Tile_X1Y3_WW4BEG[4] ,
    \Tile_X1Y3_WW4BEG[3] ,
    \Tile_X1Y3_WW4BEG[2] ,
    \Tile_X1Y3_WW4BEG[1] ,
    \Tile_X1Y3_WW4BEG[0] }),
    .WW4END({\Tile_X2Y3_WW4BEG[15] ,
    \Tile_X2Y3_WW4BEG[14] ,
    \Tile_X2Y3_WW4BEG[13] ,
    \Tile_X2Y3_WW4BEG[12] ,
    \Tile_X2Y3_WW4BEG[11] ,
    \Tile_X2Y3_WW4BEG[10] ,
    \Tile_X2Y3_WW4BEG[9] ,
    \Tile_X2Y3_WW4BEG[8] ,
    \Tile_X2Y3_WW4BEG[7] ,
    \Tile_X2Y3_WW4BEG[6] ,
    \Tile_X2Y3_WW4BEG[5] ,
    \Tile_X2Y3_WW4BEG[4] ,
    \Tile_X2Y3_WW4BEG[3] ,
    \Tile_X2Y3_WW4BEG[2] ,
    \Tile_X2Y3_WW4BEG[1] ,
    \Tile_X2Y3_WW4BEG[0] }));
 LUT4AB Tile_X1Y4_LUT4AB (.Ci(Tile_X1Y5_Co),
    .Co(Tile_X1Y4_Co),
    .UserCLK(Tile_X1Y5_UserCLKo),
    .UserCLKo(Tile_X1Y4_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X1Y4_E1BEG[3] ,
    \Tile_X1Y4_E1BEG[2] ,
    \Tile_X1Y4_E1BEG[1] ,
    \Tile_X1Y4_E1BEG[0] }),
    .E1END({\Tile_X0Y4_E1BEG[3] ,
    \Tile_X0Y4_E1BEG[2] ,
    \Tile_X0Y4_E1BEG[1] ,
    \Tile_X0Y4_E1BEG[0] }),
    .E2BEG({\Tile_X1Y4_E2BEG[7] ,
    \Tile_X1Y4_E2BEG[6] ,
    \Tile_X1Y4_E2BEG[5] ,
    \Tile_X1Y4_E2BEG[4] ,
    \Tile_X1Y4_E2BEG[3] ,
    \Tile_X1Y4_E2BEG[2] ,
    \Tile_X1Y4_E2BEG[1] ,
    \Tile_X1Y4_E2BEG[0] }),
    .E2BEGb({\Tile_X1Y4_E2BEGb[7] ,
    \Tile_X1Y4_E2BEGb[6] ,
    \Tile_X1Y4_E2BEGb[5] ,
    \Tile_X1Y4_E2BEGb[4] ,
    \Tile_X1Y4_E2BEGb[3] ,
    \Tile_X1Y4_E2BEGb[2] ,
    \Tile_X1Y4_E2BEGb[1] ,
    \Tile_X1Y4_E2BEGb[0] }),
    .E2END({\Tile_X0Y4_E2BEGb[7] ,
    \Tile_X0Y4_E2BEGb[6] ,
    \Tile_X0Y4_E2BEGb[5] ,
    \Tile_X0Y4_E2BEGb[4] ,
    \Tile_X0Y4_E2BEGb[3] ,
    \Tile_X0Y4_E2BEGb[2] ,
    \Tile_X0Y4_E2BEGb[1] ,
    \Tile_X0Y4_E2BEGb[0] }),
    .E2MID({\Tile_X0Y4_E2BEG[7] ,
    \Tile_X0Y4_E2BEG[6] ,
    \Tile_X0Y4_E2BEG[5] ,
    \Tile_X0Y4_E2BEG[4] ,
    \Tile_X0Y4_E2BEG[3] ,
    \Tile_X0Y4_E2BEG[2] ,
    \Tile_X0Y4_E2BEG[1] ,
    \Tile_X0Y4_E2BEG[0] }),
    .E6BEG({\Tile_X1Y4_E6BEG[11] ,
    \Tile_X1Y4_E6BEG[10] ,
    \Tile_X1Y4_E6BEG[9] ,
    \Tile_X1Y4_E6BEG[8] ,
    \Tile_X1Y4_E6BEG[7] ,
    \Tile_X1Y4_E6BEG[6] ,
    \Tile_X1Y4_E6BEG[5] ,
    \Tile_X1Y4_E6BEG[4] ,
    \Tile_X1Y4_E6BEG[3] ,
    \Tile_X1Y4_E6BEG[2] ,
    \Tile_X1Y4_E6BEG[1] ,
    \Tile_X1Y4_E6BEG[0] }),
    .E6END({\Tile_X0Y4_E6BEG[11] ,
    \Tile_X0Y4_E6BEG[10] ,
    \Tile_X0Y4_E6BEG[9] ,
    \Tile_X0Y4_E6BEG[8] ,
    \Tile_X0Y4_E6BEG[7] ,
    \Tile_X0Y4_E6BEG[6] ,
    \Tile_X0Y4_E6BEG[5] ,
    \Tile_X0Y4_E6BEG[4] ,
    \Tile_X0Y4_E6BEG[3] ,
    \Tile_X0Y4_E6BEG[2] ,
    \Tile_X0Y4_E6BEG[1] ,
    \Tile_X0Y4_E6BEG[0] }),
    .EE4BEG({\Tile_X1Y4_EE4BEG[15] ,
    \Tile_X1Y4_EE4BEG[14] ,
    \Tile_X1Y4_EE4BEG[13] ,
    \Tile_X1Y4_EE4BEG[12] ,
    \Tile_X1Y4_EE4BEG[11] ,
    \Tile_X1Y4_EE4BEG[10] ,
    \Tile_X1Y4_EE4BEG[9] ,
    \Tile_X1Y4_EE4BEG[8] ,
    \Tile_X1Y4_EE4BEG[7] ,
    \Tile_X1Y4_EE4BEG[6] ,
    \Tile_X1Y4_EE4BEG[5] ,
    \Tile_X1Y4_EE4BEG[4] ,
    \Tile_X1Y4_EE4BEG[3] ,
    \Tile_X1Y4_EE4BEG[2] ,
    \Tile_X1Y4_EE4BEG[1] ,
    \Tile_X1Y4_EE4BEG[0] }),
    .EE4END({\Tile_X0Y4_EE4BEG[15] ,
    \Tile_X0Y4_EE4BEG[14] ,
    \Tile_X0Y4_EE4BEG[13] ,
    \Tile_X0Y4_EE4BEG[12] ,
    \Tile_X0Y4_EE4BEG[11] ,
    \Tile_X0Y4_EE4BEG[10] ,
    \Tile_X0Y4_EE4BEG[9] ,
    \Tile_X0Y4_EE4BEG[8] ,
    \Tile_X0Y4_EE4BEG[7] ,
    \Tile_X0Y4_EE4BEG[6] ,
    \Tile_X0Y4_EE4BEG[5] ,
    \Tile_X0Y4_EE4BEG[4] ,
    \Tile_X0Y4_EE4BEG[3] ,
    \Tile_X0Y4_EE4BEG[2] ,
    \Tile_X0Y4_EE4BEG[1] ,
    \Tile_X0Y4_EE4BEG[0] }),
    .FrameData({\Tile_X0Y4_FrameData_O[31] ,
    \Tile_X0Y4_FrameData_O[30] ,
    \Tile_X0Y4_FrameData_O[29] ,
    \Tile_X0Y4_FrameData_O[28] ,
    \Tile_X0Y4_FrameData_O[27] ,
    \Tile_X0Y4_FrameData_O[26] ,
    \Tile_X0Y4_FrameData_O[25] ,
    \Tile_X0Y4_FrameData_O[24] ,
    \Tile_X0Y4_FrameData_O[23] ,
    \Tile_X0Y4_FrameData_O[22] ,
    \Tile_X0Y4_FrameData_O[21] ,
    \Tile_X0Y4_FrameData_O[20] ,
    \Tile_X0Y4_FrameData_O[19] ,
    \Tile_X0Y4_FrameData_O[18] ,
    \Tile_X0Y4_FrameData_O[17] ,
    \Tile_X0Y4_FrameData_O[16] ,
    \Tile_X0Y4_FrameData_O[15] ,
    \Tile_X0Y4_FrameData_O[14] ,
    \Tile_X0Y4_FrameData_O[13] ,
    \Tile_X0Y4_FrameData_O[12] ,
    \Tile_X0Y4_FrameData_O[11] ,
    \Tile_X0Y4_FrameData_O[10] ,
    \Tile_X0Y4_FrameData_O[9] ,
    \Tile_X0Y4_FrameData_O[8] ,
    \Tile_X0Y4_FrameData_O[7] ,
    \Tile_X0Y4_FrameData_O[6] ,
    \Tile_X0Y4_FrameData_O[5] ,
    \Tile_X0Y4_FrameData_O[4] ,
    \Tile_X0Y4_FrameData_O[3] ,
    \Tile_X0Y4_FrameData_O[2] ,
    \Tile_X0Y4_FrameData_O[1] ,
    \Tile_X0Y4_FrameData_O[0] }),
    .FrameData_O({\Tile_X1Y4_FrameData_O[31] ,
    \Tile_X1Y4_FrameData_O[30] ,
    \Tile_X1Y4_FrameData_O[29] ,
    \Tile_X1Y4_FrameData_O[28] ,
    \Tile_X1Y4_FrameData_O[27] ,
    \Tile_X1Y4_FrameData_O[26] ,
    \Tile_X1Y4_FrameData_O[25] ,
    \Tile_X1Y4_FrameData_O[24] ,
    \Tile_X1Y4_FrameData_O[23] ,
    \Tile_X1Y4_FrameData_O[22] ,
    \Tile_X1Y4_FrameData_O[21] ,
    \Tile_X1Y4_FrameData_O[20] ,
    \Tile_X1Y4_FrameData_O[19] ,
    \Tile_X1Y4_FrameData_O[18] ,
    \Tile_X1Y4_FrameData_O[17] ,
    \Tile_X1Y4_FrameData_O[16] ,
    \Tile_X1Y4_FrameData_O[15] ,
    \Tile_X1Y4_FrameData_O[14] ,
    \Tile_X1Y4_FrameData_O[13] ,
    \Tile_X1Y4_FrameData_O[12] ,
    \Tile_X1Y4_FrameData_O[11] ,
    \Tile_X1Y4_FrameData_O[10] ,
    \Tile_X1Y4_FrameData_O[9] ,
    \Tile_X1Y4_FrameData_O[8] ,
    \Tile_X1Y4_FrameData_O[7] ,
    \Tile_X1Y4_FrameData_O[6] ,
    \Tile_X1Y4_FrameData_O[5] ,
    \Tile_X1Y4_FrameData_O[4] ,
    \Tile_X1Y4_FrameData_O[3] ,
    \Tile_X1Y4_FrameData_O[2] ,
    \Tile_X1Y4_FrameData_O[1] ,
    \Tile_X1Y4_FrameData_O[0] }),
    .FrameStrobe({\Tile_X1Y5_FrameStrobe_O[19] ,
    \Tile_X1Y5_FrameStrobe_O[18] ,
    \Tile_X1Y5_FrameStrobe_O[17] ,
    \Tile_X1Y5_FrameStrobe_O[16] ,
    \Tile_X1Y5_FrameStrobe_O[15] ,
    \Tile_X1Y5_FrameStrobe_O[14] ,
    \Tile_X1Y5_FrameStrobe_O[13] ,
    \Tile_X1Y5_FrameStrobe_O[12] ,
    \Tile_X1Y5_FrameStrobe_O[11] ,
    \Tile_X1Y5_FrameStrobe_O[10] ,
    \Tile_X1Y5_FrameStrobe_O[9] ,
    \Tile_X1Y5_FrameStrobe_O[8] ,
    \Tile_X1Y5_FrameStrobe_O[7] ,
    \Tile_X1Y5_FrameStrobe_O[6] ,
    \Tile_X1Y5_FrameStrobe_O[5] ,
    \Tile_X1Y5_FrameStrobe_O[4] ,
    \Tile_X1Y5_FrameStrobe_O[3] ,
    \Tile_X1Y5_FrameStrobe_O[2] ,
    \Tile_X1Y5_FrameStrobe_O[1] ,
    \Tile_X1Y5_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X1Y4_FrameStrobe_O[19] ,
    \Tile_X1Y4_FrameStrobe_O[18] ,
    \Tile_X1Y4_FrameStrobe_O[17] ,
    \Tile_X1Y4_FrameStrobe_O[16] ,
    \Tile_X1Y4_FrameStrobe_O[15] ,
    \Tile_X1Y4_FrameStrobe_O[14] ,
    \Tile_X1Y4_FrameStrobe_O[13] ,
    \Tile_X1Y4_FrameStrobe_O[12] ,
    \Tile_X1Y4_FrameStrobe_O[11] ,
    \Tile_X1Y4_FrameStrobe_O[10] ,
    \Tile_X1Y4_FrameStrobe_O[9] ,
    \Tile_X1Y4_FrameStrobe_O[8] ,
    \Tile_X1Y4_FrameStrobe_O[7] ,
    \Tile_X1Y4_FrameStrobe_O[6] ,
    \Tile_X1Y4_FrameStrobe_O[5] ,
    \Tile_X1Y4_FrameStrobe_O[4] ,
    \Tile_X1Y4_FrameStrobe_O[3] ,
    \Tile_X1Y4_FrameStrobe_O[2] ,
    \Tile_X1Y4_FrameStrobe_O[1] ,
    \Tile_X1Y4_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X1Y4_N1BEG[3] ,
    \Tile_X1Y4_N1BEG[2] ,
    \Tile_X1Y4_N1BEG[1] ,
    \Tile_X1Y4_N1BEG[0] }),
    .N1END({\Tile_X1Y5_N1BEG[3] ,
    \Tile_X1Y5_N1BEG[2] ,
    \Tile_X1Y5_N1BEG[1] ,
    \Tile_X1Y5_N1BEG[0] }),
    .N2BEG({\Tile_X1Y4_N2BEG[7] ,
    \Tile_X1Y4_N2BEG[6] ,
    \Tile_X1Y4_N2BEG[5] ,
    \Tile_X1Y4_N2BEG[4] ,
    \Tile_X1Y4_N2BEG[3] ,
    \Tile_X1Y4_N2BEG[2] ,
    \Tile_X1Y4_N2BEG[1] ,
    \Tile_X1Y4_N2BEG[0] }),
    .N2BEGb({\Tile_X1Y4_N2BEGb[7] ,
    \Tile_X1Y4_N2BEGb[6] ,
    \Tile_X1Y4_N2BEGb[5] ,
    \Tile_X1Y4_N2BEGb[4] ,
    \Tile_X1Y4_N2BEGb[3] ,
    \Tile_X1Y4_N2BEGb[2] ,
    \Tile_X1Y4_N2BEGb[1] ,
    \Tile_X1Y4_N2BEGb[0] }),
    .N2END({\Tile_X1Y5_N2BEGb[7] ,
    \Tile_X1Y5_N2BEGb[6] ,
    \Tile_X1Y5_N2BEGb[5] ,
    \Tile_X1Y5_N2BEGb[4] ,
    \Tile_X1Y5_N2BEGb[3] ,
    \Tile_X1Y5_N2BEGb[2] ,
    \Tile_X1Y5_N2BEGb[1] ,
    \Tile_X1Y5_N2BEGb[0] }),
    .N2MID({\Tile_X1Y5_N2BEG[7] ,
    \Tile_X1Y5_N2BEG[6] ,
    \Tile_X1Y5_N2BEG[5] ,
    \Tile_X1Y5_N2BEG[4] ,
    \Tile_X1Y5_N2BEG[3] ,
    \Tile_X1Y5_N2BEG[2] ,
    \Tile_X1Y5_N2BEG[1] ,
    \Tile_X1Y5_N2BEG[0] }),
    .N4BEG({\Tile_X1Y4_N4BEG[15] ,
    \Tile_X1Y4_N4BEG[14] ,
    \Tile_X1Y4_N4BEG[13] ,
    \Tile_X1Y4_N4BEG[12] ,
    \Tile_X1Y4_N4BEG[11] ,
    \Tile_X1Y4_N4BEG[10] ,
    \Tile_X1Y4_N4BEG[9] ,
    \Tile_X1Y4_N4BEG[8] ,
    \Tile_X1Y4_N4BEG[7] ,
    \Tile_X1Y4_N4BEG[6] ,
    \Tile_X1Y4_N4BEG[5] ,
    \Tile_X1Y4_N4BEG[4] ,
    \Tile_X1Y4_N4BEG[3] ,
    \Tile_X1Y4_N4BEG[2] ,
    \Tile_X1Y4_N4BEG[1] ,
    \Tile_X1Y4_N4BEG[0] }),
    .N4END({\Tile_X1Y5_N4BEG[15] ,
    \Tile_X1Y5_N4BEG[14] ,
    \Tile_X1Y5_N4BEG[13] ,
    \Tile_X1Y5_N4BEG[12] ,
    \Tile_X1Y5_N4BEG[11] ,
    \Tile_X1Y5_N4BEG[10] ,
    \Tile_X1Y5_N4BEG[9] ,
    \Tile_X1Y5_N4BEG[8] ,
    \Tile_X1Y5_N4BEG[7] ,
    \Tile_X1Y5_N4BEG[6] ,
    \Tile_X1Y5_N4BEG[5] ,
    \Tile_X1Y5_N4BEG[4] ,
    \Tile_X1Y5_N4BEG[3] ,
    \Tile_X1Y5_N4BEG[2] ,
    \Tile_X1Y5_N4BEG[1] ,
    \Tile_X1Y5_N4BEG[0] }),
    .NN4BEG({\Tile_X1Y4_NN4BEG[15] ,
    \Tile_X1Y4_NN4BEG[14] ,
    \Tile_X1Y4_NN4BEG[13] ,
    \Tile_X1Y4_NN4BEG[12] ,
    \Tile_X1Y4_NN4BEG[11] ,
    \Tile_X1Y4_NN4BEG[10] ,
    \Tile_X1Y4_NN4BEG[9] ,
    \Tile_X1Y4_NN4BEG[8] ,
    \Tile_X1Y4_NN4BEG[7] ,
    \Tile_X1Y4_NN4BEG[6] ,
    \Tile_X1Y4_NN4BEG[5] ,
    \Tile_X1Y4_NN4BEG[4] ,
    \Tile_X1Y4_NN4BEG[3] ,
    \Tile_X1Y4_NN4BEG[2] ,
    \Tile_X1Y4_NN4BEG[1] ,
    \Tile_X1Y4_NN4BEG[0] }),
    .NN4END({\Tile_X1Y5_NN4BEG[15] ,
    \Tile_X1Y5_NN4BEG[14] ,
    \Tile_X1Y5_NN4BEG[13] ,
    \Tile_X1Y5_NN4BEG[12] ,
    \Tile_X1Y5_NN4BEG[11] ,
    \Tile_X1Y5_NN4BEG[10] ,
    \Tile_X1Y5_NN4BEG[9] ,
    \Tile_X1Y5_NN4BEG[8] ,
    \Tile_X1Y5_NN4BEG[7] ,
    \Tile_X1Y5_NN4BEG[6] ,
    \Tile_X1Y5_NN4BEG[5] ,
    \Tile_X1Y5_NN4BEG[4] ,
    \Tile_X1Y5_NN4BEG[3] ,
    \Tile_X1Y5_NN4BEG[2] ,
    \Tile_X1Y5_NN4BEG[1] ,
    \Tile_X1Y5_NN4BEG[0] }),
    .S1BEG({\Tile_X1Y4_S1BEG[3] ,
    \Tile_X1Y4_S1BEG[2] ,
    \Tile_X1Y4_S1BEG[1] ,
    \Tile_X1Y4_S1BEG[0] }),
    .S1END({\Tile_X1Y3_S1BEG[3] ,
    \Tile_X1Y3_S1BEG[2] ,
    \Tile_X1Y3_S1BEG[1] ,
    \Tile_X1Y3_S1BEG[0] }),
    .S2BEG({\Tile_X1Y4_S2BEG[7] ,
    \Tile_X1Y4_S2BEG[6] ,
    \Tile_X1Y4_S2BEG[5] ,
    \Tile_X1Y4_S2BEG[4] ,
    \Tile_X1Y4_S2BEG[3] ,
    \Tile_X1Y4_S2BEG[2] ,
    \Tile_X1Y4_S2BEG[1] ,
    \Tile_X1Y4_S2BEG[0] }),
    .S2BEGb({\Tile_X1Y4_S2BEGb[7] ,
    \Tile_X1Y4_S2BEGb[6] ,
    \Tile_X1Y4_S2BEGb[5] ,
    \Tile_X1Y4_S2BEGb[4] ,
    \Tile_X1Y4_S2BEGb[3] ,
    \Tile_X1Y4_S2BEGb[2] ,
    \Tile_X1Y4_S2BEGb[1] ,
    \Tile_X1Y4_S2BEGb[0] }),
    .S2END({\Tile_X1Y3_S2BEGb[7] ,
    \Tile_X1Y3_S2BEGb[6] ,
    \Tile_X1Y3_S2BEGb[5] ,
    \Tile_X1Y3_S2BEGb[4] ,
    \Tile_X1Y3_S2BEGb[3] ,
    \Tile_X1Y3_S2BEGb[2] ,
    \Tile_X1Y3_S2BEGb[1] ,
    \Tile_X1Y3_S2BEGb[0] }),
    .S2MID({\Tile_X1Y3_S2BEG[7] ,
    \Tile_X1Y3_S2BEG[6] ,
    \Tile_X1Y3_S2BEG[5] ,
    \Tile_X1Y3_S2BEG[4] ,
    \Tile_X1Y3_S2BEG[3] ,
    \Tile_X1Y3_S2BEG[2] ,
    \Tile_X1Y3_S2BEG[1] ,
    \Tile_X1Y3_S2BEG[0] }),
    .S4BEG({\Tile_X1Y4_S4BEG[15] ,
    \Tile_X1Y4_S4BEG[14] ,
    \Tile_X1Y4_S4BEG[13] ,
    \Tile_X1Y4_S4BEG[12] ,
    \Tile_X1Y4_S4BEG[11] ,
    \Tile_X1Y4_S4BEG[10] ,
    \Tile_X1Y4_S4BEG[9] ,
    \Tile_X1Y4_S4BEG[8] ,
    \Tile_X1Y4_S4BEG[7] ,
    \Tile_X1Y4_S4BEG[6] ,
    \Tile_X1Y4_S4BEG[5] ,
    \Tile_X1Y4_S4BEG[4] ,
    \Tile_X1Y4_S4BEG[3] ,
    \Tile_X1Y4_S4BEG[2] ,
    \Tile_X1Y4_S4BEG[1] ,
    \Tile_X1Y4_S4BEG[0] }),
    .S4END({\Tile_X1Y3_S4BEG[15] ,
    \Tile_X1Y3_S4BEG[14] ,
    \Tile_X1Y3_S4BEG[13] ,
    \Tile_X1Y3_S4BEG[12] ,
    \Tile_X1Y3_S4BEG[11] ,
    \Tile_X1Y3_S4BEG[10] ,
    \Tile_X1Y3_S4BEG[9] ,
    \Tile_X1Y3_S4BEG[8] ,
    \Tile_X1Y3_S4BEG[7] ,
    \Tile_X1Y3_S4BEG[6] ,
    \Tile_X1Y3_S4BEG[5] ,
    \Tile_X1Y3_S4BEG[4] ,
    \Tile_X1Y3_S4BEG[3] ,
    \Tile_X1Y3_S4BEG[2] ,
    \Tile_X1Y3_S4BEG[1] ,
    \Tile_X1Y3_S4BEG[0] }),
    .SS4BEG({\Tile_X1Y4_SS4BEG[15] ,
    \Tile_X1Y4_SS4BEG[14] ,
    \Tile_X1Y4_SS4BEG[13] ,
    \Tile_X1Y4_SS4BEG[12] ,
    \Tile_X1Y4_SS4BEG[11] ,
    \Tile_X1Y4_SS4BEG[10] ,
    \Tile_X1Y4_SS4BEG[9] ,
    \Tile_X1Y4_SS4BEG[8] ,
    \Tile_X1Y4_SS4BEG[7] ,
    \Tile_X1Y4_SS4BEG[6] ,
    \Tile_X1Y4_SS4BEG[5] ,
    \Tile_X1Y4_SS4BEG[4] ,
    \Tile_X1Y4_SS4BEG[3] ,
    \Tile_X1Y4_SS4BEG[2] ,
    \Tile_X1Y4_SS4BEG[1] ,
    \Tile_X1Y4_SS4BEG[0] }),
    .SS4END({\Tile_X1Y3_SS4BEG[15] ,
    \Tile_X1Y3_SS4BEG[14] ,
    \Tile_X1Y3_SS4BEG[13] ,
    \Tile_X1Y3_SS4BEG[12] ,
    \Tile_X1Y3_SS4BEG[11] ,
    \Tile_X1Y3_SS4BEG[10] ,
    \Tile_X1Y3_SS4BEG[9] ,
    \Tile_X1Y3_SS4BEG[8] ,
    \Tile_X1Y3_SS4BEG[7] ,
    \Tile_X1Y3_SS4BEG[6] ,
    \Tile_X1Y3_SS4BEG[5] ,
    \Tile_X1Y3_SS4BEG[4] ,
    \Tile_X1Y3_SS4BEG[3] ,
    \Tile_X1Y3_SS4BEG[2] ,
    \Tile_X1Y3_SS4BEG[1] ,
    \Tile_X1Y3_SS4BEG[0] }),
    .W1BEG({\Tile_X1Y4_W1BEG[3] ,
    \Tile_X1Y4_W1BEG[2] ,
    \Tile_X1Y4_W1BEG[1] ,
    \Tile_X1Y4_W1BEG[0] }),
    .W1END({\Tile_X2Y4_W1BEG[3] ,
    \Tile_X2Y4_W1BEG[2] ,
    \Tile_X2Y4_W1BEG[1] ,
    \Tile_X2Y4_W1BEG[0] }),
    .W2BEG({\Tile_X1Y4_W2BEG[7] ,
    \Tile_X1Y4_W2BEG[6] ,
    \Tile_X1Y4_W2BEG[5] ,
    \Tile_X1Y4_W2BEG[4] ,
    \Tile_X1Y4_W2BEG[3] ,
    \Tile_X1Y4_W2BEG[2] ,
    \Tile_X1Y4_W2BEG[1] ,
    \Tile_X1Y4_W2BEG[0] }),
    .W2BEGb({\Tile_X1Y4_W2BEGb[7] ,
    \Tile_X1Y4_W2BEGb[6] ,
    \Tile_X1Y4_W2BEGb[5] ,
    \Tile_X1Y4_W2BEGb[4] ,
    \Tile_X1Y4_W2BEGb[3] ,
    \Tile_X1Y4_W2BEGb[2] ,
    \Tile_X1Y4_W2BEGb[1] ,
    \Tile_X1Y4_W2BEGb[0] }),
    .W2END({\Tile_X2Y4_W2BEGb[7] ,
    \Tile_X2Y4_W2BEGb[6] ,
    \Tile_X2Y4_W2BEGb[5] ,
    \Tile_X2Y4_W2BEGb[4] ,
    \Tile_X2Y4_W2BEGb[3] ,
    \Tile_X2Y4_W2BEGb[2] ,
    \Tile_X2Y4_W2BEGb[1] ,
    \Tile_X2Y4_W2BEGb[0] }),
    .W2MID({\Tile_X2Y4_W2BEG[7] ,
    \Tile_X2Y4_W2BEG[6] ,
    \Tile_X2Y4_W2BEG[5] ,
    \Tile_X2Y4_W2BEG[4] ,
    \Tile_X2Y4_W2BEG[3] ,
    \Tile_X2Y4_W2BEG[2] ,
    \Tile_X2Y4_W2BEG[1] ,
    \Tile_X2Y4_W2BEG[0] }),
    .W6BEG({\Tile_X1Y4_W6BEG[11] ,
    \Tile_X1Y4_W6BEG[10] ,
    \Tile_X1Y4_W6BEG[9] ,
    \Tile_X1Y4_W6BEG[8] ,
    \Tile_X1Y4_W6BEG[7] ,
    \Tile_X1Y4_W6BEG[6] ,
    \Tile_X1Y4_W6BEG[5] ,
    \Tile_X1Y4_W6BEG[4] ,
    \Tile_X1Y4_W6BEG[3] ,
    \Tile_X1Y4_W6BEG[2] ,
    \Tile_X1Y4_W6BEG[1] ,
    \Tile_X1Y4_W6BEG[0] }),
    .W6END({\Tile_X2Y4_W6BEG[11] ,
    \Tile_X2Y4_W6BEG[10] ,
    \Tile_X2Y4_W6BEG[9] ,
    \Tile_X2Y4_W6BEG[8] ,
    \Tile_X2Y4_W6BEG[7] ,
    \Tile_X2Y4_W6BEG[6] ,
    \Tile_X2Y4_W6BEG[5] ,
    \Tile_X2Y4_W6BEG[4] ,
    \Tile_X2Y4_W6BEG[3] ,
    \Tile_X2Y4_W6BEG[2] ,
    \Tile_X2Y4_W6BEG[1] ,
    \Tile_X2Y4_W6BEG[0] }),
    .WW4BEG({\Tile_X1Y4_WW4BEG[15] ,
    \Tile_X1Y4_WW4BEG[14] ,
    \Tile_X1Y4_WW4BEG[13] ,
    \Tile_X1Y4_WW4BEG[12] ,
    \Tile_X1Y4_WW4BEG[11] ,
    \Tile_X1Y4_WW4BEG[10] ,
    \Tile_X1Y4_WW4BEG[9] ,
    \Tile_X1Y4_WW4BEG[8] ,
    \Tile_X1Y4_WW4BEG[7] ,
    \Tile_X1Y4_WW4BEG[6] ,
    \Tile_X1Y4_WW4BEG[5] ,
    \Tile_X1Y4_WW4BEG[4] ,
    \Tile_X1Y4_WW4BEG[3] ,
    \Tile_X1Y4_WW4BEG[2] ,
    \Tile_X1Y4_WW4BEG[1] ,
    \Tile_X1Y4_WW4BEG[0] }),
    .WW4END({\Tile_X2Y4_WW4BEG[15] ,
    \Tile_X2Y4_WW4BEG[14] ,
    \Tile_X2Y4_WW4BEG[13] ,
    \Tile_X2Y4_WW4BEG[12] ,
    \Tile_X2Y4_WW4BEG[11] ,
    \Tile_X2Y4_WW4BEG[10] ,
    \Tile_X2Y4_WW4BEG[9] ,
    \Tile_X2Y4_WW4BEG[8] ,
    \Tile_X2Y4_WW4BEG[7] ,
    \Tile_X2Y4_WW4BEG[6] ,
    \Tile_X2Y4_WW4BEG[5] ,
    \Tile_X2Y4_WW4BEG[4] ,
    \Tile_X2Y4_WW4BEG[3] ,
    \Tile_X2Y4_WW4BEG[2] ,
    \Tile_X2Y4_WW4BEG[1] ,
    \Tile_X2Y4_WW4BEG[0] }));
 LUT4AB Tile_X1Y5_LUT4AB (.Ci(Tile_X1Y6_Co),
    .Co(Tile_X1Y5_Co),
    .UserCLK(Tile_X1Y6_UserCLKo),
    .UserCLKo(Tile_X1Y5_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X1Y5_E1BEG[3] ,
    \Tile_X1Y5_E1BEG[2] ,
    \Tile_X1Y5_E1BEG[1] ,
    \Tile_X1Y5_E1BEG[0] }),
    .E1END({\Tile_X0Y5_E1BEG[3] ,
    \Tile_X0Y5_E1BEG[2] ,
    \Tile_X0Y5_E1BEG[1] ,
    \Tile_X0Y5_E1BEG[0] }),
    .E2BEG({\Tile_X1Y5_E2BEG[7] ,
    \Tile_X1Y5_E2BEG[6] ,
    \Tile_X1Y5_E2BEG[5] ,
    \Tile_X1Y5_E2BEG[4] ,
    \Tile_X1Y5_E2BEG[3] ,
    \Tile_X1Y5_E2BEG[2] ,
    \Tile_X1Y5_E2BEG[1] ,
    \Tile_X1Y5_E2BEG[0] }),
    .E2BEGb({\Tile_X1Y5_E2BEGb[7] ,
    \Tile_X1Y5_E2BEGb[6] ,
    \Tile_X1Y5_E2BEGb[5] ,
    \Tile_X1Y5_E2BEGb[4] ,
    \Tile_X1Y5_E2BEGb[3] ,
    \Tile_X1Y5_E2BEGb[2] ,
    \Tile_X1Y5_E2BEGb[1] ,
    \Tile_X1Y5_E2BEGb[0] }),
    .E2END({\Tile_X0Y5_E2BEGb[7] ,
    \Tile_X0Y5_E2BEGb[6] ,
    \Tile_X0Y5_E2BEGb[5] ,
    \Tile_X0Y5_E2BEGb[4] ,
    \Tile_X0Y5_E2BEGb[3] ,
    \Tile_X0Y5_E2BEGb[2] ,
    \Tile_X0Y5_E2BEGb[1] ,
    \Tile_X0Y5_E2BEGb[0] }),
    .E2MID({\Tile_X0Y5_E2BEG[7] ,
    \Tile_X0Y5_E2BEG[6] ,
    \Tile_X0Y5_E2BEG[5] ,
    \Tile_X0Y5_E2BEG[4] ,
    \Tile_X0Y5_E2BEG[3] ,
    \Tile_X0Y5_E2BEG[2] ,
    \Tile_X0Y5_E2BEG[1] ,
    \Tile_X0Y5_E2BEG[0] }),
    .E6BEG({\Tile_X1Y5_E6BEG[11] ,
    \Tile_X1Y5_E6BEG[10] ,
    \Tile_X1Y5_E6BEG[9] ,
    \Tile_X1Y5_E6BEG[8] ,
    \Tile_X1Y5_E6BEG[7] ,
    \Tile_X1Y5_E6BEG[6] ,
    \Tile_X1Y5_E6BEG[5] ,
    \Tile_X1Y5_E6BEG[4] ,
    \Tile_X1Y5_E6BEG[3] ,
    \Tile_X1Y5_E6BEG[2] ,
    \Tile_X1Y5_E6BEG[1] ,
    \Tile_X1Y5_E6BEG[0] }),
    .E6END({\Tile_X0Y5_E6BEG[11] ,
    \Tile_X0Y5_E6BEG[10] ,
    \Tile_X0Y5_E6BEG[9] ,
    \Tile_X0Y5_E6BEG[8] ,
    \Tile_X0Y5_E6BEG[7] ,
    \Tile_X0Y5_E6BEG[6] ,
    \Tile_X0Y5_E6BEG[5] ,
    \Tile_X0Y5_E6BEG[4] ,
    \Tile_X0Y5_E6BEG[3] ,
    \Tile_X0Y5_E6BEG[2] ,
    \Tile_X0Y5_E6BEG[1] ,
    \Tile_X0Y5_E6BEG[0] }),
    .EE4BEG({\Tile_X1Y5_EE4BEG[15] ,
    \Tile_X1Y5_EE4BEG[14] ,
    \Tile_X1Y5_EE4BEG[13] ,
    \Tile_X1Y5_EE4BEG[12] ,
    \Tile_X1Y5_EE4BEG[11] ,
    \Tile_X1Y5_EE4BEG[10] ,
    \Tile_X1Y5_EE4BEG[9] ,
    \Tile_X1Y5_EE4BEG[8] ,
    \Tile_X1Y5_EE4BEG[7] ,
    \Tile_X1Y5_EE4BEG[6] ,
    \Tile_X1Y5_EE4BEG[5] ,
    \Tile_X1Y5_EE4BEG[4] ,
    \Tile_X1Y5_EE4BEG[3] ,
    \Tile_X1Y5_EE4BEG[2] ,
    \Tile_X1Y5_EE4BEG[1] ,
    \Tile_X1Y5_EE4BEG[0] }),
    .EE4END({\Tile_X0Y5_EE4BEG[15] ,
    \Tile_X0Y5_EE4BEG[14] ,
    \Tile_X0Y5_EE4BEG[13] ,
    \Tile_X0Y5_EE4BEG[12] ,
    \Tile_X0Y5_EE4BEG[11] ,
    \Tile_X0Y5_EE4BEG[10] ,
    \Tile_X0Y5_EE4BEG[9] ,
    \Tile_X0Y5_EE4BEG[8] ,
    \Tile_X0Y5_EE4BEG[7] ,
    \Tile_X0Y5_EE4BEG[6] ,
    \Tile_X0Y5_EE4BEG[5] ,
    \Tile_X0Y5_EE4BEG[4] ,
    \Tile_X0Y5_EE4BEG[3] ,
    \Tile_X0Y5_EE4BEG[2] ,
    \Tile_X0Y5_EE4BEG[1] ,
    \Tile_X0Y5_EE4BEG[0] }),
    .FrameData({\Tile_X0Y5_FrameData_O[31] ,
    \Tile_X0Y5_FrameData_O[30] ,
    \Tile_X0Y5_FrameData_O[29] ,
    \Tile_X0Y5_FrameData_O[28] ,
    \Tile_X0Y5_FrameData_O[27] ,
    \Tile_X0Y5_FrameData_O[26] ,
    \Tile_X0Y5_FrameData_O[25] ,
    \Tile_X0Y5_FrameData_O[24] ,
    \Tile_X0Y5_FrameData_O[23] ,
    \Tile_X0Y5_FrameData_O[22] ,
    \Tile_X0Y5_FrameData_O[21] ,
    \Tile_X0Y5_FrameData_O[20] ,
    \Tile_X0Y5_FrameData_O[19] ,
    \Tile_X0Y5_FrameData_O[18] ,
    \Tile_X0Y5_FrameData_O[17] ,
    \Tile_X0Y5_FrameData_O[16] ,
    \Tile_X0Y5_FrameData_O[15] ,
    \Tile_X0Y5_FrameData_O[14] ,
    \Tile_X0Y5_FrameData_O[13] ,
    \Tile_X0Y5_FrameData_O[12] ,
    \Tile_X0Y5_FrameData_O[11] ,
    \Tile_X0Y5_FrameData_O[10] ,
    \Tile_X0Y5_FrameData_O[9] ,
    \Tile_X0Y5_FrameData_O[8] ,
    \Tile_X0Y5_FrameData_O[7] ,
    \Tile_X0Y5_FrameData_O[6] ,
    \Tile_X0Y5_FrameData_O[5] ,
    \Tile_X0Y5_FrameData_O[4] ,
    \Tile_X0Y5_FrameData_O[3] ,
    \Tile_X0Y5_FrameData_O[2] ,
    \Tile_X0Y5_FrameData_O[1] ,
    \Tile_X0Y5_FrameData_O[0] }),
    .FrameData_O({\Tile_X1Y5_FrameData_O[31] ,
    \Tile_X1Y5_FrameData_O[30] ,
    \Tile_X1Y5_FrameData_O[29] ,
    \Tile_X1Y5_FrameData_O[28] ,
    \Tile_X1Y5_FrameData_O[27] ,
    \Tile_X1Y5_FrameData_O[26] ,
    \Tile_X1Y5_FrameData_O[25] ,
    \Tile_X1Y5_FrameData_O[24] ,
    \Tile_X1Y5_FrameData_O[23] ,
    \Tile_X1Y5_FrameData_O[22] ,
    \Tile_X1Y5_FrameData_O[21] ,
    \Tile_X1Y5_FrameData_O[20] ,
    \Tile_X1Y5_FrameData_O[19] ,
    \Tile_X1Y5_FrameData_O[18] ,
    \Tile_X1Y5_FrameData_O[17] ,
    \Tile_X1Y5_FrameData_O[16] ,
    \Tile_X1Y5_FrameData_O[15] ,
    \Tile_X1Y5_FrameData_O[14] ,
    \Tile_X1Y5_FrameData_O[13] ,
    \Tile_X1Y5_FrameData_O[12] ,
    \Tile_X1Y5_FrameData_O[11] ,
    \Tile_X1Y5_FrameData_O[10] ,
    \Tile_X1Y5_FrameData_O[9] ,
    \Tile_X1Y5_FrameData_O[8] ,
    \Tile_X1Y5_FrameData_O[7] ,
    \Tile_X1Y5_FrameData_O[6] ,
    \Tile_X1Y5_FrameData_O[5] ,
    \Tile_X1Y5_FrameData_O[4] ,
    \Tile_X1Y5_FrameData_O[3] ,
    \Tile_X1Y5_FrameData_O[2] ,
    \Tile_X1Y5_FrameData_O[1] ,
    \Tile_X1Y5_FrameData_O[0] }),
    .FrameStrobe({\Tile_X1Y6_FrameStrobe_O[19] ,
    \Tile_X1Y6_FrameStrobe_O[18] ,
    \Tile_X1Y6_FrameStrobe_O[17] ,
    \Tile_X1Y6_FrameStrobe_O[16] ,
    \Tile_X1Y6_FrameStrobe_O[15] ,
    \Tile_X1Y6_FrameStrobe_O[14] ,
    \Tile_X1Y6_FrameStrobe_O[13] ,
    \Tile_X1Y6_FrameStrobe_O[12] ,
    \Tile_X1Y6_FrameStrobe_O[11] ,
    \Tile_X1Y6_FrameStrobe_O[10] ,
    \Tile_X1Y6_FrameStrobe_O[9] ,
    \Tile_X1Y6_FrameStrobe_O[8] ,
    \Tile_X1Y6_FrameStrobe_O[7] ,
    \Tile_X1Y6_FrameStrobe_O[6] ,
    \Tile_X1Y6_FrameStrobe_O[5] ,
    \Tile_X1Y6_FrameStrobe_O[4] ,
    \Tile_X1Y6_FrameStrobe_O[3] ,
    \Tile_X1Y6_FrameStrobe_O[2] ,
    \Tile_X1Y6_FrameStrobe_O[1] ,
    \Tile_X1Y6_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X1Y5_FrameStrobe_O[19] ,
    \Tile_X1Y5_FrameStrobe_O[18] ,
    \Tile_X1Y5_FrameStrobe_O[17] ,
    \Tile_X1Y5_FrameStrobe_O[16] ,
    \Tile_X1Y5_FrameStrobe_O[15] ,
    \Tile_X1Y5_FrameStrobe_O[14] ,
    \Tile_X1Y5_FrameStrobe_O[13] ,
    \Tile_X1Y5_FrameStrobe_O[12] ,
    \Tile_X1Y5_FrameStrobe_O[11] ,
    \Tile_X1Y5_FrameStrobe_O[10] ,
    \Tile_X1Y5_FrameStrobe_O[9] ,
    \Tile_X1Y5_FrameStrobe_O[8] ,
    \Tile_X1Y5_FrameStrobe_O[7] ,
    \Tile_X1Y5_FrameStrobe_O[6] ,
    \Tile_X1Y5_FrameStrobe_O[5] ,
    \Tile_X1Y5_FrameStrobe_O[4] ,
    \Tile_X1Y5_FrameStrobe_O[3] ,
    \Tile_X1Y5_FrameStrobe_O[2] ,
    \Tile_X1Y5_FrameStrobe_O[1] ,
    \Tile_X1Y5_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X1Y5_N1BEG[3] ,
    \Tile_X1Y5_N1BEG[2] ,
    \Tile_X1Y5_N1BEG[1] ,
    \Tile_X1Y5_N1BEG[0] }),
    .N1END({\Tile_X1Y6_N1BEG[3] ,
    \Tile_X1Y6_N1BEG[2] ,
    \Tile_X1Y6_N1BEG[1] ,
    \Tile_X1Y6_N1BEG[0] }),
    .N2BEG({\Tile_X1Y5_N2BEG[7] ,
    \Tile_X1Y5_N2BEG[6] ,
    \Tile_X1Y5_N2BEG[5] ,
    \Tile_X1Y5_N2BEG[4] ,
    \Tile_X1Y5_N2BEG[3] ,
    \Tile_X1Y5_N2BEG[2] ,
    \Tile_X1Y5_N2BEG[1] ,
    \Tile_X1Y5_N2BEG[0] }),
    .N2BEGb({\Tile_X1Y5_N2BEGb[7] ,
    \Tile_X1Y5_N2BEGb[6] ,
    \Tile_X1Y5_N2BEGb[5] ,
    \Tile_X1Y5_N2BEGb[4] ,
    \Tile_X1Y5_N2BEGb[3] ,
    \Tile_X1Y5_N2BEGb[2] ,
    \Tile_X1Y5_N2BEGb[1] ,
    \Tile_X1Y5_N2BEGb[0] }),
    .N2END({\Tile_X1Y6_N2BEGb[7] ,
    \Tile_X1Y6_N2BEGb[6] ,
    \Tile_X1Y6_N2BEGb[5] ,
    \Tile_X1Y6_N2BEGb[4] ,
    \Tile_X1Y6_N2BEGb[3] ,
    \Tile_X1Y6_N2BEGb[2] ,
    \Tile_X1Y6_N2BEGb[1] ,
    \Tile_X1Y6_N2BEGb[0] }),
    .N2MID({\Tile_X1Y6_N2BEG[7] ,
    \Tile_X1Y6_N2BEG[6] ,
    \Tile_X1Y6_N2BEG[5] ,
    \Tile_X1Y6_N2BEG[4] ,
    \Tile_X1Y6_N2BEG[3] ,
    \Tile_X1Y6_N2BEG[2] ,
    \Tile_X1Y6_N2BEG[1] ,
    \Tile_X1Y6_N2BEG[0] }),
    .N4BEG({\Tile_X1Y5_N4BEG[15] ,
    \Tile_X1Y5_N4BEG[14] ,
    \Tile_X1Y5_N4BEG[13] ,
    \Tile_X1Y5_N4BEG[12] ,
    \Tile_X1Y5_N4BEG[11] ,
    \Tile_X1Y5_N4BEG[10] ,
    \Tile_X1Y5_N4BEG[9] ,
    \Tile_X1Y5_N4BEG[8] ,
    \Tile_X1Y5_N4BEG[7] ,
    \Tile_X1Y5_N4BEG[6] ,
    \Tile_X1Y5_N4BEG[5] ,
    \Tile_X1Y5_N4BEG[4] ,
    \Tile_X1Y5_N4BEG[3] ,
    \Tile_X1Y5_N4BEG[2] ,
    \Tile_X1Y5_N4BEG[1] ,
    \Tile_X1Y5_N4BEG[0] }),
    .N4END({\Tile_X1Y6_N4BEG[15] ,
    \Tile_X1Y6_N4BEG[14] ,
    \Tile_X1Y6_N4BEG[13] ,
    \Tile_X1Y6_N4BEG[12] ,
    \Tile_X1Y6_N4BEG[11] ,
    \Tile_X1Y6_N4BEG[10] ,
    \Tile_X1Y6_N4BEG[9] ,
    \Tile_X1Y6_N4BEG[8] ,
    \Tile_X1Y6_N4BEG[7] ,
    \Tile_X1Y6_N4BEG[6] ,
    \Tile_X1Y6_N4BEG[5] ,
    \Tile_X1Y6_N4BEG[4] ,
    \Tile_X1Y6_N4BEG[3] ,
    \Tile_X1Y6_N4BEG[2] ,
    \Tile_X1Y6_N4BEG[1] ,
    \Tile_X1Y6_N4BEG[0] }),
    .NN4BEG({\Tile_X1Y5_NN4BEG[15] ,
    \Tile_X1Y5_NN4BEG[14] ,
    \Tile_X1Y5_NN4BEG[13] ,
    \Tile_X1Y5_NN4BEG[12] ,
    \Tile_X1Y5_NN4BEG[11] ,
    \Tile_X1Y5_NN4BEG[10] ,
    \Tile_X1Y5_NN4BEG[9] ,
    \Tile_X1Y5_NN4BEG[8] ,
    \Tile_X1Y5_NN4BEG[7] ,
    \Tile_X1Y5_NN4BEG[6] ,
    \Tile_X1Y5_NN4BEG[5] ,
    \Tile_X1Y5_NN4BEG[4] ,
    \Tile_X1Y5_NN4BEG[3] ,
    \Tile_X1Y5_NN4BEG[2] ,
    \Tile_X1Y5_NN4BEG[1] ,
    \Tile_X1Y5_NN4BEG[0] }),
    .NN4END({\Tile_X1Y6_NN4BEG[15] ,
    \Tile_X1Y6_NN4BEG[14] ,
    \Tile_X1Y6_NN4BEG[13] ,
    \Tile_X1Y6_NN4BEG[12] ,
    \Tile_X1Y6_NN4BEG[11] ,
    \Tile_X1Y6_NN4BEG[10] ,
    \Tile_X1Y6_NN4BEG[9] ,
    \Tile_X1Y6_NN4BEG[8] ,
    \Tile_X1Y6_NN4BEG[7] ,
    \Tile_X1Y6_NN4BEG[6] ,
    \Tile_X1Y6_NN4BEG[5] ,
    \Tile_X1Y6_NN4BEG[4] ,
    \Tile_X1Y6_NN4BEG[3] ,
    \Tile_X1Y6_NN4BEG[2] ,
    \Tile_X1Y6_NN4BEG[1] ,
    \Tile_X1Y6_NN4BEG[0] }),
    .S1BEG({\Tile_X1Y5_S1BEG[3] ,
    \Tile_X1Y5_S1BEG[2] ,
    \Tile_X1Y5_S1BEG[1] ,
    \Tile_X1Y5_S1BEG[0] }),
    .S1END({\Tile_X1Y4_S1BEG[3] ,
    \Tile_X1Y4_S1BEG[2] ,
    \Tile_X1Y4_S1BEG[1] ,
    \Tile_X1Y4_S1BEG[0] }),
    .S2BEG({\Tile_X1Y5_S2BEG[7] ,
    \Tile_X1Y5_S2BEG[6] ,
    \Tile_X1Y5_S2BEG[5] ,
    \Tile_X1Y5_S2BEG[4] ,
    \Tile_X1Y5_S2BEG[3] ,
    \Tile_X1Y5_S2BEG[2] ,
    \Tile_X1Y5_S2BEG[1] ,
    \Tile_X1Y5_S2BEG[0] }),
    .S2BEGb({\Tile_X1Y5_S2BEGb[7] ,
    \Tile_X1Y5_S2BEGb[6] ,
    \Tile_X1Y5_S2BEGb[5] ,
    \Tile_X1Y5_S2BEGb[4] ,
    \Tile_X1Y5_S2BEGb[3] ,
    \Tile_X1Y5_S2BEGb[2] ,
    \Tile_X1Y5_S2BEGb[1] ,
    \Tile_X1Y5_S2BEGb[0] }),
    .S2END({\Tile_X1Y4_S2BEGb[7] ,
    \Tile_X1Y4_S2BEGb[6] ,
    \Tile_X1Y4_S2BEGb[5] ,
    \Tile_X1Y4_S2BEGb[4] ,
    \Tile_X1Y4_S2BEGb[3] ,
    \Tile_X1Y4_S2BEGb[2] ,
    \Tile_X1Y4_S2BEGb[1] ,
    \Tile_X1Y4_S2BEGb[0] }),
    .S2MID({\Tile_X1Y4_S2BEG[7] ,
    \Tile_X1Y4_S2BEG[6] ,
    \Tile_X1Y4_S2BEG[5] ,
    \Tile_X1Y4_S2BEG[4] ,
    \Tile_X1Y4_S2BEG[3] ,
    \Tile_X1Y4_S2BEG[2] ,
    \Tile_X1Y4_S2BEG[1] ,
    \Tile_X1Y4_S2BEG[0] }),
    .S4BEG({\Tile_X1Y5_S4BEG[15] ,
    \Tile_X1Y5_S4BEG[14] ,
    \Tile_X1Y5_S4BEG[13] ,
    \Tile_X1Y5_S4BEG[12] ,
    \Tile_X1Y5_S4BEG[11] ,
    \Tile_X1Y5_S4BEG[10] ,
    \Tile_X1Y5_S4BEG[9] ,
    \Tile_X1Y5_S4BEG[8] ,
    \Tile_X1Y5_S4BEG[7] ,
    \Tile_X1Y5_S4BEG[6] ,
    \Tile_X1Y5_S4BEG[5] ,
    \Tile_X1Y5_S4BEG[4] ,
    \Tile_X1Y5_S4BEG[3] ,
    \Tile_X1Y5_S4BEG[2] ,
    \Tile_X1Y5_S4BEG[1] ,
    \Tile_X1Y5_S4BEG[0] }),
    .S4END({\Tile_X1Y4_S4BEG[15] ,
    \Tile_X1Y4_S4BEG[14] ,
    \Tile_X1Y4_S4BEG[13] ,
    \Tile_X1Y4_S4BEG[12] ,
    \Tile_X1Y4_S4BEG[11] ,
    \Tile_X1Y4_S4BEG[10] ,
    \Tile_X1Y4_S4BEG[9] ,
    \Tile_X1Y4_S4BEG[8] ,
    \Tile_X1Y4_S4BEG[7] ,
    \Tile_X1Y4_S4BEG[6] ,
    \Tile_X1Y4_S4BEG[5] ,
    \Tile_X1Y4_S4BEG[4] ,
    \Tile_X1Y4_S4BEG[3] ,
    \Tile_X1Y4_S4BEG[2] ,
    \Tile_X1Y4_S4BEG[1] ,
    \Tile_X1Y4_S4BEG[0] }),
    .SS4BEG({\Tile_X1Y5_SS4BEG[15] ,
    \Tile_X1Y5_SS4BEG[14] ,
    \Tile_X1Y5_SS4BEG[13] ,
    \Tile_X1Y5_SS4BEG[12] ,
    \Tile_X1Y5_SS4BEG[11] ,
    \Tile_X1Y5_SS4BEG[10] ,
    \Tile_X1Y5_SS4BEG[9] ,
    \Tile_X1Y5_SS4BEG[8] ,
    \Tile_X1Y5_SS4BEG[7] ,
    \Tile_X1Y5_SS4BEG[6] ,
    \Tile_X1Y5_SS4BEG[5] ,
    \Tile_X1Y5_SS4BEG[4] ,
    \Tile_X1Y5_SS4BEG[3] ,
    \Tile_X1Y5_SS4BEG[2] ,
    \Tile_X1Y5_SS4BEG[1] ,
    \Tile_X1Y5_SS4BEG[0] }),
    .SS4END({\Tile_X1Y4_SS4BEG[15] ,
    \Tile_X1Y4_SS4BEG[14] ,
    \Tile_X1Y4_SS4BEG[13] ,
    \Tile_X1Y4_SS4BEG[12] ,
    \Tile_X1Y4_SS4BEG[11] ,
    \Tile_X1Y4_SS4BEG[10] ,
    \Tile_X1Y4_SS4BEG[9] ,
    \Tile_X1Y4_SS4BEG[8] ,
    \Tile_X1Y4_SS4BEG[7] ,
    \Tile_X1Y4_SS4BEG[6] ,
    \Tile_X1Y4_SS4BEG[5] ,
    \Tile_X1Y4_SS4BEG[4] ,
    \Tile_X1Y4_SS4BEG[3] ,
    \Tile_X1Y4_SS4BEG[2] ,
    \Tile_X1Y4_SS4BEG[1] ,
    \Tile_X1Y4_SS4BEG[0] }),
    .W1BEG({\Tile_X1Y5_W1BEG[3] ,
    \Tile_X1Y5_W1BEG[2] ,
    \Tile_X1Y5_W1BEG[1] ,
    \Tile_X1Y5_W1BEG[0] }),
    .W1END({\Tile_X2Y5_W1BEG[3] ,
    \Tile_X2Y5_W1BEG[2] ,
    \Tile_X2Y5_W1BEG[1] ,
    \Tile_X2Y5_W1BEG[0] }),
    .W2BEG({\Tile_X1Y5_W2BEG[7] ,
    \Tile_X1Y5_W2BEG[6] ,
    \Tile_X1Y5_W2BEG[5] ,
    \Tile_X1Y5_W2BEG[4] ,
    \Tile_X1Y5_W2BEG[3] ,
    \Tile_X1Y5_W2BEG[2] ,
    \Tile_X1Y5_W2BEG[1] ,
    \Tile_X1Y5_W2BEG[0] }),
    .W2BEGb({\Tile_X1Y5_W2BEGb[7] ,
    \Tile_X1Y5_W2BEGb[6] ,
    \Tile_X1Y5_W2BEGb[5] ,
    \Tile_X1Y5_W2BEGb[4] ,
    \Tile_X1Y5_W2BEGb[3] ,
    \Tile_X1Y5_W2BEGb[2] ,
    \Tile_X1Y5_W2BEGb[1] ,
    \Tile_X1Y5_W2BEGb[0] }),
    .W2END({\Tile_X2Y5_W2BEGb[7] ,
    \Tile_X2Y5_W2BEGb[6] ,
    \Tile_X2Y5_W2BEGb[5] ,
    \Tile_X2Y5_W2BEGb[4] ,
    \Tile_X2Y5_W2BEGb[3] ,
    \Tile_X2Y5_W2BEGb[2] ,
    \Tile_X2Y5_W2BEGb[1] ,
    \Tile_X2Y5_W2BEGb[0] }),
    .W2MID({\Tile_X2Y5_W2BEG[7] ,
    \Tile_X2Y5_W2BEG[6] ,
    \Tile_X2Y5_W2BEG[5] ,
    \Tile_X2Y5_W2BEG[4] ,
    \Tile_X2Y5_W2BEG[3] ,
    \Tile_X2Y5_W2BEG[2] ,
    \Tile_X2Y5_W2BEG[1] ,
    \Tile_X2Y5_W2BEG[0] }),
    .W6BEG({\Tile_X1Y5_W6BEG[11] ,
    \Tile_X1Y5_W6BEG[10] ,
    \Tile_X1Y5_W6BEG[9] ,
    \Tile_X1Y5_W6BEG[8] ,
    \Tile_X1Y5_W6BEG[7] ,
    \Tile_X1Y5_W6BEG[6] ,
    \Tile_X1Y5_W6BEG[5] ,
    \Tile_X1Y5_W6BEG[4] ,
    \Tile_X1Y5_W6BEG[3] ,
    \Tile_X1Y5_W6BEG[2] ,
    \Tile_X1Y5_W6BEG[1] ,
    \Tile_X1Y5_W6BEG[0] }),
    .W6END({\Tile_X2Y5_W6BEG[11] ,
    \Tile_X2Y5_W6BEG[10] ,
    \Tile_X2Y5_W6BEG[9] ,
    \Tile_X2Y5_W6BEG[8] ,
    \Tile_X2Y5_W6BEG[7] ,
    \Tile_X2Y5_W6BEG[6] ,
    \Tile_X2Y5_W6BEG[5] ,
    \Tile_X2Y5_W6BEG[4] ,
    \Tile_X2Y5_W6BEG[3] ,
    \Tile_X2Y5_W6BEG[2] ,
    \Tile_X2Y5_W6BEG[1] ,
    \Tile_X2Y5_W6BEG[0] }),
    .WW4BEG({\Tile_X1Y5_WW4BEG[15] ,
    \Tile_X1Y5_WW4BEG[14] ,
    \Tile_X1Y5_WW4BEG[13] ,
    \Tile_X1Y5_WW4BEG[12] ,
    \Tile_X1Y5_WW4BEG[11] ,
    \Tile_X1Y5_WW4BEG[10] ,
    \Tile_X1Y5_WW4BEG[9] ,
    \Tile_X1Y5_WW4BEG[8] ,
    \Tile_X1Y5_WW4BEG[7] ,
    \Tile_X1Y5_WW4BEG[6] ,
    \Tile_X1Y5_WW4BEG[5] ,
    \Tile_X1Y5_WW4BEG[4] ,
    \Tile_X1Y5_WW4BEG[3] ,
    \Tile_X1Y5_WW4BEG[2] ,
    \Tile_X1Y5_WW4BEG[1] ,
    \Tile_X1Y5_WW4BEG[0] }),
    .WW4END({\Tile_X2Y5_WW4BEG[15] ,
    \Tile_X2Y5_WW4BEG[14] ,
    \Tile_X2Y5_WW4BEG[13] ,
    \Tile_X2Y5_WW4BEG[12] ,
    \Tile_X2Y5_WW4BEG[11] ,
    \Tile_X2Y5_WW4BEG[10] ,
    \Tile_X2Y5_WW4BEG[9] ,
    \Tile_X2Y5_WW4BEG[8] ,
    \Tile_X2Y5_WW4BEG[7] ,
    \Tile_X2Y5_WW4BEG[6] ,
    \Tile_X2Y5_WW4BEG[5] ,
    \Tile_X2Y5_WW4BEG[4] ,
    \Tile_X2Y5_WW4BEG[3] ,
    \Tile_X2Y5_WW4BEG[2] ,
    \Tile_X2Y5_WW4BEG[1] ,
    \Tile_X2Y5_WW4BEG[0] }));
 LUT4AB Tile_X1Y6_LUT4AB (.Ci(Tile_X1Y7_Co),
    .Co(Tile_X1Y6_Co),
    .UserCLK(Tile_X1Y7_UserCLKo),
    .UserCLKo(Tile_X1Y6_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X1Y6_E1BEG[3] ,
    \Tile_X1Y6_E1BEG[2] ,
    \Tile_X1Y6_E1BEG[1] ,
    \Tile_X1Y6_E1BEG[0] }),
    .E1END({\Tile_X0Y6_E1BEG[3] ,
    \Tile_X0Y6_E1BEG[2] ,
    \Tile_X0Y6_E1BEG[1] ,
    \Tile_X0Y6_E1BEG[0] }),
    .E2BEG({\Tile_X1Y6_E2BEG[7] ,
    \Tile_X1Y6_E2BEG[6] ,
    \Tile_X1Y6_E2BEG[5] ,
    \Tile_X1Y6_E2BEG[4] ,
    \Tile_X1Y6_E2BEG[3] ,
    \Tile_X1Y6_E2BEG[2] ,
    \Tile_X1Y6_E2BEG[1] ,
    \Tile_X1Y6_E2BEG[0] }),
    .E2BEGb({\Tile_X1Y6_E2BEGb[7] ,
    \Tile_X1Y6_E2BEGb[6] ,
    \Tile_X1Y6_E2BEGb[5] ,
    \Tile_X1Y6_E2BEGb[4] ,
    \Tile_X1Y6_E2BEGb[3] ,
    \Tile_X1Y6_E2BEGb[2] ,
    \Tile_X1Y6_E2BEGb[1] ,
    \Tile_X1Y6_E2BEGb[0] }),
    .E2END({\Tile_X0Y6_E2BEGb[7] ,
    \Tile_X0Y6_E2BEGb[6] ,
    \Tile_X0Y6_E2BEGb[5] ,
    \Tile_X0Y6_E2BEGb[4] ,
    \Tile_X0Y6_E2BEGb[3] ,
    \Tile_X0Y6_E2BEGb[2] ,
    \Tile_X0Y6_E2BEGb[1] ,
    \Tile_X0Y6_E2BEGb[0] }),
    .E2MID({\Tile_X0Y6_E2BEG[7] ,
    \Tile_X0Y6_E2BEG[6] ,
    \Tile_X0Y6_E2BEG[5] ,
    \Tile_X0Y6_E2BEG[4] ,
    \Tile_X0Y6_E2BEG[3] ,
    \Tile_X0Y6_E2BEG[2] ,
    \Tile_X0Y6_E2BEG[1] ,
    \Tile_X0Y6_E2BEG[0] }),
    .E6BEG({\Tile_X1Y6_E6BEG[11] ,
    \Tile_X1Y6_E6BEG[10] ,
    \Tile_X1Y6_E6BEG[9] ,
    \Tile_X1Y6_E6BEG[8] ,
    \Tile_X1Y6_E6BEG[7] ,
    \Tile_X1Y6_E6BEG[6] ,
    \Tile_X1Y6_E6BEG[5] ,
    \Tile_X1Y6_E6BEG[4] ,
    \Tile_X1Y6_E6BEG[3] ,
    \Tile_X1Y6_E6BEG[2] ,
    \Tile_X1Y6_E6BEG[1] ,
    \Tile_X1Y6_E6BEG[0] }),
    .E6END({\Tile_X0Y6_E6BEG[11] ,
    \Tile_X0Y6_E6BEG[10] ,
    \Tile_X0Y6_E6BEG[9] ,
    \Tile_X0Y6_E6BEG[8] ,
    \Tile_X0Y6_E6BEG[7] ,
    \Tile_X0Y6_E6BEG[6] ,
    \Tile_X0Y6_E6BEG[5] ,
    \Tile_X0Y6_E6BEG[4] ,
    \Tile_X0Y6_E6BEG[3] ,
    \Tile_X0Y6_E6BEG[2] ,
    \Tile_X0Y6_E6BEG[1] ,
    \Tile_X0Y6_E6BEG[0] }),
    .EE4BEG({\Tile_X1Y6_EE4BEG[15] ,
    \Tile_X1Y6_EE4BEG[14] ,
    \Tile_X1Y6_EE4BEG[13] ,
    \Tile_X1Y6_EE4BEG[12] ,
    \Tile_X1Y6_EE4BEG[11] ,
    \Tile_X1Y6_EE4BEG[10] ,
    \Tile_X1Y6_EE4BEG[9] ,
    \Tile_X1Y6_EE4BEG[8] ,
    \Tile_X1Y6_EE4BEG[7] ,
    \Tile_X1Y6_EE4BEG[6] ,
    \Tile_X1Y6_EE4BEG[5] ,
    \Tile_X1Y6_EE4BEG[4] ,
    \Tile_X1Y6_EE4BEG[3] ,
    \Tile_X1Y6_EE4BEG[2] ,
    \Tile_X1Y6_EE4BEG[1] ,
    \Tile_X1Y6_EE4BEG[0] }),
    .EE4END({\Tile_X0Y6_EE4BEG[15] ,
    \Tile_X0Y6_EE4BEG[14] ,
    \Tile_X0Y6_EE4BEG[13] ,
    \Tile_X0Y6_EE4BEG[12] ,
    \Tile_X0Y6_EE4BEG[11] ,
    \Tile_X0Y6_EE4BEG[10] ,
    \Tile_X0Y6_EE4BEG[9] ,
    \Tile_X0Y6_EE4BEG[8] ,
    \Tile_X0Y6_EE4BEG[7] ,
    \Tile_X0Y6_EE4BEG[6] ,
    \Tile_X0Y6_EE4BEG[5] ,
    \Tile_X0Y6_EE4BEG[4] ,
    \Tile_X0Y6_EE4BEG[3] ,
    \Tile_X0Y6_EE4BEG[2] ,
    \Tile_X0Y6_EE4BEG[1] ,
    \Tile_X0Y6_EE4BEG[0] }),
    .FrameData({\Tile_X0Y6_FrameData_O[31] ,
    \Tile_X0Y6_FrameData_O[30] ,
    \Tile_X0Y6_FrameData_O[29] ,
    \Tile_X0Y6_FrameData_O[28] ,
    \Tile_X0Y6_FrameData_O[27] ,
    \Tile_X0Y6_FrameData_O[26] ,
    \Tile_X0Y6_FrameData_O[25] ,
    \Tile_X0Y6_FrameData_O[24] ,
    \Tile_X0Y6_FrameData_O[23] ,
    \Tile_X0Y6_FrameData_O[22] ,
    \Tile_X0Y6_FrameData_O[21] ,
    \Tile_X0Y6_FrameData_O[20] ,
    \Tile_X0Y6_FrameData_O[19] ,
    \Tile_X0Y6_FrameData_O[18] ,
    \Tile_X0Y6_FrameData_O[17] ,
    \Tile_X0Y6_FrameData_O[16] ,
    \Tile_X0Y6_FrameData_O[15] ,
    \Tile_X0Y6_FrameData_O[14] ,
    \Tile_X0Y6_FrameData_O[13] ,
    \Tile_X0Y6_FrameData_O[12] ,
    \Tile_X0Y6_FrameData_O[11] ,
    \Tile_X0Y6_FrameData_O[10] ,
    \Tile_X0Y6_FrameData_O[9] ,
    \Tile_X0Y6_FrameData_O[8] ,
    \Tile_X0Y6_FrameData_O[7] ,
    \Tile_X0Y6_FrameData_O[6] ,
    \Tile_X0Y6_FrameData_O[5] ,
    \Tile_X0Y6_FrameData_O[4] ,
    \Tile_X0Y6_FrameData_O[3] ,
    \Tile_X0Y6_FrameData_O[2] ,
    \Tile_X0Y6_FrameData_O[1] ,
    \Tile_X0Y6_FrameData_O[0] }),
    .FrameData_O({\Tile_X1Y6_FrameData_O[31] ,
    \Tile_X1Y6_FrameData_O[30] ,
    \Tile_X1Y6_FrameData_O[29] ,
    \Tile_X1Y6_FrameData_O[28] ,
    \Tile_X1Y6_FrameData_O[27] ,
    \Tile_X1Y6_FrameData_O[26] ,
    \Tile_X1Y6_FrameData_O[25] ,
    \Tile_X1Y6_FrameData_O[24] ,
    \Tile_X1Y6_FrameData_O[23] ,
    \Tile_X1Y6_FrameData_O[22] ,
    \Tile_X1Y6_FrameData_O[21] ,
    \Tile_X1Y6_FrameData_O[20] ,
    \Tile_X1Y6_FrameData_O[19] ,
    \Tile_X1Y6_FrameData_O[18] ,
    \Tile_X1Y6_FrameData_O[17] ,
    \Tile_X1Y6_FrameData_O[16] ,
    \Tile_X1Y6_FrameData_O[15] ,
    \Tile_X1Y6_FrameData_O[14] ,
    \Tile_X1Y6_FrameData_O[13] ,
    \Tile_X1Y6_FrameData_O[12] ,
    \Tile_X1Y6_FrameData_O[11] ,
    \Tile_X1Y6_FrameData_O[10] ,
    \Tile_X1Y6_FrameData_O[9] ,
    \Tile_X1Y6_FrameData_O[8] ,
    \Tile_X1Y6_FrameData_O[7] ,
    \Tile_X1Y6_FrameData_O[6] ,
    \Tile_X1Y6_FrameData_O[5] ,
    \Tile_X1Y6_FrameData_O[4] ,
    \Tile_X1Y6_FrameData_O[3] ,
    \Tile_X1Y6_FrameData_O[2] ,
    \Tile_X1Y6_FrameData_O[1] ,
    \Tile_X1Y6_FrameData_O[0] }),
    .FrameStrobe({\Tile_X1Y7_FrameStrobe_O[19] ,
    \Tile_X1Y7_FrameStrobe_O[18] ,
    \Tile_X1Y7_FrameStrobe_O[17] ,
    \Tile_X1Y7_FrameStrobe_O[16] ,
    \Tile_X1Y7_FrameStrobe_O[15] ,
    \Tile_X1Y7_FrameStrobe_O[14] ,
    \Tile_X1Y7_FrameStrobe_O[13] ,
    \Tile_X1Y7_FrameStrobe_O[12] ,
    \Tile_X1Y7_FrameStrobe_O[11] ,
    \Tile_X1Y7_FrameStrobe_O[10] ,
    \Tile_X1Y7_FrameStrobe_O[9] ,
    \Tile_X1Y7_FrameStrobe_O[8] ,
    \Tile_X1Y7_FrameStrobe_O[7] ,
    \Tile_X1Y7_FrameStrobe_O[6] ,
    \Tile_X1Y7_FrameStrobe_O[5] ,
    \Tile_X1Y7_FrameStrobe_O[4] ,
    \Tile_X1Y7_FrameStrobe_O[3] ,
    \Tile_X1Y7_FrameStrobe_O[2] ,
    \Tile_X1Y7_FrameStrobe_O[1] ,
    \Tile_X1Y7_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X1Y6_FrameStrobe_O[19] ,
    \Tile_X1Y6_FrameStrobe_O[18] ,
    \Tile_X1Y6_FrameStrobe_O[17] ,
    \Tile_X1Y6_FrameStrobe_O[16] ,
    \Tile_X1Y6_FrameStrobe_O[15] ,
    \Tile_X1Y6_FrameStrobe_O[14] ,
    \Tile_X1Y6_FrameStrobe_O[13] ,
    \Tile_X1Y6_FrameStrobe_O[12] ,
    \Tile_X1Y6_FrameStrobe_O[11] ,
    \Tile_X1Y6_FrameStrobe_O[10] ,
    \Tile_X1Y6_FrameStrobe_O[9] ,
    \Tile_X1Y6_FrameStrobe_O[8] ,
    \Tile_X1Y6_FrameStrobe_O[7] ,
    \Tile_X1Y6_FrameStrobe_O[6] ,
    \Tile_X1Y6_FrameStrobe_O[5] ,
    \Tile_X1Y6_FrameStrobe_O[4] ,
    \Tile_X1Y6_FrameStrobe_O[3] ,
    \Tile_X1Y6_FrameStrobe_O[2] ,
    \Tile_X1Y6_FrameStrobe_O[1] ,
    \Tile_X1Y6_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X1Y6_N1BEG[3] ,
    \Tile_X1Y6_N1BEG[2] ,
    \Tile_X1Y6_N1BEG[1] ,
    \Tile_X1Y6_N1BEG[0] }),
    .N1END({\Tile_X1Y7_N1BEG[3] ,
    \Tile_X1Y7_N1BEG[2] ,
    \Tile_X1Y7_N1BEG[1] ,
    \Tile_X1Y7_N1BEG[0] }),
    .N2BEG({\Tile_X1Y6_N2BEG[7] ,
    \Tile_X1Y6_N2BEG[6] ,
    \Tile_X1Y6_N2BEG[5] ,
    \Tile_X1Y6_N2BEG[4] ,
    \Tile_X1Y6_N2BEG[3] ,
    \Tile_X1Y6_N2BEG[2] ,
    \Tile_X1Y6_N2BEG[1] ,
    \Tile_X1Y6_N2BEG[0] }),
    .N2BEGb({\Tile_X1Y6_N2BEGb[7] ,
    \Tile_X1Y6_N2BEGb[6] ,
    \Tile_X1Y6_N2BEGb[5] ,
    \Tile_X1Y6_N2BEGb[4] ,
    \Tile_X1Y6_N2BEGb[3] ,
    \Tile_X1Y6_N2BEGb[2] ,
    \Tile_X1Y6_N2BEGb[1] ,
    \Tile_X1Y6_N2BEGb[0] }),
    .N2END({\Tile_X1Y7_N2BEGb[7] ,
    \Tile_X1Y7_N2BEGb[6] ,
    \Tile_X1Y7_N2BEGb[5] ,
    \Tile_X1Y7_N2BEGb[4] ,
    \Tile_X1Y7_N2BEGb[3] ,
    \Tile_X1Y7_N2BEGb[2] ,
    \Tile_X1Y7_N2BEGb[1] ,
    \Tile_X1Y7_N2BEGb[0] }),
    .N2MID({\Tile_X1Y7_N2BEG[7] ,
    \Tile_X1Y7_N2BEG[6] ,
    \Tile_X1Y7_N2BEG[5] ,
    \Tile_X1Y7_N2BEG[4] ,
    \Tile_X1Y7_N2BEG[3] ,
    \Tile_X1Y7_N2BEG[2] ,
    \Tile_X1Y7_N2BEG[1] ,
    \Tile_X1Y7_N2BEG[0] }),
    .N4BEG({\Tile_X1Y6_N4BEG[15] ,
    \Tile_X1Y6_N4BEG[14] ,
    \Tile_X1Y6_N4BEG[13] ,
    \Tile_X1Y6_N4BEG[12] ,
    \Tile_X1Y6_N4BEG[11] ,
    \Tile_X1Y6_N4BEG[10] ,
    \Tile_X1Y6_N4BEG[9] ,
    \Tile_X1Y6_N4BEG[8] ,
    \Tile_X1Y6_N4BEG[7] ,
    \Tile_X1Y6_N4BEG[6] ,
    \Tile_X1Y6_N4BEG[5] ,
    \Tile_X1Y6_N4BEG[4] ,
    \Tile_X1Y6_N4BEG[3] ,
    \Tile_X1Y6_N4BEG[2] ,
    \Tile_X1Y6_N4BEG[1] ,
    \Tile_X1Y6_N4BEG[0] }),
    .N4END({\Tile_X1Y7_N4BEG[15] ,
    \Tile_X1Y7_N4BEG[14] ,
    \Tile_X1Y7_N4BEG[13] ,
    \Tile_X1Y7_N4BEG[12] ,
    \Tile_X1Y7_N4BEG[11] ,
    \Tile_X1Y7_N4BEG[10] ,
    \Tile_X1Y7_N4BEG[9] ,
    \Tile_X1Y7_N4BEG[8] ,
    \Tile_X1Y7_N4BEG[7] ,
    \Tile_X1Y7_N4BEG[6] ,
    \Tile_X1Y7_N4BEG[5] ,
    \Tile_X1Y7_N4BEG[4] ,
    \Tile_X1Y7_N4BEG[3] ,
    \Tile_X1Y7_N4BEG[2] ,
    \Tile_X1Y7_N4BEG[1] ,
    \Tile_X1Y7_N4BEG[0] }),
    .NN4BEG({\Tile_X1Y6_NN4BEG[15] ,
    \Tile_X1Y6_NN4BEG[14] ,
    \Tile_X1Y6_NN4BEG[13] ,
    \Tile_X1Y6_NN4BEG[12] ,
    \Tile_X1Y6_NN4BEG[11] ,
    \Tile_X1Y6_NN4BEG[10] ,
    \Tile_X1Y6_NN4BEG[9] ,
    \Tile_X1Y6_NN4BEG[8] ,
    \Tile_X1Y6_NN4BEG[7] ,
    \Tile_X1Y6_NN4BEG[6] ,
    \Tile_X1Y6_NN4BEG[5] ,
    \Tile_X1Y6_NN4BEG[4] ,
    \Tile_X1Y6_NN4BEG[3] ,
    \Tile_X1Y6_NN4BEG[2] ,
    \Tile_X1Y6_NN4BEG[1] ,
    \Tile_X1Y6_NN4BEG[0] }),
    .NN4END({\Tile_X1Y7_NN4BEG[15] ,
    \Tile_X1Y7_NN4BEG[14] ,
    \Tile_X1Y7_NN4BEG[13] ,
    \Tile_X1Y7_NN4BEG[12] ,
    \Tile_X1Y7_NN4BEG[11] ,
    \Tile_X1Y7_NN4BEG[10] ,
    \Tile_X1Y7_NN4BEG[9] ,
    \Tile_X1Y7_NN4BEG[8] ,
    \Tile_X1Y7_NN4BEG[7] ,
    \Tile_X1Y7_NN4BEG[6] ,
    \Tile_X1Y7_NN4BEG[5] ,
    \Tile_X1Y7_NN4BEG[4] ,
    \Tile_X1Y7_NN4BEG[3] ,
    \Tile_X1Y7_NN4BEG[2] ,
    \Tile_X1Y7_NN4BEG[1] ,
    \Tile_X1Y7_NN4BEG[0] }),
    .S1BEG({\Tile_X1Y6_S1BEG[3] ,
    \Tile_X1Y6_S1BEG[2] ,
    \Tile_X1Y6_S1BEG[1] ,
    \Tile_X1Y6_S1BEG[0] }),
    .S1END({\Tile_X1Y5_S1BEG[3] ,
    \Tile_X1Y5_S1BEG[2] ,
    \Tile_X1Y5_S1BEG[1] ,
    \Tile_X1Y5_S1BEG[0] }),
    .S2BEG({\Tile_X1Y6_S2BEG[7] ,
    \Tile_X1Y6_S2BEG[6] ,
    \Tile_X1Y6_S2BEG[5] ,
    \Tile_X1Y6_S2BEG[4] ,
    \Tile_X1Y6_S2BEG[3] ,
    \Tile_X1Y6_S2BEG[2] ,
    \Tile_X1Y6_S2BEG[1] ,
    \Tile_X1Y6_S2BEG[0] }),
    .S2BEGb({\Tile_X1Y6_S2BEGb[7] ,
    \Tile_X1Y6_S2BEGb[6] ,
    \Tile_X1Y6_S2BEGb[5] ,
    \Tile_X1Y6_S2BEGb[4] ,
    \Tile_X1Y6_S2BEGb[3] ,
    \Tile_X1Y6_S2BEGb[2] ,
    \Tile_X1Y6_S2BEGb[1] ,
    \Tile_X1Y6_S2BEGb[0] }),
    .S2END({\Tile_X1Y5_S2BEGb[7] ,
    \Tile_X1Y5_S2BEGb[6] ,
    \Tile_X1Y5_S2BEGb[5] ,
    \Tile_X1Y5_S2BEGb[4] ,
    \Tile_X1Y5_S2BEGb[3] ,
    \Tile_X1Y5_S2BEGb[2] ,
    \Tile_X1Y5_S2BEGb[1] ,
    \Tile_X1Y5_S2BEGb[0] }),
    .S2MID({\Tile_X1Y5_S2BEG[7] ,
    \Tile_X1Y5_S2BEG[6] ,
    \Tile_X1Y5_S2BEG[5] ,
    \Tile_X1Y5_S2BEG[4] ,
    \Tile_X1Y5_S2BEG[3] ,
    \Tile_X1Y5_S2BEG[2] ,
    \Tile_X1Y5_S2BEG[1] ,
    \Tile_X1Y5_S2BEG[0] }),
    .S4BEG({\Tile_X1Y6_S4BEG[15] ,
    \Tile_X1Y6_S4BEG[14] ,
    \Tile_X1Y6_S4BEG[13] ,
    \Tile_X1Y6_S4BEG[12] ,
    \Tile_X1Y6_S4BEG[11] ,
    \Tile_X1Y6_S4BEG[10] ,
    \Tile_X1Y6_S4BEG[9] ,
    \Tile_X1Y6_S4BEG[8] ,
    \Tile_X1Y6_S4BEG[7] ,
    \Tile_X1Y6_S4BEG[6] ,
    \Tile_X1Y6_S4BEG[5] ,
    \Tile_X1Y6_S4BEG[4] ,
    \Tile_X1Y6_S4BEG[3] ,
    \Tile_X1Y6_S4BEG[2] ,
    \Tile_X1Y6_S4BEG[1] ,
    \Tile_X1Y6_S4BEG[0] }),
    .S4END({\Tile_X1Y5_S4BEG[15] ,
    \Tile_X1Y5_S4BEG[14] ,
    \Tile_X1Y5_S4BEG[13] ,
    \Tile_X1Y5_S4BEG[12] ,
    \Tile_X1Y5_S4BEG[11] ,
    \Tile_X1Y5_S4BEG[10] ,
    \Tile_X1Y5_S4BEG[9] ,
    \Tile_X1Y5_S4BEG[8] ,
    \Tile_X1Y5_S4BEG[7] ,
    \Tile_X1Y5_S4BEG[6] ,
    \Tile_X1Y5_S4BEG[5] ,
    \Tile_X1Y5_S4BEG[4] ,
    \Tile_X1Y5_S4BEG[3] ,
    \Tile_X1Y5_S4BEG[2] ,
    \Tile_X1Y5_S4BEG[1] ,
    \Tile_X1Y5_S4BEG[0] }),
    .SS4BEG({\Tile_X1Y6_SS4BEG[15] ,
    \Tile_X1Y6_SS4BEG[14] ,
    \Tile_X1Y6_SS4BEG[13] ,
    \Tile_X1Y6_SS4BEG[12] ,
    \Tile_X1Y6_SS4BEG[11] ,
    \Tile_X1Y6_SS4BEG[10] ,
    \Tile_X1Y6_SS4BEG[9] ,
    \Tile_X1Y6_SS4BEG[8] ,
    \Tile_X1Y6_SS4BEG[7] ,
    \Tile_X1Y6_SS4BEG[6] ,
    \Tile_X1Y6_SS4BEG[5] ,
    \Tile_X1Y6_SS4BEG[4] ,
    \Tile_X1Y6_SS4BEG[3] ,
    \Tile_X1Y6_SS4BEG[2] ,
    \Tile_X1Y6_SS4BEG[1] ,
    \Tile_X1Y6_SS4BEG[0] }),
    .SS4END({\Tile_X1Y5_SS4BEG[15] ,
    \Tile_X1Y5_SS4BEG[14] ,
    \Tile_X1Y5_SS4BEG[13] ,
    \Tile_X1Y5_SS4BEG[12] ,
    \Tile_X1Y5_SS4BEG[11] ,
    \Tile_X1Y5_SS4BEG[10] ,
    \Tile_X1Y5_SS4BEG[9] ,
    \Tile_X1Y5_SS4BEG[8] ,
    \Tile_X1Y5_SS4BEG[7] ,
    \Tile_X1Y5_SS4BEG[6] ,
    \Tile_X1Y5_SS4BEG[5] ,
    \Tile_X1Y5_SS4BEG[4] ,
    \Tile_X1Y5_SS4BEG[3] ,
    \Tile_X1Y5_SS4BEG[2] ,
    \Tile_X1Y5_SS4BEG[1] ,
    \Tile_X1Y5_SS4BEG[0] }),
    .W1BEG({\Tile_X1Y6_W1BEG[3] ,
    \Tile_X1Y6_W1BEG[2] ,
    \Tile_X1Y6_W1BEG[1] ,
    \Tile_X1Y6_W1BEG[0] }),
    .W1END({\Tile_X2Y6_W1BEG[3] ,
    \Tile_X2Y6_W1BEG[2] ,
    \Tile_X2Y6_W1BEG[1] ,
    \Tile_X2Y6_W1BEG[0] }),
    .W2BEG({\Tile_X1Y6_W2BEG[7] ,
    \Tile_X1Y6_W2BEG[6] ,
    \Tile_X1Y6_W2BEG[5] ,
    \Tile_X1Y6_W2BEG[4] ,
    \Tile_X1Y6_W2BEG[3] ,
    \Tile_X1Y6_W2BEG[2] ,
    \Tile_X1Y6_W2BEG[1] ,
    \Tile_X1Y6_W2BEG[0] }),
    .W2BEGb({\Tile_X1Y6_W2BEGb[7] ,
    \Tile_X1Y6_W2BEGb[6] ,
    \Tile_X1Y6_W2BEGb[5] ,
    \Tile_X1Y6_W2BEGb[4] ,
    \Tile_X1Y6_W2BEGb[3] ,
    \Tile_X1Y6_W2BEGb[2] ,
    \Tile_X1Y6_W2BEGb[1] ,
    \Tile_X1Y6_W2BEGb[0] }),
    .W2END({\Tile_X2Y6_W2BEGb[7] ,
    \Tile_X2Y6_W2BEGb[6] ,
    \Tile_X2Y6_W2BEGb[5] ,
    \Tile_X2Y6_W2BEGb[4] ,
    \Tile_X2Y6_W2BEGb[3] ,
    \Tile_X2Y6_W2BEGb[2] ,
    \Tile_X2Y6_W2BEGb[1] ,
    \Tile_X2Y6_W2BEGb[0] }),
    .W2MID({\Tile_X2Y6_W2BEG[7] ,
    \Tile_X2Y6_W2BEG[6] ,
    \Tile_X2Y6_W2BEG[5] ,
    \Tile_X2Y6_W2BEG[4] ,
    \Tile_X2Y6_W2BEG[3] ,
    \Tile_X2Y6_W2BEG[2] ,
    \Tile_X2Y6_W2BEG[1] ,
    \Tile_X2Y6_W2BEG[0] }),
    .W6BEG({\Tile_X1Y6_W6BEG[11] ,
    \Tile_X1Y6_W6BEG[10] ,
    \Tile_X1Y6_W6BEG[9] ,
    \Tile_X1Y6_W6BEG[8] ,
    \Tile_X1Y6_W6BEG[7] ,
    \Tile_X1Y6_W6BEG[6] ,
    \Tile_X1Y6_W6BEG[5] ,
    \Tile_X1Y6_W6BEG[4] ,
    \Tile_X1Y6_W6BEG[3] ,
    \Tile_X1Y6_W6BEG[2] ,
    \Tile_X1Y6_W6BEG[1] ,
    \Tile_X1Y6_W6BEG[0] }),
    .W6END({\Tile_X2Y6_W6BEG[11] ,
    \Tile_X2Y6_W6BEG[10] ,
    \Tile_X2Y6_W6BEG[9] ,
    \Tile_X2Y6_W6BEG[8] ,
    \Tile_X2Y6_W6BEG[7] ,
    \Tile_X2Y6_W6BEG[6] ,
    \Tile_X2Y6_W6BEG[5] ,
    \Tile_X2Y6_W6BEG[4] ,
    \Tile_X2Y6_W6BEG[3] ,
    \Tile_X2Y6_W6BEG[2] ,
    \Tile_X2Y6_W6BEG[1] ,
    \Tile_X2Y6_W6BEG[0] }),
    .WW4BEG({\Tile_X1Y6_WW4BEG[15] ,
    \Tile_X1Y6_WW4BEG[14] ,
    \Tile_X1Y6_WW4BEG[13] ,
    \Tile_X1Y6_WW4BEG[12] ,
    \Tile_X1Y6_WW4BEG[11] ,
    \Tile_X1Y6_WW4BEG[10] ,
    \Tile_X1Y6_WW4BEG[9] ,
    \Tile_X1Y6_WW4BEG[8] ,
    \Tile_X1Y6_WW4BEG[7] ,
    \Tile_X1Y6_WW4BEG[6] ,
    \Tile_X1Y6_WW4BEG[5] ,
    \Tile_X1Y6_WW4BEG[4] ,
    \Tile_X1Y6_WW4BEG[3] ,
    \Tile_X1Y6_WW4BEG[2] ,
    \Tile_X1Y6_WW4BEG[1] ,
    \Tile_X1Y6_WW4BEG[0] }),
    .WW4END({\Tile_X2Y6_WW4BEG[15] ,
    \Tile_X2Y6_WW4BEG[14] ,
    \Tile_X2Y6_WW4BEG[13] ,
    \Tile_X2Y6_WW4BEG[12] ,
    \Tile_X2Y6_WW4BEG[11] ,
    \Tile_X2Y6_WW4BEG[10] ,
    \Tile_X2Y6_WW4BEG[9] ,
    \Tile_X2Y6_WW4BEG[8] ,
    \Tile_X2Y6_WW4BEG[7] ,
    \Tile_X2Y6_WW4BEG[6] ,
    \Tile_X2Y6_WW4BEG[5] ,
    \Tile_X2Y6_WW4BEG[4] ,
    \Tile_X2Y6_WW4BEG[3] ,
    \Tile_X2Y6_WW4BEG[2] ,
    \Tile_X2Y6_WW4BEG[1] ,
    \Tile_X2Y6_WW4BEG[0] }));
 LUT4AB Tile_X1Y7_LUT4AB (.Ci(Tile_X1Y8_Co),
    .Co(Tile_X1Y7_Co),
    .UserCLK(Tile_X1Y8_UserCLKo),
    .UserCLKo(Tile_X1Y7_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X1Y7_E1BEG[3] ,
    \Tile_X1Y7_E1BEG[2] ,
    \Tile_X1Y7_E1BEG[1] ,
    \Tile_X1Y7_E1BEG[0] }),
    .E1END({\Tile_X0Y7_E1BEG[3] ,
    \Tile_X0Y7_E1BEG[2] ,
    \Tile_X0Y7_E1BEG[1] ,
    \Tile_X0Y7_E1BEG[0] }),
    .E2BEG({\Tile_X1Y7_E2BEG[7] ,
    \Tile_X1Y7_E2BEG[6] ,
    \Tile_X1Y7_E2BEG[5] ,
    \Tile_X1Y7_E2BEG[4] ,
    \Tile_X1Y7_E2BEG[3] ,
    \Tile_X1Y7_E2BEG[2] ,
    \Tile_X1Y7_E2BEG[1] ,
    \Tile_X1Y7_E2BEG[0] }),
    .E2BEGb({\Tile_X1Y7_E2BEGb[7] ,
    \Tile_X1Y7_E2BEGb[6] ,
    \Tile_X1Y7_E2BEGb[5] ,
    \Tile_X1Y7_E2BEGb[4] ,
    \Tile_X1Y7_E2BEGb[3] ,
    \Tile_X1Y7_E2BEGb[2] ,
    \Tile_X1Y7_E2BEGb[1] ,
    \Tile_X1Y7_E2BEGb[0] }),
    .E2END({\Tile_X0Y7_E2BEGb[7] ,
    \Tile_X0Y7_E2BEGb[6] ,
    \Tile_X0Y7_E2BEGb[5] ,
    \Tile_X0Y7_E2BEGb[4] ,
    \Tile_X0Y7_E2BEGb[3] ,
    \Tile_X0Y7_E2BEGb[2] ,
    \Tile_X0Y7_E2BEGb[1] ,
    \Tile_X0Y7_E2BEGb[0] }),
    .E2MID({\Tile_X0Y7_E2BEG[7] ,
    \Tile_X0Y7_E2BEG[6] ,
    \Tile_X0Y7_E2BEG[5] ,
    \Tile_X0Y7_E2BEG[4] ,
    \Tile_X0Y7_E2BEG[3] ,
    \Tile_X0Y7_E2BEG[2] ,
    \Tile_X0Y7_E2BEG[1] ,
    \Tile_X0Y7_E2BEG[0] }),
    .E6BEG({\Tile_X1Y7_E6BEG[11] ,
    \Tile_X1Y7_E6BEG[10] ,
    \Tile_X1Y7_E6BEG[9] ,
    \Tile_X1Y7_E6BEG[8] ,
    \Tile_X1Y7_E6BEG[7] ,
    \Tile_X1Y7_E6BEG[6] ,
    \Tile_X1Y7_E6BEG[5] ,
    \Tile_X1Y7_E6BEG[4] ,
    \Tile_X1Y7_E6BEG[3] ,
    \Tile_X1Y7_E6BEG[2] ,
    \Tile_X1Y7_E6BEG[1] ,
    \Tile_X1Y7_E6BEG[0] }),
    .E6END({\Tile_X0Y7_E6BEG[11] ,
    \Tile_X0Y7_E6BEG[10] ,
    \Tile_X0Y7_E6BEG[9] ,
    \Tile_X0Y7_E6BEG[8] ,
    \Tile_X0Y7_E6BEG[7] ,
    \Tile_X0Y7_E6BEG[6] ,
    \Tile_X0Y7_E6BEG[5] ,
    \Tile_X0Y7_E6BEG[4] ,
    \Tile_X0Y7_E6BEG[3] ,
    \Tile_X0Y7_E6BEG[2] ,
    \Tile_X0Y7_E6BEG[1] ,
    \Tile_X0Y7_E6BEG[0] }),
    .EE4BEG({\Tile_X1Y7_EE4BEG[15] ,
    \Tile_X1Y7_EE4BEG[14] ,
    \Tile_X1Y7_EE4BEG[13] ,
    \Tile_X1Y7_EE4BEG[12] ,
    \Tile_X1Y7_EE4BEG[11] ,
    \Tile_X1Y7_EE4BEG[10] ,
    \Tile_X1Y7_EE4BEG[9] ,
    \Tile_X1Y7_EE4BEG[8] ,
    \Tile_X1Y7_EE4BEG[7] ,
    \Tile_X1Y7_EE4BEG[6] ,
    \Tile_X1Y7_EE4BEG[5] ,
    \Tile_X1Y7_EE4BEG[4] ,
    \Tile_X1Y7_EE4BEG[3] ,
    \Tile_X1Y7_EE4BEG[2] ,
    \Tile_X1Y7_EE4BEG[1] ,
    \Tile_X1Y7_EE4BEG[0] }),
    .EE4END({\Tile_X0Y7_EE4BEG[15] ,
    \Tile_X0Y7_EE4BEG[14] ,
    \Tile_X0Y7_EE4BEG[13] ,
    \Tile_X0Y7_EE4BEG[12] ,
    \Tile_X0Y7_EE4BEG[11] ,
    \Tile_X0Y7_EE4BEG[10] ,
    \Tile_X0Y7_EE4BEG[9] ,
    \Tile_X0Y7_EE4BEG[8] ,
    \Tile_X0Y7_EE4BEG[7] ,
    \Tile_X0Y7_EE4BEG[6] ,
    \Tile_X0Y7_EE4BEG[5] ,
    \Tile_X0Y7_EE4BEG[4] ,
    \Tile_X0Y7_EE4BEG[3] ,
    \Tile_X0Y7_EE4BEG[2] ,
    \Tile_X0Y7_EE4BEG[1] ,
    \Tile_X0Y7_EE4BEG[0] }),
    .FrameData({\Tile_X0Y7_FrameData_O[31] ,
    \Tile_X0Y7_FrameData_O[30] ,
    \Tile_X0Y7_FrameData_O[29] ,
    \Tile_X0Y7_FrameData_O[28] ,
    \Tile_X0Y7_FrameData_O[27] ,
    \Tile_X0Y7_FrameData_O[26] ,
    \Tile_X0Y7_FrameData_O[25] ,
    \Tile_X0Y7_FrameData_O[24] ,
    \Tile_X0Y7_FrameData_O[23] ,
    \Tile_X0Y7_FrameData_O[22] ,
    \Tile_X0Y7_FrameData_O[21] ,
    \Tile_X0Y7_FrameData_O[20] ,
    \Tile_X0Y7_FrameData_O[19] ,
    \Tile_X0Y7_FrameData_O[18] ,
    \Tile_X0Y7_FrameData_O[17] ,
    \Tile_X0Y7_FrameData_O[16] ,
    \Tile_X0Y7_FrameData_O[15] ,
    \Tile_X0Y7_FrameData_O[14] ,
    \Tile_X0Y7_FrameData_O[13] ,
    \Tile_X0Y7_FrameData_O[12] ,
    \Tile_X0Y7_FrameData_O[11] ,
    \Tile_X0Y7_FrameData_O[10] ,
    \Tile_X0Y7_FrameData_O[9] ,
    \Tile_X0Y7_FrameData_O[8] ,
    \Tile_X0Y7_FrameData_O[7] ,
    \Tile_X0Y7_FrameData_O[6] ,
    \Tile_X0Y7_FrameData_O[5] ,
    \Tile_X0Y7_FrameData_O[4] ,
    \Tile_X0Y7_FrameData_O[3] ,
    \Tile_X0Y7_FrameData_O[2] ,
    \Tile_X0Y7_FrameData_O[1] ,
    \Tile_X0Y7_FrameData_O[0] }),
    .FrameData_O({\Tile_X1Y7_FrameData_O[31] ,
    \Tile_X1Y7_FrameData_O[30] ,
    \Tile_X1Y7_FrameData_O[29] ,
    \Tile_X1Y7_FrameData_O[28] ,
    \Tile_X1Y7_FrameData_O[27] ,
    \Tile_X1Y7_FrameData_O[26] ,
    \Tile_X1Y7_FrameData_O[25] ,
    \Tile_X1Y7_FrameData_O[24] ,
    \Tile_X1Y7_FrameData_O[23] ,
    \Tile_X1Y7_FrameData_O[22] ,
    \Tile_X1Y7_FrameData_O[21] ,
    \Tile_X1Y7_FrameData_O[20] ,
    \Tile_X1Y7_FrameData_O[19] ,
    \Tile_X1Y7_FrameData_O[18] ,
    \Tile_X1Y7_FrameData_O[17] ,
    \Tile_X1Y7_FrameData_O[16] ,
    \Tile_X1Y7_FrameData_O[15] ,
    \Tile_X1Y7_FrameData_O[14] ,
    \Tile_X1Y7_FrameData_O[13] ,
    \Tile_X1Y7_FrameData_O[12] ,
    \Tile_X1Y7_FrameData_O[11] ,
    \Tile_X1Y7_FrameData_O[10] ,
    \Tile_X1Y7_FrameData_O[9] ,
    \Tile_X1Y7_FrameData_O[8] ,
    \Tile_X1Y7_FrameData_O[7] ,
    \Tile_X1Y7_FrameData_O[6] ,
    \Tile_X1Y7_FrameData_O[5] ,
    \Tile_X1Y7_FrameData_O[4] ,
    \Tile_X1Y7_FrameData_O[3] ,
    \Tile_X1Y7_FrameData_O[2] ,
    \Tile_X1Y7_FrameData_O[1] ,
    \Tile_X1Y7_FrameData_O[0] }),
    .FrameStrobe({\Tile_X1Y8_FrameStrobe_O[19] ,
    \Tile_X1Y8_FrameStrobe_O[18] ,
    \Tile_X1Y8_FrameStrobe_O[17] ,
    \Tile_X1Y8_FrameStrobe_O[16] ,
    \Tile_X1Y8_FrameStrobe_O[15] ,
    \Tile_X1Y8_FrameStrobe_O[14] ,
    \Tile_X1Y8_FrameStrobe_O[13] ,
    \Tile_X1Y8_FrameStrobe_O[12] ,
    \Tile_X1Y8_FrameStrobe_O[11] ,
    \Tile_X1Y8_FrameStrobe_O[10] ,
    \Tile_X1Y8_FrameStrobe_O[9] ,
    \Tile_X1Y8_FrameStrobe_O[8] ,
    \Tile_X1Y8_FrameStrobe_O[7] ,
    \Tile_X1Y8_FrameStrobe_O[6] ,
    \Tile_X1Y8_FrameStrobe_O[5] ,
    \Tile_X1Y8_FrameStrobe_O[4] ,
    \Tile_X1Y8_FrameStrobe_O[3] ,
    \Tile_X1Y8_FrameStrobe_O[2] ,
    \Tile_X1Y8_FrameStrobe_O[1] ,
    \Tile_X1Y8_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X1Y7_FrameStrobe_O[19] ,
    \Tile_X1Y7_FrameStrobe_O[18] ,
    \Tile_X1Y7_FrameStrobe_O[17] ,
    \Tile_X1Y7_FrameStrobe_O[16] ,
    \Tile_X1Y7_FrameStrobe_O[15] ,
    \Tile_X1Y7_FrameStrobe_O[14] ,
    \Tile_X1Y7_FrameStrobe_O[13] ,
    \Tile_X1Y7_FrameStrobe_O[12] ,
    \Tile_X1Y7_FrameStrobe_O[11] ,
    \Tile_X1Y7_FrameStrobe_O[10] ,
    \Tile_X1Y7_FrameStrobe_O[9] ,
    \Tile_X1Y7_FrameStrobe_O[8] ,
    \Tile_X1Y7_FrameStrobe_O[7] ,
    \Tile_X1Y7_FrameStrobe_O[6] ,
    \Tile_X1Y7_FrameStrobe_O[5] ,
    \Tile_X1Y7_FrameStrobe_O[4] ,
    \Tile_X1Y7_FrameStrobe_O[3] ,
    \Tile_X1Y7_FrameStrobe_O[2] ,
    \Tile_X1Y7_FrameStrobe_O[1] ,
    \Tile_X1Y7_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X1Y7_N1BEG[3] ,
    \Tile_X1Y7_N1BEG[2] ,
    \Tile_X1Y7_N1BEG[1] ,
    \Tile_X1Y7_N1BEG[0] }),
    .N1END({\Tile_X1Y8_N1BEG[3] ,
    \Tile_X1Y8_N1BEG[2] ,
    \Tile_X1Y8_N1BEG[1] ,
    \Tile_X1Y8_N1BEG[0] }),
    .N2BEG({\Tile_X1Y7_N2BEG[7] ,
    \Tile_X1Y7_N2BEG[6] ,
    \Tile_X1Y7_N2BEG[5] ,
    \Tile_X1Y7_N2BEG[4] ,
    \Tile_X1Y7_N2BEG[3] ,
    \Tile_X1Y7_N2BEG[2] ,
    \Tile_X1Y7_N2BEG[1] ,
    \Tile_X1Y7_N2BEG[0] }),
    .N2BEGb({\Tile_X1Y7_N2BEGb[7] ,
    \Tile_X1Y7_N2BEGb[6] ,
    \Tile_X1Y7_N2BEGb[5] ,
    \Tile_X1Y7_N2BEGb[4] ,
    \Tile_X1Y7_N2BEGb[3] ,
    \Tile_X1Y7_N2BEGb[2] ,
    \Tile_X1Y7_N2BEGb[1] ,
    \Tile_X1Y7_N2BEGb[0] }),
    .N2END({\Tile_X1Y8_N2BEGb[7] ,
    \Tile_X1Y8_N2BEGb[6] ,
    \Tile_X1Y8_N2BEGb[5] ,
    \Tile_X1Y8_N2BEGb[4] ,
    \Tile_X1Y8_N2BEGb[3] ,
    \Tile_X1Y8_N2BEGb[2] ,
    \Tile_X1Y8_N2BEGb[1] ,
    \Tile_X1Y8_N2BEGb[0] }),
    .N2MID({\Tile_X1Y8_N2BEG[7] ,
    \Tile_X1Y8_N2BEG[6] ,
    \Tile_X1Y8_N2BEG[5] ,
    \Tile_X1Y8_N2BEG[4] ,
    \Tile_X1Y8_N2BEG[3] ,
    \Tile_X1Y8_N2BEG[2] ,
    \Tile_X1Y8_N2BEG[1] ,
    \Tile_X1Y8_N2BEG[0] }),
    .N4BEG({\Tile_X1Y7_N4BEG[15] ,
    \Tile_X1Y7_N4BEG[14] ,
    \Tile_X1Y7_N4BEG[13] ,
    \Tile_X1Y7_N4BEG[12] ,
    \Tile_X1Y7_N4BEG[11] ,
    \Tile_X1Y7_N4BEG[10] ,
    \Tile_X1Y7_N4BEG[9] ,
    \Tile_X1Y7_N4BEG[8] ,
    \Tile_X1Y7_N4BEG[7] ,
    \Tile_X1Y7_N4BEG[6] ,
    \Tile_X1Y7_N4BEG[5] ,
    \Tile_X1Y7_N4BEG[4] ,
    \Tile_X1Y7_N4BEG[3] ,
    \Tile_X1Y7_N4BEG[2] ,
    \Tile_X1Y7_N4BEG[1] ,
    \Tile_X1Y7_N4BEG[0] }),
    .N4END({\Tile_X1Y8_N4BEG[15] ,
    \Tile_X1Y8_N4BEG[14] ,
    \Tile_X1Y8_N4BEG[13] ,
    \Tile_X1Y8_N4BEG[12] ,
    \Tile_X1Y8_N4BEG[11] ,
    \Tile_X1Y8_N4BEG[10] ,
    \Tile_X1Y8_N4BEG[9] ,
    \Tile_X1Y8_N4BEG[8] ,
    \Tile_X1Y8_N4BEG[7] ,
    \Tile_X1Y8_N4BEG[6] ,
    \Tile_X1Y8_N4BEG[5] ,
    \Tile_X1Y8_N4BEG[4] ,
    \Tile_X1Y8_N4BEG[3] ,
    \Tile_X1Y8_N4BEG[2] ,
    \Tile_X1Y8_N4BEG[1] ,
    \Tile_X1Y8_N4BEG[0] }),
    .NN4BEG({\Tile_X1Y7_NN4BEG[15] ,
    \Tile_X1Y7_NN4BEG[14] ,
    \Tile_X1Y7_NN4BEG[13] ,
    \Tile_X1Y7_NN4BEG[12] ,
    \Tile_X1Y7_NN4BEG[11] ,
    \Tile_X1Y7_NN4BEG[10] ,
    \Tile_X1Y7_NN4BEG[9] ,
    \Tile_X1Y7_NN4BEG[8] ,
    \Tile_X1Y7_NN4BEG[7] ,
    \Tile_X1Y7_NN4BEG[6] ,
    \Tile_X1Y7_NN4BEG[5] ,
    \Tile_X1Y7_NN4BEG[4] ,
    \Tile_X1Y7_NN4BEG[3] ,
    \Tile_X1Y7_NN4BEG[2] ,
    \Tile_X1Y7_NN4BEG[1] ,
    \Tile_X1Y7_NN4BEG[0] }),
    .NN4END({\Tile_X1Y8_NN4BEG[15] ,
    \Tile_X1Y8_NN4BEG[14] ,
    \Tile_X1Y8_NN4BEG[13] ,
    \Tile_X1Y8_NN4BEG[12] ,
    \Tile_X1Y8_NN4BEG[11] ,
    \Tile_X1Y8_NN4BEG[10] ,
    \Tile_X1Y8_NN4BEG[9] ,
    \Tile_X1Y8_NN4BEG[8] ,
    \Tile_X1Y8_NN4BEG[7] ,
    \Tile_X1Y8_NN4BEG[6] ,
    \Tile_X1Y8_NN4BEG[5] ,
    \Tile_X1Y8_NN4BEG[4] ,
    \Tile_X1Y8_NN4BEG[3] ,
    \Tile_X1Y8_NN4BEG[2] ,
    \Tile_X1Y8_NN4BEG[1] ,
    \Tile_X1Y8_NN4BEG[0] }),
    .S1BEG({\Tile_X1Y7_S1BEG[3] ,
    \Tile_X1Y7_S1BEG[2] ,
    \Tile_X1Y7_S1BEG[1] ,
    \Tile_X1Y7_S1BEG[0] }),
    .S1END({\Tile_X1Y6_S1BEG[3] ,
    \Tile_X1Y6_S1BEG[2] ,
    \Tile_X1Y6_S1BEG[1] ,
    \Tile_X1Y6_S1BEG[0] }),
    .S2BEG({\Tile_X1Y7_S2BEG[7] ,
    \Tile_X1Y7_S2BEG[6] ,
    \Tile_X1Y7_S2BEG[5] ,
    \Tile_X1Y7_S2BEG[4] ,
    \Tile_X1Y7_S2BEG[3] ,
    \Tile_X1Y7_S2BEG[2] ,
    \Tile_X1Y7_S2BEG[1] ,
    \Tile_X1Y7_S2BEG[0] }),
    .S2BEGb({\Tile_X1Y7_S2BEGb[7] ,
    \Tile_X1Y7_S2BEGb[6] ,
    \Tile_X1Y7_S2BEGb[5] ,
    \Tile_X1Y7_S2BEGb[4] ,
    \Tile_X1Y7_S2BEGb[3] ,
    \Tile_X1Y7_S2BEGb[2] ,
    \Tile_X1Y7_S2BEGb[1] ,
    \Tile_X1Y7_S2BEGb[0] }),
    .S2END({\Tile_X1Y6_S2BEGb[7] ,
    \Tile_X1Y6_S2BEGb[6] ,
    \Tile_X1Y6_S2BEGb[5] ,
    \Tile_X1Y6_S2BEGb[4] ,
    \Tile_X1Y6_S2BEGb[3] ,
    \Tile_X1Y6_S2BEGb[2] ,
    \Tile_X1Y6_S2BEGb[1] ,
    \Tile_X1Y6_S2BEGb[0] }),
    .S2MID({\Tile_X1Y6_S2BEG[7] ,
    \Tile_X1Y6_S2BEG[6] ,
    \Tile_X1Y6_S2BEG[5] ,
    \Tile_X1Y6_S2BEG[4] ,
    \Tile_X1Y6_S2BEG[3] ,
    \Tile_X1Y6_S2BEG[2] ,
    \Tile_X1Y6_S2BEG[1] ,
    \Tile_X1Y6_S2BEG[0] }),
    .S4BEG({\Tile_X1Y7_S4BEG[15] ,
    \Tile_X1Y7_S4BEG[14] ,
    \Tile_X1Y7_S4BEG[13] ,
    \Tile_X1Y7_S4BEG[12] ,
    \Tile_X1Y7_S4BEG[11] ,
    \Tile_X1Y7_S4BEG[10] ,
    \Tile_X1Y7_S4BEG[9] ,
    \Tile_X1Y7_S4BEG[8] ,
    \Tile_X1Y7_S4BEG[7] ,
    \Tile_X1Y7_S4BEG[6] ,
    \Tile_X1Y7_S4BEG[5] ,
    \Tile_X1Y7_S4BEG[4] ,
    \Tile_X1Y7_S4BEG[3] ,
    \Tile_X1Y7_S4BEG[2] ,
    \Tile_X1Y7_S4BEG[1] ,
    \Tile_X1Y7_S4BEG[0] }),
    .S4END({\Tile_X1Y6_S4BEG[15] ,
    \Tile_X1Y6_S4BEG[14] ,
    \Tile_X1Y6_S4BEG[13] ,
    \Tile_X1Y6_S4BEG[12] ,
    \Tile_X1Y6_S4BEG[11] ,
    \Tile_X1Y6_S4BEG[10] ,
    \Tile_X1Y6_S4BEG[9] ,
    \Tile_X1Y6_S4BEG[8] ,
    \Tile_X1Y6_S4BEG[7] ,
    \Tile_X1Y6_S4BEG[6] ,
    \Tile_X1Y6_S4BEG[5] ,
    \Tile_X1Y6_S4BEG[4] ,
    \Tile_X1Y6_S4BEG[3] ,
    \Tile_X1Y6_S4BEG[2] ,
    \Tile_X1Y6_S4BEG[1] ,
    \Tile_X1Y6_S4BEG[0] }),
    .SS4BEG({\Tile_X1Y7_SS4BEG[15] ,
    \Tile_X1Y7_SS4BEG[14] ,
    \Tile_X1Y7_SS4BEG[13] ,
    \Tile_X1Y7_SS4BEG[12] ,
    \Tile_X1Y7_SS4BEG[11] ,
    \Tile_X1Y7_SS4BEG[10] ,
    \Tile_X1Y7_SS4BEG[9] ,
    \Tile_X1Y7_SS4BEG[8] ,
    \Tile_X1Y7_SS4BEG[7] ,
    \Tile_X1Y7_SS4BEG[6] ,
    \Tile_X1Y7_SS4BEG[5] ,
    \Tile_X1Y7_SS4BEG[4] ,
    \Tile_X1Y7_SS4BEG[3] ,
    \Tile_X1Y7_SS4BEG[2] ,
    \Tile_X1Y7_SS4BEG[1] ,
    \Tile_X1Y7_SS4BEG[0] }),
    .SS4END({\Tile_X1Y6_SS4BEG[15] ,
    \Tile_X1Y6_SS4BEG[14] ,
    \Tile_X1Y6_SS4BEG[13] ,
    \Tile_X1Y6_SS4BEG[12] ,
    \Tile_X1Y6_SS4BEG[11] ,
    \Tile_X1Y6_SS4BEG[10] ,
    \Tile_X1Y6_SS4BEG[9] ,
    \Tile_X1Y6_SS4BEG[8] ,
    \Tile_X1Y6_SS4BEG[7] ,
    \Tile_X1Y6_SS4BEG[6] ,
    \Tile_X1Y6_SS4BEG[5] ,
    \Tile_X1Y6_SS4BEG[4] ,
    \Tile_X1Y6_SS4BEG[3] ,
    \Tile_X1Y6_SS4BEG[2] ,
    \Tile_X1Y6_SS4BEG[1] ,
    \Tile_X1Y6_SS4BEG[0] }),
    .W1BEG({\Tile_X1Y7_W1BEG[3] ,
    \Tile_X1Y7_W1BEG[2] ,
    \Tile_X1Y7_W1BEG[1] ,
    \Tile_X1Y7_W1BEG[0] }),
    .W1END({\Tile_X2Y7_W1BEG[3] ,
    \Tile_X2Y7_W1BEG[2] ,
    \Tile_X2Y7_W1BEG[1] ,
    \Tile_X2Y7_W1BEG[0] }),
    .W2BEG({\Tile_X1Y7_W2BEG[7] ,
    \Tile_X1Y7_W2BEG[6] ,
    \Tile_X1Y7_W2BEG[5] ,
    \Tile_X1Y7_W2BEG[4] ,
    \Tile_X1Y7_W2BEG[3] ,
    \Tile_X1Y7_W2BEG[2] ,
    \Tile_X1Y7_W2BEG[1] ,
    \Tile_X1Y7_W2BEG[0] }),
    .W2BEGb({\Tile_X1Y7_W2BEGb[7] ,
    \Tile_X1Y7_W2BEGb[6] ,
    \Tile_X1Y7_W2BEGb[5] ,
    \Tile_X1Y7_W2BEGb[4] ,
    \Tile_X1Y7_W2BEGb[3] ,
    \Tile_X1Y7_W2BEGb[2] ,
    \Tile_X1Y7_W2BEGb[1] ,
    \Tile_X1Y7_W2BEGb[0] }),
    .W2END({\Tile_X2Y7_W2BEGb[7] ,
    \Tile_X2Y7_W2BEGb[6] ,
    \Tile_X2Y7_W2BEGb[5] ,
    \Tile_X2Y7_W2BEGb[4] ,
    \Tile_X2Y7_W2BEGb[3] ,
    \Tile_X2Y7_W2BEGb[2] ,
    \Tile_X2Y7_W2BEGb[1] ,
    \Tile_X2Y7_W2BEGb[0] }),
    .W2MID({\Tile_X2Y7_W2BEG[7] ,
    \Tile_X2Y7_W2BEG[6] ,
    \Tile_X2Y7_W2BEG[5] ,
    \Tile_X2Y7_W2BEG[4] ,
    \Tile_X2Y7_W2BEG[3] ,
    \Tile_X2Y7_W2BEG[2] ,
    \Tile_X2Y7_W2BEG[1] ,
    \Tile_X2Y7_W2BEG[0] }),
    .W6BEG({\Tile_X1Y7_W6BEG[11] ,
    \Tile_X1Y7_W6BEG[10] ,
    \Tile_X1Y7_W6BEG[9] ,
    \Tile_X1Y7_W6BEG[8] ,
    \Tile_X1Y7_W6BEG[7] ,
    \Tile_X1Y7_W6BEG[6] ,
    \Tile_X1Y7_W6BEG[5] ,
    \Tile_X1Y7_W6BEG[4] ,
    \Tile_X1Y7_W6BEG[3] ,
    \Tile_X1Y7_W6BEG[2] ,
    \Tile_X1Y7_W6BEG[1] ,
    \Tile_X1Y7_W6BEG[0] }),
    .W6END({\Tile_X2Y7_W6BEG[11] ,
    \Tile_X2Y7_W6BEG[10] ,
    \Tile_X2Y7_W6BEG[9] ,
    \Tile_X2Y7_W6BEG[8] ,
    \Tile_X2Y7_W6BEG[7] ,
    \Tile_X2Y7_W6BEG[6] ,
    \Tile_X2Y7_W6BEG[5] ,
    \Tile_X2Y7_W6BEG[4] ,
    \Tile_X2Y7_W6BEG[3] ,
    \Tile_X2Y7_W6BEG[2] ,
    \Tile_X2Y7_W6BEG[1] ,
    \Tile_X2Y7_W6BEG[0] }),
    .WW4BEG({\Tile_X1Y7_WW4BEG[15] ,
    \Tile_X1Y7_WW4BEG[14] ,
    \Tile_X1Y7_WW4BEG[13] ,
    \Tile_X1Y7_WW4BEG[12] ,
    \Tile_X1Y7_WW4BEG[11] ,
    \Tile_X1Y7_WW4BEG[10] ,
    \Tile_X1Y7_WW4BEG[9] ,
    \Tile_X1Y7_WW4BEG[8] ,
    \Tile_X1Y7_WW4BEG[7] ,
    \Tile_X1Y7_WW4BEG[6] ,
    \Tile_X1Y7_WW4BEG[5] ,
    \Tile_X1Y7_WW4BEG[4] ,
    \Tile_X1Y7_WW4BEG[3] ,
    \Tile_X1Y7_WW4BEG[2] ,
    \Tile_X1Y7_WW4BEG[1] ,
    \Tile_X1Y7_WW4BEG[0] }),
    .WW4END({\Tile_X2Y7_WW4BEG[15] ,
    \Tile_X2Y7_WW4BEG[14] ,
    \Tile_X2Y7_WW4BEG[13] ,
    \Tile_X2Y7_WW4BEG[12] ,
    \Tile_X2Y7_WW4BEG[11] ,
    \Tile_X2Y7_WW4BEG[10] ,
    \Tile_X2Y7_WW4BEG[9] ,
    \Tile_X2Y7_WW4BEG[8] ,
    \Tile_X2Y7_WW4BEG[7] ,
    \Tile_X2Y7_WW4BEG[6] ,
    \Tile_X2Y7_WW4BEG[5] ,
    \Tile_X2Y7_WW4BEG[4] ,
    \Tile_X2Y7_WW4BEG[3] ,
    \Tile_X2Y7_WW4BEG[2] ,
    \Tile_X2Y7_WW4BEG[1] ,
    \Tile_X2Y7_WW4BEG[0] }));
 LUT4AB Tile_X1Y8_LUT4AB (.Ci(Tile_X1Y9_Co),
    .Co(Tile_X1Y8_Co),
    .UserCLK(Tile_X1Y9_UserCLKo),
    .UserCLKo(Tile_X1Y8_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X1Y8_E1BEG[3] ,
    \Tile_X1Y8_E1BEG[2] ,
    \Tile_X1Y8_E1BEG[1] ,
    \Tile_X1Y8_E1BEG[0] }),
    .E1END({\Tile_X0Y8_E1BEG[3] ,
    \Tile_X0Y8_E1BEG[2] ,
    \Tile_X0Y8_E1BEG[1] ,
    \Tile_X0Y8_E1BEG[0] }),
    .E2BEG({\Tile_X1Y8_E2BEG[7] ,
    \Tile_X1Y8_E2BEG[6] ,
    \Tile_X1Y8_E2BEG[5] ,
    \Tile_X1Y8_E2BEG[4] ,
    \Tile_X1Y8_E2BEG[3] ,
    \Tile_X1Y8_E2BEG[2] ,
    \Tile_X1Y8_E2BEG[1] ,
    \Tile_X1Y8_E2BEG[0] }),
    .E2BEGb({\Tile_X1Y8_E2BEGb[7] ,
    \Tile_X1Y8_E2BEGb[6] ,
    \Tile_X1Y8_E2BEGb[5] ,
    \Tile_X1Y8_E2BEGb[4] ,
    \Tile_X1Y8_E2BEGb[3] ,
    \Tile_X1Y8_E2BEGb[2] ,
    \Tile_X1Y8_E2BEGb[1] ,
    \Tile_X1Y8_E2BEGb[0] }),
    .E2END({\Tile_X0Y8_E2BEGb[7] ,
    \Tile_X0Y8_E2BEGb[6] ,
    \Tile_X0Y8_E2BEGb[5] ,
    \Tile_X0Y8_E2BEGb[4] ,
    \Tile_X0Y8_E2BEGb[3] ,
    \Tile_X0Y8_E2BEGb[2] ,
    \Tile_X0Y8_E2BEGb[1] ,
    \Tile_X0Y8_E2BEGb[0] }),
    .E2MID({\Tile_X0Y8_E2BEG[7] ,
    \Tile_X0Y8_E2BEG[6] ,
    \Tile_X0Y8_E2BEG[5] ,
    \Tile_X0Y8_E2BEG[4] ,
    \Tile_X0Y8_E2BEG[3] ,
    \Tile_X0Y8_E2BEG[2] ,
    \Tile_X0Y8_E2BEG[1] ,
    \Tile_X0Y8_E2BEG[0] }),
    .E6BEG({\Tile_X1Y8_E6BEG[11] ,
    \Tile_X1Y8_E6BEG[10] ,
    \Tile_X1Y8_E6BEG[9] ,
    \Tile_X1Y8_E6BEG[8] ,
    \Tile_X1Y8_E6BEG[7] ,
    \Tile_X1Y8_E6BEG[6] ,
    \Tile_X1Y8_E6BEG[5] ,
    \Tile_X1Y8_E6BEG[4] ,
    \Tile_X1Y8_E6BEG[3] ,
    \Tile_X1Y8_E6BEG[2] ,
    \Tile_X1Y8_E6BEG[1] ,
    \Tile_X1Y8_E6BEG[0] }),
    .E6END({\Tile_X0Y8_E6BEG[11] ,
    \Tile_X0Y8_E6BEG[10] ,
    \Tile_X0Y8_E6BEG[9] ,
    \Tile_X0Y8_E6BEG[8] ,
    \Tile_X0Y8_E6BEG[7] ,
    \Tile_X0Y8_E6BEG[6] ,
    \Tile_X0Y8_E6BEG[5] ,
    \Tile_X0Y8_E6BEG[4] ,
    \Tile_X0Y8_E6BEG[3] ,
    \Tile_X0Y8_E6BEG[2] ,
    \Tile_X0Y8_E6BEG[1] ,
    \Tile_X0Y8_E6BEG[0] }),
    .EE4BEG({\Tile_X1Y8_EE4BEG[15] ,
    \Tile_X1Y8_EE4BEG[14] ,
    \Tile_X1Y8_EE4BEG[13] ,
    \Tile_X1Y8_EE4BEG[12] ,
    \Tile_X1Y8_EE4BEG[11] ,
    \Tile_X1Y8_EE4BEG[10] ,
    \Tile_X1Y8_EE4BEG[9] ,
    \Tile_X1Y8_EE4BEG[8] ,
    \Tile_X1Y8_EE4BEG[7] ,
    \Tile_X1Y8_EE4BEG[6] ,
    \Tile_X1Y8_EE4BEG[5] ,
    \Tile_X1Y8_EE4BEG[4] ,
    \Tile_X1Y8_EE4BEG[3] ,
    \Tile_X1Y8_EE4BEG[2] ,
    \Tile_X1Y8_EE4BEG[1] ,
    \Tile_X1Y8_EE4BEG[0] }),
    .EE4END({\Tile_X0Y8_EE4BEG[15] ,
    \Tile_X0Y8_EE4BEG[14] ,
    \Tile_X0Y8_EE4BEG[13] ,
    \Tile_X0Y8_EE4BEG[12] ,
    \Tile_X0Y8_EE4BEG[11] ,
    \Tile_X0Y8_EE4BEG[10] ,
    \Tile_X0Y8_EE4BEG[9] ,
    \Tile_X0Y8_EE4BEG[8] ,
    \Tile_X0Y8_EE4BEG[7] ,
    \Tile_X0Y8_EE4BEG[6] ,
    \Tile_X0Y8_EE4BEG[5] ,
    \Tile_X0Y8_EE4BEG[4] ,
    \Tile_X0Y8_EE4BEG[3] ,
    \Tile_X0Y8_EE4BEG[2] ,
    \Tile_X0Y8_EE4BEG[1] ,
    \Tile_X0Y8_EE4BEG[0] }),
    .FrameData({\Tile_X0Y8_FrameData_O[31] ,
    \Tile_X0Y8_FrameData_O[30] ,
    \Tile_X0Y8_FrameData_O[29] ,
    \Tile_X0Y8_FrameData_O[28] ,
    \Tile_X0Y8_FrameData_O[27] ,
    \Tile_X0Y8_FrameData_O[26] ,
    \Tile_X0Y8_FrameData_O[25] ,
    \Tile_X0Y8_FrameData_O[24] ,
    \Tile_X0Y8_FrameData_O[23] ,
    \Tile_X0Y8_FrameData_O[22] ,
    \Tile_X0Y8_FrameData_O[21] ,
    \Tile_X0Y8_FrameData_O[20] ,
    \Tile_X0Y8_FrameData_O[19] ,
    \Tile_X0Y8_FrameData_O[18] ,
    \Tile_X0Y8_FrameData_O[17] ,
    \Tile_X0Y8_FrameData_O[16] ,
    \Tile_X0Y8_FrameData_O[15] ,
    \Tile_X0Y8_FrameData_O[14] ,
    \Tile_X0Y8_FrameData_O[13] ,
    \Tile_X0Y8_FrameData_O[12] ,
    \Tile_X0Y8_FrameData_O[11] ,
    \Tile_X0Y8_FrameData_O[10] ,
    \Tile_X0Y8_FrameData_O[9] ,
    \Tile_X0Y8_FrameData_O[8] ,
    \Tile_X0Y8_FrameData_O[7] ,
    \Tile_X0Y8_FrameData_O[6] ,
    \Tile_X0Y8_FrameData_O[5] ,
    \Tile_X0Y8_FrameData_O[4] ,
    \Tile_X0Y8_FrameData_O[3] ,
    \Tile_X0Y8_FrameData_O[2] ,
    \Tile_X0Y8_FrameData_O[1] ,
    \Tile_X0Y8_FrameData_O[0] }),
    .FrameData_O({\Tile_X1Y8_FrameData_O[31] ,
    \Tile_X1Y8_FrameData_O[30] ,
    \Tile_X1Y8_FrameData_O[29] ,
    \Tile_X1Y8_FrameData_O[28] ,
    \Tile_X1Y8_FrameData_O[27] ,
    \Tile_X1Y8_FrameData_O[26] ,
    \Tile_X1Y8_FrameData_O[25] ,
    \Tile_X1Y8_FrameData_O[24] ,
    \Tile_X1Y8_FrameData_O[23] ,
    \Tile_X1Y8_FrameData_O[22] ,
    \Tile_X1Y8_FrameData_O[21] ,
    \Tile_X1Y8_FrameData_O[20] ,
    \Tile_X1Y8_FrameData_O[19] ,
    \Tile_X1Y8_FrameData_O[18] ,
    \Tile_X1Y8_FrameData_O[17] ,
    \Tile_X1Y8_FrameData_O[16] ,
    \Tile_X1Y8_FrameData_O[15] ,
    \Tile_X1Y8_FrameData_O[14] ,
    \Tile_X1Y8_FrameData_O[13] ,
    \Tile_X1Y8_FrameData_O[12] ,
    \Tile_X1Y8_FrameData_O[11] ,
    \Tile_X1Y8_FrameData_O[10] ,
    \Tile_X1Y8_FrameData_O[9] ,
    \Tile_X1Y8_FrameData_O[8] ,
    \Tile_X1Y8_FrameData_O[7] ,
    \Tile_X1Y8_FrameData_O[6] ,
    \Tile_X1Y8_FrameData_O[5] ,
    \Tile_X1Y8_FrameData_O[4] ,
    \Tile_X1Y8_FrameData_O[3] ,
    \Tile_X1Y8_FrameData_O[2] ,
    \Tile_X1Y8_FrameData_O[1] ,
    \Tile_X1Y8_FrameData_O[0] }),
    .FrameStrobe({\Tile_X1Y9_FrameStrobe_O[19] ,
    \Tile_X1Y9_FrameStrobe_O[18] ,
    \Tile_X1Y9_FrameStrobe_O[17] ,
    \Tile_X1Y9_FrameStrobe_O[16] ,
    \Tile_X1Y9_FrameStrobe_O[15] ,
    \Tile_X1Y9_FrameStrobe_O[14] ,
    \Tile_X1Y9_FrameStrobe_O[13] ,
    \Tile_X1Y9_FrameStrobe_O[12] ,
    \Tile_X1Y9_FrameStrobe_O[11] ,
    \Tile_X1Y9_FrameStrobe_O[10] ,
    \Tile_X1Y9_FrameStrobe_O[9] ,
    \Tile_X1Y9_FrameStrobe_O[8] ,
    \Tile_X1Y9_FrameStrobe_O[7] ,
    \Tile_X1Y9_FrameStrobe_O[6] ,
    \Tile_X1Y9_FrameStrobe_O[5] ,
    \Tile_X1Y9_FrameStrobe_O[4] ,
    \Tile_X1Y9_FrameStrobe_O[3] ,
    \Tile_X1Y9_FrameStrobe_O[2] ,
    \Tile_X1Y9_FrameStrobe_O[1] ,
    \Tile_X1Y9_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X1Y8_FrameStrobe_O[19] ,
    \Tile_X1Y8_FrameStrobe_O[18] ,
    \Tile_X1Y8_FrameStrobe_O[17] ,
    \Tile_X1Y8_FrameStrobe_O[16] ,
    \Tile_X1Y8_FrameStrobe_O[15] ,
    \Tile_X1Y8_FrameStrobe_O[14] ,
    \Tile_X1Y8_FrameStrobe_O[13] ,
    \Tile_X1Y8_FrameStrobe_O[12] ,
    \Tile_X1Y8_FrameStrobe_O[11] ,
    \Tile_X1Y8_FrameStrobe_O[10] ,
    \Tile_X1Y8_FrameStrobe_O[9] ,
    \Tile_X1Y8_FrameStrobe_O[8] ,
    \Tile_X1Y8_FrameStrobe_O[7] ,
    \Tile_X1Y8_FrameStrobe_O[6] ,
    \Tile_X1Y8_FrameStrobe_O[5] ,
    \Tile_X1Y8_FrameStrobe_O[4] ,
    \Tile_X1Y8_FrameStrobe_O[3] ,
    \Tile_X1Y8_FrameStrobe_O[2] ,
    \Tile_X1Y8_FrameStrobe_O[1] ,
    \Tile_X1Y8_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X1Y8_N1BEG[3] ,
    \Tile_X1Y8_N1BEG[2] ,
    \Tile_X1Y8_N1BEG[1] ,
    \Tile_X1Y8_N1BEG[0] }),
    .N1END({\Tile_X1Y9_N1BEG[3] ,
    \Tile_X1Y9_N1BEG[2] ,
    \Tile_X1Y9_N1BEG[1] ,
    \Tile_X1Y9_N1BEG[0] }),
    .N2BEG({\Tile_X1Y8_N2BEG[7] ,
    \Tile_X1Y8_N2BEG[6] ,
    \Tile_X1Y8_N2BEG[5] ,
    \Tile_X1Y8_N2BEG[4] ,
    \Tile_X1Y8_N2BEG[3] ,
    \Tile_X1Y8_N2BEG[2] ,
    \Tile_X1Y8_N2BEG[1] ,
    \Tile_X1Y8_N2BEG[0] }),
    .N2BEGb({\Tile_X1Y8_N2BEGb[7] ,
    \Tile_X1Y8_N2BEGb[6] ,
    \Tile_X1Y8_N2BEGb[5] ,
    \Tile_X1Y8_N2BEGb[4] ,
    \Tile_X1Y8_N2BEGb[3] ,
    \Tile_X1Y8_N2BEGb[2] ,
    \Tile_X1Y8_N2BEGb[1] ,
    \Tile_X1Y8_N2BEGb[0] }),
    .N2END({\Tile_X1Y9_N2BEGb[7] ,
    \Tile_X1Y9_N2BEGb[6] ,
    \Tile_X1Y9_N2BEGb[5] ,
    \Tile_X1Y9_N2BEGb[4] ,
    \Tile_X1Y9_N2BEGb[3] ,
    \Tile_X1Y9_N2BEGb[2] ,
    \Tile_X1Y9_N2BEGb[1] ,
    \Tile_X1Y9_N2BEGb[0] }),
    .N2MID({\Tile_X1Y9_N2BEG[7] ,
    \Tile_X1Y9_N2BEG[6] ,
    \Tile_X1Y9_N2BEG[5] ,
    \Tile_X1Y9_N2BEG[4] ,
    \Tile_X1Y9_N2BEG[3] ,
    \Tile_X1Y9_N2BEG[2] ,
    \Tile_X1Y9_N2BEG[1] ,
    \Tile_X1Y9_N2BEG[0] }),
    .N4BEG({\Tile_X1Y8_N4BEG[15] ,
    \Tile_X1Y8_N4BEG[14] ,
    \Tile_X1Y8_N4BEG[13] ,
    \Tile_X1Y8_N4BEG[12] ,
    \Tile_X1Y8_N4BEG[11] ,
    \Tile_X1Y8_N4BEG[10] ,
    \Tile_X1Y8_N4BEG[9] ,
    \Tile_X1Y8_N4BEG[8] ,
    \Tile_X1Y8_N4BEG[7] ,
    \Tile_X1Y8_N4BEG[6] ,
    \Tile_X1Y8_N4BEG[5] ,
    \Tile_X1Y8_N4BEG[4] ,
    \Tile_X1Y8_N4BEG[3] ,
    \Tile_X1Y8_N4BEG[2] ,
    \Tile_X1Y8_N4BEG[1] ,
    \Tile_X1Y8_N4BEG[0] }),
    .N4END({\Tile_X1Y9_N4BEG[15] ,
    \Tile_X1Y9_N4BEG[14] ,
    \Tile_X1Y9_N4BEG[13] ,
    \Tile_X1Y9_N4BEG[12] ,
    \Tile_X1Y9_N4BEG[11] ,
    \Tile_X1Y9_N4BEG[10] ,
    \Tile_X1Y9_N4BEG[9] ,
    \Tile_X1Y9_N4BEG[8] ,
    \Tile_X1Y9_N4BEG[7] ,
    \Tile_X1Y9_N4BEG[6] ,
    \Tile_X1Y9_N4BEG[5] ,
    \Tile_X1Y9_N4BEG[4] ,
    \Tile_X1Y9_N4BEG[3] ,
    \Tile_X1Y9_N4BEG[2] ,
    \Tile_X1Y9_N4BEG[1] ,
    \Tile_X1Y9_N4BEG[0] }),
    .NN4BEG({\Tile_X1Y8_NN4BEG[15] ,
    \Tile_X1Y8_NN4BEG[14] ,
    \Tile_X1Y8_NN4BEG[13] ,
    \Tile_X1Y8_NN4BEG[12] ,
    \Tile_X1Y8_NN4BEG[11] ,
    \Tile_X1Y8_NN4BEG[10] ,
    \Tile_X1Y8_NN4BEG[9] ,
    \Tile_X1Y8_NN4BEG[8] ,
    \Tile_X1Y8_NN4BEG[7] ,
    \Tile_X1Y8_NN4BEG[6] ,
    \Tile_X1Y8_NN4BEG[5] ,
    \Tile_X1Y8_NN4BEG[4] ,
    \Tile_X1Y8_NN4BEG[3] ,
    \Tile_X1Y8_NN4BEG[2] ,
    \Tile_X1Y8_NN4BEG[1] ,
    \Tile_X1Y8_NN4BEG[0] }),
    .NN4END({\Tile_X1Y9_NN4BEG[15] ,
    \Tile_X1Y9_NN4BEG[14] ,
    \Tile_X1Y9_NN4BEG[13] ,
    \Tile_X1Y9_NN4BEG[12] ,
    \Tile_X1Y9_NN4BEG[11] ,
    \Tile_X1Y9_NN4BEG[10] ,
    \Tile_X1Y9_NN4BEG[9] ,
    \Tile_X1Y9_NN4BEG[8] ,
    \Tile_X1Y9_NN4BEG[7] ,
    \Tile_X1Y9_NN4BEG[6] ,
    \Tile_X1Y9_NN4BEG[5] ,
    \Tile_X1Y9_NN4BEG[4] ,
    \Tile_X1Y9_NN4BEG[3] ,
    \Tile_X1Y9_NN4BEG[2] ,
    \Tile_X1Y9_NN4BEG[1] ,
    \Tile_X1Y9_NN4BEG[0] }),
    .S1BEG({\Tile_X1Y8_S1BEG[3] ,
    \Tile_X1Y8_S1BEG[2] ,
    \Tile_X1Y8_S1BEG[1] ,
    \Tile_X1Y8_S1BEG[0] }),
    .S1END({\Tile_X1Y7_S1BEG[3] ,
    \Tile_X1Y7_S1BEG[2] ,
    \Tile_X1Y7_S1BEG[1] ,
    \Tile_X1Y7_S1BEG[0] }),
    .S2BEG({\Tile_X1Y8_S2BEG[7] ,
    \Tile_X1Y8_S2BEG[6] ,
    \Tile_X1Y8_S2BEG[5] ,
    \Tile_X1Y8_S2BEG[4] ,
    \Tile_X1Y8_S2BEG[3] ,
    \Tile_X1Y8_S2BEG[2] ,
    \Tile_X1Y8_S2BEG[1] ,
    \Tile_X1Y8_S2BEG[0] }),
    .S2BEGb({\Tile_X1Y8_S2BEGb[7] ,
    \Tile_X1Y8_S2BEGb[6] ,
    \Tile_X1Y8_S2BEGb[5] ,
    \Tile_X1Y8_S2BEGb[4] ,
    \Tile_X1Y8_S2BEGb[3] ,
    \Tile_X1Y8_S2BEGb[2] ,
    \Tile_X1Y8_S2BEGb[1] ,
    \Tile_X1Y8_S2BEGb[0] }),
    .S2END({\Tile_X1Y7_S2BEGb[7] ,
    \Tile_X1Y7_S2BEGb[6] ,
    \Tile_X1Y7_S2BEGb[5] ,
    \Tile_X1Y7_S2BEGb[4] ,
    \Tile_X1Y7_S2BEGb[3] ,
    \Tile_X1Y7_S2BEGb[2] ,
    \Tile_X1Y7_S2BEGb[1] ,
    \Tile_X1Y7_S2BEGb[0] }),
    .S2MID({\Tile_X1Y7_S2BEG[7] ,
    \Tile_X1Y7_S2BEG[6] ,
    \Tile_X1Y7_S2BEG[5] ,
    \Tile_X1Y7_S2BEG[4] ,
    \Tile_X1Y7_S2BEG[3] ,
    \Tile_X1Y7_S2BEG[2] ,
    \Tile_X1Y7_S2BEG[1] ,
    \Tile_X1Y7_S2BEG[0] }),
    .S4BEG({\Tile_X1Y8_S4BEG[15] ,
    \Tile_X1Y8_S4BEG[14] ,
    \Tile_X1Y8_S4BEG[13] ,
    \Tile_X1Y8_S4BEG[12] ,
    \Tile_X1Y8_S4BEG[11] ,
    \Tile_X1Y8_S4BEG[10] ,
    \Tile_X1Y8_S4BEG[9] ,
    \Tile_X1Y8_S4BEG[8] ,
    \Tile_X1Y8_S4BEG[7] ,
    \Tile_X1Y8_S4BEG[6] ,
    \Tile_X1Y8_S4BEG[5] ,
    \Tile_X1Y8_S4BEG[4] ,
    \Tile_X1Y8_S4BEG[3] ,
    \Tile_X1Y8_S4BEG[2] ,
    \Tile_X1Y8_S4BEG[1] ,
    \Tile_X1Y8_S4BEG[0] }),
    .S4END({\Tile_X1Y7_S4BEG[15] ,
    \Tile_X1Y7_S4BEG[14] ,
    \Tile_X1Y7_S4BEG[13] ,
    \Tile_X1Y7_S4BEG[12] ,
    \Tile_X1Y7_S4BEG[11] ,
    \Tile_X1Y7_S4BEG[10] ,
    \Tile_X1Y7_S4BEG[9] ,
    \Tile_X1Y7_S4BEG[8] ,
    \Tile_X1Y7_S4BEG[7] ,
    \Tile_X1Y7_S4BEG[6] ,
    \Tile_X1Y7_S4BEG[5] ,
    \Tile_X1Y7_S4BEG[4] ,
    \Tile_X1Y7_S4BEG[3] ,
    \Tile_X1Y7_S4BEG[2] ,
    \Tile_X1Y7_S4BEG[1] ,
    \Tile_X1Y7_S4BEG[0] }),
    .SS4BEG({\Tile_X1Y8_SS4BEG[15] ,
    \Tile_X1Y8_SS4BEG[14] ,
    \Tile_X1Y8_SS4BEG[13] ,
    \Tile_X1Y8_SS4BEG[12] ,
    \Tile_X1Y8_SS4BEG[11] ,
    \Tile_X1Y8_SS4BEG[10] ,
    \Tile_X1Y8_SS4BEG[9] ,
    \Tile_X1Y8_SS4BEG[8] ,
    \Tile_X1Y8_SS4BEG[7] ,
    \Tile_X1Y8_SS4BEG[6] ,
    \Tile_X1Y8_SS4BEG[5] ,
    \Tile_X1Y8_SS4BEG[4] ,
    \Tile_X1Y8_SS4BEG[3] ,
    \Tile_X1Y8_SS4BEG[2] ,
    \Tile_X1Y8_SS4BEG[1] ,
    \Tile_X1Y8_SS4BEG[0] }),
    .SS4END({\Tile_X1Y7_SS4BEG[15] ,
    \Tile_X1Y7_SS4BEG[14] ,
    \Tile_X1Y7_SS4BEG[13] ,
    \Tile_X1Y7_SS4BEG[12] ,
    \Tile_X1Y7_SS4BEG[11] ,
    \Tile_X1Y7_SS4BEG[10] ,
    \Tile_X1Y7_SS4BEG[9] ,
    \Tile_X1Y7_SS4BEG[8] ,
    \Tile_X1Y7_SS4BEG[7] ,
    \Tile_X1Y7_SS4BEG[6] ,
    \Tile_X1Y7_SS4BEG[5] ,
    \Tile_X1Y7_SS4BEG[4] ,
    \Tile_X1Y7_SS4BEG[3] ,
    \Tile_X1Y7_SS4BEG[2] ,
    \Tile_X1Y7_SS4BEG[1] ,
    \Tile_X1Y7_SS4BEG[0] }),
    .W1BEG({\Tile_X1Y8_W1BEG[3] ,
    \Tile_X1Y8_W1BEG[2] ,
    \Tile_X1Y8_W1BEG[1] ,
    \Tile_X1Y8_W1BEG[0] }),
    .W1END({\Tile_X2Y8_W1BEG[3] ,
    \Tile_X2Y8_W1BEG[2] ,
    \Tile_X2Y8_W1BEG[1] ,
    \Tile_X2Y8_W1BEG[0] }),
    .W2BEG({\Tile_X1Y8_W2BEG[7] ,
    \Tile_X1Y8_W2BEG[6] ,
    \Tile_X1Y8_W2BEG[5] ,
    \Tile_X1Y8_W2BEG[4] ,
    \Tile_X1Y8_W2BEG[3] ,
    \Tile_X1Y8_W2BEG[2] ,
    \Tile_X1Y8_W2BEG[1] ,
    \Tile_X1Y8_W2BEG[0] }),
    .W2BEGb({\Tile_X1Y8_W2BEGb[7] ,
    \Tile_X1Y8_W2BEGb[6] ,
    \Tile_X1Y8_W2BEGb[5] ,
    \Tile_X1Y8_W2BEGb[4] ,
    \Tile_X1Y8_W2BEGb[3] ,
    \Tile_X1Y8_W2BEGb[2] ,
    \Tile_X1Y8_W2BEGb[1] ,
    \Tile_X1Y8_W2BEGb[0] }),
    .W2END({\Tile_X2Y8_W2BEGb[7] ,
    \Tile_X2Y8_W2BEGb[6] ,
    \Tile_X2Y8_W2BEGb[5] ,
    \Tile_X2Y8_W2BEGb[4] ,
    \Tile_X2Y8_W2BEGb[3] ,
    \Tile_X2Y8_W2BEGb[2] ,
    \Tile_X2Y8_W2BEGb[1] ,
    \Tile_X2Y8_W2BEGb[0] }),
    .W2MID({\Tile_X2Y8_W2BEG[7] ,
    \Tile_X2Y8_W2BEG[6] ,
    \Tile_X2Y8_W2BEG[5] ,
    \Tile_X2Y8_W2BEG[4] ,
    \Tile_X2Y8_W2BEG[3] ,
    \Tile_X2Y8_W2BEG[2] ,
    \Tile_X2Y8_W2BEG[1] ,
    \Tile_X2Y8_W2BEG[0] }),
    .W6BEG({\Tile_X1Y8_W6BEG[11] ,
    \Tile_X1Y8_W6BEG[10] ,
    \Tile_X1Y8_W6BEG[9] ,
    \Tile_X1Y8_W6BEG[8] ,
    \Tile_X1Y8_W6BEG[7] ,
    \Tile_X1Y8_W6BEG[6] ,
    \Tile_X1Y8_W6BEG[5] ,
    \Tile_X1Y8_W6BEG[4] ,
    \Tile_X1Y8_W6BEG[3] ,
    \Tile_X1Y8_W6BEG[2] ,
    \Tile_X1Y8_W6BEG[1] ,
    \Tile_X1Y8_W6BEG[0] }),
    .W6END({\Tile_X2Y8_W6BEG[11] ,
    \Tile_X2Y8_W6BEG[10] ,
    \Tile_X2Y8_W6BEG[9] ,
    \Tile_X2Y8_W6BEG[8] ,
    \Tile_X2Y8_W6BEG[7] ,
    \Tile_X2Y8_W6BEG[6] ,
    \Tile_X2Y8_W6BEG[5] ,
    \Tile_X2Y8_W6BEG[4] ,
    \Tile_X2Y8_W6BEG[3] ,
    \Tile_X2Y8_W6BEG[2] ,
    \Tile_X2Y8_W6BEG[1] ,
    \Tile_X2Y8_W6BEG[0] }),
    .WW4BEG({\Tile_X1Y8_WW4BEG[15] ,
    \Tile_X1Y8_WW4BEG[14] ,
    \Tile_X1Y8_WW4BEG[13] ,
    \Tile_X1Y8_WW4BEG[12] ,
    \Tile_X1Y8_WW4BEG[11] ,
    \Tile_X1Y8_WW4BEG[10] ,
    \Tile_X1Y8_WW4BEG[9] ,
    \Tile_X1Y8_WW4BEG[8] ,
    \Tile_X1Y8_WW4BEG[7] ,
    \Tile_X1Y8_WW4BEG[6] ,
    \Tile_X1Y8_WW4BEG[5] ,
    \Tile_X1Y8_WW4BEG[4] ,
    \Tile_X1Y8_WW4BEG[3] ,
    \Tile_X1Y8_WW4BEG[2] ,
    \Tile_X1Y8_WW4BEG[1] ,
    \Tile_X1Y8_WW4BEG[0] }),
    .WW4END({\Tile_X2Y8_WW4BEG[15] ,
    \Tile_X2Y8_WW4BEG[14] ,
    \Tile_X2Y8_WW4BEG[13] ,
    \Tile_X2Y8_WW4BEG[12] ,
    \Tile_X2Y8_WW4BEG[11] ,
    \Tile_X2Y8_WW4BEG[10] ,
    \Tile_X2Y8_WW4BEG[9] ,
    \Tile_X2Y8_WW4BEG[8] ,
    \Tile_X2Y8_WW4BEG[7] ,
    \Tile_X2Y8_WW4BEG[6] ,
    \Tile_X2Y8_WW4BEG[5] ,
    \Tile_X2Y8_WW4BEG[4] ,
    \Tile_X2Y8_WW4BEG[3] ,
    \Tile_X2Y8_WW4BEG[2] ,
    \Tile_X2Y8_WW4BEG[1] ,
    \Tile_X2Y8_WW4BEG[0] }));
 S_IO4 Tile_X1Y9_S_IO4 (.A_I_top(Tile_X1Y9_A_I_top),
    .A_O_top(Tile_X1Y9_A_O_top),
    .A_T_top(Tile_X1Y9_A_T_top),
    .B_I_top(Tile_X1Y9_B_I_top),
    .B_O_top(Tile_X1Y9_B_O_top),
    .B_T_top(Tile_X1Y9_B_T_top),
    .C_I_top(Tile_X1Y9_C_I_top),
    .C_O_top(Tile_X1Y9_C_O_top),
    .C_T_top(Tile_X1Y9_C_T_top),
    .Co(Tile_X1Y9_Co),
    .D_I_top(Tile_X1Y9_D_I_top),
    .D_O_top(Tile_X1Y9_D_O_top),
    .D_T_top(Tile_X1Y9_D_T_top),
    .UserCLK(UserCLK),
    .UserCLKo(Tile_X1Y9_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .FrameData({\Tile_X0Y9_FrameData_O[31] ,
    \Tile_X0Y9_FrameData_O[30] ,
    \Tile_X0Y9_FrameData_O[29] ,
    \Tile_X0Y9_FrameData_O[28] ,
    \Tile_X0Y9_FrameData_O[27] ,
    \Tile_X0Y9_FrameData_O[26] ,
    \Tile_X0Y9_FrameData_O[25] ,
    \Tile_X0Y9_FrameData_O[24] ,
    \Tile_X0Y9_FrameData_O[23] ,
    \Tile_X0Y9_FrameData_O[22] ,
    \Tile_X0Y9_FrameData_O[21] ,
    \Tile_X0Y9_FrameData_O[20] ,
    \Tile_X0Y9_FrameData_O[19] ,
    \Tile_X0Y9_FrameData_O[18] ,
    \Tile_X0Y9_FrameData_O[17] ,
    \Tile_X0Y9_FrameData_O[16] ,
    \Tile_X0Y9_FrameData_O[15] ,
    \Tile_X0Y9_FrameData_O[14] ,
    \Tile_X0Y9_FrameData_O[13] ,
    \Tile_X0Y9_FrameData_O[12] ,
    \Tile_X0Y9_FrameData_O[11] ,
    \Tile_X0Y9_FrameData_O[10] ,
    \Tile_X0Y9_FrameData_O[9] ,
    \Tile_X0Y9_FrameData_O[8] ,
    \Tile_X0Y9_FrameData_O[7] ,
    \Tile_X0Y9_FrameData_O[6] ,
    \Tile_X0Y9_FrameData_O[5] ,
    \Tile_X0Y9_FrameData_O[4] ,
    \Tile_X0Y9_FrameData_O[3] ,
    \Tile_X0Y9_FrameData_O[2] ,
    \Tile_X0Y9_FrameData_O[1] ,
    \Tile_X0Y9_FrameData_O[0] }),
    .FrameData_O({\Tile_X1Y9_FrameData_O[31] ,
    \Tile_X1Y9_FrameData_O[30] ,
    \Tile_X1Y9_FrameData_O[29] ,
    \Tile_X1Y9_FrameData_O[28] ,
    \Tile_X1Y9_FrameData_O[27] ,
    \Tile_X1Y9_FrameData_O[26] ,
    \Tile_X1Y9_FrameData_O[25] ,
    \Tile_X1Y9_FrameData_O[24] ,
    \Tile_X1Y9_FrameData_O[23] ,
    \Tile_X1Y9_FrameData_O[22] ,
    \Tile_X1Y9_FrameData_O[21] ,
    \Tile_X1Y9_FrameData_O[20] ,
    \Tile_X1Y9_FrameData_O[19] ,
    \Tile_X1Y9_FrameData_O[18] ,
    \Tile_X1Y9_FrameData_O[17] ,
    \Tile_X1Y9_FrameData_O[16] ,
    \Tile_X1Y9_FrameData_O[15] ,
    \Tile_X1Y9_FrameData_O[14] ,
    \Tile_X1Y9_FrameData_O[13] ,
    \Tile_X1Y9_FrameData_O[12] ,
    \Tile_X1Y9_FrameData_O[11] ,
    \Tile_X1Y9_FrameData_O[10] ,
    \Tile_X1Y9_FrameData_O[9] ,
    \Tile_X1Y9_FrameData_O[8] ,
    \Tile_X1Y9_FrameData_O[7] ,
    \Tile_X1Y9_FrameData_O[6] ,
    \Tile_X1Y9_FrameData_O[5] ,
    \Tile_X1Y9_FrameData_O[4] ,
    \Tile_X1Y9_FrameData_O[3] ,
    \Tile_X1Y9_FrameData_O[2] ,
    \Tile_X1Y9_FrameData_O[1] ,
    \Tile_X1Y9_FrameData_O[0] }),
    .FrameStrobe({FrameStrobe[39],
    FrameStrobe[38],
    FrameStrobe[37],
    FrameStrobe[36],
    FrameStrobe[35],
    FrameStrobe[34],
    FrameStrobe[33],
    FrameStrobe[32],
    FrameStrobe[31],
    FrameStrobe[30],
    FrameStrobe[29],
    FrameStrobe[28],
    FrameStrobe[27],
    FrameStrobe[26],
    FrameStrobe[25],
    FrameStrobe[24],
    FrameStrobe[23],
    FrameStrobe[22],
    FrameStrobe[21],
    FrameStrobe[20]}),
    .FrameStrobe_O({\Tile_X1Y9_FrameStrobe_O[19] ,
    \Tile_X1Y9_FrameStrobe_O[18] ,
    \Tile_X1Y9_FrameStrobe_O[17] ,
    \Tile_X1Y9_FrameStrobe_O[16] ,
    \Tile_X1Y9_FrameStrobe_O[15] ,
    \Tile_X1Y9_FrameStrobe_O[14] ,
    \Tile_X1Y9_FrameStrobe_O[13] ,
    \Tile_X1Y9_FrameStrobe_O[12] ,
    \Tile_X1Y9_FrameStrobe_O[11] ,
    \Tile_X1Y9_FrameStrobe_O[10] ,
    \Tile_X1Y9_FrameStrobe_O[9] ,
    \Tile_X1Y9_FrameStrobe_O[8] ,
    \Tile_X1Y9_FrameStrobe_O[7] ,
    \Tile_X1Y9_FrameStrobe_O[6] ,
    \Tile_X1Y9_FrameStrobe_O[5] ,
    \Tile_X1Y9_FrameStrobe_O[4] ,
    \Tile_X1Y9_FrameStrobe_O[3] ,
    \Tile_X1Y9_FrameStrobe_O[2] ,
    \Tile_X1Y9_FrameStrobe_O[1] ,
    \Tile_X1Y9_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X1Y9_N1BEG[3] ,
    \Tile_X1Y9_N1BEG[2] ,
    \Tile_X1Y9_N1BEG[1] ,
    \Tile_X1Y9_N1BEG[0] }),
    .N2BEG({\Tile_X1Y9_N2BEG[7] ,
    \Tile_X1Y9_N2BEG[6] ,
    \Tile_X1Y9_N2BEG[5] ,
    \Tile_X1Y9_N2BEG[4] ,
    \Tile_X1Y9_N2BEG[3] ,
    \Tile_X1Y9_N2BEG[2] ,
    \Tile_X1Y9_N2BEG[1] ,
    \Tile_X1Y9_N2BEG[0] }),
    .N2BEGb({\Tile_X1Y9_N2BEGb[7] ,
    \Tile_X1Y9_N2BEGb[6] ,
    \Tile_X1Y9_N2BEGb[5] ,
    \Tile_X1Y9_N2BEGb[4] ,
    \Tile_X1Y9_N2BEGb[3] ,
    \Tile_X1Y9_N2BEGb[2] ,
    \Tile_X1Y9_N2BEGb[1] ,
    \Tile_X1Y9_N2BEGb[0] }),
    .N4BEG({\Tile_X1Y9_N4BEG[15] ,
    \Tile_X1Y9_N4BEG[14] ,
    \Tile_X1Y9_N4BEG[13] ,
    \Tile_X1Y9_N4BEG[12] ,
    \Tile_X1Y9_N4BEG[11] ,
    \Tile_X1Y9_N4BEG[10] ,
    \Tile_X1Y9_N4BEG[9] ,
    \Tile_X1Y9_N4BEG[8] ,
    \Tile_X1Y9_N4BEG[7] ,
    \Tile_X1Y9_N4BEG[6] ,
    \Tile_X1Y9_N4BEG[5] ,
    \Tile_X1Y9_N4BEG[4] ,
    \Tile_X1Y9_N4BEG[3] ,
    \Tile_X1Y9_N4BEG[2] ,
    \Tile_X1Y9_N4BEG[1] ,
    \Tile_X1Y9_N4BEG[0] }),
    .NN4BEG({\Tile_X1Y9_NN4BEG[15] ,
    \Tile_X1Y9_NN4BEG[14] ,
    \Tile_X1Y9_NN4BEG[13] ,
    \Tile_X1Y9_NN4BEG[12] ,
    \Tile_X1Y9_NN4BEG[11] ,
    \Tile_X1Y9_NN4BEG[10] ,
    \Tile_X1Y9_NN4BEG[9] ,
    \Tile_X1Y9_NN4BEG[8] ,
    \Tile_X1Y9_NN4BEG[7] ,
    \Tile_X1Y9_NN4BEG[6] ,
    \Tile_X1Y9_NN4BEG[5] ,
    \Tile_X1Y9_NN4BEG[4] ,
    \Tile_X1Y9_NN4BEG[3] ,
    \Tile_X1Y9_NN4BEG[2] ,
    \Tile_X1Y9_NN4BEG[1] ,
    \Tile_X1Y9_NN4BEG[0] }),
    .S1END({\Tile_X1Y8_S1BEG[3] ,
    \Tile_X1Y8_S1BEG[2] ,
    \Tile_X1Y8_S1BEG[1] ,
    \Tile_X1Y8_S1BEG[0] }),
    .S2END({\Tile_X1Y8_S2BEGb[7] ,
    \Tile_X1Y8_S2BEGb[6] ,
    \Tile_X1Y8_S2BEGb[5] ,
    \Tile_X1Y8_S2BEGb[4] ,
    \Tile_X1Y8_S2BEGb[3] ,
    \Tile_X1Y8_S2BEGb[2] ,
    \Tile_X1Y8_S2BEGb[1] ,
    \Tile_X1Y8_S2BEGb[0] }),
    .S2MID({\Tile_X1Y8_S2BEG[7] ,
    \Tile_X1Y8_S2BEG[6] ,
    \Tile_X1Y8_S2BEG[5] ,
    \Tile_X1Y8_S2BEG[4] ,
    \Tile_X1Y8_S2BEG[3] ,
    \Tile_X1Y8_S2BEG[2] ,
    \Tile_X1Y8_S2BEG[1] ,
    \Tile_X1Y8_S2BEG[0] }),
    .S4END({\Tile_X1Y8_S4BEG[15] ,
    \Tile_X1Y8_S4BEG[14] ,
    \Tile_X1Y8_S4BEG[13] ,
    \Tile_X1Y8_S4BEG[12] ,
    \Tile_X1Y8_S4BEG[11] ,
    \Tile_X1Y8_S4BEG[10] ,
    \Tile_X1Y8_S4BEG[9] ,
    \Tile_X1Y8_S4BEG[8] ,
    \Tile_X1Y8_S4BEG[7] ,
    \Tile_X1Y8_S4BEG[6] ,
    \Tile_X1Y8_S4BEG[5] ,
    \Tile_X1Y8_S4BEG[4] ,
    \Tile_X1Y8_S4BEG[3] ,
    \Tile_X1Y8_S4BEG[2] ,
    \Tile_X1Y8_S4BEG[1] ,
    \Tile_X1Y8_S4BEG[0] }),
    .SS4END({\Tile_X1Y8_SS4BEG[15] ,
    \Tile_X1Y8_SS4BEG[14] ,
    \Tile_X1Y8_SS4BEG[13] ,
    \Tile_X1Y8_SS4BEG[12] ,
    \Tile_X1Y8_SS4BEG[11] ,
    \Tile_X1Y8_SS4BEG[10] ,
    \Tile_X1Y8_SS4BEG[9] ,
    \Tile_X1Y8_SS4BEG[8] ,
    \Tile_X1Y8_SS4BEG[7] ,
    \Tile_X1Y8_SS4BEG[6] ,
    \Tile_X1Y8_SS4BEG[5] ,
    \Tile_X1Y8_SS4BEG[4] ,
    \Tile_X1Y8_SS4BEG[3] ,
    \Tile_X1Y8_SS4BEG[2] ,
    \Tile_X1Y8_SS4BEG[1] ,
    \Tile_X1Y8_SS4BEG[0] }));
 N_IO4 Tile_X2Y0_N_IO4 (.A_I_top(Tile_X2Y0_A_I_top),
    .A_O_top(Tile_X2Y0_A_O_top),
    .A_T_top(Tile_X2Y0_A_T_top),
    .B_I_top(Tile_X2Y0_B_I_top),
    .B_O_top(Tile_X2Y0_B_O_top),
    .B_T_top(Tile_X2Y0_B_T_top),
    .C_I_top(Tile_X2Y0_C_I_top),
    .C_O_top(Tile_X2Y0_C_O_top),
    .C_T_top(Tile_X2Y0_C_T_top),
    .Ci(Tile_X2Y1_Co),
    .D_I_top(Tile_X2Y0_D_I_top),
    .D_O_top(Tile_X2Y0_D_O_top),
    .D_T_top(Tile_X2Y0_D_T_top),
    .UserCLK(Tile_X2Y1_UserCLKo),
    .UserCLKo(Tile_X2Y0_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .FrameData({\Tile_X1Y0_FrameData_O[31] ,
    \Tile_X1Y0_FrameData_O[30] ,
    \Tile_X1Y0_FrameData_O[29] ,
    \Tile_X1Y0_FrameData_O[28] ,
    \Tile_X1Y0_FrameData_O[27] ,
    \Tile_X1Y0_FrameData_O[26] ,
    \Tile_X1Y0_FrameData_O[25] ,
    \Tile_X1Y0_FrameData_O[24] ,
    \Tile_X1Y0_FrameData_O[23] ,
    \Tile_X1Y0_FrameData_O[22] ,
    \Tile_X1Y0_FrameData_O[21] ,
    \Tile_X1Y0_FrameData_O[20] ,
    \Tile_X1Y0_FrameData_O[19] ,
    \Tile_X1Y0_FrameData_O[18] ,
    \Tile_X1Y0_FrameData_O[17] ,
    \Tile_X1Y0_FrameData_O[16] ,
    \Tile_X1Y0_FrameData_O[15] ,
    \Tile_X1Y0_FrameData_O[14] ,
    \Tile_X1Y0_FrameData_O[13] ,
    \Tile_X1Y0_FrameData_O[12] ,
    \Tile_X1Y0_FrameData_O[11] ,
    \Tile_X1Y0_FrameData_O[10] ,
    \Tile_X1Y0_FrameData_O[9] ,
    \Tile_X1Y0_FrameData_O[8] ,
    \Tile_X1Y0_FrameData_O[7] ,
    \Tile_X1Y0_FrameData_O[6] ,
    \Tile_X1Y0_FrameData_O[5] ,
    \Tile_X1Y0_FrameData_O[4] ,
    \Tile_X1Y0_FrameData_O[3] ,
    \Tile_X1Y0_FrameData_O[2] ,
    \Tile_X1Y0_FrameData_O[1] ,
    \Tile_X1Y0_FrameData_O[0] }),
    .FrameData_O({\Tile_X2Y0_FrameData_O[31] ,
    \Tile_X2Y0_FrameData_O[30] ,
    \Tile_X2Y0_FrameData_O[29] ,
    \Tile_X2Y0_FrameData_O[28] ,
    \Tile_X2Y0_FrameData_O[27] ,
    \Tile_X2Y0_FrameData_O[26] ,
    \Tile_X2Y0_FrameData_O[25] ,
    \Tile_X2Y0_FrameData_O[24] ,
    \Tile_X2Y0_FrameData_O[23] ,
    \Tile_X2Y0_FrameData_O[22] ,
    \Tile_X2Y0_FrameData_O[21] ,
    \Tile_X2Y0_FrameData_O[20] ,
    \Tile_X2Y0_FrameData_O[19] ,
    \Tile_X2Y0_FrameData_O[18] ,
    \Tile_X2Y0_FrameData_O[17] ,
    \Tile_X2Y0_FrameData_O[16] ,
    \Tile_X2Y0_FrameData_O[15] ,
    \Tile_X2Y0_FrameData_O[14] ,
    \Tile_X2Y0_FrameData_O[13] ,
    \Tile_X2Y0_FrameData_O[12] ,
    \Tile_X2Y0_FrameData_O[11] ,
    \Tile_X2Y0_FrameData_O[10] ,
    \Tile_X2Y0_FrameData_O[9] ,
    \Tile_X2Y0_FrameData_O[8] ,
    \Tile_X2Y0_FrameData_O[7] ,
    \Tile_X2Y0_FrameData_O[6] ,
    \Tile_X2Y0_FrameData_O[5] ,
    \Tile_X2Y0_FrameData_O[4] ,
    \Tile_X2Y0_FrameData_O[3] ,
    \Tile_X2Y0_FrameData_O[2] ,
    \Tile_X2Y0_FrameData_O[1] ,
    \Tile_X2Y0_FrameData_O[0] }),
    .FrameStrobe({\Tile_X2Y1_FrameStrobe_O[19] ,
    \Tile_X2Y1_FrameStrobe_O[18] ,
    \Tile_X2Y1_FrameStrobe_O[17] ,
    \Tile_X2Y1_FrameStrobe_O[16] ,
    \Tile_X2Y1_FrameStrobe_O[15] ,
    \Tile_X2Y1_FrameStrobe_O[14] ,
    \Tile_X2Y1_FrameStrobe_O[13] ,
    \Tile_X2Y1_FrameStrobe_O[12] ,
    \Tile_X2Y1_FrameStrobe_O[11] ,
    \Tile_X2Y1_FrameStrobe_O[10] ,
    \Tile_X2Y1_FrameStrobe_O[9] ,
    \Tile_X2Y1_FrameStrobe_O[8] ,
    \Tile_X2Y1_FrameStrobe_O[7] ,
    \Tile_X2Y1_FrameStrobe_O[6] ,
    \Tile_X2Y1_FrameStrobe_O[5] ,
    \Tile_X2Y1_FrameStrobe_O[4] ,
    \Tile_X2Y1_FrameStrobe_O[3] ,
    \Tile_X2Y1_FrameStrobe_O[2] ,
    \Tile_X2Y1_FrameStrobe_O[1] ,
    \Tile_X2Y1_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X2Y0_FrameStrobe_O[19] ,
    \Tile_X2Y0_FrameStrobe_O[18] ,
    \Tile_X2Y0_FrameStrobe_O[17] ,
    \Tile_X2Y0_FrameStrobe_O[16] ,
    \Tile_X2Y0_FrameStrobe_O[15] ,
    \Tile_X2Y0_FrameStrobe_O[14] ,
    \Tile_X2Y0_FrameStrobe_O[13] ,
    \Tile_X2Y0_FrameStrobe_O[12] ,
    \Tile_X2Y0_FrameStrobe_O[11] ,
    \Tile_X2Y0_FrameStrobe_O[10] ,
    \Tile_X2Y0_FrameStrobe_O[9] ,
    \Tile_X2Y0_FrameStrobe_O[8] ,
    \Tile_X2Y0_FrameStrobe_O[7] ,
    \Tile_X2Y0_FrameStrobe_O[6] ,
    \Tile_X2Y0_FrameStrobe_O[5] ,
    \Tile_X2Y0_FrameStrobe_O[4] ,
    \Tile_X2Y0_FrameStrobe_O[3] ,
    \Tile_X2Y0_FrameStrobe_O[2] ,
    \Tile_X2Y0_FrameStrobe_O[1] ,
    \Tile_X2Y0_FrameStrobe_O[0] }),
    .N1END({\Tile_X2Y1_N1BEG[3] ,
    \Tile_X2Y1_N1BEG[2] ,
    \Tile_X2Y1_N1BEG[1] ,
    \Tile_X2Y1_N1BEG[0] }),
    .N2END({\Tile_X2Y1_N2BEGb[7] ,
    \Tile_X2Y1_N2BEGb[6] ,
    \Tile_X2Y1_N2BEGb[5] ,
    \Tile_X2Y1_N2BEGb[4] ,
    \Tile_X2Y1_N2BEGb[3] ,
    \Tile_X2Y1_N2BEGb[2] ,
    \Tile_X2Y1_N2BEGb[1] ,
    \Tile_X2Y1_N2BEGb[0] }),
    .N2MID({\Tile_X2Y1_N2BEG[7] ,
    \Tile_X2Y1_N2BEG[6] ,
    \Tile_X2Y1_N2BEG[5] ,
    \Tile_X2Y1_N2BEG[4] ,
    \Tile_X2Y1_N2BEG[3] ,
    \Tile_X2Y1_N2BEG[2] ,
    \Tile_X2Y1_N2BEG[1] ,
    \Tile_X2Y1_N2BEG[0] }),
    .N4END({\Tile_X2Y1_N4BEG[15] ,
    \Tile_X2Y1_N4BEG[14] ,
    \Tile_X2Y1_N4BEG[13] ,
    \Tile_X2Y1_N4BEG[12] ,
    \Tile_X2Y1_N4BEG[11] ,
    \Tile_X2Y1_N4BEG[10] ,
    \Tile_X2Y1_N4BEG[9] ,
    \Tile_X2Y1_N4BEG[8] ,
    \Tile_X2Y1_N4BEG[7] ,
    \Tile_X2Y1_N4BEG[6] ,
    \Tile_X2Y1_N4BEG[5] ,
    \Tile_X2Y1_N4BEG[4] ,
    \Tile_X2Y1_N4BEG[3] ,
    \Tile_X2Y1_N4BEG[2] ,
    \Tile_X2Y1_N4BEG[1] ,
    \Tile_X2Y1_N4BEG[0] }),
    .NN4END({\Tile_X2Y1_NN4BEG[15] ,
    \Tile_X2Y1_NN4BEG[14] ,
    \Tile_X2Y1_NN4BEG[13] ,
    \Tile_X2Y1_NN4BEG[12] ,
    \Tile_X2Y1_NN4BEG[11] ,
    \Tile_X2Y1_NN4BEG[10] ,
    \Tile_X2Y1_NN4BEG[9] ,
    \Tile_X2Y1_NN4BEG[8] ,
    \Tile_X2Y1_NN4BEG[7] ,
    \Tile_X2Y1_NN4BEG[6] ,
    \Tile_X2Y1_NN4BEG[5] ,
    \Tile_X2Y1_NN4BEG[4] ,
    \Tile_X2Y1_NN4BEG[3] ,
    \Tile_X2Y1_NN4BEG[2] ,
    \Tile_X2Y1_NN4BEG[1] ,
    \Tile_X2Y1_NN4BEG[0] }),
    .S1BEG({\Tile_X2Y0_S1BEG[3] ,
    \Tile_X2Y0_S1BEG[2] ,
    \Tile_X2Y0_S1BEG[1] ,
    \Tile_X2Y0_S1BEG[0] }),
    .S2BEG({\Tile_X2Y0_S2BEG[7] ,
    \Tile_X2Y0_S2BEG[6] ,
    \Tile_X2Y0_S2BEG[5] ,
    \Tile_X2Y0_S2BEG[4] ,
    \Tile_X2Y0_S2BEG[3] ,
    \Tile_X2Y0_S2BEG[2] ,
    \Tile_X2Y0_S2BEG[1] ,
    \Tile_X2Y0_S2BEG[0] }),
    .S2BEGb({\Tile_X2Y0_S2BEGb[7] ,
    \Tile_X2Y0_S2BEGb[6] ,
    \Tile_X2Y0_S2BEGb[5] ,
    \Tile_X2Y0_S2BEGb[4] ,
    \Tile_X2Y0_S2BEGb[3] ,
    \Tile_X2Y0_S2BEGb[2] ,
    \Tile_X2Y0_S2BEGb[1] ,
    \Tile_X2Y0_S2BEGb[0] }),
    .S4BEG({\Tile_X2Y0_S4BEG[15] ,
    \Tile_X2Y0_S4BEG[14] ,
    \Tile_X2Y0_S4BEG[13] ,
    \Tile_X2Y0_S4BEG[12] ,
    \Tile_X2Y0_S4BEG[11] ,
    \Tile_X2Y0_S4BEG[10] ,
    \Tile_X2Y0_S4BEG[9] ,
    \Tile_X2Y0_S4BEG[8] ,
    \Tile_X2Y0_S4BEG[7] ,
    \Tile_X2Y0_S4BEG[6] ,
    \Tile_X2Y0_S4BEG[5] ,
    \Tile_X2Y0_S4BEG[4] ,
    \Tile_X2Y0_S4BEG[3] ,
    \Tile_X2Y0_S4BEG[2] ,
    \Tile_X2Y0_S4BEG[1] ,
    \Tile_X2Y0_S4BEG[0] }),
    .SS4BEG({\Tile_X2Y0_SS4BEG[15] ,
    \Tile_X2Y0_SS4BEG[14] ,
    \Tile_X2Y0_SS4BEG[13] ,
    \Tile_X2Y0_SS4BEG[12] ,
    \Tile_X2Y0_SS4BEG[11] ,
    \Tile_X2Y0_SS4BEG[10] ,
    \Tile_X2Y0_SS4BEG[9] ,
    \Tile_X2Y0_SS4BEG[8] ,
    \Tile_X2Y0_SS4BEG[7] ,
    \Tile_X2Y0_SS4BEG[6] ,
    \Tile_X2Y0_SS4BEG[5] ,
    \Tile_X2Y0_SS4BEG[4] ,
    \Tile_X2Y0_SS4BEG[3] ,
    \Tile_X2Y0_SS4BEG[2] ,
    \Tile_X2Y0_SS4BEG[1] ,
    \Tile_X2Y0_SS4BEG[0] }));
 LUT4AB Tile_X2Y1_LUT4AB (.Ci(Tile_X2Y2_Co),
    .Co(Tile_X2Y1_Co),
    .UserCLK(Tile_X2Y2_UserCLKo),
    .UserCLKo(Tile_X2Y1_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X2Y1_E1BEG[3] ,
    \Tile_X2Y1_E1BEG[2] ,
    \Tile_X2Y1_E1BEG[1] ,
    \Tile_X2Y1_E1BEG[0] }),
    .E1END({\Tile_X1Y1_E1BEG[3] ,
    \Tile_X1Y1_E1BEG[2] ,
    \Tile_X1Y1_E1BEG[1] ,
    \Tile_X1Y1_E1BEG[0] }),
    .E2BEG({\Tile_X2Y1_E2BEG[7] ,
    \Tile_X2Y1_E2BEG[6] ,
    \Tile_X2Y1_E2BEG[5] ,
    \Tile_X2Y1_E2BEG[4] ,
    \Tile_X2Y1_E2BEG[3] ,
    \Tile_X2Y1_E2BEG[2] ,
    \Tile_X2Y1_E2BEG[1] ,
    \Tile_X2Y1_E2BEG[0] }),
    .E2BEGb({\Tile_X2Y1_E2BEGb[7] ,
    \Tile_X2Y1_E2BEGb[6] ,
    \Tile_X2Y1_E2BEGb[5] ,
    \Tile_X2Y1_E2BEGb[4] ,
    \Tile_X2Y1_E2BEGb[3] ,
    \Tile_X2Y1_E2BEGb[2] ,
    \Tile_X2Y1_E2BEGb[1] ,
    \Tile_X2Y1_E2BEGb[0] }),
    .E2END({\Tile_X1Y1_E2BEGb[7] ,
    \Tile_X1Y1_E2BEGb[6] ,
    \Tile_X1Y1_E2BEGb[5] ,
    \Tile_X1Y1_E2BEGb[4] ,
    \Tile_X1Y1_E2BEGb[3] ,
    \Tile_X1Y1_E2BEGb[2] ,
    \Tile_X1Y1_E2BEGb[1] ,
    \Tile_X1Y1_E2BEGb[0] }),
    .E2MID({\Tile_X1Y1_E2BEG[7] ,
    \Tile_X1Y1_E2BEG[6] ,
    \Tile_X1Y1_E2BEG[5] ,
    \Tile_X1Y1_E2BEG[4] ,
    \Tile_X1Y1_E2BEG[3] ,
    \Tile_X1Y1_E2BEG[2] ,
    \Tile_X1Y1_E2BEG[1] ,
    \Tile_X1Y1_E2BEG[0] }),
    .E6BEG({\Tile_X2Y1_E6BEG[11] ,
    \Tile_X2Y1_E6BEG[10] ,
    \Tile_X2Y1_E6BEG[9] ,
    \Tile_X2Y1_E6BEG[8] ,
    \Tile_X2Y1_E6BEG[7] ,
    \Tile_X2Y1_E6BEG[6] ,
    \Tile_X2Y1_E6BEG[5] ,
    \Tile_X2Y1_E6BEG[4] ,
    \Tile_X2Y1_E6BEG[3] ,
    \Tile_X2Y1_E6BEG[2] ,
    \Tile_X2Y1_E6BEG[1] ,
    \Tile_X2Y1_E6BEG[0] }),
    .E6END({\Tile_X1Y1_E6BEG[11] ,
    \Tile_X1Y1_E6BEG[10] ,
    \Tile_X1Y1_E6BEG[9] ,
    \Tile_X1Y1_E6BEG[8] ,
    \Tile_X1Y1_E6BEG[7] ,
    \Tile_X1Y1_E6BEG[6] ,
    \Tile_X1Y1_E6BEG[5] ,
    \Tile_X1Y1_E6BEG[4] ,
    \Tile_X1Y1_E6BEG[3] ,
    \Tile_X1Y1_E6BEG[2] ,
    \Tile_X1Y1_E6BEG[1] ,
    \Tile_X1Y1_E6BEG[0] }),
    .EE4BEG({\Tile_X2Y1_EE4BEG[15] ,
    \Tile_X2Y1_EE4BEG[14] ,
    \Tile_X2Y1_EE4BEG[13] ,
    \Tile_X2Y1_EE4BEG[12] ,
    \Tile_X2Y1_EE4BEG[11] ,
    \Tile_X2Y1_EE4BEG[10] ,
    \Tile_X2Y1_EE4BEG[9] ,
    \Tile_X2Y1_EE4BEG[8] ,
    \Tile_X2Y1_EE4BEG[7] ,
    \Tile_X2Y1_EE4BEG[6] ,
    \Tile_X2Y1_EE4BEG[5] ,
    \Tile_X2Y1_EE4BEG[4] ,
    \Tile_X2Y1_EE4BEG[3] ,
    \Tile_X2Y1_EE4BEG[2] ,
    \Tile_X2Y1_EE4BEG[1] ,
    \Tile_X2Y1_EE4BEG[0] }),
    .EE4END({\Tile_X1Y1_EE4BEG[15] ,
    \Tile_X1Y1_EE4BEG[14] ,
    \Tile_X1Y1_EE4BEG[13] ,
    \Tile_X1Y1_EE4BEG[12] ,
    \Tile_X1Y1_EE4BEG[11] ,
    \Tile_X1Y1_EE4BEG[10] ,
    \Tile_X1Y1_EE4BEG[9] ,
    \Tile_X1Y1_EE4BEG[8] ,
    \Tile_X1Y1_EE4BEG[7] ,
    \Tile_X1Y1_EE4BEG[6] ,
    \Tile_X1Y1_EE4BEG[5] ,
    \Tile_X1Y1_EE4BEG[4] ,
    \Tile_X1Y1_EE4BEG[3] ,
    \Tile_X1Y1_EE4BEG[2] ,
    \Tile_X1Y1_EE4BEG[1] ,
    \Tile_X1Y1_EE4BEG[0] }),
    .FrameData({\Tile_X1Y1_FrameData_O[31] ,
    \Tile_X1Y1_FrameData_O[30] ,
    \Tile_X1Y1_FrameData_O[29] ,
    \Tile_X1Y1_FrameData_O[28] ,
    \Tile_X1Y1_FrameData_O[27] ,
    \Tile_X1Y1_FrameData_O[26] ,
    \Tile_X1Y1_FrameData_O[25] ,
    \Tile_X1Y1_FrameData_O[24] ,
    \Tile_X1Y1_FrameData_O[23] ,
    \Tile_X1Y1_FrameData_O[22] ,
    \Tile_X1Y1_FrameData_O[21] ,
    \Tile_X1Y1_FrameData_O[20] ,
    \Tile_X1Y1_FrameData_O[19] ,
    \Tile_X1Y1_FrameData_O[18] ,
    \Tile_X1Y1_FrameData_O[17] ,
    \Tile_X1Y1_FrameData_O[16] ,
    \Tile_X1Y1_FrameData_O[15] ,
    \Tile_X1Y1_FrameData_O[14] ,
    \Tile_X1Y1_FrameData_O[13] ,
    \Tile_X1Y1_FrameData_O[12] ,
    \Tile_X1Y1_FrameData_O[11] ,
    \Tile_X1Y1_FrameData_O[10] ,
    \Tile_X1Y1_FrameData_O[9] ,
    \Tile_X1Y1_FrameData_O[8] ,
    \Tile_X1Y1_FrameData_O[7] ,
    \Tile_X1Y1_FrameData_O[6] ,
    \Tile_X1Y1_FrameData_O[5] ,
    \Tile_X1Y1_FrameData_O[4] ,
    \Tile_X1Y1_FrameData_O[3] ,
    \Tile_X1Y1_FrameData_O[2] ,
    \Tile_X1Y1_FrameData_O[1] ,
    \Tile_X1Y1_FrameData_O[0] }),
    .FrameData_O({\Tile_X2Y1_FrameData_O[31] ,
    \Tile_X2Y1_FrameData_O[30] ,
    \Tile_X2Y1_FrameData_O[29] ,
    \Tile_X2Y1_FrameData_O[28] ,
    \Tile_X2Y1_FrameData_O[27] ,
    \Tile_X2Y1_FrameData_O[26] ,
    \Tile_X2Y1_FrameData_O[25] ,
    \Tile_X2Y1_FrameData_O[24] ,
    \Tile_X2Y1_FrameData_O[23] ,
    \Tile_X2Y1_FrameData_O[22] ,
    \Tile_X2Y1_FrameData_O[21] ,
    \Tile_X2Y1_FrameData_O[20] ,
    \Tile_X2Y1_FrameData_O[19] ,
    \Tile_X2Y1_FrameData_O[18] ,
    \Tile_X2Y1_FrameData_O[17] ,
    \Tile_X2Y1_FrameData_O[16] ,
    \Tile_X2Y1_FrameData_O[15] ,
    \Tile_X2Y1_FrameData_O[14] ,
    \Tile_X2Y1_FrameData_O[13] ,
    \Tile_X2Y1_FrameData_O[12] ,
    \Tile_X2Y1_FrameData_O[11] ,
    \Tile_X2Y1_FrameData_O[10] ,
    \Tile_X2Y1_FrameData_O[9] ,
    \Tile_X2Y1_FrameData_O[8] ,
    \Tile_X2Y1_FrameData_O[7] ,
    \Tile_X2Y1_FrameData_O[6] ,
    \Tile_X2Y1_FrameData_O[5] ,
    \Tile_X2Y1_FrameData_O[4] ,
    \Tile_X2Y1_FrameData_O[3] ,
    \Tile_X2Y1_FrameData_O[2] ,
    \Tile_X2Y1_FrameData_O[1] ,
    \Tile_X2Y1_FrameData_O[0] }),
    .FrameStrobe({\Tile_X2Y2_FrameStrobe_O[19] ,
    \Tile_X2Y2_FrameStrobe_O[18] ,
    \Tile_X2Y2_FrameStrobe_O[17] ,
    \Tile_X2Y2_FrameStrobe_O[16] ,
    \Tile_X2Y2_FrameStrobe_O[15] ,
    \Tile_X2Y2_FrameStrobe_O[14] ,
    \Tile_X2Y2_FrameStrobe_O[13] ,
    \Tile_X2Y2_FrameStrobe_O[12] ,
    \Tile_X2Y2_FrameStrobe_O[11] ,
    \Tile_X2Y2_FrameStrobe_O[10] ,
    \Tile_X2Y2_FrameStrobe_O[9] ,
    \Tile_X2Y2_FrameStrobe_O[8] ,
    \Tile_X2Y2_FrameStrobe_O[7] ,
    \Tile_X2Y2_FrameStrobe_O[6] ,
    \Tile_X2Y2_FrameStrobe_O[5] ,
    \Tile_X2Y2_FrameStrobe_O[4] ,
    \Tile_X2Y2_FrameStrobe_O[3] ,
    \Tile_X2Y2_FrameStrobe_O[2] ,
    \Tile_X2Y2_FrameStrobe_O[1] ,
    \Tile_X2Y2_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X2Y1_FrameStrobe_O[19] ,
    \Tile_X2Y1_FrameStrobe_O[18] ,
    \Tile_X2Y1_FrameStrobe_O[17] ,
    \Tile_X2Y1_FrameStrobe_O[16] ,
    \Tile_X2Y1_FrameStrobe_O[15] ,
    \Tile_X2Y1_FrameStrobe_O[14] ,
    \Tile_X2Y1_FrameStrobe_O[13] ,
    \Tile_X2Y1_FrameStrobe_O[12] ,
    \Tile_X2Y1_FrameStrobe_O[11] ,
    \Tile_X2Y1_FrameStrobe_O[10] ,
    \Tile_X2Y1_FrameStrobe_O[9] ,
    \Tile_X2Y1_FrameStrobe_O[8] ,
    \Tile_X2Y1_FrameStrobe_O[7] ,
    \Tile_X2Y1_FrameStrobe_O[6] ,
    \Tile_X2Y1_FrameStrobe_O[5] ,
    \Tile_X2Y1_FrameStrobe_O[4] ,
    \Tile_X2Y1_FrameStrobe_O[3] ,
    \Tile_X2Y1_FrameStrobe_O[2] ,
    \Tile_X2Y1_FrameStrobe_O[1] ,
    \Tile_X2Y1_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X2Y1_N1BEG[3] ,
    \Tile_X2Y1_N1BEG[2] ,
    \Tile_X2Y1_N1BEG[1] ,
    \Tile_X2Y1_N1BEG[0] }),
    .N1END({\Tile_X2Y2_N1BEG[3] ,
    \Tile_X2Y2_N1BEG[2] ,
    \Tile_X2Y2_N1BEG[1] ,
    \Tile_X2Y2_N1BEG[0] }),
    .N2BEG({\Tile_X2Y1_N2BEG[7] ,
    \Tile_X2Y1_N2BEG[6] ,
    \Tile_X2Y1_N2BEG[5] ,
    \Tile_X2Y1_N2BEG[4] ,
    \Tile_X2Y1_N2BEG[3] ,
    \Tile_X2Y1_N2BEG[2] ,
    \Tile_X2Y1_N2BEG[1] ,
    \Tile_X2Y1_N2BEG[0] }),
    .N2BEGb({\Tile_X2Y1_N2BEGb[7] ,
    \Tile_X2Y1_N2BEGb[6] ,
    \Tile_X2Y1_N2BEGb[5] ,
    \Tile_X2Y1_N2BEGb[4] ,
    \Tile_X2Y1_N2BEGb[3] ,
    \Tile_X2Y1_N2BEGb[2] ,
    \Tile_X2Y1_N2BEGb[1] ,
    \Tile_X2Y1_N2BEGb[0] }),
    .N2END({\Tile_X2Y2_N2BEGb[7] ,
    \Tile_X2Y2_N2BEGb[6] ,
    \Tile_X2Y2_N2BEGb[5] ,
    \Tile_X2Y2_N2BEGb[4] ,
    \Tile_X2Y2_N2BEGb[3] ,
    \Tile_X2Y2_N2BEGb[2] ,
    \Tile_X2Y2_N2BEGb[1] ,
    \Tile_X2Y2_N2BEGb[0] }),
    .N2MID({\Tile_X2Y2_N2BEG[7] ,
    \Tile_X2Y2_N2BEG[6] ,
    \Tile_X2Y2_N2BEG[5] ,
    \Tile_X2Y2_N2BEG[4] ,
    \Tile_X2Y2_N2BEG[3] ,
    \Tile_X2Y2_N2BEG[2] ,
    \Tile_X2Y2_N2BEG[1] ,
    \Tile_X2Y2_N2BEG[0] }),
    .N4BEG({\Tile_X2Y1_N4BEG[15] ,
    \Tile_X2Y1_N4BEG[14] ,
    \Tile_X2Y1_N4BEG[13] ,
    \Tile_X2Y1_N4BEG[12] ,
    \Tile_X2Y1_N4BEG[11] ,
    \Tile_X2Y1_N4BEG[10] ,
    \Tile_X2Y1_N4BEG[9] ,
    \Tile_X2Y1_N4BEG[8] ,
    \Tile_X2Y1_N4BEG[7] ,
    \Tile_X2Y1_N4BEG[6] ,
    \Tile_X2Y1_N4BEG[5] ,
    \Tile_X2Y1_N4BEG[4] ,
    \Tile_X2Y1_N4BEG[3] ,
    \Tile_X2Y1_N4BEG[2] ,
    \Tile_X2Y1_N4BEG[1] ,
    \Tile_X2Y1_N4BEG[0] }),
    .N4END({\Tile_X2Y2_N4BEG[15] ,
    \Tile_X2Y2_N4BEG[14] ,
    \Tile_X2Y2_N4BEG[13] ,
    \Tile_X2Y2_N4BEG[12] ,
    \Tile_X2Y2_N4BEG[11] ,
    \Tile_X2Y2_N4BEG[10] ,
    \Tile_X2Y2_N4BEG[9] ,
    \Tile_X2Y2_N4BEG[8] ,
    \Tile_X2Y2_N4BEG[7] ,
    \Tile_X2Y2_N4BEG[6] ,
    \Tile_X2Y2_N4BEG[5] ,
    \Tile_X2Y2_N4BEG[4] ,
    \Tile_X2Y2_N4BEG[3] ,
    \Tile_X2Y2_N4BEG[2] ,
    \Tile_X2Y2_N4BEG[1] ,
    \Tile_X2Y2_N4BEG[0] }),
    .NN4BEG({\Tile_X2Y1_NN4BEG[15] ,
    \Tile_X2Y1_NN4BEG[14] ,
    \Tile_X2Y1_NN4BEG[13] ,
    \Tile_X2Y1_NN4BEG[12] ,
    \Tile_X2Y1_NN4BEG[11] ,
    \Tile_X2Y1_NN4BEG[10] ,
    \Tile_X2Y1_NN4BEG[9] ,
    \Tile_X2Y1_NN4BEG[8] ,
    \Tile_X2Y1_NN4BEG[7] ,
    \Tile_X2Y1_NN4BEG[6] ,
    \Tile_X2Y1_NN4BEG[5] ,
    \Tile_X2Y1_NN4BEG[4] ,
    \Tile_X2Y1_NN4BEG[3] ,
    \Tile_X2Y1_NN4BEG[2] ,
    \Tile_X2Y1_NN4BEG[1] ,
    \Tile_X2Y1_NN4BEG[0] }),
    .NN4END({\Tile_X2Y2_NN4BEG[15] ,
    \Tile_X2Y2_NN4BEG[14] ,
    \Tile_X2Y2_NN4BEG[13] ,
    \Tile_X2Y2_NN4BEG[12] ,
    \Tile_X2Y2_NN4BEG[11] ,
    \Tile_X2Y2_NN4BEG[10] ,
    \Tile_X2Y2_NN4BEG[9] ,
    \Tile_X2Y2_NN4BEG[8] ,
    \Tile_X2Y2_NN4BEG[7] ,
    \Tile_X2Y2_NN4BEG[6] ,
    \Tile_X2Y2_NN4BEG[5] ,
    \Tile_X2Y2_NN4BEG[4] ,
    \Tile_X2Y2_NN4BEG[3] ,
    \Tile_X2Y2_NN4BEG[2] ,
    \Tile_X2Y2_NN4BEG[1] ,
    \Tile_X2Y2_NN4BEG[0] }),
    .S1BEG({\Tile_X2Y1_S1BEG[3] ,
    \Tile_X2Y1_S1BEG[2] ,
    \Tile_X2Y1_S1BEG[1] ,
    \Tile_X2Y1_S1BEG[0] }),
    .S1END({\Tile_X2Y0_S1BEG[3] ,
    \Tile_X2Y0_S1BEG[2] ,
    \Tile_X2Y0_S1BEG[1] ,
    \Tile_X2Y0_S1BEG[0] }),
    .S2BEG({\Tile_X2Y1_S2BEG[7] ,
    \Tile_X2Y1_S2BEG[6] ,
    \Tile_X2Y1_S2BEG[5] ,
    \Tile_X2Y1_S2BEG[4] ,
    \Tile_X2Y1_S2BEG[3] ,
    \Tile_X2Y1_S2BEG[2] ,
    \Tile_X2Y1_S2BEG[1] ,
    \Tile_X2Y1_S2BEG[0] }),
    .S2BEGb({\Tile_X2Y1_S2BEGb[7] ,
    \Tile_X2Y1_S2BEGb[6] ,
    \Tile_X2Y1_S2BEGb[5] ,
    \Tile_X2Y1_S2BEGb[4] ,
    \Tile_X2Y1_S2BEGb[3] ,
    \Tile_X2Y1_S2BEGb[2] ,
    \Tile_X2Y1_S2BEGb[1] ,
    \Tile_X2Y1_S2BEGb[0] }),
    .S2END({\Tile_X2Y0_S2BEGb[7] ,
    \Tile_X2Y0_S2BEGb[6] ,
    \Tile_X2Y0_S2BEGb[5] ,
    \Tile_X2Y0_S2BEGb[4] ,
    \Tile_X2Y0_S2BEGb[3] ,
    \Tile_X2Y0_S2BEGb[2] ,
    \Tile_X2Y0_S2BEGb[1] ,
    \Tile_X2Y0_S2BEGb[0] }),
    .S2MID({\Tile_X2Y0_S2BEG[7] ,
    \Tile_X2Y0_S2BEG[6] ,
    \Tile_X2Y0_S2BEG[5] ,
    \Tile_X2Y0_S2BEG[4] ,
    \Tile_X2Y0_S2BEG[3] ,
    \Tile_X2Y0_S2BEG[2] ,
    \Tile_X2Y0_S2BEG[1] ,
    \Tile_X2Y0_S2BEG[0] }),
    .S4BEG({\Tile_X2Y1_S4BEG[15] ,
    \Tile_X2Y1_S4BEG[14] ,
    \Tile_X2Y1_S4BEG[13] ,
    \Tile_X2Y1_S4BEG[12] ,
    \Tile_X2Y1_S4BEG[11] ,
    \Tile_X2Y1_S4BEG[10] ,
    \Tile_X2Y1_S4BEG[9] ,
    \Tile_X2Y1_S4BEG[8] ,
    \Tile_X2Y1_S4BEG[7] ,
    \Tile_X2Y1_S4BEG[6] ,
    \Tile_X2Y1_S4BEG[5] ,
    \Tile_X2Y1_S4BEG[4] ,
    \Tile_X2Y1_S4BEG[3] ,
    \Tile_X2Y1_S4BEG[2] ,
    \Tile_X2Y1_S4BEG[1] ,
    \Tile_X2Y1_S4BEG[0] }),
    .S4END({\Tile_X2Y0_S4BEG[15] ,
    \Tile_X2Y0_S4BEG[14] ,
    \Tile_X2Y0_S4BEG[13] ,
    \Tile_X2Y0_S4BEG[12] ,
    \Tile_X2Y0_S4BEG[11] ,
    \Tile_X2Y0_S4BEG[10] ,
    \Tile_X2Y0_S4BEG[9] ,
    \Tile_X2Y0_S4BEG[8] ,
    \Tile_X2Y0_S4BEG[7] ,
    \Tile_X2Y0_S4BEG[6] ,
    \Tile_X2Y0_S4BEG[5] ,
    \Tile_X2Y0_S4BEG[4] ,
    \Tile_X2Y0_S4BEG[3] ,
    \Tile_X2Y0_S4BEG[2] ,
    \Tile_X2Y0_S4BEG[1] ,
    \Tile_X2Y0_S4BEG[0] }),
    .SS4BEG({\Tile_X2Y1_SS4BEG[15] ,
    \Tile_X2Y1_SS4BEG[14] ,
    \Tile_X2Y1_SS4BEG[13] ,
    \Tile_X2Y1_SS4BEG[12] ,
    \Tile_X2Y1_SS4BEG[11] ,
    \Tile_X2Y1_SS4BEG[10] ,
    \Tile_X2Y1_SS4BEG[9] ,
    \Tile_X2Y1_SS4BEG[8] ,
    \Tile_X2Y1_SS4BEG[7] ,
    \Tile_X2Y1_SS4BEG[6] ,
    \Tile_X2Y1_SS4BEG[5] ,
    \Tile_X2Y1_SS4BEG[4] ,
    \Tile_X2Y1_SS4BEG[3] ,
    \Tile_X2Y1_SS4BEG[2] ,
    \Tile_X2Y1_SS4BEG[1] ,
    \Tile_X2Y1_SS4BEG[0] }),
    .SS4END({\Tile_X2Y0_SS4BEG[15] ,
    \Tile_X2Y0_SS4BEG[14] ,
    \Tile_X2Y0_SS4BEG[13] ,
    \Tile_X2Y0_SS4BEG[12] ,
    \Tile_X2Y0_SS4BEG[11] ,
    \Tile_X2Y0_SS4BEG[10] ,
    \Tile_X2Y0_SS4BEG[9] ,
    \Tile_X2Y0_SS4BEG[8] ,
    \Tile_X2Y0_SS4BEG[7] ,
    \Tile_X2Y0_SS4BEG[6] ,
    \Tile_X2Y0_SS4BEG[5] ,
    \Tile_X2Y0_SS4BEG[4] ,
    \Tile_X2Y0_SS4BEG[3] ,
    \Tile_X2Y0_SS4BEG[2] ,
    \Tile_X2Y0_SS4BEG[1] ,
    \Tile_X2Y0_SS4BEG[0] }),
    .W1BEG({\Tile_X2Y1_W1BEG[3] ,
    \Tile_X2Y1_W1BEG[2] ,
    \Tile_X2Y1_W1BEG[1] ,
    \Tile_X2Y1_W1BEG[0] }),
    .W1END({\Tile_X3Y1_W1BEG[3] ,
    \Tile_X3Y1_W1BEG[2] ,
    \Tile_X3Y1_W1BEG[1] ,
    \Tile_X3Y1_W1BEG[0] }),
    .W2BEG({\Tile_X2Y1_W2BEG[7] ,
    \Tile_X2Y1_W2BEG[6] ,
    \Tile_X2Y1_W2BEG[5] ,
    \Tile_X2Y1_W2BEG[4] ,
    \Tile_X2Y1_W2BEG[3] ,
    \Tile_X2Y1_W2BEG[2] ,
    \Tile_X2Y1_W2BEG[1] ,
    \Tile_X2Y1_W2BEG[0] }),
    .W2BEGb({\Tile_X2Y1_W2BEGb[7] ,
    \Tile_X2Y1_W2BEGb[6] ,
    \Tile_X2Y1_W2BEGb[5] ,
    \Tile_X2Y1_W2BEGb[4] ,
    \Tile_X2Y1_W2BEGb[3] ,
    \Tile_X2Y1_W2BEGb[2] ,
    \Tile_X2Y1_W2BEGb[1] ,
    \Tile_X2Y1_W2BEGb[0] }),
    .W2END({\Tile_X3Y1_W2BEGb[7] ,
    \Tile_X3Y1_W2BEGb[6] ,
    \Tile_X3Y1_W2BEGb[5] ,
    \Tile_X3Y1_W2BEGb[4] ,
    \Tile_X3Y1_W2BEGb[3] ,
    \Tile_X3Y1_W2BEGb[2] ,
    \Tile_X3Y1_W2BEGb[1] ,
    \Tile_X3Y1_W2BEGb[0] }),
    .W2MID({\Tile_X3Y1_W2BEG[7] ,
    \Tile_X3Y1_W2BEG[6] ,
    \Tile_X3Y1_W2BEG[5] ,
    \Tile_X3Y1_W2BEG[4] ,
    \Tile_X3Y1_W2BEG[3] ,
    \Tile_X3Y1_W2BEG[2] ,
    \Tile_X3Y1_W2BEG[1] ,
    \Tile_X3Y1_W2BEG[0] }),
    .W6BEG({\Tile_X2Y1_W6BEG[11] ,
    \Tile_X2Y1_W6BEG[10] ,
    \Tile_X2Y1_W6BEG[9] ,
    \Tile_X2Y1_W6BEG[8] ,
    \Tile_X2Y1_W6BEG[7] ,
    \Tile_X2Y1_W6BEG[6] ,
    \Tile_X2Y1_W6BEG[5] ,
    \Tile_X2Y1_W6BEG[4] ,
    \Tile_X2Y1_W6BEG[3] ,
    \Tile_X2Y1_W6BEG[2] ,
    \Tile_X2Y1_W6BEG[1] ,
    \Tile_X2Y1_W6BEG[0] }),
    .W6END({\Tile_X3Y1_W6BEG[11] ,
    \Tile_X3Y1_W6BEG[10] ,
    \Tile_X3Y1_W6BEG[9] ,
    \Tile_X3Y1_W6BEG[8] ,
    \Tile_X3Y1_W6BEG[7] ,
    \Tile_X3Y1_W6BEG[6] ,
    \Tile_X3Y1_W6BEG[5] ,
    \Tile_X3Y1_W6BEG[4] ,
    \Tile_X3Y1_W6BEG[3] ,
    \Tile_X3Y1_W6BEG[2] ,
    \Tile_X3Y1_W6BEG[1] ,
    \Tile_X3Y1_W6BEG[0] }),
    .WW4BEG({\Tile_X2Y1_WW4BEG[15] ,
    \Tile_X2Y1_WW4BEG[14] ,
    \Tile_X2Y1_WW4BEG[13] ,
    \Tile_X2Y1_WW4BEG[12] ,
    \Tile_X2Y1_WW4BEG[11] ,
    \Tile_X2Y1_WW4BEG[10] ,
    \Tile_X2Y1_WW4BEG[9] ,
    \Tile_X2Y1_WW4BEG[8] ,
    \Tile_X2Y1_WW4BEG[7] ,
    \Tile_X2Y1_WW4BEG[6] ,
    \Tile_X2Y1_WW4BEG[5] ,
    \Tile_X2Y1_WW4BEG[4] ,
    \Tile_X2Y1_WW4BEG[3] ,
    \Tile_X2Y1_WW4BEG[2] ,
    \Tile_X2Y1_WW4BEG[1] ,
    \Tile_X2Y1_WW4BEG[0] }),
    .WW4END({\Tile_X3Y1_WW4BEG[15] ,
    \Tile_X3Y1_WW4BEG[14] ,
    \Tile_X3Y1_WW4BEG[13] ,
    \Tile_X3Y1_WW4BEG[12] ,
    \Tile_X3Y1_WW4BEG[11] ,
    \Tile_X3Y1_WW4BEG[10] ,
    \Tile_X3Y1_WW4BEG[9] ,
    \Tile_X3Y1_WW4BEG[8] ,
    \Tile_X3Y1_WW4BEG[7] ,
    \Tile_X3Y1_WW4BEG[6] ,
    \Tile_X3Y1_WW4BEG[5] ,
    \Tile_X3Y1_WW4BEG[4] ,
    \Tile_X3Y1_WW4BEG[3] ,
    \Tile_X3Y1_WW4BEG[2] ,
    \Tile_X3Y1_WW4BEG[1] ,
    \Tile_X3Y1_WW4BEG[0] }));
 LUT4AB Tile_X2Y2_LUT4AB (.Ci(Tile_X2Y3_Co),
    .Co(Tile_X2Y2_Co),
    .UserCLK(Tile_X2Y3_UserCLKo),
    .UserCLKo(Tile_X2Y2_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X2Y2_E1BEG[3] ,
    \Tile_X2Y2_E1BEG[2] ,
    \Tile_X2Y2_E1BEG[1] ,
    \Tile_X2Y2_E1BEG[0] }),
    .E1END({\Tile_X1Y2_E1BEG[3] ,
    \Tile_X1Y2_E1BEG[2] ,
    \Tile_X1Y2_E1BEG[1] ,
    \Tile_X1Y2_E1BEG[0] }),
    .E2BEG({\Tile_X2Y2_E2BEG[7] ,
    \Tile_X2Y2_E2BEG[6] ,
    \Tile_X2Y2_E2BEG[5] ,
    \Tile_X2Y2_E2BEG[4] ,
    \Tile_X2Y2_E2BEG[3] ,
    \Tile_X2Y2_E2BEG[2] ,
    \Tile_X2Y2_E2BEG[1] ,
    \Tile_X2Y2_E2BEG[0] }),
    .E2BEGb({\Tile_X2Y2_E2BEGb[7] ,
    \Tile_X2Y2_E2BEGb[6] ,
    \Tile_X2Y2_E2BEGb[5] ,
    \Tile_X2Y2_E2BEGb[4] ,
    \Tile_X2Y2_E2BEGb[3] ,
    \Tile_X2Y2_E2BEGb[2] ,
    \Tile_X2Y2_E2BEGb[1] ,
    \Tile_X2Y2_E2BEGb[0] }),
    .E2END({\Tile_X1Y2_E2BEGb[7] ,
    \Tile_X1Y2_E2BEGb[6] ,
    \Tile_X1Y2_E2BEGb[5] ,
    \Tile_X1Y2_E2BEGb[4] ,
    \Tile_X1Y2_E2BEGb[3] ,
    \Tile_X1Y2_E2BEGb[2] ,
    \Tile_X1Y2_E2BEGb[1] ,
    \Tile_X1Y2_E2BEGb[0] }),
    .E2MID({\Tile_X1Y2_E2BEG[7] ,
    \Tile_X1Y2_E2BEG[6] ,
    \Tile_X1Y2_E2BEG[5] ,
    \Tile_X1Y2_E2BEG[4] ,
    \Tile_X1Y2_E2BEG[3] ,
    \Tile_X1Y2_E2BEG[2] ,
    \Tile_X1Y2_E2BEG[1] ,
    \Tile_X1Y2_E2BEG[0] }),
    .E6BEG({\Tile_X2Y2_E6BEG[11] ,
    \Tile_X2Y2_E6BEG[10] ,
    \Tile_X2Y2_E6BEG[9] ,
    \Tile_X2Y2_E6BEG[8] ,
    \Tile_X2Y2_E6BEG[7] ,
    \Tile_X2Y2_E6BEG[6] ,
    \Tile_X2Y2_E6BEG[5] ,
    \Tile_X2Y2_E6BEG[4] ,
    \Tile_X2Y2_E6BEG[3] ,
    \Tile_X2Y2_E6BEG[2] ,
    \Tile_X2Y2_E6BEG[1] ,
    \Tile_X2Y2_E6BEG[0] }),
    .E6END({\Tile_X1Y2_E6BEG[11] ,
    \Tile_X1Y2_E6BEG[10] ,
    \Tile_X1Y2_E6BEG[9] ,
    \Tile_X1Y2_E6BEG[8] ,
    \Tile_X1Y2_E6BEG[7] ,
    \Tile_X1Y2_E6BEG[6] ,
    \Tile_X1Y2_E6BEG[5] ,
    \Tile_X1Y2_E6BEG[4] ,
    \Tile_X1Y2_E6BEG[3] ,
    \Tile_X1Y2_E6BEG[2] ,
    \Tile_X1Y2_E6BEG[1] ,
    \Tile_X1Y2_E6BEG[0] }),
    .EE4BEG({\Tile_X2Y2_EE4BEG[15] ,
    \Tile_X2Y2_EE4BEG[14] ,
    \Tile_X2Y2_EE4BEG[13] ,
    \Tile_X2Y2_EE4BEG[12] ,
    \Tile_X2Y2_EE4BEG[11] ,
    \Tile_X2Y2_EE4BEG[10] ,
    \Tile_X2Y2_EE4BEG[9] ,
    \Tile_X2Y2_EE4BEG[8] ,
    \Tile_X2Y2_EE4BEG[7] ,
    \Tile_X2Y2_EE4BEG[6] ,
    \Tile_X2Y2_EE4BEG[5] ,
    \Tile_X2Y2_EE4BEG[4] ,
    \Tile_X2Y2_EE4BEG[3] ,
    \Tile_X2Y2_EE4BEG[2] ,
    \Tile_X2Y2_EE4BEG[1] ,
    \Tile_X2Y2_EE4BEG[0] }),
    .EE4END({\Tile_X1Y2_EE4BEG[15] ,
    \Tile_X1Y2_EE4BEG[14] ,
    \Tile_X1Y2_EE4BEG[13] ,
    \Tile_X1Y2_EE4BEG[12] ,
    \Tile_X1Y2_EE4BEG[11] ,
    \Tile_X1Y2_EE4BEG[10] ,
    \Tile_X1Y2_EE4BEG[9] ,
    \Tile_X1Y2_EE4BEG[8] ,
    \Tile_X1Y2_EE4BEG[7] ,
    \Tile_X1Y2_EE4BEG[6] ,
    \Tile_X1Y2_EE4BEG[5] ,
    \Tile_X1Y2_EE4BEG[4] ,
    \Tile_X1Y2_EE4BEG[3] ,
    \Tile_X1Y2_EE4BEG[2] ,
    \Tile_X1Y2_EE4BEG[1] ,
    \Tile_X1Y2_EE4BEG[0] }),
    .FrameData({\Tile_X1Y2_FrameData_O[31] ,
    \Tile_X1Y2_FrameData_O[30] ,
    \Tile_X1Y2_FrameData_O[29] ,
    \Tile_X1Y2_FrameData_O[28] ,
    \Tile_X1Y2_FrameData_O[27] ,
    \Tile_X1Y2_FrameData_O[26] ,
    \Tile_X1Y2_FrameData_O[25] ,
    \Tile_X1Y2_FrameData_O[24] ,
    \Tile_X1Y2_FrameData_O[23] ,
    \Tile_X1Y2_FrameData_O[22] ,
    \Tile_X1Y2_FrameData_O[21] ,
    \Tile_X1Y2_FrameData_O[20] ,
    \Tile_X1Y2_FrameData_O[19] ,
    \Tile_X1Y2_FrameData_O[18] ,
    \Tile_X1Y2_FrameData_O[17] ,
    \Tile_X1Y2_FrameData_O[16] ,
    \Tile_X1Y2_FrameData_O[15] ,
    \Tile_X1Y2_FrameData_O[14] ,
    \Tile_X1Y2_FrameData_O[13] ,
    \Tile_X1Y2_FrameData_O[12] ,
    \Tile_X1Y2_FrameData_O[11] ,
    \Tile_X1Y2_FrameData_O[10] ,
    \Tile_X1Y2_FrameData_O[9] ,
    \Tile_X1Y2_FrameData_O[8] ,
    \Tile_X1Y2_FrameData_O[7] ,
    \Tile_X1Y2_FrameData_O[6] ,
    \Tile_X1Y2_FrameData_O[5] ,
    \Tile_X1Y2_FrameData_O[4] ,
    \Tile_X1Y2_FrameData_O[3] ,
    \Tile_X1Y2_FrameData_O[2] ,
    \Tile_X1Y2_FrameData_O[1] ,
    \Tile_X1Y2_FrameData_O[0] }),
    .FrameData_O({\Tile_X2Y2_FrameData_O[31] ,
    \Tile_X2Y2_FrameData_O[30] ,
    \Tile_X2Y2_FrameData_O[29] ,
    \Tile_X2Y2_FrameData_O[28] ,
    \Tile_X2Y2_FrameData_O[27] ,
    \Tile_X2Y2_FrameData_O[26] ,
    \Tile_X2Y2_FrameData_O[25] ,
    \Tile_X2Y2_FrameData_O[24] ,
    \Tile_X2Y2_FrameData_O[23] ,
    \Tile_X2Y2_FrameData_O[22] ,
    \Tile_X2Y2_FrameData_O[21] ,
    \Tile_X2Y2_FrameData_O[20] ,
    \Tile_X2Y2_FrameData_O[19] ,
    \Tile_X2Y2_FrameData_O[18] ,
    \Tile_X2Y2_FrameData_O[17] ,
    \Tile_X2Y2_FrameData_O[16] ,
    \Tile_X2Y2_FrameData_O[15] ,
    \Tile_X2Y2_FrameData_O[14] ,
    \Tile_X2Y2_FrameData_O[13] ,
    \Tile_X2Y2_FrameData_O[12] ,
    \Tile_X2Y2_FrameData_O[11] ,
    \Tile_X2Y2_FrameData_O[10] ,
    \Tile_X2Y2_FrameData_O[9] ,
    \Tile_X2Y2_FrameData_O[8] ,
    \Tile_X2Y2_FrameData_O[7] ,
    \Tile_X2Y2_FrameData_O[6] ,
    \Tile_X2Y2_FrameData_O[5] ,
    \Tile_X2Y2_FrameData_O[4] ,
    \Tile_X2Y2_FrameData_O[3] ,
    \Tile_X2Y2_FrameData_O[2] ,
    \Tile_X2Y2_FrameData_O[1] ,
    \Tile_X2Y2_FrameData_O[0] }),
    .FrameStrobe({\Tile_X2Y3_FrameStrobe_O[19] ,
    \Tile_X2Y3_FrameStrobe_O[18] ,
    \Tile_X2Y3_FrameStrobe_O[17] ,
    \Tile_X2Y3_FrameStrobe_O[16] ,
    \Tile_X2Y3_FrameStrobe_O[15] ,
    \Tile_X2Y3_FrameStrobe_O[14] ,
    \Tile_X2Y3_FrameStrobe_O[13] ,
    \Tile_X2Y3_FrameStrobe_O[12] ,
    \Tile_X2Y3_FrameStrobe_O[11] ,
    \Tile_X2Y3_FrameStrobe_O[10] ,
    \Tile_X2Y3_FrameStrobe_O[9] ,
    \Tile_X2Y3_FrameStrobe_O[8] ,
    \Tile_X2Y3_FrameStrobe_O[7] ,
    \Tile_X2Y3_FrameStrobe_O[6] ,
    \Tile_X2Y3_FrameStrobe_O[5] ,
    \Tile_X2Y3_FrameStrobe_O[4] ,
    \Tile_X2Y3_FrameStrobe_O[3] ,
    \Tile_X2Y3_FrameStrobe_O[2] ,
    \Tile_X2Y3_FrameStrobe_O[1] ,
    \Tile_X2Y3_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X2Y2_FrameStrobe_O[19] ,
    \Tile_X2Y2_FrameStrobe_O[18] ,
    \Tile_X2Y2_FrameStrobe_O[17] ,
    \Tile_X2Y2_FrameStrobe_O[16] ,
    \Tile_X2Y2_FrameStrobe_O[15] ,
    \Tile_X2Y2_FrameStrobe_O[14] ,
    \Tile_X2Y2_FrameStrobe_O[13] ,
    \Tile_X2Y2_FrameStrobe_O[12] ,
    \Tile_X2Y2_FrameStrobe_O[11] ,
    \Tile_X2Y2_FrameStrobe_O[10] ,
    \Tile_X2Y2_FrameStrobe_O[9] ,
    \Tile_X2Y2_FrameStrobe_O[8] ,
    \Tile_X2Y2_FrameStrobe_O[7] ,
    \Tile_X2Y2_FrameStrobe_O[6] ,
    \Tile_X2Y2_FrameStrobe_O[5] ,
    \Tile_X2Y2_FrameStrobe_O[4] ,
    \Tile_X2Y2_FrameStrobe_O[3] ,
    \Tile_X2Y2_FrameStrobe_O[2] ,
    \Tile_X2Y2_FrameStrobe_O[1] ,
    \Tile_X2Y2_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X2Y2_N1BEG[3] ,
    \Tile_X2Y2_N1BEG[2] ,
    \Tile_X2Y2_N1BEG[1] ,
    \Tile_X2Y2_N1BEG[0] }),
    .N1END({\Tile_X2Y3_N1BEG[3] ,
    \Tile_X2Y3_N1BEG[2] ,
    \Tile_X2Y3_N1BEG[1] ,
    \Tile_X2Y3_N1BEG[0] }),
    .N2BEG({\Tile_X2Y2_N2BEG[7] ,
    \Tile_X2Y2_N2BEG[6] ,
    \Tile_X2Y2_N2BEG[5] ,
    \Tile_X2Y2_N2BEG[4] ,
    \Tile_X2Y2_N2BEG[3] ,
    \Tile_X2Y2_N2BEG[2] ,
    \Tile_X2Y2_N2BEG[1] ,
    \Tile_X2Y2_N2BEG[0] }),
    .N2BEGb({\Tile_X2Y2_N2BEGb[7] ,
    \Tile_X2Y2_N2BEGb[6] ,
    \Tile_X2Y2_N2BEGb[5] ,
    \Tile_X2Y2_N2BEGb[4] ,
    \Tile_X2Y2_N2BEGb[3] ,
    \Tile_X2Y2_N2BEGb[2] ,
    \Tile_X2Y2_N2BEGb[1] ,
    \Tile_X2Y2_N2BEGb[0] }),
    .N2END({\Tile_X2Y3_N2BEGb[7] ,
    \Tile_X2Y3_N2BEGb[6] ,
    \Tile_X2Y3_N2BEGb[5] ,
    \Tile_X2Y3_N2BEGb[4] ,
    \Tile_X2Y3_N2BEGb[3] ,
    \Tile_X2Y3_N2BEGb[2] ,
    \Tile_X2Y3_N2BEGb[1] ,
    \Tile_X2Y3_N2BEGb[0] }),
    .N2MID({\Tile_X2Y3_N2BEG[7] ,
    \Tile_X2Y3_N2BEG[6] ,
    \Tile_X2Y3_N2BEG[5] ,
    \Tile_X2Y3_N2BEG[4] ,
    \Tile_X2Y3_N2BEG[3] ,
    \Tile_X2Y3_N2BEG[2] ,
    \Tile_X2Y3_N2BEG[1] ,
    \Tile_X2Y3_N2BEG[0] }),
    .N4BEG({\Tile_X2Y2_N4BEG[15] ,
    \Tile_X2Y2_N4BEG[14] ,
    \Tile_X2Y2_N4BEG[13] ,
    \Tile_X2Y2_N4BEG[12] ,
    \Tile_X2Y2_N4BEG[11] ,
    \Tile_X2Y2_N4BEG[10] ,
    \Tile_X2Y2_N4BEG[9] ,
    \Tile_X2Y2_N4BEG[8] ,
    \Tile_X2Y2_N4BEG[7] ,
    \Tile_X2Y2_N4BEG[6] ,
    \Tile_X2Y2_N4BEG[5] ,
    \Tile_X2Y2_N4BEG[4] ,
    \Tile_X2Y2_N4BEG[3] ,
    \Tile_X2Y2_N4BEG[2] ,
    \Tile_X2Y2_N4BEG[1] ,
    \Tile_X2Y2_N4BEG[0] }),
    .N4END({\Tile_X2Y3_N4BEG[15] ,
    \Tile_X2Y3_N4BEG[14] ,
    \Tile_X2Y3_N4BEG[13] ,
    \Tile_X2Y3_N4BEG[12] ,
    \Tile_X2Y3_N4BEG[11] ,
    \Tile_X2Y3_N4BEG[10] ,
    \Tile_X2Y3_N4BEG[9] ,
    \Tile_X2Y3_N4BEG[8] ,
    \Tile_X2Y3_N4BEG[7] ,
    \Tile_X2Y3_N4BEG[6] ,
    \Tile_X2Y3_N4BEG[5] ,
    \Tile_X2Y3_N4BEG[4] ,
    \Tile_X2Y3_N4BEG[3] ,
    \Tile_X2Y3_N4BEG[2] ,
    \Tile_X2Y3_N4BEG[1] ,
    \Tile_X2Y3_N4BEG[0] }),
    .NN4BEG({\Tile_X2Y2_NN4BEG[15] ,
    \Tile_X2Y2_NN4BEG[14] ,
    \Tile_X2Y2_NN4BEG[13] ,
    \Tile_X2Y2_NN4BEG[12] ,
    \Tile_X2Y2_NN4BEG[11] ,
    \Tile_X2Y2_NN4BEG[10] ,
    \Tile_X2Y2_NN4BEG[9] ,
    \Tile_X2Y2_NN4BEG[8] ,
    \Tile_X2Y2_NN4BEG[7] ,
    \Tile_X2Y2_NN4BEG[6] ,
    \Tile_X2Y2_NN4BEG[5] ,
    \Tile_X2Y2_NN4BEG[4] ,
    \Tile_X2Y2_NN4BEG[3] ,
    \Tile_X2Y2_NN4BEG[2] ,
    \Tile_X2Y2_NN4BEG[1] ,
    \Tile_X2Y2_NN4BEG[0] }),
    .NN4END({\Tile_X2Y3_NN4BEG[15] ,
    \Tile_X2Y3_NN4BEG[14] ,
    \Tile_X2Y3_NN4BEG[13] ,
    \Tile_X2Y3_NN4BEG[12] ,
    \Tile_X2Y3_NN4BEG[11] ,
    \Tile_X2Y3_NN4BEG[10] ,
    \Tile_X2Y3_NN4BEG[9] ,
    \Tile_X2Y3_NN4BEG[8] ,
    \Tile_X2Y3_NN4BEG[7] ,
    \Tile_X2Y3_NN4BEG[6] ,
    \Tile_X2Y3_NN4BEG[5] ,
    \Tile_X2Y3_NN4BEG[4] ,
    \Tile_X2Y3_NN4BEG[3] ,
    \Tile_X2Y3_NN4BEG[2] ,
    \Tile_X2Y3_NN4BEG[1] ,
    \Tile_X2Y3_NN4BEG[0] }),
    .S1BEG({\Tile_X2Y2_S1BEG[3] ,
    \Tile_X2Y2_S1BEG[2] ,
    \Tile_X2Y2_S1BEG[1] ,
    \Tile_X2Y2_S1BEG[0] }),
    .S1END({\Tile_X2Y1_S1BEG[3] ,
    \Tile_X2Y1_S1BEG[2] ,
    \Tile_X2Y1_S1BEG[1] ,
    \Tile_X2Y1_S1BEG[0] }),
    .S2BEG({\Tile_X2Y2_S2BEG[7] ,
    \Tile_X2Y2_S2BEG[6] ,
    \Tile_X2Y2_S2BEG[5] ,
    \Tile_X2Y2_S2BEG[4] ,
    \Tile_X2Y2_S2BEG[3] ,
    \Tile_X2Y2_S2BEG[2] ,
    \Tile_X2Y2_S2BEG[1] ,
    \Tile_X2Y2_S2BEG[0] }),
    .S2BEGb({\Tile_X2Y2_S2BEGb[7] ,
    \Tile_X2Y2_S2BEGb[6] ,
    \Tile_X2Y2_S2BEGb[5] ,
    \Tile_X2Y2_S2BEGb[4] ,
    \Tile_X2Y2_S2BEGb[3] ,
    \Tile_X2Y2_S2BEGb[2] ,
    \Tile_X2Y2_S2BEGb[1] ,
    \Tile_X2Y2_S2BEGb[0] }),
    .S2END({\Tile_X2Y1_S2BEGb[7] ,
    \Tile_X2Y1_S2BEGb[6] ,
    \Tile_X2Y1_S2BEGb[5] ,
    \Tile_X2Y1_S2BEGb[4] ,
    \Tile_X2Y1_S2BEGb[3] ,
    \Tile_X2Y1_S2BEGb[2] ,
    \Tile_X2Y1_S2BEGb[1] ,
    \Tile_X2Y1_S2BEGb[0] }),
    .S2MID({\Tile_X2Y1_S2BEG[7] ,
    \Tile_X2Y1_S2BEG[6] ,
    \Tile_X2Y1_S2BEG[5] ,
    \Tile_X2Y1_S2BEG[4] ,
    \Tile_X2Y1_S2BEG[3] ,
    \Tile_X2Y1_S2BEG[2] ,
    \Tile_X2Y1_S2BEG[1] ,
    \Tile_X2Y1_S2BEG[0] }),
    .S4BEG({\Tile_X2Y2_S4BEG[15] ,
    \Tile_X2Y2_S4BEG[14] ,
    \Tile_X2Y2_S4BEG[13] ,
    \Tile_X2Y2_S4BEG[12] ,
    \Tile_X2Y2_S4BEG[11] ,
    \Tile_X2Y2_S4BEG[10] ,
    \Tile_X2Y2_S4BEG[9] ,
    \Tile_X2Y2_S4BEG[8] ,
    \Tile_X2Y2_S4BEG[7] ,
    \Tile_X2Y2_S4BEG[6] ,
    \Tile_X2Y2_S4BEG[5] ,
    \Tile_X2Y2_S4BEG[4] ,
    \Tile_X2Y2_S4BEG[3] ,
    \Tile_X2Y2_S4BEG[2] ,
    \Tile_X2Y2_S4BEG[1] ,
    \Tile_X2Y2_S4BEG[0] }),
    .S4END({\Tile_X2Y1_S4BEG[15] ,
    \Tile_X2Y1_S4BEG[14] ,
    \Tile_X2Y1_S4BEG[13] ,
    \Tile_X2Y1_S4BEG[12] ,
    \Tile_X2Y1_S4BEG[11] ,
    \Tile_X2Y1_S4BEG[10] ,
    \Tile_X2Y1_S4BEG[9] ,
    \Tile_X2Y1_S4BEG[8] ,
    \Tile_X2Y1_S4BEG[7] ,
    \Tile_X2Y1_S4BEG[6] ,
    \Tile_X2Y1_S4BEG[5] ,
    \Tile_X2Y1_S4BEG[4] ,
    \Tile_X2Y1_S4BEG[3] ,
    \Tile_X2Y1_S4BEG[2] ,
    \Tile_X2Y1_S4BEG[1] ,
    \Tile_X2Y1_S4BEG[0] }),
    .SS4BEG({\Tile_X2Y2_SS4BEG[15] ,
    \Tile_X2Y2_SS4BEG[14] ,
    \Tile_X2Y2_SS4BEG[13] ,
    \Tile_X2Y2_SS4BEG[12] ,
    \Tile_X2Y2_SS4BEG[11] ,
    \Tile_X2Y2_SS4BEG[10] ,
    \Tile_X2Y2_SS4BEG[9] ,
    \Tile_X2Y2_SS4BEG[8] ,
    \Tile_X2Y2_SS4BEG[7] ,
    \Tile_X2Y2_SS4BEG[6] ,
    \Tile_X2Y2_SS4BEG[5] ,
    \Tile_X2Y2_SS4BEG[4] ,
    \Tile_X2Y2_SS4BEG[3] ,
    \Tile_X2Y2_SS4BEG[2] ,
    \Tile_X2Y2_SS4BEG[1] ,
    \Tile_X2Y2_SS4BEG[0] }),
    .SS4END({\Tile_X2Y1_SS4BEG[15] ,
    \Tile_X2Y1_SS4BEG[14] ,
    \Tile_X2Y1_SS4BEG[13] ,
    \Tile_X2Y1_SS4BEG[12] ,
    \Tile_X2Y1_SS4BEG[11] ,
    \Tile_X2Y1_SS4BEG[10] ,
    \Tile_X2Y1_SS4BEG[9] ,
    \Tile_X2Y1_SS4BEG[8] ,
    \Tile_X2Y1_SS4BEG[7] ,
    \Tile_X2Y1_SS4BEG[6] ,
    \Tile_X2Y1_SS4BEG[5] ,
    \Tile_X2Y1_SS4BEG[4] ,
    \Tile_X2Y1_SS4BEG[3] ,
    \Tile_X2Y1_SS4BEG[2] ,
    \Tile_X2Y1_SS4BEG[1] ,
    \Tile_X2Y1_SS4BEG[0] }),
    .W1BEG({\Tile_X2Y2_W1BEG[3] ,
    \Tile_X2Y2_W1BEG[2] ,
    \Tile_X2Y2_W1BEG[1] ,
    \Tile_X2Y2_W1BEG[0] }),
    .W1END({\Tile_X3Y2_W1BEG[3] ,
    \Tile_X3Y2_W1BEG[2] ,
    \Tile_X3Y2_W1BEG[1] ,
    \Tile_X3Y2_W1BEG[0] }),
    .W2BEG({\Tile_X2Y2_W2BEG[7] ,
    \Tile_X2Y2_W2BEG[6] ,
    \Tile_X2Y2_W2BEG[5] ,
    \Tile_X2Y2_W2BEG[4] ,
    \Tile_X2Y2_W2BEG[3] ,
    \Tile_X2Y2_W2BEG[2] ,
    \Tile_X2Y2_W2BEG[1] ,
    \Tile_X2Y2_W2BEG[0] }),
    .W2BEGb({\Tile_X2Y2_W2BEGb[7] ,
    \Tile_X2Y2_W2BEGb[6] ,
    \Tile_X2Y2_W2BEGb[5] ,
    \Tile_X2Y2_W2BEGb[4] ,
    \Tile_X2Y2_W2BEGb[3] ,
    \Tile_X2Y2_W2BEGb[2] ,
    \Tile_X2Y2_W2BEGb[1] ,
    \Tile_X2Y2_W2BEGb[0] }),
    .W2END({\Tile_X3Y2_W2BEGb[7] ,
    \Tile_X3Y2_W2BEGb[6] ,
    \Tile_X3Y2_W2BEGb[5] ,
    \Tile_X3Y2_W2BEGb[4] ,
    \Tile_X3Y2_W2BEGb[3] ,
    \Tile_X3Y2_W2BEGb[2] ,
    \Tile_X3Y2_W2BEGb[1] ,
    \Tile_X3Y2_W2BEGb[0] }),
    .W2MID({\Tile_X3Y2_W2BEG[7] ,
    \Tile_X3Y2_W2BEG[6] ,
    \Tile_X3Y2_W2BEG[5] ,
    \Tile_X3Y2_W2BEG[4] ,
    \Tile_X3Y2_W2BEG[3] ,
    \Tile_X3Y2_W2BEG[2] ,
    \Tile_X3Y2_W2BEG[1] ,
    \Tile_X3Y2_W2BEG[0] }),
    .W6BEG({\Tile_X2Y2_W6BEG[11] ,
    \Tile_X2Y2_W6BEG[10] ,
    \Tile_X2Y2_W6BEG[9] ,
    \Tile_X2Y2_W6BEG[8] ,
    \Tile_X2Y2_W6BEG[7] ,
    \Tile_X2Y2_W6BEG[6] ,
    \Tile_X2Y2_W6BEG[5] ,
    \Tile_X2Y2_W6BEG[4] ,
    \Tile_X2Y2_W6BEG[3] ,
    \Tile_X2Y2_W6BEG[2] ,
    \Tile_X2Y2_W6BEG[1] ,
    \Tile_X2Y2_W6BEG[0] }),
    .W6END({\Tile_X3Y2_W6BEG[11] ,
    \Tile_X3Y2_W6BEG[10] ,
    \Tile_X3Y2_W6BEG[9] ,
    \Tile_X3Y2_W6BEG[8] ,
    \Tile_X3Y2_W6BEG[7] ,
    \Tile_X3Y2_W6BEG[6] ,
    \Tile_X3Y2_W6BEG[5] ,
    \Tile_X3Y2_W6BEG[4] ,
    \Tile_X3Y2_W6BEG[3] ,
    \Tile_X3Y2_W6BEG[2] ,
    \Tile_X3Y2_W6BEG[1] ,
    \Tile_X3Y2_W6BEG[0] }),
    .WW4BEG({\Tile_X2Y2_WW4BEG[15] ,
    \Tile_X2Y2_WW4BEG[14] ,
    \Tile_X2Y2_WW4BEG[13] ,
    \Tile_X2Y2_WW4BEG[12] ,
    \Tile_X2Y2_WW4BEG[11] ,
    \Tile_X2Y2_WW4BEG[10] ,
    \Tile_X2Y2_WW4BEG[9] ,
    \Tile_X2Y2_WW4BEG[8] ,
    \Tile_X2Y2_WW4BEG[7] ,
    \Tile_X2Y2_WW4BEG[6] ,
    \Tile_X2Y2_WW4BEG[5] ,
    \Tile_X2Y2_WW4BEG[4] ,
    \Tile_X2Y2_WW4BEG[3] ,
    \Tile_X2Y2_WW4BEG[2] ,
    \Tile_X2Y2_WW4BEG[1] ,
    \Tile_X2Y2_WW4BEG[0] }),
    .WW4END({\Tile_X3Y2_WW4BEG[15] ,
    \Tile_X3Y2_WW4BEG[14] ,
    \Tile_X3Y2_WW4BEG[13] ,
    \Tile_X3Y2_WW4BEG[12] ,
    \Tile_X3Y2_WW4BEG[11] ,
    \Tile_X3Y2_WW4BEG[10] ,
    \Tile_X3Y2_WW4BEG[9] ,
    \Tile_X3Y2_WW4BEG[8] ,
    \Tile_X3Y2_WW4BEG[7] ,
    \Tile_X3Y2_WW4BEG[6] ,
    \Tile_X3Y2_WW4BEG[5] ,
    \Tile_X3Y2_WW4BEG[4] ,
    \Tile_X3Y2_WW4BEG[3] ,
    \Tile_X3Y2_WW4BEG[2] ,
    \Tile_X3Y2_WW4BEG[1] ,
    \Tile_X3Y2_WW4BEG[0] }));
 LUT4AB Tile_X2Y3_LUT4AB (.Ci(Tile_X2Y4_Co),
    .Co(Tile_X2Y3_Co),
    .UserCLK(Tile_X2Y4_UserCLKo),
    .UserCLKo(Tile_X2Y3_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X2Y3_E1BEG[3] ,
    \Tile_X2Y3_E1BEG[2] ,
    \Tile_X2Y3_E1BEG[1] ,
    \Tile_X2Y3_E1BEG[0] }),
    .E1END({\Tile_X1Y3_E1BEG[3] ,
    \Tile_X1Y3_E1BEG[2] ,
    \Tile_X1Y3_E1BEG[1] ,
    \Tile_X1Y3_E1BEG[0] }),
    .E2BEG({\Tile_X2Y3_E2BEG[7] ,
    \Tile_X2Y3_E2BEG[6] ,
    \Tile_X2Y3_E2BEG[5] ,
    \Tile_X2Y3_E2BEG[4] ,
    \Tile_X2Y3_E2BEG[3] ,
    \Tile_X2Y3_E2BEG[2] ,
    \Tile_X2Y3_E2BEG[1] ,
    \Tile_X2Y3_E2BEG[0] }),
    .E2BEGb({\Tile_X2Y3_E2BEGb[7] ,
    \Tile_X2Y3_E2BEGb[6] ,
    \Tile_X2Y3_E2BEGb[5] ,
    \Tile_X2Y3_E2BEGb[4] ,
    \Tile_X2Y3_E2BEGb[3] ,
    \Tile_X2Y3_E2BEGb[2] ,
    \Tile_X2Y3_E2BEGb[1] ,
    \Tile_X2Y3_E2BEGb[0] }),
    .E2END({\Tile_X1Y3_E2BEGb[7] ,
    \Tile_X1Y3_E2BEGb[6] ,
    \Tile_X1Y3_E2BEGb[5] ,
    \Tile_X1Y3_E2BEGb[4] ,
    \Tile_X1Y3_E2BEGb[3] ,
    \Tile_X1Y3_E2BEGb[2] ,
    \Tile_X1Y3_E2BEGb[1] ,
    \Tile_X1Y3_E2BEGb[0] }),
    .E2MID({\Tile_X1Y3_E2BEG[7] ,
    \Tile_X1Y3_E2BEG[6] ,
    \Tile_X1Y3_E2BEG[5] ,
    \Tile_X1Y3_E2BEG[4] ,
    \Tile_X1Y3_E2BEG[3] ,
    \Tile_X1Y3_E2BEG[2] ,
    \Tile_X1Y3_E2BEG[1] ,
    \Tile_X1Y3_E2BEG[0] }),
    .E6BEG({\Tile_X2Y3_E6BEG[11] ,
    \Tile_X2Y3_E6BEG[10] ,
    \Tile_X2Y3_E6BEG[9] ,
    \Tile_X2Y3_E6BEG[8] ,
    \Tile_X2Y3_E6BEG[7] ,
    \Tile_X2Y3_E6BEG[6] ,
    \Tile_X2Y3_E6BEG[5] ,
    \Tile_X2Y3_E6BEG[4] ,
    \Tile_X2Y3_E6BEG[3] ,
    \Tile_X2Y3_E6BEG[2] ,
    \Tile_X2Y3_E6BEG[1] ,
    \Tile_X2Y3_E6BEG[0] }),
    .E6END({\Tile_X1Y3_E6BEG[11] ,
    \Tile_X1Y3_E6BEG[10] ,
    \Tile_X1Y3_E6BEG[9] ,
    \Tile_X1Y3_E6BEG[8] ,
    \Tile_X1Y3_E6BEG[7] ,
    \Tile_X1Y3_E6BEG[6] ,
    \Tile_X1Y3_E6BEG[5] ,
    \Tile_X1Y3_E6BEG[4] ,
    \Tile_X1Y3_E6BEG[3] ,
    \Tile_X1Y3_E6BEG[2] ,
    \Tile_X1Y3_E6BEG[1] ,
    \Tile_X1Y3_E6BEG[0] }),
    .EE4BEG({\Tile_X2Y3_EE4BEG[15] ,
    \Tile_X2Y3_EE4BEG[14] ,
    \Tile_X2Y3_EE4BEG[13] ,
    \Tile_X2Y3_EE4BEG[12] ,
    \Tile_X2Y3_EE4BEG[11] ,
    \Tile_X2Y3_EE4BEG[10] ,
    \Tile_X2Y3_EE4BEG[9] ,
    \Tile_X2Y3_EE4BEG[8] ,
    \Tile_X2Y3_EE4BEG[7] ,
    \Tile_X2Y3_EE4BEG[6] ,
    \Tile_X2Y3_EE4BEG[5] ,
    \Tile_X2Y3_EE4BEG[4] ,
    \Tile_X2Y3_EE4BEG[3] ,
    \Tile_X2Y3_EE4BEG[2] ,
    \Tile_X2Y3_EE4BEG[1] ,
    \Tile_X2Y3_EE4BEG[0] }),
    .EE4END({\Tile_X1Y3_EE4BEG[15] ,
    \Tile_X1Y3_EE4BEG[14] ,
    \Tile_X1Y3_EE4BEG[13] ,
    \Tile_X1Y3_EE4BEG[12] ,
    \Tile_X1Y3_EE4BEG[11] ,
    \Tile_X1Y3_EE4BEG[10] ,
    \Tile_X1Y3_EE4BEG[9] ,
    \Tile_X1Y3_EE4BEG[8] ,
    \Tile_X1Y3_EE4BEG[7] ,
    \Tile_X1Y3_EE4BEG[6] ,
    \Tile_X1Y3_EE4BEG[5] ,
    \Tile_X1Y3_EE4BEG[4] ,
    \Tile_X1Y3_EE4BEG[3] ,
    \Tile_X1Y3_EE4BEG[2] ,
    \Tile_X1Y3_EE4BEG[1] ,
    \Tile_X1Y3_EE4BEG[0] }),
    .FrameData({\Tile_X1Y3_FrameData_O[31] ,
    \Tile_X1Y3_FrameData_O[30] ,
    \Tile_X1Y3_FrameData_O[29] ,
    \Tile_X1Y3_FrameData_O[28] ,
    \Tile_X1Y3_FrameData_O[27] ,
    \Tile_X1Y3_FrameData_O[26] ,
    \Tile_X1Y3_FrameData_O[25] ,
    \Tile_X1Y3_FrameData_O[24] ,
    \Tile_X1Y3_FrameData_O[23] ,
    \Tile_X1Y3_FrameData_O[22] ,
    \Tile_X1Y3_FrameData_O[21] ,
    \Tile_X1Y3_FrameData_O[20] ,
    \Tile_X1Y3_FrameData_O[19] ,
    \Tile_X1Y3_FrameData_O[18] ,
    \Tile_X1Y3_FrameData_O[17] ,
    \Tile_X1Y3_FrameData_O[16] ,
    \Tile_X1Y3_FrameData_O[15] ,
    \Tile_X1Y3_FrameData_O[14] ,
    \Tile_X1Y3_FrameData_O[13] ,
    \Tile_X1Y3_FrameData_O[12] ,
    \Tile_X1Y3_FrameData_O[11] ,
    \Tile_X1Y3_FrameData_O[10] ,
    \Tile_X1Y3_FrameData_O[9] ,
    \Tile_X1Y3_FrameData_O[8] ,
    \Tile_X1Y3_FrameData_O[7] ,
    \Tile_X1Y3_FrameData_O[6] ,
    \Tile_X1Y3_FrameData_O[5] ,
    \Tile_X1Y3_FrameData_O[4] ,
    \Tile_X1Y3_FrameData_O[3] ,
    \Tile_X1Y3_FrameData_O[2] ,
    \Tile_X1Y3_FrameData_O[1] ,
    \Tile_X1Y3_FrameData_O[0] }),
    .FrameData_O({\Tile_X2Y3_FrameData_O[31] ,
    \Tile_X2Y3_FrameData_O[30] ,
    \Tile_X2Y3_FrameData_O[29] ,
    \Tile_X2Y3_FrameData_O[28] ,
    \Tile_X2Y3_FrameData_O[27] ,
    \Tile_X2Y3_FrameData_O[26] ,
    \Tile_X2Y3_FrameData_O[25] ,
    \Tile_X2Y3_FrameData_O[24] ,
    \Tile_X2Y3_FrameData_O[23] ,
    \Tile_X2Y3_FrameData_O[22] ,
    \Tile_X2Y3_FrameData_O[21] ,
    \Tile_X2Y3_FrameData_O[20] ,
    \Tile_X2Y3_FrameData_O[19] ,
    \Tile_X2Y3_FrameData_O[18] ,
    \Tile_X2Y3_FrameData_O[17] ,
    \Tile_X2Y3_FrameData_O[16] ,
    \Tile_X2Y3_FrameData_O[15] ,
    \Tile_X2Y3_FrameData_O[14] ,
    \Tile_X2Y3_FrameData_O[13] ,
    \Tile_X2Y3_FrameData_O[12] ,
    \Tile_X2Y3_FrameData_O[11] ,
    \Tile_X2Y3_FrameData_O[10] ,
    \Tile_X2Y3_FrameData_O[9] ,
    \Tile_X2Y3_FrameData_O[8] ,
    \Tile_X2Y3_FrameData_O[7] ,
    \Tile_X2Y3_FrameData_O[6] ,
    \Tile_X2Y3_FrameData_O[5] ,
    \Tile_X2Y3_FrameData_O[4] ,
    \Tile_X2Y3_FrameData_O[3] ,
    \Tile_X2Y3_FrameData_O[2] ,
    \Tile_X2Y3_FrameData_O[1] ,
    \Tile_X2Y3_FrameData_O[0] }),
    .FrameStrobe({\Tile_X2Y4_FrameStrobe_O[19] ,
    \Tile_X2Y4_FrameStrobe_O[18] ,
    \Tile_X2Y4_FrameStrobe_O[17] ,
    \Tile_X2Y4_FrameStrobe_O[16] ,
    \Tile_X2Y4_FrameStrobe_O[15] ,
    \Tile_X2Y4_FrameStrobe_O[14] ,
    \Tile_X2Y4_FrameStrobe_O[13] ,
    \Tile_X2Y4_FrameStrobe_O[12] ,
    \Tile_X2Y4_FrameStrobe_O[11] ,
    \Tile_X2Y4_FrameStrobe_O[10] ,
    \Tile_X2Y4_FrameStrobe_O[9] ,
    \Tile_X2Y4_FrameStrobe_O[8] ,
    \Tile_X2Y4_FrameStrobe_O[7] ,
    \Tile_X2Y4_FrameStrobe_O[6] ,
    \Tile_X2Y4_FrameStrobe_O[5] ,
    \Tile_X2Y4_FrameStrobe_O[4] ,
    \Tile_X2Y4_FrameStrobe_O[3] ,
    \Tile_X2Y4_FrameStrobe_O[2] ,
    \Tile_X2Y4_FrameStrobe_O[1] ,
    \Tile_X2Y4_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X2Y3_FrameStrobe_O[19] ,
    \Tile_X2Y3_FrameStrobe_O[18] ,
    \Tile_X2Y3_FrameStrobe_O[17] ,
    \Tile_X2Y3_FrameStrobe_O[16] ,
    \Tile_X2Y3_FrameStrobe_O[15] ,
    \Tile_X2Y3_FrameStrobe_O[14] ,
    \Tile_X2Y3_FrameStrobe_O[13] ,
    \Tile_X2Y3_FrameStrobe_O[12] ,
    \Tile_X2Y3_FrameStrobe_O[11] ,
    \Tile_X2Y3_FrameStrobe_O[10] ,
    \Tile_X2Y3_FrameStrobe_O[9] ,
    \Tile_X2Y3_FrameStrobe_O[8] ,
    \Tile_X2Y3_FrameStrobe_O[7] ,
    \Tile_X2Y3_FrameStrobe_O[6] ,
    \Tile_X2Y3_FrameStrobe_O[5] ,
    \Tile_X2Y3_FrameStrobe_O[4] ,
    \Tile_X2Y3_FrameStrobe_O[3] ,
    \Tile_X2Y3_FrameStrobe_O[2] ,
    \Tile_X2Y3_FrameStrobe_O[1] ,
    \Tile_X2Y3_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X2Y3_N1BEG[3] ,
    \Tile_X2Y3_N1BEG[2] ,
    \Tile_X2Y3_N1BEG[1] ,
    \Tile_X2Y3_N1BEG[0] }),
    .N1END({\Tile_X2Y4_N1BEG[3] ,
    \Tile_X2Y4_N1BEG[2] ,
    \Tile_X2Y4_N1BEG[1] ,
    \Tile_X2Y4_N1BEG[0] }),
    .N2BEG({\Tile_X2Y3_N2BEG[7] ,
    \Tile_X2Y3_N2BEG[6] ,
    \Tile_X2Y3_N2BEG[5] ,
    \Tile_X2Y3_N2BEG[4] ,
    \Tile_X2Y3_N2BEG[3] ,
    \Tile_X2Y3_N2BEG[2] ,
    \Tile_X2Y3_N2BEG[1] ,
    \Tile_X2Y3_N2BEG[0] }),
    .N2BEGb({\Tile_X2Y3_N2BEGb[7] ,
    \Tile_X2Y3_N2BEGb[6] ,
    \Tile_X2Y3_N2BEGb[5] ,
    \Tile_X2Y3_N2BEGb[4] ,
    \Tile_X2Y3_N2BEGb[3] ,
    \Tile_X2Y3_N2BEGb[2] ,
    \Tile_X2Y3_N2BEGb[1] ,
    \Tile_X2Y3_N2BEGb[0] }),
    .N2END({\Tile_X2Y4_N2BEGb[7] ,
    \Tile_X2Y4_N2BEGb[6] ,
    \Tile_X2Y4_N2BEGb[5] ,
    \Tile_X2Y4_N2BEGb[4] ,
    \Tile_X2Y4_N2BEGb[3] ,
    \Tile_X2Y4_N2BEGb[2] ,
    \Tile_X2Y4_N2BEGb[1] ,
    \Tile_X2Y4_N2BEGb[0] }),
    .N2MID({\Tile_X2Y4_N2BEG[7] ,
    \Tile_X2Y4_N2BEG[6] ,
    \Tile_X2Y4_N2BEG[5] ,
    \Tile_X2Y4_N2BEG[4] ,
    \Tile_X2Y4_N2BEG[3] ,
    \Tile_X2Y4_N2BEG[2] ,
    \Tile_X2Y4_N2BEG[1] ,
    \Tile_X2Y4_N2BEG[0] }),
    .N4BEG({\Tile_X2Y3_N4BEG[15] ,
    \Tile_X2Y3_N4BEG[14] ,
    \Tile_X2Y3_N4BEG[13] ,
    \Tile_X2Y3_N4BEG[12] ,
    \Tile_X2Y3_N4BEG[11] ,
    \Tile_X2Y3_N4BEG[10] ,
    \Tile_X2Y3_N4BEG[9] ,
    \Tile_X2Y3_N4BEG[8] ,
    \Tile_X2Y3_N4BEG[7] ,
    \Tile_X2Y3_N4BEG[6] ,
    \Tile_X2Y3_N4BEG[5] ,
    \Tile_X2Y3_N4BEG[4] ,
    \Tile_X2Y3_N4BEG[3] ,
    \Tile_X2Y3_N4BEG[2] ,
    \Tile_X2Y3_N4BEG[1] ,
    \Tile_X2Y3_N4BEG[0] }),
    .N4END({\Tile_X2Y4_N4BEG[15] ,
    \Tile_X2Y4_N4BEG[14] ,
    \Tile_X2Y4_N4BEG[13] ,
    \Tile_X2Y4_N4BEG[12] ,
    \Tile_X2Y4_N4BEG[11] ,
    \Tile_X2Y4_N4BEG[10] ,
    \Tile_X2Y4_N4BEG[9] ,
    \Tile_X2Y4_N4BEG[8] ,
    \Tile_X2Y4_N4BEG[7] ,
    \Tile_X2Y4_N4BEG[6] ,
    \Tile_X2Y4_N4BEG[5] ,
    \Tile_X2Y4_N4BEG[4] ,
    \Tile_X2Y4_N4BEG[3] ,
    \Tile_X2Y4_N4BEG[2] ,
    \Tile_X2Y4_N4BEG[1] ,
    \Tile_X2Y4_N4BEG[0] }),
    .NN4BEG({\Tile_X2Y3_NN4BEG[15] ,
    \Tile_X2Y3_NN4BEG[14] ,
    \Tile_X2Y3_NN4BEG[13] ,
    \Tile_X2Y3_NN4BEG[12] ,
    \Tile_X2Y3_NN4BEG[11] ,
    \Tile_X2Y3_NN4BEG[10] ,
    \Tile_X2Y3_NN4BEG[9] ,
    \Tile_X2Y3_NN4BEG[8] ,
    \Tile_X2Y3_NN4BEG[7] ,
    \Tile_X2Y3_NN4BEG[6] ,
    \Tile_X2Y3_NN4BEG[5] ,
    \Tile_X2Y3_NN4BEG[4] ,
    \Tile_X2Y3_NN4BEG[3] ,
    \Tile_X2Y3_NN4BEG[2] ,
    \Tile_X2Y3_NN4BEG[1] ,
    \Tile_X2Y3_NN4BEG[0] }),
    .NN4END({\Tile_X2Y4_NN4BEG[15] ,
    \Tile_X2Y4_NN4BEG[14] ,
    \Tile_X2Y4_NN4BEG[13] ,
    \Tile_X2Y4_NN4BEG[12] ,
    \Tile_X2Y4_NN4BEG[11] ,
    \Tile_X2Y4_NN4BEG[10] ,
    \Tile_X2Y4_NN4BEG[9] ,
    \Tile_X2Y4_NN4BEG[8] ,
    \Tile_X2Y4_NN4BEG[7] ,
    \Tile_X2Y4_NN4BEG[6] ,
    \Tile_X2Y4_NN4BEG[5] ,
    \Tile_X2Y4_NN4BEG[4] ,
    \Tile_X2Y4_NN4BEG[3] ,
    \Tile_X2Y4_NN4BEG[2] ,
    \Tile_X2Y4_NN4BEG[1] ,
    \Tile_X2Y4_NN4BEG[0] }),
    .S1BEG({\Tile_X2Y3_S1BEG[3] ,
    \Tile_X2Y3_S1BEG[2] ,
    \Tile_X2Y3_S1BEG[1] ,
    \Tile_X2Y3_S1BEG[0] }),
    .S1END({\Tile_X2Y2_S1BEG[3] ,
    \Tile_X2Y2_S1BEG[2] ,
    \Tile_X2Y2_S1BEG[1] ,
    \Tile_X2Y2_S1BEG[0] }),
    .S2BEG({\Tile_X2Y3_S2BEG[7] ,
    \Tile_X2Y3_S2BEG[6] ,
    \Tile_X2Y3_S2BEG[5] ,
    \Tile_X2Y3_S2BEG[4] ,
    \Tile_X2Y3_S2BEG[3] ,
    \Tile_X2Y3_S2BEG[2] ,
    \Tile_X2Y3_S2BEG[1] ,
    \Tile_X2Y3_S2BEG[0] }),
    .S2BEGb({\Tile_X2Y3_S2BEGb[7] ,
    \Tile_X2Y3_S2BEGb[6] ,
    \Tile_X2Y3_S2BEGb[5] ,
    \Tile_X2Y3_S2BEGb[4] ,
    \Tile_X2Y3_S2BEGb[3] ,
    \Tile_X2Y3_S2BEGb[2] ,
    \Tile_X2Y3_S2BEGb[1] ,
    \Tile_X2Y3_S2BEGb[0] }),
    .S2END({\Tile_X2Y2_S2BEGb[7] ,
    \Tile_X2Y2_S2BEGb[6] ,
    \Tile_X2Y2_S2BEGb[5] ,
    \Tile_X2Y2_S2BEGb[4] ,
    \Tile_X2Y2_S2BEGb[3] ,
    \Tile_X2Y2_S2BEGb[2] ,
    \Tile_X2Y2_S2BEGb[1] ,
    \Tile_X2Y2_S2BEGb[0] }),
    .S2MID({\Tile_X2Y2_S2BEG[7] ,
    \Tile_X2Y2_S2BEG[6] ,
    \Tile_X2Y2_S2BEG[5] ,
    \Tile_X2Y2_S2BEG[4] ,
    \Tile_X2Y2_S2BEG[3] ,
    \Tile_X2Y2_S2BEG[2] ,
    \Tile_X2Y2_S2BEG[1] ,
    \Tile_X2Y2_S2BEG[0] }),
    .S4BEG({\Tile_X2Y3_S4BEG[15] ,
    \Tile_X2Y3_S4BEG[14] ,
    \Tile_X2Y3_S4BEG[13] ,
    \Tile_X2Y3_S4BEG[12] ,
    \Tile_X2Y3_S4BEG[11] ,
    \Tile_X2Y3_S4BEG[10] ,
    \Tile_X2Y3_S4BEG[9] ,
    \Tile_X2Y3_S4BEG[8] ,
    \Tile_X2Y3_S4BEG[7] ,
    \Tile_X2Y3_S4BEG[6] ,
    \Tile_X2Y3_S4BEG[5] ,
    \Tile_X2Y3_S4BEG[4] ,
    \Tile_X2Y3_S4BEG[3] ,
    \Tile_X2Y3_S4BEG[2] ,
    \Tile_X2Y3_S4BEG[1] ,
    \Tile_X2Y3_S4BEG[0] }),
    .S4END({\Tile_X2Y2_S4BEG[15] ,
    \Tile_X2Y2_S4BEG[14] ,
    \Tile_X2Y2_S4BEG[13] ,
    \Tile_X2Y2_S4BEG[12] ,
    \Tile_X2Y2_S4BEG[11] ,
    \Tile_X2Y2_S4BEG[10] ,
    \Tile_X2Y2_S4BEG[9] ,
    \Tile_X2Y2_S4BEG[8] ,
    \Tile_X2Y2_S4BEG[7] ,
    \Tile_X2Y2_S4BEG[6] ,
    \Tile_X2Y2_S4BEG[5] ,
    \Tile_X2Y2_S4BEG[4] ,
    \Tile_X2Y2_S4BEG[3] ,
    \Tile_X2Y2_S4BEG[2] ,
    \Tile_X2Y2_S4BEG[1] ,
    \Tile_X2Y2_S4BEG[0] }),
    .SS4BEG({\Tile_X2Y3_SS4BEG[15] ,
    \Tile_X2Y3_SS4BEG[14] ,
    \Tile_X2Y3_SS4BEG[13] ,
    \Tile_X2Y3_SS4BEG[12] ,
    \Tile_X2Y3_SS4BEG[11] ,
    \Tile_X2Y3_SS4BEG[10] ,
    \Tile_X2Y3_SS4BEG[9] ,
    \Tile_X2Y3_SS4BEG[8] ,
    \Tile_X2Y3_SS4BEG[7] ,
    \Tile_X2Y3_SS4BEG[6] ,
    \Tile_X2Y3_SS4BEG[5] ,
    \Tile_X2Y3_SS4BEG[4] ,
    \Tile_X2Y3_SS4BEG[3] ,
    \Tile_X2Y3_SS4BEG[2] ,
    \Tile_X2Y3_SS4BEG[1] ,
    \Tile_X2Y3_SS4BEG[0] }),
    .SS4END({\Tile_X2Y2_SS4BEG[15] ,
    \Tile_X2Y2_SS4BEG[14] ,
    \Tile_X2Y2_SS4BEG[13] ,
    \Tile_X2Y2_SS4BEG[12] ,
    \Tile_X2Y2_SS4BEG[11] ,
    \Tile_X2Y2_SS4BEG[10] ,
    \Tile_X2Y2_SS4BEG[9] ,
    \Tile_X2Y2_SS4BEG[8] ,
    \Tile_X2Y2_SS4BEG[7] ,
    \Tile_X2Y2_SS4BEG[6] ,
    \Tile_X2Y2_SS4BEG[5] ,
    \Tile_X2Y2_SS4BEG[4] ,
    \Tile_X2Y2_SS4BEG[3] ,
    \Tile_X2Y2_SS4BEG[2] ,
    \Tile_X2Y2_SS4BEG[1] ,
    \Tile_X2Y2_SS4BEG[0] }),
    .W1BEG({\Tile_X2Y3_W1BEG[3] ,
    \Tile_X2Y3_W1BEG[2] ,
    \Tile_X2Y3_W1BEG[1] ,
    \Tile_X2Y3_W1BEG[0] }),
    .W1END({\Tile_X3Y3_W1BEG[3] ,
    \Tile_X3Y3_W1BEG[2] ,
    \Tile_X3Y3_W1BEG[1] ,
    \Tile_X3Y3_W1BEG[0] }),
    .W2BEG({\Tile_X2Y3_W2BEG[7] ,
    \Tile_X2Y3_W2BEG[6] ,
    \Tile_X2Y3_W2BEG[5] ,
    \Tile_X2Y3_W2BEG[4] ,
    \Tile_X2Y3_W2BEG[3] ,
    \Tile_X2Y3_W2BEG[2] ,
    \Tile_X2Y3_W2BEG[1] ,
    \Tile_X2Y3_W2BEG[0] }),
    .W2BEGb({\Tile_X2Y3_W2BEGb[7] ,
    \Tile_X2Y3_W2BEGb[6] ,
    \Tile_X2Y3_W2BEGb[5] ,
    \Tile_X2Y3_W2BEGb[4] ,
    \Tile_X2Y3_W2BEGb[3] ,
    \Tile_X2Y3_W2BEGb[2] ,
    \Tile_X2Y3_W2BEGb[1] ,
    \Tile_X2Y3_W2BEGb[0] }),
    .W2END({\Tile_X3Y3_W2BEGb[7] ,
    \Tile_X3Y3_W2BEGb[6] ,
    \Tile_X3Y3_W2BEGb[5] ,
    \Tile_X3Y3_W2BEGb[4] ,
    \Tile_X3Y3_W2BEGb[3] ,
    \Tile_X3Y3_W2BEGb[2] ,
    \Tile_X3Y3_W2BEGb[1] ,
    \Tile_X3Y3_W2BEGb[0] }),
    .W2MID({\Tile_X3Y3_W2BEG[7] ,
    \Tile_X3Y3_W2BEG[6] ,
    \Tile_X3Y3_W2BEG[5] ,
    \Tile_X3Y3_W2BEG[4] ,
    \Tile_X3Y3_W2BEG[3] ,
    \Tile_X3Y3_W2BEG[2] ,
    \Tile_X3Y3_W2BEG[1] ,
    \Tile_X3Y3_W2BEG[0] }),
    .W6BEG({\Tile_X2Y3_W6BEG[11] ,
    \Tile_X2Y3_W6BEG[10] ,
    \Tile_X2Y3_W6BEG[9] ,
    \Tile_X2Y3_W6BEG[8] ,
    \Tile_X2Y3_W6BEG[7] ,
    \Tile_X2Y3_W6BEG[6] ,
    \Tile_X2Y3_W6BEG[5] ,
    \Tile_X2Y3_W6BEG[4] ,
    \Tile_X2Y3_W6BEG[3] ,
    \Tile_X2Y3_W6BEG[2] ,
    \Tile_X2Y3_W6BEG[1] ,
    \Tile_X2Y3_W6BEG[0] }),
    .W6END({\Tile_X3Y3_W6BEG[11] ,
    \Tile_X3Y3_W6BEG[10] ,
    \Tile_X3Y3_W6BEG[9] ,
    \Tile_X3Y3_W6BEG[8] ,
    \Tile_X3Y3_W6BEG[7] ,
    \Tile_X3Y3_W6BEG[6] ,
    \Tile_X3Y3_W6BEG[5] ,
    \Tile_X3Y3_W6BEG[4] ,
    \Tile_X3Y3_W6BEG[3] ,
    \Tile_X3Y3_W6BEG[2] ,
    \Tile_X3Y3_W6BEG[1] ,
    \Tile_X3Y3_W6BEG[0] }),
    .WW4BEG({\Tile_X2Y3_WW4BEG[15] ,
    \Tile_X2Y3_WW4BEG[14] ,
    \Tile_X2Y3_WW4BEG[13] ,
    \Tile_X2Y3_WW4BEG[12] ,
    \Tile_X2Y3_WW4BEG[11] ,
    \Tile_X2Y3_WW4BEG[10] ,
    \Tile_X2Y3_WW4BEG[9] ,
    \Tile_X2Y3_WW4BEG[8] ,
    \Tile_X2Y3_WW4BEG[7] ,
    \Tile_X2Y3_WW4BEG[6] ,
    \Tile_X2Y3_WW4BEG[5] ,
    \Tile_X2Y3_WW4BEG[4] ,
    \Tile_X2Y3_WW4BEG[3] ,
    \Tile_X2Y3_WW4BEG[2] ,
    \Tile_X2Y3_WW4BEG[1] ,
    \Tile_X2Y3_WW4BEG[0] }),
    .WW4END({\Tile_X3Y3_WW4BEG[15] ,
    \Tile_X3Y3_WW4BEG[14] ,
    \Tile_X3Y3_WW4BEG[13] ,
    \Tile_X3Y3_WW4BEG[12] ,
    \Tile_X3Y3_WW4BEG[11] ,
    \Tile_X3Y3_WW4BEG[10] ,
    \Tile_X3Y3_WW4BEG[9] ,
    \Tile_X3Y3_WW4BEG[8] ,
    \Tile_X3Y3_WW4BEG[7] ,
    \Tile_X3Y3_WW4BEG[6] ,
    \Tile_X3Y3_WW4BEG[5] ,
    \Tile_X3Y3_WW4BEG[4] ,
    \Tile_X3Y3_WW4BEG[3] ,
    \Tile_X3Y3_WW4BEG[2] ,
    \Tile_X3Y3_WW4BEG[1] ,
    \Tile_X3Y3_WW4BEG[0] }));
 LUT4AB Tile_X2Y4_LUT4AB (.Ci(Tile_X2Y5_Co),
    .Co(Tile_X2Y4_Co),
    .UserCLK(Tile_X2Y5_UserCLKo),
    .UserCLKo(Tile_X2Y4_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X2Y4_E1BEG[3] ,
    \Tile_X2Y4_E1BEG[2] ,
    \Tile_X2Y4_E1BEG[1] ,
    \Tile_X2Y4_E1BEG[0] }),
    .E1END({\Tile_X1Y4_E1BEG[3] ,
    \Tile_X1Y4_E1BEG[2] ,
    \Tile_X1Y4_E1BEG[1] ,
    \Tile_X1Y4_E1BEG[0] }),
    .E2BEG({\Tile_X2Y4_E2BEG[7] ,
    \Tile_X2Y4_E2BEG[6] ,
    \Tile_X2Y4_E2BEG[5] ,
    \Tile_X2Y4_E2BEG[4] ,
    \Tile_X2Y4_E2BEG[3] ,
    \Tile_X2Y4_E2BEG[2] ,
    \Tile_X2Y4_E2BEG[1] ,
    \Tile_X2Y4_E2BEG[0] }),
    .E2BEGb({\Tile_X2Y4_E2BEGb[7] ,
    \Tile_X2Y4_E2BEGb[6] ,
    \Tile_X2Y4_E2BEGb[5] ,
    \Tile_X2Y4_E2BEGb[4] ,
    \Tile_X2Y4_E2BEGb[3] ,
    \Tile_X2Y4_E2BEGb[2] ,
    \Tile_X2Y4_E2BEGb[1] ,
    \Tile_X2Y4_E2BEGb[0] }),
    .E2END({\Tile_X1Y4_E2BEGb[7] ,
    \Tile_X1Y4_E2BEGb[6] ,
    \Tile_X1Y4_E2BEGb[5] ,
    \Tile_X1Y4_E2BEGb[4] ,
    \Tile_X1Y4_E2BEGb[3] ,
    \Tile_X1Y4_E2BEGb[2] ,
    \Tile_X1Y4_E2BEGb[1] ,
    \Tile_X1Y4_E2BEGb[0] }),
    .E2MID({\Tile_X1Y4_E2BEG[7] ,
    \Tile_X1Y4_E2BEG[6] ,
    \Tile_X1Y4_E2BEG[5] ,
    \Tile_X1Y4_E2BEG[4] ,
    \Tile_X1Y4_E2BEG[3] ,
    \Tile_X1Y4_E2BEG[2] ,
    \Tile_X1Y4_E2BEG[1] ,
    \Tile_X1Y4_E2BEG[0] }),
    .E6BEG({\Tile_X2Y4_E6BEG[11] ,
    \Tile_X2Y4_E6BEG[10] ,
    \Tile_X2Y4_E6BEG[9] ,
    \Tile_X2Y4_E6BEG[8] ,
    \Tile_X2Y4_E6BEG[7] ,
    \Tile_X2Y4_E6BEG[6] ,
    \Tile_X2Y4_E6BEG[5] ,
    \Tile_X2Y4_E6BEG[4] ,
    \Tile_X2Y4_E6BEG[3] ,
    \Tile_X2Y4_E6BEG[2] ,
    \Tile_X2Y4_E6BEG[1] ,
    \Tile_X2Y4_E6BEG[0] }),
    .E6END({\Tile_X1Y4_E6BEG[11] ,
    \Tile_X1Y4_E6BEG[10] ,
    \Tile_X1Y4_E6BEG[9] ,
    \Tile_X1Y4_E6BEG[8] ,
    \Tile_X1Y4_E6BEG[7] ,
    \Tile_X1Y4_E6BEG[6] ,
    \Tile_X1Y4_E6BEG[5] ,
    \Tile_X1Y4_E6BEG[4] ,
    \Tile_X1Y4_E6BEG[3] ,
    \Tile_X1Y4_E6BEG[2] ,
    \Tile_X1Y4_E6BEG[1] ,
    \Tile_X1Y4_E6BEG[0] }),
    .EE4BEG({\Tile_X2Y4_EE4BEG[15] ,
    \Tile_X2Y4_EE4BEG[14] ,
    \Tile_X2Y4_EE4BEG[13] ,
    \Tile_X2Y4_EE4BEG[12] ,
    \Tile_X2Y4_EE4BEG[11] ,
    \Tile_X2Y4_EE4BEG[10] ,
    \Tile_X2Y4_EE4BEG[9] ,
    \Tile_X2Y4_EE4BEG[8] ,
    \Tile_X2Y4_EE4BEG[7] ,
    \Tile_X2Y4_EE4BEG[6] ,
    \Tile_X2Y4_EE4BEG[5] ,
    \Tile_X2Y4_EE4BEG[4] ,
    \Tile_X2Y4_EE4BEG[3] ,
    \Tile_X2Y4_EE4BEG[2] ,
    \Tile_X2Y4_EE4BEG[1] ,
    \Tile_X2Y4_EE4BEG[0] }),
    .EE4END({\Tile_X1Y4_EE4BEG[15] ,
    \Tile_X1Y4_EE4BEG[14] ,
    \Tile_X1Y4_EE4BEG[13] ,
    \Tile_X1Y4_EE4BEG[12] ,
    \Tile_X1Y4_EE4BEG[11] ,
    \Tile_X1Y4_EE4BEG[10] ,
    \Tile_X1Y4_EE4BEG[9] ,
    \Tile_X1Y4_EE4BEG[8] ,
    \Tile_X1Y4_EE4BEG[7] ,
    \Tile_X1Y4_EE4BEG[6] ,
    \Tile_X1Y4_EE4BEG[5] ,
    \Tile_X1Y4_EE4BEG[4] ,
    \Tile_X1Y4_EE4BEG[3] ,
    \Tile_X1Y4_EE4BEG[2] ,
    \Tile_X1Y4_EE4BEG[1] ,
    \Tile_X1Y4_EE4BEG[0] }),
    .FrameData({\Tile_X1Y4_FrameData_O[31] ,
    \Tile_X1Y4_FrameData_O[30] ,
    \Tile_X1Y4_FrameData_O[29] ,
    \Tile_X1Y4_FrameData_O[28] ,
    \Tile_X1Y4_FrameData_O[27] ,
    \Tile_X1Y4_FrameData_O[26] ,
    \Tile_X1Y4_FrameData_O[25] ,
    \Tile_X1Y4_FrameData_O[24] ,
    \Tile_X1Y4_FrameData_O[23] ,
    \Tile_X1Y4_FrameData_O[22] ,
    \Tile_X1Y4_FrameData_O[21] ,
    \Tile_X1Y4_FrameData_O[20] ,
    \Tile_X1Y4_FrameData_O[19] ,
    \Tile_X1Y4_FrameData_O[18] ,
    \Tile_X1Y4_FrameData_O[17] ,
    \Tile_X1Y4_FrameData_O[16] ,
    \Tile_X1Y4_FrameData_O[15] ,
    \Tile_X1Y4_FrameData_O[14] ,
    \Tile_X1Y4_FrameData_O[13] ,
    \Tile_X1Y4_FrameData_O[12] ,
    \Tile_X1Y4_FrameData_O[11] ,
    \Tile_X1Y4_FrameData_O[10] ,
    \Tile_X1Y4_FrameData_O[9] ,
    \Tile_X1Y4_FrameData_O[8] ,
    \Tile_X1Y4_FrameData_O[7] ,
    \Tile_X1Y4_FrameData_O[6] ,
    \Tile_X1Y4_FrameData_O[5] ,
    \Tile_X1Y4_FrameData_O[4] ,
    \Tile_X1Y4_FrameData_O[3] ,
    \Tile_X1Y4_FrameData_O[2] ,
    \Tile_X1Y4_FrameData_O[1] ,
    \Tile_X1Y4_FrameData_O[0] }),
    .FrameData_O({\Tile_X2Y4_FrameData_O[31] ,
    \Tile_X2Y4_FrameData_O[30] ,
    \Tile_X2Y4_FrameData_O[29] ,
    \Tile_X2Y4_FrameData_O[28] ,
    \Tile_X2Y4_FrameData_O[27] ,
    \Tile_X2Y4_FrameData_O[26] ,
    \Tile_X2Y4_FrameData_O[25] ,
    \Tile_X2Y4_FrameData_O[24] ,
    \Tile_X2Y4_FrameData_O[23] ,
    \Tile_X2Y4_FrameData_O[22] ,
    \Tile_X2Y4_FrameData_O[21] ,
    \Tile_X2Y4_FrameData_O[20] ,
    \Tile_X2Y4_FrameData_O[19] ,
    \Tile_X2Y4_FrameData_O[18] ,
    \Tile_X2Y4_FrameData_O[17] ,
    \Tile_X2Y4_FrameData_O[16] ,
    \Tile_X2Y4_FrameData_O[15] ,
    \Tile_X2Y4_FrameData_O[14] ,
    \Tile_X2Y4_FrameData_O[13] ,
    \Tile_X2Y4_FrameData_O[12] ,
    \Tile_X2Y4_FrameData_O[11] ,
    \Tile_X2Y4_FrameData_O[10] ,
    \Tile_X2Y4_FrameData_O[9] ,
    \Tile_X2Y4_FrameData_O[8] ,
    \Tile_X2Y4_FrameData_O[7] ,
    \Tile_X2Y4_FrameData_O[6] ,
    \Tile_X2Y4_FrameData_O[5] ,
    \Tile_X2Y4_FrameData_O[4] ,
    \Tile_X2Y4_FrameData_O[3] ,
    \Tile_X2Y4_FrameData_O[2] ,
    \Tile_X2Y4_FrameData_O[1] ,
    \Tile_X2Y4_FrameData_O[0] }),
    .FrameStrobe({\Tile_X2Y5_FrameStrobe_O[19] ,
    \Tile_X2Y5_FrameStrobe_O[18] ,
    \Tile_X2Y5_FrameStrobe_O[17] ,
    \Tile_X2Y5_FrameStrobe_O[16] ,
    \Tile_X2Y5_FrameStrobe_O[15] ,
    \Tile_X2Y5_FrameStrobe_O[14] ,
    \Tile_X2Y5_FrameStrobe_O[13] ,
    \Tile_X2Y5_FrameStrobe_O[12] ,
    \Tile_X2Y5_FrameStrobe_O[11] ,
    \Tile_X2Y5_FrameStrobe_O[10] ,
    \Tile_X2Y5_FrameStrobe_O[9] ,
    \Tile_X2Y5_FrameStrobe_O[8] ,
    \Tile_X2Y5_FrameStrobe_O[7] ,
    \Tile_X2Y5_FrameStrobe_O[6] ,
    \Tile_X2Y5_FrameStrobe_O[5] ,
    \Tile_X2Y5_FrameStrobe_O[4] ,
    \Tile_X2Y5_FrameStrobe_O[3] ,
    \Tile_X2Y5_FrameStrobe_O[2] ,
    \Tile_X2Y5_FrameStrobe_O[1] ,
    \Tile_X2Y5_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X2Y4_FrameStrobe_O[19] ,
    \Tile_X2Y4_FrameStrobe_O[18] ,
    \Tile_X2Y4_FrameStrobe_O[17] ,
    \Tile_X2Y4_FrameStrobe_O[16] ,
    \Tile_X2Y4_FrameStrobe_O[15] ,
    \Tile_X2Y4_FrameStrobe_O[14] ,
    \Tile_X2Y4_FrameStrobe_O[13] ,
    \Tile_X2Y4_FrameStrobe_O[12] ,
    \Tile_X2Y4_FrameStrobe_O[11] ,
    \Tile_X2Y4_FrameStrobe_O[10] ,
    \Tile_X2Y4_FrameStrobe_O[9] ,
    \Tile_X2Y4_FrameStrobe_O[8] ,
    \Tile_X2Y4_FrameStrobe_O[7] ,
    \Tile_X2Y4_FrameStrobe_O[6] ,
    \Tile_X2Y4_FrameStrobe_O[5] ,
    \Tile_X2Y4_FrameStrobe_O[4] ,
    \Tile_X2Y4_FrameStrobe_O[3] ,
    \Tile_X2Y4_FrameStrobe_O[2] ,
    \Tile_X2Y4_FrameStrobe_O[1] ,
    \Tile_X2Y4_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X2Y4_N1BEG[3] ,
    \Tile_X2Y4_N1BEG[2] ,
    \Tile_X2Y4_N1BEG[1] ,
    \Tile_X2Y4_N1BEG[0] }),
    .N1END({\Tile_X2Y5_N1BEG[3] ,
    \Tile_X2Y5_N1BEG[2] ,
    \Tile_X2Y5_N1BEG[1] ,
    \Tile_X2Y5_N1BEG[0] }),
    .N2BEG({\Tile_X2Y4_N2BEG[7] ,
    \Tile_X2Y4_N2BEG[6] ,
    \Tile_X2Y4_N2BEG[5] ,
    \Tile_X2Y4_N2BEG[4] ,
    \Tile_X2Y4_N2BEG[3] ,
    \Tile_X2Y4_N2BEG[2] ,
    \Tile_X2Y4_N2BEG[1] ,
    \Tile_X2Y4_N2BEG[0] }),
    .N2BEGb({\Tile_X2Y4_N2BEGb[7] ,
    \Tile_X2Y4_N2BEGb[6] ,
    \Tile_X2Y4_N2BEGb[5] ,
    \Tile_X2Y4_N2BEGb[4] ,
    \Tile_X2Y4_N2BEGb[3] ,
    \Tile_X2Y4_N2BEGb[2] ,
    \Tile_X2Y4_N2BEGb[1] ,
    \Tile_X2Y4_N2BEGb[0] }),
    .N2END({\Tile_X2Y5_N2BEGb[7] ,
    \Tile_X2Y5_N2BEGb[6] ,
    \Tile_X2Y5_N2BEGb[5] ,
    \Tile_X2Y5_N2BEGb[4] ,
    \Tile_X2Y5_N2BEGb[3] ,
    \Tile_X2Y5_N2BEGb[2] ,
    \Tile_X2Y5_N2BEGb[1] ,
    \Tile_X2Y5_N2BEGb[0] }),
    .N2MID({\Tile_X2Y5_N2BEG[7] ,
    \Tile_X2Y5_N2BEG[6] ,
    \Tile_X2Y5_N2BEG[5] ,
    \Tile_X2Y5_N2BEG[4] ,
    \Tile_X2Y5_N2BEG[3] ,
    \Tile_X2Y5_N2BEG[2] ,
    \Tile_X2Y5_N2BEG[1] ,
    \Tile_X2Y5_N2BEG[0] }),
    .N4BEG({\Tile_X2Y4_N4BEG[15] ,
    \Tile_X2Y4_N4BEG[14] ,
    \Tile_X2Y4_N4BEG[13] ,
    \Tile_X2Y4_N4BEG[12] ,
    \Tile_X2Y4_N4BEG[11] ,
    \Tile_X2Y4_N4BEG[10] ,
    \Tile_X2Y4_N4BEG[9] ,
    \Tile_X2Y4_N4BEG[8] ,
    \Tile_X2Y4_N4BEG[7] ,
    \Tile_X2Y4_N4BEG[6] ,
    \Tile_X2Y4_N4BEG[5] ,
    \Tile_X2Y4_N4BEG[4] ,
    \Tile_X2Y4_N4BEG[3] ,
    \Tile_X2Y4_N4BEG[2] ,
    \Tile_X2Y4_N4BEG[1] ,
    \Tile_X2Y4_N4BEG[0] }),
    .N4END({\Tile_X2Y5_N4BEG[15] ,
    \Tile_X2Y5_N4BEG[14] ,
    \Tile_X2Y5_N4BEG[13] ,
    \Tile_X2Y5_N4BEG[12] ,
    \Tile_X2Y5_N4BEG[11] ,
    \Tile_X2Y5_N4BEG[10] ,
    \Tile_X2Y5_N4BEG[9] ,
    \Tile_X2Y5_N4BEG[8] ,
    \Tile_X2Y5_N4BEG[7] ,
    \Tile_X2Y5_N4BEG[6] ,
    \Tile_X2Y5_N4BEG[5] ,
    \Tile_X2Y5_N4BEG[4] ,
    \Tile_X2Y5_N4BEG[3] ,
    \Tile_X2Y5_N4BEG[2] ,
    \Tile_X2Y5_N4BEG[1] ,
    \Tile_X2Y5_N4BEG[0] }),
    .NN4BEG({\Tile_X2Y4_NN4BEG[15] ,
    \Tile_X2Y4_NN4BEG[14] ,
    \Tile_X2Y4_NN4BEG[13] ,
    \Tile_X2Y4_NN4BEG[12] ,
    \Tile_X2Y4_NN4BEG[11] ,
    \Tile_X2Y4_NN4BEG[10] ,
    \Tile_X2Y4_NN4BEG[9] ,
    \Tile_X2Y4_NN4BEG[8] ,
    \Tile_X2Y4_NN4BEG[7] ,
    \Tile_X2Y4_NN4BEG[6] ,
    \Tile_X2Y4_NN4BEG[5] ,
    \Tile_X2Y4_NN4BEG[4] ,
    \Tile_X2Y4_NN4BEG[3] ,
    \Tile_X2Y4_NN4BEG[2] ,
    \Tile_X2Y4_NN4BEG[1] ,
    \Tile_X2Y4_NN4BEG[0] }),
    .NN4END({\Tile_X2Y5_NN4BEG[15] ,
    \Tile_X2Y5_NN4BEG[14] ,
    \Tile_X2Y5_NN4BEG[13] ,
    \Tile_X2Y5_NN4BEG[12] ,
    \Tile_X2Y5_NN4BEG[11] ,
    \Tile_X2Y5_NN4BEG[10] ,
    \Tile_X2Y5_NN4BEG[9] ,
    \Tile_X2Y5_NN4BEG[8] ,
    \Tile_X2Y5_NN4BEG[7] ,
    \Tile_X2Y5_NN4BEG[6] ,
    \Tile_X2Y5_NN4BEG[5] ,
    \Tile_X2Y5_NN4BEG[4] ,
    \Tile_X2Y5_NN4BEG[3] ,
    \Tile_X2Y5_NN4BEG[2] ,
    \Tile_X2Y5_NN4BEG[1] ,
    \Tile_X2Y5_NN4BEG[0] }),
    .S1BEG({\Tile_X2Y4_S1BEG[3] ,
    \Tile_X2Y4_S1BEG[2] ,
    \Tile_X2Y4_S1BEG[1] ,
    \Tile_X2Y4_S1BEG[0] }),
    .S1END({\Tile_X2Y3_S1BEG[3] ,
    \Tile_X2Y3_S1BEG[2] ,
    \Tile_X2Y3_S1BEG[1] ,
    \Tile_X2Y3_S1BEG[0] }),
    .S2BEG({\Tile_X2Y4_S2BEG[7] ,
    \Tile_X2Y4_S2BEG[6] ,
    \Tile_X2Y4_S2BEG[5] ,
    \Tile_X2Y4_S2BEG[4] ,
    \Tile_X2Y4_S2BEG[3] ,
    \Tile_X2Y4_S2BEG[2] ,
    \Tile_X2Y4_S2BEG[1] ,
    \Tile_X2Y4_S2BEG[0] }),
    .S2BEGb({\Tile_X2Y4_S2BEGb[7] ,
    \Tile_X2Y4_S2BEGb[6] ,
    \Tile_X2Y4_S2BEGb[5] ,
    \Tile_X2Y4_S2BEGb[4] ,
    \Tile_X2Y4_S2BEGb[3] ,
    \Tile_X2Y4_S2BEGb[2] ,
    \Tile_X2Y4_S2BEGb[1] ,
    \Tile_X2Y4_S2BEGb[0] }),
    .S2END({\Tile_X2Y3_S2BEGb[7] ,
    \Tile_X2Y3_S2BEGb[6] ,
    \Tile_X2Y3_S2BEGb[5] ,
    \Tile_X2Y3_S2BEGb[4] ,
    \Tile_X2Y3_S2BEGb[3] ,
    \Tile_X2Y3_S2BEGb[2] ,
    \Tile_X2Y3_S2BEGb[1] ,
    \Tile_X2Y3_S2BEGb[0] }),
    .S2MID({\Tile_X2Y3_S2BEG[7] ,
    \Tile_X2Y3_S2BEG[6] ,
    \Tile_X2Y3_S2BEG[5] ,
    \Tile_X2Y3_S2BEG[4] ,
    \Tile_X2Y3_S2BEG[3] ,
    \Tile_X2Y3_S2BEG[2] ,
    \Tile_X2Y3_S2BEG[1] ,
    \Tile_X2Y3_S2BEG[0] }),
    .S4BEG({\Tile_X2Y4_S4BEG[15] ,
    \Tile_X2Y4_S4BEG[14] ,
    \Tile_X2Y4_S4BEG[13] ,
    \Tile_X2Y4_S4BEG[12] ,
    \Tile_X2Y4_S4BEG[11] ,
    \Tile_X2Y4_S4BEG[10] ,
    \Tile_X2Y4_S4BEG[9] ,
    \Tile_X2Y4_S4BEG[8] ,
    \Tile_X2Y4_S4BEG[7] ,
    \Tile_X2Y4_S4BEG[6] ,
    \Tile_X2Y4_S4BEG[5] ,
    \Tile_X2Y4_S4BEG[4] ,
    \Tile_X2Y4_S4BEG[3] ,
    \Tile_X2Y4_S4BEG[2] ,
    \Tile_X2Y4_S4BEG[1] ,
    \Tile_X2Y4_S4BEG[0] }),
    .S4END({\Tile_X2Y3_S4BEG[15] ,
    \Tile_X2Y3_S4BEG[14] ,
    \Tile_X2Y3_S4BEG[13] ,
    \Tile_X2Y3_S4BEG[12] ,
    \Tile_X2Y3_S4BEG[11] ,
    \Tile_X2Y3_S4BEG[10] ,
    \Tile_X2Y3_S4BEG[9] ,
    \Tile_X2Y3_S4BEG[8] ,
    \Tile_X2Y3_S4BEG[7] ,
    \Tile_X2Y3_S4BEG[6] ,
    \Tile_X2Y3_S4BEG[5] ,
    \Tile_X2Y3_S4BEG[4] ,
    \Tile_X2Y3_S4BEG[3] ,
    \Tile_X2Y3_S4BEG[2] ,
    \Tile_X2Y3_S4BEG[1] ,
    \Tile_X2Y3_S4BEG[0] }),
    .SS4BEG({\Tile_X2Y4_SS4BEG[15] ,
    \Tile_X2Y4_SS4BEG[14] ,
    \Tile_X2Y4_SS4BEG[13] ,
    \Tile_X2Y4_SS4BEG[12] ,
    \Tile_X2Y4_SS4BEG[11] ,
    \Tile_X2Y4_SS4BEG[10] ,
    \Tile_X2Y4_SS4BEG[9] ,
    \Tile_X2Y4_SS4BEG[8] ,
    \Tile_X2Y4_SS4BEG[7] ,
    \Tile_X2Y4_SS4BEG[6] ,
    \Tile_X2Y4_SS4BEG[5] ,
    \Tile_X2Y4_SS4BEG[4] ,
    \Tile_X2Y4_SS4BEG[3] ,
    \Tile_X2Y4_SS4BEG[2] ,
    \Tile_X2Y4_SS4BEG[1] ,
    \Tile_X2Y4_SS4BEG[0] }),
    .SS4END({\Tile_X2Y3_SS4BEG[15] ,
    \Tile_X2Y3_SS4BEG[14] ,
    \Tile_X2Y3_SS4BEG[13] ,
    \Tile_X2Y3_SS4BEG[12] ,
    \Tile_X2Y3_SS4BEG[11] ,
    \Tile_X2Y3_SS4BEG[10] ,
    \Tile_X2Y3_SS4BEG[9] ,
    \Tile_X2Y3_SS4BEG[8] ,
    \Tile_X2Y3_SS4BEG[7] ,
    \Tile_X2Y3_SS4BEG[6] ,
    \Tile_X2Y3_SS4BEG[5] ,
    \Tile_X2Y3_SS4BEG[4] ,
    \Tile_X2Y3_SS4BEG[3] ,
    \Tile_X2Y3_SS4BEG[2] ,
    \Tile_X2Y3_SS4BEG[1] ,
    \Tile_X2Y3_SS4BEG[0] }),
    .W1BEG({\Tile_X2Y4_W1BEG[3] ,
    \Tile_X2Y4_W1BEG[2] ,
    \Tile_X2Y4_W1BEG[1] ,
    \Tile_X2Y4_W1BEG[0] }),
    .W1END({\Tile_X3Y4_W1BEG[3] ,
    \Tile_X3Y4_W1BEG[2] ,
    \Tile_X3Y4_W1BEG[1] ,
    \Tile_X3Y4_W1BEG[0] }),
    .W2BEG({\Tile_X2Y4_W2BEG[7] ,
    \Tile_X2Y4_W2BEG[6] ,
    \Tile_X2Y4_W2BEG[5] ,
    \Tile_X2Y4_W2BEG[4] ,
    \Tile_X2Y4_W2BEG[3] ,
    \Tile_X2Y4_W2BEG[2] ,
    \Tile_X2Y4_W2BEG[1] ,
    \Tile_X2Y4_W2BEG[0] }),
    .W2BEGb({\Tile_X2Y4_W2BEGb[7] ,
    \Tile_X2Y4_W2BEGb[6] ,
    \Tile_X2Y4_W2BEGb[5] ,
    \Tile_X2Y4_W2BEGb[4] ,
    \Tile_X2Y4_W2BEGb[3] ,
    \Tile_X2Y4_W2BEGb[2] ,
    \Tile_X2Y4_W2BEGb[1] ,
    \Tile_X2Y4_W2BEGb[0] }),
    .W2END({\Tile_X3Y4_W2BEGb[7] ,
    \Tile_X3Y4_W2BEGb[6] ,
    \Tile_X3Y4_W2BEGb[5] ,
    \Tile_X3Y4_W2BEGb[4] ,
    \Tile_X3Y4_W2BEGb[3] ,
    \Tile_X3Y4_W2BEGb[2] ,
    \Tile_X3Y4_W2BEGb[1] ,
    \Tile_X3Y4_W2BEGb[0] }),
    .W2MID({\Tile_X3Y4_W2BEG[7] ,
    \Tile_X3Y4_W2BEG[6] ,
    \Tile_X3Y4_W2BEG[5] ,
    \Tile_X3Y4_W2BEG[4] ,
    \Tile_X3Y4_W2BEG[3] ,
    \Tile_X3Y4_W2BEG[2] ,
    \Tile_X3Y4_W2BEG[1] ,
    \Tile_X3Y4_W2BEG[0] }),
    .W6BEG({\Tile_X2Y4_W6BEG[11] ,
    \Tile_X2Y4_W6BEG[10] ,
    \Tile_X2Y4_W6BEG[9] ,
    \Tile_X2Y4_W6BEG[8] ,
    \Tile_X2Y4_W6BEG[7] ,
    \Tile_X2Y4_W6BEG[6] ,
    \Tile_X2Y4_W6BEG[5] ,
    \Tile_X2Y4_W6BEG[4] ,
    \Tile_X2Y4_W6BEG[3] ,
    \Tile_X2Y4_W6BEG[2] ,
    \Tile_X2Y4_W6BEG[1] ,
    \Tile_X2Y4_W6BEG[0] }),
    .W6END({\Tile_X3Y4_W6BEG[11] ,
    \Tile_X3Y4_W6BEG[10] ,
    \Tile_X3Y4_W6BEG[9] ,
    \Tile_X3Y4_W6BEG[8] ,
    \Tile_X3Y4_W6BEG[7] ,
    \Tile_X3Y4_W6BEG[6] ,
    \Tile_X3Y4_W6BEG[5] ,
    \Tile_X3Y4_W6BEG[4] ,
    \Tile_X3Y4_W6BEG[3] ,
    \Tile_X3Y4_W6BEG[2] ,
    \Tile_X3Y4_W6BEG[1] ,
    \Tile_X3Y4_W6BEG[0] }),
    .WW4BEG({\Tile_X2Y4_WW4BEG[15] ,
    \Tile_X2Y4_WW4BEG[14] ,
    \Tile_X2Y4_WW4BEG[13] ,
    \Tile_X2Y4_WW4BEG[12] ,
    \Tile_X2Y4_WW4BEG[11] ,
    \Tile_X2Y4_WW4BEG[10] ,
    \Tile_X2Y4_WW4BEG[9] ,
    \Tile_X2Y4_WW4BEG[8] ,
    \Tile_X2Y4_WW4BEG[7] ,
    \Tile_X2Y4_WW4BEG[6] ,
    \Tile_X2Y4_WW4BEG[5] ,
    \Tile_X2Y4_WW4BEG[4] ,
    \Tile_X2Y4_WW4BEG[3] ,
    \Tile_X2Y4_WW4BEG[2] ,
    \Tile_X2Y4_WW4BEG[1] ,
    \Tile_X2Y4_WW4BEG[0] }),
    .WW4END({\Tile_X3Y4_WW4BEG[15] ,
    \Tile_X3Y4_WW4BEG[14] ,
    \Tile_X3Y4_WW4BEG[13] ,
    \Tile_X3Y4_WW4BEG[12] ,
    \Tile_X3Y4_WW4BEG[11] ,
    \Tile_X3Y4_WW4BEG[10] ,
    \Tile_X3Y4_WW4BEG[9] ,
    \Tile_X3Y4_WW4BEG[8] ,
    \Tile_X3Y4_WW4BEG[7] ,
    \Tile_X3Y4_WW4BEG[6] ,
    \Tile_X3Y4_WW4BEG[5] ,
    \Tile_X3Y4_WW4BEG[4] ,
    \Tile_X3Y4_WW4BEG[3] ,
    \Tile_X3Y4_WW4BEG[2] ,
    \Tile_X3Y4_WW4BEG[1] ,
    \Tile_X3Y4_WW4BEG[0] }));
 LUT4AB Tile_X2Y5_LUT4AB (.Ci(Tile_X2Y6_Co),
    .Co(Tile_X2Y5_Co),
    .UserCLK(Tile_X2Y6_UserCLKo),
    .UserCLKo(Tile_X2Y5_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X2Y5_E1BEG[3] ,
    \Tile_X2Y5_E1BEG[2] ,
    \Tile_X2Y5_E1BEG[1] ,
    \Tile_X2Y5_E1BEG[0] }),
    .E1END({\Tile_X1Y5_E1BEG[3] ,
    \Tile_X1Y5_E1BEG[2] ,
    \Tile_X1Y5_E1BEG[1] ,
    \Tile_X1Y5_E1BEG[0] }),
    .E2BEG({\Tile_X2Y5_E2BEG[7] ,
    \Tile_X2Y5_E2BEG[6] ,
    \Tile_X2Y5_E2BEG[5] ,
    \Tile_X2Y5_E2BEG[4] ,
    \Tile_X2Y5_E2BEG[3] ,
    \Tile_X2Y5_E2BEG[2] ,
    \Tile_X2Y5_E2BEG[1] ,
    \Tile_X2Y5_E2BEG[0] }),
    .E2BEGb({\Tile_X2Y5_E2BEGb[7] ,
    \Tile_X2Y5_E2BEGb[6] ,
    \Tile_X2Y5_E2BEGb[5] ,
    \Tile_X2Y5_E2BEGb[4] ,
    \Tile_X2Y5_E2BEGb[3] ,
    \Tile_X2Y5_E2BEGb[2] ,
    \Tile_X2Y5_E2BEGb[1] ,
    \Tile_X2Y5_E2BEGb[0] }),
    .E2END({\Tile_X1Y5_E2BEGb[7] ,
    \Tile_X1Y5_E2BEGb[6] ,
    \Tile_X1Y5_E2BEGb[5] ,
    \Tile_X1Y5_E2BEGb[4] ,
    \Tile_X1Y5_E2BEGb[3] ,
    \Tile_X1Y5_E2BEGb[2] ,
    \Tile_X1Y5_E2BEGb[1] ,
    \Tile_X1Y5_E2BEGb[0] }),
    .E2MID({\Tile_X1Y5_E2BEG[7] ,
    \Tile_X1Y5_E2BEG[6] ,
    \Tile_X1Y5_E2BEG[5] ,
    \Tile_X1Y5_E2BEG[4] ,
    \Tile_X1Y5_E2BEG[3] ,
    \Tile_X1Y5_E2BEG[2] ,
    \Tile_X1Y5_E2BEG[1] ,
    \Tile_X1Y5_E2BEG[0] }),
    .E6BEG({\Tile_X2Y5_E6BEG[11] ,
    \Tile_X2Y5_E6BEG[10] ,
    \Tile_X2Y5_E6BEG[9] ,
    \Tile_X2Y5_E6BEG[8] ,
    \Tile_X2Y5_E6BEG[7] ,
    \Tile_X2Y5_E6BEG[6] ,
    \Tile_X2Y5_E6BEG[5] ,
    \Tile_X2Y5_E6BEG[4] ,
    \Tile_X2Y5_E6BEG[3] ,
    \Tile_X2Y5_E6BEG[2] ,
    \Tile_X2Y5_E6BEG[1] ,
    \Tile_X2Y5_E6BEG[0] }),
    .E6END({\Tile_X1Y5_E6BEG[11] ,
    \Tile_X1Y5_E6BEG[10] ,
    \Tile_X1Y5_E6BEG[9] ,
    \Tile_X1Y5_E6BEG[8] ,
    \Tile_X1Y5_E6BEG[7] ,
    \Tile_X1Y5_E6BEG[6] ,
    \Tile_X1Y5_E6BEG[5] ,
    \Tile_X1Y5_E6BEG[4] ,
    \Tile_X1Y5_E6BEG[3] ,
    \Tile_X1Y5_E6BEG[2] ,
    \Tile_X1Y5_E6BEG[1] ,
    \Tile_X1Y5_E6BEG[0] }),
    .EE4BEG({\Tile_X2Y5_EE4BEG[15] ,
    \Tile_X2Y5_EE4BEG[14] ,
    \Tile_X2Y5_EE4BEG[13] ,
    \Tile_X2Y5_EE4BEG[12] ,
    \Tile_X2Y5_EE4BEG[11] ,
    \Tile_X2Y5_EE4BEG[10] ,
    \Tile_X2Y5_EE4BEG[9] ,
    \Tile_X2Y5_EE4BEG[8] ,
    \Tile_X2Y5_EE4BEG[7] ,
    \Tile_X2Y5_EE4BEG[6] ,
    \Tile_X2Y5_EE4BEG[5] ,
    \Tile_X2Y5_EE4BEG[4] ,
    \Tile_X2Y5_EE4BEG[3] ,
    \Tile_X2Y5_EE4BEG[2] ,
    \Tile_X2Y5_EE4BEG[1] ,
    \Tile_X2Y5_EE4BEG[0] }),
    .EE4END({\Tile_X1Y5_EE4BEG[15] ,
    \Tile_X1Y5_EE4BEG[14] ,
    \Tile_X1Y5_EE4BEG[13] ,
    \Tile_X1Y5_EE4BEG[12] ,
    \Tile_X1Y5_EE4BEG[11] ,
    \Tile_X1Y5_EE4BEG[10] ,
    \Tile_X1Y5_EE4BEG[9] ,
    \Tile_X1Y5_EE4BEG[8] ,
    \Tile_X1Y5_EE4BEG[7] ,
    \Tile_X1Y5_EE4BEG[6] ,
    \Tile_X1Y5_EE4BEG[5] ,
    \Tile_X1Y5_EE4BEG[4] ,
    \Tile_X1Y5_EE4BEG[3] ,
    \Tile_X1Y5_EE4BEG[2] ,
    \Tile_X1Y5_EE4BEG[1] ,
    \Tile_X1Y5_EE4BEG[0] }),
    .FrameData({\Tile_X1Y5_FrameData_O[31] ,
    \Tile_X1Y5_FrameData_O[30] ,
    \Tile_X1Y5_FrameData_O[29] ,
    \Tile_X1Y5_FrameData_O[28] ,
    \Tile_X1Y5_FrameData_O[27] ,
    \Tile_X1Y5_FrameData_O[26] ,
    \Tile_X1Y5_FrameData_O[25] ,
    \Tile_X1Y5_FrameData_O[24] ,
    \Tile_X1Y5_FrameData_O[23] ,
    \Tile_X1Y5_FrameData_O[22] ,
    \Tile_X1Y5_FrameData_O[21] ,
    \Tile_X1Y5_FrameData_O[20] ,
    \Tile_X1Y5_FrameData_O[19] ,
    \Tile_X1Y5_FrameData_O[18] ,
    \Tile_X1Y5_FrameData_O[17] ,
    \Tile_X1Y5_FrameData_O[16] ,
    \Tile_X1Y5_FrameData_O[15] ,
    \Tile_X1Y5_FrameData_O[14] ,
    \Tile_X1Y5_FrameData_O[13] ,
    \Tile_X1Y5_FrameData_O[12] ,
    \Tile_X1Y5_FrameData_O[11] ,
    \Tile_X1Y5_FrameData_O[10] ,
    \Tile_X1Y5_FrameData_O[9] ,
    \Tile_X1Y5_FrameData_O[8] ,
    \Tile_X1Y5_FrameData_O[7] ,
    \Tile_X1Y5_FrameData_O[6] ,
    \Tile_X1Y5_FrameData_O[5] ,
    \Tile_X1Y5_FrameData_O[4] ,
    \Tile_X1Y5_FrameData_O[3] ,
    \Tile_X1Y5_FrameData_O[2] ,
    \Tile_X1Y5_FrameData_O[1] ,
    \Tile_X1Y5_FrameData_O[0] }),
    .FrameData_O({\Tile_X2Y5_FrameData_O[31] ,
    \Tile_X2Y5_FrameData_O[30] ,
    \Tile_X2Y5_FrameData_O[29] ,
    \Tile_X2Y5_FrameData_O[28] ,
    \Tile_X2Y5_FrameData_O[27] ,
    \Tile_X2Y5_FrameData_O[26] ,
    \Tile_X2Y5_FrameData_O[25] ,
    \Tile_X2Y5_FrameData_O[24] ,
    \Tile_X2Y5_FrameData_O[23] ,
    \Tile_X2Y5_FrameData_O[22] ,
    \Tile_X2Y5_FrameData_O[21] ,
    \Tile_X2Y5_FrameData_O[20] ,
    \Tile_X2Y5_FrameData_O[19] ,
    \Tile_X2Y5_FrameData_O[18] ,
    \Tile_X2Y5_FrameData_O[17] ,
    \Tile_X2Y5_FrameData_O[16] ,
    \Tile_X2Y5_FrameData_O[15] ,
    \Tile_X2Y5_FrameData_O[14] ,
    \Tile_X2Y5_FrameData_O[13] ,
    \Tile_X2Y5_FrameData_O[12] ,
    \Tile_X2Y5_FrameData_O[11] ,
    \Tile_X2Y5_FrameData_O[10] ,
    \Tile_X2Y5_FrameData_O[9] ,
    \Tile_X2Y5_FrameData_O[8] ,
    \Tile_X2Y5_FrameData_O[7] ,
    \Tile_X2Y5_FrameData_O[6] ,
    \Tile_X2Y5_FrameData_O[5] ,
    \Tile_X2Y5_FrameData_O[4] ,
    \Tile_X2Y5_FrameData_O[3] ,
    \Tile_X2Y5_FrameData_O[2] ,
    \Tile_X2Y5_FrameData_O[1] ,
    \Tile_X2Y5_FrameData_O[0] }),
    .FrameStrobe({\Tile_X2Y6_FrameStrobe_O[19] ,
    \Tile_X2Y6_FrameStrobe_O[18] ,
    \Tile_X2Y6_FrameStrobe_O[17] ,
    \Tile_X2Y6_FrameStrobe_O[16] ,
    \Tile_X2Y6_FrameStrobe_O[15] ,
    \Tile_X2Y6_FrameStrobe_O[14] ,
    \Tile_X2Y6_FrameStrobe_O[13] ,
    \Tile_X2Y6_FrameStrobe_O[12] ,
    \Tile_X2Y6_FrameStrobe_O[11] ,
    \Tile_X2Y6_FrameStrobe_O[10] ,
    \Tile_X2Y6_FrameStrobe_O[9] ,
    \Tile_X2Y6_FrameStrobe_O[8] ,
    \Tile_X2Y6_FrameStrobe_O[7] ,
    \Tile_X2Y6_FrameStrobe_O[6] ,
    \Tile_X2Y6_FrameStrobe_O[5] ,
    \Tile_X2Y6_FrameStrobe_O[4] ,
    \Tile_X2Y6_FrameStrobe_O[3] ,
    \Tile_X2Y6_FrameStrobe_O[2] ,
    \Tile_X2Y6_FrameStrobe_O[1] ,
    \Tile_X2Y6_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X2Y5_FrameStrobe_O[19] ,
    \Tile_X2Y5_FrameStrobe_O[18] ,
    \Tile_X2Y5_FrameStrobe_O[17] ,
    \Tile_X2Y5_FrameStrobe_O[16] ,
    \Tile_X2Y5_FrameStrobe_O[15] ,
    \Tile_X2Y5_FrameStrobe_O[14] ,
    \Tile_X2Y5_FrameStrobe_O[13] ,
    \Tile_X2Y5_FrameStrobe_O[12] ,
    \Tile_X2Y5_FrameStrobe_O[11] ,
    \Tile_X2Y5_FrameStrobe_O[10] ,
    \Tile_X2Y5_FrameStrobe_O[9] ,
    \Tile_X2Y5_FrameStrobe_O[8] ,
    \Tile_X2Y5_FrameStrobe_O[7] ,
    \Tile_X2Y5_FrameStrobe_O[6] ,
    \Tile_X2Y5_FrameStrobe_O[5] ,
    \Tile_X2Y5_FrameStrobe_O[4] ,
    \Tile_X2Y5_FrameStrobe_O[3] ,
    \Tile_X2Y5_FrameStrobe_O[2] ,
    \Tile_X2Y5_FrameStrobe_O[1] ,
    \Tile_X2Y5_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X2Y5_N1BEG[3] ,
    \Tile_X2Y5_N1BEG[2] ,
    \Tile_X2Y5_N1BEG[1] ,
    \Tile_X2Y5_N1BEG[0] }),
    .N1END({\Tile_X2Y6_N1BEG[3] ,
    \Tile_X2Y6_N1BEG[2] ,
    \Tile_X2Y6_N1BEG[1] ,
    \Tile_X2Y6_N1BEG[0] }),
    .N2BEG({\Tile_X2Y5_N2BEG[7] ,
    \Tile_X2Y5_N2BEG[6] ,
    \Tile_X2Y5_N2BEG[5] ,
    \Tile_X2Y5_N2BEG[4] ,
    \Tile_X2Y5_N2BEG[3] ,
    \Tile_X2Y5_N2BEG[2] ,
    \Tile_X2Y5_N2BEG[1] ,
    \Tile_X2Y5_N2BEG[0] }),
    .N2BEGb({\Tile_X2Y5_N2BEGb[7] ,
    \Tile_X2Y5_N2BEGb[6] ,
    \Tile_X2Y5_N2BEGb[5] ,
    \Tile_X2Y5_N2BEGb[4] ,
    \Tile_X2Y5_N2BEGb[3] ,
    \Tile_X2Y5_N2BEGb[2] ,
    \Tile_X2Y5_N2BEGb[1] ,
    \Tile_X2Y5_N2BEGb[0] }),
    .N2END({\Tile_X2Y6_N2BEGb[7] ,
    \Tile_X2Y6_N2BEGb[6] ,
    \Tile_X2Y6_N2BEGb[5] ,
    \Tile_X2Y6_N2BEGb[4] ,
    \Tile_X2Y6_N2BEGb[3] ,
    \Tile_X2Y6_N2BEGb[2] ,
    \Tile_X2Y6_N2BEGb[1] ,
    \Tile_X2Y6_N2BEGb[0] }),
    .N2MID({\Tile_X2Y6_N2BEG[7] ,
    \Tile_X2Y6_N2BEG[6] ,
    \Tile_X2Y6_N2BEG[5] ,
    \Tile_X2Y6_N2BEG[4] ,
    \Tile_X2Y6_N2BEG[3] ,
    \Tile_X2Y6_N2BEG[2] ,
    \Tile_X2Y6_N2BEG[1] ,
    \Tile_X2Y6_N2BEG[0] }),
    .N4BEG({\Tile_X2Y5_N4BEG[15] ,
    \Tile_X2Y5_N4BEG[14] ,
    \Tile_X2Y5_N4BEG[13] ,
    \Tile_X2Y5_N4BEG[12] ,
    \Tile_X2Y5_N4BEG[11] ,
    \Tile_X2Y5_N4BEG[10] ,
    \Tile_X2Y5_N4BEG[9] ,
    \Tile_X2Y5_N4BEG[8] ,
    \Tile_X2Y5_N4BEG[7] ,
    \Tile_X2Y5_N4BEG[6] ,
    \Tile_X2Y5_N4BEG[5] ,
    \Tile_X2Y5_N4BEG[4] ,
    \Tile_X2Y5_N4BEG[3] ,
    \Tile_X2Y5_N4BEG[2] ,
    \Tile_X2Y5_N4BEG[1] ,
    \Tile_X2Y5_N4BEG[0] }),
    .N4END({\Tile_X2Y6_N4BEG[15] ,
    \Tile_X2Y6_N4BEG[14] ,
    \Tile_X2Y6_N4BEG[13] ,
    \Tile_X2Y6_N4BEG[12] ,
    \Tile_X2Y6_N4BEG[11] ,
    \Tile_X2Y6_N4BEG[10] ,
    \Tile_X2Y6_N4BEG[9] ,
    \Tile_X2Y6_N4BEG[8] ,
    \Tile_X2Y6_N4BEG[7] ,
    \Tile_X2Y6_N4BEG[6] ,
    \Tile_X2Y6_N4BEG[5] ,
    \Tile_X2Y6_N4BEG[4] ,
    \Tile_X2Y6_N4BEG[3] ,
    \Tile_X2Y6_N4BEG[2] ,
    \Tile_X2Y6_N4BEG[1] ,
    \Tile_X2Y6_N4BEG[0] }),
    .NN4BEG({\Tile_X2Y5_NN4BEG[15] ,
    \Tile_X2Y5_NN4BEG[14] ,
    \Tile_X2Y5_NN4BEG[13] ,
    \Tile_X2Y5_NN4BEG[12] ,
    \Tile_X2Y5_NN4BEG[11] ,
    \Tile_X2Y5_NN4BEG[10] ,
    \Tile_X2Y5_NN4BEG[9] ,
    \Tile_X2Y5_NN4BEG[8] ,
    \Tile_X2Y5_NN4BEG[7] ,
    \Tile_X2Y5_NN4BEG[6] ,
    \Tile_X2Y5_NN4BEG[5] ,
    \Tile_X2Y5_NN4BEG[4] ,
    \Tile_X2Y5_NN4BEG[3] ,
    \Tile_X2Y5_NN4BEG[2] ,
    \Tile_X2Y5_NN4BEG[1] ,
    \Tile_X2Y5_NN4BEG[0] }),
    .NN4END({\Tile_X2Y6_NN4BEG[15] ,
    \Tile_X2Y6_NN4BEG[14] ,
    \Tile_X2Y6_NN4BEG[13] ,
    \Tile_X2Y6_NN4BEG[12] ,
    \Tile_X2Y6_NN4BEG[11] ,
    \Tile_X2Y6_NN4BEG[10] ,
    \Tile_X2Y6_NN4BEG[9] ,
    \Tile_X2Y6_NN4BEG[8] ,
    \Tile_X2Y6_NN4BEG[7] ,
    \Tile_X2Y6_NN4BEG[6] ,
    \Tile_X2Y6_NN4BEG[5] ,
    \Tile_X2Y6_NN4BEG[4] ,
    \Tile_X2Y6_NN4BEG[3] ,
    \Tile_X2Y6_NN4BEG[2] ,
    \Tile_X2Y6_NN4BEG[1] ,
    \Tile_X2Y6_NN4BEG[0] }),
    .S1BEG({\Tile_X2Y5_S1BEG[3] ,
    \Tile_X2Y5_S1BEG[2] ,
    \Tile_X2Y5_S1BEG[1] ,
    \Tile_X2Y5_S1BEG[0] }),
    .S1END({\Tile_X2Y4_S1BEG[3] ,
    \Tile_X2Y4_S1BEG[2] ,
    \Tile_X2Y4_S1BEG[1] ,
    \Tile_X2Y4_S1BEG[0] }),
    .S2BEG({\Tile_X2Y5_S2BEG[7] ,
    \Tile_X2Y5_S2BEG[6] ,
    \Tile_X2Y5_S2BEG[5] ,
    \Tile_X2Y5_S2BEG[4] ,
    \Tile_X2Y5_S2BEG[3] ,
    \Tile_X2Y5_S2BEG[2] ,
    \Tile_X2Y5_S2BEG[1] ,
    \Tile_X2Y5_S2BEG[0] }),
    .S2BEGb({\Tile_X2Y5_S2BEGb[7] ,
    \Tile_X2Y5_S2BEGb[6] ,
    \Tile_X2Y5_S2BEGb[5] ,
    \Tile_X2Y5_S2BEGb[4] ,
    \Tile_X2Y5_S2BEGb[3] ,
    \Tile_X2Y5_S2BEGb[2] ,
    \Tile_X2Y5_S2BEGb[1] ,
    \Tile_X2Y5_S2BEGb[0] }),
    .S2END({\Tile_X2Y4_S2BEGb[7] ,
    \Tile_X2Y4_S2BEGb[6] ,
    \Tile_X2Y4_S2BEGb[5] ,
    \Tile_X2Y4_S2BEGb[4] ,
    \Tile_X2Y4_S2BEGb[3] ,
    \Tile_X2Y4_S2BEGb[2] ,
    \Tile_X2Y4_S2BEGb[1] ,
    \Tile_X2Y4_S2BEGb[0] }),
    .S2MID({\Tile_X2Y4_S2BEG[7] ,
    \Tile_X2Y4_S2BEG[6] ,
    \Tile_X2Y4_S2BEG[5] ,
    \Tile_X2Y4_S2BEG[4] ,
    \Tile_X2Y4_S2BEG[3] ,
    \Tile_X2Y4_S2BEG[2] ,
    \Tile_X2Y4_S2BEG[1] ,
    \Tile_X2Y4_S2BEG[0] }),
    .S4BEG({\Tile_X2Y5_S4BEG[15] ,
    \Tile_X2Y5_S4BEG[14] ,
    \Tile_X2Y5_S4BEG[13] ,
    \Tile_X2Y5_S4BEG[12] ,
    \Tile_X2Y5_S4BEG[11] ,
    \Tile_X2Y5_S4BEG[10] ,
    \Tile_X2Y5_S4BEG[9] ,
    \Tile_X2Y5_S4BEG[8] ,
    \Tile_X2Y5_S4BEG[7] ,
    \Tile_X2Y5_S4BEG[6] ,
    \Tile_X2Y5_S4BEG[5] ,
    \Tile_X2Y5_S4BEG[4] ,
    \Tile_X2Y5_S4BEG[3] ,
    \Tile_X2Y5_S4BEG[2] ,
    \Tile_X2Y5_S4BEG[1] ,
    \Tile_X2Y5_S4BEG[0] }),
    .S4END({\Tile_X2Y4_S4BEG[15] ,
    \Tile_X2Y4_S4BEG[14] ,
    \Tile_X2Y4_S4BEG[13] ,
    \Tile_X2Y4_S4BEG[12] ,
    \Tile_X2Y4_S4BEG[11] ,
    \Tile_X2Y4_S4BEG[10] ,
    \Tile_X2Y4_S4BEG[9] ,
    \Tile_X2Y4_S4BEG[8] ,
    \Tile_X2Y4_S4BEG[7] ,
    \Tile_X2Y4_S4BEG[6] ,
    \Tile_X2Y4_S4BEG[5] ,
    \Tile_X2Y4_S4BEG[4] ,
    \Tile_X2Y4_S4BEG[3] ,
    \Tile_X2Y4_S4BEG[2] ,
    \Tile_X2Y4_S4BEG[1] ,
    \Tile_X2Y4_S4BEG[0] }),
    .SS4BEG({\Tile_X2Y5_SS4BEG[15] ,
    \Tile_X2Y5_SS4BEG[14] ,
    \Tile_X2Y5_SS4BEG[13] ,
    \Tile_X2Y5_SS4BEG[12] ,
    \Tile_X2Y5_SS4BEG[11] ,
    \Tile_X2Y5_SS4BEG[10] ,
    \Tile_X2Y5_SS4BEG[9] ,
    \Tile_X2Y5_SS4BEG[8] ,
    \Tile_X2Y5_SS4BEG[7] ,
    \Tile_X2Y5_SS4BEG[6] ,
    \Tile_X2Y5_SS4BEG[5] ,
    \Tile_X2Y5_SS4BEG[4] ,
    \Tile_X2Y5_SS4BEG[3] ,
    \Tile_X2Y5_SS4BEG[2] ,
    \Tile_X2Y5_SS4BEG[1] ,
    \Tile_X2Y5_SS4BEG[0] }),
    .SS4END({\Tile_X2Y4_SS4BEG[15] ,
    \Tile_X2Y4_SS4BEG[14] ,
    \Tile_X2Y4_SS4BEG[13] ,
    \Tile_X2Y4_SS4BEG[12] ,
    \Tile_X2Y4_SS4BEG[11] ,
    \Tile_X2Y4_SS4BEG[10] ,
    \Tile_X2Y4_SS4BEG[9] ,
    \Tile_X2Y4_SS4BEG[8] ,
    \Tile_X2Y4_SS4BEG[7] ,
    \Tile_X2Y4_SS4BEG[6] ,
    \Tile_X2Y4_SS4BEG[5] ,
    \Tile_X2Y4_SS4BEG[4] ,
    \Tile_X2Y4_SS4BEG[3] ,
    \Tile_X2Y4_SS4BEG[2] ,
    \Tile_X2Y4_SS4BEG[1] ,
    \Tile_X2Y4_SS4BEG[0] }),
    .W1BEG({\Tile_X2Y5_W1BEG[3] ,
    \Tile_X2Y5_W1BEG[2] ,
    \Tile_X2Y5_W1BEG[1] ,
    \Tile_X2Y5_W1BEG[0] }),
    .W1END({\Tile_X3Y5_W1BEG[3] ,
    \Tile_X3Y5_W1BEG[2] ,
    \Tile_X3Y5_W1BEG[1] ,
    \Tile_X3Y5_W1BEG[0] }),
    .W2BEG({\Tile_X2Y5_W2BEG[7] ,
    \Tile_X2Y5_W2BEG[6] ,
    \Tile_X2Y5_W2BEG[5] ,
    \Tile_X2Y5_W2BEG[4] ,
    \Tile_X2Y5_W2BEG[3] ,
    \Tile_X2Y5_W2BEG[2] ,
    \Tile_X2Y5_W2BEG[1] ,
    \Tile_X2Y5_W2BEG[0] }),
    .W2BEGb({\Tile_X2Y5_W2BEGb[7] ,
    \Tile_X2Y5_W2BEGb[6] ,
    \Tile_X2Y5_W2BEGb[5] ,
    \Tile_X2Y5_W2BEGb[4] ,
    \Tile_X2Y5_W2BEGb[3] ,
    \Tile_X2Y5_W2BEGb[2] ,
    \Tile_X2Y5_W2BEGb[1] ,
    \Tile_X2Y5_W2BEGb[0] }),
    .W2END({\Tile_X3Y5_W2BEGb[7] ,
    \Tile_X3Y5_W2BEGb[6] ,
    \Tile_X3Y5_W2BEGb[5] ,
    \Tile_X3Y5_W2BEGb[4] ,
    \Tile_X3Y5_W2BEGb[3] ,
    \Tile_X3Y5_W2BEGb[2] ,
    \Tile_X3Y5_W2BEGb[1] ,
    \Tile_X3Y5_W2BEGb[0] }),
    .W2MID({\Tile_X3Y5_W2BEG[7] ,
    \Tile_X3Y5_W2BEG[6] ,
    \Tile_X3Y5_W2BEG[5] ,
    \Tile_X3Y5_W2BEG[4] ,
    \Tile_X3Y5_W2BEG[3] ,
    \Tile_X3Y5_W2BEG[2] ,
    \Tile_X3Y5_W2BEG[1] ,
    \Tile_X3Y5_W2BEG[0] }),
    .W6BEG({\Tile_X2Y5_W6BEG[11] ,
    \Tile_X2Y5_W6BEG[10] ,
    \Tile_X2Y5_W6BEG[9] ,
    \Tile_X2Y5_W6BEG[8] ,
    \Tile_X2Y5_W6BEG[7] ,
    \Tile_X2Y5_W6BEG[6] ,
    \Tile_X2Y5_W6BEG[5] ,
    \Tile_X2Y5_W6BEG[4] ,
    \Tile_X2Y5_W6BEG[3] ,
    \Tile_X2Y5_W6BEG[2] ,
    \Tile_X2Y5_W6BEG[1] ,
    \Tile_X2Y5_W6BEG[0] }),
    .W6END({\Tile_X3Y5_W6BEG[11] ,
    \Tile_X3Y5_W6BEG[10] ,
    \Tile_X3Y5_W6BEG[9] ,
    \Tile_X3Y5_W6BEG[8] ,
    \Tile_X3Y5_W6BEG[7] ,
    \Tile_X3Y5_W6BEG[6] ,
    \Tile_X3Y5_W6BEG[5] ,
    \Tile_X3Y5_W6BEG[4] ,
    \Tile_X3Y5_W6BEG[3] ,
    \Tile_X3Y5_W6BEG[2] ,
    \Tile_X3Y5_W6BEG[1] ,
    \Tile_X3Y5_W6BEG[0] }),
    .WW4BEG({\Tile_X2Y5_WW4BEG[15] ,
    \Tile_X2Y5_WW4BEG[14] ,
    \Tile_X2Y5_WW4BEG[13] ,
    \Tile_X2Y5_WW4BEG[12] ,
    \Tile_X2Y5_WW4BEG[11] ,
    \Tile_X2Y5_WW4BEG[10] ,
    \Tile_X2Y5_WW4BEG[9] ,
    \Tile_X2Y5_WW4BEG[8] ,
    \Tile_X2Y5_WW4BEG[7] ,
    \Tile_X2Y5_WW4BEG[6] ,
    \Tile_X2Y5_WW4BEG[5] ,
    \Tile_X2Y5_WW4BEG[4] ,
    \Tile_X2Y5_WW4BEG[3] ,
    \Tile_X2Y5_WW4BEG[2] ,
    \Tile_X2Y5_WW4BEG[1] ,
    \Tile_X2Y5_WW4BEG[0] }),
    .WW4END({\Tile_X3Y5_WW4BEG[15] ,
    \Tile_X3Y5_WW4BEG[14] ,
    \Tile_X3Y5_WW4BEG[13] ,
    \Tile_X3Y5_WW4BEG[12] ,
    \Tile_X3Y5_WW4BEG[11] ,
    \Tile_X3Y5_WW4BEG[10] ,
    \Tile_X3Y5_WW4BEG[9] ,
    \Tile_X3Y5_WW4BEG[8] ,
    \Tile_X3Y5_WW4BEG[7] ,
    \Tile_X3Y5_WW4BEG[6] ,
    \Tile_X3Y5_WW4BEG[5] ,
    \Tile_X3Y5_WW4BEG[4] ,
    \Tile_X3Y5_WW4BEG[3] ,
    \Tile_X3Y5_WW4BEG[2] ,
    \Tile_X3Y5_WW4BEG[1] ,
    \Tile_X3Y5_WW4BEG[0] }));
 LUT4AB Tile_X2Y6_LUT4AB (.Ci(Tile_X2Y7_Co),
    .Co(Tile_X2Y6_Co),
    .UserCLK(Tile_X2Y7_UserCLKo),
    .UserCLKo(Tile_X2Y6_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X2Y6_E1BEG[3] ,
    \Tile_X2Y6_E1BEG[2] ,
    \Tile_X2Y6_E1BEG[1] ,
    \Tile_X2Y6_E1BEG[0] }),
    .E1END({\Tile_X1Y6_E1BEG[3] ,
    \Tile_X1Y6_E1BEG[2] ,
    \Tile_X1Y6_E1BEG[1] ,
    \Tile_X1Y6_E1BEG[0] }),
    .E2BEG({\Tile_X2Y6_E2BEG[7] ,
    \Tile_X2Y6_E2BEG[6] ,
    \Tile_X2Y6_E2BEG[5] ,
    \Tile_X2Y6_E2BEG[4] ,
    \Tile_X2Y6_E2BEG[3] ,
    \Tile_X2Y6_E2BEG[2] ,
    \Tile_X2Y6_E2BEG[1] ,
    \Tile_X2Y6_E2BEG[0] }),
    .E2BEGb({\Tile_X2Y6_E2BEGb[7] ,
    \Tile_X2Y6_E2BEGb[6] ,
    \Tile_X2Y6_E2BEGb[5] ,
    \Tile_X2Y6_E2BEGb[4] ,
    \Tile_X2Y6_E2BEGb[3] ,
    \Tile_X2Y6_E2BEGb[2] ,
    \Tile_X2Y6_E2BEGb[1] ,
    \Tile_X2Y6_E2BEGb[0] }),
    .E2END({\Tile_X1Y6_E2BEGb[7] ,
    \Tile_X1Y6_E2BEGb[6] ,
    \Tile_X1Y6_E2BEGb[5] ,
    \Tile_X1Y6_E2BEGb[4] ,
    \Tile_X1Y6_E2BEGb[3] ,
    \Tile_X1Y6_E2BEGb[2] ,
    \Tile_X1Y6_E2BEGb[1] ,
    \Tile_X1Y6_E2BEGb[0] }),
    .E2MID({\Tile_X1Y6_E2BEG[7] ,
    \Tile_X1Y6_E2BEG[6] ,
    \Tile_X1Y6_E2BEG[5] ,
    \Tile_X1Y6_E2BEG[4] ,
    \Tile_X1Y6_E2BEG[3] ,
    \Tile_X1Y6_E2BEG[2] ,
    \Tile_X1Y6_E2BEG[1] ,
    \Tile_X1Y6_E2BEG[0] }),
    .E6BEG({\Tile_X2Y6_E6BEG[11] ,
    \Tile_X2Y6_E6BEG[10] ,
    \Tile_X2Y6_E6BEG[9] ,
    \Tile_X2Y6_E6BEG[8] ,
    \Tile_X2Y6_E6BEG[7] ,
    \Tile_X2Y6_E6BEG[6] ,
    \Tile_X2Y6_E6BEG[5] ,
    \Tile_X2Y6_E6BEG[4] ,
    \Tile_X2Y6_E6BEG[3] ,
    \Tile_X2Y6_E6BEG[2] ,
    \Tile_X2Y6_E6BEG[1] ,
    \Tile_X2Y6_E6BEG[0] }),
    .E6END({\Tile_X1Y6_E6BEG[11] ,
    \Tile_X1Y6_E6BEG[10] ,
    \Tile_X1Y6_E6BEG[9] ,
    \Tile_X1Y6_E6BEG[8] ,
    \Tile_X1Y6_E6BEG[7] ,
    \Tile_X1Y6_E6BEG[6] ,
    \Tile_X1Y6_E6BEG[5] ,
    \Tile_X1Y6_E6BEG[4] ,
    \Tile_X1Y6_E6BEG[3] ,
    \Tile_X1Y6_E6BEG[2] ,
    \Tile_X1Y6_E6BEG[1] ,
    \Tile_X1Y6_E6BEG[0] }),
    .EE4BEG({\Tile_X2Y6_EE4BEG[15] ,
    \Tile_X2Y6_EE4BEG[14] ,
    \Tile_X2Y6_EE4BEG[13] ,
    \Tile_X2Y6_EE4BEG[12] ,
    \Tile_X2Y6_EE4BEG[11] ,
    \Tile_X2Y6_EE4BEG[10] ,
    \Tile_X2Y6_EE4BEG[9] ,
    \Tile_X2Y6_EE4BEG[8] ,
    \Tile_X2Y6_EE4BEG[7] ,
    \Tile_X2Y6_EE4BEG[6] ,
    \Tile_X2Y6_EE4BEG[5] ,
    \Tile_X2Y6_EE4BEG[4] ,
    \Tile_X2Y6_EE4BEG[3] ,
    \Tile_X2Y6_EE4BEG[2] ,
    \Tile_X2Y6_EE4BEG[1] ,
    \Tile_X2Y6_EE4BEG[0] }),
    .EE4END({\Tile_X1Y6_EE4BEG[15] ,
    \Tile_X1Y6_EE4BEG[14] ,
    \Tile_X1Y6_EE4BEG[13] ,
    \Tile_X1Y6_EE4BEG[12] ,
    \Tile_X1Y6_EE4BEG[11] ,
    \Tile_X1Y6_EE4BEG[10] ,
    \Tile_X1Y6_EE4BEG[9] ,
    \Tile_X1Y6_EE4BEG[8] ,
    \Tile_X1Y6_EE4BEG[7] ,
    \Tile_X1Y6_EE4BEG[6] ,
    \Tile_X1Y6_EE4BEG[5] ,
    \Tile_X1Y6_EE4BEG[4] ,
    \Tile_X1Y6_EE4BEG[3] ,
    \Tile_X1Y6_EE4BEG[2] ,
    \Tile_X1Y6_EE4BEG[1] ,
    \Tile_X1Y6_EE4BEG[0] }),
    .FrameData({\Tile_X1Y6_FrameData_O[31] ,
    \Tile_X1Y6_FrameData_O[30] ,
    \Tile_X1Y6_FrameData_O[29] ,
    \Tile_X1Y6_FrameData_O[28] ,
    \Tile_X1Y6_FrameData_O[27] ,
    \Tile_X1Y6_FrameData_O[26] ,
    \Tile_X1Y6_FrameData_O[25] ,
    \Tile_X1Y6_FrameData_O[24] ,
    \Tile_X1Y6_FrameData_O[23] ,
    \Tile_X1Y6_FrameData_O[22] ,
    \Tile_X1Y6_FrameData_O[21] ,
    \Tile_X1Y6_FrameData_O[20] ,
    \Tile_X1Y6_FrameData_O[19] ,
    \Tile_X1Y6_FrameData_O[18] ,
    \Tile_X1Y6_FrameData_O[17] ,
    \Tile_X1Y6_FrameData_O[16] ,
    \Tile_X1Y6_FrameData_O[15] ,
    \Tile_X1Y6_FrameData_O[14] ,
    \Tile_X1Y6_FrameData_O[13] ,
    \Tile_X1Y6_FrameData_O[12] ,
    \Tile_X1Y6_FrameData_O[11] ,
    \Tile_X1Y6_FrameData_O[10] ,
    \Tile_X1Y6_FrameData_O[9] ,
    \Tile_X1Y6_FrameData_O[8] ,
    \Tile_X1Y6_FrameData_O[7] ,
    \Tile_X1Y6_FrameData_O[6] ,
    \Tile_X1Y6_FrameData_O[5] ,
    \Tile_X1Y6_FrameData_O[4] ,
    \Tile_X1Y6_FrameData_O[3] ,
    \Tile_X1Y6_FrameData_O[2] ,
    \Tile_X1Y6_FrameData_O[1] ,
    \Tile_X1Y6_FrameData_O[0] }),
    .FrameData_O({\Tile_X2Y6_FrameData_O[31] ,
    \Tile_X2Y6_FrameData_O[30] ,
    \Tile_X2Y6_FrameData_O[29] ,
    \Tile_X2Y6_FrameData_O[28] ,
    \Tile_X2Y6_FrameData_O[27] ,
    \Tile_X2Y6_FrameData_O[26] ,
    \Tile_X2Y6_FrameData_O[25] ,
    \Tile_X2Y6_FrameData_O[24] ,
    \Tile_X2Y6_FrameData_O[23] ,
    \Tile_X2Y6_FrameData_O[22] ,
    \Tile_X2Y6_FrameData_O[21] ,
    \Tile_X2Y6_FrameData_O[20] ,
    \Tile_X2Y6_FrameData_O[19] ,
    \Tile_X2Y6_FrameData_O[18] ,
    \Tile_X2Y6_FrameData_O[17] ,
    \Tile_X2Y6_FrameData_O[16] ,
    \Tile_X2Y6_FrameData_O[15] ,
    \Tile_X2Y6_FrameData_O[14] ,
    \Tile_X2Y6_FrameData_O[13] ,
    \Tile_X2Y6_FrameData_O[12] ,
    \Tile_X2Y6_FrameData_O[11] ,
    \Tile_X2Y6_FrameData_O[10] ,
    \Tile_X2Y6_FrameData_O[9] ,
    \Tile_X2Y6_FrameData_O[8] ,
    \Tile_X2Y6_FrameData_O[7] ,
    \Tile_X2Y6_FrameData_O[6] ,
    \Tile_X2Y6_FrameData_O[5] ,
    \Tile_X2Y6_FrameData_O[4] ,
    \Tile_X2Y6_FrameData_O[3] ,
    \Tile_X2Y6_FrameData_O[2] ,
    \Tile_X2Y6_FrameData_O[1] ,
    \Tile_X2Y6_FrameData_O[0] }),
    .FrameStrobe({\Tile_X2Y7_FrameStrobe_O[19] ,
    \Tile_X2Y7_FrameStrobe_O[18] ,
    \Tile_X2Y7_FrameStrobe_O[17] ,
    \Tile_X2Y7_FrameStrobe_O[16] ,
    \Tile_X2Y7_FrameStrobe_O[15] ,
    \Tile_X2Y7_FrameStrobe_O[14] ,
    \Tile_X2Y7_FrameStrobe_O[13] ,
    \Tile_X2Y7_FrameStrobe_O[12] ,
    \Tile_X2Y7_FrameStrobe_O[11] ,
    \Tile_X2Y7_FrameStrobe_O[10] ,
    \Tile_X2Y7_FrameStrobe_O[9] ,
    \Tile_X2Y7_FrameStrobe_O[8] ,
    \Tile_X2Y7_FrameStrobe_O[7] ,
    \Tile_X2Y7_FrameStrobe_O[6] ,
    \Tile_X2Y7_FrameStrobe_O[5] ,
    \Tile_X2Y7_FrameStrobe_O[4] ,
    \Tile_X2Y7_FrameStrobe_O[3] ,
    \Tile_X2Y7_FrameStrobe_O[2] ,
    \Tile_X2Y7_FrameStrobe_O[1] ,
    \Tile_X2Y7_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X2Y6_FrameStrobe_O[19] ,
    \Tile_X2Y6_FrameStrobe_O[18] ,
    \Tile_X2Y6_FrameStrobe_O[17] ,
    \Tile_X2Y6_FrameStrobe_O[16] ,
    \Tile_X2Y6_FrameStrobe_O[15] ,
    \Tile_X2Y6_FrameStrobe_O[14] ,
    \Tile_X2Y6_FrameStrobe_O[13] ,
    \Tile_X2Y6_FrameStrobe_O[12] ,
    \Tile_X2Y6_FrameStrobe_O[11] ,
    \Tile_X2Y6_FrameStrobe_O[10] ,
    \Tile_X2Y6_FrameStrobe_O[9] ,
    \Tile_X2Y6_FrameStrobe_O[8] ,
    \Tile_X2Y6_FrameStrobe_O[7] ,
    \Tile_X2Y6_FrameStrobe_O[6] ,
    \Tile_X2Y6_FrameStrobe_O[5] ,
    \Tile_X2Y6_FrameStrobe_O[4] ,
    \Tile_X2Y6_FrameStrobe_O[3] ,
    \Tile_X2Y6_FrameStrobe_O[2] ,
    \Tile_X2Y6_FrameStrobe_O[1] ,
    \Tile_X2Y6_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X2Y6_N1BEG[3] ,
    \Tile_X2Y6_N1BEG[2] ,
    \Tile_X2Y6_N1BEG[1] ,
    \Tile_X2Y6_N1BEG[0] }),
    .N1END({\Tile_X2Y7_N1BEG[3] ,
    \Tile_X2Y7_N1BEG[2] ,
    \Tile_X2Y7_N1BEG[1] ,
    \Tile_X2Y7_N1BEG[0] }),
    .N2BEG({\Tile_X2Y6_N2BEG[7] ,
    \Tile_X2Y6_N2BEG[6] ,
    \Tile_X2Y6_N2BEG[5] ,
    \Tile_X2Y6_N2BEG[4] ,
    \Tile_X2Y6_N2BEG[3] ,
    \Tile_X2Y6_N2BEG[2] ,
    \Tile_X2Y6_N2BEG[1] ,
    \Tile_X2Y6_N2BEG[0] }),
    .N2BEGb({\Tile_X2Y6_N2BEGb[7] ,
    \Tile_X2Y6_N2BEGb[6] ,
    \Tile_X2Y6_N2BEGb[5] ,
    \Tile_X2Y6_N2BEGb[4] ,
    \Tile_X2Y6_N2BEGb[3] ,
    \Tile_X2Y6_N2BEGb[2] ,
    \Tile_X2Y6_N2BEGb[1] ,
    \Tile_X2Y6_N2BEGb[0] }),
    .N2END({\Tile_X2Y7_N2BEGb[7] ,
    \Tile_X2Y7_N2BEGb[6] ,
    \Tile_X2Y7_N2BEGb[5] ,
    \Tile_X2Y7_N2BEGb[4] ,
    \Tile_X2Y7_N2BEGb[3] ,
    \Tile_X2Y7_N2BEGb[2] ,
    \Tile_X2Y7_N2BEGb[1] ,
    \Tile_X2Y7_N2BEGb[0] }),
    .N2MID({\Tile_X2Y7_N2BEG[7] ,
    \Tile_X2Y7_N2BEG[6] ,
    \Tile_X2Y7_N2BEG[5] ,
    \Tile_X2Y7_N2BEG[4] ,
    \Tile_X2Y7_N2BEG[3] ,
    \Tile_X2Y7_N2BEG[2] ,
    \Tile_X2Y7_N2BEG[1] ,
    \Tile_X2Y7_N2BEG[0] }),
    .N4BEG({\Tile_X2Y6_N4BEG[15] ,
    \Tile_X2Y6_N4BEG[14] ,
    \Tile_X2Y6_N4BEG[13] ,
    \Tile_X2Y6_N4BEG[12] ,
    \Tile_X2Y6_N4BEG[11] ,
    \Tile_X2Y6_N4BEG[10] ,
    \Tile_X2Y6_N4BEG[9] ,
    \Tile_X2Y6_N4BEG[8] ,
    \Tile_X2Y6_N4BEG[7] ,
    \Tile_X2Y6_N4BEG[6] ,
    \Tile_X2Y6_N4BEG[5] ,
    \Tile_X2Y6_N4BEG[4] ,
    \Tile_X2Y6_N4BEG[3] ,
    \Tile_X2Y6_N4BEG[2] ,
    \Tile_X2Y6_N4BEG[1] ,
    \Tile_X2Y6_N4BEG[0] }),
    .N4END({\Tile_X2Y7_N4BEG[15] ,
    \Tile_X2Y7_N4BEG[14] ,
    \Tile_X2Y7_N4BEG[13] ,
    \Tile_X2Y7_N4BEG[12] ,
    \Tile_X2Y7_N4BEG[11] ,
    \Tile_X2Y7_N4BEG[10] ,
    \Tile_X2Y7_N4BEG[9] ,
    \Tile_X2Y7_N4BEG[8] ,
    \Tile_X2Y7_N4BEG[7] ,
    \Tile_X2Y7_N4BEG[6] ,
    \Tile_X2Y7_N4BEG[5] ,
    \Tile_X2Y7_N4BEG[4] ,
    \Tile_X2Y7_N4BEG[3] ,
    \Tile_X2Y7_N4BEG[2] ,
    \Tile_X2Y7_N4BEG[1] ,
    \Tile_X2Y7_N4BEG[0] }),
    .NN4BEG({\Tile_X2Y6_NN4BEG[15] ,
    \Tile_X2Y6_NN4BEG[14] ,
    \Tile_X2Y6_NN4BEG[13] ,
    \Tile_X2Y6_NN4BEG[12] ,
    \Tile_X2Y6_NN4BEG[11] ,
    \Tile_X2Y6_NN4BEG[10] ,
    \Tile_X2Y6_NN4BEG[9] ,
    \Tile_X2Y6_NN4BEG[8] ,
    \Tile_X2Y6_NN4BEG[7] ,
    \Tile_X2Y6_NN4BEG[6] ,
    \Tile_X2Y6_NN4BEG[5] ,
    \Tile_X2Y6_NN4BEG[4] ,
    \Tile_X2Y6_NN4BEG[3] ,
    \Tile_X2Y6_NN4BEG[2] ,
    \Tile_X2Y6_NN4BEG[1] ,
    \Tile_X2Y6_NN4BEG[0] }),
    .NN4END({\Tile_X2Y7_NN4BEG[15] ,
    \Tile_X2Y7_NN4BEG[14] ,
    \Tile_X2Y7_NN4BEG[13] ,
    \Tile_X2Y7_NN4BEG[12] ,
    \Tile_X2Y7_NN4BEG[11] ,
    \Tile_X2Y7_NN4BEG[10] ,
    \Tile_X2Y7_NN4BEG[9] ,
    \Tile_X2Y7_NN4BEG[8] ,
    \Tile_X2Y7_NN4BEG[7] ,
    \Tile_X2Y7_NN4BEG[6] ,
    \Tile_X2Y7_NN4BEG[5] ,
    \Tile_X2Y7_NN4BEG[4] ,
    \Tile_X2Y7_NN4BEG[3] ,
    \Tile_X2Y7_NN4BEG[2] ,
    \Tile_X2Y7_NN4BEG[1] ,
    \Tile_X2Y7_NN4BEG[0] }),
    .S1BEG({\Tile_X2Y6_S1BEG[3] ,
    \Tile_X2Y6_S1BEG[2] ,
    \Tile_X2Y6_S1BEG[1] ,
    \Tile_X2Y6_S1BEG[0] }),
    .S1END({\Tile_X2Y5_S1BEG[3] ,
    \Tile_X2Y5_S1BEG[2] ,
    \Tile_X2Y5_S1BEG[1] ,
    \Tile_X2Y5_S1BEG[0] }),
    .S2BEG({\Tile_X2Y6_S2BEG[7] ,
    \Tile_X2Y6_S2BEG[6] ,
    \Tile_X2Y6_S2BEG[5] ,
    \Tile_X2Y6_S2BEG[4] ,
    \Tile_X2Y6_S2BEG[3] ,
    \Tile_X2Y6_S2BEG[2] ,
    \Tile_X2Y6_S2BEG[1] ,
    \Tile_X2Y6_S2BEG[0] }),
    .S2BEGb({\Tile_X2Y6_S2BEGb[7] ,
    \Tile_X2Y6_S2BEGb[6] ,
    \Tile_X2Y6_S2BEGb[5] ,
    \Tile_X2Y6_S2BEGb[4] ,
    \Tile_X2Y6_S2BEGb[3] ,
    \Tile_X2Y6_S2BEGb[2] ,
    \Tile_X2Y6_S2BEGb[1] ,
    \Tile_X2Y6_S2BEGb[0] }),
    .S2END({\Tile_X2Y5_S2BEGb[7] ,
    \Tile_X2Y5_S2BEGb[6] ,
    \Tile_X2Y5_S2BEGb[5] ,
    \Tile_X2Y5_S2BEGb[4] ,
    \Tile_X2Y5_S2BEGb[3] ,
    \Tile_X2Y5_S2BEGb[2] ,
    \Tile_X2Y5_S2BEGb[1] ,
    \Tile_X2Y5_S2BEGb[0] }),
    .S2MID({\Tile_X2Y5_S2BEG[7] ,
    \Tile_X2Y5_S2BEG[6] ,
    \Tile_X2Y5_S2BEG[5] ,
    \Tile_X2Y5_S2BEG[4] ,
    \Tile_X2Y5_S2BEG[3] ,
    \Tile_X2Y5_S2BEG[2] ,
    \Tile_X2Y5_S2BEG[1] ,
    \Tile_X2Y5_S2BEG[0] }),
    .S4BEG({\Tile_X2Y6_S4BEG[15] ,
    \Tile_X2Y6_S4BEG[14] ,
    \Tile_X2Y6_S4BEG[13] ,
    \Tile_X2Y6_S4BEG[12] ,
    \Tile_X2Y6_S4BEG[11] ,
    \Tile_X2Y6_S4BEG[10] ,
    \Tile_X2Y6_S4BEG[9] ,
    \Tile_X2Y6_S4BEG[8] ,
    \Tile_X2Y6_S4BEG[7] ,
    \Tile_X2Y6_S4BEG[6] ,
    \Tile_X2Y6_S4BEG[5] ,
    \Tile_X2Y6_S4BEG[4] ,
    \Tile_X2Y6_S4BEG[3] ,
    \Tile_X2Y6_S4BEG[2] ,
    \Tile_X2Y6_S4BEG[1] ,
    \Tile_X2Y6_S4BEG[0] }),
    .S4END({\Tile_X2Y5_S4BEG[15] ,
    \Tile_X2Y5_S4BEG[14] ,
    \Tile_X2Y5_S4BEG[13] ,
    \Tile_X2Y5_S4BEG[12] ,
    \Tile_X2Y5_S4BEG[11] ,
    \Tile_X2Y5_S4BEG[10] ,
    \Tile_X2Y5_S4BEG[9] ,
    \Tile_X2Y5_S4BEG[8] ,
    \Tile_X2Y5_S4BEG[7] ,
    \Tile_X2Y5_S4BEG[6] ,
    \Tile_X2Y5_S4BEG[5] ,
    \Tile_X2Y5_S4BEG[4] ,
    \Tile_X2Y5_S4BEG[3] ,
    \Tile_X2Y5_S4BEG[2] ,
    \Tile_X2Y5_S4BEG[1] ,
    \Tile_X2Y5_S4BEG[0] }),
    .SS4BEG({\Tile_X2Y6_SS4BEG[15] ,
    \Tile_X2Y6_SS4BEG[14] ,
    \Tile_X2Y6_SS4BEG[13] ,
    \Tile_X2Y6_SS4BEG[12] ,
    \Tile_X2Y6_SS4BEG[11] ,
    \Tile_X2Y6_SS4BEG[10] ,
    \Tile_X2Y6_SS4BEG[9] ,
    \Tile_X2Y6_SS4BEG[8] ,
    \Tile_X2Y6_SS4BEG[7] ,
    \Tile_X2Y6_SS4BEG[6] ,
    \Tile_X2Y6_SS4BEG[5] ,
    \Tile_X2Y6_SS4BEG[4] ,
    \Tile_X2Y6_SS4BEG[3] ,
    \Tile_X2Y6_SS4BEG[2] ,
    \Tile_X2Y6_SS4BEG[1] ,
    \Tile_X2Y6_SS4BEG[0] }),
    .SS4END({\Tile_X2Y5_SS4BEG[15] ,
    \Tile_X2Y5_SS4BEG[14] ,
    \Tile_X2Y5_SS4BEG[13] ,
    \Tile_X2Y5_SS4BEG[12] ,
    \Tile_X2Y5_SS4BEG[11] ,
    \Tile_X2Y5_SS4BEG[10] ,
    \Tile_X2Y5_SS4BEG[9] ,
    \Tile_X2Y5_SS4BEG[8] ,
    \Tile_X2Y5_SS4BEG[7] ,
    \Tile_X2Y5_SS4BEG[6] ,
    \Tile_X2Y5_SS4BEG[5] ,
    \Tile_X2Y5_SS4BEG[4] ,
    \Tile_X2Y5_SS4BEG[3] ,
    \Tile_X2Y5_SS4BEG[2] ,
    \Tile_X2Y5_SS4BEG[1] ,
    \Tile_X2Y5_SS4BEG[0] }),
    .W1BEG({\Tile_X2Y6_W1BEG[3] ,
    \Tile_X2Y6_W1BEG[2] ,
    \Tile_X2Y6_W1BEG[1] ,
    \Tile_X2Y6_W1BEG[0] }),
    .W1END({\Tile_X3Y6_W1BEG[3] ,
    \Tile_X3Y6_W1BEG[2] ,
    \Tile_X3Y6_W1BEG[1] ,
    \Tile_X3Y6_W1BEG[0] }),
    .W2BEG({\Tile_X2Y6_W2BEG[7] ,
    \Tile_X2Y6_W2BEG[6] ,
    \Tile_X2Y6_W2BEG[5] ,
    \Tile_X2Y6_W2BEG[4] ,
    \Tile_X2Y6_W2BEG[3] ,
    \Tile_X2Y6_W2BEG[2] ,
    \Tile_X2Y6_W2BEG[1] ,
    \Tile_X2Y6_W2BEG[0] }),
    .W2BEGb({\Tile_X2Y6_W2BEGb[7] ,
    \Tile_X2Y6_W2BEGb[6] ,
    \Tile_X2Y6_W2BEGb[5] ,
    \Tile_X2Y6_W2BEGb[4] ,
    \Tile_X2Y6_W2BEGb[3] ,
    \Tile_X2Y6_W2BEGb[2] ,
    \Tile_X2Y6_W2BEGb[1] ,
    \Tile_X2Y6_W2BEGb[0] }),
    .W2END({\Tile_X3Y6_W2BEGb[7] ,
    \Tile_X3Y6_W2BEGb[6] ,
    \Tile_X3Y6_W2BEGb[5] ,
    \Tile_X3Y6_W2BEGb[4] ,
    \Tile_X3Y6_W2BEGb[3] ,
    \Tile_X3Y6_W2BEGb[2] ,
    \Tile_X3Y6_W2BEGb[1] ,
    \Tile_X3Y6_W2BEGb[0] }),
    .W2MID({\Tile_X3Y6_W2BEG[7] ,
    \Tile_X3Y6_W2BEG[6] ,
    \Tile_X3Y6_W2BEG[5] ,
    \Tile_X3Y6_W2BEG[4] ,
    \Tile_X3Y6_W2BEG[3] ,
    \Tile_X3Y6_W2BEG[2] ,
    \Tile_X3Y6_W2BEG[1] ,
    \Tile_X3Y6_W2BEG[0] }),
    .W6BEG({\Tile_X2Y6_W6BEG[11] ,
    \Tile_X2Y6_W6BEG[10] ,
    \Tile_X2Y6_W6BEG[9] ,
    \Tile_X2Y6_W6BEG[8] ,
    \Tile_X2Y6_W6BEG[7] ,
    \Tile_X2Y6_W6BEG[6] ,
    \Tile_X2Y6_W6BEG[5] ,
    \Tile_X2Y6_W6BEG[4] ,
    \Tile_X2Y6_W6BEG[3] ,
    \Tile_X2Y6_W6BEG[2] ,
    \Tile_X2Y6_W6BEG[1] ,
    \Tile_X2Y6_W6BEG[0] }),
    .W6END({\Tile_X3Y6_W6BEG[11] ,
    \Tile_X3Y6_W6BEG[10] ,
    \Tile_X3Y6_W6BEG[9] ,
    \Tile_X3Y6_W6BEG[8] ,
    \Tile_X3Y6_W6BEG[7] ,
    \Tile_X3Y6_W6BEG[6] ,
    \Tile_X3Y6_W6BEG[5] ,
    \Tile_X3Y6_W6BEG[4] ,
    \Tile_X3Y6_W6BEG[3] ,
    \Tile_X3Y6_W6BEG[2] ,
    \Tile_X3Y6_W6BEG[1] ,
    \Tile_X3Y6_W6BEG[0] }),
    .WW4BEG({\Tile_X2Y6_WW4BEG[15] ,
    \Tile_X2Y6_WW4BEG[14] ,
    \Tile_X2Y6_WW4BEG[13] ,
    \Tile_X2Y6_WW4BEG[12] ,
    \Tile_X2Y6_WW4BEG[11] ,
    \Tile_X2Y6_WW4BEG[10] ,
    \Tile_X2Y6_WW4BEG[9] ,
    \Tile_X2Y6_WW4BEG[8] ,
    \Tile_X2Y6_WW4BEG[7] ,
    \Tile_X2Y6_WW4BEG[6] ,
    \Tile_X2Y6_WW4BEG[5] ,
    \Tile_X2Y6_WW4BEG[4] ,
    \Tile_X2Y6_WW4BEG[3] ,
    \Tile_X2Y6_WW4BEG[2] ,
    \Tile_X2Y6_WW4BEG[1] ,
    \Tile_X2Y6_WW4BEG[0] }),
    .WW4END({\Tile_X3Y6_WW4BEG[15] ,
    \Tile_X3Y6_WW4BEG[14] ,
    \Tile_X3Y6_WW4BEG[13] ,
    \Tile_X3Y6_WW4BEG[12] ,
    \Tile_X3Y6_WW4BEG[11] ,
    \Tile_X3Y6_WW4BEG[10] ,
    \Tile_X3Y6_WW4BEG[9] ,
    \Tile_X3Y6_WW4BEG[8] ,
    \Tile_X3Y6_WW4BEG[7] ,
    \Tile_X3Y6_WW4BEG[6] ,
    \Tile_X3Y6_WW4BEG[5] ,
    \Tile_X3Y6_WW4BEG[4] ,
    \Tile_X3Y6_WW4BEG[3] ,
    \Tile_X3Y6_WW4BEG[2] ,
    \Tile_X3Y6_WW4BEG[1] ,
    \Tile_X3Y6_WW4BEG[0] }));
 LUT4AB Tile_X2Y7_LUT4AB (.Ci(Tile_X2Y8_Co),
    .Co(Tile_X2Y7_Co),
    .UserCLK(Tile_X2Y8_UserCLKo),
    .UserCLKo(Tile_X2Y7_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X2Y7_E1BEG[3] ,
    \Tile_X2Y7_E1BEG[2] ,
    \Tile_X2Y7_E1BEG[1] ,
    \Tile_X2Y7_E1BEG[0] }),
    .E1END({\Tile_X1Y7_E1BEG[3] ,
    \Tile_X1Y7_E1BEG[2] ,
    \Tile_X1Y7_E1BEG[1] ,
    \Tile_X1Y7_E1BEG[0] }),
    .E2BEG({\Tile_X2Y7_E2BEG[7] ,
    \Tile_X2Y7_E2BEG[6] ,
    \Tile_X2Y7_E2BEG[5] ,
    \Tile_X2Y7_E2BEG[4] ,
    \Tile_X2Y7_E2BEG[3] ,
    \Tile_X2Y7_E2BEG[2] ,
    \Tile_X2Y7_E2BEG[1] ,
    \Tile_X2Y7_E2BEG[0] }),
    .E2BEGb({\Tile_X2Y7_E2BEGb[7] ,
    \Tile_X2Y7_E2BEGb[6] ,
    \Tile_X2Y7_E2BEGb[5] ,
    \Tile_X2Y7_E2BEGb[4] ,
    \Tile_X2Y7_E2BEGb[3] ,
    \Tile_X2Y7_E2BEGb[2] ,
    \Tile_X2Y7_E2BEGb[1] ,
    \Tile_X2Y7_E2BEGb[0] }),
    .E2END({\Tile_X1Y7_E2BEGb[7] ,
    \Tile_X1Y7_E2BEGb[6] ,
    \Tile_X1Y7_E2BEGb[5] ,
    \Tile_X1Y7_E2BEGb[4] ,
    \Tile_X1Y7_E2BEGb[3] ,
    \Tile_X1Y7_E2BEGb[2] ,
    \Tile_X1Y7_E2BEGb[1] ,
    \Tile_X1Y7_E2BEGb[0] }),
    .E2MID({\Tile_X1Y7_E2BEG[7] ,
    \Tile_X1Y7_E2BEG[6] ,
    \Tile_X1Y7_E2BEG[5] ,
    \Tile_X1Y7_E2BEG[4] ,
    \Tile_X1Y7_E2BEG[3] ,
    \Tile_X1Y7_E2BEG[2] ,
    \Tile_X1Y7_E2BEG[1] ,
    \Tile_X1Y7_E2BEG[0] }),
    .E6BEG({\Tile_X2Y7_E6BEG[11] ,
    \Tile_X2Y7_E6BEG[10] ,
    \Tile_X2Y7_E6BEG[9] ,
    \Tile_X2Y7_E6BEG[8] ,
    \Tile_X2Y7_E6BEG[7] ,
    \Tile_X2Y7_E6BEG[6] ,
    \Tile_X2Y7_E6BEG[5] ,
    \Tile_X2Y7_E6BEG[4] ,
    \Tile_X2Y7_E6BEG[3] ,
    \Tile_X2Y7_E6BEG[2] ,
    \Tile_X2Y7_E6BEG[1] ,
    \Tile_X2Y7_E6BEG[0] }),
    .E6END({\Tile_X1Y7_E6BEG[11] ,
    \Tile_X1Y7_E6BEG[10] ,
    \Tile_X1Y7_E6BEG[9] ,
    \Tile_X1Y7_E6BEG[8] ,
    \Tile_X1Y7_E6BEG[7] ,
    \Tile_X1Y7_E6BEG[6] ,
    \Tile_X1Y7_E6BEG[5] ,
    \Tile_X1Y7_E6BEG[4] ,
    \Tile_X1Y7_E6BEG[3] ,
    \Tile_X1Y7_E6BEG[2] ,
    \Tile_X1Y7_E6BEG[1] ,
    \Tile_X1Y7_E6BEG[0] }),
    .EE4BEG({\Tile_X2Y7_EE4BEG[15] ,
    \Tile_X2Y7_EE4BEG[14] ,
    \Tile_X2Y7_EE4BEG[13] ,
    \Tile_X2Y7_EE4BEG[12] ,
    \Tile_X2Y7_EE4BEG[11] ,
    \Tile_X2Y7_EE4BEG[10] ,
    \Tile_X2Y7_EE4BEG[9] ,
    \Tile_X2Y7_EE4BEG[8] ,
    \Tile_X2Y7_EE4BEG[7] ,
    \Tile_X2Y7_EE4BEG[6] ,
    \Tile_X2Y7_EE4BEG[5] ,
    \Tile_X2Y7_EE4BEG[4] ,
    \Tile_X2Y7_EE4BEG[3] ,
    \Tile_X2Y7_EE4BEG[2] ,
    \Tile_X2Y7_EE4BEG[1] ,
    \Tile_X2Y7_EE4BEG[0] }),
    .EE4END({\Tile_X1Y7_EE4BEG[15] ,
    \Tile_X1Y7_EE4BEG[14] ,
    \Tile_X1Y7_EE4BEG[13] ,
    \Tile_X1Y7_EE4BEG[12] ,
    \Tile_X1Y7_EE4BEG[11] ,
    \Tile_X1Y7_EE4BEG[10] ,
    \Tile_X1Y7_EE4BEG[9] ,
    \Tile_X1Y7_EE4BEG[8] ,
    \Tile_X1Y7_EE4BEG[7] ,
    \Tile_X1Y7_EE4BEG[6] ,
    \Tile_X1Y7_EE4BEG[5] ,
    \Tile_X1Y7_EE4BEG[4] ,
    \Tile_X1Y7_EE4BEG[3] ,
    \Tile_X1Y7_EE4BEG[2] ,
    \Tile_X1Y7_EE4BEG[1] ,
    \Tile_X1Y7_EE4BEG[0] }),
    .FrameData({\Tile_X1Y7_FrameData_O[31] ,
    \Tile_X1Y7_FrameData_O[30] ,
    \Tile_X1Y7_FrameData_O[29] ,
    \Tile_X1Y7_FrameData_O[28] ,
    \Tile_X1Y7_FrameData_O[27] ,
    \Tile_X1Y7_FrameData_O[26] ,
    \Tile_X1Y7_FrameData_O[25] ,
    \Tile_X1Y7_FrameData_O[24] ,
    \Tile_X1Y7_FrameData_O[23] ,
    \Tile_X1Y7_FrameData_O[22] ,
    \Tile_X1Y7_FrameData_O[21] ,
    \Tile_X1Y7_FrameData_O[20] ,
    \Tile_X1Y7_FrameData_O[19] ,
    \Tile_X1Y7_FrameData_O[18] ,
    \Tile_X1Y7_FrameData_O[17] ,
    \Tile_X1Y7_FrameData_O[16] ,
    \Tile_X1Y7_FrameData_O[15] ,
    \Tile_X1Y7_FrameData_O[14] ,
    \Tile_X1Y7_FrameData_O[13] ,
    \Tile_X1Y7_FrameData_O[12] ,
    \Tile_X1Y7_FrameData_O[11] ,
    \Tile_X1Y7_FrameData_O[10] ,
    \Tile_X1Y7_FrameData_O[9] ,
    \Tile_X1Y7_FrameData_O[8] ,
    \Tile_X1Y7_FrameData_O[7] ,
    \Tile_X1Y7_FrameData_O[6] ,
    \Tile_X1Y7_FrameData_O[5] ,
    \Tile_X1Y7_FrameData_O[4] ,
    \Tile_X1Y7_FrameData_O[3] ,
    \Tile_X1Y7_FrameData_O[2] ,
    \Tile_X1Y7_FrameData_O[1] ,
    \Tile_X1Y7_FrameData_O[0] }),
    .FrameData_O({\Tile_X2Y7_FrameData_O[31] ,
    \Tile_X2Y7_FrameData_O[30] ,
    \Tile_X2Y7_FrameData_O[29] ,
    \Tile_X2Y7_FrameData_O[28] ,
    \Tile_X2Y7_FrameData_O[27] ,
    \Tile_X2Y7_FrameData_O[26] ,
    \Tile_X2Y7_FrameData_O[25] ,
    \Tile_X2Y7_FrameData_O[24] ,
    \Tile_X2Y7_FrameData_O[23] ,
    \Tile_X2Y7_FrameData_O[22] ,
    \Tile_X2Y7_FrameData_O[21] ,
    \Tile_X2Y7_FrameData_O[20] ,
    \Tile_X2Y7_FrameData_O[19] ,
    \Tile_X2Y7_FrameData_O[18] ,
    \Tile_X2Y7_FrameData_O[17] ,
    \Tile_X2Y7_FrameData_O[16] ,
    \Tile_X2Y7_FrameData_O[15] ,
    \Tile_X2Y7_FrameData_O[14] ,
    \Tile_X2Y7_FrameData_O[13] ,
    \Tile_X2Y7_FrameData_O[12] ,
    \Tile_X2Y7_FrameData_O[11] ,
    \Tile_X2Y7_FrameData_O[10] ,
    \Tile_X2Y7_FrameData_O[9] ,
    \Tile_X2Y7_FrameData_O[8] ,
    \Tile_X2Y7_FrameData_O[7] ,
    \Tile_X2Y7_FrameData_O[6] ,
    \Tile_X2Y7_FrameData_O[5] ,
    \Tile_X2Y7_FrameData_O[4] ,
    \Tile_X2Y7_FrameData_O[3] ,
    \Tile_X2Y7_FrameData_O[2] ,
    \Tile_X2Y7_FrameData_O[1] ,
    \Tile_X2Y7_FrameData_O[0] }),
    .FrameStrobe({\Tile_X2Y8_FrameStrobe_O[19] ,
    \Tile_X2Y8_FrameStrobe_O[18] ,
    \Tile_X2Y8_FrameStrobe_O[17] ,
    \Tile_X2Y8_FrameStrobe_O[16] ,
    \Tile_X2Y8_FrameStrobe_O[15] ,
    \Tile_X2Y8_FrameStrobe_O[14] ,
    \Tile_X2Y8_FrameStrobe_O[13] ,
    \Tile_X2Y8_FrameStrobe_O[12] ,
    \Tile_X2Y8_FrameStrobe_O[11] ,
    \Tile_X2Y8_FrameStrobe_O[10] ,
    \Tile_X2Y8_FrameStrobe_O[9] ,
    \Tile_X2Y8_FrameStrobe_O[8] ,
    \Tile_X2Y8_FrameStrobe_O[7] ,
    \Tile_X2Y8_FrameStrobe_O[6] ,
    \Tile_X2Y8_FrameStrobe_O[5] ,
    \Tile_X2Y8_FrameStrobe_O[4] ,
    \Tile_X2Y8_FrameStrobe_O[3] ,
    \Tile_X2Y8_FrameStrobe_O[2] ,
    \Tile_X2Y8_FrameStrobe_O[1] ,
    \Tile_X2Y8_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X2Y7_FrameStrobe_O[19] ,
    \Tile_X2Y7_FrameStrobe_O[18] ,
    \Tile_X2Y7_FrameStrobe_O[17] ,
    \Tile_X2Y7_FrameStrobe_O[16] ,
    \Tile_X2Y7_FrameStrobe_O[15] ,
    \Tile_X2Y7_FrameStrobe_O[14] ,
    \Tile_X2Y7_FrameStrobe_O[13] ,
    \Tile_X2Y7_FrameStrobe_O[12] ,
    \Tile_X2Y7_FrameStrobe_O[11] ,
    \Tile_X2Y7_FrameStrobe_O[10] ,
    \Tile_X2Y7_FrameStrobe_O[9] ,
    \Tile_X2Y7_FrameStrobe_O[8] ,
    \Tile_X2Y7_FrameStrobe_O[7] ,
    \Tile_X2Y7_FrameStrobe_O[6] ,
    \Tile_X2Y7_FrameStrobe_O[5] ,
    \Tile_X2Y7_FrameStrobe_O[4] ,
    \Tile_X2Y7_FrameStrobe_O[3] ,
    \Tile_X2Y7_FrameStrobe_O[2] ,
    \Tile_X2Y7_FrameStrobe_O[1] ,
    \Tile_X2Y7_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X2Y7_N1BEG[3] ,
    \Tile_X2Y7_N1BEG[2] ,
    \Tile_X2Y7_N1BEG[1] ,
    \Tile_X2Y7_N1BEG[0] }),
    .N1END({\Tile_X2Y8_N1BEG[3] ,
    \Tile_X2Y8_N1BEG[2] ,
    \Tile_X2Y8_N1BEG[1] ,
    \Tile_X2Y8_N1BEG[0] }),
    .N2BEG({\Tile_X2Y7_N2BEG[7] ,
    \Tile_X2Y7_N2BEG[6] ,
    \Tile_X2Y7_N2BEG[5] ,
    \Tile_X2Y7_N2BEG[4] ,
    \Tile_X2Y7_N2BEG[3] ,
    \Tile_X2Y7_N2BEG[2] ,
    \Tile_X2Y7_N2BEG[1] ,
    \Tile_X2Y7_N2BEG[0] }),
    .N2BEGb({\Tile_X2Y7_N2BEGb[7] ,
    \Tile_X2Y7_N2BEGb[6] ,
    \Tile_X2Y7_N2BEGb[5] ,
    \Tile_X2Y7_N2BEGb[4] ,
    \Tile_X2Y7_N2BEGb[3] ,
    \Tile_X2Y7_N2BEGb[2] ,
    \Tile_X2Y7_N2BEGb[1] ,
    \Tile_X2Y7_N2BEGb[0] }),
    .N2END({\Tile_X2Y8_N2BEGb[7] ,
    \Tile_X2Y8_N2BEGb[6] ,
    \Tile_X2Y8_N2BEGb[5] ,
    \Tile_X2Y8_N2BEGb[4] ,
    \Tile_X2Y8_N2BEGb[3] ,
    \Tile_X2Y8_N2BEGb[2] ,
    \Tile_X2Y8_N2BEGb[1] ,
    \Tile_X2Y8_N2BEGb[0] }),
    .N2MID({\Tile_X2Y8_N2BEG[7] ,
    \Tile_X2Y8_N2BEG[6] ,
    \Tile_X2Y8_N2BEG[5] ,
    \Tile_X2Y8_N2BEG[4] ,
    \Tile_X2Y8_N2BEG[3] ,
    \Tile_X2Y8_N2BEG[2] ,
    \Tile_X2Y8_N2BEG[1] ,
    \Tile_X2Y8_N2BEG[0] }),
    .N4BEG({\Tile_X2Y7_N4BEG[15] ,
    \Tile_X2Y7_N4BEG[14] ,
    \Tile_X2Y7_N4BEG[13] ,
    \Tile_X2Y7_N4BEG[12] ,
    \Tile_X2Y7_N4BEG[11] ,
    \Tile_X2Y7_N4BEG[10] ,
    \Tile_X2Y7_N4BEG[9] ,
    \Tile_X2Y7_N4BEG[8] ,
    \Tile_X2Y7_N4BEG[7] ,
    \Tile_X2Y7_N4BEG[6] ,
    \Tile_X2Y7_N4BEG[5] ,
    \Tile_X2Y7_N4BEG[4] ,
    \Tile_X2Y7_N4BEG[3] ,
    \Tile_X2Y7_N4BEG[2] ,
    \Tile_X2Y7_N4BEG[1] ,
    \Tile_X2Y7_N4BEG[0] }),
    .N4END({\Tile_X2Y8_N4BEG[15] ,
    \Tile_X2Y8_N4BEG[14] ,
    \Tile_X2Y8_N4BEG[13] ,
    \Tile_X2Y8_N4BEG[12] ,
    \Tile_X2Y8_N4BEG[11] ,
    \Tile_X2Y8_N4BEG[10] ,
    \Tile_X2Y8_N4BEG[9] ,
    \Tile_X2Y8_N4BEG[8] ,
    \Tile_X2Y8_N4BEG[7] ,
    \Tile_X2Y8_N4BEG[6] ,
    \Tile_X2Y8_N4BEG[5] ,
    \Tile_X2Y8_N4BEG[4] ,
    \Tile_X2Y8_N4BEG[3] ,
    \Tile_X2Y8_N4BEG[2] ,
    \Tile_X2Y8_N4BEG[1] ,
    \Tile_X2Y8_N4BEG[0] }),
    .NN4BEG({\Tile_X2Y7_NN4BEG[15] ,
    \Tile_X2Y7_NN4BEG[14] ,
    \Tile_X2Y7_NN4BEG[13] ,
    \Tile_X2Y7_NN4BEG[12] ,
    \Tile_X2Y7_NN4BEG[11] ,
    \Tile_X2Y7_NN4BEG[10] ,
    \Tile_X2Y7_NN4BEG[9] ,
    \Tile_X2Y7_NN4BEG[8] ,
    \Tile_X2Y7_NN4BEG[7] ,
    \Tile_X2Y7_NN4BEG[6] ,
    \Tile_X2Y7_NN4BEG[5] ,
    \Tile_X2Y7_NN4BEG[4] ,
    \Tile_X2Y7_NN4BEG[3] ,
    \Tile_X2Y7_NN4BEG[2] ,
    \Tile_X2Y7_NN4BEG[1] ,
    \Tile_X2Y7_NN4BEG[0] }),
    .NN4END({\Tile_X2Y8_NN4BEG[15] ,
    \Tile_X2Y8_NN4BEG[14] ,
    \Tile_X2Y8_NN4BEG[13] ,
    \Tile_X2Y8_NN4BEG[12] ,
    \Tile_X2Y8_NN4BEG[11] ,
    \Tile_X2Y8_NN4BEG[10] ,
    \Tile_X2Y8_NN4BEG[9] ,
    \Tile_X2Y8_NN4BEG[8] ,
    \Tile_X2Y8_NN4BEG[7] ,
    \Tile_X2Y8_NN4BEG[6] ,
    \Tile_X2Y8_NN4BEG[5] ,
    \Tile_X2Y8_NN4BEG[4] ,
    \Tile_X2Y8_NN4BEG[3] ,
    \Tile_X2Y8_NN4BEG[2] ,
    \Tile_X2Y8_NN4BEG[1] ,
    \Tile_X2Y8_NN4BEG[0] }),
    .S1BEG({\Tile_X2Y7_S1BEG[3] ,
    \Tile_X2Y7_S1BEG[2] ,
    \Tile_X2Y7_S1BEG[1] ,
    \Tile_X2Y7_S1BEG[0] }),
    .S1END({\Tile_X2Y6_S1BEG[3] ,
    \Tile_X2Y6_S1BEG[2] ,
    \Tile_X2Y6_S1BEG[1] ,
    \Tile_X2Y6_S1BEG[0] }),
    .S2BEG({\Tile_X2Y7_S2BEG[7] ,
    \Tile_X2Y7_S2BEG[6] ,
    \Tile_X2Y7_S2BEG[5] ,
    \Tile_X2Y7_S2BEG[4] ,
    \Tile_X2Y7_S2BEG[3] ,
    \Tile_X2Y7_S2BEG[2] ,
    \Tile_X2Y7_S2BEG[1] ,
    \Tile_X2Y7_S2BEG[0] }),
    .S2BEGb({\Tile_X2Y7_S2BEGb[7] ,
    \Tile_X2Y7_S2BEGb[6] ,
    \Tile_X2Y7_S2BEGb[5] ,
    \Tile_X2Y7_S2BEGb[4] ,
    \Tile_X2Y7_S2BEGb[3] ,
    \Tile_X2Y7_S2BEGb[2] ,
    \Tile_X2Y7_S2BEGb[1] ,
    \Tile_X2Y7_S2BEGb[0] }),
    .S2END({\Tile_X2Y6_S2BEGb[7] ,
    \Tile_X2Y6_S2BEGb[6] ,
    \Tile_X2Y6_S2BEGb[5] ,
    \Tile_X2Y6_S2BEGb[4] ,
    \Tile_X2Y6_S2BEGb[3] ,
    \Tile_X2Y6_S2BEGb[2] ,
    \Tile_X2Y6_S2BEGb[1] ,
    \Tile_X2Y6_S2BEGb[0] }),
    .S2MID({\Tile_X2Y6_S2BEG[7] ,
    \Tile_X2Y6_S2BEG[6] ,
    \Tile_X2Y6_S2BEG[5] ,
    \Tile_X2Y6_S2BEG[4] ,
    \Tile_X2Y6_S2BEG[3] ,
    \Tile_X2Y6_S2BEG[2] ,
    \Tile_X2Y6_S2BEG[1] ,
    \Tile_X2Y6_S2BEG[0] }),
    .S4BEG({\Tile_X2Y7_S4BEG[15] ,
    \Tile_X2Y7_S4BEG[14] ,
    \Tile_X2Y7_S4BEG[13] ,
    \Tile_X2Y7_S4BEG[12] ,
    \Tile_X2Y7_S4BEG[11] ,
    \Tile_X2Y7_S4BEG[10] ,
    \Tile_X2Y7_S4BEG[9] ,
    \Tile_X2Y7_S4BEG[8] ,
    \Tile_X2Y7_S4BEG[7] ,
    \Tile_X2Y7_S4BEG[6] ,
    \Tile_X2Y7_S4BEG[5] ,
    \Tile_X2Y7_S4BEG[4] ,
    \Tile_X2Y7_S4BEG[3] ,
    \Tile_X2Y7_S4BEG[2] ,
    \Tile_X2Y7_S4BEG[1] ,
    \Tile_X2Y7_S4BEG[0] }),
    .S4END({\Tile_X2Y6_S4BEG[15] ,
    \Tile_X2Y6_S4BEG[14] ,
    \Tile_X2Y6_S4BEG[13] ,
    \Tile_X2Y6_S4BEG[12] ,
    \Tile_X2Y6_S4BEG[11] ,
    \Tile_X2Y6_S4BEG[10] ,
    \Tile_X2Y6_S4BEG[9] ,
    \Tile_X2Y6_S4BEG[8] ,
    \Tile_X2Y6_S4BEG[7] ,
    \Tile_X2Y6_S4BEG[6] ,
    \Tile_X2Y6_S4BEG[5] ,
    \Tile_X2Y6_S4BEG[4] ,
    \Tile_X2Y6_S4BEG[3] ,
    \Tile_X2Y6_S4BEG[2] ,
    \Tile_X2Y6_S4BEG[1] ,
    \Tile_X2Y6_S4BEG[0] }),
    .SS4BEG({\Tile_X2Y7_SS4BEG[15] ,
    \Tile_X2Y7_SS4BEG[14] ,
    \Tile_X2Y7_SS4BEG[13] ,
    \Tile_X2Y7_SS4BEG[12] ,
    \Tile_X2Y7_SS4BEG[11] ,
    \Tile_X2Y7_SS4BEG[10] ,
    \Tile_X2Y7_SS4BEG[9] ,
    \Tile_X2Y7_SS4BEG[8] ,
    \Tile_X2Y7_SS4BEG[7] ,
    \Tile_X2Y7_SS4BEG[6] ,
    \Tile_X2Y7_SS4BEG[5] ,
    \Tile_X2Y7_SS4BEG[4] ,
    \Tile_X2Y7_SS4BEG[3] ,
    \Tile_X2Y7_SS4BEG[2] ,
    \Tile_X2Y7_SS4BEG[1] ,
    \Tile_X2Y7_SS4BEG[0] }),
    .SS4END({\Tile_X2Y6_SS4BEG[15] ,
    \Tile_X2Y6_SS4BEG[14] ,
    \Tile_X2Y6_SS4BEG[13] ,
    \Tile_X2Y6_SS4BEG[12] ,
    \Tile_X2Y6_SS4BEG[11] ,
    \Tile_X2Y6_SS4BEG[10] ,
    \Tile_X2Y6_SS4BEG[9] ,
    \Tile_X2Y6_SS4BEG[8] ,
    \Tile_X2Y6_SS4BEG[7] ,
    \Tile_X2Y6_SS4BEG[6] ,
    \Tile_X2Y6_SS4BEG[5] ,
    \Tile_X2Y6_SS4BEG[4] ,
    \Tile_X2Y6_SS4BEG[3] ,
    \Tile_X2Y6_SS4BEG[2] ,
    \Tile_X2Y6_SS4BEG[1] ,
    \Tile_X2Y6_SS4BEG[0] }),
    .W1BEG({\Tile_X2Y7_W1BEG[3] ,
    \Tile_X2Y7_W1BEG[2] ,
    \Tile_X2Y7_W1BEG[1] ,
    \Tile_X2Y7_W1BEG[0] }),
    .W1END({\Tile_X3Y7_W1BEG[3] ,
    \Tile_X3Y7_W1BEG[2] ,
    \Tile_X3Y7_W1BEG[1] ,
    \Tile_X3Y7_W1BEG[0] }),
    .W2BEG({\Tile_X2Y7_W2BEG[7] ,
    \Tile_X2Y7_W2BEG[6] ,
    \Tile_X2Y7_W2BEG[5] ,
    \Tile_X2Y7_W2BEG[4] ,
    \Tile_X2Y7_W2BEG[3] ,
    \Tile_X2Y7_W2BEG[2] ,
    \Tile_X2Y7_W2BEG[1] ,
    \Tile_X2Y7_W2BEG[0] }),
    .W2BEGb({\Tile_X2Y7_W2BEGb[7] ,
    \Tile_X2Y7_W2BEGb[6] ,
    \Tile_X2Y7_W2BEGb[5] ,
    \Tile_X2Y7_W2BEGb[4] ,
    \Tile_X2Y7_W2BEGb[3] ,
    \Tile_X2Y7_W2BEGb[2] ,
    \Tile_X2Y7_W2BEGb[1] ,
    \Tile_X2Y7_W2BEGb[0] }),
    .W2END({\Tile_X3Y7_W2BEGb[7] ,
    \Tile_X3Y7_W2BEGb[6] ,
    \Tile_X3Y7_W2BEGb[5] ,
    \Tile_X3Y7_W2BEGb[4] ,
    \Tile_X3Y7_W2BEGb[3] ,
    \Tile_X3Y7_W2BEGb[2] ,
    \Tile_X3Y7_W2BEGb[1] ,
    \Tile_X3Y7_W2BEGb[0] }),
    .W2MID({\Tile_X3Y7_W2BEG[7] ,
    \Tile_X3Y7_W2BEG[6] ,
    \Tile_X3Y7_W2BEG[5] ,
    \Tile_X3Y7_W2BEG[4] ,
    \Tile_X3Y7_W2BEG[3] ,
    \Tile_X3Y7_W2BEG[2] ,
    \Tile_X3Y7_W2BEG[1] ,
    \Tile_X3Y7_W2BEG[0] }),
    .W6BEG({\Tile_X2Y7_W6BEG[11] ,
    \Tile_X2Y7_W6BEG[10] ,
    \Tile_X2Y7_W6BEG[9] ,
    \Tile_X2Y7_W6BEG[8] ,
    \Tile_X2Y7_W6BEG[7] ,
    \Tile_X2Y7_W6BEG[6] ,
    \Tile_X2Y7_W6BEG[5] ,
    \Tile_X2Y7_W6BEG[4] ,
    \Tile_X2Y7_W6BEG[3] ,
    \Tile_X2Y7_W6BEG[2] ,
    \Tile_X2Y7_W6BEG[1] ,
    \Tile_X2Y7_W6BEG[0] }),
    .W6END({\Tile_X3Y7_W6BEG[11] ,
    \Tile_X3Y7_W6BEG[10] ,
    \Tile_X3Y7_W6BEG[9] ,
    \Tile_X3Y7_W6BEG[8] ,
    \Tile_X3Y7_W6BEG[7] ,
    \Tile_X3Y7_W6BEG[6] ,
    \Tile_X3Y7_W6BEG[5] ,
    \Tile_X3Y7_W6BEG[4] ,
    \Tile_X3Y7_W6BEG[3] ,
    \Tile_X3Y7_W6BEG[2] ,
    \Tile_X3Y7_W6BEG[1] ,
    \Tile_X3Y7_W6BEG[0] }),
    .WW4BEG({\Tile_X2Y7_WW4BEG[15] ,
    \Tile_X2Y7_WW4BEG[14] ,
    \Tile_X2Y7_WW4BEG[13] ,
    \Tile_X2Y7_WW4BEG[12] ,
    \Tile_X2Y7_WW4BEG[11] ,
    \Tile_X2Y7_WW4BEG[10] ,
    \Tile_X2Y7_WW4BEG[9] ,
    \Tile_X2Y7_WW4BEG[8] ,
    \Tile_X2Y7_WW4BEG[7] ,
    \Tile_X2Y7_WW4BEG[6] ,
    \Tile_X2Y7_WW4BEG[5] ,
    \Tile_X2Y7_WW4BEG[4] ,
    \Tile_X2Y7_WW4BEG[3] ,
    \Tile_X2Y7_WW4BEG[2] ,
    \Tile_X2Y7_WW4BEG[1] ,
    \Tile_X2Y7_WW4BEG[0] }),
    .WW4END({\Tile_X3Y7_WW4BEG[15] ,
    \Tile_X3Y7_WW4BEG[14] ,
    \Tile_X3Y7_WW4BEG[13] ,
    \Tile_X3Y7_WW4BEG[12] ,
    \Tile_X3Y7_WW4BEG[11] ,
    \Tile_X3Y7_WW4BEG[10] ,
    \Tile_X3Y7_WW4BEG[9] ,
    \Tile_X3Y7_WW4BEG[8] ,
    \Tile_X3Y7_WW4BEG[7] ,
    \Tile_X3Y7_WW4BEG[6] ,
    \Tile_X3Y7_WW4BEG[5] ,
    \Tile_X3Y7_WW4BEG[4] ,
    \Tile_X3Y7_WW4BEG[3] ,
    \Tile_X3Y7_WW4BEG[2] ,
    \Tile_X3Y7_WW4BEG[1] ,
    \Tile_X3Y7_WW4BEG[0] }));
 LUT4AB Tile_X2Y8_LUT4AB (.Ci(Tile_X2Y9_Co),
    .Co(Tile_X2Y8_Co),
    .UserCLK(Tile_X2Y9_UserCLKo),
    .UserCLKo(Tile_X2Y8_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X2Y8_E1BEG[3] ,
    \Tile_X2Y8_E1BEG[2] ,
    \Tile_X2Y8_E1BEG[1] ,
    \Tile_X2Y8_E1BEG[0] }),
    .E1END({\Tile_X1Y8_E1BEG[3] ,
    \Tile_X1Y8_E1BEG[2] ,
    \Tile_X1Y8_E1BEG[1] ,
    \Tile_X1Y8_E1BEG[0] }),
    .E2BEG({\Tile_X2Y8_E2BEG[7] ,
    \Tile_X2Y8_E2BEG[6] ,
    \Tile_X2Y8_E2BEG[5] ,
    \Tile_X2Y8_E2BEG[4] ,
    \Tile_X2Y8_E2BEG[3] ,
    \Tile_X2Y8_E2BEG[2] ,
    \Tile_X2Y8_E2BEG[1] ,
    \Tile_X2Y8_E2BEG[0] }),
    .E2BEGb({\Tile_X2Y8_E2BEGb[7] ,
    \Tile_X2Y8_E2BEGb[6] ,
    \Tile_X2Y8_E2BEGb[5] ,
    \Tile_X2Y8_E2BEGb[4] ,
    \Tile_X2Y8_E2BEGb[3] ,
    \Tile_X2Y8_E2BEGb[2] ,
    \Tile_X2Y8_E2BEGb[1] ,
    \Tile_X2Y8_E2BEGb[0] }),
    .E2END({\Tile_X1Y8_E2BEGb[7] ,
    \Tile_X1Y8_E2BEGb[6] ,
    \Tile_X1Y8_E2BEGb[5] ,
    \Tile_X1Y8_E2BEGb[4] ,
    \Tile_X1Y8_E2BEGb[3] ,
    \Tile_X1Y8_E2BEGb[2] ,
    \Tile_X1Y8_E2BEGb[1] ,
    \Tile_X1Y8_E2BEGb[0] }),
    .E2MID({\Tile_X1Y8_E2BEG[7] ,
    \Tile_X1Y8_E2BEG[6] ,
    \Tile_X1Y8_E2BEG[5] ,
    \Tile_X1Y8_E2BEG[4] ,
    \Tile_X1Y8_E2BEG[3] ,
    \Tile_X1Y8_E2BEG[2] ,
    \Tile_X1Y8_E2BEG[1] ,
    \Tile_X1Y8_E2BEG[0] }),
    .E6BEG({\Tile_X2Y8_E6BEG[11] ,
    \Tile_X2Y8_E6BEG[10] ,
    \Tile_X2Y8_E6BEG[9] ,
    \Tile_X2Y8_E6BEG[8] ,
    \Tile_X2Y8_E6BEG[7] ,
    \Tile_X2Y8_E6BEG[6] ,
    \Tile_X2Y8_E6BEG[5] ,
    \Tile_X2Y8_E6BEG[4] ,
    \Tile_X2Y8_E6BEG[3] ,
    \Tile_X2Y8_E6BEG[2] ,
    \Tile_X2Y8_E6BEG[1] ,
    \Tile_X2Y8_E6BEG[0] }),
    .E6END({\Tile_X1Y8_E6BEG[11] ,
    \Tile_X1Y8_E6BEG[10] ,
    \Tile_X1Y8_E6BEG[9] ,
    \Tile_X1Y8_E6BEG[8] ,
    \Tile_X1Y8_E6BEG[7] ,
    \Tile_X1Y8_E6BEG[6] ,
    \Tile_X1Y8_E6BEG[5] ,
    \Tile_X1Y8_E6BEG[4] ,
    \Tile_X1Y8_E6BEG[3] ,
    \Tile_X1Y8_E6BEG[2] ,
    \Tile_X1Y8_E6BEG[1] ,
    \Tile_X1Y8_E6BEG[0] }),
    .EE4BEG({\Tile_X2Y8_EE4BEG[15] ,
    \Tile_X2Y8_EE4BEG[14] ,
    \Tile_X2Y8_EE4BEG[13] ,
    \Tile_X2Y8_EE4BEG[12] ,
    \Tile_X2Y8_EE4BEG[11] ,
    \Tile_X2Y8_EE4BEG[10] ,
    \Tile_X2Y8_EE4BEG[9] ,
    \Tile_X2Y8_EE4BEG[8] ,
    \Tile_X2Y8_EE4BEG[7] ,
    \Tile_X2Y8_EE4BEG[6] ,
    \Tile_X2Y8_EE4BEG[5] ,
    \Tile_X2Y8_EE4BEG[4] ,
    \Tile_X2Y8_EE4BEG[3] ,
    \Tile_X2Y8_EE4BEG[2] ,
    \Tile_X2Y8_EE4BEG[1] ,
    \Tile_X2Y8_EE4BEG[0] }),
    .EE4END({\Tile_X1Y8_EE4BEG[15] ,
    \Tile_X1Y8_EE4BEG[14] ,
    \Tile_X1Y8_EE4BEG[13] ,
    \Tile_X1Y8_EE4BEG[12] ,
    \Tile_X1Y8_EE4BEG[11] ,
    \Tile_X1Y8_EE4BEG[10] ,
    \Tile_X1Y8_EE4BEG[9] ,
    \Tile_X1Y8_EE4BEG[8] ,
    \Tile_X1Y8_EE4BEG[7] ,
    \Tile_X1Y8_EE4BEG[6] ,
    \Tile_X1Y8_EE4BEG[5] ,
    \Tile_X1Y8_EE4BEG[4] ,
    \Tile_X1Y8_EE4BEG[3] ,
    \Tile_X1Y8_EE4BEG[2] ,
    \Tile_X1Y8_EE4BEG[1] ,
    \Tile_X1Y8_EE4BEG[0] }),
    .FrameData({\Tile_X1Y8_FrameData_O[31] ,
    \Tile_X1Y8_FrameData_O[30] ,
    \Tile_X1Y8_FrameData_O[29] ,
    \Tile_X1Y8_FrameData_O[28] ,
    \Tile_X1Y8_FrameData_O[27] ,
    \Tile_X1Y8_FrameData_O[26] ,
    \Tile_X1Y8_FrameData_O[25] ,
    \Tile_X1Y8_FrameData_O[24] ,
    \Tile_X1Y8_FrameData_O[23] ,
    \Tile_X1Y8_FrameData_O[22] ,
    \Tile_X1Y8_FrameData_O[21] ,
    \Tile_X1Y8_FrameData_O[20] ,
    \Tile_X1Y8_FrameData_O[19] ,
    \Tile_X1Y8_FrameData_O[18] ,
    \Tile_X1Y8_FrameData_O[17] ,
    \Tile_X1Y8_FrameData_O[16] ,
    \Tile_X1Y8_FrameData_O[15] ,
    \Tile_X1Y8_FrameData_O[14] ,
    \Tile_X1Y8_FrameData_O[13] ,
    \Tile_X1Y8_FrameData_O[12] ,
    \Tile_X1Y8_FrameData_O[11] ,
    \Tile_X1Y8_FrameData_O[10] ,
    \Tile_X1Y8_FrameData_O[9] ,
    \Tile_X1Y8_FrameData_O[8] ,
    \Tile_X1Y8_FrameData_O[7] ,
    \Tile_X1Y8_FrameData_O[6] ,
    \Tile_X1Y8_FrameData_O[5] ,
    \Tile_X1Y8_FrameData_O[4] ,
    \Tile_X1Y8_FrameData_O[3] ,
    \Tile_X1Y8_FrameData_O[2] ,
    \Tile_X1Y8_FrameData_O[1] ,
    \Tile_X1Y8_FrameData_O[0] }),
    .FrameData_O({\Tile_X2Y8_FrameData_O[31] ,
    \Tile_X2Y8_FrameData_O[30] ,
    \Tile_X2Y8_FrameData_O[29] ,
    \Tile_X2Y8_FrameData_O[28] ,
    \Tile_X2Y8_FrameData_O[27] ,
    \Tile_X2Y8_FrameData_O[26] ,
    \Tile_X2Y8_FrameData_O[25] ,
    \Tile_X2Y8_FrameData_O[24] ,
    \Tile_X2Y8_FrameData_O[23] ,
    \Tile_X2Y8_FrameData_O[22] ,
    \Tile_X2Y8_FrameData_O[21] ,
    \Tile_X2Y8_FrameData_O[20] ,
    \Tile_X2Y8_FrameData_O[19] ,
    \Tile_X2Y8_FrameData_O[18] ,
    \Tile_X2Y8_FrameData_O[17] ,
    \Tile_X2Y8_FrameData_O[16] ,
    \Tile_X2Y8_FrameData_O[15] ,
    \Tile_X2Y8_FrameData_O[14] ,
    \Tile_X2Y8_FrameData_O[13] ,
    \Tile_X2Y8_FrameData_O[12] ,
    \Tile_X2Y8_FrameData_O[11] ,
    \Tile_X2Y8_FrameData_O[10] ,
    \Tile_X2Y8_FrameData_O[9] ,
    \Tile_X2Y8_FrameData_O[8] ,
    \Tile_X2Y8_FrameData_O[7] ,
    \Tile_X2Y8_FrameData_O[6] ,
    \Tile_X2Y8_FrameData_O[5] ,
    \Tile_X2Y8_FrameData_O[4] ,
    \Tile_X2Y8_FrameData_O[3] ,
    \Tile_X2Y8_FrameData_O[2] ,
    \Tile_X2Y8_FrameData_O[1] ,
    \Tile_X2Y8_FrameData_O[0] }),
    .FrameStrobe({\Tile_X2Y9_FrameStrobe_O[19] ,
    \Tile_X2Y9_FrameStrobe_O[18] ,
    \Tile_X2Y9_FrameStrobe_O[17] ,
    \Tile_X2Y9_FrameStrobe_O[16] ,
    \Tile_X2Y9_FrameStrobe_O[15] ,
    \Tile_X2Y9_FrameStrobe_O[14] ,
    \Tile_X2Y9_FrameStrobe_O[13] ,
    \Tile_X2Y9_FrameStrobe_O[12] ,
    \Tile_X2Y9_FrameStrobe_O[11] ,
    \Tile_X2Y9_FrameStrobe_O[10] ,
    \Tile_X2Y9_FrameStrobe_O[9] ,
    \Tile_X2Y9_FrameStrobe_O[8] ,
    \Tile_X2Y9_FrameStrobe_O[7] ,
    \Tile_X2Y9_FrameStrobe_O[6] ,
    \Tile_X2Y9_FrameStrobe_O[5] ,
    \Tile_X2Y9_FrameStrobe_O[4] ,
    \Tile_X2Y9_FrameStrobe_O[3] ,
    \Tile_X2Y9_FrameStrobe_O[2] ,
    \Tile_X2Y9_FrameStrobe_O[1] ,
    \Tile_X2Y9_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X2Y8_FrameStrobe_O[19] ,
    \Tile_X2Y8_FrameStrobe_O[18] ,
    \Tile_X2Y8_FrameStrobe_O[17] ,
    \Tile_X2Y8_FrameStrobe_O[16] ,
    \Tile_X2Y8_FrameStrobe_O[15] ,
    \Tile_X2Y8_FrameStrobe_O[14] ,
    \Tile_X2Y8_FrameStrobe_O[13] ,
    \Tile_X2Y8_FrameStrobe_O[12] ,
    \Tile_X2Y8_FrameStrobe_O[11] ,
    \Tile_X2Y8_FrameStrobe_O[10] ,
    \Tile_X2Y8_FrameStrobe_O[9] ,
    \Tile_X2Y8_FrameStrobe_O[8] ,
    \Tile_X2Y8_FrameStrobe_O[7] ,
    \Tile_X2Y8_FrameStrobe_O[6] ,
    \Tile_X2Y8_FrameStrobe_O[5] ,
    \Tile_X2Y8_FrameStrobe_O[4] ,
    \Tile_X2Y8_FrameStrobe_O[3] ,
    \Tile_X2Y8_FrameStrobe_O[2] ,
    \Tile_X2Y8_FrameStrobe_O[1] ,
    \Tile_X2Y8_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X2Y8_N1BEG[3] ,
    \Tile_X2Y8_N1BEG[2] ,
    \Tile_X2Y8_N1BEG[1] ,
    \Tile_X2Y8_N1BEG[0] }),
    .N1END({\Tile_X2Y9_N1BEG[3] ,
    \Tile_X2Y9_N1BEG[2] ,
    \Tile_X2Y9_N1BEG[1] ,
    \Tile_X2Y9_N1BEG[0] }),
    .N2BEG({\Tile_X2Y8_N2BEG[7] ,
    \Tile_X2Y8_N2BEG[6] ,
    \Tile_X2Y8_N2BEG[5] ,
    \Tile_X2Y8_N2BEG[4] ,
    \Tile_X2Y8_N2BEG[3] ,
    \Tile_X2Y8_N2BEG[2] ,
    \Tile_X2Y8_N2BEG[1] ,
    \Tile_X2Y8_N2BEG[0] }),
    .N2BEGb({\Tile_X2Y8_N2BEGb[7] ,
    \Tile_X2Y8_N2BEGb[6] ,
    \Tile_X2Y8_N2BEGb[5] ,
    \Tile_X2Y8_N2BEGb[4] ,
    \Tile_X2Y8_N2BEGb[3] ,
    \Tile_X2Y8_N2BEGb[2] ,
    \Tile_X2Y8_N2BEGb[1] ,
    \Tile_X2Y8_N2BEGb[0] }),
    .N2END({\Tile_X2Y9_N2BEGb[7] ,
    \Tile_X2Y9_N2BEGb[6] ,
    \Tile_X2Y9_N2BEGb[5] ,
    \Tile_X2Y9_N2BEGb[4] ,
    \Tile_X2Y9_N2BEGb[3] ,
    \Tile_X2Y9_N2BEGb[2] ,
    \Tile_X2Y9_N2BEGb[1] ,
    \Tile_X2Y9_N2BEGb[0] }),
    .N2MID({\Tile_X2Y9_N2BEG[7] ,
    \Tile_X2Y9_N2BEG[6] ,
    \Tile_X2Y9_N2BEG[5] ,
    \Tile_X2Y9_N2BEG[4] ,
    \Tile_X2Y9_N2BEG[3] ,
    \Tile_X2Y9_N2BEG[2] ,
    \Tile_X2Y9_N2BEG[1] ,
    \Tile_X2Y9_N2BEG[0] }),
    .N4BEG({\Tile_X2Y8_N4BEG[15] ,
    \Tile_X2Y8_N4BEG[14] ,
    \Tile_X2Y8_N4BEG[13] ,
    \Tile_X2Y8_N4BEG[12] ,
    \Tile_X2Y8_N4BEG[11] ,
    \Tile_X2Y8_N4BEG[10] ,
    \Tile_X2Y8_N4BEG[9] ,
    \Tile_X2Y8_N4BEG[8] ,
    \Tile_X2Y8_N4BEG[7] ,
    \Tile_X2Y8_N4BEG[6] ,
    \Tile_X2Y8_N4BEG[5] ,
    \Tile_X2Y8_N4BEG[4] ,
    \Tile_X2Y8_N4BEG[3] ,
    \Tile_X2Y8_N4BEG[2] ,
    \Tile_X2Y8_N4BEG[1] ,
    \Tile_X2Y8_N4BEG[0] }),
    .N4END({\Tile_X2Y9_N4BEG[15] ,
    \Tile_X2Y9_N4BEG[14] ,
    \Tile_X2Y9_N4BEG[13] ,
    \Tile_X2Y9_N4BEG[12] ,
    \Tile_X2Y9_N4BEG[11] ,
    \Tile_X2Y9_N4BEG[10] ,
    \Tile_X2Y9_N4BEG[9] ,
    \Tile_X2Y9_N4BEG[8] ,
    \Tile_X2Y9_N4BEG[7] ,
    \Tile_X2Y9_N4BEG[6] ,
    \Tile_X2Y9_N4BEG[5] ,
    \Tile_X2Y9_N4BEG[4] ,
    \Tile_X2Y9_N4BEG[3] ,
    \Tile_X2Y9_N4BEG[2] ,
    \Tile_X2Y9_N4BEG[1] ,
    \Tile_X2Y9_N4BEG[0] }),
    .NN4BEG({\Tile_X2Y8_NN4BEG[15] ,
    \Tile_X2Y8_NN4BEG[14] ,
    \Tile_X2Y8_NN4BEG[13] ,
    \Tile_X2Y8_NN4BEG[12] ,
    \Tile_X2Y8_NN4BEG[11] ,
    \Tile_X2Y8_NN4BEG[10] ,
    \Tile_X2Y8_NN4BEG[9] ,
    \Tile_X2Y8_NN4BEG[8] ,
    \Tile_X2Y8_NN4BEG[7] ,
    \Tile_X2Y8_NN4BEG[6] ,
    \Tile_X2Y8_NN4BEG[5] ,
    \Tile_X2Y8_NN4BEG[4] ,
    \Tile_X2Y8_NN4BEG[3] ,
    \Tile_X2Y8_NN4BEG[2] ,
    \Tile_X2Y8_NN4BEG[1] ,
    \Tile_X2Y8_NN4BEG[0] }),
    .NN4END({\Tile_X2Y9_NN4BEG[15] ,
    \Tile_X2Y9_NN4BEG[14] ,
    \Tile_X2Y9_NN4BEG[13] ,
    \Tile_X2Y9_NN4BEG[12] ,
    \Tile_X2Y9_NN4BEG[11] ,
    \Tile_X2Y9_NN4BEG[10] ,
    \Tile_X2Y9_NN4BEG[9] ,
    \Tile_X2Y9_NN4BEG[8] ,
    \Tile_X2Y9_NN4BEG[7] ,
    \Tile_X2Y9_NN4BEG[6] ,
    \Tile_X2Y9_NN4BEG[5] ,
    \Tile_X2Y9_NN4BEG[4] ,
    \Tile_X2Y9_NN4BEG[3] ,
    \Tile_X2Y9_NN4BEG[2] ,
    \Tile_X2Y9_NN4BEG[1] ,
    \Tile_X2Y9_NN4BEG[0] }),
    .S1BEG({\Tile_X2Y8_S1BEG[3] ,
    \Tile_X2Y8_S1BEG[2] ,
    \Tile_X2Y8_S1BEG[1] ,
    \Tile_X2Y8_S1BEG[0] }),
    .S1END({\Tile_X2Y7_S1BEG[3] ,
    \Tile_X2Y7_S1BEG[2] ,
    \Tile_X2Y7_S1BEG[1] ,
    \Tile_X2Y7_S1BEG[0] }),
    .S2BEG({\Tile_X2Y8_S2BEG[7] ,
    \Tile_X2Y8_S2BEG[6] ,
    \Tile_X2Y8_S2BEG[5] ,
    \Tile_X2Y8_S2BEG[4] ,
    \Tile_X2Y8_S2BEG[3] ,
    \Tile_X2Y8_S2BEG[2] ,
    \Tile_X2Y8_S2BEG[1] ,
    \Tile_X2Y8_S2BEG[0] }),
    .S2BEGb({\Tile_X2Y8_S2BEGb[7] ,
    \Tile_X2Y8_S2BEGb[6] ,
    \Tile_X2Y8_S2BEGb[5] ,
    \Tile_X2Y8_S2BEGb[4] ,
    \Tile_X2Y8_S2BEGb[3] ,
    \Tile_X2Y8_S2BEGb[2] ,
    \Tile_X2Y8_S2BEGb[1] ,
    \Tile_X2Y8_S2BEGb[0] }),
    .S2END({\Tile_X2Y7_S2BEGb[7] ,
    \Tile_X2Y7_S2BEGb[6] ,
    \Tile_X2Y7_S2BEGb[5] ,
    \Tile_X2Y7_S2BEGb[4] ,
    \Tile_X2Y7_S2BEGb[3] ,
    \Tile_X2Y7_S2BEGb[2] ,
    \Tile_X2Y7_S2BEGb[1] ,
    \Tile_X2Y7_S2BEGb[0] }),
    .S2MID({\Tile_X2Y7_S2BEG[7] ,
    \Tile_X2Y7_S2BEG[6] ,
    \Tile_X2Y7_S2BEG[5] ,
    \Tile_X2Y7_S2BEG[4] ,
    \Tile_X2Y7_S2BEG[3] ,
    \Tile_X2Y7_S2BEG[2] ,
    \Tile_X2Y7_S2BEG[1] ,
    \Tile_X2Y7_S2BEG[0] }),
    .S4BEG({\Tile_X2Y8_S4BEG[15] ,
    \Tile_X2Y8_S4BEG[14] ,
    \Tile_X2Y8_S4BEG[13] ,
    \Tile_X2Y8_S4BEG[12] ,
    \Tile_X2Y8_S4BEG[11] ,
    \Tile_X2Y8_S4BEG[10] ,
    \Tile_X2Y8_S4BEG[9] ,
    \Tile_X2Y8_S4BEG[8] ,
    \Tile_X2Y8_S4BEG[7] ,
    \Tile_X2Y8_S4BEG[6] ,
    \Tile_X2Y8_S4BEG[5] ,
    \Tile_X2Y8_S4BEG[4] ,
    \Tile_X2Y8_S4BEG[3] ,
    \Tile_X2Y8_S4BEG[2] ,
    \Tile_X2Y8_S4BEG[1] ,
    \Tile_X2Y8_S4BEG[0] }),
    .S4END({\Tile_X2Y7_S4BEG[15] ,
    \Tile_X2Y7_S4BEG[14] ,
    \Tile_X2Y7_S4BEG[13] ,
    \Tile_X2Y7_S4BEG[12] ,
    \Tile_X2Y7_S4BEG[11] ,
    \Tile_X2Y7_S4BEG[10] ,
    \Tile_X2Y7_S4BEG[9] ,
    \Tile_X2Y7_S4BEG[8] ,
    \Tile_X2Y7_S4BEG[7] ,
    \Tile_X2Y7_S4BEG[6] ,
    \Tile_X2Y7_S4BEG[5] ,
    \Tile_X2Y7_S4BEG[4] ,
    \Tile_X2Y7_S4BEG[3] ,
    \Tile_X2Y7_S4BEG[2] ,
    \Tile_X2Y7_S4BEG[1] ,
    \Tile_X2Y7_S4BEG[0] }),
    .SS4BEG({\Tile_X2Y8_SS4BEG[15] ,
    \Tile_X2Y8_SS4BEG[14] ,
    \Tile_X2Y8_SS4BEG[13] ,
    \Tile_X2Y8_SS4BEG[12] ,
    \Tile_X2Y8_SS4BEG[11] ,
    \Tile_X2Y8_SS4BEG[10] ,
    \Tile_X2Y8_SS4BEG[9] ,
    \Tile_X2Y8_SS4BEG[8] ,
    \Tile_X2Y8_SS4BEG[7] ,
    \Tile_X2Y8_SS4BEG[6] ,
    \Tile_X2Y8_SS4BEG[5] ,
    \Tile_X2Y8_SS4BEG[4] ,
    \Tile_X2Y8_SS4BEG[3] ,
    \Tile_X2Y8_SS4BEG[2] ,
    \Tile_X2Y8_SS4BEG[1] ,
    \Tile_X2Y8_SS4BEG[0] }),
    .SS4END({\Tile_X2Y7_SS4BEG[15] ,
    \Tile_X2Y7_SS4BEG[14] ,
    \Tile_X2Y7_SS4BEG[13] ,
    \Tile_X2Y7_SS4BEG[12] ,
    \Tile_X2Y7_SS4BEG[11] ,
    \Tile_X2Y7_SS4BEG[10] ,
    \Tile_X2Y7_SS4BEG[9] ,
    \Tile_X2Y7_SS4BEG[8] ,
    \Tile_X2Y7_SS4BEG[7] ,
    \Tile_X2Y7_SS4BEG[6] ,
    \Tile_X2Y7_SS4BEG[5] ,
    \Tile_X2Y7_SS4BEG[4] ,
    \Tile_X2Y7_SS4BEG[3] ,
    \Tile_X2Y7_SS4BEG[2] ,
    \Tile_X2Y7_SS4BEG[1] ,
    \Tile_X2Y7_SS4BEG[0] }),
    .W1BEG({\Tile_X2Y8_W1BEG[3] ,
    \Tile_X2Y8_W1BEG[2] ,
    \Tile_X2Y8_W1BEG[1] ,
    \Tile_X2Y8_W1BEG[0] }),
    .W1END({\Tile_X3Y8_W1BEG[3] ,
    \Tile_X3Y8_W1BEG[2] ,
    \Tile_X3Y8_W1BEG[1] ,
    \Tile_X3Y8_W1BEG[0] }),
    .W2BEG({\Tile_X2Y8_W2BEG[7] ,
    \Tile_X2Y8_W2BEG[6] ,
    \Tile_X2Y8_W2BEG[5] ,
    \Tile_X2Y8_W2BEG[4] ,
    \Tile_X2Y8_W2BEG[3] ,
    \Tile_X2Y8_W2BEG[2] ,
    \Tile_X2Y8_W2BEG[1] ,
    \Tile_X2Y8_W2BEG[0] }),
    .W2BEGb({\Tile_X2Y8_W2BEGb[7] ,
    \Tile_X2Y8_W2BEGb[6] ,
    \Tile_X2Y8_W2BEGb[5] ,
    \Tile_X2Y8_W2BEGb[4] ,
    \Tile_X2Y8_W2BEGb[3] ,
    \Tile_X2Y8_W2BEGb[2] ,
    \Tile_X2Y8_W2BEGb[1] ,
    \Tile_X2Y8_W2BEGb[0] }),
    .W2END({\Tile_X3Y8_W2BEGb[7] ,
    \Tile_X3Y8_W2BEGb[6] ,
    \Tile_X3Y8_W2BEGb[5] ,
    \Tile_X3Y8_W2BEGb[4] ,
    \Tile_X3Y8_W2BEGb[3] ,
    \Tile_X3Y8_W2BEGb[2] ,
    \Tile_X3Y8_W2BEGb[1] ,
    \Tile_X3Y8_W2BEGb[0] }),
    .W2MID({\Tile_X3Y8_W2BEG[7] ,
    \Tile_X3Y8_W2BEG[6] ,
    \Tile_X3Y8_W2BEG[5] ,
    \Tile_X3Y8_W2BEG[4] ,
    \Tile_X3Y8_W2BEG[3] ,
    \Tile_X3Y8_W2BEG[2] ,
    \Tile_X3Y8_W2BEG[1] ,
    \Tile_X3Y8_W2BEG[0] }),
    .W6BEG({\Tile_X2Y8_W6BEG[11] ,
    \Tile_X2Y8_W6BEG[10] ,
    \Tile_X2Y8_W6BEG[9] ,
    \Tile_X2Y8_W6BEG[8] ,
    \Tile_X2Y8_W6BEG[7] ,
    \Tile_X2Y8_W6BEG[6] ,
    \Tile_X2Y8_W6BEG[5] ,
    \Tile_X2Y8_W6BEG[4] ,
    \Tile_X2Y8_W6BEG[3] ,
    \Tile_X2Y8_W6BEG[2] ,
    \Tile_X2Y8_W6BEG[1] ,
    \Tile_X2Y8_W6BEG[0] }),
    .W6END({\Tile_X3Y8_W6BEG[11] ,
    \Tile_X3Y8_W6BEG[10] ,
    \Tile_X3Y8_W6BEG[9] ,
    \Tile_X3Y8_W6BEG[8] ,
    \Tile_X3Y8_W6BEG[7] ,
    \Tile_X3Y8_W6BEG[6] ,
    \Tile_X3Y8_W6BEG[5] ,
    \Tile_X3Y8_W6BEG[4] ,
    \Tile_X3Y8_W6BEG[3] ,
    \Tile_X3Y8_W6BEG[2] ,
    \Tile_X3Y8_W6BEG[1] ,
    \Tile_X3Y8_W6BEG[0] }),
    .WW4BEG({\Tile_X2Y8_WW4BEG[15] ,
    \Tile_X2Y8_WW4BEG[14] ,
    \Tile_X2Y8_WW4BEG[13] ,
    \Tile_X2Y8_WW4BEG[12] ,
    \Tile_X2Y8_WW4BEG[11] ,
    \Tile_X2Y8_WW4BEG[10] ,
    \Tile_X2Y8_WW4BEG[9] ,
    \Tile_X2Y8_WW4BEG[8] ,
    \Tile_X2Y8_WW4BEG[7] ,
    \Tile_X2Y8_WW4BEG[6] ,
    \Tile_X2Y8_WW4BEG[5] ,
    \Tile_X2Y8_WW4BEG[4] ,
    \Tile_X2Y8_WW4BEG[3] ,
    \Tile_X2Y8_WW4BEG[2] ,
    \Tile_X2Y8_WW4BEG[1] ,
    \Tile_X2Y8_WW4BEG[0] }),
    .WW4END({\Tile_X3Y8_WW4BEG[15] ,
    \Tile_X3Y8_WW4BEG[14] ,
    \Tile_X3Y8_WW4BEG[13] ,
    \Tile_X3Y8_WW4BEG[12] ,
    \Tile_X3Y8_WW4BEG[11] ,
    \Tile_X3Y8_WW4BEG[10] ,
    \Tile_X3Y8_WW4BEG[9] ,
    \Tile_X3Y8_WW4BEG[8] ,
    \Tile_X3Y8_WW4BEG[7] ,
    \Tile_X3Y8_WW4BEG[6] ,
    \Tile_X3Y8_WW4BEG[5] ,
    \Tile_X3Y8_WW4BEG[4] ,
    \Tile_X3Y8_WW4BEG[3] ,
    \Tile_X3Y8_WW4BEG[2] ,
    \Tile_X3Y8_WW4BEG[1] ,
    \Tile_X3Y8_WW4BEG[0] }));
 S_IO4 Tile_X2Y9_S_IO4 (.A_I_top(Tile_X2Y9_A_I_top),
    .A_O_top(Tile_X2Y9_A_O_top),
    .A_T_top(Tile_X2Y9_A_T_top),
    .B_I_top(Tile_X2Y9_B_I_top),
    .B_O_top(Tile_X2Y9_B_O_top),
    .B_T_top(Tile_X2Y9_B_T_top),
    .C_I_top(Tile_X2Y9_C_I_top),
    .C_O_top(Tile_X2Y9_C_O_top),
    .C_T_top(Tile_X2Y9_C_T_top),
    .Co(Tile_X2Y9_Co),
    .D_I_top(Tile_X2Y9_D_I_top),
    .D_O_top(Tile_X2Y9_D_O_top),
    .D_T_top(Tile_X2Y9_D_T_top),
    .UserCLK(UserCLK),
    .UserCLKo(Tile_X2Y9_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .FrameData({\Tile_X1Y9_FrameData_O[31] ,
    \Tile_X1Y9_FrameData_O[30] ,
    \Tile_X1Y9_FrameData_O[29] ,
    \Tile_X1Y9_FrameData_O[28] ,
    \Tile_X1Y9_FrameData_O[27] ,
    \Tile_X1Y9_FrameData_O[26] ,
    \Tile_X1Y9_FrameData_O[25] ,
    \Tile_X1Y9_FrameData_O[24] ,
    \Tile_X1Y9_FrameData_O[23] ,
    \Tile_X1Y9_FrameData_O[22] ,
    \Tile_X1Y9_FrameData_O[21] ,
    \Tile_X1Y9_FrameData_O[20] ,
    \Tile_X1Y9_FrameData_O[19] ,
    \Tile_X1Y9_FrameData_O[18] ,
    \Tile_X1Y9_FrameData_O[17] ,
    \Tile_X1Y9_FrameData_O[16] ,
    \Tile_X1Y9_FrameData_O[15] ,
    \Tile_X1Y9_FrameData_O[14] ,
    \Tile_X1Y9_FrameData_O[13] ,
    \Tile_X1Y9_FrameData_O[12] ,
    \Tile_X1Y9_FrameData_O[11] ,
    \Tile_X1Y9_FrameData_O[10] ,
    \Tile_X1Y9_FrameData_O[9] ,
    \Tile_X1Y9_FrameData_O[8] ,
    \Tile_X1Y9_FrameData_O[7] ,
    \Tile_X1Y9_FrameData_O[6] ,
    \Tile_X1Y9_FrameData_O[5] ,
    \Tile_X1Y9_FrameData_O[4] ,
    \Tile_X1Y9_FrameData_O[3] ,
    \Tile_X1Y9_FrameData_O[2] ,
    \Tile_X1Y9_FrameData_O[1] ,
    \Tile_X1Y9_FrameData_O[0] }),
    .FrameData_O({\Tile_X2Y9_FrameData_O[31] ,
    \Tile_X2Y9_FrameData_O[30] ,
    \Tile_X2Y9_FrameData_O[29] ,
    \Tile_X2Y9_FrameData_O[28] ,
    \Tile_X2Y9_FrameData_O[27] ,
    \Tile_X2Y9_FrameData_O[26] ,
    \Tile_X2Y9_FrameData_O[25] ,
    \Tile_X2Y9_FrameData_O[24] ,
    \Tile_X2Y9_FrameData_O[23] ,
    \Tile_X2Y9_FrameData_O[22] ,
    \Tile_X2Y9_FrameData_O[21] ,
    \Tile_X2Y9_FrameData_O[20] ,
    \Tile_X2Y9_FrameData_O[19] ,
    \Tile_X2Y9_FrameData_O[18] ,
    \Tile_X2Y9_FrameData_O[17] ,
    \Tile_X2Y9_FrameData_O[16] ,
    \Tile_X2Y9_FrameData_O[15] ,
    \Tile_X2Y9_FrameData_O[14] ,
    \Tile_X2Y9_FrameData_O[13] ,
    \Tile_X2Y9_FrameData_O[12] ,
    \Tile_X2Y9_FrameData_O[11] ,
    \Tile_X2Y9_FrameData_O[10] ,
    \Tile_X2Y9_FrameData_O[9] ,
    \Tile_X2Y9_FrameData_O[8] ,
    \Tile_X2Y9_FrameData_O[7] ,
    \Tile_X2Y9_FrameData_O[6] ,
    \Tile_X2Y9_FrameData_O[5] ,
    \Tile_X2Y9_FrameData_O[4] ,
    \Tile_X2Y9_FrameData_O[3] ,
    \Tile_X2Y9_FrameData_O[2] ,
    \Tile_X2Y9_FrameData_O[1] ,
    \Tile_X2Y9_FrameData_O[0] }),
    .FrameStrobe({FrameStrobe[59],
    FrameStrobe[58],
    FrameStrobe[57],
    FrameStrobe[56],
    FrameStrobe[55],
    FrameStrobe[54],
    FrameStrobe[53],
    FrameStrobe[52],
    FrameStrobe[51],
    FrameStrobe[50],
    FrameStrobe[49],
    FrameStrobe[48],
    FrameStrobe[47],
    FrameStrobe[46],
    FrameStrobe[45],
    FrameStrobe[44],
    FrameStrobe[43],
    FrameStrobe[42],
    FrameStrobe[41],
    FrameStrobe[40]}),
    .FrameStrobe_O({\Tile_X2Y9_FrameStrobe_O[19] ,
    \Tile_X2Y9_FrameStrobe_O[18] ,
    \Tile_X2Y9_FrameStrobe_O[17] ,
    \Tile_X2Y9_FrameStrobe_O[16] ,
    \Tile_X2Y9_FrameStrobe_O[15] ,
    \Tile_X2Y9_FrameStrobe_O[14] ,
    \Tile_X2Y9_FrameStrobe_O[13] ,
    \Tile_X2Y9_FrameStrobe_O[12] ,
    \Tile_X2Y9_FrameStrobe_O[11] ,
    \Tile_X2Y9_FrameStrobe_O[10] ,
    \Tile_X2Y9_FrameStrobe_O[9] ,
    \Tile_X2Y9_FrameStrobe_O[8] ,
    \Tile_X2Y9_FrameStrobe_O[7] ,
    \Tile_X2Y9_FrameStrobe_O[6] ,
    \Tile_X2Y9_FrameStrobe_O[5] ,
    \Tile_X2Y9_FrameStrobe_O[4] ,
    \Tile_X2Y9_FrameStrobe_O[3] ,
    \Tile_X2Y9_FrameStrobe_O[2] ,
    \Tile_X2Y9_FrameStrobe_O[1] ,
    \Tile_X2Y9_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X2Y9_N1BEG[3] ,
    \Tile_X2Y9_N1BEG[2] ,
    \Tile_X2Y9_N1BEG[1] ,
    \Tile_X2Y9_N1BEG[0] }),
    .N2BEG({\Tile_X2Y9_N2BEG[7] ,
    \Tile_X2Y9_N2BEG[6] ,
    \Tile_X2Y9_N2BEG[5] ,
    \Tile_X2Y9_N2BEG[4] ,
    \Tile_X2Y9_N2BEG[3] ,
    \Tile_X2Y9_N2BEG[2] ,
    \Tile_X2Y9_N2BEG[1] ,
    \Tile_X2Y9_N2BEG[0] }),
    .N2BEGb({\Tile_X2Y9_N2BEGb[7] ,
    \Tile_X2Y9_N2BEGb[6] ,
    \Tile_X2Y9_N2BEGb[5] ,
    \Tile_X2Y9_N2BEGb[4] ,
    \Tile_X2Y9_N2BEGb[3] ,
    \Tile_X2Y9_N2BEGb[2] ,
    \Tile_X2Y9_N2BEGb[1] ,
    \Tile_X2Y9_N2BEGb[0] }),
    .N4BEG({\Tile_X2Y9_N4BEG[15] ,
    \Tile_X2Y9_N4BEG[14] ,
    \Tile_X2Y9_N4BEG[13] ,
    \Tile_X2Y9_N4BEG[12] ,
    \Tile_X2Y9_N4BEG[11] ,
    \Tile_X2Y9_N4BEG[10] ,
    \Tile_X2Y9_N4BEG[9] ,
    \Tile_X2Y9_N4BEG[8] ,
    \Tile_X2Y9_N4BEG[7] ,
    \Tile_X2Y9_N4BEG[6] ,
    \Tile_X2Y9_N4BEG[5] ,
    \Tile_X2Y9_N4BEG[4] ,
    \Tile_X2Y9_N4BEG[3] ,
    \Tile_X2Y9_N4BEG[2] ,
    \Tile_X2Y9_N4BEG[1] ,
    \Tile_X2Y9_N4BEG[0] }),
    .NN4BEG({\Tile_X2Y9_NN4BEG[15] ,
    \Tile_X2Y9_NN4BEG[14] ,
    \Tile_X2Y9_NN4BEG[13] ,
    \Tile_X2Y9_NN4BEG[12] ,
    \Tile_X2Y9_NN4BEG[11] ,
    \Tile_X2Y9_NN4BEG[10] ,
    \Tile_X2Y9_NN4BEG[9] ,
    \Tile_X2Y9_NN4BEG[8] ,
    \Tile_X2Y9_NN4BEG[7] ,
    \Tile_X2Y9_NN4BEG[6] ,
    \Tile_X2Y9_NN4BEG[5] ,
    \Tile_X2Y9_NN4BEG[4] ,
    \Tile_X2Y9_NN4BEG[3] ,
    \Tile_X2Y9_NN4BEG[2] ,
    \Tile_X2Y9_NN4BEG[1] ,
    \Tile_X2Y9_NN4BEG[0] }),
    .S1END({\Tile_X2Y8_S1BEG[3] ,
    \Tile_X2Y8_S1BEG[2] ,
    \Tile_X2Y8_S1BEG[1] ,
    \Tile_X2Y8_S1BEG[0] }),
    .S2END({\Tile_X2Y8_S2BEGb[7] ,
    \Tile_X2Y8_S2BEGb[6] ,
    \Tile_X2Y8_S2BEGb[5] ,
    \Tile_X2Y8_S2BEGb[4] ,
    \Tile_X2Y8_S2BEGb[3] ,
    \Tile_X2Y8_S2BEGb[2] ,
    \Tile_X2Y8_S2BEGb[1] ,
    \Tile_X2Y8_S2BEGb[0] }),
    .S2MID({\Tile_X2Y8_S2BEG[7] ,
    \Tile_X2Y8_S2BEG[6] ,
    \Tile_X2Y8_S2BEG[5] ,
    \Tile_X2Y8_S2BEG[4] ,
    \Tile_X2Y8_S2BEG[3] ,
    \Tile_X2Y8_S2BEG[2] ,
    \Tile_X2Y8_S2BEG[1] ,
    \Tile_X2Y8_S2BEG[0] }),
    .S4END({\Tile_X2Y8_S4BEG[15] ,
    \Tile_X2Y8_S4BEG[14] ,
    \Tile_X2Y8_S4BEG[13] ,
    \Tile_X2Y8_S4BEG[12] ,
    \Tile_X2Y8_S4BEG[11] ,
    \Tile_X2Y8_S4BEG[10] ,
    \Tile_X2Y8_S4BEG[9] ,
    \Tile_X2Y8_S4BEG[8] ,
    \Tile_X2Y8_S4BEG[7] ,
    \Tile_X2Y8_S4BEG[6] ,
    \Tile_X2Y8_S4BEG[5] ,
    \Tile_X2Y8_S4BEG[4] ,
    \Tile_X2Y8_S4BEG[3] ,
    \Tile_X2Y8_S4BEG[2] ,
    \Tile_X2Y8_S4BEG[1] ,
    \Tile_X2Y8_S4BEG[0] }),
    .SS4END({\Tile_X2Y8_SS4BEG[15] ,
    \Tile_X2Y8_SS4BEG[14] ,
    \Tile_X2Y8_SS4BEG[13] ,
    \Tile_X2Y8_SS4BEG[12] ,
    \Tile_X2Y8_SS4BEG[11] ,
    \Tile_X2Y8_SS4BEG[10] ,
    \Tile_X2Y8_SS4BEG[9] ,
    \Tile_X2Y8_SS4BEG[8] ,
    \Tile_X2Y8_SS4BEG[7] ,
    \Tile_X2Y8_SS4BEG[6] ,
    \Tile_X2Y8_SS4BEG[5] ,
    \Tile_X2Y8_SS4BEG[4] ,
    \Tile_X2Y8_SS4BEG[3] ,
    \Tile_X2Y8_SS4BEG[2] ,
    \Tile_X2Y8_SS4BEG[1] ,
    \Tile_X2Y8_SS4BEG[0] }));
 N_IO4 Tile_X3Y0_N_IO4 (.A_I_top(Tile_X3Y0_A_I_top),
    .A_O_top(Tile_X3Y0_A_O_top),
    .A_T_top(Tile_X3Y0_A_T_top),
    .B_I_top(Tile_X3Y0_B_I_top),
    .B_O_top(Tile_X3Y0_B_O_top),
    .B_T_top(Tile_X3Y0_B_T_top),
    .C_I_top(Tile_X3Y0_C_I_top),
    .C_O_top(Tile_X3Y0_C_O_top),
    .C_T_top(Tile_X3Y0_C_T_top),
    .Ci(Tile_X3Y1_Co),
    .D_I_top(Tile_X3Y0_D_I_top),
    .D_O_top(Tile_X3Y0_D_O_top),
    .D_T_top(Tile_X3Y0_D_T_top),
    .UserCLK(Tile_X3Y1_UserCLKo),
    .UserCLKo(Tile_X3Y0_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .FrameData({\Tile_X2Y0_FrameData_O[31] ,
    \Tile_X2Y0_FrameData_O[30] ,
    \Tile_X2Y0_FrameData_O[29] ,
    \Tile_X2Y0_FrameData_O[28] ,
    \Tile_X2Y0_FrameData_O[27] ,
    \Tile_X2Y0_FrameData_O[26] ,
    \Tile_X2Y0_FrameData_O[25] ,
    \Tile_X2Y0_FrameData_O[24] ,
    \Tile_X2Y0_FrameData_O[23] ,
    \Tile_X2Y0_FrameData_O[22] ,
    \Tile_X2Y0_FrameData_O[21] ,
    \Tile_X2Y0_FrameData_O[20] ,
    \Tile_X2Y0_FrameData_O[19] ,
    \Tile_X2Y0_FrameData_O[18] ,
    \Tile_X2Y0_FrameData_O[17] ,
    \Tile_X2Y0_FrameData_O[16] ,
    \Tile_X2Y0_FrameData_O[15] ,
    \Tile_X2Y0_FrameData_O[14] ,
    \Tile_X2Y0_FrameData_O[13] ,
    \Tile_X2Y0_FrameData_O[12] ,
    \Tile_X2Y0_FrameData_O[11] ,
    \Tile_X2Y0_FrameData_O[10] ,
    \Tile_X2Y0_FrameData_O[9] ,
    \Tile_X2Y0_FrameData_O[8] ,
    \Tile_X2Y0_FrameData_O[7] ,
    \Tile_X2Y0_FrameData_O[6] ,
    \Tile_X2Y0_FrameData_O[5] ,
    \Tile_X2Y0_FrameData_O[4] ,
    \Tile_X2Y0_FrameData_O[3] ,
    \Tile_X2Y0_FrameData_O[2] ,
    \Tile_X2Y0_FrameData_O[1] ,
    \Tile_X2Y0_FrameData_O[0] }),
    .FrameData_O({\Tile_X3Y0_FrameData_O[31] ,
    \Tile_X3Y0_FrameData_O[30] ,
    \Tile_X3Y0_FrameData_O[29] ,
    \Tile_X3Y0_FrameData_O[28] ,
    \Tile_X3Y0_FrameData_O[27] ,
    \Tile_X3Y0_FrameData_O[26] ,
    \Tile_X3Y0_FrameData_O[25] ,
    \Tile_X3Y0_FrameData_O[24] ,
    \Tile_X3Y0_FrameData_O[23] ,
    \Tile_X3Y0_FrameData_O[22] ,
    \Tile_X3Y0_FrameData_O[21] ,
    \Tile_X3Y0_FrameData_O[20] ,
    \Tile_X3Y0_FrameData_O[19] ,
    \Tile_X3Y0_FrameData_O[18] ,
    \Tile_X3Y0_FrameData_O[17] ,
    \Tile_X3Y0_FrameData_O[16] ,
    \Tile_X3Y0_FrameData_O[15] ,
    \Tile_X3Y0_FrameData_O[14] ,
    \Tile_X3Y0_FrameData_O[13] ,
    \Tile_X3Y0_FrameData_O[12] ,
    \Tile_X3Y0_FrameData_O[11] ,
    \Tile_X3Y0_FrameData_O[10] ,
    \Tile_X3Y0_FrameData_O[9] ,
    \Tile_X3Y0_FrameData_O[8] ,
    \Tile_X3Y0_FrameData_O[7] ,
    \Tile_X3Y0_FrameData_O[6] ,
    \Tile_X3Y0_FrameData_O[5] ,
    \Tile_X3Y0_FrameData_O[4] ,
    \Tile_X3Y0_FrameData_O[3] ,
    \Tile_X3Y0_FrameData_O[2] ,
    \Tile_X3Y0_FrameData_O[1] ,
    \Tile_X3Y0_FrameData_O[0] }),
    .FrameStrobe({\Tile_X3Y1_FrameStrobe_O[19] ,
    \Tile_X3Y1_FrameStrobe_O[18] ,
    \Tile_X3Y1_FrameStrobe_O[17] ,
    \Tile_X3Y1_FrameStrobe_O[16] ,
    \Tile_X3Y1_FrameStrobe_O[15] ,
    \Tile_X3Y1_FrameStrobe_O[14] ,
    \Tile_X3Y1_FrameStrobe_O[13] ,
    \Tile_X3Y1_FrameStrobe_O[12] ,
    \Tile_X3Y1_FrameStrobe_O[11] ,
    \Tile_X3Y1_FrameStrobe_O[10] ,
    \Tile_X3Y1_FrameStrobe_O[9] ,
    \Tile_X3Y1_FrameStrobe_O[8] ,
    \Tile_X3Y1_FrameStrobe_O[7] ,
    \Tile_X3Y1_FrameStrobe_O[6] ,
    \Tile_X3Y1_FrameStrobe_O[5] ,
    \Tile_X3Y1_FrameStrobe_O[4] ,
    \Tile_X3Y1_FrameStrobe_O[3] ,
    \Tile_X3Y1_FrameStrobe_O[2] ,
    \Tile_X3Y1_FrameStrobe_O[1] ,
    \Tile_X3Y1_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X3Y0_FrameStrobe_O[19] ,
    \Tile_X3Y0_FrameStrobe_O[18] ,
    \Tile_X3Y0_FrameStrobe_O[17] ,
    \Tile_X3Y0_FrameStrobe_O[16] ,
    \Tile_X3Y0_FrameStrobe_O[15] ,
    \Tile_X3Y0_FrameStrobe_O[14] ,
    \Tile_X3Y0_FrameStrobe_O[13] ,
    \Tile_X3Y0_FrameStrobe_O[12] ,
    \Tile_X3Y0_FrameStrobe_O[11] ,
    \Tile_X3Y0_FrameStrobe_O[10] ,
    \Tile_X3Y0_FrameStrobe_O[9] ,
    \Tile_X3Y0_FrameStrobe_O[8] ,
    \Tile_X3Y0_FrameStrobe_O[7] ,
    \Tile_X3Y0_FrameStrobe_O[6] ,
    \Tile_X3Y0_FrameStrobe_O[5] ,
    \Tile_X3Y0_FrameStrobe_O[4] ,
    \Tile_X3Y0_FrameStrobe_O[3] ,
    \Tile_X3Y0_FrameStrobe_O[2] ,
    \Tile_X3Y0_FrameStrobe_O[1] ,
    \Tile_X3Y0_FrameStrobe_O[0] }),
    .N1END({\Tile_X3Y1_N1BEG[3] ,
    \Tile_X3Y1_N1BEG[2] ,
    \Tile_X3Y1_N1BEG[1] ,
    \Tile_X3Y1_N1BEG[0] }),
    .N2END({\Tile_X3Y1_N2BEGb[7] ,
    \Tile_X3Y1_N2BEGb[6] ,
    \Tile_X3Y1_N2BEGb[5] ,
    \Tile_X3Y1_N2BEGb[4] ,
    \Tile_X3Y1_N2BEGb[3] ,
    \Tile_X3Y1_N2BEGb[2] ,
    \Tile_X3Y1_N2BEGb[1] ,
    \Tile_X3Y1_N2BEGb[0] }),
    .N2MID({\Tile_X3Y1_N2BEG[7] ,
    \Tile_X3Y1_N2BEG[6] ,
    \Tile_X3Y1_N2BEG[5] ,
    \Tile_X3Y1_N2BEG[4] ,
    \Tile_X3Y1_N2BEG[3] ,
    \Tile_X3Y1_N2BEG[2] ,
    \Tile_X3Y1_N2BEG[1] ,
    \Tile_X3Y1_N2BEG[0] }),
    .N4END({\Tile_X3Y1_N4BEG[15] ,
    \Tile_X3Y1_N4BEG[14] ,
    \Tile_X3Y1_N4BEG[13] ,
    \Tile_X3Y1_N4BEG[12] ,
    \Tile_X3Y1_N4BEG[11] ,
    \Tile_X3Y1_N4BEG[10] ,
    \Tile_X3Y1_N4BEG[9] ,
    \Tile_X3Y1_N4BEG[8] ,
    \Tile_X3Y1_N4BEG[7] ,
    \Tile_X3Y1_N4BEG[6] ,
    \Tile_X3Y1_N4BEG[5] ,
    \Tile_X3Y1_N4BEG[4] ,
    \Tile_X3Y1_N4BEG[3] ,
    \Tile_X3Y1_N4BEG[2] ,
    \Tile_X3Y1_N4BEG[1] ,
    \Tile_X3Y1_N4BEG[0] }),
    .NN4END({\Tile_X3Y1_NN4BEG[15] ,
    \Tile_X3Y1_NN4BEG[14] ,
    \Tile_X3Y1_NN4BEG[13] ,
    \Tile_X3Y1_NN4BEG[12] ,
    \Tile_X3Y1_NN4BEG[11] ,
    \Tile_X3Y1_NN4BEG[10] ,
    \Tile_X3Y1_NN4BEG[9] ,
    \Tile_X3Y1_NN4BEG[8] ,
    \Tile_X3Y1_NN4BEG[7] ,
    \Tile_X3Y1_NN4BEG[6] ,
    \Tile_X3Y1_NN4BEG[5] ,
    \Tile_X3Y1_NN4BEG[4] ,
    \Tile_X3Y1_NN4BEG[3] ,
    \Tile_X3Y1_NN4BEG[2] ,
    \Tile_X3Y1_NN4BEG[1] ,
    \Tile_X3Y1_NN4BEG[0] }),
    .S1BEG({\Tile_X3Y0_S1BEG[3] ,
    \Tile_X3Y0_S1BEG[2] ,
    \Tile_X3Y0_S1BEG[1] ,
    \Tile_X3Y0_S1BEG[0] }),
    .S2BEG({\Tile_X3Y0_S2BEG[7] ,
    \Tile_X3Y0_S2BEG[6] ,
    \Tile_X3Y0_S2BEG[5] ,
    \Tile_X3Y0_S2BEG[4] ,
    \Tile_X3Y0_S2BEG[3] ,
    \Tile_X3Y0_S2BEG[2] ,
    \Tile_X3Y0_S2BEG[1] ,
    \Tile_X3Y0_S2BEG[0] }),
    .S2BEGb({\Tile_X3Y0_S2BEGb[7] ,
    \Tile_X3Y0_S2BEGb[6] ,
    \Tile_X3Y0_S2BEGb[5] ,
    \Tile_X3Y0_S2BEGb[4] ,
    \Tile_X3Y0_S2BEGb[3] ,
    \Tile_X3Y0_S2BEGb[2] ,
    \Tile_X3Y0_S2BEGb[1] ,
    \Tile_X3Y0_S2BEGb[0] }),
    .S4BEG({\Tile_X3Y0_S4BEG[15] ,
    \Tile_X3Y0_S4BEG[14] ,
    \Tile_X3Y0_S4BEG[13] ,
    \Tile_X3Y0_S4BEG[12] ,
    \Tile_X3Y0_S4BEG[11] ,
    \Tile_X3Y0_S4BEG[10] ,
    \Tile_X3Y0_S4BEG[9] ,
    \Tile_X3Y0_S4BEG[8] ,
    \Tile_X3Y0_S4BEG[7] ,
    \Tile_X3Y0_S4BEG[6] ,
    \Tile_X3Y0_S4BEG[5] ,
    \Tile_X3Y0_S4BEG[4] ,
    \Tile_X3Y0_S4BEG[3] ,
    \Tile_X3Y0_S4BEG[2] ,
    \Tile_X3Y0_S4BEG[1] ,
    \Tile_X3Y0_S4BEG[0] }),
    .SS4BEG({\Tile_X3Y0_SS4BEG[15] ,
    \Tile_X3Y0_SS4BEG[14] ,
    \Tile_X3Y0_SS4BEG[13] ,
    \Tile_X3Y0_SS4BEG[12] ,
    \Tile_X3Y0_SS4BEG[11] ,
    \Tile_X3Y0_SS4BEG[10] ,
    \Tile_X3Y0_SS4BEG[9] ,
    \Tile_X3Y0_SS4BEG[8] ,
    \Tile_X3Y0_SS4BEG[7] ,
    \Tile_X3Y0_SS4BEG[6] ,
    \Tile_X3Y0_SS4BEG[5] ,
    \Tile_X3Y0_SS4BEG[4] ,
    \Tile_X3Y0_SS4BEG[3] ,
    \Tile_X3Y0_SS4BEG[2] ,
    \Tile_X3Y0_SS4BEG[1] ,
    \Tile_X3Y0_SS4BEG[0] }));
 LUT4AB Tile_X3Y1_LUT4AB (.Ci(Tile_X3Y2_Co),
    .Co(Tile_X3Y1_Co),
    .UserCLK(Tile_X3Y2_UserCLKo),
    .UserCLKo(Tile_X3Y1_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X3Y1_E1BEG[3] ,
    \Tile_X3Y1_E1BEG[2] ,
    \Tile_X3Y1_E1BEG[1] ,
    \Tile_X3Y1_E1BEG[0] }),
    .E1END({\Tile_X2Y1_E1BEG[3] ,
    \Tile_X2Y1_E1BEG[2] ,
    \Tile_X2Y1_E1BEG[1] ,
    \Tile_X2Y1_E1BEG[0] }),
    .E2BEG({\Tile_X3Y1_E2BEG[7] ,
    \Tile_X3Y1_E2BEG[6] ,
    \Tile_X3Y1_E2BEG[5] ,
    \Tile_X3Y1_E2BEG[4] ,
    \Tile_X3Y1_E2BEG[3] ,
    \Tile_X3Y1_E2BEG[2] ,
    \Tile_X3Y1_E2BEG[1] ,
    \Tile_X3Y1_E2BEG[0] }),
    .E2BEGb({\Tile_X3Y1_E2BEGb[7] ,
    \Tile_X3Y1_E2BEGb[6] ,
    \Tile_X3Y1_E2BEGb[5] ,
    \Tile_X3Y1_E2BEGb[4] ,
    \Tile_X3Y1_E2BEGb[3] ,
    \Tile_X3Y1_E2BEGb[2] ,
    \Tile_X3Y1_E2BEGb[1] ,
    \Tile_X3Y1_E2BEGb[0] }),
    .E2END({\Tile_X2Y1_E2BEGb[7] ,
    \Tile_X2Y1_E2BEGb[6] ,
    \Tile_X2Y1_E2BEGb[5] ,
    \Tile_X2Y1_E2BEGb[4] ,
    \Tile_X2Y1_E2BEGb[3] ,
    \Tile_X2Y1_E2BEGb[2] ,
    \Tile_X2Y1_E2BEGb[1] ,
    \Tile_X2Y1_E2BEGb[0] }),
    .E2MID({\Tile_X2Y1_E2BEG[7] ,
    \Tile_X2Y1_E2BEG[6] ,
    \Tile_X2Y1_E2BEG[5] ,
    \Tile_X2Y1_E2BEG[4] ,
    \Tile_X2Y1_E2BEG[3] ,
    \Tile_X2Y1_E2BEG[2] ,
    \Tile_X2Y1_E2BEG[1] ,
    \Tile_X2Y1_E2BEG[0] }),
    .E6BEG({\Tile_X3Y1_E6BEG[11] ,
    \Tile_X3Y1_E6BEG[10] ,
    \Tile_X3Y1_E6BEG[9] ,
    \Tile_X3Y1_E6BEG[8] ,
    \Tile_X3Y1_E6BEG[7] ,
    \Tile_X3Y1_E6BEG[6] ,
    \Tile_X3Y1_E6BEG[5] ,
    \Tile_X3Y1_E6BEG[4] ,
    \Tile_X3Y1_E6BEG[3] ,
    \Tile_X3Y1_E6BEG[2] ,
    \Tile_X3Y1_E6BEG[1] ,
    \Tile_X3Y1_E6BEG[0] }),
    .E6END({\Tile_X2Y1_E6BEG[11] ,
    \Tile_X2Y1_E6BEG[10] ,
    \Tile_X2Y1_E6BEG[9] ,
    \Tile_X2Y1_E6BEG[8] ,
    \Tile_X2Y1_E6BEG[7] ,
    \Tile_X2Y1_E6BEG[6] ,
    \Tile_X2Y1_E6BEG[5] ,
    \Tile_X2Y1_E6BEG[4] ,
    \Tile_X2Y1_E6BEG[3] ,
    \Tile_X2Y1_E6BEG[2] ,
    \Tile_X2Y1_E6BEG[1] ,
    \Tile_X2Y1_E6BEG[0] }),
    .EE4BEG({\Tile_X3Y1_EE4BEG[15] ,
    \Tile_X3Y1_EE4BEG[14] ,
    \Tile_X3Y1_EE4BEG[13] ,
    \Tile_X3Y1_EE4BEG[12] ,
    \Tile_X3Y1_EE4BEG[11] ,
    \Tile_X3Y1_EE4BEG[10] ,
    \Tile_X3Y1_EE4BEG[9] ,
    \Tile_X3Y1_EE4BEG[8] ,
    \Tile_X3Y1_EE4BEG[7] ,
    \Tile_X3Y1_EE4BEG[6] ,
    \Tile_X3Y1_EE4BEG[5] ,
    \Tile_X3Y1_EE4BEG[4] ,
    \Tile_X3Y1_EE4BEG[3] ,
    \Tile_X3Y1_EE4BEG[2] ,
    \Tile_X3Y1_EE4BEG[1] ,
    \Tile_X3Y1_EE4BEG[0] }),
    .EE4END({\Tile_X2Y1_EE4BEG[15] ,
    \Tile_X2Y1_EE4BEG[14] ,
    \Tile_X2Y1_EE4BEG[13] ,
    \Tile_X2Y1_EE4BEG[12] ,
    \Tile_X2Y1_EE4BEG[11] ,
    \Tile_X2Y1_EE4BEG[10] ,
    \Tile_X2Y1_EE4BEG[9] ,
    \Tile_X2Y1_EE4BEG[8] ,
    \Tile_X2Y1_EE4BEG[7] ,
    \Tile_X2Y1_EE4BEG[6] ,
    \Tile_X2Y1_EE4BEG[5] ,
    \Tile_X2Y1_EE4BEG[4] ,
    \Tile_X2Y1_EE4BEG[3] ,
    \Tile_X2Y1_EE4BEG[2] ,
    \Tile_X2Y1_EE4BEG[1] ,
    \Tile_X2Y1_EE4BEG[0] }),
    .FrameData({\Tile_X2Y1_FrameData_O[31] ,
    \Tile_X2Y1_FrameData_O[30] ,
    \Tile_X2Y1_FrameData_O[29] ,
    \Tile_X2Y1_FrameData_O[28] ,
    \Tile_X2Y1_FrameData_O[27] ,
    \Tile_X2Y1_FrameData_O[26] ,
    \Tile_X2Y1_FrameData_O[25] ,
    \Tile_X2Y1_FrameData_O[24] ,
    \Tile_X2Y1_FrameData_O[23] ,
    \Tile_X2Y1_FrameData_O[22] ,
    \Tile_X2Y1_FrameData_O[21] ,
    \Tile_X2Y1_FrameData_O[20] ,
    \Tile_X2Y1_FrameData_O[19] ,
    \Tile_X2Y1_FrameData_O[18] ,
    \Tile_X2Y1_FrameData_O[17] ,
    \Tile_X2Y1_FrameData_O[16] ,
    \Tile_X2Y1_FrameData_O[15] ,
    \Tile_X2Y1_FrameData_O[14] ,
    \Tile_X2Y1_FrameData_O[13] ,
    \Tile_X2Y1_FrameData_O[12] ,
    \Tile_X2Y1_FrameData_O[11] ,
    \Tile_X2Y1_FrameData_O[10] ,
    \Tile_X2Y1_FrameData_O[9] ,
    \Tile_X2Y1_FrameData_O[8] ,
    \Tile_X2Y1_FrameData_O[7] ,
    \Tile_X2Y1_FrameData_O[6] ,
    \Tile_X2Y1_FrameData_O[5] ,
    \Tile_X2Y1_FrameData_O[4] ,
    \Tile_X2Y1_FrameData_O[3] ,
    \Tile_X2Y1_FrameData_O[2] ,
    \Tile_X2Y1_FrameData_O[1] ,
    \Tile_X2Y1_FrameData_O[0] }),
    .FrameData_O({\Tile_X3Y1_FrameData_O[31] ,
    \Tile_X3Y1_FrameData_O[30] ,
    \Tile_X3Y1_FrameData_O[29] ,
    \Tile_X3Y1_FrameData_O[28] ,
    \Tile_X3Y1_FrameData_O[27] ,
    \Tile_X3Y1_FrameData_O[26] ,
    \Tile_X3Y1_FrameData_O[25] ,
    \Tile_X3Y1_FrameData_O[24] ,
    \Tile_X3Y1_FrameData_O[23] ,
    \Tile_X3Y1_FrameData_O[22] ,
    \Tile_X3Y1_FrameData_O[21] ,
    \Tile_X3Y1_FrameData_O[20] ,
    \Tile_X3Y1_FrameData_O[19] ,
    \Tile_X3Y1_FrameData_O[18] ,
    \Tile_X3Y1_FrameData_O[17] ,
    \Tile_X3Y1_FrameData_O[16] ,
    \Tile_X3Y1_FrameData_O[15] ,
    \Tile_X3Y1_FrameData_O[14] ,
    \Tile_X3Y1_FrameData_O[13] ,
    \Tile_X3Y1_FrameData_O[12] ,
    \Tile_X3Y1_FrameData_O[11] ,
    \Tile_X3Y1_FrameData_O[10] ,
    \Tile_X3Y1_FrameData_O[9] ,
    \Tile_X3Y1_FrameData_O[8] ,
    \Tile_X3Y1_FrameData_O[7] ,
    \Tile_X3Y1_FrameData_O[6] ,
    \Tile_X3Y1_FrameData_O[5] ,
    \Tile_X3Y1_FrameData_O[4] ,
    \Tile_X3Y1_FrameData_O[3] ,
    \Tile_X3Y1_FrameData_O[2] ,
    \Tile_X3Y1_FrameData_O[1] ,
    \Tile_X3Y1_FrameData_O[0] }),
    .FrameStrobe({\Tile_X3Y2_FrameStrobe_O[19] ,
    \Tile_X3Y2_FrameStrobe_O[18] ,
    \Tile_X3Y2_FrameStrobe_O[17] ,
    \Tile_X3Y2_FrameStrobe_O[16] ,
    \Tile_X3Y2_FrameStrobe_O[15] ,
    \Tile_X3Y2_FrameStrobe_O[14] ,
    \Tile_X3Y2_FrameStrobe_O[13] ,
    \Tile_X3Y2_FrameStrobe_O[12] ,
    \Tile_X3Y2_FrameStrobe_O[11] ,
    \Tile_X3Y2_FrameStrobe_O[10] ,
    \Tile_X3Y2_FrameStrobe_O[9] ,
    \Tile_X3Y2_FrameStrobe_O[8] ,
    \Tile_X3Y2_FrameStrobe_O[7] ,
    \Tile_X3Y2_FrameStrobe_O[6] ,
    \Tile_X3Y2_FrameStrobe_O[5] ,
    \Tile_X3Y2_FrameStrobe_O[4] ,
    \Tile_X3Y2_FrameStrobe_O[3] ,
    \Tile_X3Y2_FrameStrobe_O[2] ,
    \Tile_X3Y2_FrameStrobe_O[1] ,
    \Tile_X3Y2_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X3Y1_FrameStrobe_O[19] ,
    \Tile_X3Y1_FrameStrobe_O[18] ,
    \Tile_X3Y1_FrameStrobe_O[17] ,
    \Tile_X3Y1_FrameStrobe_O[16] ,
    \Tile_X3Y1_FrameStrobe_O[15] ,
    \Tile_X3Y1_FrameStrobe_O[14] ,
    \Tile_X3Y1_FrameStrobe_O[13] ,
    \Tile_X3Y1_FrameStrobe_O[12] ,
    \Tile_X3Y1_FrameStrobe_O[11] ,
    \Tile_X3Y1_FrameStrobe_O[10] ,
    \Tile_X3Y1_FrameStrobe_O[9] ,
    \Tile_X3Y1_FrameStrobe_O[8] ,
    \Tile_X3Y1_FrameStrobe_O[7] ,
    \Tile_X3Y1_FrameStrobe_O[6] ,
    \Tile_X3Y1_FrameStrobe_O[5] ,
    \Tile_X3Y1_FrameStrobe_O[4] ,
    \Tile_X3Y1_FrameStrobe_O[3] ,
    \Tile_X3Y1_FrameStrobe_O[2] ,
    \Tile_X3Y1_FrameStrobe_O[1] ,
    \Tile_X3Y1_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X3Y1_N1BEG[3] ,
    \Tile_X3Y1_N1BEG[2] ,
    \Tile_X3Y1_N1BEG[1] ,
    \Tile_X3Y1_N1BEG[0] }),
    .N1END({\Tile_X3Y2_N1BEG[3] ,
    \Tile_X3Y2_N1BEG[2] ,
    \Tile_X3Y2_N1BEG[1] ,
    \Tile_X3Y2_N1BEG[0] }),
    .N2BEG({\Tile_X3Y1_N2BEG[7] ,
    \Tile_X3Y1_N2BEG[6] ,
    \Tile_X3Y1_N2BEG[5] ,
    \Tile_X3Y1_N2BEG[4] ,
    \Tile_X3Y1_N2BEG[3] ,
    \Tile_X3Y1_N2BEG[2] ,
    \Tile_X3Y1_N2BEG[1] ,
    \Tile_X3Y1_N2BEG[0] }),
    .N2BEGb({\Tile_X3Y1_N2BEGb[7] ,
    \Tile_X3Y1_N2BEGb[6] ,
    \Tile_X3Y1_N2BEGb[5] ,
    \Tile_X3Y1_N2BEGb[4] ,
    \Tile_X3Y1_N2BEGb[3] ,
    \Tile_X3Y1_N2BEGb[2] ,
    \Tile_X3Y1_N2BEGb[1] ,
    \Tile_X3Y1_N2BEGb[0] }),
    .N2END({\Tile_X3Y2_N2BEGb[7] ,
    \Tile_X3Y2_N2BEGb[6] ,
    \Tile_X3Y2_N2BEGb[5] ,
    \Tile_X3Y2_N2BEGb[4] ,
    \Tile_X3Y2_N2BEGb[3] ,
    \Tile_X3Y2_N2BEGb[2] ,
    \Tile_X3Y2_N2BEGb[1] ,
    \Tile_X3Y2_N2BEGb[0] }),
    .N2MID({\Tile_X3Y2_N2BEG[7] ,
    \Tile_X3Y2_N2BEG[6] ,
    \Tile_X3Y2_N2BEG[5] ,
    \Tile_X3Y2_N2BEG[4] ,
    \Tile_X3Y2_N2BEG[3] ,
    \Tile_X3Y2_N2BEG[2] ,
    \Tile_X3Y2_N2BEG[1] ,
    \Tile_X3Y2_N2BEG[0] }),
    .N4BEG({\Tile_X3Y1_N4BEG[15] ,
    \Tile_X3Y1_N4BEG[14] ,
    \Tile_X3Y1_N4BEG[13] ,
    \Tile_X3Y1_N4BEG[12] ,
    \Tile_X3Y1_N4BEG[11] ,
    \Tile_X3Y1_N4BEG[10] ,
    \Tile_X3Y1_N4BEG[9] ,
    \Tile_X3Y1_N4BEG[8] ,
    \Tile_X3Y1_N4BEG[7] ,
    \Tile_X3Y1_N4BEG[6] ,
    \Tile_X3Y1_N4BEG[5] ,
    \Tile_X3Y1_N4BEG[4] ,
    \Tile_X3Y1_N4BEG[3] ,
    \Tile_X3Y1_N4BEG[2] ,
    \Tile_X3Y1_N4BEG[1] ,
    \Tile_X3Y1_N4BEG[0] }),
    .N4END({\Tile_X3Y2_N4BEG[15] ,
    \Tile_X3Y2_N4BEG[14] ,
    \Tile_X3Y2_N4BEG[13] ,
    \Tile_X3Y2_N4BEG[12] ,
    \Tile_X3Y2_N4BEG[11] ,
    \Tile_X3Y2_N4BEG[10] ,
    \Tile_X3Y2_N4BEG[9] ,
    \Tile_X3Y2_N4BEG[8] ,
    \Tile_X3Y2_N4BEG[7] ,
    \Tile_X3Y2_N4BEG[6] ,
    \Tile_X3Y2_N4BEG[5] ,
    \Tile_X3Y2_N4BEG[4] ,
    \Tile_X3Y2_N4BEG[3] ,
    \Tile_X3Y2_N4BEG[2] ,
    \Tile_X3Y2_N4BEG[1] ,
    \Tile_X3Y2_N4BEG[0] }),
    .NN4BEG({\Tile_X3Y1_NN4BEG[15] ,
    \Tile_X3Y1_NN4BEG[14] ,
    \Tile_X3Y1_NN4BEG[13] ,
    \Tile_X3Y1_NN4BEG[12] ,
    \Tile_X3Y1_NN4BEG[11] ,
    \Tile_X3Y1_NN4BEG[10] ,
    \Tile_X3Y1_NN4BEG[9] ,
    \Tile_X3Y1_NN4BEG[8] ,
    \Tile_X3Y1_NN4BEG[7] ,
    \Tile_X3Y1_NN4BEG[6] ,
    \Tile_X3Y1_NN4BEG[5] ,
    \Tile_X3Y1_NN4BEG[4] ,
    \Tile_X3Y1_NN4BEG[3] ,
    \Tile_X3Y1_NN4BEG[2] ,
    \Tile_X3Y1_NN4BEG[1] ,
    \Tile_X3Y1_NN4BEG[0] }),
    .NN4END({\Tile_X3Y2_NN4BEG[15] ,
    \Tile_X3Y2_NN4BEG[14] ,
    \Tile_X3Y2_NN4BEG[13] ,
    \Tile_X3Y2_NN4BEG[12] ,
    \Tile_X3Y2_NN4BEG[11] ,
    \Tile_X3Y2_NN4BEG[10] ,
    \Tile_X3Y2_NN4BEG[9] ,
    \Tile_X3Y2_NN4BEG[8] ,
    \Tile_X3Y2_NN4BEG[7] ,
    \Tile_X3Y2_NN4BEG[6] ,
    \Tile_X3Y2_NN4BEG[5] ,
    \Tile_X3Y2_NN4BEG[4] ,
    \Tile_X3Y2_NN4BEG[3] ,
    \Tile_X3Y2_NN4BEG[2] ,
    \Tile_X3Y2_NN4BEG[1] ,
    \Tile_X3Y2_NN4BEG[0] }),
    .S1BEG({\Tile_X3Y1_S1BEG[3] ,
    \Tile_X3Y1_S1BEG[2] ,
    \Tile_X3Y1_S1BEG[1] ,
    \Tile_X3Y1_S1BEG[0] }),
    .S1END({\Tile_X3Y0_S1BEG[3] ,
    \Tile_X3Y0_S1BEG[2] ,
    \Tile_X3Y0_S1BEG[1] ,
    \Tile_X3Y0_S1BEG[0] }),
    .S2BEG({\Tile_X3Y1_S2BEG[7] ,
    \Tile_X3Y1_S2BEG[6] ,
    \Tile_X3Y1_S2BEG[5] ,
    \Tile_X3Y1_S2BEG[4] ,
    \Tile_X3Y1_S2BEG[3] ,
    \Tile_X3Y1_S2BEG[2] ,
    \Tile_X3Y1_S2BEG[1] ,
    \Tile_X3Y1_S2BEG[0] }),
    .S2BEGb({\Tile_X3Y1_S2BEGb[7] ,
    \Tile_X3Y1_S2BEGb[6] ,
    \Tile_X3Y1_S2BEGb[5] ,
    \Tile_X3Y1_S2BEGb[4] ,
    \Tile_X3Y1_S2BEGb[3] ,
    \Tile_X3Y1_S2BEGb[2] ,
    \Tile_X3Y1_S2BEGb[1] ,
    \Tile_X3Y1_S2BEGb[0] }),
    .S2END({\Tile_X3Y0_S2BEGb[7] ,
    \Tile_X3Y0_S2BEGb[6] ,
    \Tile_X3Y0_S2BEGb[5] ,
    \Tile_X3Y0_S2BEGb[4] ,
    \Tile_X3Y0_S2BEGb[3] ,
    \Tile_X3Y0_S2BEGb[2] ,
    \Tile_X3Y0_S2BEGb[1] ,
    \Tile_X3Y0_S2BEGb[0] }),
    .S2MID({\Tile_X3Y0_S2BEG[7] ,
    \Tile_X3Y0_S2BEG[6] ,
    \Tile_X3Y0_S2BEG[5] ,
    \Tile_X3Y0_S2BEG[4] ,
    \Tile_X3Y0_S2BEG[3] ,
    \Tile_X3Y0_S2BEG[2] ,
    \Tile_X3Y0_S2BEG[1] ,
    \Tile_X3Y0_S2BEG[0] }),
    .S4BEG({\Tile_X3Y1_S4BEG[15] ,
    \Tile_X3Y1_S4BEG[14] ,
    \Tile_X3Y1_S4BEG[13] ,
    \Tile_X3Y1_S4BEG[12] ,
    \Tile_X3Y1_S4BEG[11] ,
    \Tile_X3Y1_S4BEG[10] ,
    \Tile_X3Y1_S4BEG[9] ,
    \Tile_X3Y1_S4BEG[8] ,
    \Tile_X3Y1_S4BEG[7] ,
    \Tile_X3Y1_S4BEG[6] ,
    \Tile_X3Y1_S4BEG[5] ,
    \Tile_X3Y1_S4BEG[4] ,
    \Tile_X3Y1_S4BEG[3] ,
    \Tile_X3Y1_S4BEG[2] ,
    \Tile_X3Y1_S4BEG[1] ,
    \Tile_X3Y1_S4BEG[0] }),
    .S4END({\Tile_X3Y0_S4BEG[15] ,
    \Tile_X3Y0_S4BEG[14] ,
    \Tile_X3Y0_S4BEG[13] ,
    \Tile_X3Y0_S4BEG[12] ,
    \Tile_X3Y0_S4BEG[11] ,
    \Tile_X3Y0_S4BEG[10] ,
    \Tile_X3Y0_S4BEG[9] ,
    \Tile_X3Y0_S4BEG[8] ,
    \Tile_X3Y0_S4BEG[7] ,
    \Tile_X3Y0_S4BEG[6] ,
    \Tile_X3Y0_S4BEG[5] ,
    \Tile_X3Y0_S4BEG[4] ,
    \Tile_X3Y0_S4BEG[3] ,
    \Tile_X3Y0_S4BEG[2] ,
    \Tile_X3Y0_S4BEG[1] ,
    \Tile_X3Y0_S4BEG[0] }),
    .SS4BEG({\Tile_X3Y1_SS4BEG[15] ,
    \Tile_X3Y1_SS4BEG[14] ,
    \Tile_X3Y1_SS4BEG[13] ,
    \Tile_X3Y1_SS4BEG[12] ,
    \Tile_X3Y1_SS4BEG[11] ,
    \Tile_X3Y1_SS4BEG[10] ,
    \Tile_X3Y1_SS4BEG[9] ,
    \Tile_X3Y1_SS4BEG[8] ,
    \Tile_X3Y1_SS4BEG[7] ,
    \Tile_X3Y1_SS4BEG[6] ,
    \Tile_X3Y1_SS4BEG[5] ,
    \Tile_X3Y1_SS4BEG[4] ,
    \Tile_X3Y1_SS4BEG[3] ,
    \Tile_X3Y1_SS4BEG[2] ,
    \Tile_X3Y1_SS4BEG[1] ,
    \Tile_X3Y1_SS4BEG[0] }),
    .SS4END({\Tile_X3Y0_SS4BEG[15] ,
    \Tile_X3Y0_SS4BEG[14] ,
    \Tile_X3Y0_SS4BEG[13] ,
    \Tile_X3Y0_SS4BEG[12] ,
    \Tile_X3Y0_SS4BEG[11] ,
    \Tile_X3Y0_SS4BEG[10] ,
    \Tile_X3Y0_SS4BEG[9] ,
    \Tile_X3Y0_SS4BEG[8] ,
    \Tile_X3Y0_SS4BEG[7] ,
    \Tile_X3Y0_SS4BEG[6] ,
    \Tile_X3Y0_SS4BEG[5] ,
    \Tile_X3Y0_SS4BEG[4] ,
    \Tile_X3Y0_SS4BEG[3] ,
    \Tile_X3Y0_SS4BEG[2] ,
    \Tile_X3Y0_SS4BEG[1] ,
    \Tile_X3Y0_SS4BEG[0] }),
    .W1BEG({\Tile_X3Y1_W1BEG[3] ,
    \Tile_X3Y1_W1BEG[2] ,
    \Tile_X3Y1_W1BEG[1] ,
    \Tile_X3Y1_W1BEG[0] }),
    .W1END({\Tile_X4Y1_W1BEG[3] ,
    \Tile_X4Y1_W1BEG[2] ,
    \Tile_X4Y1_W1BEG[1] ,
    \Tile_X4Y1_W1BEG[0] }),
    .W2BEG({\Tile_X3Y1_W2BEG[7] ,
    \Tile_X3Y1_W2BEG[6] ,
    \Tile_X3Y1_W2BEG[5] ,
    \Tile_X3Y1_W2BEG[4] ,
    \Tile_X3Y1_W2BEG[3] ,
    \Tile_X3Y1_W2BEG[2] ,
    \Tile_X3Y1_W2BEG[1] ,
    \Tile_X3Y1_W2BEG[0] }),
    .W2BEGb({\Tile_X3Y1_W2BEGb[7] ,
    \Tile_X3Y1_W2BEGb[6] ,
    \Tile_X3Y1_W2BEGb[5] ,
    \Tile_X3Y1_W2BEGb[4] ,
    \Tile_X3Y1_W2BEGb[3] ,
    \Tile_X3Y1_W2BEGb[2] ,
    \Tile_X3Y1_W2BEGb[1] ,
    \Tile_X3Y1_W2BEGb[0] }),
    .W2END({\Tile_X4Y1_W2BEGb[7] ,
    \Tile_X4Y1_W2BEGb[6] ,
    \Tile_X4Y1_W2BEGb[5] ,
    \Tile_X4Y1_W2BEGb[4] ,
    \Tile_X4Y1_W2BEGb[3] ,
    \Tile_X4Y1_W2BEGb[2] ,
    \Tile_X4Y1_W2BEGb[1] ,
    \Tile_X4Y1_W2BEGb[0] }),
    .W2MID({\Tile_X4Y1_W2BEG[7] ,
    \Tile_X4Y1_W2BEG[6] ,
    \Tile_X4Y1_W2BEG[5] ,
    \Tile_X4Y1_W2BEG[4] ,
    \Tile_X4Y1_W2BEG[3] ,
    \Tile_X4Y1_W2BEG[2] ,
    \Tile_X4Y1_W2BEG[1] ,
    \Tile_X4Y1_W2BEG[0] }),
    .W6BEG({\Tile_X3Y1_W6BEG[11] ,
    \Tile_X3Y1_W6BEG[10] ,
    \Tile_X3Y1_W6BEG[9] ,
    \Tile_X3Y1_W6BEG[8] ,
    \Tile_X3Y1_W6BEG[7] ,
    \Tile_X3Y1_W6BEG[6] ,
    \Tile_X3Y1_W6BEG[5] ,
    \Tile_X3Y1_W6BEG[4] ,
    \Tile_X3Y1_W6BEG[3] ,
    \Tile_X3Y1_W6BEG[2] ,
    \Tile_X3Y1_W6BEG[1] ,
    \Tile_X3Y1_W6BEG[0] }),
    .W6END({\Tile_X4Y1_W6BEG[11] ,
    \Tile_X4Y1_W6BEG[10] ,
    \Tile_X4Y1_W6BEG[9] ,
    \Tile_X4Y1_W6BEG[8] ,
    \Tile_X4Y1_W6BEG[7] ,
    \Tile_X4Y1_W6BEG[6] ,
    \Tile_X4Y1_W6BEG[5] ,
    \Tile_X4Y1_W6BEG[4] ,
    \Tile_X4Y1_W6BEG[3] ,
    \Tile_X4Y1_W6BEG[2] ,
    \Tile_X4Y1_W6BEG[1] ,
    \Tile_X4Y1_W6BEG[0] }),
    .WW4BEG({\Tile_X3Y1_WW4BEG[15] ,
    \Tile_X3Y1_WW4BEG[14] ,
    \Tile_X3Y1_WW4BEG[13] ,
    \Tile_X3Y1_WW4BEG[12] ,
    \Tile_X3Y1_WW4BEG[11] ,
    \Tile_X3Y1_WW4BEG[10] ,
    \Tile_X3Y1_WW4BEG[9] ,
    \Tile_X3Y1_WW4BEG[8] ,
    \Tile_X3Y1_WW4BEG[7] ,
    \Tile_X3Y1_WW4BEG[6] ,
    \Tile_X3Y1_WW4BEG[5] ,
    \Tile_X3Y1_WW4BEG[4] ,
    \Tile_X3Y1_WW4BEG[3] ,
    \Tile_X3Y1_WW4BEG[2] ,
    \Tile_X3Y1_WW4BEG[1] ,
    \Tile_X3Y1_WW4BEG[0] }),
    .WW4END({\Tile_X4Y1_WW4BEG[15] ,
    \Tile_X4Y1_WW4BEG[14] ,
    \Tile_X4Y1_WW4BEG[13] ,
    \Tile_X4Y1_WW4BEG[12] ,
    \Tile_X4Y1_WW4BEG[11] ,
    \Tile_X4Y1_WW4BEG[10] ,
    \Tile_X4Y1_WW4BEG[9] ,
    \Tile_X4Y1_WW4BEG[8] ,
    \Tile_X4Y1_WW4BEG[7] ,
    \Tile_X4Y1_WW4BEG[6] ,
    \Tile_X4Y1_WW4BEG[5] ,
    \Tile_X4Y1_WW4BEG[4] ,
    \Tile_X4Y1_WW4BEG[3] ,
    \Tile_X4Y1_WW4BEG[2] ,
    \Tile_X4Y1_WW4BEG[1] ,
    \Tile_X4Y1_WW4BEG[0] }));
 LUT4AB Tile_X3Y2_LUT4AB (.Ci(Tile_X3Y3_Co),
    .Co(Tile_X3Y2_Co),
    .UserCLK(Tile_X3Y3_UserCLKo),
    .UserCLKo(Tile_X3Y2_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X3Y2_E1BEG[3] ,
    \Tile_X3Y2_E1BEG[2] ,
    \Tile_X3Y2_E1BEG[1] ,
    \Tile_X3Y2_E1BEG[0] }),
    .E1END({\Tile_X2Y2_E1BEG[3] ,
    \Tile_X2Y2_E1BEG[2] ,
    \Tile_X2Y2_E1BEG[1] ,
    \Tile_X2Y2_E1BEG[0] }),
    .E2BEG({\Tile_X3Y2_E2BEG[7] ,
    \Tile_X3Y2_E2BEG[6] ,
    \Tile_X3Y2_E2BEG[5] ,
    \Tile_X3Y2_E2BEG[4] ,
    \Tile_X3Y2_E2BEG[3] ,
    \Tile_X3Y2_E2BEG[2] ,
    \Tile_X3Y2_E2BEG[1] ,
    \Tile_X3Y2_E2BEG[0] }),
    .E2BEGb({\Tile_X3Y2_E2BEGb[7] ,
    \Tile_X3Y2_E2BEGb[6] ,
    \Tile_X3Y2_E2BEGb[5] ,
    \Tile_X3Y2_E2BEGb[4] ,
    \Tile_X3Y2_E2BEGb[3] ,
    \Tile_X3Y2_E2BEGb[2] ,
    \Tile_X3Y2_E2BEGb[1] ,
    \Tile_X3Y2_E2BEGb[0] }),
    .E2END({\Tile_X2Y2_E2BEGb[7] ,
    \Tile_X2Y2_E2BEGb[6] ,
    \Tile_X2Y2_E2BEGb[5] ,
    \Tile_X2Y2_E2BEGb[4] ,
    \Tile_X2Y2_E2BEGb[3] ,
    \Tile_X2Y2_E2BEGb[2] ,
    \Tile_X2Y2_E2BEGb[1] ,
    \Tile_X2Y2_E2BEGb[0] }),
    .E2MID({\Tile_X2Y2_E2BEG[7] ,
    \Tile_X2Y2_E2BEG[6] ,
    \Tile_X2Y2_E2BEG[5] ,
    \Tile_X2Y2_E2BEG[4] ,
    \Tile_X2Y2_E2BEG[3] ,
    \Tile_X2Y2_E2BEG[2] ,
    \Tile_X2Y2_E2BEG[1] ,
    \Tile_X2Y2_E2BEG[0] }),
    .E6BEG({\Tile_X3Y2_E6BEG[11] ,
    \Tile_X3Y2_E6BEG[10] ,
    \Tile_X3Y2_E6BEG[9] ,
    \Tile_X3Y2_E6BEG[8] ,
    \Tile_X3Y2_E6BEG[7] ,
    \Tile_X3Y2_E6BEG[6] ,
    \Tile_X3Y2_E6BEG[5] ,
    \Tile_X3Y2_E6BEG[4] ,
    \Tile_X3Y2_E6BEG[3] ,
    \Tile_X3Y2_E6BEG[2] ,
    \Tile_X3Y2_E6BEG[1] ,
    \Tile_X3Y2_E6BEG[0] }),
    .E6END({\Tile_X2Y2_E6BEG[11] ,
    \Tile_X2Y2_E6BEG[10] ,
    \Tile_X2Y2_E6BEG[9] ,
    \Tile_X2Y2_E6BEG[8] ,
    \Tile_X2Y2_E6BEG[7] ,
    \Tile_X2Y2_E6BEG[6] ,
    \Tile_X2Y2_E6BEG[5] ,
    \Tile_X2Y2_E6BEG[4] ,
    \Tile_X2Y2_E6BEG[3] ,
    \Tile_X2Y2_E6BEG[2] ,
    \Tile_X2Y2_E6BEG[1] ,
    \Tile_X2Y2_E6BEG[0] }),
    .EE4BEG({\Tile_X3Y2_EE4BEG[15] ,
    \Tile_X3Y2_EE4BEG[14] ,
    \Tile_X3Y2_EE4BEG[13] ,
    \Tile_X3Y2_EE4BEG[12] ,
    \Tile_X3Y2_EE4BEG[11] ,
    \Tile_X3Y2_EE4BEG[10] ,
    \Tile_X3Y2_EE4BEG[9] ,
    \Tile_X3Y2_EE4BEG[8] ,
    \Tile_X3Y2_EE4BEG[7] ,
    \Tile_X3Y2_EE4BEG[6] ,
    \Tile_X3Y2_EE4BEG[5] ,
    \Tile_X3Y2_EE4BEG[4] ,
    \Tile_X3Y2_EE4BEG[3] ,
    \Tile_X3Y2_EE4BEG[2] ,
    \Tile_X3Y2_EE4BEG[1] ,
    \Tile_X3Y2_EE4BEG[0] }),
    .EE4END({\Tile_X2Y2_EE4BEG[15] ,
    \Tile_X2Y2_EE4BEG[14] ,
    \Tile_X2Y2_EE4BEG[13] ,
    \Tile_X2Y2_EE4BEG[12] ,
    \Tile_X2Y2_EE4BEG[11] ,
    \Tile_X2Y2_EE4BEG[10] ,
    \Tile_X2Y2_EE4BEG[9] ,
    \Tile_X2Y2_EE4BEG[8] ,
    \Tile_X2Y2_EE4BEG[7] ,
    \Tile_X2Y2_EE4BEG[6] ,
    \Tile_X2Y2_EE4BEG[5] ,
    \Tile_X2Y2_EE4BEG[4] ,
    \Tile_X2Y2_EE4BEG[3] ,
    \Tile_X2Y2_EE4BEG[2] ,
    \Tile_X2Y2_EE4BEG[1] ,
    \Tile_X2Y2_EE4BEG[0] }),
    .FrameData({\Tile_X2Y2_FrameData_O[31] ,
    \Tile_X2Y2_FrameData_O[30] ,
    \Tile_X2Y2_FrameData_O[29] ,
    \Tile_X2Y2_FrameData_O[28] ,
    \Tile_X2Y2_FrameData_O[27] ,
    \Tile_X2Y2_FrameData_O[26] ,
    \Tile_X2Y2_FrameData_O[25] ,
    \Tile_X2Y2_FrameData_O[24] ,
    \Tile_X2Y2_FrameData_O[23] ,
    \Tile_X2Y2_FrameData_O[22] ,
    \Tile_X2Y2_FrameData_O[21] ,
    \Tile_X2Y2_FrameData_O[20] ,
    \Tile_X2Y2_FrameData_O[19] ,
    \Tile_X2Y2_FrameData_O[18] ,
    \Tile_X2Y2_FrameData_O[17] ,
    \Tile_X2Y2_FrameData_O[16] ,
    \Tile_X2Y2_FrameData_O[15] ,
    \Tile_X2Y2_FrameData_O[14] ,
    \Tile_X2Y2_FrameData_O[13] ,
    \Tile_X2Y2_FrameData_O[12] ,
    \Tile_X2Y2_FrameData_O[11] ,
    \Tile_X2Y2_FrameData_O[10] ,
    \Tile_X2Y2_FrameData_O[9] ,
    \Tile_X2Y2_FrameData_O[8] ,
    \Tile_X2Y2_FrameData_O[7] ,
    \Tile_X2Y2_FrameData_O[6] ,
    \Tile_X2Y2_FrameData_O[5] ,
    \Tile_X2Y2_FrameData_O[4] ,
    \Tile_X2Y2_FrameData_O[3] ,
    \Tile_X2Y2_FrameData_O[2] ,
    \Tile_X2Y2_FrameData_O[1] ,
    \Tile_X2Y2_FrameData_O[0] }),
    .FrameData_O({\Tile_X3Y2_FrameData_O[31] ,
    \Tile_X3Y2_FrameData_O[30] ,
    \Tile_X3Y2_FrameData_O[29] ,
    \Tile_X3Y2_FrameData_O[28] ,
    \Tile_X3Y2_FrameData_O[27] ,
    \Tile_X3Y2_FrameData_O[26] ,
    \Tile_X3Y2_FrameData_O[25] ,
    \Tile_X3Y2_FrameData_O[24] ,
    \Tile_X3Y2_FrameData_O[23] ,
    \Tile_X3Y2_FrameData_O[22] ,
    \Tile_X3Y2_FrameData_O[21] ,
    \Tile_X3Y2_FrameData_O[20] ,
    \Tile_X3Y2_FrameData_O[19] ,
    \Tile_X3Y2_FrameData_O[18] ,
    \Tile_X3Y2_FrameData_O[17] ,
    \Tile_X3Y2_FrameData_O[16] ,
    \Tile_X3Y2_FrameData_O[15] ,
    \Tile_X3Y2_FrameData_O[14] ,
    \Tile_X3Y2_FrameData_O[13] ,
    \Tile_X3Y2_FrameData_O[12] ,
    \Tile_X3Y2_FrameData_O[11] ,
    \Tile_X3Y2_FrameData_O[10] ,
    \Tile_X3Y2_FrameData_O[9] ,
    \Tile_X3Y2_FrameData_O[8] ,
    \Tile_X3Y2_FrameData_O[7] ,
    \Tile_X3Y2_FrameData_O[6] ,
    \Tile_X3Y2_FrameData_O[5] ,
    \Tile_X3Y2_FrameData_O[4] ,
    \Tile_X3Y2_FrameData_O[3] ,
    \Tile_X3Y2_FrameData_O[2] ,
    \Tile_X3Y2_FrameData_O[1] ,
    \Tile_X3Y2_FrameData_O[0] }),
    .FrameStrobe({\Tile_X3Y3_FrameStrobe_O[19] ,
    \Tile_X3Y3_FrameStrobe_O[18] ,
    \Tile_X3Y3_FrameStrobe_O[17] ,
    \Tile_X3Y3_FrameStrobe_O[16] ,
    \Tile_X3Y3_FrameStrobe_O[15] ,
    \Tile_X3Y3_FrameStrobe_O[14] ,
    \Tile_X3Y3_FrameStrobe_O[13] ,
    \Tile_X3Y3_FrameStrobe_O[12] ,
    \Tile_X3Y3_FrameStrobe_O[11] ,
    \Tile_X3Y3_FrameStrobe_O[10] ,
    \Tile_X3Y3_FrameStrobe_O[9] ,
    \Tile_X3Y3_FrameStrobe_O[8] ,
    \Tile_X3Y3_FrameStrobe_O[7] ,
    \Tile_X3Y3_FrameStrobe_O[6] ,
    \Tile_X3Y3_FrameStrobe_O[5] ,
    \Tile_X3Y3_FrameStrobe_O[4] ,
    \Tile_X3Y3_FrameStrobe_O[3] ,
    \Tile_X3Y3_FrameStrobe_O[2] ,
    \Tile_X3Y3_FrameStrobe_O[1] ,
    \Tile_X3Y3_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X3Y2_FrameStrobe_O[19] ,
    \Tile_X3Y2_FrameStrobe_O[18] ,
    \Tile_X3Y2_FrameStrobe_O[17] ,
    \Tile_X3Y2_FrameStrobe_O[16] ,
    \Tile_X3Y2_FrameStrobe_O[15] ,
    \Tile_X3Y2_FrameStrobe_O[14] ,
    \Tile_X3Y2_FrameStrobe_O[13] ,
    \Tile_X3Y2_FrameStrobe_O[12] ,
    \Tile_X3Y2_FrameStrobe_O[11] ,
    \Tile_X3Y2_FrameStrobe_O[10] ,
    \Tile_X3Y2_FrameStrobe_O[9] ,
    \Tile_X3Y2_FrameStrobe_O[8] ,
    \Tile_X3Y2_FrameStrobe_O[7] ,
    \Tile_X3Y2_FrameStrobe_O[6] ,
    \Tile_X3Y2_FrameStrobe_O[5] ,
    \Tile_X3Y2_FrameStrobe_O[4] ,
    \Tile_X3Y2_FrameStrobe_O[3] ,
    \Tile_X3Y2_FrameStrobe_O[2] ,
    \Tile_X3Y2_FrameStrobe_O[1] ,
    \Tile_X3Y2_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X3Y2_N1BEG[3] ,
    \Tile_X3Y2_N1BEG[2] ,
    \Tile_X3Y2_N1BEG[1] ,
    \Tile_X3Y2_N1BEG[0] }),
    .N1END({\Tile_X3Y3_N1BEG[3] ,
    \Tile_X3Y3_N1BEG[2] ,
    \Tile_X3Y3_N1BEG[1] ,
    \Tile_X3Y3_N1BEG[0] }),
    .N2BEG({\Tile_X3Y2_N2BEG[7] ,
    \Tile_X3Y2_N2BEG[6] ,
    \Tile_X3Y2_N2BEG[5] ,
    \Tile_X3Y2_N2BEG[4] ,
    \Tile_X3Y2_N2BEG[3] ,
    \Tile_X3Y2_N2BEG[2] ,
    \Tile_X3Y2_N2BEG[1] ,
    \Tile_X3Y2_N2BEG[0] }),
    .N2BEGb({\Tile_X3Y2_N2BEGb[7] ,
    \Tile_X3Y2_N2BEGb[6] ,
    \Tile_X3Y2_N2BEGb[5] ,
    \Tile_X3Y2_N2BEGb[4] ,
    \Tile_X3Y2_N2BEGb[3] ,
    \Tile_X3Y2_N2BEGb[2] ,
    \Tile_X3Y2_N2BEGb[1] ,
    \Tile_X3Y2_N2BEGb[0] }),
    .N2END({\Tile_X3Y3_N2BEGb[7] ,
    \Tile_X3Y3_N2BEGb[6] ,
    \Tile_X3Y3_N2BEGb[5] ,
    \Tile_X3Y3_N2BEGb[4] ,
    \Tile_X3Y3_N2BEGb[3] ,
    \Tile_X3Y3_N2BEGb[2] ,
    \Tile_X3Y3_N2BEGb[1] ,
    \Tile_X3Y3_N2BEGb[0] }),
    .N2MID({\Tile_X3Y3_N2BEG[7] ,
    \Tile_X3Y3_N2BEG[6] ,
    \Tile_X3Y3_N2BEG[5] ,
    \Tile_X3Y3_N2BEG[4] ,
    \Tile_X3Y3_N2BEG[3] ,
    \Tile_X3Y3_N2BEG[2] ,
    \Tile_X3Y3_N2BEG[1] ,
    \Tile_X3Y3_N2BEG[0] }),
    .N4BEG({\Tile_X3Y2_N4BEG[15] ,
    \Tile_X3Y2_N4BEG[14] ,
    \Tile_X3Y2_N4BEG[13] ,
    \Tile_X3Y2_N4BEG[12] ,
    \Tile_X3Y2_N4BEG[11] ,
    \Tile_X3Y2_N4BEG[10] ,
    \Tile_X3Y2_N4BEG[9] ,
    \Tile_X3Y2_N4BEG[8] ,
    \Tile_X3Y2_N4BEG[7] ,
    \Tile_X3Y2_N4BEG[6] ,
    \Tile_X3Y2_N4BEG[5] ,
    \Tile_X3Y2_N4BEG[4] ,
    \Tile_X3Y2_N4BEG[3] ,
    \Tile_X3Y2_N4BEG[2] ,
    \Tile_X3Y2_N4BEG[1] ,
    \Tile_X3Y2_N4BEG[0] }),
    .N4END({\Tile_X3Y3_N4BEG[15] ,
    \Tile_X3Y3_N4BEG[14] ,
    \Tile_X3Y3_N4BEG[13] ,
    \Tile_X3Y3_N4BEG[12] ,
    \Tile_X3Y3_N4BEG[11] ,
    \Tile_X3Y3_N4BEG[10] ,
    \Tile_X3Y3_N4BEG[9] ,
    \Tile_X3Y3_N4BEG[8] ,
    \Tile_X3Y3_N4BEG[7] ,
    \Tile_X3Y3_N4BEG[6] ,
    \Tile_X3Y3_N4BEG[5] ,
    \Tile_X3Y3_N4BEG[4] ,
    \Tile_X3Y3_N4BEG[3] ,
    \Tile_X3Y3_N4BEG[2] ,
    \Tile_X3Y3_N4BEG[1] ,
    \Tile_X3Y3_N4BEG[0] }),
    .NN4BEG({\Tile_X3Y2_NN4BEG[15] ,
    \Tile_X3Y2_NN4BEG[14] ,
    \Tile_X3Y2_NN4BEG[13] ,
    \Tile_X3Y2_NN4BEG[12] ,
    \Tile_X3Y2_NN4BEG[11] ,
    \Tile_X3Y2_NN4BEG[10] ,
    \Tile_X3Y2_NN4BEG[9] ,
    \Tile_X3Y2_NN4BEG[8] ,
    \Tile_X3Y2_NN4BEG[7] ,
    \Tile_X3Y2_NN4BEG[6] ,
    \Tile_X3Y2_NN4BEG[5] ,
    \Tile_X3Y2_NN4BEG[4] ,
    \Tile_X3Y2_NN4BEG[3] ,
    \Tile_X3Y2_NN4BEG[2] ,
    \Tile_X3Y2_NN4BEG[1] ,
    \Tile_X3Y2_NN4BEG[0] }),
    .NN4END({\Tile_X3Y3_NN4BEG[15] ,
    \Tile_X3Y3_NN4BEG[14] ,
    \Tile_X3Y3_NN4BEG[13] ,
    \Tile_X3Y3_NN4BEG[12] ,
    \Tile_X3Y3_NN4BEG[11] ,
    \Tile_X3Y3_NN4BEG[10] ,
    \Tile_X3Y3_NN4BEG[9] ,
    \Tile_X3Y3_NN4BEG[8] ,
    \Tile_X3Y3_NN4BEG[7] ,
    \Tile_X3Y3_NN4BEG[6] ,
    \Tile_X3Y3_NN4BEG[5] ,
    \Tile_X3Y3_NN4BEG[4] ,
    \Tile_X3Y3_NN4BEG[3] ,
    \Tile_X3Y3_NN4BEG[2] ,
    \Tile_X3Y3_NN4BEG[1] ,
    \Tile_X3Y3_NN4BEG[0] }),
    .S1BEG({\Tile_X3Y2_S1BEG[3] ,
    \Tile_X3Y2_S1BEG[2] ,
    \Tile_X3Y2_S1BEG[1] ,
    \Tile_X3Y2_S1BEG[0] }),
    .S1END({\Tile_X3Y1_S1BEG[3] ,
    \Tile_X3Y1_S1BEG[2] ,
    \Tile_X3Y1_S1BEG[1] ,
    \Tile_X3Y1_S1BEG[0] }),
    .S2BEG({\Tile_X3Y2_S2BEG[7] ,
    \Tile_X3Y2_S2BEG[6] ,
    \Tile_X3Y2_S2BEG[5] ,
    \Tile_X3Y2_S2BEG[4] ,
    \Tile_X3Y2_S2BEG[3] ,
    \Tile_X3Y2_S2BEG[2] ,
    \Tile_X3Y2_S2BEG[1] ,
    \Tile_X3Y2_S2BEG[0] }),
    .S2BEGb({\Tile_X3Y2_S2BEGb[7] ,
    \Tile_X3Y2_S2BEGb[6] ,
    \Tile_X3Y2_S2BEGb[5] ,
    \Tile_X3Y2_S2BEGb[4] ,
    \Tile_X3Y2_S2BEGb[3] ,
    \Tile_X3Y2_S2BEGb[2] ,
    \Tile_X3Y2_S2BEGb[1] ,
    \Tile_X3Y2_S2BEGb[0] }),
    .S2END({\Tile_X3Y1_S2BEGb[7] ,
    \Tile_X3Y1_S2BEGb[6] ,
    \Tile_X3Y1_S2BEGb[5] ,
    \Tile_X3Y1_S2BEGb[4] ,
    \Tile_X3Y1_S2BEGb[3] ,
    \Tile_X3Y1_S2BEGb[2] ,
    \Tile_X3Y1_S2BEGb[1] ,
    \Tile_X3Y1_S2BEGb[0] }),
    .S2MID({\Tile_X3Y1_S2BEG[7] ,
    \Tile_X3Y1_S2BEG[6] ,
    \Tile_X3Y1_S2BEG[5] ,
    \Tile_X3Y1_S2BEG[4] ,
    \Tile_X3Y1_S2BEG[3] ,
    \Tile_X3Y1_S2BEG[2] ,
    \Tile_X3Y1_S2BEG[1] ,
    \Tile_X3Y1_S2BEG[0] }),
    .S4BEG({\Tile_X3Y2_S4BEG[15] ,
    \Tile_X3Y2_S4BEG[14] ,
    \Tile_X3Y2_S4BEG[13] ,
    \Tile_X3Y2_S4BEG[12] ,
    \Tile_X3Y2_S4BEG[11] ,
    \Tile_X3Y2_S4BEG[10] ,
    \Tile_X3Y2_S4BEG[9] ,
    \Tile_X3Y2_S4BEG[8] ,
    \Tile_X3Y2_S4BEG[7] ,
    \Tile_X3Y2_S4BEG[6] ,
    \Tile_X3Y2_S4BEG[5] ,
    \Tile_X3Y2_S4BEG[4] ,
    \Tile_X3Y2_S4BEG[3] ,
    \Tile_X3Y2_S4BEG[2] ,
    \Tile_X3Y2_S4BEG[1] ,
    \Tile_X3Y2_S4BEG[0] }),
    .S4END({\Tile_X3Y1_S4BEG[15] ,
    \Tile_X3Y1_S4BEG[14] ,
    \Tile_X3Y1_S4BEG[13] ,
    \Tile_X3Y1_S4BEG[12] ,
    \Tile_X3Y1_S4BEG[11] ,
    \Tile_X3Y1_S4BEG[10] ,
    \Tile_X3Y1_S4BEG[9] ,
    \Tile_X3Y1_S4BEG[8] ,
    \Tile_X3Y1_S4BEG[7] ,
    \Tile_X3Y1_S4BEG[6] ,
    \Tile_X3Y1_S4BEG[5] ,
    \Tile_X3Y1_S4BEG[4] ,
    \Tile_X3Y1_S4BEG[3] ,
    \Tile_X3Y1_S4BEG[2] ,
    \Tile_X3Y1_S4BEG[1] ,
    \Tile_X3Y1_S4BEG[0] }),
    .SS4BEG({\Tile_X3Y2_SS4BEG[15] ,
    \Tile_X3Y2_SS4BEG[14] ,
    \Tile_X3Y2_SS4BEG[13] ,
    \Tile_X3Y2_SS4BEG[12] ,
    \Tile_X3Y2_SS4BEG[11] ,
    \Tile_X3Y2_SS4BEG[10] ,
    \Tile_X3Y2_SS4BEG[9] ,
    \Tile_X3Y2_SS4BEG[8] ,
    \Tile_X3Y2_SS4BEG[7] ,
    \Tile_X3Y2_SS4BEG[6] ,
    \Tile_X3Y2_SS4BEG[5] ,
    \Tile_X3Y2_SS4BEG[4] ,
    \Tile_X3Y2_SS4BEG[3] ,
    \Tile_X3Y2_SS4BEG[2] ,
    \Tile_X3Y2_SS4BEG[1] ,
    \Tile_X3Y2_SS4BEG[0] }),
    .SS4END({\Tile_X3Y1_SS4BEG[15] ,
    \Tile_X3Y1_SS4BEG[14] ,
    \Tile_X3Y1_SS4BEG[13] ,
    \Tile_X3Y1_SS4BEG[12] ,
    \Tile_X3Y1_SS4BEG[11] ,
    \Tile_X3Y1_SS4BEG[10] ,
    \Tile_X3Y1_SS4BEG[9] ,
    \Tile_X3Y1_SS4BEG[8] ,
    \Tile_X3Y1_SS4BEG[7] ,
    \Tile_X3Y1_SS4BEG[6] ,
    \Tile_X3Y1_SS4BEG[5] ,
    \Tile_X3Y1_SS4BEG[4] ,
    \Tile_X3Y1_SS4BEG[3] ,
    \Tile_X3Y1_SS4BEG[2] ,
    \Tile_X3Y1_SS4BEG[1] ,
    \Tile_X3Y1_SS4BEG[0] }),
    .W1BEG({\Tile_X3Y2_W1BEG[3] ,
    \Tile_X3Y2_W1BEG[2] ,
    \Tile_X3Y2_W1BEG[1] ,
    \Tile_X3Y2_W1BEG[0] }),
    .W1END({\Tile_X4Y2_W1BEG[3] ,
    \Tile_X4Y2_W1BEG[2] ,
    \Tile_X4Y2_W1BEG[1] ,
    \Tile_X4Y2_W1BEG[0] }),
    .W2BEG({\Tile_X3Y2_W2BEG[7] ,
    \Tile_X3Y2_W2BEG[6] ,
    \Tile_X3Y2_W2BEG[5] ,
    \Tile_X3Y2_W2BEG[4] ,
    \Tile_X3Y2_W2BEG[3] ,
    \Tile_X3Y2_W2BEG[2] ,
    \Tile_X3Y2_W2BEG[1] ,
    \Tile_X3Y2_W2BEG[0] }),
    .W2BEGb({\Tile_X3Y2_W2BEGb[7] ,
    \Tile_X3Y2_W2BEGb[6] ,
    \Tile_X3Y2_W2BEGb[5] ,
    \Tile_X3Y2_W2BEGb[4] ,
    \Tile_X3Y2_W2BEGb[3] ,
    \Tile_X3Y2_W2BEGb[2] ,
    \Tile_X3Y2_W2BEGb[1] ,
    \Tile_X3Y2_W2BEGb[0] }),
    .W2END({\Tile_X4Y2_W2BEGb[7] ,
    \Tile_X4Y2_W2BEGb[6] ,
    \Tile_X4Y2_W2BEGb[5] ,
    \Tile_X4Y2_W2BEGb[4] ,
    \Tile_X4Y2_W2BEGb[3] ,
    \Tile_X4Y2_W2BEGb[2] ,
    \Tile_X4Y2_W2BEGb[1] ,
    \Tile_X4Y2_W2BEGb[0] }),
    .W2MID({\Tile_X4Y2_W2BEG[7] ,
    \Tile_X4Y2_W2BEG[6] ,
    \Tile_X4Y2_W2BEG[5] ,
    \Tile_X4Y2_W2BEG[4] ,
    \Tile_X4Y2_W2BEG[3] ,
    \Tile_X4Y2_W2BEG[2] ,
    \Tile_X4Y2_W2BEG[1] ,
    \Tile_X4Y2_W2BEG[0] }),
    .W6BEG({\Tile_X3Y2_W6BEG[11] ,
    \Tile_X3Y2_W6BEG[10] ,
    \Tile_X3Y2_W6BEG[9] ,
    \Tile_X3Y2_W6BEG[8] ,
    \Tile_X3Y2_W6BEG[7] ,
    \Tile_X3Y2_W6BEG[6] ,
    \Tile_X3Y2_W6BEG[5] ,
    \Tile_X3Y2_W6BEG[4] ,
    \Tile_X3Y2_W6BEG[3] ,
    \Tile_X3Y2_W6BEG[2] ,
    \Tile_X3Y2_W6BEG[1] ,
    \Tile_X3Y2_W6BEG[0] }),
    .W6END({\Tile_X4Y2_W6BEG[11] ,
    \Tile_X4Y2_W6BEG[10] ,
    \Tile_X4Y2_W6BEG[9] ,
    \Tile_X4Y2_W6BEG[8] ,
    \Tile_X4Y2_W6BEG[7] ,
    \Tile_X4Y2_W6BEG[6] ,
    \Tile_X4Y2_W6BEG[5] ,
    \Tile_X4Y2_W6BEG[4] ,
    \Tile_X4Y2_W6BEG[3] ,
    \Tile_X4Y2_W6BEG[2] ,
    \Tile_X4Y2_W6BEG[1] ,
    \Tile_X4Y2_W6BEG[0] }),
    .WW4BEG({\Tile_X3Y2_WW4BEG[15] ,
    \Tile_X3Y2_WW4BEG[14] ,
    \Tile_X3Y2_WW4BEG[13] ,
    \Tile_X3Y2_WW4BEG[12] ,
    \Tile_X3Y2_WW4BEG[11] ,
    \Tile_X3Y2_WW4BEG[10] ,
    \Tile_X3Y2_WW4BEG[9] ,
    \Tile_X3Y2_WW4BEG[8] ,
    \Tile_X3Y2_WW4BEG[7] ,
    \Tile_X3Y2_WW4BEG[6] ,
    \Tile_X3Y2_WW4BEG[5] ,
    \Tile_X3Y2_WW4BEG[4] ,
    \Tile_X3Y2_WW4BEG[3] ,
    \Tile_X3Y2_WW4BEG[2] ,
    \Tile_X3Y2_WW4BEG[1] ,
    \Tile_X3Y2_WW4BEG[0] }),
    .WW4END({\Tile_X4Y2_WW4BEG[15] ,
    \Tile_X4Y2_WW4BEG[14] ,
    \Tile_X4Y2_WW4BEG[13] ,
    \Tile_X4Y2_WW4BEG[12] ,
    \Tile_X4Y2_WW4BEG[11] ,
    \Tile_X4Y2_WW4BEG[10] ,
    \Tile_X4Y2_WW4BEG[9] ,
    \Tile_X4Y2_WW4BEG[8] ,
    \Tile_X4Y2_WW4BEG[7] ,
    \Tile_X4Y2_WW4BEG[6] ,
    \Tile_X4Y2_WW4BEG[5] ,
    \Tile_X4Y2_WW4BEG[4] ,
    \Tile_X4Y2_WW4BEG[3] ,
    \Tile_X4Y2_WW4BEG[2] ,
    \Tile_X4Y2_WW4BEG[1] ,
    \Tile_X4Y2_WW4BEG[0] }));
 LUT4AB Tile_X3Y3_LUT4AB (.Ci(Tile_X3Y4_Co),
    .Co(Tile_X3Y3_Co),
    .UserCLK(Tile_X3Y4_UserCLKo),
    .UserCLKo(Tile_X3Y3_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X3Y3_E1BEG[3] ,
    \Tile_X3Y3_E1BEG[2] ,
    \Tile_X3Y3_E1BEG[1] ,
    \Tile_X3Y3_E1BEG[0] }),
    .E1END({\Tile_X2Y3_E1BEG[3] ,
    \Tile_X2Y3_E1BEG[2] ,
    \Tile_X2Y3_E1BEG[1] ,
    \Tile_X2Y3_E1BEG[0] }),
    .E2BEG({\Tile_X3Y3_E2BEG[7] ,
    \Tile_X3Y3_E2BEG[6] ,
    \Tile_X3Y3_E2BEG[5] ,
    \Tile_X3Y3_E2BEG[4] ,
    \Tile_X3Y3_E2BEG[3] ,
    \Tile_X3Y3_E2BEG[2] ,
    \Tile_X3Y3_E2BEG[1] ,
    \Tile_X3Y3_E2BEG[0] }),
    .E2BEGb({\Tile_X3Y3_E2BEGb[7] ,
    \Tile_X3Y3_E2BEGb[6] ,
    \Tile_X3Y3_E2BEGb[5] ,
    \Tile_X3Y3_E2BEGb[4] ,
    \Tile_X3Y3_E2BEGb[3] ,
    \Tile_X3Y3_E2BEGb[2] ,
    \Tile_X3Y3_E2BEGb[1] ,
    \Tile_X3Y3_E2BEGb[0] }),
    .E2END({\Tile_X2Y3_E2BEGb[7] ,
    \Tile_X2Y3_E2BEGb[6] ,
    \Tile_X2Y3_E2BEGb[5] ,
    \Tile_X2Y3_E2BEGb[4] ,
    \Tile_X2Y3_E2BEGb[3] ,
    \Tile_X2Y3_E2BEGb[2] ,
    \Tile_X2Y3_E2BEGb[1] ,
    \Tile_X2Y3_E2BEGb[0] }),
    .E2MID({\Tile_X2Y3_E2BEG[7] ,
    \Tile_X2Y3_E2BEG[6] ,
    \Tile_X2Y3_E2BEG[5] ,
    \Tile_X2Y3_E2BEG[4] ,
    \Tile_X2Y3_E2BEG[3] ,
    \Tile_X2Y3_E2BEG[2] ,
    \Tile_X2Y3_E2BEG[1] ,
    \Tile_X2Y3_E2BEG[0] }),
    .E6BEG({\Tile_X3Y3_E6BEG[11] ,
    \Tile_X3Y3_E6BEG[10] ,
    \Tile_X3Y3_E6BEG[9] ,
    \Tile_X3Y3_E6BEG[8] ,
    \Tile_X3Y3_E6BEG[7] ,
    \Tile_X3Y3_E6BEG[6] ,
    \Tile_X3Y3_E6BEG[5] ,
    \Tile_X3Y3_E6BEG[4] ,
    \Tile_X3Y3_E6BEG[3] ,
    \Tile_X3Y3_E6BEG[2] ,
    \Tile_X3Y3_E6BEG[1] ,
    \Tile_X3Y3_E6BEG[0] }),
    .E6END({\Tile_X2Y3_E6BEG[11] ,
    \Tile_X2Y3_E6BEG[10] ,
    \Tile_X2Y3_E6BEG[9] ,
    \Tile_X2Y3_E6BEG[8] ,
    \Tile_X2Y3_E6BEG[7] ,
    \Tile_X2Y3_E6BEG[6] ,
    \Tile_X2Y3_E6BEG[5] ,
    \Tile_X2Y3_E6BEG[4] ,
    \Tile_X2Y3_E6BEG[3] ,
    \Tile_X2Y3_E6BEG[2] ,
    \Tile_X2Y3_E6BEG[1] ,
    \Tile_X2Y3_E6BEG[0] }),
    .EE4BEG({\Tile_X3Y3_EE4BEG[15] ,
    \Tile_X3Y3_EE4BEG[14] ,
    \Tile_X3Y3_EE4BEG[13] ,
    \Tile_X3Y3_EE4BEG[12] ,
    \Tile_X3Y3_EE4BEG[11] ,
    \Tile_X3Y3_EE4BEG[10] ,
    \Tile_X3Y3_EE4BEG[9] ,
    \Tile_X3Y3_EE4BEG[8] ,
    \Tile_X3Y3_EE4BEG[7] ,
    \Tile_X3Y3_EE4BEG[6] ,
    \Tile_X3Y3_EE4BEG[5] ,
    \Tile_X3Y3_EE4BEG[4] ,
    \Tile_X3Y3_EE4BEG[3] ,
    \Tile_X3Y3_EE4BEG[2] ,
    \Tile_X3Y3_EE4BEG[1] ,
    \Tile_X3Y3_EE4BEG[0] }),
    .EE4END({\Tile_X2Y3_EE4BEG[15] ,
    \Tile_X2Y3_EE4BEG[14] ,
    \Tile_X2Y3_EE4BEG[13] ,
    \Tile_X2Y3_EE4BEG[12] ,
    \Tile_X2Y3_EE4BEG[11] ,
    \Tile_X2Y3_EE4BEG[10] ,
    \Tile_X2Y3_EE4BEG[9] ,
    \Tile_X2Y3_EE4BEG[8] ,
    \Tile_X2Y3_EE4BEG[7] ,
    \Tile_X2Y3_EE4BEG[6] ,
    \Tile_X2Y3_EE4BEG[5] ,
    \Tile_X2Y3_EE4BEG[4] ,
    \Tile_X2Y3_EE4BEG[3] ,
    \Tile_X2Y3_EE4BEG[2] ,
    \Tile_X2Y3_EE4BEG[1] ,
    \Tile_X2Y3_EE4BEG[0] }),
    .FrameData({\Tile_X2Y3_FrameData_O[31] ,
    \Tile_X2Y3_FrameData_O[30] ,
    \Tile_X2Y3_FrameData_O[29] ,
    \Tile_X2Y3_FrameData_O[28] ,
    \Tile_X2Y3_FrameData_O[27] ,
    \Tile_X2Y3_FrameData_O[26] ,
    \Tile_X2Y3_FrameData_O[25] ,
    \Tile_X2Y3_FrameData_O[24] ,
    \Tile_X2Y3_FrameData_O[23] ,
    \Tile_X2Y3_FrameData_O[22] ,
    \Tile_X2Y3_FrameData_O[21] ,
    \Tile_X2Y3_FrameData_O[20] ,
    \Tile_X2Y3_FrameData_O[19] ,
    \Tile_X2Y3_FrameData_O[18] ,
    \Tile_X2Y3_FrameData_O[17] ,
    \Tile_X2Y3_FrameData_O[16] ,
    \Tile_X2Y3_FrameData_O[15] ,
    \Tile_X2Y3_FrameData_O[14] ,
    \Tile_X2Y3_FrameData_O[13] ,
    \Tile_X2Y3_FrameData_O[12] ,
    \Tile_X2Y3_FrameData_O[11] ,
    \Tile_X2Y3_FrameData_O[10] ,
    \Tile_X2Y3_FrameData_O[9] ,
    \Tile_X2Y3_FrameData_O[8] ,
    \Tile_X2Y3_FrameData_O[7] ,
    \Tile_X2Y3_FrameData_O[6] ,
    \Tile_X2Y3_FrameData_O[5] ,
    \Tile_X2Y3_FrameData_O[4] ,
    \Tile_X2Y3_FrameData_O[3] ,
    \Tile_X2Y3_FrameData_O[2] ,
    \Tile_X2Y3_FrameData_O[1] ,
    \Tile_X2Y3_FrameData_O[0] }),
    .FrameData_O({\Tile_X3Y3_FrameData_O[31] ,
    \Tile_X3Y3_FrameData_O[30] ,
    \Tile_X3Y3_FrameData_O[29] ,
    \Tile_X3Y3_FrameData_O[28] ,
    \Tile_X3Y3_FrameData_O[27] ,
    \Tile_X3Y3_FrameData_O[26] ,
    \Tile_X3Y3_FrameData_O[25] ,
    \Tile_X3Y3_FrameData_O[24] ,
    \Tile_X3Y3_FrameData_O[23] ,
    \Tile_X3Y3_FrameData_O[22] ,
    \Tile_X3Y3_FrameData_O[21] ,
    \Tile_X3Y3_FrameData_O[20] ,
    \Tile_X3Y3_FrameData_O[19] ,
    \Tile_X3Y3_FrameData_O[18] ,
    \Tile_X3Y3_FrameData_O[17] ,
    \Tile_X3Y3_FrameData_O[16] ,
    \Tile_X3Y3_FrameData_O[15] ,
    \Tile_X3Y3_FrameData_O[14] ,
    \Tile_X3Y3_FrameData_O[13] ,
    \Tile_X3Y3_FrameData_O[12] ,
    \Tile_X3Y3_FrameData_O[11] ,
    \Tile_X3Y3_FrameData_O[10] ,
    \Tile_X3Y3_FrameData_O[9] ,
    \Tile_X3Y3_FrameData_O[8] ,
    \Tile_X3Y3_FrameData_O[7] ,
    \Tile_X3Y3_FrameData_O[6] ,
    \Tile_X3Y3_FrameData_O[5] ,
    \Tile_X3Y3_FrameData_O[4] ,
    \Tile_X3Y3_FrameData_O[3] ,
    \Tile_X3Y3_FrameData_O[2] ,
    \Tile_X3Y3_FrameData_O[1] ,
    \Tile_X3Y3_FrameData_O[0] }),
    .FrameStrobe({\Tile_X3Y4_FrameStrobe_O[19] ,
    \Tile_X3Y4_FrameStrobe_O[18] ,
    \Tile_X3Y4_FrameStrobe_O[17] ,
    \Tile_X3Y4_FrameStrobe_O[16] ,
    \Tile_X3Y4_FrameStrobe_O[15] ,
    \Tile_X3Y4_FrameStrobe_O[14] ,
    \Tile_X3Y4_FrameStrobe_O[13] ,
    \Tile_X3Y4_FrameStrobe_O[12] ,
    \Tile_X3Y4_FrameStrobe_O[11] ,
    \Tile_X3Y4_FrameStrobe_O[10] ,
    \Tile_X3Y4_FrameStrobe_O[9] ,
    \Tile_X3Y4_FrameStrobe_O[8] ,
    \Tile_X3Y4_FrameStrobe_O[7] ,
    \Tile_X3Y4_FrameStrobe_O[6] ,
    \Tile_X3Y4_FrameStrobe_O[5] ,
    \Tile_X3Y4_FrameStrobe_O[4] ,
    \Tile_X3Y4_FrameStrobe_O[3] ,
    \Tile_X3Y4_FrameStrobe_O[2] ,
    \Tile_X3Y4_FrameStrobe_O[1] ,
    \Tile_X3Y4_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X3Y3_FrameStrobe_O[19] ,
    \Tile_X3Y3_FrameStrobe_O[18] ,
    \Tile_X3Y3_FrameStrobe_O[17] ,
    \Tile_X3Y3_FrameStrobe_O[16] ,
    \Tile_X3Y3_FrameStrobe_O[15] ,
    \Tile_X3Y3_FrameStrobe_O[14] ,
    \Tile_X3Y3_FrameStrobe_O[13] ,
    \Tile_X3Y3_FrameStrobe_O[12] ,
    \Tile_X3Y3_FrameStrobe_O[11] ,
    \Tile_X3Y3_FrameStrobe_O[10] ,
    \Tile_X3Y3_FrameStrobe_O[9] ,
    \Tile_X3Y3_FrameStrobe_O[8] ,
    \Tile_X3Y3_FrameStrobe_O[7] ,
    \Tile_X3Y3_FrameStrobe_O[6] ,
    \Tile_X3Y3_FrameStrobe_O[5] ,
    \Tile_X3Y3_FrameStrobe_O[4] ,
    \Tile_X3Y3_FrameStrobe_O[3] ,
    \Tile_X3Y3_FrameStrobe_O[2] ,
    \Tile_X3Y3_FrameStrobe_O[1] ,
    \Tile_X3Y3_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X3Y3_N1BEG[3] ,
    \Tile_X3Y3_N1BEG[2] ,
    \Tile_X3Y3_N1BEG[1] ,
    \Tile_X3Y3_N1BEG[0] }),
    .N1END({\Tile_X3Y4_N1BEG[3] ,
    \Tile_X3Y4_N1BEG[2] ,
    \Tile_X3Y4_N1BEG[1] ,
    \Tile_X3Y4_N1BEG[0] }),
    .N2BEG({\Tile_X3Y3_N2BEG[7] ,
    \Tile_X3Y3_N2BEG[6] ,
    \Tile_X3Y3_N2BEG[5] ,
    \Tile_X3Y3_N2BEG[4] ,
    \Tile_X3Y3_N2BEG[3] ,
    \Tile_X3Y3_N2BEG[2] ,
    \Tile_X3Y3_N2BEG[1] ,
    \Tile_X3Y3_N2BEG[0] }),
    .N2BEGb({\Tile_X3Y3_N2BEGb[7] ,
    \Tile_X3Y3_N2BEGb[6] ,
    \Tile_X3Y3_N2BEGb[5] ,
    \Tile_X3Y3_N2BEGb[4] ,
    \Tile_X3Y3_N2BEGb[3] ,
    \Tile_X3Y3_N2BEGb[2] ,
    \Tile_X3Y3_N2BEGb[1] ,
    \Tile_X3Y3_N2BEGb[0] }),
    .N2END({\Tile_X3Y4_N2BEGb[7] ,
    \Tile_X3Y4_N2BEGb[6] ,
    \Tile_X3Y4_N2BEGb[5] ,
    \Tile_X3Y4_N2BEGb[4] ,
    \Tile_X3Y4_N2BEGb[3] ,
    \Tile_X3Y4_N2BEGb[2] ,
    \Tile_X3Y4_N2BEGb[1] ,
    \Tile_X3Y4_N2BEGb[0] }),
    .N2MID({\Tile_X3Y4_N2BEG[7] ,
    \Tile_X3Y4_N2BEG[6] ,
    \Tile_X3Y4_N2BEG[5] ,
    \Tile_X3Y4_N2BEG[4] ,
    \Tile_X3Y4_N2BEG[3] ,
    \Tile_X3Y4_N2BEG[2] ,
    \Tile_X3Y4_N2BEG[1] ,
    \Tile_X3Y4_N2BEG[0] }),
    .N4BEG({\Tile_X3Y3_N4BEG[15] ,
    \Tile_X3Y3_N4BEG[14] ,
    \Tile_X3Y3_N4BEG[13] ,
    \Tile_X3Y3_N4BEG[12] ,
    \Tile_X3Y3_N4BEG[11] ,
    \Tile_X3Y3_N4BEG[10] ,
    \Tile_X3Y3_N4BEG[9] ,
    \Tile_X3Y3_N4BEG[8] ,
    \Tile_X3Y3_N4BEG[7] ,
    \Tile_X3Y3_N4BEG[6] ,
    \Tile_X3Y3_N4BEG[5] ,
    \Tile_X3Y3_N4BEG[4] ,
    \Tile_X3Y3_N4BEG[3] ,
    \Tile_X3Y3_N4BEG[2] ,
    \Tile_X3Y3_N4BEG[1] ,
    \Tile_X3Y3_N4BEG[0] }),
    .N4END({\Tile_X3Y4_N4BEG[15] ,
    \Tile_X3Y4_N4BEG[14] ,
    \Tile_X3Y4_N4BEG[13] ,
    \Tile_X3Y4_N4BEG[12] ,
    \Tile_X3Y4_N4BEG[11] ,
    \Tile_X3Y4_N4BEG[10] ,
    \Tile_X3Y4_N4BEG[9] ,
    \Tile_X3Y4_N4BEG[8] ,
    \Tile_X3Y4_N4BEG[7] ,
    \Tile_X3Y4_N4BEG[6] ,
    \Tile_X3Y4_N4BEG[5] ,
    \Tile_X3Y4_N4BEG[4] ,
    \Tile_X3Y4_N4BEG[3] ,
    \Tile_X3Y4_N4BEG[2] ,
    \Tile_X3Y4_N4BEG[1] ,
    \Tile_X3Y4_N4BEG[0] }),
    .NN4BEG({\Tile_X3Y3_NN4BEG[15] ,
    \Tile_X3Y3_NN4BEG[14] ,
    \Tile_X3Y3_NN4BEG[13] ,
    \Tile_X3Y3_NN4BEG[12] ,
    \Tile_X3Y3_NN4BEG[11] ,
    \Tile_X3Y3_NN4BEG[10] ,
    \Tile_X3Y3_NN4BEG[9] ,
    \Tile_X3Y3_NN4BEG[8] ,
    \Tile_X3Y3_NN4BEG[7] ,
    \Tile_X3Y3_NN4BEG[6] ,
    \Tile_X3Y3_NN4BEG[5] ,
    \Tile_X3Y3_NN4BEG[4] ,
    \Tile_X3Y3_NN4BEG[3] ,
    \Tile_X3Y3_NN4BEG[2] ,
    \Tile_X3Y3_NN4BEG[1] ,
    \Tile_X3Y3_NN4BEG[0] }),
    .NN4END({\Tile_X3Y4_NN4BEG[15] ,
    \Tile_X3Y4_NN4BEG[14] ,
    \Tile_X3Y4_NN4BEG[13] ,
    \Tile_X3Y4_NN4BEG[12] ,
    \Tile_X3Y4_NN4BEG[11] ,
    \Tile_X3Y4_NN4BEG[10] ,
    \Tile_X3Y4_NN4BEG[9] ,
    \Tile_X3Y4_NN4BEG[8] ,
    \Tile_X3Y4_NN4BEG[7] ,
    \Tile_X3Y4_NN4BEG[6] ,
    \Tile_X3Y4_NN4BEG[5] ,
    \Tile_X3Y4_NN4BEG[4] ,
    \Tile_X3Y4_NN4BEG[3] ,
    \Tile_X3Y4_NN4BEG[2] ,
    \Tile_X3Y4_NN4BEG[1] ,
    \Tile_X3Y4_NN4BEG[0] }),
    .S1BEG({\Tile_X3Y3_S1BEG[3] ,
    \Tile_X3Y3_S1BEG[2] ,
    \Tile_X3Y3_S1BEG[1] ,
    \Tile_X3Y3_S1BEG[0] }),
    .S1END({\Tile_X3Y2_S1BEG[3] ,
    \Tile_X3Y2_S1BEG[2] ,
    \Tile_X3Y2_S1BEG[1] ,
    \Tile_X3Y2_S1BEG[0] }),
    .S2BEG({\Tile_X3Y3_S2BEG[7] ,
    \Tile_X3Y3_S2BEG[6] ,
    \Tile_X3Y3_S2BEG[5] ,
    \Tile_X3Y3_S2BEG[4] ,
    \Tile_X3Y3_S2BEG[3] ,
    \Tile_X3Y3_S2BEG[2] ,
    \Tile_X3Y3_S2BEG[1] ,
    \Tile_X3Y3_S2BEG[0] }),
    .S2BEGb({\Tile_X3Y3_S2BEGb[7] ,
    \Tile_X3Y3_S2BEGb[6] ,
    \Tile_X3Y3_S2BEGb[5] ,
    \Tile_X3Y3_S2BEGb[4] ,
    \Tile_X3Y3_S2BEGb[3] ,
    \Tile_X3Y3_S2BEGb[2] ,
    \Tile_X3Y3_S2BEGb[1] ,
    \Tile_X3Y3_S2BEGb[0] }),
    .S2END({\Tile_X3Y2_S2BEGb[7] ,
    \Tile_X3Y2_S2BEGb[6] ,
    \Tile_X3Y2_S2BEGb[5] ,
    \Tile_X3Y2_S2BEGb[4] ,
    \Tile_X3Y2_S2BEGb[3] ,
    \Tile_X3Y2_S2BEGb[2] ,
    \Tile_X3Y2_S2BEGb[1] ,
    \Tile_X3Y2_S2BEGb[0] }),
    .S2MID({\Tile_X3Y2_S2BEG[7] ,
    \Tile_X3Y2_S2BEG[6] ,
    \Tile_X3Y2_S2BEG[5] ,
    \Tile_X3Y2_S2BEG[4] ,
    \Tile_X3Y2_S2BEG[3] ,
    \Tile_X3Y2_S2BEG[2] ,
    \Tile_X3Y2_S2BEG[1] ,
    \Tile_X3Y2_S2BEG[0] }),
    .S4BEG({\Tile_X3Y3_S4BEG[15] ,
    \Tile_X3Y3_S4BEG[14] ,
    \Tile_X3Y3_S4BEG[13] ,
    \Tile_X3Y3_S4BEG[12] ,
    \Tile_X3Y3_S4BEG[11] ,
    \Tile_X3Y3_S4BEG[10] ,
    \Tile_X3Y3_S4BEG[9] ,
    \Tile_X3Y3_S4BEG[8] ,
    \Tile_X3Y3_S4BEG[7] ,
    \Tile_X3Y3_S4BEG[6] ,
    \Tile_X3Y3_S4BEG[5] ,
    \Tile_X3Y3_S4BEG[4] ,
    \Tile_X3Y3_S4BEG[3] ,
    \Tile_X3Y3_S4BEG[2] ,
    \Tile_X3Y3_S4BEG[1] ,
    \Tile_X3Y3_S4BEG[0] }),
    .S4END({\Tile_X3Y2_S4BEG[15] ,
    \Tile_X3Y2_S4BEG[14] ,
    \Tile_X3Y2_S4BEG[13] ,
    \Tile_X3Y2_S4BEG[12] ,
    \Tile_X3Y2_S4BEG[11] ,
    \Tile_X3Y2_S4BEG[10] ,
    \Tile_X3Y2_S4BEG[9] ,
    \Tile_X3Y2_S4BEG[8] ,
    \Tile_X3Y2_S4BEG[7] ,
    \Tile_X3Y2_S4BEG[6] ,
    \Tile_X3Y2_S4BEG[5] ,
    \Tile_X3Y2_S4BEG[4] ,
    \Tile_X3Y2_S4BEG[3] ,
    \Tile_X3Y2_S4BEG[2] ,
    \Tile_X3Y2_S4BEG[1] ,
    \Tile_X3Y2_S4BEG[0] }),
    .SS4BEG({\Tile_X3Y3_SS4BEG[15] ,
    \Tile_X3Y3_SS4BEG[14] ,
    \Tile_X3Y3_SS4BEG[13] ,
    \Tile_X3Y3_SS4BEG[12] ,
    \Tile_X3Y3_SS4BEG[11] ,
    \Tile_X3Y3_SS4BEG[10] ,
    \Tile_X3Y3_SS4BEG[9] ,
    \Tile_X3Y3_SS4BEG[8] ,
    \Tile_X3Y3_SS4BEG[7] ,
    \Tile_X3Y3_SS4BEG[6] ,
    \Tile_X3Y3_SS4BEG[5] ,
    \Tile_X3Y3_SS4BEG[4] ,
    \Tile_X3Y3_SS4BEG[3] ,
    \Tile_X3Y3_SS4BEG[2] ,
    \Tile_X3Y3_SS4BEG[1] ,
    \Tile_X3Y3_SS4BEG[0] }),
    .SS4END({\Tile_X3Y2_SS4BEG[15] ,
    \Tile_X3Y2_SS4BEG[14] ,
    \Tile_X3Y2_SS4BEG[13] ,
    \Tile_X3Y2_SS4BEG[12] ,
    \Tile_X3Y2_SS4BEG[11] ,
    \Tile_X3Y2_SS4BEG[10] ,
    \Tile_X3Y2_SS4BEG[9] ,
    \Tile_X3Y2_SS4BEG[8] ,
    \Tile_X3Y2_SS4BEG[7] ,
    \Tile_X3Y2_SS4BEG[6] ,
    \Tile_X3Y2_SS4BEG[5] ,
    \Tile_X3Y2_SS4BEG[4] ,
    \Tile_X3Y2_SS4BEG[3] ,
    \Tile_X3Y2_SS4BEG[2] ,
    \Tile_X3Y2_SS4BEG[1] ,
    \Tile_X3Y2_SS4BEG[0] }),
    .W1BEG({\Tile_X3Y3_W1BEG[3] ,
    \Tile_X3Y3_W1BEG[2] ,
    \Tile_X3Y3_W1BEG[1] ,
    \Tile_X3Y3_W1BEG[0] }),
    .W1END({\Tile_X4Y3_W1BEG[3] ,
    \Tile_X4Y3_W1BEG[2] ,
    \Tile_X4Y3_W1BEG[1] ,
    \Tile_X4Y3_W1BEG[0] }),
    .W2BEG({\Tile_X3Y3_W2BEG[7] ,
    \Tile_X3Y3_W2BEG[6] ,
    \Tile_X3Y3_W2BEG[5] ,
    \Tile_X3Y3_W2BEG[4] ,
    \Tile_X3Y3_W2BEG[3] ,
    \Tile_X3Y3_W2BEG[2] ,
    \Tile_X3Y3_W2BEG[1] ,
    \Tile_X3Y3_W2BEG[0] }),
    .W2BEGb({\Tile_X3Y3_W2BEGb[7] ,
    \Tile_X3Y3_W2BEGb[6] ,
    \Tile_X3Y3_W2BEGb[5] ,
    \Tile_X3Y3_W2BEGb[4] ,
    \Tile_X3Y3_W2BEGb[3] ,
    \Tile_X3Y3_W2BEGb[2] ,
    \Tile_X3Y3_W2BEGb[1] ,
    \Tile_X3Y3_W2BEGb[0] }),
    .W2END({\Tile_X4Y3_W2BEGb[7] ,
    \Tile_X4Y3_W2BEGb[6] ,
    \Tile_X4Y3_W2BEGb[5] ,
    \Tile_X4Y3_W2BEGb[4] ,
    \Tile_X4Y3_W2BEGb[3] ,
    \Tile_X4Y3_W2BEGb[2] ,
    \Tile_X4Y3_W2BEGb[1] ,
    \Tile_X4Y3_W2BEGb[0] }),
    .W2MID({\Tile_X4Y3_W2BEG[7] ,
    \Tile_X4Y3_W2BEG[6] ,
    \Tile_X4Y3_W2BEG[5] ,
    \Tile_X4Y3_W2BEG[4] ,
    \Tile_X4Y3_W2BEG[3] ,
    \Tile_X4Y3_W2BEG[2] ,
    \Tile_X4Y3_W2BEG[1] ,
    \Tile_X4Y3_W2BEG[0] }),
    .W6BEG({\Tile_X3Y3_W6BEG[11] ,
    \Tile_X3Y3_W6BEG[10] ,
    \Tile_X3Y3_W6BEG[9] ,
    \Tile_X3Y3_W6BEG[8] ,
    \Tile_X3Y3_W6BEG[7] ,
    \Tile_X3Y3_W6BEG[6] ,
    \Tile_X3Y3_W6BEG[5] ,
    \Tile_X3Y3_W6BEG[4] ,
    \Tile_X3Y3_W6BEG[3] ,
    \Tile_X3Y3_W6BEG[2] ,
    \Tile_X3Y3_W6BEG[1] ,
    \Tile_X3Y3_W6BEG[0] }),
    .W6END({\Tile_X4Y3_W6BEG[11] ,
    \Tile_X4Y3_W6BEG[10] ,
    \Tile_X4Y3_W6BEG[9] ,
    \Tile_X4Y3_W6BEG[8] ,
    \Tile_X4Y3_W6BEG[7] ,
    \Tile_X4Y3_W6BEG[6] ,
    \Tile_X4Y3_W6BEG[5] ,
    \Tile_X4Y3_W6BEG[4] ,
    \Tile_X4Y3_W6BEG[3] ,
    \Tile_X4Y3_W6BEG[2] ,
    \Tile_X4Y3_W6BEG[1] ,
    \Tile_X4Y3_W6BEG[0] }),
    .WW4BEG({\Tile_X3Y3_WW4BEG[15] ,
    \Tile_X3Y3_WW4BEG[14] ,
    \Tile_X3Y3_WW4BEG[13] ,
    \Tile_X3Y3_WW4BEG[12] ,
    \Tile_X3Y3_WW4BEG[11] ,
    \Tile_X3Y3_WW4BEG[10] ,
    \Tile_X3Y3_WW4BEG[9] ,
    \Tile_X3Y3_WW4BEG[8] ,
    \Tile_X3Y3_WW4BEG[7] ,
    \Tile_X3Y3_WW4BEG[6] ,
    \Tile_X3Y3_WW4BEG[5] ,
    \Tile_X3Y3_WW4BEG[4] ,
    \Tile_X3Y3_WW4BEG[3] ,
    \Tile_X3Y3_WW4BEG[2] ,
    \Tile_X3Y3_WW4BEG[1] ,
    \Tile_X3Y3_WW4BEG[0] }),
    .WW4END({\Tile_X4Y3_WW4BEG[15] ,
    \Tile_X4Y3_WW4BEG[14] ,
    \Tile_X4Y3_WW4BEG[13] ,
    \Tile_X4Y3_WW4BEG[12] ,
    \Tile_X4Y3_WW4BEG[11] ,
    \Tile_X4Y3_WW4BEG[10] ,
    \Tile_X4Y3_WW4BEG[9] ,
    \Tile_X4Y3_WW4BEG[8] ,
    \Tile_X4Y3_WW4BEG[7] ,
    \Tile_X4Y3_WW4BEG[6] ,
    \Tile_X4Y3_WW4BEG[5] ,
    \Tile_X4Y3_WW4BEG[4] ,
    \Tile_X4Y3_WW4BEG[3] ,
    \Tile_X4Y3_WW4BEG[2] ,
    \Tile_X4Y3_WW4BEG[1] ,
    \Tile_X4Y3_WW4BEG[0] }));
 LUT4AB Tile_X3Y4_LUT4AB (.Ci(Tile_X3Y5_Co),
    .Co(Tile_X3Y4_Co),
    .UserCLK(Tile_X3Y5_UserCLKo),
    .UserCLKo(Tile_X3Y4_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X3Y4_E1BEG[3] ,
    \Tile_X3Y4_E1BEG[2] ,
    \Tile_X3Y4_E1BEG[1] ,
    \Tile_X3Y4_E1BEG[0] }),
    .E1END({\Tile_X2Y4_E1BEG[3] ,
    \Tile_X2Y4_E1BEG[2] ,
    \Tile_X2Y4_E1BEG[1] ,
    \Tile_X2Y4_E1BEG[0] }),
    .E2BEG({\Tile_X3Y4_E2BEG[7] ,
    \Tile_X3Y4_E2BEG[6] ,
    \Tile_X3Y4_E2BEG[5] ,
    \Tile_X3Y4_E2BEG[4] ,
    \Tile_X3Y4_E2BEG[3] ,
    \Tile_X3Y4_E2BEG[2] ,
    \Tile_X3Y4_E2BEG[1] ,
    \Tile_X3Y4_E2BEG[0] }),
    .E2BEGb({\Tile_X3Y4_E2BEGb[7] ,
    \Tile_X3Y4_E2BEGb[6] ,
    \Tile_X3Y4_E2BEGb[5] ,
    \Tile_X3Y4_E2BEGb[4] ,
    \Tile_X3Y4_E2BEGb[3] ,
    \Tile_X3Y4_E2BEGb[2] ,
    \Tile_X3Y4_E2BEGb[1] ,
    \Tile_X3Y4_E2BEGb[0] }),
    .E2END({\Tile_X2Y4_E2BEGb[7] ,
    \Tile_X2Y4_E2BEGb[6] ,
    \Tile_X2Y4_E2BEGb[5] ,
    \Tile_X2Y4_E2BEGb[4] ,
    \Tile_X2Y4_E2BEGb[3] ,
    \Tile_X2Y4_E2BEGb[2] ,
    \Tile_X2Y4_E2BEGb[1] ,
    \Tile_X2Y4_E2BEGb[0] }),
    .E2MID({\Tile_X2Y4_E2BEG[7] ,
    \Tile_X2Y4_E2BEG[6] ,
    \Tile_X2Y4_E2BEG[5] ,
    \Tile_X2Y4_E2BEG[4] ,
    \Tile_X2Y4_E2BEG[3] ,
    \Tile_X2Y4_E2BEG[2] ,
    \Tile_X2Y4_E2BEG[1] ,
    \Tile_X2Y4_E2BEG[0] }),
    .E6BEG({\Tile_X3Y4_E6BEG[11] ,
    \Tile_X3Y4_E6BEG[10] ,
    \Tile_X3Y4_E6BEG[9] ,
    \Tile_X3Y4_E6BEG[8] ,
    \Tile_X3Y4_E6BEG[7] ,
    \Tile_X3Y4_E6BEG[6] ,
    \Tile_X3Y4_E6BEG[5] ,
    \Tile_X3Y4_E6BEG[4] ,
    \Tile_X3Y4_E6BEG[3] ,
    \Tile_X3Y4_E6BEG[2] ,
    \Tile_X3Y4_E6BEG[1] ,
    \Tile_X3Y4_E6BEG[0] }),
    .E6END({\Tile_X2Y4_E6BEG[11] ,
    \Tile_X2Y4_E6BEG[10] ,
    \Tile_X2Y4_E6BEG[9] ,
    \Tile_X2Y4_E6BEG[8] ,
    \Tile_X2Y4_E6BEG[7] ,
    \Tile_X2Y4_E6BEG[6] ,
    \Tile_X2Y4_E6BEG[5] ,
    \Tile_X2Y4_E6BEG[4] ,
    \Tile_X2Y4_E6BEG[3] ,
    \Tile_X2Y4_E6BEG[2] ,
    \Tile_X2Y4_E6BEG[1] ,
    \Tile_X2Y4_E6BEG[0] }),
    .EE4BEG({\Tile_X3Y4_EE4BEG[15] ,
    \Tile_X3Y4_EE4BEG[14] ,
    \Tile_X3Y4_EE4BEG[13] ,
    \Tile_X3Y4_EE4BEG[12] ,
    \Tile_X3Y4_EE4BEG[11] ,
    \Tile_X3Y4_EE4BEG[10] ,
    \Tile_X3Y4_EE4BEG[9] ,
    \Tile_X3Y4_EE4BEG[8] ,
    \Tile_X3Y4_EE4BEG[7] ,
    \Tile_X3Y4_EE4BEG[6] ,
    \Tile_X3Y4_EE4BEG[5] ,
    \Tile_X3Y4_EE4BEG[4] ,
    \Tile_X3Y4_EE4BEG[3] ,
    \Tile_X3Y4_EE4BEG[2] ,
    \Tile_X3Y4_EE4BEG[1] ,
    \Tile_X3Y4_EE4BEG[0] }),
    .EE4END({\Tile_X2Y4_EE4BEG[15] ,
    \Tile_X2Y4_EE4BEG[14] ,
    \Tile_X2Y4_EE4BEG[13] ,
    \Tile_X2Y4_EE4BEG[12] ,
    \Tile_X2Y4_EE4BEG[11] ,
    \Tile_X2Y4_EE4BEG[10] ,
    \Tile_X2Y4_EE4BEG[9] ,
    \Tile_X2Y4_EE4BEG[8] ,
    \Tile_X2Y4_EE4BEG[7] ,
    \Tile_X2Y4_EE4BEG[6] ,
    \Tile_X2Y4_EE4BEG[5] ,
    \Tile_X2Y4_EE4BEG[4] ,
    \Tile_X2Y4_EE4BEG[3] ,
    \Tile_X2Y4_EE4BEG[2] ,
    \Tile_X2Y4_EE4BEG[1] ,
    \Tile_X2Y4_EE4BEG[0] }),
    .FrameData({\Tile_X2Y4_FrameData_O[31] ,
    \Tile_X2Y4_FrameData_O[30] ,
    \Tile_X2Y4_FrameData_O[29] ,
    \Tile_X2Y4_FrameData_O[28] ,
    \Tile_X2Y4_FrameData_O[27] ,
    \Tile_X2Y4_FrameData_O[26] ,
    \Tile_X2Y4_FrameData_O[25] ,
    \Tile_X2Y4_FrameData_O[24] ,
    \Tile_X2Y4_FrameData_O[23] ,
    \Tile_X2Y4_FrameData_O[22] ,
    \Tile_X2Y4_FrameData_O[21] ,
    \Tile_X2Y4_FrameData_O[20] ,
    \Tile_X2Y4_FrameData_O[19] ,
    \Tile_X2Y4_FrameData_O[18] ,
    \Tile_X2Y4_FrameData_O[17] ,
    \Tile_X2Y4_FrameData_O[16] ,
    \Tile_X2Y4_FrameData_O[15] ,
    \Tile_X2Y4_FrameData_O[14] ,
    \Tile_X2Y4_FrameData_O[13] ,
    \Tile_X2Y4_FrameData_O[12] ,
    \Tile_X2Y4_FrameData_O[11] ,
    \Tile_X2Y4_FrameData_O[10] ,
    \Tile_X2Y4_FrameData_O[9] ,
    \Tile_X2Y4_FrameData_O[8] ,
    \Tile_X2Y4_FrameData_O[7] ,
    \Tile_X2Y4_FrameData_O[6] ,
    \Tile_X2Y4_FrameData_O[5] ,
    \Tile_X2Y4_FrameData_O[4] ,
    \Tile_X2Y4_FrameData_O[3] ,
    \Tile_X2Y4_FrameData_O[2] ,
    \Tile_X2Y4_FrameData_O[1] ,
    \Tile_X2Y4_FrameData_O[0] }),
    .FrameData_O({\Tile_X3Y4_FrameData_O[31] ,
    \Tile_X3Y4_FrameData_O[30] ,
    \Tile_X3Y4_FrameData_O[29] ,
    \Tile_X3Y4_FrameData_O[28] ,
    \Tile_X3Y4_FrameData_O[27] ,
    \Tile_X3Y4_FrameData_O[26] ,
    \Tile_X3Y4_FrameData_O[25] ,
    \Tile_X3Y4_FrameData_O[24] ,
    \Tile_X3Y4_FrameData_O[23] ,
    \Tile_X3Y4_FrameData_O[22] ,
    \Tile_X3Y4_FrameData_O[21] ,
    \Tile_X3Y4_FrameData_O[20] ,
    \Tile_X3Y4_FrameData_O[19] ,
    \Tile_X3Y4_FrameData_O[18] ,
    \Tile_X3Y4_FrameData_O[17] ,
    \Tile_X3Y4_FrameData_O[16] ,
    \Tile_X3Y4_FrameData_O[15] ,
    \Tile_X3Y4_FrameData_O[14] ,
    \Tile_X3Y4_FrameData_O[13] ,
    \Tile_X3Y4_FrameData_O[12] ,
    \Tile_X3Y4_FrameData_O[11] ,
    \Tile_X3Y4_FrameData_O[10] ,
    \Tile_X3Y4_FrameData_O[9] ,
    \Tile_X3Y4_FrameData_O[8] ,
    \Tile_X3Y4_FrameData_O[7] ,
    \Tile_X3Y4_FrameData_O[6] ,
    \Tile_X3Y4_FrameData_O[5] ,
    \Tile_X3Y4_FrameData_O[4] ,
    \Tile_X3Y4_FrameData_O[3] ,
    \Tile_X3Y4_FrameData_O[2] ,
    \Tile_X3Y4_FrameData_O[1] ,
    \Tile_X3Y4_FrameData_O[0] }),
    .FrameStrobe({\Tile_X3Y5_FrameStrobe_O[19] ,
    \Tile_X3Y5_FrameStrobe_O[18] ,
    \Tile_X3Y5_FrameStrobe_O[17] ,
    \Tile_X3Y5_FrameStrobe_O[16] ,
    \Tile_X3Y5_FrameStrobe_O[15] ,
    \Tile_X3Y5_FrameStrobe_O[14] ,
    \Tile_X3Y5_FrameStrobe_O[13] ,
    \Tile_X3Y5_FrameStrobe_O[12] ,
    \Tile_X3Y5_FrameStrobe_O[11] ,
    \Tile_X3Y5_FrameStrobe_O[10] ,
    \Tile_X3Y5_FrameStrobe_O[9] ,
    \Tile_X3Y5_FrameStrobe_O[8] ,
    \Tile_X3Y5_FrameStrobe_O[7] ,
    \Tile_X3Y5_FrameStrobe_O[6] ,
    \Tile_X3Y5_FrameStrobe_O[5] ,
    \Tile_X3Y5_FrameStrobe_O[4] ,
    \Tile_X3Y5_FrameStrobe_O[3] ,
    \Tile_X3Y5_FrameStrobe_O[2] ,
    \Tile_X3Y5_FrameStrobe_O[1] ,
    \Tile_X3Y5_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X3Y4_FrameStrobe_O[19] ,
    \Tile_X3Y4_FrameStrobe_O[18] ,
    \Tile_X3Y4_FrameStrobe_O[17] ,
    \Tile_X3Y4_FrameStrobe_O[16] ,
    \Tile_X3Y4_FrameStrobe_O[15] ,
    \Tile_X3Y4_FrameStrobe_O[14] ,
    \Tile_X3Y4_FrameStrobe_O[13] ,
    \Tile_X3Y4_FrameStrobe_O[12] ,
    \Tile_X3Y4_FrameStrobe_O[11] ,
    \Tile_X3Y4_FrameStrobe_O[10] ,
    \Tile_X3Y4_FrameStrobe_O[9] ,
    \Tile_X3Y4_FrameStrobe_O[8] ,
    \Tile_X3Y4_FrameStrobe_O[7] ,
    \Tile_X3Y4_FrameStrobe_O[6] ,
    \Tile_X3Y4_FrameStrobe_O[5] ,
    \Tile_X3Y4_FrameStrobe_O[4] ,
    \Tile_X3Y4_FrameStrobe_O[3] ,
    \Tile_X3Y4_FrameStrobe_O[2] ,
    \Tile_X3Y4_FrameStrobe_O[1] ,
    \Tile_X3Y4_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X3Y4_N1BEG[3] ,
    \Tile_X3Y4_N1BEG[2] ,
    \Tile_X3Y4_N1BEG[1] ,
    \Tile_X3Y4_N1BEG[0] }),
    .N1END({\Tile_X3Y5_N1BEG[3] ,
    \Tile_X3Y5_N1BEG[2] ,
    \Tile_X3Y5_N1BEG[1] ,
    \Tile_X3Y5_N1BEG[0] }),
    .N2BEG({\Tile_X3Y4_N2BEG[7] ,
    \Tile_X3Y4_N2BEG[6] ,
    \Tile_X3Y4_N2BEG[5] ,
    \Tile_X3Y4_N2BEG[4] ,
    \Tile_X3Y4_N2BEG[3] ,
    \Tile_X3Y4_N2BEG[2] ,
    \Tile_X3Y4_N2BEG[1] ,
    \Tile_X3Y4_N2BEG[0] }),
    .N2BEGb({\Tile_X3Y4_N2BEGb[7] ,
    \Tile_X3Y4_N2BEGb[6] ,
    \Tile_X3Y4_N2BEGb[5] ,
    \Tile_X3Y4_N2BEGb[4] ,
    \Tile_X3Y4_N2BEGb[3] ,
    \Tile_X3Y4_N2BEGb[2] ,
    \Tile_X3Y4_N2BEGb[1] ,
    \Tile_X3Y4_N2BEGb[0] }),
    .N2END({\Tile_X3Y5_N2BEGb[7] ,
    \Tile_X3Y5_N2BEGb[6] ,
    \Tile_X3Y5_N2BEGb[5] ,
    \Tile_X3Y5_N2BEGb[4] ,
    \Tile_X3Y5_N2BEGb[3] ,
    \Tile_X3Y5_N2BEGb[2] ,
    \Tile_X3Y5_N2BEGb[1] ,
    \Tile_X3Y5_N2BEGb[0] }),
    .N2MID({\Tile_X3Y5_N2BEG[7] ,
    \Tile_X3Y5_N2BEG[6] ,
    \Tile_X3Y5_N2BEG[5] ,
    \Tile_X3Y5_N2BEG[4] ,
    \Tile_X3Y5_N2BEG[3] ,
    \Tile_X3Y5_N2BEG[2] ,
    \Tile_X3Y5_N2BEG[1] ,
    \Tile_X3Y5_N2BEG[0] }),
    .N4BEG({\Tile_X3Y4_N4BEG[15] ,
    \Tile_X3Y4_N4BEG[14] ,
    \Tile_X3Y4_N4BEG[13] ,
    \Tile_X3Y4_N4BEG[12] ,
    \Tile_X3Y4_N4BEG[11] ,
    \Tile_X3Y4_N4BEG[10] ,
    \Tile_X3Y4_N4BEG[9] ,
    \Tile_X3Y4_N4BEG[8] ,
    \Tile_X3Y4_N4BEG[7] ,
    \Tile_X3Y4_N4BEG[6] ,
    \Tile_X3Y4_N4BEG[5] ,
    \Tile_X3Y4_N4BEG[4] ,
    \Tile_X3Y4_N4BEG[3] ,
    \Tile_X3Y4_N4BEG[2] ,
    \Tile_X3Y4_N4BEG[1] ,
    \Tile_X3Y4_N4BEG[0] }),
    .N4END({\Tile_X3Y5_N4BEG[15] ,
    \Tile_X3Y5_N4BEG[14] ,
    \Tile_X3Y5_N4BEG[13] ,
    \Tile_X3Y5_N4BEG[12] ,
    \Tile_X3Y5_N4BEG[11] ,
    \Tile_X3Y5_N4BEG[10] ,
    \Tile_X3Y5_N4BEG[9] ,
    \Tile_X3Y5_N4BEG[8] ,
    \Tile_X3Y5_N4BEG[7] ,
    \Tile_X3Y5_N4BEG[6] ,
    \Tile_X3Y5_N4BEG[5] ,
    \Tile_X3Y5_N4BEG[4] ,
    \Tile_X3Y5_N4BEG[3] ,
    \Tile_X3Y5_N4BEG[2] ,
    \Tile_X3Y5_N4BEG[1] ,
    \Tile_X3Y5_N4BEG[0] }),
    .NN4BEG({\Tile_X3Y4_NN4BEG[15] ,
    \Tile_X3Y4_NN4BEG[14] ,
    \Tile_X3Y4_NN4BEG[13] ,
    \Tile_X3Y4_NN4BEG[12] ,
    \Tile_X3Y4_NN4BEG[11] ,
    \Tile_X3Y4_NN4BEG[10] ,
    \Tile_X3Y4_NN4BEG[9] ,
    \Tile_X3Y4_NN4BEG[8] ,
    \Tile_X3Y4_NN4BEG[7] ,
    \Tile_X3Y4_NN4BEG[6] ,
    \Tile_X3Y4_NN4BEG[5] ,
    \Tile_X3Y4_NN4BEG[4] ,
    \Tile_X3Y4_NN4BEG[3] ,
    \Tile_X3Y4_NN4BEG[2] ,
    \Tile_X3Y4_NN4BEG[1] ,
    \Tile_X3Y4_NN4BEG[0] }),
    .NN4END({\Tile_X3Y5_NN4BEG[15] ,
    \Tile_X3Y5_NN4BEG[14] ,
    \Tile_X3Y5_NN4BEG[13] ,
    \Tile_X3Y5_NN4BEG[12] ,
    \Tile_X3Y5_NN4BEG[11] ,
    \Tile_X3Y5_NN4BEG[10] ,
    \Tile_X3Y5_NN4BEG[9] ,
    \Tile_X3Y5_NN4BEG[8] ,
    \Tile_X3Y5_NN4BEG[7] ,
    \Tile_X3Y5_NN4BEG[6] ,
    \Tile_X3Y5_NN4BEG[5] ,
    \Tile_X3Y5_NN4BEG[4] ,
    \Tile_X3Y5_NN4BEG[3] ,
    \Tile_X3Y5_NN4BEG[2] ,
    \Tile_X3Y5_NN4BEG[1] ,
    \Tile_X3Y5_NN4BEG[0] }),
    .S1BEG({\Tile_X3Y4_S1BEG[3] ,
    \Tile_X3Y4_S1BEG[2] ,
    \Tile_X3Y4_S1BEG[1] ,
    \Tile_X3Y4_S1BEG[0] }),
    .S1END({\Tile_X3Y3_S1BEG[3] ,
    \Tile_X3Y3_S1BEG[2] ,
    \Tile_X3Y3_S1BEG[1] ,
    \Tile_X3Y3_S1BEG[0] }),
    .S2BEG({\Tile_X3Y4_S2BEG[7] ,
    \Tile_X3Y4_S2BEG[6] ,
    \Tile_X3Y4_S2BEG[5] ,
    \Tile_X3Y4_S2BEG[4] ,
    \Tile_X3Y4_S2BEG[3] ,
    \Tile_X3Y4_S2BEG[2] ,
    \Tile_X3Y4_S2BEG[1] ,
    \Tile_X3Y4_S2BEG[0] }),
    .S2BEGb({\Tile_X3Y4_S2BEGb[7] ,
    \Tile_X3Y4_S2BEGb[6] ,
    \Tile_X3Y4_S2BEGb[5] ,
    \Tile_X3Y4_S2BEGb[4] ,
    \Tile_X3Y4_S2BEGb[3] ,
    \Tile_X3Y4_S2BEGb[2] ,
    \Tile_X3Y4_S2BEGb[1] ,
    \Tile_X3Y4_S2BEGb[0] }),
    .S2END({\Tile_X3Y3_S2BEGb[7] ,
    \Tile_X3Y3_S2BEGb[6] ,
    \Tile_X3Y3_S2BEGb[5] ,
    \Tile_X3Y3_S2BEGb[4] ,
    \Tile_X3Y3_S2BEGb[3] ,
    \Tile_X3Y3_S2BEGb[2] ,
    \Tile_X3Y3_S2BEGb[1] ,
    \Tile_X3Y3_S2BEGb[0] }),
    .S2MID({\Tile_X3Y3_S2BEG[7] ,
    \Tile_X3Y3_S2BEG[6] ,
    \Tile_X3Y3_S2BEG[5] ,
    \Tile_X3Y3_S2BEG[4] ,
    \Tile_X3Y3_S2BEG[3] ,
    \Tile_X3Y3_S2BEG[2] ,
    \Tile_X3Y3_S2BEG[1] ,
    \Tile_X3Y3_S2BEG[0] }),
    .S4BEG({\Tile_X3Y4_S4BEG[15] ,
    \Tile_X3Y4_S4BEG[14] ,
    \Tile_X3Y4_S4BEG[13] ,
    \Tile_X3Y4_S4BEG[12] ,
    \Tile_X3Y4_S4BEG[11] ,
    \Tile_X3Y4_S4BEG[10] ,
    \Tile_X3Y4_S4BEG[9] ,
    \Tile_X3Y4_S4BEG[8] ,
    \Tile_X3Y4_S4BEG[7] ,
    \Tile_X3Y4_S4BEG[6] ,
    \Tile_X3Y4_S4BEG[5] ,
    \Tile_X3Y4_S4BEG[4] ,
    \Tile_X3Y4_S4BEG[3] ,
    \Tile_X3Y4_S4BEG[2] ,
    \Tile_X3Y4_S4BEG[1] ,
    \Tile_X3Y4_S4BEG[0] }),
    .S4END({\Tile_X3Y3_S4BEG[15] ,
    \Tile_X3Y3_S4BEG[14] ,
    \Tile_X3Y3_S4BEG[13] ,
    \Tile_X3Y3_S4BEG[12] ,
    \Tile_X3Y3_S4BEG[11] ,
    \Tile_X3Y3_S4BEG[10] ,
    \Tile_X3Y3_S4BEG[9] ,
    \Tile_X3Y3_S4BEG[8] ,
    \Tile_X3Y3_S4BEG[7] ,
    \Tile_X3Y3_S4BEG[6] ,
    \Tile_X3Y3_S4BEG[5] ,
    \Tile_X3Y3_S4BEG[4] ,
    \Tile_X3Y3_S4BEG[3] ,
    \Tile_X3Y3_S4BEG[2] ,
    \Tile_X3Y3_S4BEG[1] ,
    \Tile_X3Y3_S4BEG[0] }),
    .SS4BEG({\Tile_X3Y4_SS4BEG[15] ,
    \Tile_X3Y4_SS4BEG[14] ,
    \Tile_X3Y4_SS4BEG[13] ,
    \Tile_X3Y4_SS4BEG[12] ,
    \Tile_X3Y4_SS4BEG[11] ,
    \Tile_X3Y4_SS4BEG[10] ,
    \Tile_X3Y4_SS4BEG[9] ,
    \Tile_X3Y4_SS4BEG[8] ,
    \Tile_X3Y4_SS4BEG[7] ,
    \Tile_X3Y4_SS4BEG[6] ,
    \Tile_X3Y4_SS4BEG[5] ,
    \Tile_X3Y4_SS4BEG[4] ,
    \Tile_X3Y4_SS4BEG[3] ,
    \Tile_X3Y4_SS4BEG[2] ,
    \Tile_X3Y4_SS4BEG[1] ,
    \Tile_X3Y4_SS4BEG[0] }),
    .SS4END({\Tile_X3Y3_SS4BEG[15] ,
    \Tile_X3Y3_SS4BEG[14] ,
    \Tile_X3Y3_SS4BEG[13] ,
    \Tile_X3Y3_SS4BEG[12] ,
    \Tile_X3Y3_SS4BEG[11] ,
    \Tile_X3Y3_SS4BEG[10] ,
    \Tile_X3Y3_SS4BEG[9] ,
    \Tile_X3Y3_SS4BEG[8] ,
    \Tile_X3Y3_SS4BEG[7] ,
    \Tile_X3Y3_SS4BEG[6] ,
    \Tile_X3Y3_SS4BEG[5] ,
    \Tile_X3Y3_SS4BEG[4] ,
    \Tile_X3Y3_SS4BEG[3] ,
    \Tile_X3Y3_SS4BEG[2] ,
    \Tile_X3Y3_SS4BEG[1] ,
    \Tile_X3Y3_SS4BEG[0] }),
    .W1BEG({\Tile_X3Y4_W1BEG[3] ,
    \Tile_X3Y4_W1BEG[2] ,
    \Tile_X3Y4_W1BEG[1] ,
    \Tile_X3Y4_W1BEG[0] }),
    .W1END({\Tile_X4Y4_W1BEG[3] ,
    \Tile_X4Y4_W1BEG[2] ,
    \Tile_X4Y4_W1BEG[1] ,
    \Tile_X4Y4_W1BEG[0] }),
    .W2BEG({\Tile_X3Y4_W2BEG[7] ,
    \Tile_X3Y4_W2BEG[6] ,
    \Tile_X3Y4_W2BEG[5] ,
    \Tile_X3Y4_W2BEG[4] ,
    \Tile_X3Y4_W2BEG[3] ,
    \Tile_X3Y4_W2BEG[2] ,
    \Tile_X3Y4_W2BEG[1] ,
    \Tile_X3Y4_W2BEG[0] }),
    .W2BEGb({\Tile_X3Y4_W2BEGb[7] ,
    \Tile_X3Y4_W2BEGb[6] ,
    \Tile_X3Y4_W2BEGb[5] ,
    \Tile_X3Y4_W2BEGb[4] ,
    \Tile_X3Y4_W2BEGb[3] ,
    \Tile_X3Y4_W2BEGb[2] ,
    \Tile_X3Y4_W2BEGb[1] ,
    \Tile_X3Y4_W2BEGb[0] }),
    .W2END({\Tile_X4Y4_W2BEGb[7] ,
    \Tile_X4Y4_W2BEGb[6] ,
    \Tile_X4Y4_W2BEGb[5] ,
    \Tile_X4Y4_W2BEGb[4] ,
    \Tile_X4Y4_W2BEGb[3] ,
    \Tile_X4Y4_W2BEGb[2] ,
    \Tile_X4Y4_W2BEGb[1] ,
    \Tile_X4Y4_W2BEGb[0] }),
    .W2MID({\Tile_X4Y4_W2BEG[7] ,
    \Tile_X4Y4_W2BEG[6] ,
    \Tile_X4Y4_W2BEG[5] ,
    \Tile_X4Y4_W2BEG[4] ,
    \Tile_X4Y4_W2BEG[3] ,
    \Tile_X4Y4_W2BEG[2] ,
    \Tile_X4Y4_W2BEG[1] ,
    \Tile_X4Y4_W2BEG[0] }),
    .W6BEG({\Tile_X3Y4_W6BEG[11] ,
    \Tile_X3Y4_W6BEG[10] ,
    \Tile_X3Y4_W6BEG[9] ,
    \Tile_X3Y4_W6BEG[8] ,
    \Tile_X3Y4_W6BEG[7] ,
    \Tile_X3Y4_W6BEG[6] ,
    \Tile_X3Y4_W6BEG[5] ,
    \Tile_X3Y4_W6BEG[4] ,
    \Tile_X3Y4_W6BEG[3] ,
    \Tile_X3Y4_W6BEG[2] ,
    \Tile_X3Y4_W6BEG[1] ,
    \Tile_X3Y4_W6BEG[0] }),
    .W6END({\Tile_X4Y4_W6BEG[11] ,
    \Tile_X4Y4_W6BEG[10] ,
    \Tile_X4Y4_W6BEG[9] ,
    \Tile_X4Y4_W6BEG[8] ,
    \Tile_X4Y4_W6BEG[7] ,
    \Tile_X4Y4_W6BEG[6] ,
    \Tile_X4Y4_W6BEG[5] ,
    \Tile_X4Y4_W6BEG[4] ,
    \Tile_X4Y4_W6BEG[3] ,
    \Tile_X4Y4_W6BEG[2] ,
    \Tile_X4Y4_W6BEG[1] ,
    \Tile_X4Y4_W6BEG[0] }),
    .WW4BEG({\Tile_X3Y4_WW4BEG[15] ,
    \Tile_X3Y4_WW4BEG[14] ,
    \Tile_X3Y4_WW4BEG[13] ,
    \Tile_X3Y4_WW4BEG[12] ,
    \Tile_X3Y4_WW4BEG[11] ,
    \Tile_X3Y4_WW4BEG[10] ,
    \Tile_X3Y4_WW4BEG[9] ,
    \Tile_X3Y4_WW4BEG[8] ,
    \Tile_X3Y4_WW4BEG[7] ,
    \Tile_X3Y4_WW4BEG[6] ,
    \Tile_X3Y4_WW4BEG[5] ,
    \Tile_X3Y4_WW4BEG[4] ,
    \Tile_X3Y4_WW4BEG[3] ,
    \Tile_X3Y4_WW4BEG[2] ,
    \Tile_X3Y4_WW4BEG[1] ,
    \Tile_X3Y4_WW4BEG[0] }),
    .WW4END({\Tile_X4Y4_WW4BEG[15] ,
    \Tile_X4Y4_WW4BEG[14] ,
    \Tile_X4Y4_WW4BEG[13] ,
    \Tile_X4Y4_WW4BEG[12] ,
    \Tile_X4Y4_WW4BEG[11] ,
    \Tile_X4Y4_WW4BEG[10] ,
    \Tile_X4Y4_WW4BEG[9] ,
    \Tile_X4Y4_WW4BEG[8] ,
    \Tile_X4Y4_WW4BEG[7] ,
    \Tile_X4Y4_WW4BEG[6] ,
    \Tile_X4Y4_WW4BEG[5] ,
    \Tile_X4Y4_WW4BEG[4] ,
    \Tile_X4Y4_WW4BEG[3] ,
    \Tile_X4Y4_WW4BEG[2] ,
    \Tile_X4Y4_WW4BEG[1] ,
    \Tile_X4Y4_WW4BEG[0] }));
 LUT4AB Tile_X3Y5_LUT4AB (.Ci(Tile_X3Y6_Co),
    .Co(Tile_X3Y5_Co),
    .UserCLK(Tile_X3Y6_UserCLKo),
    .UserCLKo(Tile_X3Y5_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X3Y5_E1BEG[3] ,
    \Tile_X3Y5_E1BEG[2] ,
    \Tile_X3Y5_E1BEG[1] ,
    \Tile_X3Y5_E1BEG[0] }),
    .E1END({\Tile_X2Y5_E1BEG[3] ,
    \Tile_X2Y5_E1BEG[2] ,
    \Tile_X2Y5_E1BEG[1] ,
    \Tile_X2Y5_E1BEG[0] }),
    .E2BEG({\Tile_X3Y5_E2BEG[7] ,
    \Tile_X3Y5_E2BEG[6] ,
    \Tile_X3Y5_E2BEG[5] ,
    \Tile_X3Y5_E2BEG[4] ,
    \Tile_X3Y5_E2BEG[3] ,
    \Tile_X3Y5_E2BEG[2] ,
    \Tile_X3Y5_E2BEG[1] ,
    \Tile_X3Y5_E2BEG[0] }),
    .E2BEGb({\Tile_X3Y5_E2BEGb[7] ,
    \Tile_X3Y5_E2BEGb[6] ,
    \Tile_X3Y5_E2BEGb[5] ,
    \Tile_X3Y5_E2BEGb[4] ,
    \Tile_X3Y5_E2BEGb[3] ,
    \Tile_X3Y5_E2BEGb[2] ,
    \Tile_X3Y5_E2BEGb[1] ,
    \Tile_X3Y5_E2BEGb[0] }),
    .E2END({\Tile_X2Y5_E2BEGb[7] ,
    \Tile_X2Y5_E2BEGb[6] ,
    \Tile_X2Y5_E2BEGb[5] ,
    \Tile_X2Y5_E2BEGb[4] ,
    \Tile_X2Y5_E2BEGb[3] ,
    \Tile_X2Y5_E2BEGb[2] ,
    \Tile_X2Y5_E2BEGb[1] ,
    \Tile_X2Y5_E2BEGb[0] }),
    .E2MID({\Tile_X2Y5_E2BEG[7] ,
    \Tile_X2Y5_E2BEG[6] ,
    \Tile_X2Y5_E2BEG[5] ,
    \Tile_X2Y5_E2BEG[4] ,
    \Tile_X2Y5_E2BEG[3] ,
    \Tile_X2Y5_E2BEG[2] ,
    \Tile_X2Y5_E2BEG[1] ,
    \Tile_X2Y5_E2BEG[0] }),
    .E6BEG({\Tile_X3Y5_E6BEG[11] ,
    \Tile_X3Y5_E6BEG[10] ,
    \Tile_X3Y5_E6BEG[9] ,
    \Tile_X3Y5_E6BEG[8] ,
    \Tile_X3Y5_E6BEG[7] ,
    \Tile_X3Y5_E6BEG[6] ,
    \Tile_X3Y5_E6BEG[5] ,
    \Tile_X3Y5_E6BEG[4] ,
    \Tile_X3Y5_E6BEG[3] ,
    \Tile_X3Y5_E6BEG[2] ,
    \Tile_X3Y5_E6BEG[1] ,
    \Tile_X3Y5_E6BEG[0] }),
    .E6END({\Tile_X2Y5_E6BEG[11] ,
    \Tile_X2Y5_E6BEG[10] ,
    \Tile_X2Y5_E6BEG[9] ,
    \Tile_X2Y5_E6BEG[8] ,
    \Tile_X2Y5_E6BEG[7] ,
    \Tile_X2Y5_E6BEG[6] ,
    \Tile_X2Y5_E6BEG[5] ,
    \Tile_X2Y5_E6BEG[4] ,
    \Tile_X2Y5_E6BEG[3] ,
    \Tile_X2Y5_E6BEG[2] ,
    \Tile_X2Y5_E6BEG[1] ,
    \Tile_X2Y5_E6BEG[0] }),
    .EE4BEG({\Tile_X3Y5_EE4BEG[15] ,
    \Tile_X3Y5_EE4BEG[14] ,
    \Tile_X3Y5_EE4BEG[13] ,
    \Tile_X3Y5_EE4BEG[12] ,
    \Tile_X3Y5_EE4BEG[11] ,
    \Tile_X3Y5_EE4BEG[10] ,
    \Tile_X3Y5_EE4BEG[9] ,
    \Tile_X3Y5_EE4BEG[8] ,
    \Tile_X3Y5_EE4BEG[7] ,
    \Tile_X3Y5_EE4BEG[6] ,
    \Tile_X3Y5_EE4BEG[5] ,
    \Tile_X3Y5_EE4BEG[4] ,
    \Tile_X3Y5_EE4BEG[3] ,
    \Tile_X3Y5_EE4BEG[2] ,
    \Tile_X3Y5_EE4BEG[1] ,
    \Tile_X3Y5_EE4BEG[0] }),
    .EE4END({\Tile_X2Y5_EE4BEG[15] ,
    \Tile_X2Y5_EE4BEG[14] ,
    \Tile_X2Y5_EE4BEG[13] ,
    \Tile_X2Y5_EE4BEG[12] ,
    \Tile_X2Y5_EE4BEG[11] ,
    \Tile_X2Y5_EE4BEG[10] ,
    \Tile_X2Y5_EE4BEG[9] ,
    \Tile_X2Y5_EE4BEG[8] ,
    \Tile_X2Y5_EE4BEG[7] ,
    \Tile_X2Y5_EE4BEG[6] ,
    \Tile_X2Y5_EE4BEG[5] ,
    \Tile_X2Y5_EE4BEG[4] ,
    \Tile_X2Y5_EE4BEG[3] ,
    \Tile_X2Y5_EE4BEG[2] ,
    \Tile_X2Y5_EE4BEG[1] ,
    \Tile_X2Y5_EE4BEG[0] }),
    .FrameData({\Tile_X2Y5_FrameData_O[31] ,
    \Tile_X2Y5_FrameData_O[30] ,
    \Tile_X2Y5_FrameData_O[29] ,
    \Tile_X2Y5_FrameData_O[28] ,
    \Tile_X2Y5_FrameData_O[27] ,
    \Tile_X2Y5_FrameData_O[26] ,
    \Tile_X2Y5_FrameData_O[25] ,
    \Tile_X2Y5_FrameData_O[24] ,
    \Tile_X2Y5_FrameData_O[23] ,
    \Tile_X2Y5_FrameData_O[22] ,
    \Tile_X2Y5_FrameData_O[21] ,
    \Tile_X2Y5_FrameData_O[20] ,
    \Tile_X2Y5_FrameData_O[19] ,
    \Tile_X2Y5_FrameData_O[18] ,
    \Tile_X2Y5_FrameData_O[17] ,
    \Tile_X2Y5_FrameData_O[16] ,
    \Tile_X2Y5_FrameData_O[15] ,
    \Tile_X2Y5_FrameData_O[14] ,
    \Tile_X2Y5_FrameData_O[13] ,
    \Tile_X2Y5_FrameData_O[12] ,
    \Tile_X2Y5_FrameData_O[11] ,
    \Tile_X2Y5_FrameData_O[10] ,
    \Tile_X2Y5_FrameData_O[9] ,
    \Tile_X2Y5_FrameData_O[8] ,
    \Tile_X2Y5_FrameData_O[7] ,
    \Tile_X2Y5_FrameData_O[6] ,
    \Tile_X2Y5_FrameData_O[5] ,
    \Tile_X2Y5_FrameData_O[4] ,
    \Tile_X2Y5_FrameData_O[3] ,
    \Tile_X2Y5_FrameData_O[2] ,
    \Tile_X2Y5_FrameData_O[1] ,
    \Tile_X2Y5_FrameData_O[0] }),
    .FrameData_O({\Tile_X3Y5_FrameData_O[31] ,
    \Tile_X3Y5_FrameData_O[30] ,
    \Tile_X3Y5_FrameData_O[29] ,
    \Tile_X3Y5_FrameData_O[28] ,
    \Tile_X3Y5_FrameData_O[27] ,
    \Tile_X3Y5_FrameData_O[26] ,
    \Tile_X3Y5_FrameData_O[25] ,
    \Tile_X3Y5_FrameData_O[24] ,
    \Tile_X3Y5_FrameData_O[23] ,
    \Tile_X3Y5_FrameData_O[22] ,
    \Tile_X3Y5_FrameData_O[21] ,
    \Tile_X3Y5_FrameData_O[20] ,
    \Tile_X3Y5_FrameData_O[19] ,
    \Tile_X3Y5_FrameData_O[18] ,
    \Tile_X3Y5_FrameData_O[17] ,
    \Tile_X3Y5_FrameData_O[16] ,
    \Tile_X3Y5_FrameData_O[15] ,
    \Tile_X3Y5_FrameData_O[14] ,
    \Tile_X3Y5_FrameData_O[13] ,
    \Tile_X3Y5_FrameData_O[12] ,
    \Tile_X3Y5_FrameData_O[11] ,
    \Tile_X3Y5_FrameData_O[10] ,
    \Tile_X3Y5_FrameData_O[9] ,
    \Tile_X3Y5_FrameData_O[8] ,
    \Tile_X3Y5_FrameData_O[7] ,
    \Tile_X3Y5_FrameData_O[6] ,
    \Tile_X3Y5_FrameData_O[5] ,
    \Tile_X3Y5_FrameData_O[4] ,
    \Tile_X3Y5_FrameData_O[3] ,
    \Tile_X3Y5_FrameData_O[2] ,
    \Tile_X3Y5_FrameData_O[1] ,
    \Tile_X3Y5_FrameData_O[0] }),
    .FrameStrobe({\Tile_X3Y6_FrameStrobe_O[19] ,
    \Tile_X3Y6_FrameStrobe_O[18] ,
    \Tile_X3Y6_FrameStrobe_O[17] ,
    \Tile_X3Y6_FrameStrobe_O[16] ,
    \Tile_X3Y6_FrameStrobe_O[15] ,
    \Tile_X3Y6_FrameStrobe_O[14] ,
    \Tile_X3Y6_FrameStrobe_O[13] ,
    \Tile_X3Y6_FrameStrobe_O[12] ,
    \Tile_X3Y6_FrameStrobe_O[11] ,
    \Tile_X3Y6_FrameStrobe_O[10] ,
    \Tile_X3Y6_FrameStrobe_O[9] ,
    \Tile_X3Y6_FrameStrobe_O[8] ,
    \Tile_X3Y6_FrameStrobe_O[7] ,
    \Tile_X3Y6_FrameStrobe_O[6] ,
    \Tile_X3Y6_FrameStrobe_O[5] ,
    \Tile_X3Y6_FrameStrobe_O[4] ,
    \Tile_X3Y6_FrameStrobe_O[3] ,
    \Tile_X3Y6_FrameStrobe_O[2] ,
    \Tile_X3Y6_FrameStrobe_O[1] ,
    \Tile_X3Y6_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X3Y5_FrameStrobe_O[19] ,
    \Tile_X3Y5_FrameStrobe_O[18] ,
    \Tile_X3Y5_FrameStrobe_O[17] ,
    \Tile_X3Y5_FrameStrobe_O[16] ,
    \Tile_X3Y5_FrameStrobe_O[15] ,
    \Tile_X3Y5_FrameStrobe_O[14] ,
    \Tile_X3Y5_FrameStrobe_O[13] ,
    \Tile_X3Y5_FrameStrobe_O[12] ,
    \Tile_X3Y5_FrameStrobe_O[11] ,
    \Tile_X3Y5_FrameStrobe_O[10] ,
    \Tile_X3Y5_FrameStrobe_O[9] ,
    \Tile_X3Y5_FrameStrobe_O[8] ,
    \Tile_X3Y5_FrameStrobe_O[7] ,
    \Tile_X3Y5_FrameStrobe_O[6] ,
    \Tile_X3Y5_FrameStrobe_O[5] ,
    \Tile_X3Y5_FrameStrobe_O[4] ,
    \Tile_X3Y5_FrameStrobe_O[3] ,
    \Tile_X3Y5_FrameStrobe_O[2] ,
    \Tile_X3Y5_FrameStrobe_O[1] ,
    \Tile_X3Y5_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X3Y5_N1BEG[3] ,
    \Tile_X3Y5_N1BEG[2] ,
    \Tile_X3Y5_N1BEG[1] ,
    \Tile_X3Y5_N1BEG[0] }),
    .N1END({\Tile_X3Y6_N1BEG[3] ,
    \Tile_X3Y6_N1BEG[2] ,
    \Tile_X3Y6_N1BEG[1] ,
    \Tile_X3Y6_N1BEG[0] }),
    .N2BEG({\Tile_X3Y5_N2BEG[7] ,
    \Tile_X3Y5_N2BEG[6] ,
    \Tile_X3Y5_N2BEG[5] ,
    \Tile_X3Y5_N2BEG[4] ,
    \Tile_X3Y5_N2BEG[3] ,
    \Tile_X3Y5_N2BEG[2] ,
    \Tile_X3Y5_N2BEG[1] ,
    \Tile_X3Y5_N2BEG[0] }),
    .N2BEGb({\Tile_X3Y5_N2BEGb[7] ,
    \Tile_X3Y5_N2BEGb[6] ,
    \Tile_X3Y5_N2BEGb[5] ,
    \Tile_X3Y5_N2BEGb[4] ,
    \Tile_X3Y5_N2BEGb[3] ,
    \Tile_X3Y5_N2BEGb[2] ,
    \Tile_X3Y5_N2BEGb[1] ,
    \Tile_X3Y5_N2BEGb[0] }),
    .N2END({\Tile_X3Y6_N2BEGb[7] ,
    \Tile_X3Y6_N2BEGb[6] ,
    \Tile_X3Y6_N2BEGb[5] ,
    \Tile_X3Y6_N2BEGb[4] ,
    \Tile_X3Y6_N2BEGb[3] ,
    \Tile_X3Y6_N2BEGb[2] ,
    \Tile_X3Y6_N2BEGb[1] ,
    \Tile_X3Y6_N2BEGb[0] }),
    .N2MID({\Tile_X3Y6_N2BEG[7] ,
    \Tile_X3Y6_N2BEG[6] ,
    \Tile_X3Y6_N2BEG[5] ,
    \Tile_X3Y6_N2BEG[4] ,
    \Tile_X3Y6_N2BEG[3] ,
    \Tile_X3Y6_N2BEG[2] ,
    \Tile_X3Y6_N2BEG[1] ,
    \Tile_X3Y6_N2BEG[0] }),
    .N4BEG({\Tile_X3Y5_N4BEG[15] ,
    \Tile_X3Y5_N4BEG[14] ,
    \Tile_X3Y5_N4BEG[13] ,
    \Tile_X3Y5_N4BEG[12] ,
    \Tile_X3Y5_N4BEG[11] ,
    \Tile_X3Y5_N4BEG[10] ,
    \Tile_X3Y5_N4BEG[9] ,
    \Tile_X3Y5_N4BEG[8] ,
    \Tile_X3Y5_N4BEG[7] ,
    \Tile_X3Y5_N4BEG[6] ,
    \Tile_X3Y5_N4BEG[5] ,
    \Tile_X3Y5_N4BEG[4] ,
    \Tile_X3Y5_N4BEG[3] ,
    \Tile_X3Y5_N4BEG[2] ,
    \Tile_X3Y5_N4BEG[1] ,
    \Tile_X3Y5_N4BEG[0] }),
    .N4END({\Tile_X3Y6_N4BEG[15] ,
    \Tile_X3Y6_N4BEG[14] ,
    \Tile_X3Y6_N4BEG[13] ,
    \Tile_X3Y6_N4BEG[12] ,
    \Tile_X3Y6_N4BEG[11] ,
    \Tile_X3Y6_N4BEG[10] ,
    \Tile_X3Y6_N4BEG[9] ,
    \Tile_X3Y6_N4BEG[8] ,
    \Tile_X3Y6_N4BEG[7] ,
    \Tile_X3Y6_N4BEG[6] ,
    \Tile_X3Y6_N4BEG[5] ,
    \Tile_X3Y6_N4BEG[4] ,
    \Tile_X3Y6_N4BEG[3] ,
    \Tile_X3Y6_N4BEG[2] ,
    \Tile_X3Y6_N4BEG[1] ,
    \Tile_X3Y6_N4BEG[0] }),
    .NN4BEG({\Tile_X3Y5_NN4BEG[15] ,
    \Tile_X3Y5_NN4BEG[14] ,
    \Tile_X3Y5_NN4BEG[13] ,
    \Tile_X3Y5_NN4BEG[12] ,
    \Tile_X3Y5_NN4BEG[11] ,
    \Tile_X3Y5_NN4BEG[10] ,
    \Tile_X3Y5_NN4BEG[9] ,
    \Tile_X3Y5_NN4BEG[8] ,
    \Tile_X3Y5_NN4BEG[7] ,
    \Tile_X3Y5_NN4BEG[6] ,
    \Tile_X3Y5_NN4BEG[5] ,
    \Tile_X3Y5_NN4BEG[4] ,
    \Tile_X3Y5_NN4BEG[3] ,
    \Tile_X3Y5_NN4BEG[2] ,
    \Tile_X3Y5_NN4BEG[1] ,
    \Tile_X3Y5_NN4BEG[0] }),
    .NN4END({\Tile_X3Y6_NN4BEG[15] ,
    \Tile_X3Y6_NN4BEG[14] ,
    \Tile_X3Y6_NN4BEG[13] ,
    \Tile_X3Y6_NN4BEG[12] ,
    \Tile_X3Y6_NN4BEG[11] ,
    \Tile_X3Y6_NN4BEG[10] ,
    \Tile_X3Y6_NN4BEG[9] ,
    \Tile_X3Y6_NN4BEG[8] ,
    \Tile_X3Y6_NN4BEG[7] ,
    \Tile_X3Y6_NN4BEG[6] ,
    \Tile_X3Y6_NN4BEG[5] ,
    \Tile_X3Y6_NN4BEG[4] ,
    \Tile_X3Y6_NN4BEG[3] ,
    \Tile_X3Y6_NN4BEG[2] ,
    \Tile_X3Y6_NN4BEG[1] ,
    \Tile_X3Y6_NN4BEG[0] }),
    .S1BEG({\Tile_X3Y5_S1BEG[3] ,
    \Tile_X3Y5_S1BEG[2] ,
    \Tile_X3Y5_S1BEG[1] ,
    \Tile_X3Y5_S1BEG[0] }),
    .S1END({\Tile_X3Y4_S1BEG[3] ,
    \Tile_X3Y4_S1BEG[2] ,
    \Tile_X3Y4_S1BEG[1] ,
    \Tile_X3Y4_S1BEG[0] }),
    .S2BEG({\Tile_X3Y5_S2BEG[7] ,
    \Tile_X3Y5_S2BEG[6] ,
    \Tile_X3Y5_S2BEG[5] ,
    \Tile_X3Y5_S2BEG[4] ,
    \Tile_X3Y5_S2BEG[3] ,
    \Tile_X3Y5_S2BEG[2] ,
    \Tile_X3Y5_S2BEG[1] ,
    \Tile_X3Y5_S2BEG[0] }),
    .S2BEGb({\Tile_X3Y5_S2BEGb[7] ,
    \Tile_X3Y5_S2BEGb[6] ,
    \Tile_X3Y5_S2BEGb[5] ,
    \Tile_X3Y5_S2BEGb[4] ,
    \Tile_X3Y5_S2BEGb[3] ,
    \Tile_X3Y5_S2BEGb[2] ,
    \Tile_X3Y5_S2BEGb[1] ,
    \Tile_X3Y5_S2BEGb[0] }),
    .S2END({\Tile_X3Y4_S2BEGb[7] ,
    \Tile_X3Y4_S2BEGb[6] ,
    \Tile_X3Y4_S2BEGb[5] ,
    \Tile_X3Y4_S2BEGb[4] ,
    \Tile_X3Y4_S2BEGb[3] ,
    \Tile_X3Y4_S2BEGb[2] ,
    \Tile_X3Y4_S2BEGb[1] ,
    \Tile_X3Y4_S2BEGb[0] }),
    .S2MID({\Tile_X3Y4_S2BEG[7] ,
    \Tile_X3Y4_S2BEG[6] ,
    \Tile_X3Y4_S2BEG[5] ,
    \Tile_X3Y4_S2BEG[4] ,
    \Tile_X3Y4_S2BEG[3] ,
    \Tile_X3Y4_S2BEG[2] ,
    \Tile_X3Y4_S2BEG[1] ,
    \Tile_X3Y4_S2BEG[0] }),
    .S4BEG({\Tile_X3Y5_S4BEG[15] ,
    \Tile_X3Y5_S4BEG[14] ,
    \Tile_X3Y5_S4BEG[13] ,
    \Tile_X3Y5_S4BEG[12] ,
    \Tile_X3Y5_S4BEG[11] ,
    \Tile_X3Y5_S4BEG[10] ,
    \Tile_X3Y5_S4BEG[9] ,
    \Tile_X3Y5_S4BEG[8] ,
    \Tile_X3Y5_S4BEG[7] ,
    \Tile_X3Y5_S4BEG[6] ,
    \Tile_X3Y5_S4BEG[5] ,
    \Tile_X3Y5_S4BEG[4] ,
    \Tile_X3Y5_S4BEG[3] ,
    \Tile_X3Y5_S4BEG[2] ,
    \Tile_X3Y5_S4BEG[1] ,
    \Tile_X3Y5_S4BEG[0] }),
    .S4END({\Tile_X3Y4_S4BEG[15] ,
    \Tile_X3Y4_S4BEG[14] ,
    \Tile_X3Y4_S4BEG[13] ,
    \Tile_X3Y4_S4BEG[12] ,
    \Tile_X3Y4_S4BEG[11] ,
    \Tile_X3Y4_S4BEG[10] ,
    \Tile_X3Y4_S4BEG[9] ,
    \Tile_X3Y4_S4BEG[8] ,
    \Tile_X3Y4_S4BEG[7] ,
    \Tile_X3Y4_S4BEG[6] ,
    \Tile_X3Y4_S4BEG[5] ,
    \Tile_X3Y4_S4BEG[4] ,
    \Tile_X3Y4_S4BEG[3] ,
    \Tile_X3Y4_S4BEG[2] ,
    \Tile_X3Y4_S4BEG[1] ,
    \Tile_X3Y4_S4BEG[0] }),
    .SS4BEG({\Tile_X3Y5_SS4BEG[15] ,
    \Tile_X3Y5_SS4BEG[14] ,
    \Tile_X3Y5_SS4BEG[13] ,
    \Tile_X3Y5_SS4BEG[12] ,
    \Tile_X3Y5_SS4BEG[11] ,
    \Tile_X3Y5_SS4BEG[10] ,
    \Tile_X3Y5_SS4BEG[9] ,
    \Tile_X3Y5_SS4BEG[8] ,
    \Tile_X3Y5_SS4BEG[7] ,
    \Tile_X3Y5_SS4BEG[6] ,
    \Tile_X3Y5_SS4BEG[5] ,
    \Tile_X3Y5_SS4BEG[4] ,
    \Tile_X3Y5_SS4BEG[3] ,
    \Tile_X3Y5_SS4BEG[2] ,
    \Tile_X3Y5_SS4BEG[1] ,
    \Tile_X3Y5_SS4BEG[0] }),
    .SS4END({\Tile_X3Y4_SS4BEG[15] ,
    \Tile_X3Y4_SS4BEG[14] ,
    \Tile_X3Y4_SS4BEG[13] ,
    \Tile_X3Y4_SS4BEG[12] ,
    \Tile_X3Y4_SS4BEG[11] ,
    \Tile_X3Y4_SS4BEG[10] ,
    \Tile_X3Y4_SS4BEG[9] ,
    \Tile_X3Y4_SS4BEG[8] ,
    \Tile_X3Y4_SS4BEG[7] ,
    \Tile_X3Y4_SS4BEG[6] ,
    \Tile_X3Y4_SS4BEG[5] ,
    \Tile_X3Y4_SS4BEG[4] ,
    \Tile_X3Y4_SS4BEG[3] ,
    \Tile_X3Y4_SS4BEG[2] ,
    \Tile_X3Y4_SS4BEG[1] ,
    \Tile_X3Y4_SS4BEG[0] }),
    .W1BEG({\Tile_X3Y5_W1BEG[3] ,
    \Tile_X3Y5_W1BEG[2] ,
    \Tile_X3Y5_W1BEG[1] ,
    \Tile_X3Y5_W1BEG[0] }),
    .W1END({\Tile_X4Y5_W1BEG[3] ,
    \Tile_X4Y5_W1BEG[2] ,
    \Tile_X4Y5_W1BEG[1] ,
    \Tile_X4Y5_W1BEG[0] }),
    .W2BEG({\Tile_X3Y5_W2BEG[7] ,
    \Tile_X3Y5_W2BEG[6] ,
    \Tile_X3Y5_W2BEG[5] ,
    \Tile_X3Y5_W2BEG[4] ,
    \Tile_X3Y5_W2BEG[3] ,
    \Tile_X3Y5_W2BEG[2] ,
    \Tile_X3Y5_W2BEG[1] ,
    \Tile_X3Y5_W2BEG[0] }),
    .W2BEGb({\Tile_X3Y5_W2BEGb[7] ,
    \Tile_X3Y5_W2BEGb[6] ,
    \Tile_X3Y5_W2BEGb[5] ,
    \Tile_X3Y5_W2BEGb[4] ,
    \Tile_X3Y5_W2BEGb[3] ,
    \Tile_X3Y5_W2BEGb[2] ,
    \Tile_X3Y5_W2BEGb[1] ,
    \Tile_X3Y5_W2BEGb[0] }),
    .W2END({\Tile_X4Y5_W2BEGb[7] ,
    \Tile_X4Y5_W2BEGb[6] ,
    \Tile_X4Y5_W2BEGb[5] ,
    \Tile_X4Y5_W2BEGb[4] ,
    \Tile_X4Y5_W2BEGb[3] ,
    \Tile_X4Y5_W2BEGb[2] ,
    \Tile_X4Y5_W2BEGb[1] ,
    \Tile_X4Y5_W2BEGb[0] }),
    .W2MID({\Tile_X4Y5_W2BEG[7] ,
    \Tile_X4Y5_W2BEG[6] ,
    \Tile_X4Y5_W2BEG[5] ,
    \Tile_X4Y5_W2BEG[4] ,
    \Tile_X4Y5_W2BEG[3] ,
    \Tile_X4Y5_W2BEG[2] ,
    \Tile_X4Y5_W2BEG[1] ,
    \Tile_X4Y5_W2BEG[0] }),
    .W6BEG({\Tile_X3Y5_W6BEG[11] ,
    \Tile_X3Y5_W6BEG[10] ,
    \Tile_X3Y5_W6BEG[9] ,
    \Tile_X3Y5_W6BEG[8] ,
    \Tile_X3Y5_W6BEG[7] ,
    \Tile_X3Y5_W6BEG[6] ,
    \Tile_X3Y5_W6BEG[5] ,
    \Tile_X3Y5_W6BEG[4] ,
    \Tile_X3Y5_W6BEG[3] ,
    \Tile_X3Y5_W6BEG[2] ,
    \Tile_X3Y5_W6BEG[1] ,
    \Tile_X3Y5_W6BEG[0] }),
    .W6END({\Tile_X4Y5_W6BEG[11] ,
    \Tile_X4Y5_W6BEG[10] ,
    \Tile_X4Y5_W6BEG[9] ,
    \Tile_X4Y5_W6BEG[8] ,
    \Tile_X4Y5_W6BEG[7] ,
    \Tile_X4Y5_W6BEG[6] ,
    \Tile_X4Y5_W6BEG[5] ,
    \Tile_X4Y5_W6BEG[4] ,
    \Tile_X4Y5_W6BEG[3] ,
    \Tile_X4Y5_W6BEG[2] ,
    \Tile_X4Y5_W6BEG[1] ,
    \Tile_X4Y5_W6BEG[0] }),
    .WW4BEG({\Tile_X3Y5_WW4BEG[15] ,
    \Tile_X3Y5_WW4BEG[14] ,
    \Tile_X3Y5_WW4BEG[13] ,
    \Tile_X3Y5_WW4BEG[12] ,
    \Tile_X3Y5_WW4BEG[11] ,
    \Tile_X3Y5_WW4BEG[10] ,
    \Tile_X3Y5_WW4BEG[9] ,
    \Tile_X3Y5_WW4BEG[8] ,
    \Tile_X3Y5_WW4BEG[7] ,
    \Tile_X3Y5_WW4BEG[6] ,
    \Tile_X3Y5_WW4BEG[5] ,
    \Tile_X3Y5_WW4BEG[4] ,
    \Tile_X3Y5_WW4BEG[3] ,
    \Tile_X3Y5_WW4BEG[2] ,
    \Tile_X3Y5_WW4BEG[1] ,
    \Tile_X3Y5_WW4BEG[0] }),
    .WW4END({\Tile_X4Y5_WW4BEG[15] ,
    \Tile_X4Y5_WW4BEG[14] ,
    \Tile_X4Y5_WW4BEG[13] ,
    \Tile_X4Y5_WW4BEG[12] ,
    \Tile_X4Y5_WW4BEG[11] ,
    \Tile_X4Y5_WW4BEG[10] ,
    \Tile_X4Y5_WW4BEG[9] ,
    \Tile_X4Y5_WW4BEG[8] ,
    \Tile_X4Y5_WW4BEG[7] ,
    \Tile_X4Y5_WW4BEG[6] ,
    \Tile_X4Y5_WW4BEG[5] ,
    \Tile_X4Y5_WW4BEG[4] ,
    \Tile_X4Y5_WW4BEG[3] ,
    \Tile_X4Y5_WW4BEG[2] ,
    \Tile_X4Y5_WW4BEG[1] ,
    \Tile_X4Y5_WW4BEG[0] }));
 LUT4AB Tile_X3Y6_LUT4AB (.Ci(Tile_X3Y7_Co),
    .Co(Tile_X3Y6_Co),
    .UserCLK(Tile_X3Y7_UserCLKo),
    .UserCLKo(Tile_X3Y6_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X3Y6_E1BEG[3] ,
    \Tile_X3Y6_E1BEG[2] ,
    \Tile_X3Y6_E1BEG[1] ,
    \Tile_X3Y6_E1BEG[0] }),
    .E1END({\Tile_X2Y6_E1BEG[3] ,
    \Tile_X2Y6_E1BEG[2] ,
    \Tile_X2Y6_E1BEG[1] ,
    \Tile_X2Y6_E1BEG[0] }),
    .E2BEG({\Tile_X3Y6_E2BEG[7] ,
    \Tile_X3Y6_E2BEG[6] ,
    \Tile_X3Y6_E2BEG[5] ,
    \Tile_X3Y6_E2BEG[4] ,
    \Tile_X3Y6_E2BEG[3] ,
    \Tile_X3Y6_E2BEG[2] ,
    \Tile_X3Y6_E2BEG[1] ,
    \Tile_X3Y6_E2BEG[0] }),
    .E2BEGb({\Tile_X3Y6_E2BEGb[7] ,
    \Tile_X3Y6_E2BEGb[6] ,
    \Tile_X3Y6_E2BEGb[5] ,
    \Tile_X3Y6_E2BEGb[4] ,
    \Tile_X3Y6_E2BEGb[3] ,
    \Tile_X3Y6_E2BEGb[2] ,
    \Tile_X3Y6_E2BEGb[1] ,
    \Tile_X3Y6_E2BEGb[0] }),
    .E2END({\Tile_X2Y6_E2BEGb[7] ,
    \Tile_X2Y6_E2BEGb[6] ,
    \Tile_X2Y6_E2BEGb[5] ,
    \Tile_X2Y6_E2BEGb[4] ,
    \Tile_X2Y6_E2BEGb[3] ,
    \Tile_X2Y6_E2BEGb[2] ,
    \Tile_X2Y6_E2BEGb[1] ,
    \Tile_X2Y6_E2BEGb[0] }),
    .E2MID({\Tile_X2Y6_E2BEG[7] ,
    \Tile_X2Y6_E2BEG[6] ,
    \Tile_X2Y6_E2BEG[5] ,
    \Tile_X2Y6_E2BEG[4] ,
    \Tile_X2Y6_E2BEG[3] ,
    \Tile_X2Y6_E2BEG[2] ,
    \Tile_X2Y6_E2BEG[1] ,
    \Tile_X2Y6_E2BEG[0] }),
    .E6BEG({\Tile_X3Y6_E6BEG[11] ,
    \Tile_X3Y6_E6BEG[10] ,
    \Tile_X3Y6_E6BEG[9] ,
    \Tile_X3Y6_E6BEG[8] ,
    \Tile_X3Y6_E6BEG[7] ,
    \Tile_X3Y6_E6BEG[6] ,
    \Tile_X3Y6_E6BEG[5] ,
    \Tile_X3Y6_E6BEG[4] ,
    \Tile_X3Y6_E6BEG[3] ,
    \Tile_X3Y6_E6BEG[2] ,
    \Tile_X3Y6_E6BEG[1] ,
    \Tile_X3Y6_E6BEG[0] }),
    .E6END({\Tile_X2Y6_E6BEG[11] ,
    \Tile_X2Y6_E6BEG[10] ,
    \Tile_X2Y6_E6BEG[9] ,
    \Tile_X2Y6_E6BEG[8] ,
    \Tile_X2Y6_E6BEG[7] ,
    \Tile_X2Y6_E6BEG[6] ,
    \Tile_X2Y6_E6BEG[5] ,
    \Tile_X2Y6_E6BEG[4] ,
    \Tile_X2Y6_E6BEG[3] ,
    \Tile_X2Y6_E6BEG[2] ,
    \Tile_X2Y6_E6BEG[1] ,
    \Tile_X2Y6_E6BEG[0] }),
    .EE4BEG({\Tile_X3Y6_EE4BEG[15] ,
    \Tile_X3Y6_EE4BEG[14] ,
    \Tile_X3Y6_EE4BEG[13] ,
    \Tile_X3Y6_EE4BEG[12] ,
    \Tile_X3Y6_EE4BEG[11] ,
    \Tile_X3Y6_EE4BEG[10] ,
    \Tile_X3Y6_EE4BEG[9] ,
    \Tile_X3Y6_EE4BEG[8] ,
    \Tile_X3Y6_EE4BEG[7] ,
    \Tile_X3Y6_EE4BEG[6] ,
    \Tile_X3Y6_EE4BEG[5] ,
    \Tile_X3Y6_EE4BEG[4] ,
    \Tile_X3Y6_EE4BEG[3] ,
    \Tile_X3Y6_EE4BEG[2] ,
    \Tile_X3Y6_EE4BEG[1] ,
    \Tile_X3Y6_EE4BEG[0] }),
    .EE4END({\Tile_X2Y6_EE4BEG[15] ,
    \Tile_X2Y6_EE4BEG[14] ,
    \Tile_X2Y6_EE4BEG[13] ,
    \Tile_X2Y6_EE4BEG[12] ,
    \Tile_X2Y6_EE4BEG[11] ,
    \Tile_X2Y6_EE4BEG[10] ,
    \Tile_X2Y6_EE4BEG[9] ,
    \Tile_X2Y6_EE4BEG[8] ,
    \Tile_X2Y6_EE4BEG[7] ,
    \Tile_X2Y6_EE4BEG[6] ,
    \Tile_X2Y6_EE4BEG[5] ,
    \Tile_X2Y6_EE4BEG[4] ,
    \Tile_X2Y6_EE4BEG[3] ,
    \Tile_X2Y6_EE4BEG[2] ,
    \Tile_X2Y6_EE4BEG[1] ,
    \Tile_X2Y6_EE4BEG[0] }),
    .FrameData({\Tile_X2Y6_FrameData_O[31] ,
    \Tile_X2Y6_FrameData_O[30] ,
    \Tile_X2Y6_FrameData_O[29] ,
    \Tile_X2Y6_FrameData_O[28] ,
    \Tile_X2Y6_FrameData_O[27] ,
    \Tile_X2Y6_FrameData_O[26] ,
    \Tile_X2Y6_FrameData_O[25] ,
    \Tile_X2Y6_FrameData_O[24] ,
    \Tile_X2Y6_FrameData_O[23] ,
    \Tile_X2Y6_FrameData_O[22] ,
    \Tile_X2Y6_FrameData_O[21] ,
    \Tile_X2Y6_FrameData_O[20] ,
    \Tile_X2Y6_FrameData_O[19] ,
    \Tile_X2Y6_FrameData_O[18] ,
    \Tile_X2Y6_FrameData_O[17] ,
    \Tile_X2Y6_FrameData_O[16] ,
    \Tile_X2Y6_FrameData_O[15] ,
    \Tile_X2Y6_FrameData_O[14] ,
    \Tile_X2Y6_FrameData_O[13] ,
    \Tile_X2Y6_FrameData_O[12] ,
    \Tile_X2Y6_FrameData_O[11] ,
    \Tile_X2Y6_FrameData_O[10] ,
    \Tile_X2Y6_FrameData_O[9] ,
    \Tile_X2Y6_FrameData_O[8] ,
    \Tile_X2Y6_FrameData_O[7] ,
    \Tile_X2Y6_FrameData_O[6] ,
    \Tile_X2Y6_FrameData_O[5] ,
    \Tile_X2Y6_FrameData_O[4] ,
    \Tile_X2Y6_FrameData_O[3] ,
    \Tile_X2Y6_FrameData_O[2] ,
    \Tile_X2Y6_FrameData_O[1] ,
    \Tile_X2Y6_FrameData_O[0] }),
    .FrameData_O({\Tile_X3Y6_FrameData_O[31] ,
    \Tile_X3Y6_FrameData_O[30] ,
    \Tile_X3Y6_FrameData_O[29] ,
    \Tile_X3Y6_FrameData_O[28] ,
    \Tile_X3Y6_FrameData_O[27] ,
    \Tile_X3Y6_FrameData_O[26] ,
    \Tile_X3Y6_FrameData_O[25] ,
    \Tile_X3Y6_FrameData_O[24] ,
    \Tile_X3Y6_FrameData_O[23] ,
    \Tile_X3Y6_FrameData_O[22] ,
    \Tile_X3Y6_FrameData_O[21] ,
    \Tile_X3Y6_FrameData_O[20] ,
    \Tile_X3Y6_FrameData_O[19] ,
    \Tile_X3Y6_FrameData_O[18] ,
    \Tile_X3Y6_FrameData_O[17] ,
    \Tile_X3Y6_FrameData_O[16] ,
    \Tile_X3Y6_FrameData_O[15] ,
    \Tile_X3Y6_FrameData_O[14] ,
    \Tile_X3Y6_FrameData_O[13] ,
    \Tile_X3Y6_FrameData_O[12] ,
    \Tile_X3Y6_FrameData_O[11] ,
    \Tile_X3Y6_FrameData_O[10] ,
    \Tile_X3Y6_FrameData_O[9] ,
    \Tile_X3Y6_FrameData_O[8] ,
    \Tile_X3Y6_FrameData_O[7] ,
    \Tile_X3Y6_FrameData_O[6] ,
    \Tile_X3Y6_FrameData_O[5] ,
    \Tile_X3Y6_FrameData_O[4] ,
    \Tile_X3Y6_FrameData_O[3] ,
    \Tile_X3Y6_FrameData_O[2] ,
    \Tile_X3Y6_FrameData_O[1] ,
    \Tile_X3Y6_FrameData_O[0] }),
    .FrameStrobe({\Tile_X3Y7_FrameStrobe_O[19] ,
    \Tile_X3Y7_FrameStrobe_O[18] ,
    \Tile_X3Y7_FrameStrobe_O[17] ,
    \Tile_X3Y7_FrameStrobe_O[16] ,
    \Tile_X3Y7_FrameStrobe_O[15] ,
    \Tile_X3Y7_FrameStrobe_O[14] ,
    \Tile_X3Y7_FrameStrobe_O[13] ,
    \Tile_X3Y7_FrameStrobe_O[12] ,
    \Tile_X3Y7_FrameStrobe_O[11] ,
    \Tile_X3Y7_FrameStrobe_O[10] ,
    \Tile_X3Y7_FrameStrobe_O[9] ,
    \Tile_X3Y7_FrameStrobe_O[8] ,
    \Tile_X3Y7_FrameStrobe_O[7] ,
    \Tile_X3Y7_FrameStrobe_O[6] ,
    \Tile_X3Y7_FrameStrobe_O[5] ,
    \Tile_X3Y7_FrameStrobe_O[4] ,
    \Tile_X3Y7_FrameStrobe_O[3] ,
    \Tile_X3Y7_FrameStrobe_O[2] ,
    \Tile_X3Y7_FrameStrobe_O[1] ,
    \Tile_X3Y7_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X3Y6_FrameStrobe_O[19] ,
    \Tile_X3Y6_FrameStrobe_O[18] ,
    \Tile_X3Y6_FrameStrobe_O[17] ,
    \Tile_X3Y6_FrameStrobe_O[16] ,
    \Tile_X3Y6_FrameStrobe_O[15] ,
    \Tile_X3Y6_FrameStrobe_O[14] ,
    \Tile_X3Y6_FrameStrobe_O[13] ,
    \Tile_X3Y6_FrameStrobe_O[12] ,
    \Tile_X3Y6_FrameStrobe_O[11] ,
    \Tile_X3Y6_FrameStrobe_O[10] ,
    \Tile_X3Y6_FrameStrobe_O[9] ,
    \Tile_X3Y6_FrameStrobe_O[8] ,
    \Tile_X3Y6_FrameStrobe_O[7] ,
    \Tile_X3Y6_FrameStrobe_O[6] ,
    \Tile_X3Y6_FrameStrobe_O[5] ,
    \Tile_X3Y6_FrameStrobe_O[4] ,
    \Tile_X3Y6_FrameStrobe_O[3] ,
    \Tile_X3Y6_FrameStrobe_O[2] ,
    \Tile_X3Y6_FrameStrobe_O[1] ,
    \Tile_X3Y6_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X3Y6_N1BEG[3] ,
    \Tile_X3Y6_N1BEG[2] ,
    \Tile_X3Y6_N1BEG[1] ,
    \Tile_X3Y6_N1BEG[0] }),
    .N1END({\Tile_X3Y7_N1BEG[3] ,
    \Tile_X3Y7_N1BEG[2] ,
    \Tile_X3Y7_N1BEG[1] ,
    \Tile_X3Y7_N1BEG[0] }),
    .N2BEG({\Tile_X3Y6_N2BEG[7] ,
    \Tile_X3Y6_N2BEG[6] ,
    \Tile_X3Y6_N2BEG[5] ,
    \Tile_X3Y6_N2BEG[4] ,
    \Tile_X3Y6_N2BEG[3] ,
    \Tile_X3Y6_N2BEG[2] ,
    \Tile_X3Y6_N2BEG[1] ,
    \Tile_X3Y6_N2BEG[0] }),
    .N2BEGb({\Tile_X3Y6_N2BEGb[7] ,
    \Tile_X3Y6_N2BEGb[6] ,
    \Tile_X3Y6_N2BEGb[5] ,
    \Tile_X3Y6_N2BEGb[4] ,
    \Tile_X3Y6_N2BEGb[3] ,
    \Tile_X3Y6_N2BEGb[2] ,
    \Tile_X3Y6_N2BEGb[1] ,
    \Tile_X3Y6_N2BEGb[0] }),
    .N2END({\Tile_X3Y7_N2BEGb[7] ,
    \Tile_X3Y7_N2BEGb[6] ,
    \Tile_X3Y7_N2BEGb[5] ,
    \Tile_X3Y7_N2BEGb[4] ,
    \Tile_X3Y7_N2BEGb[3] ,
    \Tile_X3Y7_N2BEGb[2] ,
    \Tile_X3Y7_N2BEGb[1] ,
    \Tile_X3Y7_N2BEGb[0] }),
    .N2MID({\Tile_X3Y7_N2BEG[7] ,
    \Tile_X3Y7_N2BEG[6] ,
    \Tile_X3Y7_N2BEG[5] ,
    \Tile_X3Y7_N2BEG[4] ,
    \Tile_X3Y7_N2BEG[3] ,
    \Tile_X3Y7_N2BEG[2] ,
    \Tile_X3Y7_N2BEG[1] ,
    \Tile_X3Y7_N2BEG[0] }),
    .N4BEG({\Tile_X3Y6_N4BEG[15] ,
    \Tile_X3Y6_N4BEG[14] ,
    \Tile_X3Y6_N4BEG[13] ,
    \Tile_X3Y6_N4BEG[12] ,
    \Tile_X3Y6_N4BEG[11] ,
    \Tile_X3Y6_N4BEG[10] ,
    \Tile_X3Y6_N4BEG[9] ,
    \Tile_X3Y6_N4BEG[8] ,
    \Tile_X3Y6_N4BEG[7] ,
    \Tile_X3Y6_N4BEG[6] ,
    \Tile_X3Y6_N4BEG[5] ,
    \Tile_X3Y6_N4BEG[4] ,
    \Tile_X3Y6_N4BEG[3] ,
    \Tile_X3Y6_N4BEG[2] ,
    \Tile_X3Y6_N4BEG[1] ,
    \Tile_X3Y6_N4BEG[0] }),
    .N4END({\Tile_X3Y7_N4BEG[15] ,
    \Tile_X3Y7_N4BEG[14] ,
    \Tile_X3Y7_N4BEG[13] ,
    \Tile_X3Y7_N4BEG[12] ,
    \Tile_X3Y7_N4BEG[11] ,
    \Tile_X3Y7_N4BEG[10] ,
    \Tile_X3Y7_N4BEG[9] ,
    \Tile_X3Y7_N4BEG[8] ,
    \Tile_X3Y7_N4BEG[7] ,
    \Tile_X3Y7_N4BEG[6] ,
    \Tile_X3Y7_N4BEG[5] ,
    \Tile_X3Y7_N4BEG[4] ,
    \Tile_X3Y7_N4BEG[3] ,
    \Tile_X3Y7_N4BEG[2] ,
    \Tile_X3Y7_N4BEG[1] ,
    \Tile_X3Y7_N4BEG[0] }),
    .NN4BEG({\Tile_X3Y6_NN4BEG[15] ,
    \Tile_X3Y6_NN4BEG[14] ,
    \Tile_X3Y6_NN4BEG[13] ,
    \Tile_X3Y6_NN4BEG[12] ,
    \Tile_X3Y6_NN4BEG[11] ,
    \Tile_X3Y6_NN4BEG[10] ,
    \Tile_X3Y6_NN4BEG[9] ,
    \Tile_X3Y6_NN4BEG[8] ,
    \Tile_X3Y6_NN4BEG[7] ,
    \Tile_X3Y6_NN4BEG[6] ,
    \Tile_X3Y6_NN4BEG[5] ,
    \Tile_X3Y6_NN4BEG[4] ,
    \Tile_X3Y6_NN4BEG[3] ,
    \Tile_X3Y6_NN4BEG[2] ,
    \Tile_X3Y6_NN4BEG[1] ,
    \Tile_X3Y6_NN4BEG[0] }),
    .NN4END({\Tile_X3Y7_NN4BEG[15] ,
    \Tile_X3Y7_NN4BEG[14] ,
    \Tile_X3Y7_NN4BEG[13] ,
    \Tile_X3Y7_NN4BEG[12] ,
    \Tile_X3Y7_NN4BEG[11] ,
    \Tile_X3Y7_NN4BEG[10] ,
    \Tile_X3Y7_NN4BEG[9] ,
    \Tile_X3Y7_NN4BEG[8] ,
    \Tile_X3Y7_NN4BEG[7] ,
    \Tile_X3Y7_NN4BEG[6] ,
    \Tile_X3Y7_NN4BEG[5] ,
    \Tile_X3Y7_NN4BEG[4] ,
    \Tile_X3Y7_NN4BEG[3] ,
    \Tile_X3Y7_NN4BEG[2] ,
    \Tile_X3Y7_NN4BEG[1] ,
    \Tile_X3Y7_NN4BEG[0] }),
    .S1BEG({\Tile_X3Y6_S1BEG[3] ,
    \Tile_X3Y6_S1BEG[2] ,
    \Tile_X3Y6_S1BEG[1] ,
    \Tile_X3Y6_S1BEG[0] }),
    .S1END({\Tile_X3Y5_S1BEG[3] ,
    \Tile_X3Y5_S1BEG[2] ,
    \Tile_X3Y5_S1BEG[1] ,
    \Tile_X3Y5_S1BEG[0] }),
    .S2BEG({\Tile_X3Y6_S2BEG[7] ,
    \Tile_X3Y6_S2BEG[6] ,
    \Tile_X3Y6_S2BEG[5] ,
    \Tile_X3Y6_S2BEG[4] ,
    \Tile_X3Y6_S2BEG[3] ,
    \Tile_X3Y6_S2BEG[2] ,
    \Tile_X3Y6_S2BEG[1] ,
    \Tile_X3Y6_S2BEG[0] }),
    .S2BEGb({\Tile_X3Y6_S2BEGb[7] ,
    \Tile_X3Y6_S2BEGb[6] ,
    \Tile_X3Y6_S2BEGb[5] ,
    \Tile_X3Y6_S2BEGb[4] ,
    \Tile_X3Y6_S2BEGb[3] ,
    \Tile_X3Y6_S2BEGb[2] ,
    \Tile_X3Y6_S2BEGb[1] ,
    \Tile_X3Y6_S2BEGb[0] }),
    .S2END({\Tile_X3Y5_S2BEGb[7] ,
    \Tile_X3Y5_S2BEGb[6] ,
    \Tile_X3Y5_S2BEGb[5] ,
    \Tile_X3Y5_S2BEGb[4] ,
    \Tile_X3Y5_S2BEGb[3] ,
    \Tile_X3Y5_S2BEGb[2] ,
    \Tile_X3Y5_S2BEGb[1] ,
    \Tile_X3Y5_S2BEGb[0] }),
    .S2MID({\Tile_X3Y5_S2BEG[7] ,
    \Tile_X3Y5_S2BEG[6] ,
    \Tile_X3Y5_S2BEG[5] ,
    \Tile_X3Y5_S2BEG[4] ,
    \Tile_X3Y5_S2BEG[3] ,
    \Tile_X3Y5_S2BEG[2] ,
    \Tile_X3Y5_S2BEG[1] ,
    \Tile_X3Y5_S2BEG[0] }),
    .S4BEG({\Tile_X3Y6_S4BEG[15] ,
    \Tile_X3Y6_S4BEG[14] ,
    \Tile_X3Y6_S4BEG[13] ,
    \Tile_X3Y6_S4BEG[12] ,
    \Tile_X3Y6_S4BEG[11] ,
    \Tile_X3Y6_S4BEG[10] ,
    \Tile_X3Y6_S4BEG[9] ,
    \Tile_X3Y6_S4BEG[8] ,
    \Tile_X3Y6_S4BEG[7] ,
    \Tile_X3Y6_S4BEG[6] ,
    \Tile_X3Y6_S4BEG[5] ,
    \Tile_X3Y6_S4BEG[4] ,
    \Tile_X3Y6_S4BEG[3] ,
    \Tile_X3Y6_S4BEG[2] ,
    \Tile_X3Y6_S4BEG[1] ,
    \Tile_X3Y6_S4BEG[0] }),
    .S4END({\Tile_X3Y5_S4BEG[15] ,
    \Tile_X3Y5_S4BEG[14] ,
    \Tile_X3Y5_S4BEG[13] ,
    \Tile_X3Y5_S4BEG[12] ,
    \Tile_X3Y5_S4BEG[11] ,
    \Tile_X3Y5_S4BEG[10] ,
    \Tile_X3Y5_S4BEG[9] ,
    \Tile_X3Y5_S4BEG[8] ,
    \Tile_X3Y5_S4BEG[7] ,
    \Tile_X3Y5_S4BEG[6] ,
    \Tile_X3Y5_S4BEG[5] ,
    \Tile_X3Y5_S4BEG[4] ,
    \Tile_X3Y5_S4BEG[3] ,
    \Tile_X3Y5_S4BEG[2] ,
    \Tile_X3Y5_S4BEG[1] ,
    \Tile_X3Y5_S4BEG[0] }),
    .SS4BEG({\Tile_X3Y6_SS4BEG[15] ,
    \Tile_X3Y6_SS4BEG[14] ,
    \Tile_X3Y6_SS4BEG[13] ,
    \Tile_X3Y6_SS4BEG[12] ,
    \Tile_X3Y6_SS4BEG[11] ,
    \Tile_X3Y6_SS4BEG[10] ,
    \Tile_X3Y6_SS4BEG[9] ,
    \Tile_X3Y6_SS4BEG[8] ,
    \Tile_X3Y6_SS4BEG[7] ,
    \Tile_X3Y6_SS4BEG[6] ,
    \Tile_X3Y6_SS4BEG[5] ,
    \Tile_X3Y6_SS4BEG[4] ,
    \Tile_X3Y6_SS4BEG[3] ,
    \Tile_X3Y6_SS4BEG[2] ,
    \Tile_X3Y6_SS4BEG[1] ,
    \Tile_X3Y6_SS4BEG[0] }),
    .SS4END({\Tile_X3Y5_SS4BEG[15] ,
    \Tile_X3Y5_SS4BEG[14] ,
    \Tile_X3Y5_SS4BEG[13] ,
    \Tile_X3Y5_SS4BEG[12] ,
    \Tile_X3Y5_SS4BEG[11] ,
    \Tile_X3Y5_SS4BEG[10] ,
    \Tile_X3Y5_SS4BEG[9] ,
    \Tile_X3Y5_SS4BEG[8] ,
    \Tile_X3Y5_SS4BEG[7] ,
    \Tile_X3Y5_SS4BEG[6] ,
    \Tile_X3Y5_SS4BEG[5] ,
    \Tile_X3Y5_SS4BEG[4] ,
    \Tile_X3Y5_SS4BEG[3] ,
    \Tile_X3Y5_SS4BEG[2] ,
    \Tile_X3Y5_SS4BEG[1] ,
    \Tile_X3Y5_SS4BEG[0] }),
    .W1BEG({\Tile_X3Y6_W1BEG[3] ,
    \Tile_X3Y6_W1BEG[2] ,
    \Tile_X3Y6_W1BEG[1] ,
    \Tile_X3Y6_W1BEG[0] }),
    .W1END({\Tile_X4Y6_W1BEG[3] ,
    \Tile_X4Y6_W1BEG[2] ,
    \Tile_X4Y6_W1BEG[1] ,
    \Tile_X4Y6_W1BEG[0] }),
    .W2BEG({\Tile_X3Y6_W2BEG[7] ,
    \Tile_X3Y6_W2BEG[6] ,
    \Tile_X3Y6_W2BEG[5] ,
    \Tile_X3Y6_W2BEG[4] ,
    \Tile_X3Y6_W2BEG[3] ,
    \Tile_X3Y6_W2BEG[2] ,
    \Tile_X3Y6_W2BEG[1] ,
    \Tile_X3Y6_W2BEG[0] }),
    .W2BEGb({\Tile_X3Y6_W2BEGb[7] ,
    \Tile_X3Y6_W2BEGb[6] ,
    \Tile_X3Y6_W2BEGb[5] ,
    \Tile_X3Y6_W2BEGb[4] ,
    \Tile_X3Y6_W2BEGb[3] ,
    \Tile_X3Y6_W2BEGb[2] ,
    \Tile_X3Y6_W2BEGb[1] ,
    \Tile_X3Y6_W2BEGb[0] }),
    .W2END({\Tile_X4Y6_W2BEGb[7] ,
    \Tile_X4Y6_W2BEGb[6] ,
    \Tile_X4Y6_W2BEGb[5] ,
    \Tile_X4Y6_W2BEGb[4] ,
    \Tile_X4Y6_W2BEGb[3] ,
    \Tile_X4Y6_W2BEGb[2] ,
    \Tile_X4Y6_W2BEGb[1] ,
    \Tile_X4Y6_W2BEGb[0] }),
    .W2MID({\Tile_X4Y6_W2BEG[7] ,
    \Tile_X4Y6_W2BEG[6] ,
    \Tile_X4Y6_W2BEG[5] ,
    \Tile_X4Y6_W2BEG[4] ,
    \Tile_X4Y6_W2BEG[3] ,
    \Tile_X4Y6_W2BEG[2] ,
    \Tile_X4Y6_W2BEG[1] ,
    \Tile_X4Y6_W2BEG[0] }),
    .W6BEG({\Tile_X3Y6_W6BEG[11] ,
    \Tile_X3Y6_W6BEG[10] ,
    \Tile_X3Y6_W6BEG[9] ,
    \Tile_X3Y6_W6BEG[8] ,
    \Tile_X3Y6_W6BEG[7] ,
    \Tile_X3Y6_W6BEG[6] ,
    \Tile_X3Y6_W6BEG[5] ,
    \Tile_X3Y6_W6BEG[4] ,
    \Tile_X3Y6_W6BEG[3] ,
    \Tile_X3Y6_W6BEG[2] ,
    \Tile_X3Y6_W6BEG[1] ,
    \Tile_X3Y6_W6BEG[0] }),
    .W6END({\Tile_X4Y6_W6BEG[11] ,
    \Tile_X4Y6_W6BEG[10] ,
    \Tile_X4Y6_W6BEG[9] ,
    \Tile_X4Y6_W6BEG[8] ,
    \Tile_X4Y6_W6BEG[7] ,
    \Tile_X4Y6_W6BEG[6] ,
    \Tile_X4Y6_W6BEG[5] ,
    \Tile_X4Y6_W6BEG[4] ,
    \Tile_X4Y6_W6BEG[3] ,
    \Tile_X4Y6_W6BEG[2] ,
    \Tile_X4Y6_W6BEG[1] ,
    \Tile_X4Y6_W6BEG[0] }),
    .WW4BEG({\Tile_X3Y6_WW4BEG[15] ,
    \Tile_X3Y6_WW4BEG[14] ,
    \Tile_X3Y6_WW4BEG[13] ,
    \Tile_X3Y6_WW4BEG[12] ,
    \Tile_X3Y6_WW4BEG[11] ,
    \Tile_X3Y6_WW4BEG[10] ,
    \Tile_X3Y6_WW4BEG[9] ,
    \Tile_X3Y6_WW4BEG[8] ,
    \Tile_X3Y6_WW4BEG[7] ,
    \Tile_X3Y6_WW4BEG[6] ,
    \Tile_X3Y6_WW4BEG[5] ,
    \Tile_X3Y6_WW4BEG[4] ,
    \Tile_X3Y6_WW4BEG[3] ,
    \Tile_X3Y6_WW4BEG[2] ,
    \Tile_X3Y6_WW4BEG[1] ,
    \Tile_X3Y6_WW4BEG[0] }),
    .WW4END({\Tile_X4Y6_WW4BEG[15] ,
    \Tile_X4Y6_WW4BEG[14] ,
    \Tile_X4Y6_WW4BEG[13] ,
    \Tile_X4Y6_WW4BEG[12] ,
    \Tile_X4Y6_WW4BEG[11] ,
    \Tile_X4Y6_WW4BEG[10] ,
    \Tile_X4Y6_WW4BEG[9] ,
    \Tile_X4Y6_WW4BEG[8] ,
    \Tile_X4Y6_WW4BEG[7] ,
    \Tile_X4Y6_WW4BEG[6] ,
    \Tile_X4Y6_WW4BEG[5] ,
    \Tile_X4Y6_WW4BEG[4] ,
    \Tile_X4Y6_WW4BEG[3] ,
    \Tile_X4Y6_WW4BEG[2] ,
    \Tile_X4Y6_WW4BEG[1] ,
    \Tile_X4Y6_WW4BEG[0] }));
 LUT4AB Tile_X3Y7_LUT4AB (.Ci(Tile_X3Y8_Co),
    .Co(Tile_X3Y7_Co),
    .UserCLK(Tile_X3Y8_UserCLKo),
    .UserCLKo(Tile_X3Y7_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X3Y7_E1BEG[3] ,
    \Tile_X3Y7_E1BEG[2] ,
    \Tile_X3Y7_E1BEG[1] ,
    \Tile_X3Y7_E1BEG[0] }),
    .E1END({\Tile_X2Y7_E1BEG[3] ,
    \Tile_X2Y7_E1BEG[2] ,
    \Tile_X2Y7_E1BEG[1] ,
    \Tile_X2Y7_E1BEG[0] }),
    .E2BEG({\Tile_X3Y7_E2BEG[7] ,
    \Tile_X3Y7_E2BEG[6] ,
    \Tile_X3Y7_E2BEG[5] ,
    \Tile_X3Y7_E2BEG[4] ,
    \Tile_X3Y7_E2BEG[3] ,
    \Tile_X3Y7_E2BEG[2] ,
    \Tile_X3Y7_E2BEG[1] ,
    \Tile_X3Y7_E2BEG[0] }),
    .E2BEGb({\Tile_X3Y7_E2BEGb[7] ,
    \Tile_X3Y7_E2BEGb[6] ,
    \Tile_X3Y7_E2BEGb[5] ,
    \Tile_X3Y7_E2BEGb[4] ,
    \Tile_X3Y7_E2BEGb[3] ,
    \Tile_X3Y7_E2BEGb[2] ,
    \Tile_X3Y7_E2BEGb[1] ,
    \Tile_X3Y7_E2BEGb[0] }),
    .E2END({\Tile_X2Y7_E2BEGb[7] ,
    \Tile_X2Y7_E2BEGb[6] ,
    \Tile_X2Y7_E2BEGb[5] ,
    \Tile_X2Y7_E2BEGb[4] ,
    \Tile_X2Y7_E2BEGb[3] ,
    \Tile_X2Y7_E2BEGb[2] ,
    \Tile_X2Y7_E2BEGb[1] ,
    \Tile_X2Y7_E2BEGb[0] }),
    .E2MID({\Tile_X2Y7_E2BEG[7] ,
    \Tile_X2Y7_E2BEG[6] ,
    \Tile_X2Y7_E2BEG[5] ,
    \Tile_X2Y7_E2BEG[4] ,
    \Tile_X2Y7_E2BEG[3] ,
    \Tile_X2Y7_E2BEG[2] ,
    \Tile_X2Y7_E2BEG[1] ,
    \Tile_X2Y7_E2BEG[0] }),
    .E6BEG({\Tile_X3Y7_E6BEG[11] ,
    \Tile_X3Y7_E6BEG[10] ,
    \Tile_X3Y7_E6BEG[9] ,
    \Tile_X3Y7_E6BEG[8] ,
    \Tile_X3Y7_E6BEG[7] ,
    \Tile_X3Y7_E6BEG[6] ,
    \Tile_X3Y7_E6BEG[5] ,
    \Tile_X3Y7_E6BEG[4] ,
    \Tile_X3Y7_E6BEG[3] ,
    \Tile_X3Y7_E6BEG[2] ,
    \Tile_X3Y7_E6BEG[1] ,
    \Tile_X3Y7_E6BEG[0] }),
    .E6END({\Tile_X2Y7_E6BEG[11] ,
    \Tile_X2Y7_E6BEG[10] ,
    \Tile_X2Y7_E6BEG[9] ,
    \Tile_X2Y7_E6BEG[8] ,
    \Tile_X2Y7_E6BEG[7] ,
    \Tile_X2Y7_E6BEG[6] ,
    \Tile_X2Y7_E6BEG[5] ,
    \Tile_X2Y7_E6BEG[4] ,
    \Tile_X2Y7_E6BEG[3] ,
    \Tile_X2Y7_E6BEG[2] ,
    \Tile_X2Y7_E6BEG[1] ,
    \Tile_X2Y7_E6BEG[0] }),
    .EE4BEG({\Tile_X3Y7_EE4BEG[15] ,
    \Tile_X3Y7_EE4BEG[14] ,
    \Tile_X3Y7_EE4BEG[13] ,
    \Tile_X3Y7_EE4BEG[12] ,
    \Tile_X3Y7_EE4BEG[11] ,
    \Tile_X3Y7_EE4BEG[10] ,
    \Tile_X3Y7_EE4BEG[9] ,
    \Tile_X3Y7_EE4BEG[8] ,
    \Tile_X3Y7_EE4BEG[7] ,
    \Tile_X3Y7_EE4BEG[6] ,
    \Tile_X3Y7_EE4BEG[5] ,
    \Tile_X3Y7_EE4BEG[4] ,
    \Tile_X3Y7_EE4BEG[3] ,
    \Tile_X3Y7_EE4BEG[2] ,
    \Tile_X3Y7_EE4BEG[1] ,
    \Tile_X3Y7_EE4BEG[0] }),
    .EE4END({\Tile_X2Y7_EE4BEG[15] ,
    \Tile_X2Y7_EE4BEG[14] ,
    \Tile_X2Y7_EE4BEG[13] ,
    \Tile_X2Y7_EE4BEG[12] ,
    \Tile_X2Y7_EE4BEG[11] ,
    \Tile_X2Y7_EE4BEG[10] ,
    \Tile_X2Y7_EE4BEG[9] ,
    \Tile_X2Y7_EE4BEG[8] ,
    \Tile_X2Y7_EE4BEG[7] ,
    \Tile_X2Y7_EE4BEG[6] ,
    \Tile_X2Y7_EE4BEG[5] ,
    \Tile_X2Y7_EE4BEG[4] ,
    \Tile_X2Y7_EE4BEG[3] ,
    \Tile_X2Y7_EE4BEG[2] ,
    \Tile_X2Y7_EE4BEG[1] ,
    \Tile_X2Y7_EE4BEG[0] }),
    .FrameData({\Tile_X2Y7_FrameData_O[31] ,
    \Tile_X2Y7_FrameData_O[30] ,
    \Tile_X2Y7_FrameData_O[29] ,
    \Tile_X2Y7_FrameData_O[28] ,
    \Tile_X2Y7_FrameData_O[27] ,
    \Tile_X2Y7_FrameData_O[26] ,
    \Tile_X2Y7_FrameData_O[25] ,
    \Tile_X2Y7_FrameData_O[24] ,
    \Tile_X2Y7_FrameData_O[23] ,
    \Tile_X2Y7_FrameData_O[22] ,
    \Tile_X2Y7_FrameData_O[21] ,
    \Tile_X2Y7_FrameData_O[20] ,
    \Tile_X2Y7_FrameData_O[19] ,
    \Tile_X2Y7_FrameData_O[18] ,
    \Tile_X2Y7_FrameData_O[17] ,
    \Tile_X2Y7_FrameData_O[16] ,
    \Tile_X2Y7_FrameData_O[15] ,
    \Tile_X2Y7_FrameData_O[14] ,
    \Tile_X2Y7_FrameData_O[13] ,
    \Tile_X2Y7_FrameData_O[12] ,
    \Tile_X2Y7_FrameData_O[11] ,
    \Tile_X2Y7_FrameData_O[10] ,
    \Tile_X2Y7_FrameData_O[9] ,
    \Tile_X2Y7_FrameData_O[8] ,
    \Tile_X2Y7_FrameData_O[7] ,
    \Tile_X2Y7_FrameData_O[6] ,
    \Tile_X2Y7_FrameData_O[5] ,
    \Tile_X2Y7_FrameData_O[4] ,
    \Tile_X2Y7_FrameData_O[3] ,
    \Tile_X2Y7_FrameData_O[2] ,
    \Tile_X2Y7_FrameData_O[1] ,
    \Tile_X2Y7_FrameData_O[0] }),
    .FrameData_O({\Tile_X3Y7_FrameData_O[31] ,
    \Tile_X3Y7_FrameData_O[30] ,
    \Tile_X3Y7_FrameData_O[29] ,
    \Tile_X3Y7_FrameData_O[28] ,
    \Tile_X3Y7_FrameData_O[27] ,
    \Tile_X3Y7_FrameData_O[26] ,
    \Tile_X3Y7_FrameData_O[25] ,
    \Tile_X3Y7_FrameData_O[24] ,
    \Tile_X3Y7_FrameData_O[23] ,
    \Tile_X3Y7_FrameData_O[22] ,
    \Tile_X3Y7_FrameData_O[21] ,
    \Tile_X3Y7_FrameData_O[20] ,
    \Tile_X3Y7_FrameData_O[19] ,
    \Tile_X3Y7_FrameData_O[18] ,
    \Tile_X3Y7_FrameData_O[17] ,
    \Tile_X3Y7_FrameData_O[16] ,
    \Tile_X3Y7_FrameData_O[15] ,
    \Tile_X3Y7_FrameData_O[14] ,
    \Tile_X3Y7_FrameData_O[13] ,
    \Tile_X3Y7_FrameData_O[12] ,
    \Tile_X3Y7_FrameData_O[11] ,
    \Tile_X3Y7_FrameData_O[10] ,
    \Tile_X3Y7_FrameData_O[9] ,
    \Tile_X3Y7_FrameData_O[8] ,
    \Tile_X3Y7_FrameData_O[7] ,
    \Tile_X3Y7_FrameData_O[6] ,
    \Tile_X3Y7_FrameData_O[5] ,
    \Tile_X3Y7_FrameData_O[4] ,
    \Tile_X3Y7_FrameData_O[3] ,
    \Tile_X3Y7_FrameData_O[2] ,
    \Tile_X3Y7_FrameData_O[1] ,
    \Tile_X3Y7_FrameData_O[0] }),
    .FrameStrobe({\Tile_X3Y8_FrameStrobe_O[19] ,
    \Tile_X3Y8_FrameStrobe_O[18] ,
    \Tile_X3Y8_FrameStrobe_O[17] ,
    \Tile_X3Y8_FrameStrobe_O[16] ,
    \Tile_X3Y8_FrameStrobe_O[15] ,
    \Tile_X3Y8_FrameStrobe_O[14] ,
    \Tile_X3Y8_FrameStrobe_O[13] ,
    \Tile_X3Y8_FrameStrobe_O[12] ,
    \Tile_X3Y8_FrameStrobe_O[11] ,
    \Tile_X3Y8_FrameStrobe_O[10] ,
    \Tile_X3Y8_FrameStrobe_O[9] ,
    \Tile_X3Y8_FrameStrobe_O[8] ,
    \Tile_X3Y8_FrameStrobe_O[7] ,
    \Tile_X3Y8_FrameStrobe_O[6] ,
    \Tile_X3Y8_FrameStrobe_O[5] ,
    \Tile_X3Y8_FrameStrobe_O[4] ,
    \Tile_X3Y8_FrameStrobe_O[3] ,
    \Tile_X3Y8_FrameStrobe_O[2] ,
    \Tile_X3Y8_FrameStrobe_O[1] ,
    \Tile_X3Y8_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X3Y7_FrameStrobe_O[19] ,
    \Tile_X3Y7_FrameStrobe_O[18] ,
    \Tile_X3Y7_FrameStrobe_O[17] ,
    \Tile_X3Y7_FrameStrobe_O[16] ,
    \Tile_X3Y7_FrameStrobe_O[15] ,
    \Tile_X3Y7_FrameStrobe_O[14] ,
    \Tile_X3Y7_FrameStrobe_O[13] ,
    \Tile_X3Y7_FrameStrobe_O[12] ,
    \Tile_X3Y7_FrameStrobe_O[11] ,
    \Tile_X3Y7_FrameStrobe_O[10] ,
    \Tile_X3Y7_FrameStrobe_O[9] ,
    \Tile_X3Y7_FrameStrobe_O[8] ,
    \Tile_X3Y7_FrameStrobe_O[7] ,
    \Tile_X3Y7_FrameStrobe_O[6] ,
    \Tile_X3Y7_FrameStrobe_O[5] ,
    \Tile_X3Y7_FrameStrobe_O[4] ,
    \Tile_X3Y7_FrameStrobe_O[3] ,
    \Tile_X3Y7_FrameStrobe_O[2] ,
    \Tile_X3Y7_FrameStrobe_O[1] ,
    \Tile_X3Y7_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X3Y7_N1BEG[3] ,
    \Tile_X3Y7_N1BEG[2] ,
    \Tile_X3Y7_N1BEG[1] ,
    \Tile_X3Y7_N1BEG[0] }),
    .N1END({\Tile_X3Y8_N1BEG[3] ,
    \Tile_X3Y8_N1BEG[2] ,
    \Tile_X3Y8_N1BEG[1] ,
    \Tile_X3Y8_N1BEG[0] }),
    .N2BEG({\Tile_X3Y7_N2BEG[7] ,
    \Tile_X3Y7_N2BEG[6] ,
    \Tile_X3Y7_N2BEG[5] ,
    \Tile_X3Y7_N2BEG[4] ,
    \Tile_X3Y7_N2BEG[3] ,
    \Tile_X3Y7_N2BEG[2] ,
    \Tile_X3Y7_N2BEG[1] ,
    \Tile_X3Y7_N2BEG[0] }),
    .N2BEGb({\Tile_X3Y7_N2BEGb[7] ,
    \Tile_X3Y7_N2BEGb[6] ,
    \Tile_X3Y7_N2BEGb[5] ,
    \Tile_X3Y7_N2BEGb[4] ,
    \Tile_X3Y7_N2BEGb[3] ,
    \Tile_X3Y7_N2BEGb[2] ,
    \Tile_X3Y7_N2BEGb[1] ,
    \Tile_X3Y7_N2BEGb[0] }),
    .N2END({\Tile_X3Y8_N2BEGb[7] ,
    \Tile_X3Y8_N2BEGb[6] ,
    \Tile_X3Y8_N2BEGb[5] ,
    \Tile_X3Y8_N2BEGb[4] ,
    \Tile_X3Y8_N2BEGb[3] ,
    \Tile_X3Y8_N2BEGb[2] ,
    \Tile_X3Y8_N2BEGb[1] ,
    \Tile_X3Y8_N2BEGb[0] }),
    .N2MID({\Tile_X3Y8_N2BEG[7] ,
    \Tile_X3Y8_N2BEG[6] ,
    \Tile_X3Y8_N2BEG[5] ,
    \Tile_X3Y8_N2BEG[4] ,
    \Tile_X3Y8_N2BEG[3] ,
    \Tile_X3Y8_N2BEG[2] ,
    \Tile_X3Y8_N2BEG[1] ,
    \Tile_X3Y8_N2BEG[0] }),
    .N4BEG({\Tile_X3Y7_N4BEG[15] ,
    \Tile_X3Y7_N4BEG[14] ,
    \Tile_X3Y7_N4BEG[13] ,
    \Tile_X3Y7_N4BEG[12] ,
    \Tile_X3Y7_N4BEG[11] ,
    \Tile_X3Y7_N4BEG[10] ,
    \Tile_X3Y7_N4BEG[9] ,
    \Tile_X3Y7_N4BEG[8] ,
    \Tile_X3Y7_N4BEG[7] ,
    \Tile_X3Y7_N4BEG[6] ,
    \Tile_X3Y7_N4BEG[5] ,
    \Tile_X3Y7_N4BEG[4] ,
    \Tile_X3Y7_N4BEG[3] ,
    \Tile_X3Y7_N4BEG[2] ,
    \Tile_X3Y7_N4BEG[1] ,
    \Tile_X3Y7_N4BEG[0] }),
    .N4END({\Tile_X3Y8_N4BEG[15] ,
    \Tile_X3Y8_N4BEG[14] ,
    \Tile_X3Y8_N4BEG[13] ,
    \Tile_X3Y8_N4BEG[12] ,
    \Tile_X3Y8_N4BEG[11] ,
    \Tile_X3Y8_N4BEG[10] ,
    \Tile_X3Y8_N4BEG[9] ,
    \Tile_X3Y8_N4BEG[8] ,
    \Tile_X3Y8_N4BEG[7] ,
    \Tile_X3Y8_N4BEG[6] ,
    \Tile_X3Y8_N4BEG[5] ,
    \Tile_X3Y8_N4BEG[4] ,
    \Tile_X3Y8_N4BEG[3] ,
    \Tile_X3Y8_N4BEG[2] ,
    \Tile_X3Y8_N4BEG[1] ,
    \Tile_X3Y8_N4BEG[0] }),
    .NN4BEG({\Tile_X3Y7_NN4BEG[15] ,
    \Tile_X3Y7_NN4BEG[14] ,
    \Tile_X3Y7_NN4BEG[13] ,
    \Tile_X3Y7_NN4BEG[12] ,
    \Tile_X3Y7_NN4BEG[11] ,
    \Tile_X3Y7_NN4BEG[10] ,
    \Tile_X3Y7_NN4BEG[9] ,
    \Tile_X3Y7_NN4BEG[8] ,
    \Tile_X3Y7_NN4BEG[7] ,
    \Tile_X3Y7_NN4BEG[6] ,
    \Tile_X3Y7_NN4BEG[5] ,
    \Tile_X3Y7_NN4BEG[4] ,
    \Tile_X3Y7_NN4BEG[3] ,
    \Tile_X3Y7_NN4BEG[2] ,
    \Tile_X3Y7_NN4BEG[1] ,
    \Tile_X3Y7_NN4BEG[0] }),
    .NN4END({\Tile_X3Y8_NN4BEG[15] ,
    \Tile_X3Y8_NN4BEG[14] ,
    \Tile_X3Y8_NN4BEG[13] ,
    \Tile_X3Y8_NN4BEG[12] ,
    \Tile_X3Y8_NN4BEG[11] ,
    \Tile_X3Y8_NN4BEG[10] ,
    \Tile_X3Y8_NN4BEG[9] ,
    \Tile_X3Y8_NN4BEG[8] ,
    \Tile_X3Y8_NN4BEG[7] ,
    \Tile_X3Y8_NN4BEG[6] ,
    \Tile_X3Y8_NN4BEG[5] ,
    \Tile_X3Y8_NN4BEG[4] ,
    \Tile_X3Y8_NN4BEG[3] ,
    \Tile_X3Y8_NN4BEG[2] ,
    \Tile_X3Y8_NN4BEG[1] ,
    \Tile_X3Y8_NN4BEG[0] }),
    .S1BEG({\Tile_X3Y7_S1BEG[3] ,
    \Tile_X3Y7_S1BEG[2] ,
    \Tile_X3Y7_S1BEG[1] ,
    \Tile_X3Y7_S1BEG[0] }),
    .S1END({\Tile_X3Y6_S1BEG[3] ,
    \Tile_X3Y6_S1BEG[2] ,
    \Tile_X3Y6_S1BEG[1] ,
    \Tile_X3Y6_S1BEG[0] }),
    .S2BEG({\Tile_X3Y7_S2BEG[7] ,
    \Tile_X3Y7_S2BEG[6] ,
    \Tile_X3Y7_S2BEG[5] ,
    \Tile_X3Y7_S2BEG[4] ,
    \Tile_X3Y7_S2BEG[3] ,
    \Tile_X3Y7_S2BEG[2] ,
    \Tile_X3Y7_S2BEG[1] ,
    \Tile_X3Y7_S2BEG[0] }),
    .S2BEGb({\Tile_X3Y7_S2BEGb[7] ,
    \Tile_X3Y7_S2BEGb[6] ,
    \Tile_X3Y7_S2BEGb[5] ,
    \Tile_X3Y7_S2BEGb[4] ,
    \Tile_X3Y7_S2BEGb[3] ,
    \Tile_X3Y7_S2BEGb[2] ,
    \Tile_X3Y7_S2BEGb[1] ,
    \Tile_X3Y7_S2BEGb[0] }),
    .S2END({\Tile_X3Y6_S2BEGb[7] ,
    \Tile_X3Y6_S2BEGb[6] ,
    \Tile_X3Y6_S2BEGb[5] ,
    \Tile_X3Y6_S2BEGb[4] ,
    \Tile_X3Y6_S2BEGb[3] ,
    \Tile_X3Y6_S2BEGb[2] ,
    \Tile_X3Y6_S2BEGb[1] ,
    \Tile_X3Y6_S2BEGb[0] }),
    .S2MID({\Tile_X3Y6_S2BEG[7] ,
    \Tile_X3Y6_S2BEG[6] ,
    \Tile_X3Y6_S2BEG[5] ,
    \Tile_X3Y6_S2BEG[4] ,
    \Tile_X3Y6_S2BEG[3] ,
    \Tile_X3Y6_S2BEG[2] ,
    \Tile_X3Y6_S2BEG[1] ,
    \Tile_X3Y6_S2BEG[0] }),
    .S4BEG({\Tile_X3Y7_S4BEG[15] ,
    \Tile_X3Y7_S4BEG[14] ,
    \Tile_X3Y7_S4BEG[13] ,
    \Tile_X3Y7_S4BEG[12] ,
    \Tile_X3Y7_S4BEG[11] ,
    \Tile_X3Y7_S4BEG[10] ,
    \Tile_X3Y7_S4BEG[9] ,
    \Tile_X3Y7_S4BEG[8] ,
    \Tile_X3Y7_S4BEG[7] ,
    \Tile_X3Y7_S4BEG[6] ,
    \Tile_X3Y7_S4BEG[5] ,
    \Tile_X3Y7_S4BEG[4] ,
    \Tile_X3Y7_S4BEG[3] ,
    \Tile_X3Y7_S4BEG[2] ,
    \Tile_X3Y7_S4BEG[1] ,
    \Tile_X3Y7_S4BEG[0] }),
    .S4END({\Tile_X3Y6_S4BEG[15] ,
    \Tile_X3Y6_S4BEG[14] ,
    \Tile_X3Y6_S4BEG[13] ,
    \Tile_X3Y6_S4BEG[12] ,
    \Tile_X3Y6_S4BEG[11] ,
    \Tile_X3Y6_S4BEG[10] ,
    \Tile_X3Y6_S4BEG[9] ,
    \Tile_X3Y6_S4BEG[8] ,
    \Tile_X3Y6_S4BEG[7] ,
    \Tile_X3Y6_S4BEG[6] ,
    \Tile_X3Y6_S4BEG[5] ,
    \Tile_X3Y6_S4BEG[4] ,
    \Tile_X3Y6_S4BEG[3] ,
    \Tile_X3Y6_S4BEG[2] ,
    \Tile_X3Y6_S4BEG[1] ,
    \Tile_X3Y6_S4BEG[0] }),
    .SS4BEG({\Tile_X3Y7_SS4BEG[15] ,
    \Tile_X3Y7_SS4BEG[14] ,
    \Tile_X3Y7_SS4BEG[13] ,
    \Tile_X3Y7_SS4BEG[12] ,
    \Tile_X3Y7_SS4BEG[11] ,
    \Tile_X3Y7_SS4BEG[10] ,
    \Tile_X3Y7_SS4BEG[9] ,
    \Tile_X3Y7_SS4BEG[8] ,
    \Tile_X3Y7_SS4BEG[7] ,
    \Tile_X3Y7_SS4BEG[6] ,
    \Tile_X3Y7_SS4BEG[5] ,
    \Tile_X3Y7_SS4BEG[4] ,
    \Tile_X3Y7_SS4BEG[3] ,
    \Tile_X3Y7_SS4BEG[2] ,
    \Tile_X3Y7_SS4BEG[1] ,
    \Tile_X3Y7_SS4BEG[0] }),
    .SS4END({\Tile_X3Y6_SS4BEG[15] ,
    \Tile_X3Y6_SS4BEG[14] ,
    \Tile_X3Y6_SS4BEG[13] ,
    \Tile_X3Y6_SS4BEG[12] ,
    \Tile_X3Y6_SS4BEG[11] ,
    \Tile_X3Y6_SS4BEG[10] ,
    \Tile_X3Y6_SS4BEG[9] ,
    \Tile_X3Y6_SS4BEG[8] ,
    \Tile_X3Y6_SS4BEG[7] ,
    \Tile_X3Y6_SS4BEG[6] ,
    \Tile_X3Y6_SS4BEG[5] ,
    \Tile_X3Y6_SS4BEG[4] ,
    \Tile_X3Y6_SS4BEG[3] ,
    \Tile_X3Y6_SS4BEG[2] ,
    \Tile_X3Y6_SS4BEG[1] ,
    \Tile_X3Y6_SS4BEG[0] }),
    .W1BEG({\Tile_X3Y7_W1BEG[3] ,
    \Tile_X3Y7_W1BEG[2] ,
    \Tile_X3Y7_W1BEG[1] ,
    \Tile_X3Y7_W1BEG[0] }),
    .W1END({\Tile_X4Y7_W1BEG[3] ,
    \Tile_X4Y7_W1BEG[2] ,
    \Tile_X4Y7_W1BEG[1] ,
    \Tile_X4Y7_W1BEG[0] }),
    .W2BEG({\Tile_X3Y7_W2BEG[7] ,
    \Tile_X3Y7_W2BEG[6] ,
    \Tile_X3Y7_W2BEG[5] ,
    \Tile_X3Y7_W2BEG[4] ,
    \Tile_X3Y7_W2BEG[3] ,
    \Tile_X3Y7_W2BEG[2] ,
    \Tile_X3Y7_W2BEG[1] ,
    \Tile_X3Y7_W2BEG[0] }),
    .W2BEGb({\Tile_X3Y7_W2BEGb[7] ,
    \Tile_X3Y7_W2BEGb[6] ,
    \Tile_X3Y7_W2BEGb[5] ,
    \Tile_X3Y7_W2BEGb[4] ,
    \Tile_X3Y7_W2BEGb[3] ,
    \Tile_X3Y7_W2BEGb[2] ,
    \Tile_X3Y7_W2BEGb[1] ,
    \Tile_X3Y7_W2BEGb[0] }),
    .W2END({\Tile_X4Y7_W2BEGb[7] ,
    \Tile_X4Y7_W2BEGb[6] ,
    \Tile_X4Y7_W2BEGb[5] ,
    \Tile_X4Y7_W2BEGb[4] ,
    \Tile_X4Y7_W2BEGb[3] ,
    \Tile_X4Y7_W2BEGb[2] ,
    \Tile_X4Y7_W2BEGb[1] ,
    \Tile_X4Y7_W2BEGb[0] }),
    .W2MID({\Tile_X4Y7_W2BEG[7] ,
    \Tile_X4Y7_W2BEG[6] ,
    \Tile_X4Y7_W2BEG[5] ,
    \Tile_X4Y7_W2BEG[4] ,
    \Tile_X4Y7_W2BEG[3] ,
    \Tile_X4Y7_W2BEG[2] ,
    \Tile_X4Y7_W2BEG[1] ,
    \Tile_X4Y7_W2BEG[0] }),
    .W6BEG({\Tile_X3Y7_W6BEG[11] ,
    \Tile_X3Y7_W6BEG[10] ,
    \Tile_X3Y7_W6BEG[9] ,
    \Tile_X3Y7_W6BEG[8] ,
    \Tile_X3Y7_W6BEG[7] ,
    \Tile_X3Y7_W6BEG[6] ,
    \Tile_X3Y7_W6BEG[5] ,
    \Tile_X3Y7_W6BEG[4] ,
    \Tile_X3Y7_W6BEG[3] ,
    \Tile_X3Y7_W6BEG[2] ,
    \Tile_X3Y7_W6BEG[1] ,
    \Tile_X3Y7_W6BEG[0] }),
    .W6END({\Tile_X4Y7_W6BEG[11] ,
    \Tile_X4Y7_W6BEG[10] ,
    \Tile_X4Y7_W6BEG[9] ,
    \Tile_X4Y7_W6BEG[8] ,
    \Tile_X4Y7_W6BEG[7] ,
    \Tile_X4Y7_W6BEG[6] ,
    \Tile_X4Y7_W6BEG[5] ,
    \Tile_X4Y7_W6BEG[4] ,
    \Tile_X4Y7_W6BEG[3] ,
    \Tile_X4Y7_W6BEG[2] ,
    \Tile_X4Y7_W6BEG[1] ,
    \Tile_X4Y7_W6BEG[0] }),
    .WW4BEG({\Tile_X3Y7_WW4BEG[15] ,
    \Tile_X3Y7_WW4BEG[14] ,
    \Tile_X3Y7_WW4BEG[13] ,
    \Tile_X3Y7_WW4BEG[12] ,
    \Tile_X3Y7_WW4BEG[11] ,
    \Tile_X3Y7_WW4BEG[10] ,
    \Tile_X3Y7_WW4BEG[9] ,
    \Tile_X3Y7_WW4BEG[8] ,
    \Tile_X3Y7_WW4BEG[7] ,
    \Tile_X3Y7_WW4BEG[6] ,
    \Tile_X3Y7_WW4BEG[5] ,
    \Tile_X3Y7_WW4BEG[4] ,
    \Tile_X3Y7_WW4BEG[3] ,
    \Tile_X3Y7_WW4BEG[2] ,
    \Tile_X3Y7_WW4BEG[1] ,
    \Tile_X3Y7_WW4BEG[0] }),
    .WW4END({\Tile_X4Y7_WW4BEG[15] ,
    \Tile_X4Y7_WW4BEG[14] ,
    \Tile_X4Y7_WW4BEG[13] ,
    \Tile_X4Y7_WW4BEG[12] ,
    \Tile_X4Y7_WW4BEG[11] ,
    \Tile_X4Y7_WW4BEG[10] ,
    \Tile_X4Y7_WW4BEG[9] ,
    \Tile_X4Y7_WW4BEG[8] ,
    \Tile_X4Y7_WW4BEG[7] ,
    \Tile_X4Y7_WW4BEG[6] ,
    \Tile_X4Y7_WW4BEG[5] ,
    \Tile_X4Y7_WW4BEG[4] ,
    \Tile_X4Y7_WW4BEG[3] ,
    \Tile_X4Y7_WW4BEG[2] ,
    \Tile_X4Y7_WW4BEG[1] ,
    \Tile_X4Y7_WW4BEG[0] }));
 LUT4AB Tile_X3Y8_LUT4AB (.Ci(Tile_X3Y9_Co),
    .Co(Tile_X3Y8_Co),
    .UserCLK(Tile_X3Y9_UserCLKo),
    .UserCLKo(Tile_X3Y8_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X3Y8_E1BEG[3] ,
    \Tile_X3Y8_E1BEG[2] ,
    \Tile_X3Y8_E1BEG[1] ,
    \Tile_X3Y8_E1BEG[0] }),
    .E1END({\Tile_X2Y8_E1BEG[3] ,
    \Tile_X2Y8_E1BEG[2] ,
    \Tile_X2Y8_E1BEG[1] ,
    \Tile_X2Y8_E1BEG[0] }),
    .E2BEG({\Tile_X3Y8_E2BEG[7] ,
    \Tile_X3Y8_E2BEG[6] ,
    \Tile_X3Y8_E2BEG[5] ,
    \Tile_X3Y8_E2BEG[4] ,
    \Tile_X3Y8_E2BEG[3] ,
    \Tile_X3Y8_E2BEG[2] ,
    \Tile_X3Y8_E2BEG[1] ,
    \Tile_X3Y8_E2BEG[0] }),
    .E2BEGb({\Tile_X3Y8_E2BEGb[7] ,
    \Tile_X3Y8_E2BEGb[6] ,
    \Tile_X3Y8_E2BEGb[5] ,
    \Tile_X3Y8_E2BEGb[4] ,
    \Tile_X3Y8_E2BEGb[3] ,
    \Tile_X3Y8_E2BEGb[2] ,
    \Tile_X3Y8_E2BEGb[1] ,
    \Tile_X3Y8_E2BEGb[0] }),
    .E2END({\Tile_X2Y8_E2BEGb[7] ,
    \Tile_X2Y8_E2BEGb[6] ,
    \Tile_X2Y8_E2BEGb[5] ,
    \Tile_X2Y8_E2BEGb[4] ,
    \Tile_X2Y8_E2BEGb[3] ,
    \Tile_X2Y8_E2BEGb[2] ,
    \Tile_X2Y8_E2BEGb[1] ,
    \Tile_X2Y8_E2BEGb[0] }),
    .E2MID({\Tile_X2Y8_E2BEG[7] ,
    \Tile_X2Y8_E2BEG[6] ,
    \Tile_X2Y8_E2BEG[5] ,
    \Tile_X2Y8_E2BEG[4] ,
    \Tile_X2Y8_E2BEG[3] ,
    \Tile_X2Y8_E2BEG[2] ,
    \Tile_X2Y8_E2BEG[1] ,
    \Tile_X2Y8_E2BEG[0] }),
    .E6BEG({\Tile_X3Y8_E6BEG[11] ,
    \Tile_X3Y8_E6BEG[10] ,
    \Tile_X3Y8_E6BEG[9] ,
    \Tile_X3Y8_E6BEG[8] ,
    \Tile_X3Y8_E6BEG[7] ,
    \Tile_X3Y8_E6BEG[6] ,
    \Tile_X3Y8_E6BEG[5] ,
    \Tile_X3Y8_E6BEG[4] ,
    \Tile_X3Y8_E6BEG[3] ,
    \Tile_X3Y8_E6BEG[2] ,
    \Tile_X3Y8_E6BEG[1] ,
    \Tile_X3Y8_E6BEG[0] }),
    .E6END({\Tile_X2Y8_E6BEG[11] ,
    \Tile_X2Y8_E6BEG[10] ,
    \Tile_X2Y8_E6BEG[9] ,
    \Tile_X2Y8_E6BEG[8] ,
    \Tile_X2Y8_E6BEG[7] ,
    \Tile_X2Y8_E6BEG[6] ,
    \Tile_X2Y8_E6BEG[5] ,
    \Tile_X2Y8_E6BEG[4] ,
    \Tile_X2Y8_E6BEG[3] ,
    \Tile_X2Y8_E6BEG[2] ,
    \Tile_X2Y8_E6BEG[1] ,
    \Tile_X2Y8_E6BEG[0] }),
    .EE4BEG({\Tile_X3Y8_EE4BEG[15] ,
    \Tile_X3Y8_EE4BEG[14] ,
    \Tile_X3Y8_EE4BEG[13] ,
    \Tile_X3Y8_EE4BEG[12] ,
    \Tile_X3Y8_EE4BEG[11] ,
    \Tile_X3Y8_EE4BEG[10] ,
    \Tile_X3Y8_EE4BEG[9] ,
    \Tile_X3Y8_EE4BEG[8] ,
    \Tile_X3Y8_EE4BEG[7] ,
    \Tile_X3Y8_EE4BEG[6] ,
    \Tile_X3Y8_EE4BEG[5] ,
    \Tile_X3Y8_EE4BEG[4] ,
    \Tile_X3Y8_EE4BEG[3] ,
    \Tile_X3Y8_EE4BEG[2] ,
    \Tile_X3Y8_EE4BEG[1] ,
    \Tile_X3Y8_EE4BEG[0] }),
    .EE4END({\Tile_X2Y8_EE4BEG[15] ,
    \Tile_X2Y8_EE4BEG[14] ,
    \Tile_X2Y8_EE4BEG[13] ,
    \Tile_X2Y8_EE4BEG[12] ,
    \Tile_X2Y8_EE4BEG[11] ,
    \Tile_X2Y8_EE4BEG[10] ,
    \Tile_X2Y8_EE4BEG[9] ,
    \Tile_X2Y8_EE4BEG[8] ,
    \Tile_X2Y8_EE4BEG[7] ,
    \Tile_X2Y8_EE4BEG[6] ,
    \Tile_X2Y8_EE4BEG[5] ,
    \Tile_X2Y8_EE4BEG[4] ,
    \Tile_X2Y8_EE4BEG[3] ,
    \Tile_X2Y8_EE4BEG[2] ,
    \Tile_X2Y8_EE4BEG[1] ,
    \Tile_X2Y8_EE4BEG[0] }),
    .FrameData({\Tile_X2Y8_FrameData_O[31] ,
    \Tile_X2Y8_FrameData_O[30] ,
    \Tile_X2Y8_FrameData_O[29] ,
    \Tile_X2Y8_FrameData_O[28] ,
    \Tile_X2Y8_FrameData_O[27] ,
    \Tile_X2Y8_FrameData_O[26] ,
    \Tile_X2Y8_FrameData_O[25] ,
    \Tile_X2Y8_FrameData_O[24] ,
    \Tile_X2Y8_FrameData_O[23] ,
    \Tile_X2Y8_FrameData_O[22] ,
    \Tile_X2Y8_FrameData_O[21] ,
    \Tile_X2Y8_FrameData_O[20] ,
    \Tile_X2Y8_FrameData_O[19] ,
    \Tile_X2Y8_FrameData_O[18] ,
    \Tile_X2Y8_FrameData_O[17] ,
    \Tile_X2Y8_FrameData_O[16] ,
    \Tile_X2Y8_FrameData_O[15] ,
    \Tile_X2Y8_FrameData_O[14] ,
    \Tile_X2Y8_FrameData_O[13] ,
    \Tile_X2Y8_FrameData_O[12] ,
    \Tile_X2Y8_FrameData_O[11] ,
    \Tile_X2Y8_FrameData_O[10] ,
    \Tile_X2Y8_FrameData_O[9] ,
    \Tile_X2Y8_FrameData_O[8] ,
    \Tile_X2Y8_FrameData_O[7] ,
    \Tile_X2Y8_FrameData_O[6] ,
    \Tile_X2Y8_FrameData_O[5] ,
    \Tile_X2Y8_FrameData_O[4] ,
    \Tile_X2Y8_FrameData_O[3] ,
    \Tile_X2Y8_FrameData_O[2] ,
    \Tile_X2Y8_FrameData_O[1] ,
    \Tile_X2Y8_FrameData_O[0] }),
    .FrameData_O({\Tile_X3Y8_FrameData_O[31] ,
    \Tile_X3Y8_FrameData_O[30] ,
    \Tile_X3Y8_FrameData_O[29] ,
    \Tile_X3Y8_FrameData_O[28] ,
    \Tile_X3Y8_FrameData_O[27] ,
    \Tile_X3Y8_FrameData_O[26] ,
    \Tile_X3Y8_FrameData_O[25] ,
    \Tile_X3Y8_FrameData_O[24] ,
    \Tile_X3Y8_FrameData_O[23] ,
    \Tile_X3Y8_FrameData_O[22] ,
    \Tile_X3Y8_FrameData_O[21] ,
    \Tile_X3Y8_FrameData_O[20] ,
    \Tile_X3Y8_FrameData_O[19] ,
    \Tile_X3Y8_FrameData_O[18] ,
    \Tile_X3Y8_FrameData_O[17] ,
    \Tile_X3Y8_FrameData_O[16] ,
    \Tile_X3Y8_FrameData_O[15] ,
    \Tile_X3Y8_FrameData_O[14] ,
    \Tile_X3Y8_FrameData_O[13] ,
    \Tile_X3Y8_FrameData_O[12] ,
    \Tile_X3Y8_FrameData_O[11] ,
    \Tile_X3Y8_FrameData_O[10] ,
    \Tile_X3Y8_FrameData_O[9] ,
    \Tile_X3Y8_FrameData_O[8] ,
    \Tile_X3Y8_FrameData_O[7] ,
    \Tile_X3Y8_FrameData_O[6] ,
    \Tile_X3Y8_FrameData_O[5] ,
    \Tile_X3Y8_FrameData_O[4] ,
    \Tile_X3Y8_FrameData_O[3] ,
    \Tile_X3Y8_FrameData_O[2] ,
    \Tile_X3Y8_FrameData_O[1] ,
    \Tile_X3Y8_FrameData_O[0] }),
    .FrameStrobe({\Tile_X3Y9_FrameStrobe_O[19] ,
    \Tile_X3Y9_FrameStrobe_O[18] ,
    \Tile_X3Y9_FrameStrobe_O[17] ,
    \Tile_X3Y9_FrameStrobe_O[16] ,
    \Tile_X3Y9_FrameStrobe_O[15] ,
    \Tile_X3Y9_FrameStrobe_O[14] ,
    \Tile_X3Y9_FrameStrobe_O[13] ,
    \Tile_X3Y9_FrameStrobe_O[12] ,
    \Tile_X3Y9_FrameStrobe_O[11] ,
    \Tile_X3Y9_FrameStrobe_O[10] ,
    \Tile_X3Y9_FrameStrobe_O[9] ,
    \Tile_X3Y9_FrameStrobe_O[8] ,
    \Tile_X3Y9_FrameStrobe_O[7] ,
    \Tile_X3Y9_FrameStrobe_O[6] ,
    \Tile_X3Y9_FrameStrobe_O[5] ,
    \Tile_X3Y9_FrameStrobe_O[4] ,
    \Tile_X3Y9_FrameStrobe_O[3] ,
    \Tile_X3Y9_FrameStrobe_O[2] ,
    \Tile_X3Y9_FrameStrobe_O[1] ,
    \Tile_X3Y9_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X3Y8_FrameStrobe_O[19] ,
    \Tile_X3Y8_FrameStrobe_O[18] ,
    \Tile_X3Y8_FrameStrobe_O[17] ,
    \Tile_X3Y8_FrameStrobe_O[16] ,
    \Tile_X3Y8_FrameStrobe_O[15] ,
    \Tile_X3Y8_FrameStrobe_O[14] ,
    \Tile_X3Y8_FrameStrobe_O[13] ,
    \Tile_X3Y8_FrameStrobe_O[12] ,
    \Tile_X3Y8_FrameStrobe_O[11] ,
    \Tile_X3Y8_FrameStrobe_O[10] ,
    \Tile_X3Y8_FrameStrobe_O[9] ,
    \Tile_X3Y8_FrameStrobe_O[8] ,
    \Tile_X3Y8_FrameStrobe_O[7] ,
    \Tile_X3Y8_FrameStrobe_O[6] ,
    \Tile_X3Y8_FrameStrobe_O[5] ,
    \Tile_X3Y8_FrameStrobe_O[4] ,
    \Tile_X3Y8_FrameStrobe_O[3] ,
    \Tile_X3Y8_FrameStrobe_O[2] ,
    \Tile_X3Y8_FrameStrobe_O[1] ,
    \Tile_X3Y8_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X3Y8_N1BEG[3] ,
    \Tile_X3Y8_N1BEG[2] ,
    \Tile_X3Y8_N1BEG[1] ,
    \Tile_X3Y8_N1BEG[0] }),
    .N1END({\Tile_X3Y9_N1BEG[3] ,
    \Tile_X3Y9_N1BEG[2] ,
    \Tile_X3Y9_N1BEG[1] ,
    \Tile_X3Y9_N1BEG[0] }),
    .N2BEG({\Tile_X3Y8_N2BEG[7] ,
    \Tile_X3Y8_N2BEG[6] ,
    \Tile_X3Y8_N2BEG[5] ,
    \Tile_X3Y8_N2BEG[4] ,
    \Tile_X3Y8_N2BEG[3] ,
    \Tile_X3Y8_N2BEG[2] ,
    \Tile_X3Y8_N2BEG[1] ,
    \Tile_X3Y8_N2BEG[0] }),
    .N2BEGb({\Tile_X3Y8_N2BEGb[7] ,
    \Tile_X3Y8_N2BEGb[6] ,
    \Tile_X3Y8_N2BEGb[5] ,
    \Tile_X3Y8_N2BEGb[4] ,
    \Tile_X3Y8_N2BEGb[3] ,
    \Tile_X3Y8_N2BEGb[2] ,
    \Tile_X3Y8_N2BEGb[1] ,
    \Tile_X3Y8_N2BEGb[0] }),
    .N2END({\Tile_X3Y9_N2BEGb[7] ,
    \Tile_X3Y9_N2BEGb[6] ,
    \Tile_X3Y9_N2BEGb[5] ,
    \Tile_X3Y9_N2BEGb[4] ,
    \Tile_X3Y9_N2BEGb[3] ,
    \Tile_X3Y9_N2BEGb[2] ,
    \Tile_X3Y9_N2BEGb[1] ,
    \Tile_X3Y9_N2BEGb[0] }),
    .N2MID({\Tile_X3Y9_N2BEG[7] ,
    \Tile_X3Y9_N2BEG[6] ,
    \Tile_X3Y9_N2BEG[5] ,
    \Tile_X3Y9_N2BEG[4] ,
    \Tile_X3Y9_N2BEG[3] ,
    \Tile_X3Y9_N2BEG[2] ,
    \Tile_X3Y9_N2BEG[1] ,
    \Tile_X3Y9_N2BEG[0] }),
    .N4BEG({\Tile_X3Y8_N4BEG[15] ,
    \Tile_X3Y8_N4BEG[14] ,
    \Tile_X3Y8_N4BEG[13] ,
    \Tile_X3Y8_N4BEG[12] ,
    \Tile_X3Y8_N4BEG[11] ,
    \Tile_X3Y8_N4BEG[10] ,
    \Tile_X3Y8_N4BEG[9] ,
    \Tile_X3Y8_N4BEG[8] ,
    \Tile_X3Y8_N4BEG[7] ,
    \Tile_X3Y8_N4BEG[6] ,
    \Tile_X3Y8_N4BEG[5] ,
    \Tile_X3Y8_N4BEG[4] ,
    \Tile_X3Y8_N4BEG[3] ,
    \Tile_X3Y8_N4BEG[2] ,
    \Tile_X3Y8_N4BEG[1] ,
    \Tile_X3Y8_N4BEG[0] }),
    .N4END({\Tile_X3Y9_N4BEG[15] ,
    \Tile_X3Y9_N4BEG[14] ,
    \Tile_X3Y9_N4BEG[13] ,
    \Tile_X3Y9_N4BEG[12] ,
    \Tile_X3Y9_N4BEG[11] ,
    \Tile_X3Y9_N4BEG[10] ,
    \Tile_X3Y9_N4BEG[9] ,
    \Tile_X3Y9_N4BEG[8] ,
    \Tile_X3Y9_N4BEG[7] ,
    \Tile_X3Y9_N4BEG[6] ,
    \Tile_X3Y9_N4BEG[5] ,
    \Tile_X3Y9_N4BEG[4] ,
    \Tile_X3Y9_N4BEG[3] ,
    \Tile_X3Y9_N4BEG[2] ,
    \Tile_X3Y9_N4BEG[1] ,
    \Tile_X3Y9_N4BEG[0] }),
    .NN4BEG({\Tile_X3Y8_NN4BEG[15] ,
    \Tile_X3Y8_NN4BEG[14] ,
    \Tile_X3Y8_NN4BEG[13] ,
    \Tile_X3Y8_NN4BEG[12] ,
    \Tile_X3Y8_NN4BEG[11] ,
    \Tile_X3Y8_NN4BEG[10] ,
    \Tile_X3Y8_NN4BEG[9] ,
    \Tile_X3Y8_NN4BEG[8] ,
    \Tile_X3Y8_NN4BEG[7] ,
    \Tile_X3Y8_NN4BEG[6] ,
    \Tile_X3Y8_NN4BEG[5] ,
    \Tile_X3Y8_NN4BEG[4] ,
    \Tile_X3Y8_NN4BEG[3] ,
    \Tile_X3Y8_NN4BEG[2] ,
    \Tile_X3Y8_NN4BEG[1] ,
    \Tile_X3Y8_NN4BEG[0] }),
    .NN4END({\Tile_X3Y9_NN4BEG[15] ,
    \Tile_X3Y9_NN4BEG[14] ,
    \Tile_X3Y9_NN4BEG[13] ,
    \Tile_X3Y9_NN4BEG[12] ,
    \Tile_X3Y9_NN4BEG[11] ,
    \Tile_X3Y9_NN4BEG[10] ,
    \Tile_X3Y9_NN4BEG[9] ,
    \Tile_X3Y9_NN4BEG[8] ,
    \Tile_X3Y9_NN4BEG[7] ,
    \Tile_X3Y9_NN4BEG[6] ,
    \Tile_X3Y9_NN4BEG[5] ,
    \Tile_X3Y9_NN4BEG[4] ,
    \Tile_X3Y9_NN4BEG[3] ,
    \Tile_X3Y9_NN4BEG[2] ,
    \Tile_X3Y9_NN4BEG[1] ,
    \Tile_X3Y9_NN4BEG[0] }),
    .S1BEG({\Tile_X3Y8_S1BEG[3] ,
    \Tile_X3Y8_S1BEG[2] ,
    \Tile_X3Y8_S1BEG[1] ,
    \Tile_X3Y8_S1BEG[0] }),
    .S1END({\Tile_X3Y7_S1BEG[3] ,
    \Tile_X3Y7_S1BEG[2] ,
    \Tile_X3Y7_S1BEG[1] ,
    \Tile_X3Y7_S1BEG[0] }),
    .S2BEG({\Tile_X3Y8_S2BEG[7] ,
    \Tile_X3Y8_S2BEG[6] ,
    \Tile_X3Y8_S2BEG[5] ,
    \Tile_X3Y8_S2BEG[4] ,
    \Tile_X3Y8_S2BEG[3] ,
    \Tile_X3Y8_S2BEG[2] ,
    \Tile_X3Y8_S2BEG[1] ,
    \Tile_X3Y8_S2BEG[0] }),
    .S2BEGb({\Tile_X3Y8_S2BEGb[7] ,
    \Tile_X3Y8_S2BEGb[6] ,
    \Tile_X3Y8_S2BEGb[5] ,
    \Tile_X3Y8_S2BEGb[4] ,
    \Tile_X3Y8_S2BEGb[3] ,
    \Tile_X3Y8_S2BEGb[2] ,
    \Tile_X3Y8_S2BEGb[1] ,
    \Tile_X3Y8_S2BEGb[0] }),
    .S2END({\Tile_X3Y7_S2BEGb[7] ,
    \Tile_X3Y7_S2BEGb[6] ,
    \Tile_X3Y7_S2BEGb[5] ,
    \Tile_X3Y7_S2BEGb[4] ,
    \Tile_X3Y7_S2BEGb[3] ,
    \Tile_X3Y7_S2BEGb[2] ,
    \Tile_X3Y7_S2BEGb[1] ,
    \Tile_X3Y7_S2BEGb[0] }),
    .S2MID({\Tile_X3Y7_S2BEG[7] ,
    \Tile_X3Y7_S2BEG[6] ,
    \Tile_X3Y7_S2BEG[5] ,
    \Tile_X3Y7_S2BEG[4] ,
    \Tile_X3Y7_S2BEG[3] ,
    \Tile_X3Y7_S2BEG[2] ,
    \Tile_X3Y7_S2BEG[1] ,
    \Tile_X3Y7_S2BEG[0] }),
    .S4BEG({\Tile_X3Y8_S4BEG[15] ,
    \Tile_X3Y8_S4BEG[14] ,
    \Tile_X3Y8_S4BEG[13] ,
    \Tile_X3Y8_S4BEG[12] ,
    \Tile_X3Y8_S4BEG[11] ,
    \Tile_X3Y8_S4BEG[10] ,
    \Tile_X3Y8_S4BEG[9] ,
    \Tile_X3Y8_S4BEG[8] ,
    \Tile_X3Y8_S4BEG[7] ,
    \Tile_X3Y8_S4BEG[6] ,
    \Tile_X3Y8_S4BEG[5] ,
    \Tile_X3Y8_S4BEG[4] ,
    \Tile_X3Y8_S4BEG[3] ,
    \Tile_X3Y8_S4BEG[2] ,
    \Tile_X3Y8_S4BEG[1] ,
    \Tile_X3Y8_S4BEG[0] }),
    .S4END({\Tile_X3Y7_S4BEG[15] ,
    \Tile_X3Y7_S4BEG[14] ,
    \Tile_X3Y7_S4BEG[13] ,
    \Tile_X3Y7_S4BEG[12] ,
    \Tile_X3Y7_S4BEG[11] ,
    \Tile_X3Y7_S4BEG[10] ,
    \Tile_X3Y7_S4BEG[9] ,
    \Tile_X3Y7_S4BEG[8] ,
    \Tile_X3Y7_S4BEG[7] ,
    \Tile_X3Y7_S4BEG[6] ,
    \Tile_X3Y7_S4BEG[5] ,
    \Tile_X3Y7_S4BEG[4] ,
    \Tile_X3Y7_S4BEG[3] ,
    \Tile_X3Y7_S4BEG[2] ,
    \Tile_X3Y7_S4BEG[1] ,
    \Tile_X3Y7_S4BEG[0] }),
    .SS4BEG({\Tile_X3Y8_SS4BEG[15] ,
    \Tile_X3Y8_SS4BEG[14] ,
    \Tile_X3Y8_SS4BEG[13] ,
    \Tile_X3Y8_SS4BEG[12] ,
    \Tile_X3Y8_SS4BEG[11] ,
    \Tile_X3Y8_SS4BEG[10] ,
    \Tile_X3Y8_SS4BEG[9] ,
    \Tile_X3Y8_SS4BEG[8] ,
    \Tile_X3Y8_SS4BEG[7] ,
    \Tile_X3Y8_SS4BEG[6] ,
    \Tile_X3Y8_SS4BEG[5] ,
    \Tile_X3Y8_SS4BEG[4] ,
    \Tile_X3Y8_SS4BEG[3] ,
    \Tile_X3Y8_SS4BEG[2] ,
    \Tile_X3Y8_SS4BEG[1] ,
    \Tile_X3Y8_SS4BEG[0] }),
    .SS4END({\Tile_X3Y7_SS4BEG[15] ,
    \Tile_X3Y7_SS4BEG[14] ,
    \Tile_X3Y7_SS4BEG[13] ,
    \Tile_X3Y7_SS4BEG[12] ,
    \Tile_X3Y7_SS4BEG[11] ,
    \Tile_X3Y7_SS4BEG[10] ,
    \Tile_X3Y7_SS4BEG[9] ,
    \Tile_X3Y7_SS4BEG[8] ,
    \Tile_X3Y7_SS4BEG[7] ,
    \Tile_X3Y7_SS4BEG[6] ,
    \Tile_X3Y7_SS4BEG[5] ,
    \Tile_X3Y7_SS4BEG[4] ,
    \Tile_X3Y7_SS4BEG[3] ,
    \Tile_X3Y7_SS4BEG[2] ,
    \Tile_X3Y7_SS4BEG[1] ,
    \Tile_X3Y7_SS4BEG[0] }),
    .W1BEG({\Tile_X3Y8_W1BEG[3] ,
    \Tile_X3Y8_W1BEG[2] ,
    \Tile_X3Y8_W1BEG[1] ,
    \Tile_X3Y8_W1BEG[0] }),
    .W1END({\Tile_X4Y8_W1BEG[3] ,
    \Tile_X4Y8_W1BEG[2] ,
    \Tile_X4Y8_W1BEG[1] ,
    \Tile_X4Y8_W1BEG[0] }),
    .W2BEG({\Tile_X3Y8_W2BEG[7] ,
    \Tile_X3Y8_W2BEG[6] ,
    \Tile_X3Y8_W2BEG[5] ,
    \Tile_X3Y8_W2BEG[4] ,
    \Tile_X3Y8_W2BEG[3] ,
    \Tile_X3Y8_W2BEG[2] ,
    \Tile_X3Y8_W2BEG[1] ,
    \Tile_X3Y8_W2BEG[0] }),
    .W2BEGb({\Tile_X3Y8_W2BEGb[7] ,
    \Tile_X3Y8_W2BEGb[6] ,
    \Tile_X3Y8_W2BEGb[5] ,
    \Tile_X3Y8_W2BEGb[4] ,
    \Tile_X3Y8_W2BEGb[3] ,
    \Tile_X3Y8_W2BEGb[2] ,
    \Tile_X3Y8_W2BEGb[1] ,
    \Tile_X3Y8_W2BEGb[0] }),
    .W2END({\Tile_X4Y8_W2BEGb[7] ,
    \Tile_X4Y8_W2BEGb[6] ,
    \Tile_X4Y8_W2BEGb[5] ,
    \Tile_X4Y8_W2BEGb[4] ,
    \Tile_X4Y8_W2BEGb[3] ,
    \Tile_X4Y8_W2BEGb[2] ,
    \Tile_X4Y8_W2BEGb[1] ,
    \Tile_X4Y8_W2BEGb[0] }),
    .W2MID({\Tile_X4Y8_W2BEG[7] ,
    \Tile_X4Y8_W2BEG[6] ,
    \Tile_X4Y8_W2BEG[5] ,
    \Tile_X4Y8_W2BEG[4] ,
    \Tile_X4Y8_W2BEG[3] ,
    \Tile_X4Y8_W2BEG[2] ,
    \Tile_X4Y8_W2BEG[1] ,
    \Tile_X4Y8_W2BEG[0] }),
    .W6BEG({\Tile_X3Y8_W6BEG[11] ,
    \Tile_X3Y8_W6BEG[10] ,
    \Tile_X3Y8_W6BEG[9] ,
    \Tile_X3Y8_W6BEG[8] ,
    \Tile_X3Y8_W6BEG[7] ,
    \Tile_X3Y8_W6BEG[6] ,
    \Tile_X3Y8_W6BEG[5] ,
    \Tile_X3Y8_W6BEG[4] ,
    \Tile_X3Y8_W6BEG[3] ,
    \Tile_X3Y8_W6BEG[2] ,
    \Tile_X3Y8_W6BEG[1] ,
    \Tile_X3Y8_W6BEG[0] }),
    .W6END({\Tile_X4Y8_W6BEG[11] ,
    \Tile_X4Y8_W6BEG[10] ,
    \Tile_X4Y8_W6BEG[9] ,
    \Tile_X4Y8_W6BEG[8] ,
    \Tile_X4Y8_W6BEG[7] ,
    \Tile_X4Y8_W6BEG[6] ,
    \Tile_X4Y8_W6BEG[5] ,
    \Tile_X4Y8_W6BEG[4] ,
    \Tile_X4Y8_W6BEG[3] ,
    \Tile_X4Y8_W6BEG[2] ,
    \Tile_X4Y8_W6BEG[1] ,
    \Tile_X4Y8_W6BEG[0] }),
    .WW4BEG({\Tile_X3Y8_WW4BEG[15] ,
    \Tile_X3Y8_WW4BEG[14] ,
    \Tile_X3Y8_WW4BEG[13] ,
    \Tile_X3Y8_WW4BEG[12] ,
    \Tile_X3Y8_WW4BEG[11] ,
    \Tile_X3Y8_WW4BEG[10] ,
    \Tile_X3Y8_WW4BEG[9] ,
    \Tile_X3Y8_WW4BEG[8] ,
    \Tile_X3Y8_WW4BEG[7] ,
    \Tile_X3Y8_WW4BEG[6] ,
    \Tile_X3Y8_WW4BEG[5] ,
    \Tile_X3Y8_WW4BEG[4] ,
    \Tile_X3Y8_WW4BEG[3] ,
    \Tile_X3Y8_WW4BEG[2] ,
    \Tile_X3Y8_WW4BEG[1] ,
    \Tile_X3Y8_WW4BEG[0] }),
    .WW4END({\Tile_X4Y8_WW4BEG[15] ,
    \Tile_X4Y8_WW4BEG[14] ,
    \Tile_X4Y8_WW4BEG[13] ,
    \Tile_X4Y8_WW4BEG[12] ,
    \Tile_X4Y8_WW4BEG[11] ,
    \Tile_X4Y8_WW4BEG[10] ,
    \Tile_X4Y8_WW4BEG[9] ,
    \Tile_X4Y8_WW4BEG[8] ,
    \Tile_X4Y8_WW4BEG[7] ,
    \Tile_X4Y8_WW4BEG[6] ,
    \Tile_X4Y8_WW4BEG[5] ,
    \Tile_X4Y8_WW4BEG[4] ,
    \Tile_X4Y8_WW4BEG[3] ,
    \Tile_X4Y8_WW4BEG[2] ,
    \Tile_X4Y8_WW4BEG[1] ,
    \Tile_X4Y8_WW4BEG[0] }));
 S_IO4 Tile_X3Y9_S_IO4 (.A_I_top(Tile_X3Y9_A_I_top),
    .A_O_top(Tile_X3Y9_A_O_top),
    .A_T_top(Tile_X3Y9_A_T_top),
    .B_I_top(Tile_X3Y9_B_I_top),
    .B_O_top(Tile_X3Y9_B_O_top),
    .B_T_top(Tile_X3Y9_B_T_top),
    .C_I_top(Tile_X3Y9_C_I_top),
    .C_O_top(Tile_X3Y9_C_O_top),
    .C_T_top(Tile_X3Y9_C_T_top),
    .Co(Tile_X3Y9_Co),
    .D_I_top(Tile_X3Y9_D_I_top),
    .D_O_top(Tile_X3Y9_D_O_top),
    .D_T_top(Tile_X3Y9_D_T_top),
    .UserCLK(UserCLK),
    .UserCLKo(Tile_X3Y9_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .FrameData({\Tile_X2Y9_FrameData_O[31] ,
    \Tile_X2Y9_FrameData_O[30] ,
    \Tile_X2Y9_FrameData_O[29] ,
    \Tile_X2Y9_FrameData_O[28] ,
    \Tile_X2Y9_FrameData_O[27] ,
    \Tile_X2Y9_FrameData_O[26] ,
    \Tile_X2Y9_FrameData_O[25] ,
    \Tile_X2Y9_FrameData_O[24] ,
    \Tile_X2Y9_FrameData_O[23] ,
    \Tile_X2Y9_FrameData_O[22] ,
    \Tile_X2Y9_FrameData_O[21] ,
    \Tile_X2Y9_FrameData_O[20] ,
    \Tile_X2Y9_FrameData_O[19] ,
    \Tile_X2Y9_FrameData_O[18] ,
    \Tile_X2Y9_FrameData_O[17] ,
    \Tile_X2Y9_FrameData_O[16] ,
    \Tile_X2Y9_FrameData_O[15] ,
    \Tile_X2Y9_FrameData_O[14] ,
    \Tile_X2Y9_FrameData_O[13] ,
    \Tile_X2Y9_FrameData_O[12] ,
    \Tile_X2Y9_FrameData_O[11] ,
    \Tile_X2Y9_FrameData_O[10] ,
    \Tile_X2Y9_FrameData_O[9] ,
    \Tile_X2Y9_FrameData_O[8] ,
    \Tile_X2Y9_FrameData_O[7] ,
    \Tile_X2Y9_FrameData_O[6] ,
    \Tile_X2Y9_FrameData_O[5] ,
    \Tile_X2Y9_FrameData_O[4] ,
    \Tile_X2Y9_FrameData_O[3] ,
    \Tile_X2Y9_FrameData_O[2] ,
    \Tile_X2Y9_FrameData_O[1] ,
    \Tile_X2Y9_FrameData_O[0] }),
    .FrameData_O({\Tile_X3Y9_FrameData_O[31] ,
    \Tile_X3Y9_FrameData_O[30] ,
    \Tile_X3Y9_FrameData_O[29] ,
    \Tile_X3Y9_FrameData_O[28] ,
    \Tile_X3Y9_FrameData_O[27] ,
    \Tile_X3Y9_FrameData_O[26] ,
    \Tile_X3Y9_FrameData_O[25] ,
    \Tile_X3Y9_FrameData_O[24] ,
    \Tile_X3Y9_FrameData_O[23] ,
    \Tile_X3Y9_FrameData_O[22] ,
    \Tile_X3Y9_FrameData_O[21] ,
    \Tile_X3Y9_FrameData_O[20] ,
    \Tile_X3Y9_FrameData_O[19] ,
    \Tile_X3Y9_FrameData_O[18] ,
    \Tile_X3Y9_FrameData_O[17] ,
    \Tile_X3Y9_FrameData_O[16] ,
    \Tile_X3Y9_FrameData_O[15] ,
    \Tile_X3Y9_FrameData_O[14] ,
    \Tile_X3Y9_FrameData_O[13] ,
    \Tile_X3Y9_FrameData_O[12] ,
    \Tile_X3Y9_FrameData_O[11] ,
    \Tile_X3Y9_FrameData_O[10] ,
    \Tile_X3Y9_FrameData_O[9] ,
    \Tile_X3Y9_FrameData_O[8] ,
    \Tile_X3Y9_FrameData_O[7] ,
    \Tile_X3Y9_FrameData_O[6] ,
    \Tile_X3Y9_FrameData_O[5] ,
    \Tile_X3Y9_FrameData_O[4] ,
    \Tile_X3Y9_FrameData_O[3] ,
    \Tile_X3Y9_FrameData_O[2] ,
    \Tile_X3Y9_FrameData_O[1] ,
    \Tile_X3Y9_FrameData_O[0] }),
    .FrameStrobe({FrameStrobe[79],
    FrameStrobe[78],
    FrameStrobe[77],
    FrameStrobe[76],
    FrameStrobe[75],
    FrameStrobe[74],
    FrameStrobe[73],
    FrameStrobe[72],
    FrameStrobe[71],
    FrameStrobe[70],
    FrameStrobe[69],
    FrameStrobe[68],
    FrameStrobe[67],
    FrameStrobe[66],
    FrameStrobe[65],
    FrameStrobe[64],
    FrameStrobe[63],
    FrameStrobe[62],
    FrameStrobe[61],
    FrameStrobe[60]}),
    .FrameStrobe_O({\Tile_X3Y9_FrameStrobe_O[19] ,
    \Tile_X3Y9_FrameStrobe_O[18] ,
    \Tile_X3Y9_FrameStrobe_O[17] ,
    \Tile_X3Y9_FrameStrobe_O[16] ,
    \Tile_X3Y9_FrameStrobe_O[15] ,
    \Tile_X3Y9_FrameStrobe_O[14] ,
    \Tile_X3Y9_FrameStrobe_O[13] ,
    \Tile_X3Y9_FrameStrobe_O[12] ,
    \Tile_X3Y9_FrameStrobe_O[11] ,
    \Tile_X3Y9_FrameStrobe_O[10] ,
    \Tile_X3Y9_FrameStrobe_O[9] ,
    \Tile_X3Y9_FrameStrobe_O[8] ,
    \Tile_X3Y9_FrameStrobe_O[7] ,
    \Tile_X3Y9_FrameStrobe_O[6] ,
    \Tile_X3Y9_FrameStrobe_O[5] ,
    \Tile_X3Y9_FrameStrobe_O[4] ,
    \Tile_X3Y9_FrameStrobe_O[3] ,
    \Tile_X3Y9_FrameStrobe_O[2] ,
    \Tile_X3Y9_FrameStrobe_O[1] ,
    \Tile_X3Y9_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X3Y9_N1BEG[3] ,
    \Tile_X3Y9_N1BEG[2] ,
    \Tile_X3Y9_N1BEG[1] ,
    \Tile_X3Y9_N1BEG[0] }),
    .N2BEG({\Tile_X3Y9_N2BEG[7] ,
    \Tile_X3Y9_N2BEG[6] ,
    \Tile_X3Y9_N2BEG[5] ,
    \Tile_X3Y9_N2BEG[4] ,
    \Tile_X3Y9_N2BEG[3] ,
    \Tile_X3Y9_N2BEG[2] ,
    \Tile_X3Y9_N2BEG[1] ,
    \Tile_X3Y9_N2BEG[0] }),
    .N2BEGb({\Tile_X3Y9_N2BEGb[7] ,
    \Tile_X3Y9_N2BEGb[6] ,
    \Tile_X3Y9_N2BEGb[5] ,
    \Tile_X3Y9_N2BEGb[4] ,
    \Tile_X3Y9_N2BEGb[3] ,
    \Tile_X3Y9_N2BEGb[2] ,
    \Tile_X3Y9_N2BEGb[1] ,
    \Tile_X3Y9_N2BEGb[0] }),
    .N4BEG({\Tile_X3Y9_N4BEG[15] ,
    \Tile_X3Y9_N4BEG[14] ,
    \Tile_X3Y9_N4BEG[13] ,
    \Tile_X3Y9_N4BEG[12] ,
    \Tile_X3Y9_N4BEG[11] ,
    \Tile_X3Y9_N4BEG[10] ,
    \Tile_X3Y9_N4BEG[9] ,
    \Tile_X3Y9_N4BEG[8] ,
    \Tile_X3Y9_N4BEG[7] ,
    \Tile_X3Y9_N4BEG[6] ,
    \Tile_X3Y9_N4BEG[5] ,
    \Tile_X3Y9_N4BEG[4] ,
    \Tile_X3Y9_N4BEG[3] ,
    \Tile_X3Y9_N4BEG[2] ,
    \Tile_X3Y9_N4BEG[1] ,
    \Tile_X3Y9_N4BEG[0] }),
    .NN4BEG({\Tile_X3Y9_NN4BEG[15] ,
    \Tile_X3Y9_NN4BEG[14] ,
    \Tile_X3Y9_NN4BEG[13] ,
    \Tile_X3Y9_NN4BEG[12] ,
    \Tile_X3Y9_NN4BEG[11] ,
    \Tile_X3Y9_NN4BEG[10] ,
    \Tile_X3Y9_NN4BEG[9] ,
    \Tile_X3Y9_NN4BEG[8] ,
    \Tile_X3Y9_NN4BEG[7] ,
    \Tile_X3Y9_NN4BEG[6] ,
    \Tile_X3Y9_NN4BEG[5] ,
    \Tile_X3Y9_NN4BEG[4] ,
    \Tile_X3Y9_NN4BEG[3] ,
    \Tile_X3Y9_NN4BEG[2] ,
    \Tile_X3Y9_NN4BEG[1] ,
    \Tile_X3Y9_NN4BEG[0] }),
    .S1END({\Tile_X3Y8_S1BEG[3] ,
    \Tile_X3Y8_S1BEG[2] ,
    \Tile_X3Y8_S1BEG[1] ,
    \Tile_X3Y8_S1BEG[0] }),
    .S2END({\Tile_X3Y8_S2BEGb[7] ,
    \Tile_X3Y8_S2BEGb[6] ,
    \Tile_X3Y8_S2BEGb[5] ,
    \Tile_X3Y8_S2BEGb[4] ,
    \Tile_X3Y8_S2BEGb[3] ,
    \Tile_X3Y8_S2BEGb[2] ,
    \Tile_X3Y8_S2BEGb[1] ,
    \Tile_X3Y8_S2BEGb[0] }),
    .S2MID({\Tile_X3Y8_S2BEG[7] ,
    \Tile_X3Y8_S2BEG[6] ,
    \Tile_X3Y8_S2BEG[5] ,
    \Tile_X3Y8_S2BEG[4] ,
    \Tile_X3Y8_S2BEG[3] ,
    \Tile_X3Y8_S2BEG[2] ,
    \Tile_X3Y8_S2BEG[1] ,
    \Tile_X3Y8_S2BEG[0] }),
    .S4END({\Tile_X3Y8_S4BEG[15] ,
    \Tile_X3Y8_S4BEG[14] ,
    \Tile_X3Y8_S4BEG[13] ,
    \Tile_X3Y8_S4BEG[12] ,
    \Tile_X3Y8_S4BEG[11] ,
    \Tile_X3Y8_S4BEG[10] ,
    \Tile_X3Y8_S4BEG[9] ,
    \Tile_X3Y8_S4BEG[8] ,
    \Tile_X3Y8_S4BEG[7] ,
    \Tile_X3Y8_S4BEG[6] ,
    \Tile_X3Y8_S4BEG[5] ,
    \Tile_X3Y8_S4BEG[4] ,
    \Tile_X3Y8_S4BEG[3] ,
    \Tile_X3Y8_S4BEG[2] ,
    \Tile_X3Y8_S4BEG[1] ,
    \Tile_X3Y8_S4BEG[0] }),
    .SS4END({\Tile_X3Y8_SS4BEG[15] ,
    \Tile_X3Y8_SS4BEG[14] ,
    \Tile_X3Y8_SS4BEG[13] ,
    \Tile_X3Y8_SS4BEG[12] ,
    \Tile_X3Y8_SS4BEG[11] ,
    \Tile_X3Y8_SS4BEG[10] ,
    \Tile_X3Y8_SS4BEG[9] ,
    \Tile_X3Y8_SS4BEG[8] ,
    \Tile_X3Y8_SS4BEG[7] ,
    \Tile_X3Y8_SS4BEG[6] ,
    \Tile_X3Y8_SS4BEG[5] ,
    \Tile_X3Y8_SS4BEG[4] ,
    \Tile_X3Y8_SS4BEG[3] ,
    \Tile_X3Y8_SS4BEG[2] ,
    \Tile_X3Y8_SS4BEG[1] ,
    \Tile_X3Y8_SS4BEG[0] }));
 N_IO4 Tile_X4Y0_N_IO4 (.A_I_top(Tile_X4Y0_A_I_top),
    .A_O_top(Tile_X4Y0_A_O_top),
    .A_T_top(Tile_X4Y0_A_T_top),
    .B_I_top(Tile_X4Y0_B_I_top),
    .B_O_top(Tile_X4Y0_B_O_top),
    .B_T_top(Tile_X4Y0_B_T_top),
    .C_I_top(Tile_X4Y0_C_I_top),
    .C_O_top(Tile_X4Y0_C_O_top),
    .C_T_top(Tile_X4Y0_C_T_top),
    .Ci(Tile_X4Y1_Co),
    .D_I_top(Tile_X4Y0_D_I_top),
    .D_O_top(Tile_X4Y0_D_O_top),
    .D_T_top(Tile_X4Y0_D_T_top),
    .UserCLK(Tile_X4Y1_UserCLKo),
    .UserCLKo(Tile_X4Y0_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .FrameData({\Tile_X3Y0_FrameData_O[31] ,
    \Tile_X3Y0_FrameData_O[30] ,
    \Tile_X3Y0_FrameData_O[29] ,
    \Tile_X3Y0_FrameData_O[28] ,
    \Tile_X3Y0_FrameData_O[27] ,
    \Tile_X3Y0_FrameData_O[26] ,
    \Tile_X3Y0_FrameData_O[25] ,
    \Tile_X3Y0_FrameData_O[24] ,
    \Tile_X3Y0_FrameData_O[23] ,
    \Tile_X3Y0_FrameData_O[22] ,
    \Tile_X3Y0_FrameData_O[21] ,
    \Tile_X3Y0_FrameData_O[20] ,
    \Tile_X3Y0_FrameData_O[19] ,
    \Tile_X3Y0_FrameData_O[18] ,
    \Tile_X3Y0_FrameData_O[17] ,
    \Tile_X3Y0_FrameData_O[16] ,
    \Tile_X3Y0_FrameData_O[15] ,
    \Tile_X3Y0_FrameData_O[14] ,
    \Tile_X3Y0_FrameData_O[13] ,
    \Tile_X3Y0_FrameData_O[12] ,
    \Tile_X3Y0_FrameData_O[11] ,
    \Tile_X3Y0_FrameData_O[10] ,
    \Tile_X3Y0_FrameData_O[9] ,
    \Tile_X3Y0_FrameData_O[8] ,
    \Tile_X3Y0_FrameData_O[7] ,
    \Tile_X3Y0_FrameData_O[6] ,
    \Tile_X3Y0_FrameData_O[5] ,
    \Tile_X3Y0_FrameData_O[4] ,
    \Tile_X3Y0_FrameData_O[3] ,
    \Tile_X3Y0_FrameData_O[2] ,
    \Tile_X3Y0_FrameData_O[1] ,
    \Tile_X3Y0_FrameData_O[0] }),
    .FrameData_O({\Tile_X4Y0_FrameData_O[31] ,
    \Tile_X4Y0_FrameData_O[30] ,
    \Tile_X4Y0_FrameData_O[29] ,
    \Tile_X4Y0_FrameData_O[28] ,
    \Tile_X4Y0_FrameData_O[27] ,
    \Tile_X4Y0_FrameData_O[26] ,
    \Tile_X4Y0_FrameData_O[25] ,
    \Tile_X4Y0_FrameData_O[24] ,
    \Tile_X4Y0_FrameData_O[23] ,
    \Tile_X4Y0_FrameData_O[22] ,
    \Tile_X4Y0_FrameData_O[21] ,
    \Tile_X4Y0_FrameData_O[20] ,
    \Tile_X4Y0_FrameData_O[19] ,
    \Tile_X4Y0_FrameData_O[18] ,
    \Tile_X4Y0_FrameData_O[17] ,
    \Tile_X4Y0_FrameData_O[16] ,
    \Tile_X4Y0_FrameData_O[15] ,
    \Tile_X4Y0_FrameData_O[14] ,
    \Tile_X4Y0_FrameData_O[13] ,
    \Tile_X4Y0_FrameData_O[12] ,
    \Tile_X4Y0_FrameData_O[11] ,
    \Tile_X4Y0_FrameData_O[10] ,
    \Tile_X4Y0_FrameData_O[9] ,
    \Tile_X4Y0_FrameData_O[8] ,
    \Tile_X4Y0_FrameData_O[7] ,
    \Tile_X4Y0_FrameData_O[6] ,
    \Tile_X4Y0_FrameData_O[5] ,
    \Tile_X4Y0_FrameData_O[4] ,
    \Tile_X4Y0_FrameData_O[3] ,
    \Tile_X4Y0_FrameData_O[2] ,
    \Tile_X4Y0_FrameData_O[1] ,
    \Tile_X4Y0_FrameData_O[0] }),
    .FrameStrobe({\Tile_X4Y1_FrameStrobe_O[19] ,
    \Tile_X4Y1_FrameStrobe_O[18] ,
    \Tile_X4Y1_FrameStrobe_O[17] ,
    \Tile_X4Y1_FrameStrobe_O[16] ,
    \Tile_X4Y1_FrameStrobe_O[15] ,
    \Tile_X4Y1_FrameStrobe_O[14] ,
    \Tile_X4Y1_FrameStrobe_O[13] ,
    \Tile_X4Y1_FrameStrobe_O[12] ,
    \Tile_X4Y1_FrameStrobe_O[11] ,
    \Tile_X4Y1_FrameStrobe_O[10] ,
    \Tile_X4Y1_FrameStrobe_O[9] ,
    \Tile_X4Y1_FrameStrobe_O[8] ,
    \Tile_X4Y1_FrameStrobe_O[7] ,
    \Tile_X4Y1_FrameStrobe_O[6] ,
    \Tile_X4Y1_FrameStrobe_O[5] ,
    \Tile_X4Y1_FrameStrobe_O[4] ,
    \Tile_X4Y1_FrameStrobe_O[3] ,
    \Tile_X4Y1_FrameStrobe_O[2] ,
    \Tile_X4Y1_FrameStrobe_O[1] ,
    \Tile_X4Y1_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X4Y0_FrameStrobe_O[19] ,
    \Tile_X4Y0_FrameStrobe_O[18] ,
    \Tile_X4Y0_FrameStrobe_O[17] ,
    \Tile_X4Y0_FrameStrobe_O[16] ,
    \Tile_X4Y0_FrameStrobe_O[15] ,
    \Tile_X4Y0_FrameStrobe_O[14] ,
    \Tile_X4Y0_FrameStrobe_O[13] ,
    \Tile_X4Y0_FrameStrobe_O[12] ,
    \Tile_X4Y0_FrameStrobe_O[11] ,
    \Tile_X4Y0_FrameStrobe_O[10] ,
    \Tile_X4Y0_FrameStrobe_O[9] ,
    \Tile_X4Y0_FrameStrobe_O[8] ,
    \Tile_X4Y0_FrameStrobe_O[7] ,
    \Tile_X4Y0_FrameStrobe_O[6] ,
    \Tile_X4Y0_FrameStrobe_O[5] ,
    \Tile_X4Y0_FrameStrobe_O[4] ,
    \Tile_X4Y0_FrameStrobe_O[3] ,
    \Tile_X4Y0_FrameStrobe_O[2] ,
    \Tile_X4Y0_FrameStrobe_O[1] ,
    \Tile_X4Y0_FrameStrobe_O[0] }),
    .N1END({\Tile_X4Y1_N1BEG[3] ,
    \Tile_X4Y1_N1BEG[2] ,
    \Tile_X4Y1_N1BEG[1] ,
    \Tile_X4Y1_N1BEG[0] }),
    .N2END({\Tile_X4Y1_N2BEGb[7] ,
    \Tile_X4Y1_N2BEGb[6] ,
    \Tile_X4Y1_N2BEGb[5] ,
    \Tile_X4Y1_N2BEGb[4] ,
    \Tile_X4Y1_N2BEGb[3] ,
    \Tile_X4Y1_N2BEGb[2] ,
    \Tile_X4Y1_N2BEGb[1] ,
    \Tile_X4Y1_N2BEGb[0] }),
    .N2MID({\Tile_X4Y1_N2BEG[7] ,
    \Tile_X4Y1_N2BEG[6] ,
    \Tile_X4Y1_N2BEG[5] ,
    \Tile_X4Y1_N2BEG[4] ,
    \Tile_X4Y1_N2BEG[3] ,
    \Tile_X4Y1_N2BEG[2] ,
    \Tile_X4Y1_N2BEG[1] ,
    \Tile_X4Y1_N2BEG[0] }),
    .N4END({\Tile_X4Y1_N4BEG[15] ,
    \Tile_X4Y1_N4BEG[14] ,
    \Tile_X4Y1_N4BEG[13] ,
    \Tile_X4Y1_N4BEG[12] ,
    \Tile_X4Y1_N4BEG[11] ,
    \Tile_X4Y1_N4BEG[10] ,
    \Tile_X4Y1_N4BEG[9] ,
    \Tile_X4Y1_N4BEG[8] ,
    \Tile_X4Y1_N4BEG[7] ,
    \Tile_X4Y1_N4BEG[6] ,
    \Tile_X4Y1_N4BEG[5] ,
    \Tile_X4Y1_N4BEG[4] ,
    \Tile_X4Y1_N4BEG[3] ,
    \Tile_X4Y1_N4BEG[2] ,
    \Tile_X4Y1_N4BEG[1] ,
    \Tile_X4Y1_N4BEG[0] }),
    .NN4END({\Tile_X4Y1_NN4BEG[15] ,
    \Tile_X4Y1_NN4BEG[14] ,
    \Tile_X4Y1_NN4BEG[13] ,
    \Tile_X4Y1_NN4BEG[12] ,
    \Tile_X4Y1_NN4BEG[11] ,
    \Tile_X4Y1_NN4BEG[10] ,
    \Tile_X4Y1_NN4BEG[9] ,
    \Tile_X4Y1_NN4BEG[8] ,
    \Tile_X4Y1_NN4BEG[7] ,
    \Tile_X4Y1_NN4BEG[6] ,
    \Tile_X4Y1_NN4BEG[5] ,
    \Tile_X4Y1_NN4BEG[4] ,
    \Tile_X4Y1_NN4BEG[3] ,
    \Tile_X4Y1_NN4BEG[2] ,
    \Tile_X4Y1_NN4BEG[1] ,
    \Tile_X4Y1_NN4BEG[0] }),
    .S1BEG({\Tile_X4Y0_S1BEG[3] ,
    \Tile_X4Y0_S1BEG[2] ,
    \Tile_X4Y0_S1BEG[1] ,
    \Tile_X4Y0_S1BEG[0] }),
    .S2BEG({\Tile_X4Y0_S2BEG[7] ,
    \Tile_X4Y0_S2BEG[6] ,
    \Tile_X4Y0_S2BEG[5] ,
    \Tile_X4Y0_S2BEG[4] ,
    \Tile_X4Y0_S2BEG[3] ,
    \Tile_X4Y0_S2BEG[2] ,
    \Tile_X4Y0_S2BEG[1] ,
    \Tile_X4Y0_S2BEG[0] }),
    .S2BEGb({\Tile_X4Y0_S2BEGb[7] ,
    \Tile_X4Y0_S2BEGb[6] ,
    \Tile_X4Y0_S2BEGb[5] ,
    \Tile_X4Y0_S2BEGb[4] ,
    \Tile_X4Y0_S2BEGb[3] ,
    \Tile_X4Y0_S2BEGb[2] ,
    \Tile_X4Y0_S2BEGb[1] ,
    \Tile_X4Y0_S2BEGb[0] }),
    .S4BEG({\Tile_X4Y0_S4BEG[15] ,
    \Tile_X4Y0_S4BEG[14] ,
    \Tile_X4Y0_S4BEG[13] ,
    \Tile_X4Y0_S4BEG[12] ,
    \Tile_X4Y0_S4BEG[11] ,
    \Tile_X4Y0_S4BEG[10] ,
    \Tile_X4Y0_S4BEG[9] ,
    \Tile_X4Y0_S4BEG[8] ,
    \Tile_X4Y0_S4BEG[7] ,
    \Tile_X4Y0_S4BEG[6] ,
    \Tile_X4Y0_S4BEG[5] ,
    \Tile_X4Y0_S4BEG[4] ,
    \Tile_X4Y0_S4BEG[3] ,
    \Tile_X4Y0_S4BEG[2] ,
    \Tile_X4Y0_S4BEG[1] ,
    \Tile_X4Y0_S4BEG[0] }),
    .SS4BEG({\Tile_X4Y0_SS4BEG[15] ,
    \Tile_X4Y0_SS4BEG[14] ,
    \Tile_X4Y0_SS4BEG[13] ,
    \Tile_X4Y0_SS4BEG[12] ,
    \Tile_X4Y0_SS4BEG[11] ,
    \Tile_X4Y0_SS4BEG[10] ,
    \Tile_X4Y0_SS4BEG[9] ,
    \Tile_X4Y0_SS4BEG[8] ,
    \Tile_X4Y0_SS4BEG[7] ,
    \Tile_X4Y0_SS4BEG[6] ,
    \Tile_X4Y0_SS4BEG[5] ,
    \Tile_X4Y0_SS4BEG[4] ,
    \Tile_X4Y0_SS4BEG[3] ,
    \Tile_X4Y0_SS4BEG[2] ,
    \Tile_X4Y0_SS4BEG[1] ,
    \Tile_X4Y0_SS4BEG[0] }));
 LUT4AB Tile_X4Y1_LUT4AB (.Ci(Tile_X4Y2_Co),
    .Co(Tile_X4Y1_Co),
    .UserCLK(Tile_X4Y2_UserCLKo),
    .UserCLKo(Tile_X4Y1_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X4Y1_E1BEG[3] ,
    \Tile_X4Y1_E1BEG[2] ,
    \Tile_X4Y1_E1BEG[1] ,
    \Tile_X4Y1_E1BEG[0] }),
    .E1END({\Tile_X3Y1_E1BEG[3] ,
    \Tile_X3Y1_E1BEG[2] ,
    \Tile_X3Y1_E1BEG[1] ,
    \Tile_X3Y1_E1BEG[0] }),
    .E2BEG({\Tile_X4Y1_E2BEG[7] ,
    \Tile_X4Y1_E2BEG[6] ,
    \Tile_X4Y1_E2BEG[5] ,
    \Tile_X4Y1_E2BEG[4] ,
    \Tile_X4Y1_E2BEG[3] ,
    \Tile_X4Y1_E2BEG[2] ,
    \Tile_X4Y1_E2BEG[1] ,
    \Tile_X4Y1_E2BEG[0] }),
    .E2BEGb({\Tile_X4Y1_E2BEGb[7] ,
    \Tile_X4Y1_E2BEGb[6] ,
    \Tile_X4Y1_E2BEGb[5] ,
    \Tile_X4Y1_E2BEGb[4] ,
    \Tile_X4Y1_E2BEGb[3] ,
    \Tile_X4Y1_E2BEGb[2] ,
    \Tile_X4Y1_E2BEGb[1] ,
    \Tile_X4Y1_E2BEGb[0] }),
    .E2END({\Tile_X3Y1_E2BEGb[7] ,
    \Tile_X3Y1_E2BEGb[6] ,
    \Tile_X3Y1_E2BEGb[5] ,
    \Tile_X3Y1_E2BEGb[4] ,
    \Tile_X3Y1_E2BEGb[3] ,
    \Tile_X3Y1_E2BEGb[2] ,
    \Tile_X3Y1_E2BEGb[1] ,
    \Tile_X3Y1_E2BEGb[0] }),
    .E2MID({\Tile_X3Y1_E2BEG[7] ,
    \Tile_X3Y1_E2BEG[6] ,
    \Tile_X3Y1_E2BEG[5] ,
    \Tile_X3Y1_E2BEG[4] ,
    \Tile_X3Y1_E2BEG[3] ,
    \Tile_X3Y1_E2BEG[2] ,
    \Tile_X3Y1_E2BEG[1] ,
    \Tile_X3Y1_E2BEG[0] }),
    .E6BEG({\Tile_X4Y1_E6BEG[11] ,
    \Tile_X4Y1_E6BEG[10] ,
    \Tile_X4Y1_E6BEG[9] ,
    \Tile_X4Y1_E6BEG[8] ,
    \Tile_X4Y1_E6BEG[7] ,
    \Tile_X4Y1_E6BEG[6] ,
    \Tile_X4Y1_E6BEG[5] ,
    \Tile_X4Y1_E6BEG[4] ,
    \Tile_X4Y1_E6BEG[3] ,
    \Tile_X4Y1_E6BEG[2] ,
    \Tile_X4Y1_E6BEG[1] ,
    \Tile_X4Y1_E6BEG[0] }),
    .E6END({\Tile_X3Y1_E6BEG[11] ,
    \Tile_X3Y1_E6BEG[10] ,
    \Tile_X3Y1_E6BEG[9] ,
    \Tile_X3Y1_E6BEG[8] ,
    \Tile_X3Y1_E6BEG[7] ,
    \Tile_X3Y1_E6BEG[6] ,
    \Tile_X3Y1_E6BEG[5] ,
    \Tile_X3Y1_E6BEG[4] ,
    \Tile_X3Y1_E6BEG[3] ,
    \Tile_X3Y1_E6BEG[2] ,
    \Tile_X3Y1_E6BEG[1] ,
    \Tile_X3Y1_E6BEG[0] }),
    .EE4BEG({\Tile_X4Y1_EE4BEG[15] ,
    \Tile_X4Y1_EE4BEG[14] ,
    \Tile_X4Y1_EE4BEG[13] ,
    \Tile_X4Y1_EE4BEG[12] ,
    \Tile_X4Y1_EE4BEG[11] ,
    \Tile_X4Y1_EE4BEG[10] ,
    \Tile_X4Y1_EE4BEG[9] ,
    \Tile_X4Y1_EE4BEG[8] ,
    \Tile_X4Y1_EE4BEG[7] ,
    \Tile_X4Y1_EE4BEG[6] ,
    \Tile_X4Y1_EE4BEG[5] ,
    \Tile_X4Y1_EE4BEG[4] ,
    \Tile_X4Y1_EE4BEG[3] ,
    \Tile_X4Y1_EE4BEG[2] ,
    \Tile_X4Y1_EE4BEG[1] ,
    \Tile_X4Y1_EE4BEG[0] }),
    .EE4END({\Tile_X3Y1_EE4BEG[15] ,
    \Tile_X3Y1_EE4BEG[14] ,
    \Tile_X3Y1_EE4BEG[13] ,
    \Tile_X3Y1_EE4BEG[12] ,
    \Tile_X3Y1_EE4BEG[11] ,
    \Tile_X3Y1_EE4BEG[10] ,
    \Tile_X3Y1_EE4BEG[9] ,
    \Tile_X3Y1_EE4BEG[8] ,
    \Tile_X3Y1_EE4BEG[7] ,
    \Tile_X3Y1_EE4BEG[6] ,
    \Tile_X3Y1_EE4BEG[5] ,
    \Tile_X3Y1_EE4BEG[4] ,
    \Tile_X3Y1_EE4BEG[3] ,
    \Tile_X3Y1_EE4BEG[2] ,
    \Tile_X3Y1_EE4BEG[1] ,
    \Tile_X3Y1_EE4BEG[0] }),
    .FrameData({\Tile_X3Y1_FrameData_O[31] ,
    \Tile_X3Y1_FrameData_O[30] ,
    \Tile_X3Y1_FrameData_O[29] ,
    \Tile_X3Y1_FrameData_O[28] ,
    \Tile_X3Y1_FrameData_O[27] ,
    \Tile_X3Y1_FrameData_O[26] ,
    \Tile_X3Y1_FrameData_O[25] ,
    \Tile_X3Y1_FrameData_O[24] ,
    \Tile_X3Y1_FrameData_O[23] ,
    \Tile_X3Y1_FrameData_O[22] ,
    \Tile_X3Y1_FrameData_O[21] ,
    \Tile_X3Y1_FrameData_O[20] ,
    \Tile_X3Y1_FrameData_O[19] ,
    \Tile_X3Y1_FrameData_O[18] ,
    \Tile_X3Y1_FrameData_O[17] ,
    \Tile_X3Y1_FrameData_O[16] ,
    \Tile_X3Y1_FrameData_O[15] ,
    \Tile_X3Y1_FrameData_O[14] ,
    \Tile_X3Y1_FrameData_O[13] ,
    \Tile_X3Y1_FrameData_O[12] ,
    \Tile_X3Y1_FrameData_O[11] ,
    \Tile_X3Y1_FrameData_O[10] ,
    \Tile_X3Y1_FrameData_O[9] ,
    \Tile_X3Y1_FrameData_O[8] ,
    \Tile_X3Y1_FrameData_O[7] ,
    \Tile_X3Y1_FrameData_O[6] ,
    \Tile_X3Y1_FrameData_O[5] ,
    \Tile_X3Y1_FrameData_O[4] ,
    \Tile_X3Y1_FrameData_O[3] ,
    \Tile_X3Y1_FrameData_O[2] ,
    \Tile_X3Y1_FrameData_O[1] ,
    \Tile_X3Y1_FrameData_O[0] }),
    .FrameData_O({\Tile_X4Y1_FrameData_O[31] ,
    \Tile_X4Y1_FrameData_O[30] ,
    \Tile_X4Y1_FrameData_O[29] ,
    \Tile_X4Y1_FrameData_O[28] ,
    \Tile_X4Y1_FrameData_O[27] ,
    \Tile_X4Y1_FrameData_O[26] ,
    \Tile_X4Y1_FrameData_O[25] ,
    \Tile_X4Y1_FrameData_O[24] ,
    \Tile_X4Y1_FrameData_O[23] ,
    \Tile_X4Y1_FrameData_O[22] ,
    \Tile_X4Y1_FrameData_O[21] ,
    \Tile_X4Y1_FrameData_O[20] ,
    \Tile_X4Y1_FrameData_O[19] ,
    \Tile_X4Y1_FrameData_O[18] ,
    \Tile_X4Y1_FrameData_O[17] ,
    \Tile_X4Y1_FrameData_O[16] ,
    \Tile_X4Y1_FrameData_O[15] ,
    \Tile_X4Y1_FrameData_O[14] ,
    \Tile_X4Y1_FrameData_O[13] ,
    \Tile_X4Y1_FrameData_O[12] ,
    \Tile_X4Y1_FrameData_O[11] ,
    \Tile_X4Y1_FrameData_O[10] ,
    \Tile_X4Y1_FrameData_O[9] ,
    \Tile_X4Y1_FrameData_O[8] ,
    \Tile_X4Y1_FrameData_O[7] ,
    \Tile_X4Y1_FrameData_O[6] ,
    \Tile_X4Y1_FrameData_O[5] ,
    \Tile_X4Y1_FrameData_O[4] ,
    \Tile_X4Y1_FrameData_O[3] ,
    \Tile_X4Y1_FrameData_O[2] ,
    \Tile_X4Y1_FrameData_O[1] ,
    \Tile_X4Y1_FrameData_O[0] }),
    .FrameStrobe({\Tile_X4Y2_FrameStrobe_O[19] ,
    \Tile_X4Y2_FrameStrobe_O[18] ,
    \Tile_X4Y2_FrameStrobe_O[17] ,
    \Tile_X4Y2_FrameStrobe_O[16] ,
    \Tile_X4Y2_FrameStrobe_O[15] ,
    \Tile_X4Y2_FrameStrobe_O[14] ,
    \Tile_X4Y2_FrameStrobe_O[13] ,
    \Tile_X4Y2_FrameStrobe_O[12] ,
    \Tile_X4Y2_FrameStrobe_O[11] ,
    \Tile_X4Y2_FrameStrobe_O[10] ,
    \Tile_X4Y2_FrameStrobe_O[9] ,
    \Tile_X4Y2_FrameStrobe_O[8] ,
    \Tile_X4Y2_FrameStrobe_O[7] ,
    \Tile_X4Y2_FrameStrobe_O[6] ,
    \Tile_X4Y2_FrameStrobe_O[5] ,
    \Tile_X4Y2_FrameStrobe_O[4] ,
    \Tile_X4Y2_FrameStrobe_O[3] ,
    \Tile_X4Y2_FrameStrobe_O[2] ,
    \Tile_X4Y2_FrameStrobe_O[1] ,
    \Tile_X4Y2_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X4Y1_FrameStrobe_O[19] ,
    \Tile_X4Y1_FrameStrobe_O[18] ,
    \Tile_X4Y1_FrameStrobe_O[17] ,
    \Tile_X4Y1_FrameStrobe_O[16] ,
    \Tile_X4Y1_FrameStrobe_O[15] ,
    \Tile_X4Y1_FrameStrobe_O[14] ,
    \Tile_X4Y1_FrameStrobe_O[13] ,
    \Tile_X4Y1_FrameStrobe_O[12] ,
    \Tile_X4Y1_FrameStrobe_O[11] ,
    \Tile_X4Y1_FrameStrobe_O[10] ,
    \Tile_X4Y1_FrameStrobe_O[9] ,
    \Tile_X4Y1_FrameStrobe_O[8] ,
    \Tile_X4Y1_FrameStrobe_O[7] ,
    \Tile_X4Y1_FrameStrobe_O[6] ,
    \Tile_X4Y1_FrameStrobe_O[5] ,
    \Tile_X4Y1_FrameStrobe_O[4] ,
    \Tile_X4Y1_FrameStrobe_O[3] ,
    \Tile_X4Y1_FrameStrobe_O[2] ,
    \Tile_X4Y1_FrameStrobe_O[1] ,
    \Tile_X4Y1_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X4Y1_N1BEG[3] ,
    \Tile_X4Y1_N1BEG[2] ,
    \Tile_X4Y1_N1BEG[1] ,
    \Tile_X4Y1_N1BEG[0] }),
    .N1END({\Tile_X4Y2_N1BEG[3] ,
    \Tile_X4Y2_N1BEG[2] ,
    \Tile_X4Y2_N1BEG[1] ,
    \Tile_X4Y2_N1BEG[0] }),
    .N2BEG({\Tile_X4Y1_N2BEG[7] ,
    \Tile_X4Y1_N2BEG[6] ,
    \Tile_X4Y1_N2BEG[5] ,
    \Tile_X4Y1_N2BEG[4] ,
    \Tile_X4Y1_N2BEG[3] ,
    \Tile_X4Y1_N2BEG[2] ,
    \Tile_X4Y1_N2BEG[1] ,
    \Tile_X4Y1_N2BEG[0] }),
    .N2BEGb({\Tile_X4Y1_N2BEGb[7] ,
    \Tile_X4Y1_N2BEGb[6] ,
    \Tile_X4Y1_N2BEGb[5] ,
    \Tile_X4Y1_N2BEGb[4] ,
    \Tile_X4Y1_N2BEGb[3] ,
    \Tile_X4Y1_N2BEGb[2] ,
    \Tile_X4Y1_N2BEGb[1] ,
    \Tile_X4Y1_N2BEGb[0] }),
    .N2END({\Tile_X4Y2_N2BEGb[7] ,
    \Tile_X4Y2_N2BEGb[6] ,
    \Tile_X4Y2_N2BEGb[5] ,
    \Tile_X4Y2_N2BEGb[4] ,
    \Tile_X4Y2_N2BEGb[3] ,
    \Tile_X4Y2_N2BEGb[2] ,
    \Tile_X4Y2_N2BEGb[1] ,
    \Tile_X4Y2_N2BEGb[0] }),
    .N2MID({\Tile_X4Y2_N2BEG[7] ,
    \Tile_X4Y2_N2BEG[6] ,
    \Tile_X4Y2_N2BEG[5] ,
    \Tile_X4Y2_N2BEG[4] ,
    \Tile_X4Y2_N2BEG[3] ,
    \Tile_X4Y2_N2BEG[2] ,
    \Tile_X4Y2_N2BEG[1] ,
    \Tile_X4Y2_N2BEG[0] }),
    .N4BEG({\Tile_X4Y1_N4BEG[15] ,
    \Tile_X4Y1_N4BEG[14] ,
    \Tile_X4Y1_N4BEG[13] ,
    \Tile_X4Y1_N4BEG[12] ,
    \Tile_X4Y1_N4BEG[11] ,
    \Tile_X4Y1_N4BEG[10] ,
    \Tile_X4Y1_N4BEG[9] ,
    \Tile_X4Y1_N4BEG[8] ,
    \Tile_X4Y1_N4BEG[7] ,
    \Tile_X4Y1_N4BEG[6] ,
    \Tile_X4Y1_N4BEG[5] ,
    \Tile_X4Y1_N4BEG[4] ,
    \Tile_X4Y1_N4BEG[3] ,
    \Tile_X4Y1_N4BEG[2] ,
    \Tile_X4Y1_N4BEG[1] ,
    \Tile_X4Y1_N4BEG[0] }),
    .N4END({\Tile_X4Y2_N4BEG[15] ,
    \Tile_X4Y2_N4BEG[14] ,
    \Tile_X4Y2_N4BEG[13] ,
    \Tile_X4Y2_N4BEG[12] ,
    \Tile_X4Y2_N4BEG[11] ,
    \Tile_X4Y2_N4BEG[10] ,
    \Tile_X4Y2_N4BEG[9] ,
    \Tile_X4Y2_N4BEG[8] ,
    \Tile_X4Y2_N4BEG[7] ,
    \Tile_X4Y2_N4BEG[6] ,
    \Tile_X4Y2_N4BEG[5] ,
    \Tile_X4Y2_N4BEG[4] ,
    \Tile_X4Y2_N4BEG[3] ,
    \Tile_X4Y2_N4BEG[2] ,
    \Tile_X4Y2_N4BEG[1] ,
    \Tile_X4Y2_N4BEG[0] }),
    .NN4BEG({\Tile_X4Y1_NN4BEG[15] ,
    \Tile_X4Y1_NN4BEG[14] ,
    \Tile_X4Y1_NN4BEG[13] ,
    \Tile_X4Y1_NN4BEG[12] ,
    \Tile_X4Y1_NN4BEG[11] ,
    \Tile_X4Y1_NN4BEG[10] ,
    \Tile_X4Y1_NN4BEG[9] ,
    \Tile_X4Y1_NN4BEG[8] ,
    \Tile_X4Y1_NN4BEG[7] ,
    \Tile_X4Y1_NN4BEG[6] ,
    \Tile_X4Y1_NN4BEG[5] ,
    \Tile_X4Y1_NN4BEG[4] ,
    \Tile_X4Y1_NN4BEG[3] ,
    \Tile_X4Y1_NN4BEG[2] ,
    \Tile_X4Y1_NN4BEG[1] ,
    \Tile_X4Y1_NN4BEG[0] }),
    .NN4END({\Tile_X4Y2_NN4BEG[15] ,
    \Tile_X4Y2_NN4BEG[14] ,
    \Tile_X4Y2_NN4BEG[13] ,
    \Tile_X4Y2_NN4BEG[12] ,
    \Tile_X4Y2_NN4BEG[11] ,
    \Tile_X4Y2_NN4BEG[10] ,
    \Tile_X4Y2_NN4BEG[9] ,
    \Tile_X4Y2_NN4BEG[8] ,
    \Tile_X4Y2_NN4BEG[7] ,
    \Tile_X4Y2_NN4BEG[6] ,
    \Tile_X4Y2_NN4BEG[5] ,
    \Tile_X4Y2_NN4BEG[4] ,
    \Tile_X4Y2_NN4BEG[3] ,
    \Tile_X4Y2_NN4BEG[2] ,
    \Tile_X4Y2_NN4BEG[1] ,
    \Tile_X4Y2_NN4BEG[0] }),
    .S1BEG({\Tile_X4Y1_S1BEG[3] ,
    \Tile_X4Y1_S1BEG[2] ,
    \Tile_X4Y1_S1BEG[1] ,
    \Tile_X4Y1_S1BEG[0] }),
    .S1END({\Tile_X4Y0_S1BEG[3] ,
    \Tile_X4Y0_S1BEG[2] ,
    \Tile_X4Y0_S1BEG[1] ,
    \Tile_X4Y0_S1BEG[0] }),
    .S2BEG({\Tile_X4Y1_S2BEG[7] ,
    \Tile_X4Y1_S2BEG[6] ,
    \Tile_X4Y1_S2BEG[5] ,
    \Tile_X4Y1_S2BEG[4] ,
    \Tile_X4Y1_S2BEG[3] ,
    \Tile_X4Y1_S2BEG[2] ,
    \Tile_X4Y1_S2BEG[1] ,
    \Tile_X4Y1_S2BEG[0] }),
    .S2BEGb({\Tile_X4Y1_S2BEGb[7] ,
    \Tile_X4Y1_S2BEGb[6] ,
    \Tile_X4Y1_S2BEGb[5] ,
    \Tile_X4Y1_S2BEGb[4] ,
    \Tile_X4Y1_S2BEGb[3] ,
    \Tile_X4Y1_S2BEGb[2] ,
    \Tile_X4Y1_S2BEGb[1] ,
    \Tile_X4Y1_S2BEGb[0] }),
    .S2END({\Tile_X4Y0_S2BEGb[7] ,
    \Tile_X4Y0_S2BEGb[6] ,
    \Tile_X4Y0_S2BEGb[5] ,
    \Tile_X4Y0_S2BEGb[4] ,
    \Tile_X4Y0_S2BEGb[3] ,
    \Tile_X4Y0_S2BEGb[2] ,
    \Tile_X4Y0_S2BEGb[1] ,
    \Tile_X4Y0_S2BEGb[0] }),
    .S2MID({\Tile_X4Y0_S2BEG[7] ,
    \Tile_X4Y0_S2BEG[6] ,
    \Tile_X4Y0_S2BEG[5] ,
    \Tile_X4Y0_S2BEG[4] ,
    \Tile_X4Y0_S2BEG[3] ,
    \Tile_X4Y0_S2BEG[2] ,
    \Tile_X4Y0_S2BEG[1] ,
    \Tile_X4Y0_S2BEG[0] }),
    .S4BEG({\Tile_X4Y1_S4BEG[15] ,
    \Tile_X4Y1_S4BEG[14] ,
    \Tile_X4Y1_S4BEG[13] ,
    \Tile_X4Y1_S4BEG[12] ,
    \Tile_X4Y1_S4BEG[11] ,
    \Tile_X4Y1_S4BEG[10] ,
    \Tile_X4Y1_S4BEG[9] ,
    \Tile_X4Y1_S4BEG[8] ,
    \Tile_X4Y1_S4BEG[7] ,
    \Tile_X4Y1_S4BEG[6] ,
    \Tile_X4Y1_S4BEG[5] ,
    \Tile_X4Y1_S4BEG[4] ,
    \Tile_X4Y1_S4BEG[3] ,
    \Tile_X4Y1_S4BEG[2] ,
    \Tile_X4Y1_S4BEG[1] ,
    \Tile_X4Y1_S4BEG[0] }),
    .S4END({\Tile_X4Y0_S4BEG[15] ,
    \Tile_X4Y0_S4BEG[14] ,
    \Tile_X4Y0_S4BEG[13] ,
    \Tile_X4Y0_S4BEG[12] ,
    \Tile_X4Y0_S4BEG[11] ,
    \Tile_X4Y0_S4BEG[10] ,
    \Tile_X4Y0_S4BEG[9] ,
    \Tile_X4Y0_S4BEG[8] ,
    \Tile_X4Y0_S4BEG[7] ,
    \Tile_X4Y0_S4BEG[6] ,
    \Tile_X4Y0_S4BEG[5] ,
    \Tile_X4Y0_S4BEG[4] ,
    \Tile_X4Y0_S4BEG[3] ,
    \Tile_X4Y0_S4BEG[2] ,
    \Tile_X4Y0_S4BEG[1] ,
    \Tile_X4Y0_S4BEG[0] }),
    .SS4BEG({\Tile_X4Y1_SS4BEG[15] ,
    \Tile_X4Y1_SS4BEG[14] ,
    \Tile_X4Y1_SS4BEG[13] ,
    \Tile_X4Y1_SS4BEG[12] ,
    \Tile_X4Y1_SS4BEG[11] ,
    \Tile_X4Y1_SS4BEG[10] ,
    \Tile_X4Y1_SS4BEG[9] ,
    \Tile_X4Y1_SS4BEG[8] ,
    \Tile_X4Y1_SS4BEG[7] ,
    \Tile_X4Y1_SS4BEG[6] ,
    \Tile_X4Y1_SS4BEG[5] ,
    \Tile_X4Y1_SS4BEG[4] ,
    \Tile_X4Y1_SS4BEG[3] ,
    \Tile_X4Y1_SS4BEG[2] ,
    \Tile_X4Y1_SS4BEG[1] ,
    \Tile_X4Y1_SS4BEG[0] }),
    .SS4END({\Tile_X4Y0_SS4BEG[15] ,
    \Tile_X4Y0_SS4BEG[14] ,
    \Tile_X4Y0_SS4BEG[13] ,
    \Tile_X4Y0_SS4BEG[12] ,
    \Tile_X4Y0_SS4BEG[11] ,
    \Tile_X4Y0_SS4BEG[10] ,
    \Tile_X4Y0_SS4BEG[9] ,
    \Tile_X4Y0_SS4BEG[8] ,
    \Tile_X4Y0_SS4BEG[7] ,
    \Tile_X4Y0_SS4BEG[6] ,
    \Tile_X4Y0_SS4BEG[5] ,
    \Tile_X4Y0_SS4BEG[4] ,
    \Tile_X4Y0_SS4BEG[3] ,
    \Tile_X4Y0_SS4BEG[2] ,
    \Tile_X4Y0_SS4BEG[1] ,
    \Tile_X4Y0_SS4BEG[0] }),
    .W1BEG({\Tile_X4Y1_W1BEG[3] ,
    \Tile_X4Y1_W1BEG[2] ,
    \Tile_X4Y1_W1BEG[1] ,
    \Tile_X4Y1_W1BEG[0] }),
    .W1END({\Tile_X5Y1_W1BEG[3] ,
    \Tile_X5Y1_W1BEG[2] ,
    \Tile_X5Y1_W1BEG[1] ,
    \Tile_X5Y1_W1BEG[0] }),
    .W2BEG({\Tile_X4Y1_W2BEG[7] ,
    \Tile_X4Y1_W2BEG[6] ,
    \Tile_X4Y1_W2BEG[5] ,
    \Tile_X4Y1_W2BEG[4] ,
    \Tile_X4Y1_W2BEG[3] ,
    \Tile_X4Y1_W2BEG[2] ,
    \Tile_X4Y1_W2BEG[1] ,
    \Tile_X4Y1_W2BEG[0] }),
    .W2BEGb({\Tile_X4Y1_W2BEGb[7] ,
    \Tile_X4Y1_W2BEGb[6] ,
    \Tile_X4Y1_W2BEGb[5] ,
    \Tile_X4Y1_W2BEGb[4] ,
    \Tile_X4Y1_W2BEGb[3] ,
    \Tile_X4Y1_W2BEGb[2] ,
    \Tile_X4Y1_W2BEGb[1] ,
    \Tile_X4Y1_W2BEGb[0] }),
    .W2END({\Tile_X5Y1_W2BEGb[7] ,
    \Tile_X5Y1_W2BEGb[6] ,
    \Tile_X5Y1_W2BEGb[5] ,
    \Tile_X5Y1_W2BEGb[4] ,
    \Tile_X5Y1_W2BEGb[3] ,
    \Tile_X5Y1_W2BEGb[2] ,
    \Tile_X5Y1_W2BEGb[1] ,
    \Tile_X5Y1_W2BEGb[0] }),
    .W2MID({\Tile_X5Y1_W2BEG[7] ,
    \Tile_X5Y1_W2BEG[6] ,
    \Tile_X5Y1_W2BEG[5] ,
    \Tile_X5Y1_W2BEG[4] ,
    \Tile_X5Y1_W2BEG[3] ,
    \Tile_X5Y1_W2BEG[2] ,
    \Tile_X5Y1_W2BEG[1] ,
    \Tile_X5Y1_W2BEG[0] }),
    .W6BEG({\Tile_X4Y1_W6BEG[11] ,
    \Tile_X4Y1_W6BEG[10] ,
    \Tile_X4Y1_W6BEG[9] ,
    \Tile_X4Y1_W6BEG[8] ,
    \Tile_X4Y1_W6BEG[7] ,
    \Tile_X4Y1_W6BEG[6] ,
    \Tile_X4Y1_W6BEG[5] ,
    \Tile_X4Y1_W6BEG[4] ,
    \Tile_X4Y1_W6BEG[3] ,
    \Tile_X4Y1_W6BEG[2] ,
    \Tile_X4Y1_W6BEG[1] ,
    \Tile_X4Y1_W6BEG[0] }),
    .W6END({\Tile_X5Y1_W6BEG[11] ,
    \Tile_X5Y1_W6BEG[10] ,
    \Tile_X5Y1_W6BEG[9] ,
    \Tile_X5Y1_W6BEG[8] ,
    \Tile_X5Y1_W6BEG[7] ,
    \Tile_X5Y1_W6BEG[6] ,
    \Tile_X5Y1_W6BEG[5] ,
    \Tile_X5Y1_W6BEG[4] ,
    \Tile_X5Y1_W6BEG[3] ,
    \Tile_X5Y1_W6BEG[2] ,
    \Tile_X5Y1_W6BEG[1] ,
    \Tile_X5Y1_W6BEG[0] }),
    .WW4BEG({\Tile_X4Y1_WW4BEG[15] ,
    \Tile_X4Y1_WW4BEG[14] ,
    \Tile_X4Y1_WW4BEG[13] ,
    \Tile_X4Y1_WW4BEG[12] ,
    \Tile_X4Y1_WW4BEG[11] ,
    \Tile_X4Y1_WW4BEG[10] ,
    \Tile_X4Y1_WW4BEG[9] ,
    \Tile_X4Y1_WW4BEG[8] ,
    \Tile_X4Y1_WW4BEG[7] ,
    \Tile_X4Y1_WW4BEG[6] ,
    \Tile_X4Y1_WW4BEG[5] ,
    \Tile_X4Y1_WW4BEG[4] ,
    \Tile_X4Y1_WW4BEG[3] ,
    \Tile_X4Y1_WW4BEG[2] ,
    \Tile_X4Y1_WW4BEG[1] ,
    \Tile_X4Y1_WW4BEG[0] }),
    .WW4END({\Tile_X5Y1_WW4BEG[15] ,
    \Tile_X5Y1_WW4BEG[14] ,
    \Tile_X5Y1_WW4BEG[13] ,
    \Tile_X5Y1_WW4BEG[12] ,
    \Tile_X5Y1_WW4BEG[11] ,
    \Tile_X5Y1_WW4BEG[10] ,
    \Tile_X5Y1_WW4BEG[9] ,
    \Tile_X5Y1_WW4BEG[8] ,
    \Tile_X5Y1_WW4BEG[7] ,
    \Tile_X5Y1_WW4BEG[6] ,
    \Tile_X5Y1_WW4BEG[5] ,
    \Tile_X5Y1_WW4BEG[4] ,
    \Tile_X5Y1_WW4BEG[3] ,
    \Tile_X5Y1_WW4BEG[2] ,
    \Tile_X5Y1_WW4BEG[1] ,
    \Tile_X5Y1_WW4BEG[0] }));
 LUT4AB Tile_X4Y2_LUT4AB (.Ci(Tile_X4Y3_Co),
    .Co(Tile_X4Y2_Co),
    .UserCLK(Tile_X4Y3_UserCLKo),
    .UserCLKo(Tile_X4Y2_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X4Y2_E1BEG[3] ,
    \Tile_X4Y2_E1BEG[2] ,
    \Tile_X4Y2_E1BEG[1] ,
    \Tile_X4Y2_E1BEG[0] }),
    .E1END({\Tile_X3Y2_E1BEG[3] ,
    \Tile_X3Y2_E1BEG[2] ,
    \Tile_X3Y2_E1BEG[1] ,
    \Tile_X3Y2_E1BEG[0] }),
    .E2BEG({\Tile_X4Y2_E2BEG[7] ,
    \Tile_X4Y2_E2BEG[6] ,
    \Tile_X4Y2_E2BEG[5] ,
    \Tile_X4Y2_E2BEG[4] ,
    \Tile_X4Y2_E2BEG[3] ,
    \Tile_X4Y2_E2BEG[2] ,
    \Tile_X4Y2_E2BEG[1] ,
    \Tile_X4Y2_E2BEG[0] }),
    .E2BEGb({\Tile_X4Y2_E2BEGb[7] ,
    \Tile_X4Y2_E2BEGb[6] ,
    \Tile_X4Y2_E2BEGb[5] ,
    \Tile_X4Y2_E2BEGb[4] ,
    \Tile_X4Y2_E2BEGb[3] ,
    \Tile_X4Y2_E2BEGb[2] ,
    \Tile_X4Y2_E2BEGb[1] ,
    \Tile_X4Y2_E2BEGb[0] }),
    .E2END({\Tile_X3Y2_E2BEGb[7] ,
    \Tile_X3Y2_E2BEGb[6] ,
    \Tile_X3Y2_E2BEGb[5] ,
    \Tile_X3Y2_E2BEGb[4] ,
    \Tile_X3Y2_E2BEGb[3] ,
    \Tile_X3Y2_E2BEGb[2] ,
    \Tile_X3Y2_E2BEGb[1] ,
    \Tile_X3Y2_E2BEGb[0] }),
    .E2MID({\Tile_X3Y2_E2BEG[7] ,
    \Tile_X3Y2_E2BEG[6] ,
    \Tile_X3Y2_E2BEG[5] ,
    \Tile_X3Y2_E2BEG[4] ,
    \Tile_X3Y2_E2BEG[3] ,
    \Tile_X3Y2_E2BEG[2] ,
    \Tile_X3Y2_E2BEG[1] ,
    \Tile_X3Y2_E2BEG[0] }),
    .E6BEG({\Tile_X4Y2_E6BEG[11] ,
    \Tile_X4Y2_E6BEG[10] ,
    \Tile_X4Y2_E6BEG[9] ,
    \Tile_X4Y2_E6BEG[8] ,
    \Tile_X4Y2_E6BEG[7] ,
    \Tile_X4Y2_E6BEG[6] ,
    \Tile_X4Y2_E6BEG[5] ,
    \Tile_X4Y2_E6BEG[4] ,
    \Tile_X4Y2_E6BEG[3] ,
    \Tile_X4Y2_E6BEG[2] ,
    \Tile_X4Y2_E6BEG[1] ,
    \Tile_X4Y2_E6BEG[0] }),
    .E6END({\Tile_X3Y2_E6BEG[11] ,
    \Tile_X3Y2_E6BEG[10] ,
    \Tile_X3Y2_E6BEG[9] ,
    \Tile_X3Y2_E6BEG[8] ,
    \Tile_X3Y2_E6BEG[7] ,
    \Tile_X3Y2_E6BEG[6] ,
    \Tile_X3Y2_E6BEG[5] ,
    \Tile_X3Y2_E6BEG[4] ,
    \Tile_X3Y2_E6BEG[3] ,
    \Tile_X3Y2_E6BEG[2] ,
    \Tile_X3Y2_E6BEG[1] ,
    \Tile_X3Y2_E6BEG[0] }),
    .EE4BEG({\Tile_X4Y2_EE4BEG[15] ,
    \Tile_X4Y2_EE4BEG[14] ,
    \Tile_X4Y2_EE4BEG[13] ,
    \Tile_X4Y2_EE4BEG[12] ,
    \Tile_X4Y2_EE4BEG[11] ,
    \Tile_X4Y2_EE4BEG[10] ,
    \Tile_X4Y2_EE4BEG[9] ,
    \Tile_X4Y2_EE4BEG[8] ,
    \Tile_X4Y2_EE4BEG[7] ,
    \Tile_X4Y2_EE4BEG[6] ,
    \Tile_X4Y2_EE4BEG[5] ,
    \Tile_X4Y2_EE4BEG[4] ,
    \Tile_X4Y2_EE4BEG[3] ,
    \Tile_X4Y2_EE4BEG[2] ,
    \Tile_X4Y2_EE4BEG[1] ,
    \Tile_X4Y2_EE4BEG[0] }),
    .EE4END({\Tile_X3Y2_EE4BEG[15] ,
    \Tile_X3Y2_EE4BEG[14] ,
    \Tile_X3Y2_EE4BEG[13] ,
    \Tile_X3Y2_EE4BEG[12] ,
    \Tile_X3Y2_EE4BEG[11] ,
    \Tile_X3Y2_EE4BEG[10] ,
    \Tile_X3Y2_EE4BEG[9] ,
    \Tile_X3Y2_EE4BEG[8] ,
    \Tile_X3Y2_EE4BEG[7] ,
    \Tile_X3Y2_EE4BEG[6] ,
    \Tile_X3Y2_EE4BEG[5] ,
    \Tile_X3Y2_EE4BEG[4] ,
    \Tile_X3Y2_EE4BEG[3] ,
    \Tile_X3Y2_EE4BEG[2] ,
    \Tile_X3Y2_EE4BEG[1] ,
    \Tile_X3Y2_EE4BEG[0] }),
    .FrameData({\Tile_X3Y2_FrameData_O[31] ,
    \Tile_X3Y2_FrameData_O[30] ,
    \Tile_X3Y2_FrameData_O[29] ,
    \Tile_X3Y2_FrameData_O[28] ,
    \Tile_X3Y2_FrameData_O[27] ,
    \Tile_X3Y2_FrameData_O[26] ,
    \Tile_X3Y2_FrameData_O[25] ,
    \Tile_X3Y2_FrameData_O[24] ,
    \Tile_X3Y2_FrameData_O[23] ,
    \Tile_X3Y2_FrameData_O[22] ,
    \Tile_X3Y2_FrameData_O[21] ,
    \Tile_X3Y2_FrameData_O[20] ,
    \Tile_X3Y2_FrameData_O[19] ,
    \Tile_X3Y2_FrameData_O[18] ,
    \Tile_X3Y2_FrameData_O[17] ,
    \Tile_X3Y2_FrameData_O[16] ,
    \Tile_X3Y2_FrameData_O[15] ,
    \Tile_X3Y2_FrameData_O[14] ,
    \Tile_X3Y2_FrameData_O[13] ,
    \Tile_X3Y2_FrameData_O[12] ,
    \Tile_X3Y2_FrameData_O[11] ,
    \Tile_X3Y2_FrameData_O[10] ,
    \Tile_X3Y2_FrameData_O[9] ,
    \Tile_X3Y2_FrameData_O[8] ,
    \Tile_X3Y2_FrameData_O[7] ,
    \Tile_X3Y2_FrameData_O[6] ,
    \Tile_X3Y2_FrameData_O[5] ,
    \Tile_X3Y2_FrameData_O[4] ,
    \Tile_X3Y2_FrameData_O[3] ,
    \Tile_X3Y2_FrameData_O[2] ,
    \Tile_X3Y2_FrameData_O[1] ,
    \Tile_X3Y2_FrameData_O[0] }),
    .FrameData_O({\Tile_X4Y2_FrameData_O[31] ,
    \Tile_X4Y2_FrameData_O[30] ,
    \Tile_X4Y2_FrameData_O[29] ,
    \Tile_X4Y2_FrameData_O[28] ,
    \Tile_X4Y2_FrameData_O[27] ,
    \Tile_X4Y2_FrameData_O[26] ,
    \Tile_X4Y2_FrameData_O[25] ,
    \Tile_X4Y2_FrameData_O[24] ,
    \Tile_X4Y2_FrameData_O[23] ,
    \Tile_X4Y2_FrameData_O[22] ,
    \Tile_X4Y2_FrameData_O[21] ,
    \Tile_X4Y2_FrameData_O[20] ,
    \Tile_X4Y2_FrameData_O[19] ,
    \Tile_X4Y2_FrameData_O[18] ,
    \Tile_X4Y2_FrameData_O[17] ,
    \Tile_X4Y2_FrameData_O[16] ,
    \Tile_X4Y2_FrameData_O[15] ,
    \Tile_X4Y2_FrameData_O[14] ,
    \Tile_X4Y2_FrameData_O[13] ,
    \Tile_X4Y2_FrameData_O[12] ,
    \Tile_X4Y2_FrameData_O[11] ,
    \Tile_X4Y2_FrameData_O[10] ,
    \Tile_X4Y2_FrameData_O[9] ,
    \Tile_X4Y2_FrameData_O[8] ,
    \Tile_X4Y2_FrameData_O[7] ,
    \Tile_X4Y2_FrameData_O[6] ,
    \Tile_X4Y2_FrameData_O[5] ,
    \Tile_X4Y2_FrameData_O[4] ,
    \Tile_X4Y2_FrameData_O[3] ,
    \Tile_X4Y2_FrameData_O[2] ,
    \Tile_X4Y2_FrameData_O[1] ,
    \Tile_X4Y2_FrameData_O[0] }),
    .FrameStrobe({\Tile_X4Y3_FrameStrobe_O[19] ,
    \Tile_X4Y3_FrameStrobe_O[18] ,
    \Tile_X4Y3_FrameStrobe_O[17] ,
    \Tile_X4Y3_FrameStrobe_O[16] ,
    \Tile_X4Y3_FrameStrobe_O[15] ,
    \Tile_X4Y3_FrameStrobe_O[14] ,
    \Tile_X4Y3_FrameStrobe_O[13] ,
    \Tile_X4Y3_FrameStrobe_O[12] ,
    \Tile_X4Y3_FrameStrobe_O[11] ,
    \Tile_X4Y3_FrameStrobe_O[10] ,
    \Tile_X4Y3_FrameStrobe_O[9] ,
    \Tile_X4Y3_FrameStrobe_O[8] ,
    \Tile_X4Y3_FrameStrobe_O[7] ,
    \Tile_X4Y3_FrameStrobe_O[6] ,
    \Tile_X4Y3_FrameStrobe_O[5] ,
    \Tile_X4Y3_FrameStrobe_O[4] ,
    \Tile_X4Y3_FrameStrobe_O[3] ,
    \Tile_X4Y3_FrameStrobe_O[2] ,
    \Tile_X4Y3_FrameStrobe_O[1] ,
    \Tile_X4Y3_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X4Y2_FrameStrobe_O[19] ,
    \Tile_X4Y2_FrameStrobe_O[18] ,
    \Tile_X4Y2_FrameStrobe_O[17] ,
    \Tile_X4Y2_FrameStrobe_O[16] ,
    \Tile_X4Y2_FrameStrobe_O[15] ,
    \Tile_X4Y2_FrameStrobe_O[14] ,
    \Tile_X4Y2_FrameStrobe_O[13] ,
    \Tile_X4Y2_FrameStrobe_O[12] ,
    \Tile_X4Y2_FrameStrobe_O[11] ,
    \Tile_X4Y2_FrameStrobe_O[10] ,
    \Tile_X4Y2_FrameStrobe_O[9] ,
    \Tile_X4Y2_FrameStrobe_O[8] ,
    \Tile_X4Y2_FrameStrobe_O[7] ,
    \Tile_X4Y2_FrameStrobe_O[6] ,
    \Tile_X4Y2_FrameStrobe_O[5] ,
    \Tile_X4Y2_FrameStrobe_O[4] ,
    \Tile_X4Y2_FrameStrobe_O[3] ,
    \Tile_X4Y2_FrameStrobe_O[2] ,
    \Tile_X4Y2_FrameStrobe_O[1] ,
    \Tile_X4Y2_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X4Y2_N1BEG[3] ,
    \Tile_X4Y2_N1BEG[2] ,
    \Tile_X4Y2_N1BEG[1] ,
    \Tile_X4Y2_N1BEG[0] }),
    .N1END({\Tile_X4Y3_N1BEG[3] ,
    \Tile_X4Y3_N1BEG[2] ,
    \Tile_X4Y3_N1BEG[1] ,
    \Tile_X4Y3_N1BEG[0] }),
    .N2BEG({\Tile_X4Y2_N2BEG[7] ,
    \Tile_X4Y2_N2BEG[6] ,
    \Tile_X4Y2_N2BEG[5] ,
    \Tile_X4Y2_N2BEG[4] ,
    \Tile_X4Y2_N2BEG[3] ,
    \Tile_X4Y2_N2BEG[2] ,
    \Tile_X4Y2_N2BEG[1] ,
    \Tile_X4Y2_N2BEG[0] }),
    .N2BEGb({\Tile_X4Y2_N2BEGb[7] ,
    \Tile_X4Y2_N2BEGb[6] ,
    \Tile_X4Y2_N2BEGb[5] ,
    \Tile_X4Y2_N2BEGb[4] ,
    \Tile_X4Y2_N2BEGb[3] ,
    \Tile_X4Y2_N2BEGb[2] ,
    \Tile_X4Y2_N2BEGb[1] ,
    \Tile_X4Y2_N2BEGb[0] }),
    .N2END({\Tile_X4Y3_N2BEGb[7] ,
    \Tile_X4Y3_N2BEGb[6] ,
    \Tile_X4Y3_N2BEGb[5] ,
    \Tile_X4Y3_N2BEGb[4] ,
    \Tile_X4Y3_N2BEGb[3] ,
    \Tile_X4Y3_N2BEGb[2] ,
    \Tile_X4Y3_N2BEGb[1] ,
    \Tile_X4Y3_N2BEGb[0] }),
    .N2MID({\Tile_X4Y3_N2BEG[7] ,
    \Tile_X4Y3_N2BEG[6] ,
    \Tile_X4Y3_N2BEG[5] ,
    \Tile_X4Y3_N2BEG[4] ,
    \Tile_X4Y3_N2BEG[3] ,
    \Tile_X4Y3_N2BEG[2] ,
    \Tile_X4Y3_N2BEG[1] ,
    \Tile_X4Y3_N2BEG[0] }),
    .N4BEG({\Tile_X4Y2_N4BEG[15] ,
    \Tile_X4Y2_N4BEG[14] ,
    \Tile_X4Y2_N4BEG[13] ,
    \Tile_X4Y2_N4BEG[12] ,
    \Tile_X4Y2_N4BEG[11] ,
    \Tile_X4Y2_N4BEG[10] ,
    \Tile_X4Y2_N4BEG[9] ,
    \Tile_X4Y2_N4BEG[8] ,
    \Tile_X4Y2_N4BEG[7] ,
    \Tile_X4Y2_N4BEG[6] ,
    \Tile_X4Y2_N4BEG[5] ,
    \Tile_X4Y2_N4BEG[4] ,
    \Tile_X4Y2_N4BEG[3] ,
    \Tile_X4Y2_N4BEG[2] ,
    \Tile_X4Y2_N4BEG[1] ,
    \Tile_X4Y2_N4BEG[0] }),
    .N4END({\Tile_X4Y3_N4BEG[15] ,
    \Tile_X4Y3_N4BEG[14] ,
    \Tile_X4Y3_N4BEG[13] ,
    \Tile_X4Y3_N4BEG[12] ,
    \Tile_X4Y3_N4BEG[11] ,
    \Tile_X4Y3_N4BEG[10] ,
    \Tile_X4Y3_N4BEG[9] ,
    \Tile_X4Y3_N4BEG[8] ,
    \Tile_X4Y3_N4BEG[7] ,
    \Tile_X4Y3_N4BEG[6] ,
    \Tile_X4Y3_N4BEG[5] ,
    \Tile_X4Y3_N4BEG[4] ,
    \Tile_X4Y3_N4BEG[3] ,
    \Tile_X4Y3_N4BEG[2] ,
    \Tile_X4Y3_N4BEG[1] ,
    \Tile_X4Y3_N4BEG[0] }),
    .NN4BEG({\Tile_X4Y2_NN4BEG[15] ,
    \Tile_X4Y2_NN4BEG[14] ,
    \Tile_X4Y2_NN4BEG[13] ,
    \Tile_X4Y2_NN4BEG[12] ,
    \Tile_X4Y2_NN4BEG[11] ,
    \Tile_X4Y2_NN4BEG[10] ,
    \Tile_X4Y2_NN4BEG[9] ,
    \Tile_X4Y2_NN4BEG[8] ,
    \Tile_X4Y2_NN4BEG[7] ,
    \Tile_X4Y2_NN4BEG[6] ,
    \Tile_X4Y2_NN4BEG[5] ,
    \Tile_X4Y2_NN4BEG[4] ,
    \Tile_X4Y2_NN4BEG[3] ,
    \Tile_X4Y2_NN4BEG[2] ,
    \Tile_X4Y2_NN4BEG[1] ,
    \Tile_X4Y2_NN4BEG[0] }),
    .NN4END({\Tile_X4Y3_NN4BEG[15] ,
    \Tile_X4Y3_NN4BEG[14] ,
    \Tile_X4Y3_NN4BEG[13] ,
    \Tile_X4Y3_NN4BEG[12] ,
    \Tile_X4Y3_NN4BEG[11] ,
    \Tile_X4Y3_NN4BEG[10] ,
    \Tile_X4Y3_NN4BEG[9] ,
    \Tile_X4Y3_NN4BEG[8] ,
    \Tile_X4Y3_NN4BEG[7] ,
    \Tile_X4Y3_NN4BEG[6] ,
    \Tile_X4Y3_NN4BEG[5] ,
    \Tile_X4Y3_NN4BEG[4] ,
    \Tile_X4Y3_NN4BEG[3] ,
    \Tile_X4Y3_NN4BEG[2] ,
    \Tile_X4Y3_NN4BEG[1] ,
    \Tile_X4Y3_NN4BEG[0] }),
    .S1BEG({\Tile_X4Y2_S1BEG[3] ,
    \Tile_X4Y2_S1BEG[2] ,
    \Tile_X4Y2_S1BEG[1] ,
    \Tile_X4Y2_S1BEG[0] }),
    .S1END({\Tile_X4Y1_S1BEG[3] ,
    \Tile_X4Y1_S1BEG[2] ,
    \Tile_X4Y1_S1BEG[1] ,
    \Tile_X4Y1_S1BEG[0] }),
    .S2BEG({\Tile_X4Y2_S2BEG[7] ,
    \Tile_X4Y2_S2BEG[6] ,
    \Tile_X4Y2_S2BEG[5] ,
    \Tile_X4Y2_S2BEG[4] ,
    \Tile_X4Y2_S2BEG[3] ,
    \Tile_X4Y2_S2BEG[2] ,
    \Tile_X4Y2_S2BEG[1] ,
    \Tile_X4Y2_S2BEG[0] }),
    .S2BEGb({\Tile_X4Y2_S2BEGb[7] ,
    \Tile_X4Y2_S2BEGb[6] ,
    \Tile_X4Y2_S2BEGb[5] ,
    \Tile_X4Y2_S2BEGb[4] ,
    \Tile_X4Y2_S2BEGb[3] ,
    \Tile_X4Y2_S2BEGb[2] ,
    \Tile_X4Y2_S2BEGb[1] ,
    \Tile_X4Y2_S2BEGb[0] }),
    .S2END({\Tile_X4Y1_S2BEGb[7] ,
    \Tile_X4Y1_S2BEGb[6] ,
    \Tile_X4Y1_S2BEGb[5] ,
    \Tile_X4Y1_S2BEGb[4] ,
    \Tile_X4Y1_S2BEGb[3] ,
    \Tile_X4Y1_S2BEGb[2] ,
    \Tile_X4Y1_S2BEGb[1] ,
    \Tile_X4Y1_S2BEGb[0] }),
    .S2MID({\Tile_X4Y1_S2BEG[7] ,
    \Tile_X4Y1_S2BEG[6] ,
    \Tile_X4Y1_S2BEG[5] ,
    \Tile_X4Y1_S2BEG[4] ,
    \Tile_X4Y1_S2BEG[3] ,
    \Tile_X4Y1_S2BEG[2] ,
    \Tile_X4Y1_S2BEG[1] ,
    \Tile_X4Y1_S2BEG[0] }),
    .S4BEG({\Tile_X4Y2_S4BEG[15] ,
    \Tile_X4Y2_S4BEG[14] ,
    \Tile_X4Y2_S4BEG[13] ,
    \Tile_X4Y2_S4BEG[12] ,
    \Tile_X4Y2_S4BEG[11] ,
    \Tile_X4Y2_S4BEG[10] ,
    \Tile_X4Y2_S4BEG[9] ,
    \Tile_X4Y2_S4BEG[8] ,
    \Tile_X4Y2_S4BEG[7] ,
    \Tile_X4Y2_S4BEG[6] ,
    \Tile_X4Y2_S4BEG[5] ,
    \Tile_X4Y2_S4BEG[4] ,
    \Tile_X4Y2_S4BEG[3] ,
    \Tile_X4Y2_S4BEG[2] ,
    \Tile_X4Y2_S4BEG[1] ,
    \Tile_X4Y2_S4BEG[0] }),
    .S4END({\Tile_X4Y1_S4BEG[15] ,
    \Tile_X4Y1_S4BEG[14] ,
    \Tile_X4Y1_S4BEG[13] ,
    \Tile_X4Y1_S4BEG[12] ,
    \Tile_X4Y1_S4BEG[11] ,
    \Tile_X4Y1_S4BEG[10] ,
    \Tile_X4Y1_S4BEG[9] ,
    \Tile_X4Y1_S4BEG[8] ,
    \Tile_X4Y1_S4BEG[7] ,
    \Tile_X4Y1_S4BEG[6] ,
    \Tile_X4Y1_S4BEG[5] ,
    \Tile_X4Y1_S4BEG[4] ,
    \Tile_X4Y1_S4BEG[3] ,
    \Tile_X4Y1_S4BEG[2] ,
    \Tile_X4Y1_S4BEG[1] ,
    \Tile_X4Y1_S4BEG[0] }),
    .SS4BEG({\Tile_X4Y2_SS4BEG[15] ,
    \Tile_X4Y2_SS4BEG[14] ,
    \Tile_X4Y2_SS4BEG[13] ,
    \Tile_X4Y2_SS4BEG[12] ,
    \Tile_X4Y2_SS4BEG[11] ,
    \Tile_X4Y2_SS4BEG[10] ,
    \Tile_X4Y2_SS4BEG[9] ,
    \Tile_X4Y2_SS4BEG[8] ,
    \Tile_X4Y2_SS4BEG[7] ,
    \Tile_X4Y2_SS4BEG[6] ,
    \Tile_X4Y2_SS4BEG[5] ,
    \Tile_X4Y2_SS4BEG[4] ,
    \Tile_X4Y2_SS4BEG[3] ,
    \Tile_X4Y2_SS4BEG[2] ,
    \Tile_X4Y2_SS4BEG[1] ,
    \Tile_X4Y2_SS4BEG[0] }),
    .SS4END({\Tile_X4Y1_SS4BEG[15] ,
    \Tile_X4Y1_SS4BEG[14] ,
    \Tile_X4Y1_SS4BEG[13] ,
    \Tile_X4Y1_SS4BEG[12] ,
    \Tile_X4Y1_SS4BEG[11] ,
    \Tile_X4Y1_SS4BEG[10] ,
    \Tile_X4Y1_SS4BEG[9] ,
    \Tile_X4Y1_SS4BEG[8] ,
    \Tile_X4Y1_SS4BEG[7] ,
    \Tile_X4Y1_SS4BEG[6] ,
    \Tile_X4Y1_SS4BEG[5] ,
    \Tile_X4Y1_SS4BEG[4] ,
    \Tile_X4Y1_SS4BEG[3] ,
    \Tile_X4Y1_SS4BEG[2] ,
    \Tile_X4Y1_SS4BEG[1] ,
    \Tile_X4Y1_SS4BEG[0] }),
    .W1BEG({\Tile_X4Y2_W1BEG[3] ,
    \Tile_X4Y2_W1BEG[2] ,
    \Tile_X4Y2_W1BEG[1] ,
    \Tile_X4Y2_W1BEG[0] }),
    .W1END({\Tile_X5Y2_W1BEG[3] ,
    \Tile_X5Y2_W1BEG[2] ,
    \Tile_X5Y2_W1BEG[1] ,
    \Tile_X5Y2_W1BEG[0] }),
    .W2BEG({\Tile_X4Y2_W2BEG[7] ,
    \Tile_X4Y2_W2BEG[6] ,
    \Tile_X4Y2_W2BEG[5] ,
    \Tile_X4Y2_W2BEG[4] ,
    \Tile_X4Y2_W2BEG[3] ,
    \Tile_X4Y2_W2BEG[2] ,
    \Tile_X4Y2_W2BEG[1] ,
    \Tile_X4Y2_W2BEG[0] }),
    .W2BEGb({\Tile_X4Y2_W2BEGb[7] ,
    \Tile_X4Y2_W2BEGb[6] ,
    \Tile_X4Y2_W2BEGb[5] ,
    \Tile_X4Y2_W2BEGb[4] ,
    \Tile_X4Y2_W2BEGb[3] ,
    \Tile_X4Y2_W2BEGb[2] ,
    \Tile_X4Y2_W2BEGb[1] ,
    \Tile_X4Y2_W2BEGb[0] }),
    .W2END({\Tile_X5Y2_W2BEGb[7] ,
    \Tile_X5Y2_W2BEGb[6] ,
    \Tile_X5Y2_W2BEGb[5] ,
    \Tile_X5Y2_W2BEGb[4] ,
    \Tile_X5Y2_W2BEGb[3] ,
    \Tile_X5Y2_W2BEGb[2] ,
    \Tile_X5Y2_W2BEGb[1] ,
    \Tile_X5Y2_W2BEGb[0] }),
    .W2MID({\Tile_X5Y2_W2BEG[7] ,
    \Tile_X5Y2_W2BEG[6] ,
    \Tile_X5Y2_W2BEG[5] ,
    \Tile_X5Y2_W2BEG[4] ,
    \Tile_X5Y2_W2BEG[3] ,
    \Tile_X5Y2_W2BEG[2] ,
    \Tile_X5Y2_W2BEG[1] ,
    \Tile_X5Y2_W2BEG[0] }),
    .W6BEG({\Tile_X4Y2_W6BEG[11] ,
    \Tile_X4Y2_W6BEG[10] ,
    \Tile_X4Y2_W6BEG[9] ,
    \Tile_X4Y2_W6BEG[8] ,
    \Tile_X4Y2_W6BEG[7] ,
    \Tile_X4Y2_W6BEG[6] ,
    \Tile_X4Y2_W6BEG[5] ,
    \Tile_X4Y2_W6BEG[4] ,
    \Tile_X4Y2_W6BEG[3] ,
    \Tile_X4Y2_W6BEG[2] ,
    \Tile_X4Y2_W6BEG[1] ,
    \Tile_X4Y2_W6BEG[0] }),
    .W6END({\Tile_X5Y2_W6BEG[11] ,
    \Tile_X5Y2_W6BEG[10] ,
    \Tile_X5Y2_W6BEG[9] ,
    \Tile_X5Y2_W6BEG[8] ,
    \Tile_X5Y2_W6BEG[7] ,
    \Tile_X5Y2_W6BEG[6] ,
    \Tile_X5Y2_W6BEG[5] ,
    \Tile_X5Y2_W6BEG[4] ,
    \Tile_X5Y2_W6BEG[3] ,
    \Tile_X5Y2_W6BEG[2] ,
    \Tile_X5Y2_W6BEG[1] ,
    \Tile_X5Y2_W6BEG[0] }),
    .WW4BEG({\Tile_X4Y2_WW4BEG[15] ,
    \Tile_X4Y2_WW4BEG[14] ,
    \Tile_X4Y2_WW4BEG[13] ,
    \Tile_X4Y2_WW4BEG[12] ,
    \Tile_X4Y2_WW4BEG[11] ,
    \Tile_X4Y2_WW4BEG[10] ,
    \Tile_X4Y2_WW4BEG[9] ,
    \Tile_X4Y2_WW4BEG[8] ,
    \Tile_X4Y2_WW4BEG[7] ,
    \Tile_X4Y2_WW4BEG[6] ,
    \Tile_X4Y2_WW4BEG[5] ,
    \Tile_X4Y2_WW4BEG[4] ,
    \Tile_X4Y2_WW4BEG[3] ,
    \Tile_X4Y2_WW4BEG[2] ,
    \Tile_X4Y2_WW4BEG[1] ,
    \Tile_X4Y2_WW4BEG[0] }),
    .WW4END({\Tile_X5Y2_WW4BEG[15] ,
    \Tile_X5Y2_WW4BEG[14] ,
    \Tile_X5Y2_WW4BEG[13] ,
    \Tile_X5Y2_WW4BEG[12] ,
    \Tile_X5Y2_WW4BEG[11] ,
    \Tile_X5Y2_WW4BEG[10] ,
    \Tile_X5Y2_WW4BEG[9] ,
    \Tile_X5Y2_WW4BEG[8] ,
    \Tile_X5Y2_WW4BEG[7] ,
    \Tile_X5Y2_WW4BEG[6] ,
    \Tile_X5Y2_WW4BEG[5] ,
    \Tile_X5Y2_WW4BEG[4] ,
    \Tile_X5Y2_WW4BEG[3] ,
    \Tile_X5Y2_WW4BEG[2] ,
    \Tile_X5Y2_WW4BEG[1] ,
    \Tile_X5Y2_WW4BEG[0] }));
 LUT4AB Tile_X4Y3_LUT4AB (.Ci(Tile_X4Y4_Co),
    .Co(Tile_X4Y3_Co),
    .UserCLK(Tile_X4Y4_UserCLKo),
    .UserCLKo(Tile_X4Y3_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X4Y3_E1BEG[3] ,
    \Tile_X4Y3_E1BEG[2] ,
    \Tile_X4Y3_E1BEG[1] ,
    \Tile_X4Y3_E1BEG[0] }),
    .E1END({\Tile_X3Y3_E1BEG[3] ,
    \Tile_X3Y3_E1BEG[2] ,
    \Tile_X3Y3_E1BEG[1] ,
    \Tile_X3Y3_E1BEG[0] }),
    .E2BEG({\Tile_X4Y3_E2BEG[7] ,
    \Tile_X4Y3_E2BEG[6] ,
    \Tile_X4Y3_E2BEG[5] ,
    \Tile_X4Y3_E2BEG[4] ,
    \Tile_X4Y3_E2BEG[3] ,
    \Tile_X4Y3_E2BEG[2] ,
    \Tile_X4Y3_E2BEG[1] ,
    \Tile_X4Y3_E2BEG[0] }),
    .E2BEGb({\Tile_X4Y3_E2BEGb[7] ,
    \Tile_X4Y3_E2BEGb[6] ,
    \Tile_X4Y3_E2BEGb[5] ,
    \Tile_X4Y3_E2BEGb[4] ,
    \Tile_X4Y3_E2BEGb[3] ,
    \Tile_X4Y3_E2BEGb[2] ,
    \Tile_X4Y3_E2BEGb[1] ,
    \Tile_X4Y3_E2BEGb[0] }),
    .E2END({\Tile_X3Y3_E2BEGb[7] ,
    \Tile_X3Y3_E2BEGb[6] ,
    \Tile_X3Y3_E2BEGb[5] ,
    \Tile_X3Y3_E2BEGb[4] ,
    \Tile_X3Y3_E2BEGb[3] ,
    \Tile_X3Y3_E2BEGb[2] ,
    \Tile_X3Y3_E2BEGb[1] ,
    \Tile_X3Y3_E2BEGb[0] }),
    .E2MID({\Tile_X3Y3_E2BEG[7] ,
    \Tile_X3Y3_E2BEG[6] ,
    \Tile_X3Y3_E2BEG[5] ,
    \Tile_X3Y3_E2BEG[4] ,
    \Tile_X3Y3_E2BEG[3] ,
    \Tile_X3Y3_E2BEG[2] ,
    \Tile_X3Y3_E2BEG[1] ,
    \Tile_X3Y3_E2BEG[0] }),
    .E6BEG({\Tile_X4Y3_E6BEG[11] ,
    \Tile_X4Y3_E6BEG[10] ,
    \Tile_X4Y3_E6BEG[9] ,
    \Tile_X4Y3_E6BEG[8] ,
    \Tile_X4Y3_E6BEG[7] ,
    \Tile_X4Y3_E6BEG[6] ,
    \Tile_X4Y3_E6BEG[5] ,
    \Tile_X4Y3_E6BEG[4] ,
    \Tile_X4Y3_E6BEG[3] ,
    \Tile_X4Y3_E6BEG[2] ,
    \Tile_X4Y3_E6BEG[1] ,
    \Tile_X4Y3_E6BEG[0] }),
    .E6END({\Tile_X3Y3_E6BEG[11] ,
    \Tile_X3Y3_E6BEG[10] ,
    \Tile_X3Y3_E6BEG[9] ,
    \Tile_X3Y3_E6BEG[8] ,
    \Tile_X3Y3_E6BEG[7] ,
    \Tile_X3Y3_E6BEG[6] ,
    \Tile_X3Y3_E6BEG[5] ,
    \Tile_X3Y3_E6BEG[4] ,
    \Tile_X3Y3_E6BEG[3] ,
    \Tile_X3Y3_E6BEG[2] ,
    \Tile_X3Y3_E6BEG[1] ,
    \Tile_X3Y3_E6BEG[0] }),
    .EE4BEG({\Tile_X4Y3_EE4BEG[15] ,
    \Tile_X4Y3_EE4BEG[14] ,
    \Tile_X4Y3_EE4BEG[13] ,
    \Tile_X4Y3_EE4BEG[12] ,
    \Tile_X4Y3_EE4BEG[11] ,
    \Tile_X4Y3_EE4BEG[10] ,
    \Tile_X4Y3_EE4BEG[9] ,
    \Tile_X4Y3_EE4BEG[8] ,
    \Tile_X4Y3_EE4BEG[7] ,
    \Tile_X4Y3_EE4BEG[6] ,
    \Tile_X4Y3_EE4BEG[5] ,
    \Tile_X4Y3_EE4BEG[4] ,
    \Tile_X4Y3_EE4BEG[3] ,
    \Tile_X4Y3_EE4BEG[2] ,
    \Tile_X4Y3_EE4BEG[1] ,
    \Tile_X4Y3_EE4BEG[0] }),
    .EE4END({\Tile_X3Y3_EE4BEG[15] ,
    \Tile_X3Y3_EE4BEG[14] ,
    \Tile_X3Y3_EE4BEG[13] ,
    \Tile_X3Y3_EE4BEG[12] ,
    \Tile_X3Y3_EE4BEG[11] ,
    \Tile_X3Y3_EE4BEG[10] ,
    \Tile_X3Y3_EE4BEG[9] ,
    \Tile_X3Y3_EE4BEG[8] ,
    \Tile_X3Y3_EE4BEG[7] ,
    \Tile_X3Y3_EE4BEG[6] ,
    \Tile_X3Y3_EE4BEG[5] ,
    \Tile_X3Y3_EE4BEG[4] ,
    \Tile_X3Y3_EE4BEG[3] ,
    \Tile_X3Y3_EE4BEG[2] ,
    \Tile_X3Y3_EE4BEG[1] ,
    \Tile_X3Y3_EE4BEG[0] }),
    .FrameData({\Tile_X3Y3_FrameData_O[31] ,
    \Tile_X3Y3_FrameData_O[30] ,
    \Tile_X3Y3_FrameData_O[29] ,
    \Tile_X3Y3_FrameData_O[28] ,
    \Tile_X3Y3_FrameData_O[27] ,
    \Tile_X3Y3_FrameData_O[26] ,
    \Tile_X3Y3_FrameData_O[25] ,
    \Tile_X3Y3_FrameData_O[24] ,
    \Tile_X3Y3_FrameData_O[23] ,
    \Tile_X3Y3_FrameData_O[22] ,
    \Tile_X3Y3_FrameData_O[21] ,
    \Tile_X3Y3_FrameData_O[20] ,
    \Tile_X3Y3_FrameData_O[19] ,
    \Tile_X3Y3_FrameData_O[18] ,
    \Tile_X3Y3_FrameData_O[17] ,
    \Tile_X3Y3_FrameData_O[16] ,
    \Tile_X3Y3_FrameData_O[15] ,
    \Tile_X3Y3_FrameData_O[14] ,
    \Tile_X3Y3_FrameData_O[13] ,
    \Tile_X3Y3_FrameData_O[12] ,
    \Tile_X3Y3_FrameData_O[11] ,
    \Tile_X3Y3_FrameData_O[10] ,
    \Tile_X3Y3_FrameData_O[9] ,
    \Tile_X3Y3_FrameData_O[8] ,
    \Tile_X3Y3_FrameData_O[7] ,
    \Tile_X3Y3_FrameData_O[6] ,
    \Tile_X3Y3_FrameData_O[5] ,
    \Tile_X3Y3_FrameData_O[4] ,
    \Tile_X3Y3_FrameData_O[3] ,
    \Tile_X3Y3_FrameData_O[2] ,
    \Tile_X3Y3_FrameData_O[1] ,
    \Tile_X3Y3_FrameData_O[0] }),
    .FrameData_O({\Tile_X4Y3_FrameData_O[31] ,
    \Tile_X4Y3_FrameData_O[30] ,
    \Tile_X4Y3_FrameData_O[29] ,
    \Tile_X4Y3_FrameData_O[28] ,
    \Tile_X4Y3_FrameData_O[27] ,
    \Tile_X4Y3_FrameData_O[26] ,
    \Tile_X4Y3_FrameData_O[25] ,
    \Tile_X4Y3_FrameData_O[24] ,
    \Tile_X4Y3_FrameData_O[23] ,
    \Tile_X4Y3_FrameData_O[22] ,
    \Tile_X4Y3_FrameData_O[21] ,
    \Tile_X4Y3_FrameData_O[20] ,
    \Tile_X4Y3_FrameData_O[19] ,
    \Tile_X4Y3_FrameData_O[18] ,
    \Tile_X4Y3_FrameData_O[17] ,
    \Tile_X4Y3_FrameData_O[16] ,
    \Tile_X4Y3_FrameData_O[15] ,
    \Tile_X4Y3_FrameData_O[14] ,
    \Tile_X4Y3_FrameData_O[13] ,
    \Tile_X4Y3_FrameData_O[12] ,
    \Tile_X4Y3_FrameData_O[11] ,
    \Tile_X4Y3_FrameData_O[10] ,
    \Tile_X4Y3_FrameData_O[9] ,
    \Tile_X4Y3_FrameData_O[8] ,
    \Tile_X4Y3_FrameData_O[7] ,
    \Tile_X4Y3_FrameData_O[6] ,
    \Tile_X4Y3_FrameData_O[5] ,
    \Tile_X4Y3_FrameData_O[4] ,
    \Tile_X4Y3_FrameData_O[3] ,
    \Tile_X4Y3_FrameData_O[2] ,
    \Tile_X4Y3_FrameData_O[1] ,
    \Tile_X4Y3_FrameData_O[0] }),
    .FrameStrobe({\Tile_X4Y4_FrameStrobe_O[19] ,
    \Tile_X4Y4_FrameStrobe_O[18] ,
    \Tile_X4Y4_FrameStrobe_O[17] ,
    \Tile_X4Y4_FrameStrobe_O[16] ,
    \Tile_X4Y4_FrameStrobe_O[15] ,
    \Tile_X4Y4_FrameStrobe_O[14] ,
    \Tile_X4Y4_FrameStrobe_O[13] ,
    \Tile_X4Y4_FrameStrobe_O[12] ,
    \Tile_X4Y4_FrameStrobe_O[11] ,
    \Tile_X4Y4_FrameStrobe_O[10] ,
    \Tile_X4Y4_FrameStrobe_O[9] ,
    \Tile_X4Y4_FrameStrobe_O[8] ,
    \Tile_X4Y4_FrameStrobe_O[7] ,
    \Tile_X4Y4_FrameStrobe_O[6] ,
    \Tile_X4Y4_FrameStrobe_O[5] ,
    \Tile_X4Y4_FrameStrobe_O[4] ,
    \Tile_X4Y4_FrameStrobe_O[3] ,
    \Tile_X4Y4_FrameStrobe_O[2] ,
    \Tile_X4Y4_FrameStrobe_O[1] ,
    \Tile_X4Y4_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X4Y3_FrameStrobe_O[19] ,
    \Tile_X4Y3_FrameStrobe_O[18] ,
    \Tile_X4Y3_FrameStrobe_O[17] ,
    \Tile_X4Y3_FrameStrobe_O[16] ,
    \Tile_X4Y3_FrameStrobe_O[15] ,
    \Tile_X4Y3_FrameStrobe_O[14] ,
    \Tile_X4Y3_FrameStrobe_O[13] ,
    \Tile_X4Y3_FrameStrobe_O[12] ,
    \Tile_X4Y3_FrameStrobe_O[11] ,
    \Tile_X4Y3_FrameStrobe_O[10] ,
    \Tile_X4Y3_FrameStrobe_O[9] ,
    \Tile_X4Y3_FrameStrobe_O[8] ,
    \Tile_X4Y3_FrameStrobe_O[7] ,
    \Tile_X4Y3_FrameStrobe_O[6] ,
    \Tile_X4Y3_FrameStrobe_O[5] ,
    \Tile_X4Y3_FrameStrobe_O[4] ,
    \Tile_X4Y3_FrameStrobe_O[3] ,
    \Tile_X4Y3_FrameStrobe_O[2] ,
    \Tile_X4Y3_FrameStrobe_O[1] ,
    \Tile_X4Y3_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X4Y3_N1BEG[3] ,
    \Tile_X4Y3_N1BEG[2] ,
    \Tile_X4Y3_N1BEG[1] ,
    \Tile_X4Y3_N1BEG[0] }),
    .N1END({\Tile_X4Y4_N1BEG[3] ,
    \Tile_X4Y4_N1BEG[2] ,
    \Tile_X4Y4_N1BEG[1] ,
    \Tile_X4Y4_N1BEG[0] }),
    .N2BEG({\Tile_X4Y3_N2BEG[7] ,
    \Tile_X4Y3_N2BEG[6] ,
    \Tile_X4Y3_N2BEG[5] ,
    \Tile_X4Y3_N2BEG[4] ,
    \Tile_X4Y3_N2BEG[3] ,
    \Tile_X4Y3_N2BEG[2] ,
    \Tile_X4Y3_N2BEG[1] ,
    \Tile_X4Y3_N2BEG[0] }),
    .N2BEGb({\Tile_X4Y3_N2BEGb[7] ,
    \Tile_X4Y3_N2BEGb[6] ,
    \Tile_X4Y3_N2BEGb[5] ,
    \Tile_X4Y3_N2BEGb[4] ,
    \Tile_X4Y3_N2BEGb[3] ,
    \Tile_X4Y3_N2BEGb[2] ,
    \Tile_X4Y3_N2BEGb[1] ,
    \Tile_X4Y3_N2BEGb[0] }),
    .N2END({\Tile_X4Y4_N2BEGb[7] ,
    \Tile_X4Y4_N2BEGb[6] ,
    \Tile_X4Y4_N2BEGb[5] ,
    \Tile_X4Y4_N2BEGb[4] ,
    \Tile_X4Y4_N2BEGb[3] ,
    \Tile_X4Y4_N2BEGb[2] ,
    \Tile_X4Y4_N2BEGb[1] ,
    \Tile_X4Y4_N2BEGb[0] }),
    .N2MID({\Tile_X4Y4_N2BEG[7] ,
    \Tile_X4Y4_N2BEG[6] ,
    \Tile_X4Y4_N2BEG[5] ,
    \Tile_X4Y4_N2BEG[4] ,
    \Tile_X4Y4_N2BEG[3] ,
    \Tile_X4Y4_N2BEG[2] ,
    \Tile_X4Y4_N2BEG[1] ,
    \Tile_X4Y4_N2BEG[0] }),
    .N4BEG({\Tile_X4Y3_N4BEG[15] ,
    \Tile_X4Y3_N4BEG[14] ,
    \Tile_X4Y3_N4BEG[13] ,
    \Tile_X4Y3_N4BEG[12] ,
    \Tile_X4Y3_N4BEG[11] ,
    \Tile_X4Y3_N4BEG[10] ,
    \Tile_X4Y3_N4BEG[9] ,
    \Tile_X4Y3_N4BEG[8] ,
    \Tile_X4Y3_N4BEG[7] ,
    \Tile_X4Y3_N4BEG[6] ,
    \Tile_X4Y3_N4BEG[5] ,
    \Tile_X4Y3_N4BEG[4] ,
    \Tile_X4Y3_N4BEG[3] ,
    \Tile_X4Y3_N4BEG[2] ,
    \Tile_X4Y3_N4BEG[1] ,
    \Tile_X4Y3_N4BEG[0] }),
    .N4END({\Tile_X4Y4_N4BEG[15] ,
    \Tile_X4Y4_N4BEG[14] ,
    \Tile_X4Y4_N4BEG[13] ,
    \Tile_X4Y4_N4BEG[12] ,
    \Tile_X4Y4_N4BEG[11] ,
    \Tile_X4Y4_N4BEG[10] ,
    \Tile_X4Y4_N4BEG[9] ,
    \Tile_X4Y4_N4BEG[8] ,
    \Tile_X4Y4_N4BEG[7] ,
    \Tile_X4Y4_N4BEG[6] ,
    \Tile_X4Y4_N4BEG[5] ,
    \Tile_X4Y4_N4BEG[4] ,
    \Tile_X4Y4_N4BEG[3] ,
    \Tile_X4Y4_N4BEG[2] ,
    \Tile_X4Y4_N4BEG[1] ,
    \Tile_X4Y4_N4BEG[0] }),
    .NN4BEG({\Tile_X4Y3_NN4BEG[15] ,
    \Tile_X4Y3_NN4BEG[14] ,
    \Tile_X4Y3_NN4BEG[13] ,
    \Tile_X4Y3_NN4BEG[12] ,
    \Tile_X4Y3_NN4BEG[11] ,
    \Tile_X4Y3_NN4BEG[10] ,
    \Tile_X4Y3_NN4BEG[9] ,
    \Tile_X4Y3_NN4BEG[8] ,
    \Tile_X4Y3_NN4BEG[7] ,
    \Tile_X4Y3_NN4BEG[6] ,
    \Tile_X4Y3_NN4BEG[5] ,
    \Tile_X4Y3_NN4BEG[4] ,
    \Tile_X4Y3_NN4BEG[3] ,
    \Tile_X4Y3_NN4BEG[2] ,
    \Tile_X4Y3_NN4BEG[1] ,
    \Tile_X4Y3_NN4BEG[0] }),
    .NN4END({\Tile_X4Y4_NN4BEG[15] ,
    \Tile_X4Y4_NN4BEG[14] ,
    \Tile_X4Y4_NN4BEG[13] ,
    \Tile_X4Y4_NN4BEG[12] ,
    \Tile_X4Y4_NN4BEG[11] ,
    \Tile_X4Y4_NN4BEG[10] ,
    \Tile_X4Y4_NN4BEG[9] ,
    \Tile_X4Y4_NN4BEG[8] ,
    \Tile_X4Y4_NN4BEG[7] ,
    \Tile_X4Y4_NN4BEG[6] ,
    \Tile_X4Y4_NN4BEG[5] ,
    \Tile_X4Y4_NN4BEG[4] ,
    \Tile_X4Y4_NN4BEG[3] ,
    \Tile_X4Y4_NN4BEG[2] ,
    \Tile_X4Y4_NN4BEG[1] ,
    \Tile_X4Y4_NN4BEG[0] }),
    .S1BEG({\Tile_X4Y3_S1BEG[3] ,
    \Tile_X4Y3_S1BEG[2] ,
    \Tile_X4Y3_S1BEG[1] ,
    \Tile_X4Y3_S1BEG[0] }),
    .S1END({\Tile_X4Y2_S1BEG[3] ,
    \Tile_X4Y2_S1BEG[2] ,
    \Tile_X4Y2_S1BEG[1] ,
    \Tile_X4Y2_S1BEG[0] }),
    .S2BEG({\Tile_X4Y3_S2BEG[7] ,
    \Tile_X4Y3_S2BEG[6] ,
    \Tile_X4Y3_S2BEG[5] ,
    \Tile_X4Y3_S2BEG[4] ,
    \Tile_X4Y3_S2BEG[3] ,
    \Tile_X4Y3_S2BEG[2] ,
    \Tile_X4Y3_S2BEG[1] ,
    \Tile_X4Y3_S2BEG[0] }),
    .S2BEGb({\Tile_X4Y3_S2BEGb[7] ,
    \Tile_X4Y3_S2BEGb[6] ,
    \Tile_X4Y3_S2BEGb[5] ,
    \Tile_X4Y3_S2BEGb[4] ,
    \Tile_X4Y3_S2BEGb[3] ,
    \Tile_X4Y3_S2BEGb[2] ,
    \Tile_X4Y3_S2BEGb[1] ,
    \Tile_X4Y3_S2BEGb[0] }),
    .S2END({\Tile_X4Y2_S2BEGb[7] ,
    \Tile_X4Y2_S2BEGb[6] ,
    \Tile_X4Y2_S2BEGb[5] ,
    \Tile_X4Y2_S2BEGb[4] ,
    \Tile_X4Y2_S2BEGb[3] ,
    \Tile_X4Y2_S2BEGb[2] ,
    \Tile_X4Y2_S2BEGb[1] ,
    \Tile_X4Y2_S2BEGb[0] }),
    .S2MID({\Tile_X4Y2_S2BEG[7] ,
    \Tile_X4Y2_S2BEG[6] ,
    \Tile_X4Y2_S2BEG[5] ,
    \Tile_X4Y2_S2BEG[4] ,
    \Tile_X4Y2_S2BEG[3] ,
    \Tile_X4Y2_S2BEG[2] ,
    \Tile_X4Y2_S2BEG[1] ,
    \Tile_X4Y2_S2BEG[0] }),
    .S4BEG({\Tile_X4Y3_S4BEG[15] ,
    \Tile_X4Y3_S4BEG[14] ,
    \Tile_X4Y3_S4BEG[13] ,
    \Tile_X4Y3_S4BEG[12] ,
    \Tile_X4Y3_S4BEG[11] ,
    \Tile_X4Y3_S4BEG[10] ,
    \Tile_X4Y3_S4BEG[9] ,
    \Tile_X4Y3_S4BEG[8] ,
    \Tile_X4Y3_S4BEG[7] ,
    \Tile_X4Y3_S4BEG[6] ,
    \Tile_X4Y3_S4BEG[5] ,
    \Tile_X4Y3_S4BEG[4] ,
    \Tile_X4Y3_S4BEG[3] ,
    \Tile_X4Y3_S4BEG[2] ,
    \Tile_X4Y3_S4BEG[1] ,
    \Tile_X4Y3_S4BEG[0] }),
    .S4END({\Tile_X4Y2_S4BEG[15] ,
    \Tile_X4Y2_S4BEG[14] ,
    \Tile_X4Y2_S4BEG[13] ,
    \Tile_X4Y2_S4BEG[12] ,
    \Tile_X4Y2_S4BEG[11] ,
    \Tile_X4Y2_S4BEG[10] ,
    \Tile_X4Y2_S4BEG[9] ,
    \Tile_X4Y2_S4BEG[8] ,
    \Tile_X4Y2_S4BEG[7] ,
    \Tile_X4Y2_S4BEG[6] ,
    \Tile_X4Y2_S4BEG[5] ,
    \Tile_X4Y2_S4BEG[4] ,
    \Tile_X4Y2_S4BEG[3] ,
    \Tile_X4Y2_S4BEG[2] ,
    \Tile_X4Y2_S4BEG[1] ,
    \Tile_X4Y2_S4BEG[0] }),
    .SS4BEG({\Tile_X4Y3_SS4BEG[15] ,
    \Tile_X4Y3_SS4BEG[14] ,
    \Tile_X4Y3_SS4BEG[13] ,
    \Tile_X4Y3_SS4BEG[12] ,
    \Tile_X4Y3_SS4BEG[11] ,
    \Tile_X4Y3_SS4BEG[10] ,
    \Tile_X4Y3_SS4BEG[9] ,
    \Tile_X4Y3_SS4BEG[8] ,
    \Tile_X4Y3_SS4BEG[7] ,
    \Tile_X4Y3_SS4BEG[6] ,
    \Tile_X4Y3_SS4BEG[5] ,
    \Tile_X4Y3_SS4BEG[4] ,
    \Tile_X4Y3_SS4BEG[3] ,
    \Tile_X4Y3_SS4BEG[2] ,
    \Tile_X4Y3_SS4BEG[1] ,
    \Tile_X4Y3_SS4BEG[0] }),
    .SS4END({\Tile_X4Y2_SS4BEG[15] ,
    \Tile_X4Y2_SS4BEG[14] ,
    \Tile_X4Y2_SS4BEG[13] ,
    \Tile_X4Y2_SS4BEG[12] ,
    \Tile_X4Y2_SS4BEG[11] ,
    \Tile_X4Y2_SS4BEG[10] ,
    \Tile_X4Y2_SS4BEG[9] ,
    \Tile_X4Y2_SS4BEG[8] ,
    \Tile_X4Y2_SS4BEG[7] ,
    \Tile_X4Y2_SS4BEG[6] ,
    \Tile_X4Y2_SS4BEG[5] ,
    \Tile_X4Y2_SS4BEG[4] ,
    \Tile_X4Y2_SS4BEG[3] ,
    \Tile_X4Y2_SS4BEG[2] ,
    \Tile_X4Y2_SS4BEG[1] ,
    \Tile_X4Y2_SS4BEG[0] }),
    .W1BEG({\Tile_X4Y3_W1BEG[3] ,
    \Tile_X4Y3_W1BEG[2] ,
    \Tile_X4Y3_W1BEG[1] ,
    \Tile_X4Y3_W1BEG[0] }),
    .W1END({\Tile_X5Y3_W1BEG[3] ,
    \Tile_X5Y3_W1BEG[2] ,
    \Tile_X5Y3_W1BEG[1] ,
    \Tile_X5Y3_W1BEG[0] }),
    .W2BEG({\Tile_X4Y3_W2BEG[7] ,
    \Tile_X4Y3_W2BEG[6] ,
    \Tile_X4Y3_W2BEG[5] ,
    \Tile_X4Y3_W2BEG[4] ,
    \Tile_X4Y3_W2BEG[3] ,
    \Tile_X4Y3_W2BEG[2] ,
    \Tile_X4Y3_W2BEG[1] ,
    \Tile_X4Y3_W2BEG[0] }),
    .W2BEGb({\Tile_X4Y3_W2BEGb[7] ,
    \Tile_X4Y3_W2BEGb[6] ,
    \Tile_X4Y3_W2BEGb[5] ,
    \Tile_X4Y3_W2BEGb[4] ,
    \Tile_X4Y3_W2BEGb[3] ,
    \Tile_X4Y3_W2BEGb[2] ,
    \Tile_X4Y3_W2BEGb[1] ,
    \Tile_X4Y3_W2BEGb[0] }),
    .W2END({\Tile_X5Y3_W2BEGb[7] ,
    \Tile_X5Y3_W2BEGb[6] ,
    \Tile_X5Y3_W2BEGb[5] ,
    \Tile_X5Y3_W2BEGb[4] ,
    \Tile_X5Y3_W2BEGb[3] ,
    \Tile_X5Y3_W2BEGb[2] ,
    \Tile_X5Y3_W2BEGb[1] ,
    \Tile_X5Y3_W2BEGb[0] }),
    .W2MID({\Tile_X5Y3_W2BEG[7] ,
    \Tile_X5Y3_W2BEG[6] ,
    \Tile_X5Y3_W2BEG[5] ,
    \Tile_X5Y3_W2BEG[4] ,
    \Tile_X5Y3_W2BEG[3] ,
    \Tile_X5Y3_W2BEG[2] ,
    \Tile_X5Y3_W2BEG[1] ,
    \Tile_X5Y3_W2BEG[0] }),
    .W6BEG({\Tile_X4Y3_W6BEG[11] ,
    \Tile_X4Y3_W6BEG[10] ,
    \Tile_X4Y3_W6BEG[9] ,
    \Tile_X4Y3_W6BEG[8] ,
    \Tile_X4Y3_W6BEG[7] ,
    \Tile_X4Y3_W6BEG[6] ,
    \Tile_X4Y3_W6BEG[5] ,
    \Tile_X4Y3_W6BEG[4] ,
    \Tile_X4Y3_W6BEG[3] ,
    \Tile_X4Y3_W6BEG[2] ,
    \Tile_X4Y3_W6BEG[1] ,
    \Tile_X4Y3_W6BEG[0] }),
    .W6END({\Tile_X5Y3_W6BEG[11] ,
    \Tile_X5Y3_W6BEG[10] ,
    \Tile_X5Y3_W6BEG[9] ,
    \Tile_X5Y3_W6BEG[8] ,
    \Tile_X5Y3_W6BEG[7] ,
    \Tile_X5Y3_W6BEG[6] ,
    \Tile_X5Y3_W6BEG[5] ,
    \Tile_X5Y3_W6BEG[4] ,
    \Tile_X5Y3_W6BEG[3] ,
    \Tile_X5Y3_W6BEG[2] ,
    \Tile_X5Y3_W6BEG[1] ,
    \Tile_X5Y3_W6BEG[0] }),
    .WW4BEG({\Tile_X4Y3_WW4BEG[15] ,
    \Tile_X4Y3_WW4BEG[14] ,
    \Tile_X4Y3_WW4BEG[13] ,
    \Tile_X4Y3_WW4BEG[12] ,
    \Tile_X4Y3_WW4BEG[11] ,
    \Tile_X4Y3_WW4BEG[10] ,
    \Tile_X4Y3_WW4BEG[9] ,
    \Tile_X4Y3_WW4BEG[8] ,
    \Tile_X4Y3_WW4BEG[7] ,
    \Tile_X4Y3_WW4BEG[6] ,
    \Tile_X4Y3_WW4BEG[5] ,
    \Tile_X4Y3_WW4BEG[4] ,
    \Tile_X4Y3_WW4BEG[3] ,
    \Tile_X4Y3_WW4BEG[2] ,
    \Tile_X4Y3_WW4BEG[1] ,
    \Tile_X4Y3_WW4BEG[0] }),
    .WW4END({\Tile_X5Y3_WW4BEG[15] ,
    \Tile_X5Y3_WW4BEG[14] ,
    \Tile_X5Y3_WW4BEG[13] ,
    \Tile_X5Y3_WW4BEG[12] ,
    \Tile_X5Y3_WW4BEG[11] ,
    \Tile_X5Y3_WW4BEG[10] ,
    \Tile_X5Y3_WW4BEG[9] ,
    \Tile_X5Y3_WW4BEG[8] ,
    \Tile_X5Y3_WW4BEG[7] ,
    \Tile_X5Y3_WW4BEG[6] ,
    \Tile_X5Y3_WW4BEG[5] ,
    \Tile_X5Y3_WW4BEG[4] ,
    \Tile_X5Y3_WW4BEG[3] ,
    \Tile_X5Y3_WW4BEG[2] ,
    \Tile_X5Y3_WW4BEG[1] ,
    \Tile_X5Y3_WW4BEG[0] }));
 LUT4AB Tile_X4Y4_LUT4AB (.Ci(Tile_X4Y5_Co),
    .Co(Tile_X4Y4_Co),
    .UserCLK(Tile_X4Y5_UserCLKo),
    .UserCLKo(Tile_X4Y4_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X4Y4_E1BEG[3] ,
    \Tile_X4Y4_E1BEG[2] ,
    \Tile_X4Y4_E1BEG[1] ,
    \Tile_X4Y4_E1BEG[0] }),
    .E1END({\Tile_X3Y4_E1BEG[3] ,
    \Tile_X3Y4_E1BEG[2] ,
    \Tile_X3Y4_E1BEG[1] ,
    \Tile_X3Y4_E1BEG[0] }),
    .E2BEG({\Tile_X4Y4_E2BEG[7] ,
    \Tile_X4Y4_E2BEG[6] ,
    \Tile_X4Y4_E2BEG[5] ,
    \Tile_X4Y4_E2BEG[4] ,
    \Tile_X4Y4_E2BEG[3] ,
    \Tile_X4Y4_E2BEG[2] ,
    \Tile_X4Y4_E2BEG[1] ,
    \Tile_X4Y4_E2BEG[0] }),
    .E2BEGb({\Tile_X4Y4_E2BEGb[7] ,
    \Tile_X4Y4_E2BEGb[6] ,
    \Tile_X4Y4_E2BEGb[5] ,
    \Tile_X4Y4_E2BEGb[4] ,
    \Tile_X4Y4_E2BEGb[3] ,
    \Tile_X4Y4_E2BEGb[2] ,
    \Tile_X4Y4_E2BEGb[1] ,
    \Tile_X4Y4_E2BEGb[0] }),
    .E2END({\Tile_X3Y4_E2BEGb[7] ,
    \Tile_X3Y4_E2BEGb[6] ,
    \Tile_X3Y4_E2BEGb[5] ,
    \Tile_X3Y4_E2BEGb[4] ,
    \Tile_X3Y4_E2BEGb[3] ,
    \Tile_X3Y4_E2BEGb[2] ,
    \Tile_X3Y4_E2BEGb[1] ,
    \Tile_X3Y4_E2BEGb[0] }),
    .E2MID({\Tile_X3Y4_E2BEG[7] ,
    \Tile_X3Y4_E2BEG[6] ,
    \Tile_X3Y4_E2BEG[5] ,
    \Tile_X3Y4_E2BEG[4] ,
    \Tile_X3Y4_E2BEG[3] ,
    \Tile_X3Y4_E2BEG[2] ,
    \Tile_X3Y4_E2BEG[1] ,
    \Tile_X3Y4_E2BEG[0] }),
    .E6BEG({\Tile_X4Y4_E6BEG[11] ,
    \Tile_X4Y4_E6BEG[10] ,
    \Tile_X4Y4_E6BEG[9] ,
    \Tile_X4Y4_E6BEG[8] ,
    \Tile_X4Y4_E6BEG[7] ,
    \Tile_X4Y4_E6BEG[6] ,
    \Tile_X4Y4_E6BEG[5] ,
    \Tile_X4Y4_E6BEG[4] ,
    \Tile_X4Y4_E6BEG[3] ,
    \Tile_X4Y4_E6BEG[2] ,
    \Tile_X4Y4_E6BEG[1] ,
    \Tile_X4Y4_E6BEG[0] }),
    .E6END({\Tile_X3Y4_E6BEG[11] ,
    \Tile_X3Y4_E6BEG[10] ,
    \Tile_X3Y4_E6BEG[9] ,
    \Tile_X3Y4_E6BEG[8] ,
    \Tile_X3Y4_E6BEG[7] ,
    \Tile_X3Y4_E6BEG[6] ,
    \Tile_X3Y4_E6BEG[5] ,
    \Tile_X3Y4_E6BEG[4] ,
    \Tile_X3Y4_E6BEG[3] ,
    \Tile_X3Y4_E6BEG[2] ,
    \Tile_X3Y4_E6BEG[1] ,
    \Tile_X3Y4_E6BEG[0] }),
    .EE4BEG({\Tile_X4Y4_EE4BEG[15] ,
    \Tile_X4Y4_EE4BEG[14] ,
    \Tile_X4Y4_EE4BEG[13] ,
    \Tile_X4Y4_EE4BEG[12] ,
    \Tile_X4Y4_EE4BEG[11] ,
    \Tile_X4Y4_EE4BEG[10] ,
    \Tile_X4Y4_EE4BEG[9] ,
    \Tile_X4Y4_EE4BEG[8] ,
    \Tile_X4Y4_EE4BEG[7] ,
    \Tile_X4Y4_EE4BEG[6] ,
    \Tile_X4Y4_EE4BEG[5] ,
    \Tile_X4Y4_EE4BEG[4] ,
    \Tile_X4Y4_EE4BEG[3] ,
    \Tile_X4Y4_EE4BEG[2] ,
    \Tile_X4Y4_EE4BEG[1] ,
    \Tile_X4Y4_EE4BEG[0] }),
    .EE4END({\Tile_X3Y4_EE4BEG[15] ,
    \Tile_X3Y4_EE4BEG[14] ,
    \Tile_X3Y4_EE4BEG[13] ,
    \Tile_X3Y4_EE4BEG[12] ,
    \Tile_X3Y4_EE4BEG[11] ,
    \Tile_X3Y4_EE4BEG[10] ,
    \Tile_X3Y4_EE4BEG[9] ,
    \Tile_X3Y4_EE4BEG[8] ,
    \Tile_X3Y4_EE4BEG[7] ,
    \Tile_X3Y4_EE4BEG[6] ,
    \Tile_X3Y4_EE4BEG[5] ,
    \Tile_X3Y4_EE4BEG[4] ,
    \Tile_X3Y4_EE4BEG[3] ,
    \Tile_X3Y4_EE4BEG[2] ,
    \Tile_X3Y4_EE4BEG[1] ,
    \Tile_X3Y4_EE4BEG[0] }),
    .FrameData({\Tile_X3Y4_FrameData_O[31] ,
    \Tile_X3Y4_FrameData_O[30] ,
    \Tile_X3Y4_FrameData_O[29] ,
    \Tile_X3Y4_FrameData_O[28] ,
    \Tile_X3Y4_FrameData_O[27] ,
    \Tile_X3Y4_FrameData_O[26] ,
    \Tile_X3Y4_FrameData_O[25] ,
    \Tile_X3Y4_FrameData_O[24] ,
    \Tile_X3Y4_FrameData_O[23] ,
    \Tile_X3Y4_FrameData_O[22] ,
    \Tile_X3Y4_FrameData_O[21] ,
    \Tile_X3Y4_FrameData_O[20] ,
    \Tile_X3Y4_FrameData_O[19] ,
    \Tile_X3Y4_FrameData_O[18] ,
    \Tile_X3Y4_FrameData_O[17] ,
    \Tile_X3Y4_FrameData_O[16] ,
    \Tile_X3Y4_FrameData_O[15] ,
    \Tile_X3Y4_FrameData_O[14] ,
    \Tile_X3Y4_FrameData_O[13] ,
    \Tile_X3Y4_FrameData_O[12] ,
    \Tile_X3Y4_FrameData_O[11] ,
    \Tile_X3Y4_FrameData_O[10] ,
    \Tile_X3Y4_FrameData_O[9] ,
    \Tile_X3Y4_FrameData_O[8] ,
    \Tile_X3Y4_FrameData_O[7] ,
    \Tile_X3Y4_FrameData_O[6] ,
    \Tile_X3Y4_FrameData_O[5] ,
    \Tile_X3Y4_FrameData_O[4] ,
    \Tile_X3Y4_FrameData_O[3] ,
    \Tile_X3Y4_FrameData_O[2] ,
    \Tile_X3Y4_FrameData_O[1] ,
    \Tile_X3Y4_FrameData_O[0] }),
    .FrameData_O({\Tile_X4Y4_FrameData_O[31] ,
    \Tile_X4Y4_FrameData_O[30] ,
    \Tile_X4Y4_FrameData_O[29] ,
    \Tile_X4Y4_FrameData_O[28] ,
    \Tile_X4Y4_FrameData_O[27] ,
    \Tile_X4Y4_FrameData_O[26] ,
    \Tile_X4Y4_FrameData_O[25] ,
    \Tile_X4Y4_FrameData_O[24] ,
    \Tile_X4Y4_FrameData_O[23] ,
    \Tile_X4Y4_FrameData_O[22] ,
    \Tile_X4Y4_FrameData_O[21] ,
    \Tile_X4Y4_FrameData_O[20] ,
    \Tile_X4Y4_FrameData_O[19] ,
    \Tile_X4Y4_FrameData_O[18] ,
    \Tile_X4Y4_FrameData_O[17] ,
    \Tile_X4Y4_FrameData_O[16] ,
    \Tile_X4Y4_FrameData_O[15] ,
    \Tile_X4Y4_FrameData_O[14] ,
    \Tile_X4Y4_FrameData_O[13] ,
    \Tile_X4Y4_FrameData_O[12] ,
    \Tile_X4Y4_FrameData_O[11] ,
    \Tile_X4Y4_FrameData_O[10] ,
    \Tile_X4Y4_FrameData_O[9] ,
    \Tile_X4Y4_FrameData_O[8] ,
    \Tile_X4Y4_FrameData_O[7] ,
    \Tile_X4Y4_FrameData_O[6] ,
    \Tile_X4Y4_FrameData_O[5] ,
    \Tile_X4Y4_FrameData_O[4] ,
    \Tile_X4Y4_FrameData_O[3] ,
    \Tile_X4Y4_FrameData_O[2] ,
    \Tile_X4Y4_FrameData_O[1] ,
    \Tile_X4Y4_FrameData_O[0] }),
    .FrameStrobe({\Tile_X4Y5_FrameStrobe_O[19] ,
    \Tile_X4Y5_FrameStrobe_O[18] ,
    \Tile_X4Y5_FrameStrobe_O[17] ,
    \Tile_X4Y5_FrameStrobe_O[16] ,
    \Tile_X4Y5_FrameStrobe_O[15] ,
    \Tile_X4Y5_FrameStrobe_O[14] ,
    \Tile_X4Y5_FrameStrobe_O[13] ,
    \Tile_X4Y5_FrameStrobe_O[12] ,
    \Tile_X4Y5_FrameStrobe_O[11] ,
    \Tile_X4Y5_FrameStrobe_O[10] ,
    \Tile_X4Y5_FrameStrobe_O[9] ,
    \Tile_X4Y5_FrameStrobe_O[8] ,
    \Tile_X4Y5_FrameStrobe_O[7] ,
    \Tile_X4Y5_FrameStrobe_O[6] ,
    \Tile_X4Y5_FrameStrobe_O[5] ,
    \Tile_X4Y5_FrameStrobe_O[4] ,
    \Tile_X4Y5_FrameStrobe_O[3] ,
    \Tile_X4Y5_FrameStrobe_O[2] ,
    \Tile_X4Y5_FrameStrobe_O[1] ,
    \Tile_X4Y5_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X4Y4_FrameStrobe_O[19] ,
    \Tile_X4Y4_FrameStrobe_O[18] ,
    \Tile_X4Y4_FrameStrobe_O[17] ,
    \Tile_X4Y4_FrameStrobe_O[16] ,
    \Tile_X4Y4_FrameStrobe_O[15] ,
    \Tile_X4Y4_FrameStrobe_O[14] ,
    \Tile_X4Y4_FrameStrobe_O[13] ,
    \Tile_X4Y4_FrameStrobe_O[12] ,
    \Tile_X4Y4_FrameStrobe_O[11] ,
    \Tile_X4Y4_FrameStrobe_O[10] ,
    \Tile_X4Y4_FrameStrobe_O[9] ,
    \Tile_X4Y4_FrameStrobe_O[8] ,
    \Tile_X4Y4_FrameStrobe_O[7] ,
    \Tile_X4Y4_FrameStrobe_O[6] ,
    \Tile_X4Y4_FrameStrobe_O[5] ,
    \Tile_X4Y4_FrameStrobe_O[4] ,
    \Tile_X4Y4_FrameStrobe_O[3] ,
    \Tile_X4Y4_FrameStrobe_O[2] ,
    \Tile_X4Y4_FrameStrobe_O[1] ,
    \Tile_X4Y4_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X4Y4_N1BEG[3] ,
    \Tile_X4Y4_N1BEG[2] ,
    \Tile_X4Y4_N1BEG[1] ,
    \Tile_X4Y4_N1BEG[0] }),
    .N1END({\Tile_X4Y5_N1BEG[3] ,
    \Tile_X4Y5_N1BEG[2] ,
    \Tile_X4Y5_N1BEG[1] ,
    \Tile_X4Y5_N1BEG[0] }),
    .N2BEG({\Tile_X4Y4_N2BEG[7] ,
    \Tile_X4Y4_N2BEG[6] ,
    \Tile_X4Y4_N2BEG[5] ,
    \Tile_X4Y4_N2BEG[4] ,
    \Tile_X4Y4_N2BEG[3] ,
    \Tile_X4Y4_N2BEG[2] ,
    \Tile_X4Y4_N2BEG[1] ,
    \Tile_X4Y4_N2BEG[0] }),
    .N2BEGb({\Tile_X4Y4_N2BEGb[7] ,
    \Tile_X4Y4_N2BEGb[6] ,
    \Tile_X4Y4_N2BEGb[5] ,
    \Tile_X4Y4_N2BEGb[4] ,
    \Tile_X4Y4_N2BEGb[3] ,
    \Tile_X4Y4_N2BEGb[2] ,
    \Tile_X4Y4_N2BEGb[1] ,
    \Tile_X4Y4_N2BEGb[0] }),
    .N2END({\Tile_X4Y5_N2BEGb[7] ,
    \Tile_X4Y5_N2BEGb[6] ,
    \Tile_X4Y5_N2BEGb[5] ,
    \Tile_X4Y5_N2BEGb[4] ,
    \Tile_X4Y5_N2BEGb[3] ,
    \Tile_X4Y5_N2BEGb[2] ,
    \Tile_X4Y5_N2BEGb[1] ,
    \Tile_X4Y5_N2BEGb[0] }),
    .N2MID({\Tile_X4Y5_N2BEG[7] ,
    \Tile_X4Y5_N2BEG[6] ,
    \Tile_X4Y5_N2BEG[5] ,
    \Tile_X4Y5_N2BEG[4] ,
    \Tile_X4Y5_N2BEG[3] ,
    \Tile_X4Y5_N2BEG[2] ,
    \Tile_X4Y5_N2BEG[1] ,
    \Tile_X4Y5_N2BEG[0] }),
    .N4BEG({\Tile_X4Y4_N4BEG[15] ,
    \Tile_X4Y4_N4BEG[14] ,
    \Tile_X4Y4_N4BEG[13] ,
    \Tile_X4Y4_N4BEG[12] ,
    \Tile_X4Y4_N4BEG[11] ,
    \Tile_X4Y4_N4BEG[10] ,
    \Tile_X4Y4_N4BEG[9] ,
    \Tile_X4Y4_N4BEG[8] ,
    \Tile_X4Y4_N4BEG[7] ,
    \Tile_X4Y4_N4BEG[6] ,
    \Tile_X4Y4_N4BEG[5] ,
    \Tile_X4Y4_N4BEG[4] ,
    \Tile_X4Y4_N4BEG[3] ,
    \Tile_X4Y4_N4BEG[2] ,
    \Tile_X4Y4_N4BEG[1] ,
    \Tile_X4Y4_N4BEG[0] }),
    .N4END({\Tile_X4Y5_N4BEG[15] ,
    \Tile_X4Y5_N4BEG[14] ,
    \Tile_X4Y5_N4BEG[13] ,
    \Tile_X4Y5_N4BEG[12] ,
    \Tile_X4Y5_N4BEG[11] ,
    \Tile_X4Y5_N4BEG[10] ,
    \Tile_X4Y5_N4BEG[9] ,
    \Tile_X4Y5_N4BEG[8] ,
    \Tile_X4Y5_N4BEG[7] ,
    \Tile_X4Y5_N4BEG[6] ,
    \Tile_X4Y5_N4BEG[5] ,
    \Tile_X4Y5_N4BEG[4] ,
    \Tile_X4Y5_N4BEG[3] ,
    \Tile_X4Y5_N4BEG[2] ,
    \Tile_X4Y5_N4BEG[1] ,
    \Tile_X4Y5_N4BEG[0] }),
    .NN4BEG({\Tile_X4Y4_NN4BEG[15] ,
    \Tile_X4Y4_NN4BEG[14] ,
    \Tile_X4Y4_NN4BEG[13] ,
    \Tile_X4Y4_NN4BEG[12] ,
    \Tile_X4Y4_NN4BEG[11] ,
    \Tile_X4Y4_NN4BEG[10] ,
    \Tile_X4Y4_NN4BEG[9] ,
    \Tile_X4Y4_NN4BEG[8] ,
    \Tile_X4Y4_NN4BEG[7] ,
    \Tile_X4Y4_NN4BEG[6] ,
    \Tile_X4Y4_NN4BEG[5] ,
    \Tile_X4Y4_NN4BEG[4] ,
    \Tile_X4Y4_NN4BEG[3] ,
    \Tile_X4Y4_NN4BEG[2] ,
    \Tile_X4Y4_NN4BEG[1] ,
    \Tile_X4Y4_NN4BEG[0] }),
    .NN4END({\Tile_X4Y5_NN4BEG[15] ,
    \Tile_X4Y5_NN4BEG[14] ,
    \Tile_X4Y5_NN4BEG[13] ,
    \Tile_X4Y5_NN4BEG[12] ,
    \Tile_X4Y5_NN4BEG[11] ,
    \Tile_X4Y5_NN4BEG[10] ,
    \Tile_X4Y5_NN4BEG[9] ,
    \Tile_X4Y5_NN4BEG[8] ,
    \Tile_X4Y5_NN4BEG[7] ,
    \Tile_X4Y5_NN4BEG[6] ,
    \Tile_X4Y5_NN4BEG[5] ,
    \Tile_X4Y5_NN4BEG[4] ,
    \Tile_X4Y5_NN4BEG[3] ,
    \Tile_X4Y5_NN4BEG[2] ,
    \Tile_X4Y5_NN4BEG[1] ,
    \Tile_X4Y5_NN4BEG[0] }),
    .S1BEG({\Tile_X4Y4_S1BEG[3] ,
    \Tile_X4Y4_S1BEG[2] ,
    \Tile_X4Y4_S1BEG[1] ,
    \Tile_X4Y4_S1BEG[0] }),
    .S1END({\Tile_X4Y3_S1BEG[3] ,
    \Tile_X4Y3_S1BEG[2] ,
    \Tile_X4Y3_S1BEG[1] ,
    \Tile_X4Y3_S1BEG[0] }),
    .S2BEG({\Tile_X4Y4_S2BEG[7] ,
    \Tile_X4Y4_S2BEG[6] ,
    \Tile_X4Y4_S2BEG[5] ,
    \Tile_X4Y4_S2BEG[4] ,
    \Tile_X4Y4_S2BEG[3] ,
    \Tile_X4Y4_S2BEG[2] ,
    \Tile_X4Y4_S2BEG[1] ,
    \Tile_X4Y4_S2BEG[0] }),
    .S2BEGb({\Tile_X4Y4_S2BEGb[7] ,
    \Tile_X4Y4_S2BEGb[6] ,
    \Tile_X4Y4_S2BEGb[5] ,
    \Tile_X4Y4_S2BEGb[4] ,
    \Tile_X4Y4_S2BEGb[3] ,
    \Tile_X4Y4_S2BEGb[2] ,
    \Tile_X4Y4_S2BEGb[1] ,
    \Tile_X4Y4_S2BEGb[0] }),
    .S2END({\Tile_X4Y3_S2BEGb[7] ,
    \Tile_X4Y3_S2BEGb[6] ,
    \Tile_X4Y3_S2BEGb[5] ,
    \Tile_X4Y3_S2BEGb[4] ,
    \Tile_X4Y3_S2BEGb[3] ,
    \Tile_X4Y3_S2BEGb[2] ,
    \Tile_X4Y3_S2BEGb[1] ,
    \Tile_X4Y3_S2BEGb[0] }),
    .S2MID({\Tile_X4Y3_S2BEG[7] ,
    \Tile_X4Y3_S2BEG[6] ,
    \Tile_X4Y3_S2BEG[5] ,
    \Tile_X4Y3_S2BEG[4] ,
    \Tile_X4Y3_S2BEG[3] ,
    \Tile_X4Y3_S2BEG[2] ,
    \Tile_X4Y3_S2BEG[1] ,
    \Tile_X4Y3_S2BEG[0] }),
    .S4BEG({\Tile_X4Y4_S4BEG[15] ,
    \Tile_X4Y4_S4BEG[14] ,
    \Tile_X4Y4_S4BEG[13] ,
    \Tile_X4Y4_S4BEG[12] ,
    \Tile_X4Y4_S4BEG[11] ,
    \Tile_X4Y4_S4BEG[10] ,
    \Tile_X4Y4_S4BEG[9] ,
    \Tile_X4Y4_S4BEG[8] ,
    \Tile_X4Y4_S4BEG[7] ,
    \Tile_X4Y4_S4BEG[6] ,
    \Tile_X4Y4_S4BEG[5] ,
    \Tile_X4Y4_S4BEG[4] ,
    \Tile_X4Y4_S4BEG[3] ,
    \Tile_X4Y4_S4BEG[2] ,
    \Tile_X4Y4_S4BEG[1] ,
    \Tile_X4Y4_S4BEG[0] }),
    .S4END({\Tile_X4Y3_S4BEG[15] ,
    \Tile_X4Y3_S4BEG[14] ,
    \Tile_X4Y3_S4BEG[13] ,
    \Tile_X4Y3_S4BEG[12] ,
    \Tile_X4Y3_S4BEG[11] ,
    \Tile_X4Y3_S4BEG[10] ,
    \Tile_X4Y3_S4BEG[9] ,
    \Tile_X4Y3_S4BEG[8] ,
    \Tile_X4Y3_S4BEG[7] ,
    \Tile_X4Y3_S4BEG[6] ,
    \Tile_X4Y3_S4BEG[5] ,
    \Tile_X4Y3_S4BEG[4] ,
    \Tile_X4Y3_S4BEG[3] ,
    \Tile_X4Y3_S4BEG[2] ,
    \Tile_X4Y3_S4BEG[1] ,
    \Tile_X4Y3_S4BEG[0] }),
    .SS4BEG({\Tile_X4Y4_SS4BEG[15] ,
    \Tile_X4Y4_SS4BEG[14] ,
    \Tile_X4Y4_SS4BEG[13] ,
    \Tile_X4Y4_SS4BEG[12] ,
    \Tile_X4Y4_SS4BEG[11] ,
    \Tile_X4Y4_SS4BEG[10] ,
    \Tile_X4Y4_SS4BEG[9] ,
    \Tile_X4Y4_SS4BEG[8] ,
    \Tile_X4Y4_SS4BEG[7] ,
    \Tile_X4Y4_SS4BEG[6] ,
    \Tile_X4Y4_SS4BEG[5] ,
    \Tile_X4Y4_SS4BEG[4] ,
    \Tile_X4Y4_SS4BEG[3] ,
    \Tile_X4Y4_SS4BEG[2] ,
    \Tile_X4Y4_SS4BEG[1] ,
    \Tile_X4Y4_SS4BEG[0] }),
    .SS4END({\Tile_X4Y3_SS4BEG[15] ,
    \Tile_X4Y3_SS4BEG[14] ,
    \Tile_X4Y3_SS4BEG[13] ,
    \Tile_X4Y3_SS4BEG[12] ,
    \Tile_X4Y3_SS4BEG[11] ,
    \Tile_X4Y3_SS4BEG[10] ,
    \Tile_X4Y3_SS4BEG[9] ,
    \Tile_X4Y3_SS4BEG[8] ,
    \Tile_X4Y3_SS4BEG[7] ,
    \Tile_X4Y3_SS4BEG[6] ,
    \Tile_X4Y3_SS4BEG[5] ,
    \Tile_X4Y3_SS4BEG[4] ,
    \Tile_X4Y3_SS4BEG[3] ,
    \Tile_X4Y3_SS4BEG[2] ,
    \Tile_X4Y3_SS4BEG[1] ,
    \Tile_X4Y3_SS4BEG[0] }),
    .W1BEG({\Tile_X4Y4_W1BEG[3] ,
    \Tile_X4Y4_W1BEG[2] ,
    \Tile_X4Y4_W1BEG[1] ,
    \Tile_X4Y4_W1BEG[0] }),
    .W1END({\Tile_X5Y4_W1BEG[3] ,
    \Tile_X5Y4_W1BEG[2] ,
    \Tile_X5Y4_W1BEG[1] ,
    \Tile_X5Y4_W1BEG[0] }),
    .W2BEG({\Tile_X4Y4_W2BEG[7] ,
    \Tile_X4Y4_W2BEG[6] ,
    \Tile_X4Y4_W2BEG[5] ,
    \Tile_X4Y4_W2BEG[4] ,
    \Tile_X4Y4_W2BEG[3] ,
    \Tile_X4Y4_W2BEG[2] ,
    \Tile_X4Y4_W2BEG[1] ,
    \Tile_X4Y4_W2BEG[0] }),
    .W2BEGb({\Tile_X4Y4_W2BEGb[7] ,
    \Tile_X4Y4_W2BEGb[6] ,
    \Tile_X4Y4_W2BEGb[5] ,
    \Tile_X4Y4_W2BEGb[4] ,
    \Tile_X4Y4_W2BEGb[3] ,
    \Tile_X4Y4_W2BEGb[2] ,
    \Tile_X4Y4_W2BEGb[1] ,
    \Tile_X4Y4_W2BEGb[0] }),
    .W2END({\Tile_X5Y4_W2BEGb[7] ,
    \Tile_X5Y4_W2BEGb[6] ,
    \Tile_X5Y4_W2BEGb[5] ,
    \Tile_X5Y4_W2BEGb[4] ,
    \Tile_X5Y4_W2BEGb[3] ,
    \Tile_X5Y4_W2BEGb[2] ,
    \Tile_X5Y4_W2BEGb[1] ,
    \Tile_X5Y4_W2BEGb[0] }),
    .W2MID({\Tile_X5Y4_W2BEG[7] ,
    \Tile_X5Y4_W2BEG[6] ,
    \Tile_X5Y4_W2BEG[5] ,
    \Tile_X5Y4_W2BEG[4] ,
    \Tile_X5Y4_W2BEG[3] ,
    \Tile_X5Y4_W2BEG[2] ,
    \Tile_X5Y4_W2BEG[1] ,
    \Tile_X5Y4_W2BEG[0] }),
    .W6BEG({\Tile_X4Y4_W6BEG[11] ,
    \Tile_X4Y4_W6BEG[10] ,
    \Tile_X4Y4_W6BEG[9] ,
    \Tile_X4Y4_W6BEG[8] ,
    \Tile_X4Y4_W6BEG[7] ,
    \Tile_X4Y4_W6BEG[6] ,
    \Tile_X4Y4_W6BEG[5] ,
    \Tile_X4Y4_W6BEG[4] ,
    \Tile_X4Y4_W6BEG[3] ,
    \Tile_X4Y4_W6BEG[2] ,
    \Tile_X4Y4_W6BEG[1] ,
    \Tile_X4Y4_W6BEG[0] }),
    .W6END({\Tile_X5Y4_W6BEG[11] ,
    \Tile_X5Y4_W6BEG[10] ,
    \Tile_X5Y4_W6BEG[9] ,
    \Tile_X5Y4_W6BEG[8] ,
    \Tile_X5Y4_W6BEG[7] ,
    \Tile_X5Y4_W6BEG[6] ,
    \Tile_X5Y4_W6BEG[5] ,
    \Tile_X5Y4_W6BEG[4] ,
    \Tile_X5Y4_W6BEG[3] ,
    \Tile_X5Y4_W6BEG[2] ,
    \Tile_X5Y4_W6BEG[1] ,
    \Tile_X5Y4_W6BEG[0] }),
    .WW4BEG({\Tile_X4Y4_WW4BEG[15] ,
    \Tile_X4Y4_WW4BEG[14] ,
    \Tile_X4Y4_WW4BEG[13] ,
    \Tile_X4Y4_WW4BEG[12] ,
    \Tile_X4Y4_WW4BEG[11] ,
    \Tile_X4Y4_WW4BEG[10] ,
    \Tile_X4Y4_WW4BEG[9] ,
    \Tile_X4Y4_WW4BEG[8] ,
    \Tile_X4Y4_WW4BEG[7] ,
    \Tile_X4Y4_WW4BEG[6] ,
    \Tile_X4Y4_WW4BEG[5] ,
    \Tile_X4Y4_WW4BEG[4] ,
    \Tile_X4Y4_WW4BEG[3] ,
    \Tile_X4Y4_WW4BEG[2] ,
    \Tile_X4Y4_WW4BEG[1] ,
    \Tile_X4Y4_WW4BEG[0] }),
    .WW4END({\Tile_X5Y4_WW4BEG[15] ,
    \Tile_X5Y4_WW4BEG[14] ,
    \Tile_X5Y4_WW4BEG[13] ,
    \Tile_X5Y4_WW4BEG[12] ,
    \Tile_X5Y4_WW4BEG[11] ,
    \Tile_X5Y4_WW4BEG[10] ,
    \Tile_X5Y4_WW4BEG[9] ,
    \Tile_X5Y4_WW4BEG[8] ,
    \Tile_X5Y4_WW4BEG[7] ,
    \Tile_X5Y4_WW4BEG[6] ,
    \Tile_X5Y4_WW4BEG[5] ,
    \Tile_X5Y4_WW4BEG[4] ,
    \Tile_X5Y4_WW4BEG[3] ,
    \Tile_X5Y4_WW4BEG[2] ,
    \Tile_X5Y4_WW4BEG[1] ,
    \Tile_X5Y4_WW4BEG[0] }));
 LUT4AB Tile_X4Y5_LUT4AB (.Ci(Tile_X4Y6_Co),
    .Co(Tile_X4Y5_Co),
    .UserCLK(Tile_X4Y6_UserCLKo),
    .UserCLKo(Tile_X4Y5_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X4Y5_E1BEG[3] ,
    \Tile_X4Y5_E1BEG[2] ,
    \Tile_X4Y5_E1BEG[1] ,
    \Tile_X4Y5_E1BEG[0] }),
    .E1END({\Tile_X3Y5_E1BEG[3] ,
    \Tile_X3Y5_E1BEG[2] ,
    \Tile_X3Y5_E1BEG[1] ,
    \Tile_X3Y5_E1BEG[0] }),
    .E2BEG({\Tile_X4Y5_E2BEG[7] ,
    \Tile_X4Y5_E2BEG[6] ,
    \Tile_X4Y5_E2BEG[5] ,
    \Tile_X4Y5_E2BEG[4] ,
    \Tile_X4Y5_E2BEG[3] ,
    \Tile_X4Y5_E2BEG[2] ,
    \Tile_X4Y5_E2BEG[1] ,
    \Tile_X4Y5_E2BEG[0] }),
    .E2BEGb({\Tile_X4Y5_E2BEGb[7] ,
    \Tile_X4Y5_E2BEGb[6] ,
    \Tile_X4Y5_E2BEGb[5] ,
    \Tile_X4Y5_E2BEGb[4] ,
    \Tile_X4Y5_E2BEGb[3] ,
    \Tile_X4Y5_E2BEGb[2] ,
    \Tile_X4Y5_E2BEGb[1] ,
    \Tile_X4Y5_E2BEGb[0] }),
    .E2END({\Tile_X3Y5_E2BEGb[7] ,
    \Tile_X3Y5_E2BEGb[6] ,
    \Tile_X3Y5_E2BEGb[5] ,
    \Tile_X3Y5_E2BEGb[4] ,
    \Tile_X3Y5_E2BEGb[3] ,
    \Tile_X3Y5_E2BEGb[2] ,
    \Tile_X3Y5_E2BEGb[1] ,
    \Tile_X3Y5_E2BEGb[0] }),
    .E2MID({\Tile_X3Y5_E2BEG[7] ,
    \Tile_X3Y5_E2BEG[6] ,
    \Tile_X3Y5_E2BEG[5] ,
    \Tile_X3Y5_E2BEG[4] ,
    \Tile_X3Y5_E2BEG[3] ,
    \Tile_X3Y5_E2BEG[2] ,
    \Tile_X3Y5_E2BEG[1] ,
    \Tile_X3Y5_E2BEG[0] }),
    .E6BEG({\Tile_X4Y5_E6BEG[11] ,
    \Tile_X4Y5_E6BEG[10] ,
    \Tile_X4Y5_E6BEG[9] ,
    \Tile_X4Y5_E6BEG[8] ,
    \Tile_X4Y5_E6BEG[7] ,
    \Tile_X4Y5_E6BEG[6] ,
    \Tile_X4Y5_E6BEG[5] ,
    \Tile_X4Y5_E6BEG[4] ,
    \Tile_X4Y5_E6BEG[3] ,
    \Tile_X4Y5_E6BEG[2] ,
    \Tile_X4Y5_E6BEG[1] ,
    \Tile_X4Y5_E6BEG[0] }),
    .E6END({\Tile_X3Y5_E6BEG[11] ,
    \Tile_X3Y5_E6BEG[10] ,
    \Tile_X3Y5_E6BEG[9] ,
    \Tile_X3Y5_E6BEG[8] ,
    \Tile_X3Y5_E6BEG[7] ,
    \Tile_X3Y5_E6BEG[6] ,
    \Tile_X3Y5_E6BEG[5] ,
    \Tile_X3Y5_E6BEG[4] ,
    \Tile_X3Y5_E6BEG[3] ,
    \Tile_X3Y5_E6BEG[2] ,
    \Tile_X3Y5_E6BEG[1] ,
    \Tile_X3Y5_E6BEG[0] }),
    .EE4BEG({\Tile_X4Y5_EE4BEG[15] ,
    \Tile_X4Y5_EE4BEG[14] ,
    \Tile_X4Y5_EE4BEG[13] ,
    \Tile_X4Y5_EE4BEG[12] ,
    \Tile_X4Y5_EE4BEG[11] ,
    \Tile_X4Y5_EE4BEG[10] ,
    \Tile_X4Y5_EE4BEG[9] ,
    \Tile_X4Y5_EE4BEG[8] ,
    \Tile_X4Y5_EE4BEG[7] ,
    \Tile_X4Y5_EE4BEG[6] ,
    \Tile_X4Y5_EE4BEG[5] ,
    \Tile_X4Y5_EE4BEG[4] ,
    \Tile_X4Y5_EE4BEG[3] ,
    \Tile_X4Y5_EE4BEG[2] ,
    \Tile_X4Y5_EE4BEG[1] ,
    \Tile_X4Y5_EE4BEG[0] }),
    .EE4END({\Tile_X3Y5_EE4BEG[15] ,
    \Tile_X3Y5_EE4BEG[14] ,
    \Tile_X3Y5_EE4BEG[13] ,
    \Tile_X3Y5_EE4BEG[12] ,
    \Tile_X3Y5_EE4BEG[11] ,
    \Tile_X3Y5_EE4BEG[10] ,
    \Tile_X3Y5_EE4BEG[9] ,
    \Tile_X3Y5_EE4BEG[8] ,
    \Tile_X3Y5_EE4BEG[7] ,
    \Tile_X3Y5_EE4BEG[6] ,
    \Tile_X3Y5_EE4BEG[5] ,
    \Tile_X3Y5_EE4BEG[4] ,
    \Tile_X3Y5_EE4BEG[3] ,
    \Tile_X3Y5_EE4BEG[2] ,
    \Tile_X3Y5_EE4BEG[1] ,
    \Tile_X3Y5_EE4BEG[0] }),
    .FrameData({\Tile_X3Y5_FrameData_O[31] ,
    \Tile_X3Y5_FrameData_O[30] ,
    \Tile_X3Y5_FrameData_O[29] ,
    \Tile_X3Y5_FrameData_O[28] ,
    \Tile_X3Y5_FrameData_O[27] ,
    \Tile_X3Y5_FrameData_O[26] ,
    \Tile_X3Y5_FrameData_O[25] ,
    \Tile_X3Y5_FrameData_O[24] ,
    \Tile_X3Y5_FrameData_O[23] ,
    \Tile_X3Y5_FrameData_O[22] ,
    \Tile_X3Y5_FrameData_O[21] ,
    \Tile_X3Y5_FrameData_O[20] ,
    \Tile_X3Y5_FrameData_O[19] ,
    \Tile_X3Y5_FrameData_O[18] ,
    \Tile_X3Y5_FrameData_O[17] ,
    \Tile_X3Y5_FrameData_O[16] ,
    \Tile_X3Y5_FrameData_O[15] ,
    \Tile_X3Y5_FrameData_O[14] ,
    \Tile_X3Y5_FrameData_O[13] ,
    \Tile_X3Y5_FrameData_O[12] ,
    \Tile_X3Y5_FrameData_O[11] ,
    \Tile_X3Y5_FrameData_O[10] ,
    \Tile_X3Y5_FrameData_O[9] ,
    \Tile_X3Y5_FrameData_O[8] ,
    \Tile_X3Y5_FrameData_O[7] ,
    \Tile_X3Y5_FrameData_O[6] ,
    \Tile_X3Y5_FrameData_O[5] ,
    \Tile_X3Y5_FrameData_O[4] ,
    \Tile_X3Y5_FrameData_O[3] ,
    \Tile_X3Y5_FrameData_O[2] ,
    \Tile_X3Y5_FrameData_O[1] ,
    \Tile_X3Y5_FrameData_O[0] }),
    .FrameData_O({\Tile_X4Y5_FrameData_O[31] ,
    \Tile_X4Y5_FrameData_O[30] ,
    \Tile_X4Y5_FrameData_O[29] ,
    \Tile_X4Y5_FrameData_O[28] ,
    \Tile_X4Y5_FrameData_O[27] ,
    \Tile_X4Y5_FrameData_O[26] ,
    \Tile_X4Y5_FrameData_O[25] ,
    \Tile_X4Y5_FrameData_O[24] ,
    \Tile_X4Y5_FrameData_O[23] ,
    \Tile_X4Y5_FrameData_O[22] ,
    \Tile_X4Y5_FrameData_O[21] ,
    \Tile_X4Y5_FrameData_O[20] ,
    \Tile_X4Y5_FrameData_O[19] ,
    \Tile_X4Y5_FrameData_O[18] ,
    \Tile_X4Y5_FrameData_O[17] ,
    \Tile_X4Y5_FrameData_O[16] ,
    \Tile_X4Y5_FrameData_O[15] ,
    \Tile_X4Y5_FrameData_O[14] ,
    \Tile_X4Y5_FrameData_O[13] ,
    \Tile_X4Y5_FrameData_O[12] ,
    \Tile_X4Y5_FrameData_O[11] ,
    \Tile_X4Y5_FrameData_O[10] ,
    \Tile_X4Y5_FrameData_O[9] ,
    \Tile_X4Y5_FrameData_O[8] ,
    \Tile_X4Y5_FrameData_O[7] ,
    \Tile_X4Y5_FrameData_O[6] ,
    \Tile_X4Y5_FrameData_O[5] ,
    \Tile_X4Y5_FrameData_O[4] ,
    \Tile_X4Y5_FrameData_O[3] ,
    \Tile_X4Y5_FrameData_O[2] ,
    \Tile_X4Y5_FrameData_O[1] ,
    \Tile_X4Y5_FrameData_O[0] }),
    .FrameStrobe({\Tile_X4Y6_FrameStrobe_O[19] ,
    \Tile_X4Y6_FrameStrobe_O[18] ,
    \Tile_X4Y6_FrameStrobe_O[17] ,
    \Tile_X4Y6_FrameStrobe_O[16] ,
    \Tile_X4Y6_FrameStrobe_O[15] ,
    \Tile_X4Y6_FrameStrobe_O[14] ,
    \Tile_X4Y6_FrameStrobe_O[13] ,
    \Tile_X4Y6_FrameStrobe_O[12] ,
    \Tile_X4Y6_FrameStrobe_O[11] ,
    \Tile_X4Y6_FrameStrobe_O[10] ,
    \Tile_X4Y6_FrameStrobe_O[9] ,
    \Tile_X4Y6_FrameStrobe_O[8] ,
    \Tile_X4Y6_FrameStrobe_O[7] ,
    \Tile_X4Y6_FrameStrobe_O[6] ,
    \Tile_X4Y6_FrameStrobe_O[5] ,
    \Tile_X4Y6_FrameStrobe_O[4] ,
    \Tile_X4Y6_FrameStrobe_O[3] ,
    \Tile_X4Y6_FrameStrobe_O[2] ,
    \Tile_X4Y6_FrameStrobe_O[1] ,
    \Tile_X4Y6_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X4Y5_FrameStrobe_O[19] ,
    \Tile_X4Y5_FrameStrobe_O[18] ,
    \Tile_X4Y5_FrameStrobe_O[17] ,
    \Tile_X4Y5_FrameStrobe_O[16] ,
    \Tile_X4Y5_FrameStrobe_O[15] ,
    \Tile_X4Y5_FrameStrobe_O[14] ,
    \Tile_X4Y5_FrameStrobe_O[13] ,
    \Tile_X4Y5_FrameStrobe_O[12] ,
    \Tile_X4Y5_FrameStrobe_O[11] ,
    \Tile_X4Y5_FrameStrobe_O[10] ,
    \Tile_X4Y5_FrameStrobe_O[9] ,
    \Tile_X4Y5_FrameStrobe_O[8] ,
    \Tile_X4Y5_FrameStrobe_O[7] ,
    \Tile_X4Y5_FrameStrobe_O[6] ,
    \Tile_X4Y5_FrameStrobe_O[5] ,
    \Tile_X4Y5_FrameStrobe_O[4] ,
    \Tile_X4Y5_FrameStrobe_O[3] ,
    \Tile_X4Y5_FrameStrobe_O[2] ,
    \Tile_X4Y5_FrameStrobe_O[1] ,
    \Tile_X4Y5_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X4Y5_N1BEG[3] ,
    \Tile_X4Y5_N1BEG[2] ,
    \Tile_X4Y5_N1BEG[1] ,
    \Tile_X4Y5_N1BEG[0] }),
    .N1END({\Tile_X4Y6_N1BEG[3] ,
    \Tile_X4Y6_N1BEG[2] ,
    \Tile_X4Y6_N1BEG[1] ,
    \Tile_X4Y6_N1BEG[0] }),
    .N2BEG({\Tile_X4Y5_N2BEG[7] ,
    \Tile_X4Y5_N2BEG[6] ,
    \Tile_X4Y5_N2BEG[5] ,
    \Tile_X4Y5_N2BEG[4] ,
    \Tile_X4Y5_N2BEG[3] ,
    \Tile_X4Y5_N2BEG[2] ,
    \Tile_X4Y5_N2BEG[1] ,
    \Tile_X4Y5_N2BEG[0] }),
    .N2BEGb({\Tile_X4Y5_N2BEGb[7] ,
    \Tile_X4Y5_N2BEGb[6] ,
    \Tile_X4Y5_N2BEGb[5] ,
    \Tile_X4Y5_N2BEGb[4] ,
    \Tile_X4Y5_N2BEGb[3] ,
    \Tile_X4Y5_N2BEGb[2] ,
    \Tile_X4Y5_N2BEGb[1] ,
    \Tile_X4Y5_N2BEGb[0] }),
    .N2END({\Tile_X4Y6_N2BEGb[7] ,
    \Tile_X4Y6_N2BEGb[6] ,
    \Tile_X4Y6_N2BEGb[5] ,
    \Tile_X4Y6_N2BEGb[4] ,
    \Tile_X4Y6_N2BEGb[3] ,
    \Tile_X4Y6_N2BEGb[2] ,
    \Tile_X4Y6_N2BEGb[1] ,
    \Tile_X4Y6_N2BEGb[0] }),
    .N2MID({\Tile_X4Y6_N2BEG[7] ,
    \Tile_X4Y6_N2BEG[6] ,
    \Tile_X4Y6_N2BEG[5] ,
    \Tile_X4Y6_N2BEG[4] ,
    \Tile_X4Y6_N2BEG[3] ,
    \Tile_X4Y6_N2BEG[2] ,
    \Tile_X4Y6_N2BEG[1] ,
    \Tile_X4Y6_N2BEG[0] }),
    .N4BEG({\Tile_X4Y5_N4BEG[15] ,
    \Tile_X4Y5_N4BEG[14] ,
    \Tile_X4Y5_N4BEG[13] ,
    \Tile_X4Y5_N4BEG[12] ,
    \Tile_X4Y5_N4BEG[11] ,
    \Tile_X4Y5_N4BEG[10] ,
    \Tile_X4Y5_N4BEG[9] ,
    \Tile_X4Y5_N4BEG[8] ,
    \Tile_X4Y5_N4BEG[7] ,
    \Tile_X4Y5_N4BEG[6] ,
    \Tile_X4Y5_N4BEG[5] ,
    \Tile_X4Y5_N4BEG[4] ,
    \Tile_X4Y5_N4BEG[3] ,
    \Tile_X4Y5_N4BEG[2] ,
    \Tile_X4Y5_N4BEG[1] ,
    \Tile_X4Y5_N4BEG[0] }),
    .N4END({\Tile_X4Y6_N4BEG[15] ,
    \Tile_X4Y6_N4BEG[14] ,
    \Tile_X4Y6_N4BEG[13] ,
    \Tile_X4Y6_N4BEG[12] ,
    \Tile_X4Y6_N4BEG[11] ,
    \Tile_X4Y6_N4BEG[10] ,
    \Tile_X4Y6_N4BEG[9] ,
    \Tile_X4Y6_N4BEG[8] ,
    \Tile_X4Y6_N4BEG[7] ,
    \Tile_X4Y6_N4BEG[6] ,
    \Tile_X4Y6_N4BEG[5] ,
    \Tile_X4Y6_N4BEG[4] ,
    \Tile_X4Y6_N4BEG[3] ,
    \Tile_X4Y6_N4BEG[2] ,
    \Tile_X4Y6_N4BEG[1] ,
    \Tile_X4Y6_N4BEG[0] }),
    .NN4BEG({\Tile_X4Y5_NN4BEG[15] ,
    \Tile_X4Y5_NN4BEG[14] ,
    \Tile_X4Y5_NN4BEG[13] ,
    \Tile_X4Y5_NN4BEG[12] ,
    \Tile_X4Y5_NN4BEG[11] ,
    \Tile_X4Y5_NN4BEG[10] ,
    \Tile_X4Y5_NN4BEG[9] ,
    \Tile_X4Y5_NN4BEG[8] ,
    \Tile_X4Y5_NN4BEG[7] ,
    \Tile_X4Y5_NN4BEG[6] ,
    \Tile_X4Y5_NN4BEG[5] ,
    \Tile_X4Y5_NN4BEG[4] ,
    \Tile_X4Y5_NN4BEG[3] ,
    \Tile_X4Y5_NN4BEG[2] ,
    \Tile_X4Y5_NN4BEG[1] ,
    \Tile_X4Y5_NN4BEG[0] }),
    .NN4END({\Tile_X4Y6_NN4BEG[15] ,
    \Tile_X4Y6_NN4BEG[14] ,
    \Tile_X4Y6_NN4BEG[13] ,
    \Tile_X4Y6_NN4BEG[12] ,
    \Tile_X4Y6_NN4BEG[11] ,
    \Tile_X4Y6_NN4BEG[10] ,
    \Tile_X4Y6_NN4BEG[9] ,
    \Tile_X4Y6_NN4BEG[8] ,
    \Tile_X4Y6_NN4BEG[7] ,
    \Tile_X4Y6_NN4BEG[6] ,
    \Tile_X4Y6_NN4BEG[5] ,
    \Tile_X4Y6_NN4BEG[4] ,
    \Tile_X4Y6_NN4BEG[3] ,
    \Tile_X4Y6_NN4BEG[2] ,
    \Tile_X4Y6_NN4BEG[1] ,
    \Tile_X4Y6_NN4BEG[0] }),
    .S1BEG({\Tile_X4Y5_S1BEG[3] ,
    \Tile_X4Y5_S1BEG[2] ,
    \Tile_X4Y5_S1BEG[1] ,
    \Tile_X4Y5_S1BEG[0] }),
    .S1END({\Tile_X4Y4_S1BEG[3] ,
    \Tile_X4Y4_S1BEG[2] ,
    \Tile_X4Y4_S1BEG[1] ,
    \Tile_X4Y4_S1BEG[0] }),
    .S2BEG({\Tile_X4Y5_S2BEG[7] ,
    \Tile_X4Y5_S2BEG[6] ,
    \Tile_X4Y5_S2BEG[5] ,
    \Tile_X4Y5_S2BEG[4] ,
    \Tile_X4Y5_S2BEG[3] ,
    \Tile_X4Y5_S2BEG[2] ,
    \Tile_X4Y5_S2BEG[1] ,
    \Tile_X4Y5_S2BEG[0] }),
    .S2BEGb({\Tile_X4Y5_S2BEGb[7] ,
    \Tile_X4Y5_S2BEGb[6] ,
    \Tile_X4Y5_S2BEGb[5] ,
    \Tile_X4Y5_S2BEGb[4] ,
    \Tile_X4Y5_S2BEGb[3] ,
    \Tile_X4Y5_S2BEGb[2] ,
    \Tile_X4Y5_S2BEGb[1] ,
    \Tile_X4Y5_S2BEGb[0] }),
    .S2END({\Tile_X4Y4_S2BEGb[7] ,
    \Tile_X4Y4_S2BEGb[6] ,
    \Tile_X4Y4_S2BEGb[5] ,
    \Tile_X4Y4_S2BEGb[4] ,
    \Tile_X4Y4_S2BEGb[3] ,
    \Tile_X4Y4_S2BEGb[2] ,
    \Tile_X4Y4_S2BEGb[1] ,
    \Tile_X4Y4_S2BEGb[0] }),
    .S2MID({\Tile_X4Y4_S2BEG[7] ,
    \Tile_X4Y4_S2BEG[6] ,
    \Tile_X4Y4_S2BEG[5] ,
    \Tile_X4Y4_S2BEG[4] ,
    \Tile_X4Y4_S2BEG[3] ,
    \Tile_X4Y4_S2BEG[2] ,
    \Tile_X4Y4_S2BEG[1] ,
    \Tile_X4Y4_S2BEG[0] }),
    .S4BEG({\Tile_X4Y5_S4BEG[15] ,
    \Tile_X4Y5_S4BEG[14] ,
    \Tile_X4Y5_S4BEG[13] ,
    \Tile_X4Y5_S4BEG[12] ,
    \Tile_X4Y5_S4BEG[11] ,
    \Tile_X4Y5_S4BEG[10] ,
    \Tile_X4Y5_S4BEG[9] ,
    \Tile_X4Y5_S4BEG[8] ,
    \Tile_X4Y5_S4BEG[7] ,
    \Tile_X4Y5_S4BEG[6] ,
    \Tile_X4Y5_S4BEG[5] ,
    \Tile_X4Y5_S4BEG[4] ,
    \Tile_X4Y5_S4BEG[3] ,
    \Tile_X4Y5_S4BEG[2] ,
    \Tile_X4Y5_S4BEG[1] ,
    \Tile_X4Y5_S4BEG[0] }),
    .S4END({\Tile_X4Y4_S4BEG[15] ,
    \Tile_X4Y4_S4BEG[14] ,
    \Tile_X4Y4_S4BEG[13] ,
    \Tile_X4Y4_S4BEG[12] ,
    \Tile_X4Y4_S4BEG[11] ,
    \Tile_X4Y4_S4BEG[10] ,
    \Tile_X4Y4_S4BEG[9] ,
    \Tile_X4Y4_S4BEG[8] ,
    \Tile_X4Y4_S4BEG[7] ,
    \Tile_X4Y4_S4BEG[6] ,
    \Tile_X4Y4_S4BEG[5] ,
    \Tile_X4Y4_S4BEG[4] ,
    \Tile_X4Y4_S4BEG[3] ,
    \Tile_X4Y4_S4BEG[2] ,
    \Tile_X4Y4_S4BEG[1] ,
    \Tile_X4Y4_S4BEG[0] }),
    .SS4BEG({\Tile_X4Y5_SS4BEG[15] ,
    \Tile_X4Y5_SS4BEG[14] ,
    \Tile_X4Y5_SS4BEG[13] ,
    \Tile_X4Y5_SS4BEG[12] ,
    \Tile_X4Y5_SS4BEG[11] ,
    \Tile_X4Y5_SS4BEG[10] ,
    \Tile_X4Y5_SS4BEG[9] ,
    \Tile_X4Y5_SS4BEG[8] ,
    \Tile_X4Y5_SS4BEG[7] ,
    \Tile_X4Y5_SS4BEG[6] ,
    \Tile_X4Y5_SS4BEG[5] ,
    \Tile_X4Y5_SS4BEG[4] ,
    \Tile_X4Y5_SS4BEG[3] ,
    \Tile_X4Y5_SS4BEG[2] ,
    \Tile_X4Y5_SS4BEG[1] ,
    \Tile_X4Y5_SS4BEG[0] }),
    .SS4END({\Tile_X4Y4_SS4BEG[15] ,
    \Tile_X4Y4_SS4BEG[14] ,
    \Tile_X4Y4_SS4BEG[13] ,
    \Tile_X4Y4_SS4BEG[12] ,
    \Tile_X4Y4_SS4BEG[11] ,
    \Tile_X4Y4_SS4BEG[10] ,
    \Tile_X4Y4_SS4BEG[9] ,
    \Tile_X4Y4_SS4BEG[8] ,
    \Tile_X4Y4_SS4BEG[7] ,
    \Tile_X4Y4_SS4BEG[6] ,
    \Tile_X4Y4_SS4BEG[5] ,
    \Tile_X4Y4_SS4BEG[4] ,
    \Tile_X4Y4_SS4BEG[3] ,
    \Tile_X4Y4_SS4BEG[2] ,
    \Tile_X4Y4_SS4BEG[1] ,
    \Tile_X4Y4_SS4BEG[0] }),
    .W1BEG({\Tile_X4Y5_W1BEG[3] ,
    \Tile_X4Y5_W1BEG[2] ,
    \Tile_X4Y5_W1BEG[1] ,
    \Tile_X4Y5_W1BEG[0] }),
    .W1END({\Tile_X5Y5_W1BEG[3] ,
    \Tile_X5Y5_W1BEG[2] ,
    \Tile_X5Y5_W1BEG[1] ,
    \Tile_X5Y5_W1BEG[0] }),
    .W2BEG({\Tile_X4Y5_W2BEG[7] ,
    \Tile_X4Y5_W2BEG[6] ,
    \Tile_X4Y5_W2BEG[5] ,
    \Tile_X4Y5_W2BEG[4] ,
    \Tile_X4Y5_W2BEG[3] ,
    \Tile_X4Y5_W2BEG[2] ,
    \Tile_X4Y5_W2BEG[1] ,
    \Tile_X4Y5_W2BEG[0] }),
    .W2BEGb({\Tile_X4Y5_W2BEGb[7] ,
    \Tile_X4Y5_W2BEGb[6] ,
    \Tile_X4Y5_W2BEGb[5] ,
    \Tile_X4Y5_W2BEGb[4] ,
    \Tile_X4Y5_W2BEGb[3] ,
    \Tile_X4Y5_W2BEGb[2] ,
    \Tile_X4Y5_W2BEGb[1] ,
    \Tile_X4Y5_W2BEGb[0] }),
    .W2END({\Tile_X5Y5_W2BEGb[7] ,
    \Tile_X5Y5_W2BEGb[6] ,
    \Tile_X5Y5_W2BEGb[5] ,
    \Tile_X5Y5_W2BEGb[4] ,
    \Tile_X5Y5_W2BEGb[3] ,
    \Tile_X5Y5_W2BEGb[2] ,
    \Tile_X5Y5_W2BEGb[1] ,
    \Tile_X5Y5_W2BEGb[0] }),
    .W2MID({\Tile_X5Y5_W2BEG[7] ,
    \Tile_X5Y5_W2BEG[6] ,
    \Tile_X5Y5_W2BEG[5] ,
    \Tile_X5Y5_W2BEG[4] ,
    \Tile_X5Y5_W2BEG[3] ,
    \Tile_X5Y5_W2BEG[2] ,
    \Tile_X5Y5_W2BEG[1] ,
    \Tile_X5Y5_W2BEG[0] }),
    .W6BEG({\Tile_X4Y5_W6BEG[11] ,
    \Tile_X4Y5_W6BEG[10] ,
    \Tile_X4Y5_W6BEG[9] ,
    \Tile_X4Y5_W6BEG[8] ,
    \Tile_X4Y5_W6BEG[7] ,
    \Tile_X4Y5_W6BEG[6] ,
    \Tile_X4Y5_W6BEG[5] ,
    \Tile_X4Y5_W6BEG[4] ,
    \Tile_X4Y5_W6BEG[3] ,
    \Tile_X4Y5_W6BEG[2] ,
    \Tile_X4Y5_W6BEG[1] ,
    \Tile_X4Y5_W6BEG[0] }),
    .W6END({\Tile_X5Y5_W6BEG[11] ,
    \Tile_X5Y5_W6BEG[10] ,
    \Tile_X5Y5_W6BEG[9] ,
    \Tile_X5Y5_W6BEG[8] ,
    \Tile_X5Y5_W6BEG[7] ,
    \Tile_X5Y5_W6BEG[6] ,
    \Tile_X5Y5_W6BEG[5] ,
    \Tile_X5Y5_W6BEG[4] ,
    \Tile_X5Y5_W6BEG[3] ,
    \Tile_X5Y5_W6BEG[2] ,
    \Tile_X5Y5_W6BEG[1] ,
    \Tile_X5Y5_W6BEG[0] }),
    .WW4BEG({\Tile_X4Y5_WW4BEG[15] ,
    \Tile_X4Y5_WW4BEG[14] ,
    \Tile_X4Y5_WW4BEG[13] ,
    \Tile_X4Y5_WW4BEG[12] ,
    \Tile_X4Y5_WW4BEG[11] ,
    \Tile_X4Y5_WW4BEG[10] ,
    \Tile_X4Y5_WW4BEG[9] ,
    \Tile_X4Y5_WW4BEG[8] ,
    \Tile_X4Y5_WW4BEG[7] ,
    \Tile_X4Y5_WW4BEG[6] ,
    \Tile_X4Y5_WW4BEG[5] ,
    \Tile_X4Y5_WW4BEG[4] ,
    \Tile_X4Y5_WW4BEG[3] ,
    \Tile_X4Y5_WW4BEG[2] ,
    \Tile_X4Y5_WW4BEG[1] ,
    \Tile_X4Y5_WW4BEG[0] }),
    .WW4END({\Tile_X5Y5_WW4BEG[15] ,
    \Tile_X5Y5_WW4BEG[14] ,
    \Tile_X5Y5_WW4BEG[13] ,
    \Tile_X5Y5_WW4BEG[12] ,
    \Tile_X5Y5_WW4BEG[11] ,
    \Tile_X5Y5_WW4BEG[10] ,
    \Tile_X5Y5_WW4BEG[9] ,
    \Tile_X5Y5_WW4BEG[8] ,
    \Tile_X5Y5_WW4BEG[7] ,
    \Tile_X5Y5_WW4BEG[6] ,
    \Tile_X5Y5_WW4BEG[5] ,
    \Tile_X5Y5_WW4BEG[4] ,
    \Tile_X5Y5_WW4BEG[3] ,
    \Tile_X5Y5_WW4BEG[2] ,
    \Tile_X5Y5_WW4BEG[1] ,
    \Tile_X5Y5_WW4BEG[0] }));
 LUT4AB Tile_X4Y6_LUT4AB (.Ci(Tile_X4Y7_Co),
    .Co(Tile_X4Y6_Co),
    .UserCLK(Tile_X4Y7_UserCLKo),
    .UserCLKo(Tile_X4Y6_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X4Y6_E1BEG[3] ,
    \Tile_X4Y6_E1BEG[2] ,
    \Tile_X4Y6_E1BEG[1] ,
    \Tile_X4Y6_E1BEG[0] }),
    .E1END({\Tile_X3Y6_E1BEG[3] ,
    \Tile_X3Y6_E1BEG[2] ,
    \Tile_X3Y6_E1BEG[1] ,
    \Tile_X3Y6_E1BEG[0] }),
    .E2BEG({\Tile_X4Y6_E2BEG[7] ,
    \Tile_X4Y6_E2BEG[6] ,
    \Tile_X4Y6_E2BEG[5] ,
    \Tile_X4Y6_E2BEG[4] ,
    \Tile_X4Y6_E2BEG[3] ,
    \Tile_X4Y6_E2BEG[2] ,
    \Tile_X4Y6_E2BEG[1] ,
    \Tile_X4Y6_E2BEG[0] }),
    .E2BEGb({\Tile_X4Y6_E2BEGb[7] ,
    \Tile_X4Y6_E2BEGb[6] ,
    \Tile_X4Y6_E2BEGb[5] ,
    \Tile_X4Y6_E2BEGb[4] ,
    \Tile_X4Y6_E2BEGb[3] ,
    \Tile_X4Y6_E2BEGb[2] ,
    \Tile_X4Y6_E2BEGb[1] ,
    \Tile_X4Y6_E2BEGb[0] }),
    .E2END({\Tile_X3Y6_E2BEGb[7] ,
    \Tile_X3Y6_E2BEGb[6] ,
    \Tile_X3Y6_E2BEGb[5] ,
    \Tile_X3Y6_E2BEGb[4] ,
    \Tile_X3Y6_E2BEGb[3] ,
    \Tile_X3Y6_E2BEGb[2] ,
    \Tile_X3Y6_E2BEGb[1] ,
    \Tile_X3Y6_E2BEGb[0] }),
    .E2MID({\Tile_X3Y6_E2BEG[7] ,
    \Tile_X3Y6_E2BEG[6] ,
    \Tile_X3Y6_E2BEG[5] ,
    \Tile_X3Y6_E2BEG[4] ,
    \Tile_X3Y6_E2BEG[3] ,
    \Tile_X3Y6_E2BEG[2] ,
    \Tile_X3Y6_E2BEG[1] ,
    \Tile_X3Y6_E2BEG[0] }),
    .E6BEG({\Tile_X4Y6_E6BEG[11] ,
    \Tile_X4Y6_E6BEG[10] ,
    \Tile_X4Y6_E6BEG[9] ,
    \Tile_X4Y6_E6BEG[8] ,
    \Tile_X4Y6_E6BEG[7] ,
    \Tile_X4Y6_E6BEG[6] ,
    \Tile_X4Y6_E6BEG[5] ,
    \Tile_X4Y6_E6BEG[4] ,
    \Tile_X4Y6_E6BEG[3] ,
    \Tile_X4Y6_E6BEG[2] ,
    \Tile_X4Y6_E6BEG[1] ,
    \Tile_X4Y6_E6BEG[0] }),
    .E6END({\Tile_X3Y6_E6BEG[11] ,
    \Tile_X3Y6_E6BEG[10] ,
    \Tile_X3Y6_E6BEG[9] ,
    \Tile_X3Y6_E6BEG[8] ,
    \Tile_X3Y6_E6BEG[7] ,
    \Tile_X3Y6_E6BEG[6] ,
    \Tile_X3Y6_E6BEG[5] ,
    \Tile_X3Y6_E6BEG[4] ,
    \Tile_X3Y6_E6BEG[3] ,
    \Tile_X3Y6_E6BEG[2] ,
    \Tile_X3Y6_E6BEG[1] ,
    \Tile_X3Y6_E6BEG[0] }),
    .EE4BEG({\Tile_X4Y6_EE4BEG[15] ,
    \Tile_X4Y6_EE4BEG[14] ,
    \Tile_X4Y6_EE4BEG[13] ,
    \Tile_X4Y6_EE4BEG[12] ,
    \Tile_X4Y6_EE4BEG[11] ,
    \Tile_X4Y6_EE4BEG[10] ,
    \Tile_X4Y6_EE4BEG[9] ,
    \Tile_X4Y6_EE4BEG[8] ,
    \Tile_X4Y6_EE4BEG[7] ,
    \Tile_X4Y6_EE4BEG[6] ,
    \Tile_X4Y6_EE4BEG[5] ,
    \Tile_X4Y6_EE4BEG[4] ,
    \Tile_X4Y6_EE4BEG[3] ,
    \Tile_X4Y6_EE4BEG[2] ,
    \Tile_X4Y6_EE4BEG[1] ,
    \Tile_X4Y6_EE4BEG[0] }),
    .EE4END({\Tile_X3Y6_EE4BEG[15] ,
    \Tile_X3Y6_EE4BEG[14] ,
    \Tile_X3Y6_EE4BEG[13] ,
    \Tile_X3Y6_EE4BEG[12] ,
    \Tile_X3Y6_EE4BEG[11] ,
    \Tile_X3Y6_EE4BEG[10] ,
    \Tile_X3Y6_EE4BEG[9] ,
    \Tile_X3Y6_EE4BEG[8] ,
    \Tile_X3Y6_EE4BEG[7] ,
    \Tile_X3Y6_EE4BEG[6] ,
    \Tile_X3Y6_EE4BEG[5] ,
    \Tile_X3Y6_EE4BEG[4] ,
    \Tile_X3Y6_EE4BEG[3] ,
    \Tile_X3Y6_EE4BEG[2] ,
    \Tile_X3Y6_EE4BEG[1] ,
    \Tile_X3Y6_EE4BEG[0] }),
    .FrameData({\Tile_X3Y6_FrameData_O[31] ,
    \Tile_X3Y6_FrameData_O[30] ,
    \Tile_X3Y6_FrameData_O[29] ,
    \Tile_X3Y6_FrameData_O[28] ,
    \Tile_X3Y6_FrameData_O[27] ,
    \Tile_X3Y6_FrameData_O[26] ,
    \Tile_X3Y6_FrameData_O[25] ,
    \Tile_X3Y6_FrameData_O[24] ,
    \Tile_X3Y6_FrameData_O[23] ,
    \Tile_X3Y6_FrameData_O[22] ,
    \Tile_X3Y6_FrameData_O[21] ,
    \Tile_X3Y6_FrameData_O[20] ,
    \Tile_X3Y6_FrameData_O[19] ,
    \Tile_X3Y6_FrameData_O[18] ,
    \Tile_X3Y6_FrameData_O[17] ,
    \Tile_X3Y6_FrameData_O[16] ,
    \Tile_X3Y6_FrameData_O[15] ,
    \Tile_X3Y6_FrameData_O[14] ,
    \Tile_X3Y6_FrameData_O[13] ,
    \Tile_X3Y6_FrameData_O[12] ,
    \Tile_X3Y6_FrameData_O[11] ,
    \Tile_X3Y6_FrameData_O[10] ,
    \Tile_X3Y6_FrameData_O[9] ,
    \Tile_X3Y6_FrameData_O[8] ,
    \Tile_X3Y6_FrameData_O[7] ,
    \Tile_X3Y6_FrameData_O[6] ,
    \Tile_X3Y6_FrameData_O[5] ,
    \Tile_X3Y6_FrameData_O[4] ,
    \Tile_X3Y6_FrameData_O[3] ,
    \Tile_X3Y6_FrameData_O[2] ,
    \Tile_X3Y6_FrameData_O[1] ,
    \Tile_X3Y6_FrameData_O[0] }),
    .FrameData_O({\Tile_X4Y6_FrameData_O[31] ,
    \Tile_X4Y6_FrameData_O[30] ,
    \Tile_X4Y6_FrameData_O[29] ,
    \Tile_X4Y6_FrameData_O[28] ,
    \Tile_X4Y6_FrameData_O[27] ,
    \Tile_X4Y6_FrameData_O[26] ,
    \Tile_X4Y6_FrameData_O[25] ,
    \Tile_X4Y6_FrameData_O[24] ,
    \Tile_X4Y6_FrameData_O[23] ,
    \Tile_X4Y6_FrameData_O[22] ,
    \Tile_X4Y6_FrameData_O[21] ,
    \Tile_X4Y6_FrameData_O[20] ,
    \Tile_X4Y6_FrameData_O[19] ,
    \Tile_X4Y6_FrameData_O[18] ,
    \Tile_X4Y6_FrameData_O[17] ,
    \Tile_X4Y6_FrameData_O[16] ,
    \Tile_X4Y6_FrameData_O[15] ,
    \Tile_X4Y6_FrameData_O[14] ,
    \Tile_X4Y6_FrameData_O[13] ,
    \Tile_X4Y6_FrameData_O[12] ,
    \Tile_X4Y6_FrameData_O[11] ,
    \Tile_X4Y6_FrameData_O[10] ,
    \Tile_X4Y6_FrameData_O[9] ,
    \Tile_X4Y6_FrameData_O[8] ,
    \Tile_X4Y6_FrameData_O[7] ,
    \Tile_X4Y6_FrameData_O[6] ,
    \Tile_X4Y6_FrameData_O[5] ,
    \Tile_X4Y6_FrameData_O[4] ,
    \Tile_X4Y6_FrameData_O[3] ,
    \Tile_X4Y6_FrameData_O[2] ,
    \Tile_X4Y6_FrameData_O[1] ,
    \Tile_X4Y6_FrameData_O[0] }),
    .FrameStrobe({\Tile_X4Y7_FrameStrobe_O[19] ,
    \Tile_X4Y7_FrameStrobe_O[18] ,
    \Tile_X4Y7_FrameStrobe_O[17] ,
    \Tile_X4Y7_FrameStrobe_O[16] ,
    \Tile_X4Y7_FrameStrobe_O[15] ,
    \Tile_X4Y7_FrameStrobe_O[14] ,
    \Tile_X4Y7_FrameStrobe_O[13] ,
    \Tile_X4Y7_FrameStrobe_O[12] ,
    \Tile_X4Y7_FrameStrobe_O[11] ,
    \Tile_X4Y7_FrameStrobe_O[10] ,
    \Tile_X4Y7_FrameStrobe_O[9] ,
    \Tile_X4Y7_FrameStrobe_O[8] ,
    \Tile_X4Y7_FrameStrobe_O[7] ,
    \Tile_X4Y7_FrameStrobe_O[6] ,
    \Tile_X4Y7_FrameStrobe_O[5] ,
    \Tile_X4Y7_FrameStrobe_O[4] ,
    \Tile_X4Y7_FrameStrobe_O[3] ,
    \Tile_X4Y7_FrameStrobe_O[2] ,
    \Tile_X4Y7_FrameStrobe_O[1] ,
    \Tile_X4Y7_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X4Y6_FrameStrobe_O[19] ,
    \Tile_X4Y6_FrameStrobe_O[18] ,
    \Tile_X4Y6_FrameStrobe_O[17] ,
    \Tile_X4Y6_FrameStrobe_O[16] ,
    \Tile_X4Y6_FrameStrobe_O[15] ,
    \Tile_X4Y6_FrameStrobe_O[14] ,
    \Tile_X4Y6_FrameStrobe_O[13] ,
    \Tile_X4Y6_FrameStrobe_O[12] ,
    \Tile_X4Y6_FrameStrobe_O[11] ,
    \Tile_X4Y6_FrameStrobe_O[10] ,
    \Tile_X4Y6_FrameStrobe_O[9] ,
    \Tile_X4Y6_FrameStrobe_O[8] ,
    \Tile_X4Y6_FrameStrobe_O[7] ,
    \Tile_X4Y6_FrameStrobe_O[6] ,
    \Tile_X4Y6_FrameStrobe_O[5] ,
    \Tile_X4Y6_FrameStrobe_O[4] ,
    \Tile_X4Y6_FrameStrobe_O[3] ,
    \Tile_X4Y6_FrameStrobe_O[2] ,
    \Tile_X4Y6_FrameStrobe_O[1] ,
    \Tile_X4Y6_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X4Y6_N1BEG[3] ,
    \Tile_X4Y6_N1BEG[2] ,
    \Tile_X4Y6_N1BEG[1] ,
    \Tile_X4Y6_N1BEG[0] }),
    .N1END({\Tile_X4Y7_N1BEG[3] ,
    \Tile_X4Y7_N1BEG[2] ,
    \Tile_X4Y7_N1BEG[1] ,
    \Tile_X4Y7_N1BEG[0] }),
    .N2BEG({\Tile_X4Y6_N2BEG[7] ,
    \Tile_X4Y6_N2BEG[6] ,
    \Tile_X4Y6_N2BEG[5] ,
    \Tile_X4Y6_N2BEG[4] ,
    \Tile_X4Y6_N2BEG[3] ,
    \Tile_X4Y6_N2BEG[2] ,
    \Tile_X4Y6_N2BEG[1] ,
    \Tile_X4Y6_N2BEG[0] }),
    .N2BEGb({\Tile_X4Y6_N2BEGb[7] ,
    \Tile_X4Y6_N2BEGb[6] ,
    \Tile_X4Y6_N2BEGb[5] ,
    \Tile_X4Y6_N2BEGb[4] ,
    \Tile_X4Y6_N2BEGb[3] ,
    \Tile_X4Y6_N2BEGb[2] ,
    \Tile_X4Y6_N2BEGb[1] ,
    \Tile_X4Y6_N2BEGb[0] }),
    .N2END({\Tile_X4Y7_N2BEGb[7] ,
    \Tile_X4Y7_N2BEGb[6] ,
    \Tile_X4Y7_N2BEGb[5] ,
    \Tile_X4Y7_N2BEGb[4] ,
    \Tile_X4Y7_N2BEGb[3] ,
    \Tile_X4Y7_N2BEGb[2] ,
    \Tile_X4Y7_N2BEGb[1] ,
    \Tile_X4Y7_N2BEGb[0] }),
    .N2MID({\Tile_X4Y7_N2BEG[7] ,
    \Tile_X4Y7_N2BEG[6] ,
    \Tile_X4Y7_N2BEG[5] ,
    \Tile_X4Y7_N2BEG[4] ,
    \Tile_X4Y7_N2BEG[3] ,
    \Tile_X4Y7_N2BEG[2] ,
    \Tile_X4Y7_N2BEG[1] ,
    \Tile_X4Y7_N2BEG[0] }),
    .N4BEG({\Tile_X4Y6_N4BEG[15] ,
    \Tile_X4Y6_N4BEG[14] ,
    \Tile_X4Y6_N4BEG[13] ,
    \Tile_X4Y6_N4BEG[12] ,
    \Tile_X4Y6_N4BEG[11] ,
    \Tile_X4Y6_N4BEG[10] ,
    \Tile_X4Y6_N4BEG[9] ,
    \Tile_X4Y6_N4BEG[8] ,
    \Tile_X4Y6_N4BEG[7] ,
    \Tile_X4Y6_N4BEG[6] ,
    \Tile_X4Y6_N4BEG[5] ,
    \Tile_X4Y6_N4BEG[4] ,
    \Tile_X4Y6_N4BEG[3] ,
    \Tile_X4Y6_N4BEG[2] ,
    \Tile_X4Y6_N4BEG[1] ,
    \Tile_X4Y6_N4BEG[0] }),
    .N4END({\Tile_X4Y7_N4BEG[15] ,
    \Tile_X4Y7_N4BEG[14] ,
    \Tile_X4Y7_N4BEG[13] ,
    \Tile_X4Y7_N4BEG[12] ,
    \Tile_X4Y7_N4BEG[11] ,
    \Tile_X4Y7_N4BEG[10] ,
    \Tile_X4Y7_N4BEG[9] ,
    \Tile_X4Y7_N4BEG[8] ,
    \Tile_X4Y7_N4BEG[7] ,
    \Tile_X4Y7_N4BEG[6] ,
    \Tile_X4Y7_N4BEG[5] ,
    \Tile_X4Y7_N4BEG[4] ,
    \Tile_X4Y7_N4BEG[3] ,
    \Tile_X4Y7_N4BEG[2] ,
    \Tile_X4Y7_N4BEG[1] ,
    \Tile_X4Y7_N4BEG[0] }),
    .NN4BEG({\Tile_X4Y6_NN4BEG[15] ,
    \Tile_X4Y6_NN4BEG[14] ,
    \Tile_X4Y6_NN4BEG[13] ,
    \Tile_X4Y6_NN4BEG[12] ,
    \Tile_X4Y6_NN4BEG[11] ,
    \Tile_X4Y6_NN4BEG[10] ,
    \Tile_X4Y6_NN4BEG[9] ,
    \Tile_X4Y6_NN4BEG[8] ,
    \Tile_X4Y6_NN4BEG[7] ,
    \Tile_X4Y6_NN4BEG[6] ,
    \Tile_X4Y6_NN4BEG[5] ,
    \Tile_X4Y6_NN4BEG[4] ,
    \Tile_X4Y6_NN4BEG[3] ,
    \Tile_X4Y6_NN4BEG[2] ,
    \Tile_X4Y6_NN4BEG[1] ,
    \Tile_X4Y6_NN4BEG[0] }),
    .NN4END({\Tile_X4Y7_NN4BEG[15] ,
    \Tile_X4Y7_NN4BEG[14] ,
    \Tile_X4Y7_NN4BEG[13] ,
    \Tile_X4Y7_NN4BEG[12] ,
    \Tile_X4Y7_NN4BEG[11] ,
    \Tile_X4Y7_NN4BEG[10] ,
    \Tile_X4Y7_NN4BEG[9] ,
    \Tile_X4Y7_NN4BEG[8] ,
    \Tile_X4Y7_NN4BEG[7] ,
    \Tile_X4Y7_NN4BEG[6] ,
    \Tile_X4Y7_NN4BEG[5] ,
    \Tile_X4Y7_NN4BEG[4] ,
    \Tile_X4Y7_NN4BEG[3] ,
    \Tile_X4Y7_NN4BEG[2] ,
    \Tile_X4Y7_NN4BEG[1] ,
    \Tile_X4Y7_NN4BEG[0] }),
    .S1BEG({\Tile_X4Y6_S1BEG[3] ,
    \Tile_X4Y6_S1BEG[2] ,
    \Tile_X4Y6_S1BEG[1] ,
    \Tile_X4Y6_S1BEG[0] }),
    .S1END({\Tile_X4Y5_S1BEG[3] ,
    \Tile_X4Y5_S1BEG[2] ,
    \Tile_X4Y5_S1BEG[1] ,
    \Tile_X4Y5_S1BEG[0] }),
    .S2BEG({\Tile_X4Y6_S2BEG[7] ,
    \Tile_X4Y6_S2BEG[6] ,
    \Tile_X4Y6_S2BEG[5] ,
    \Tile_X4Y6_S2BEG[4] ,
    \Tile_X4Y6_S2BEG[3] ,
    \Tile_X4Y6_S2BEG[2] ,
    \Tile_X4Y6_S2BEG[1] ,
    \Tile_X4Y6_S2BEG[0] }),
    .S2BEGb({\Tile_X4Y6_S2BEGb[7] ,
    \Tile_X4Y6_S2BEGb[6] ,
    \Tile_X4Y6_S2BEGb[5] ,
    \Tile_X4Y6_S2BEGb[4] ,
    \Tile_X4Y6_S2BEGb[3] ,
    \Tile_X4Y6_S2BEGb[2] ,
    \Tile_X4Y6_S2BEGb[1] ,
    \Tile_X4Y6_S2BEGb[0] }),
    .S2END({\Tile_X4Y5_S2BEGb[7] ,
    \Tile_X4Y5_S2BEGb[6] ,
    \Tile_X4Y5_S2BEGb[5] ,
    \Tile_X4Y5_S2BEGb[4] ,
    \Tile_X4Y5_S2BEGb[3] ,
    \Tile_X4Y5_S2BEGb[2] ,
    \Tile_X4Y5_S2BEGb[1] ,
    \Tile_X4Y5_S2BEGb[0] }),
    .S2MID({\Tile_X4Y5_S2BEG[7] ,
    \Tile_X4Y5_S2BEG[6] ,
    \Tile_X4Y5_S2BEG[5] ,
    \Tile_X4Y5_S2BEG[4] ,
    \Tile_X4Y5_S2BEG[3] ,
    \Tile_X4Y5_S2BEG[2] ,
    \Tile_X4Y5_S2BEG[1] ,
    \Tile_X4Y5_S2BEG[0] }),
    .S4BEG({\Tile_X4Y6_S4BEG[15] ,
    \Tile_X4Y6_S4BEG[14] ,
    \Tile_X4Y6_S4BEG[13] ,
    \Tile_X4Y6_S4BEG[12] ,
    \Tile_X4Y6_S4BEG[11] ,
    \Tile_X4Y6_S4BEG[10] ,
    \Tile_X4Y6_S4BEG[9] ,
    \Tile_X4Y6_S4BEG[8] ,
    \Tile_X4Y6_S4BEG[7] ,
    \Tile_X4Y6_S4BEG[6] ,
    \Tile_X4Y6_S4BEG[5] ,
    \Tile_X4Y6_S4BEG[4] ,
    \Tile_X4Y6_S4BEG[3] ,
    \Tile_X4Y6_S4BEG[2] ,
    \Tile_X4Y6_S4BEG[1] ,
    \Tile_X4Y6_S4BEG[0] }),
    .S4END({\Tile_X4Y5_S4BEG[15] ,
    \Tile_X4Y5_S4BEG[14] ,
    \Tile_X4Y5_S4BEG[13] ,
    \Tile_X4Y5_S4BEG[12] ,
    \Tile_X4Y5_S4BEG[11] ,
    \Tile_X4Y5_S4BEG[10] ,
    \Tile_X4Y5_S4BEG[9] ,
    \Tile_X4Y5_S4BEG[8] ,
    \Tile_X4Y5_S4BEG[7] ,
    \Tile_X4Y5_S4BEG[6] ,
    \Tile_X4Y5_S4BEG[5] ,
    \Tile_X4Y5_S4BEG[4] ,
    \Tile_X4Y5_S4BEG[3] ,
    \Tile_X4Y5_S4BEG[2] ,
    \Tile_X4Y5_S4BEG[1] ,
    \Tile_X4Y5_S4BEG[0] }),
    .SS4BEG({\Tile_X4Y6_SS4BEG[15] ,
    \Tile_X4Y6_SS4BEG[14] ,
    \Tile_X4Y6_SS4BEG[13] ,
    \Tile_X4Y6_SS4BEG[12] ,
    \Tile_X4Y6_SS4BEG[11] ,
    \Tile_X4Y6_SS4BEG[10] ,
    \Tile_X4Y6_SS4BEG[9] ,
    \Tile_X4Y6_SS4BEG[8] ,
    \Tile_X4Y6_SS4BEG[7] ,
    \Tile_X4Y6_SS4BEG[6] ,
    \Tile_X4Y6_SS4BEG[5] ,
    \Tile_X4Y6_SS4BEG[4] ,
    \Tile_X4Y6_SS4BEG[3] ,
    \Tile_X4Y6_SS4BEG[2] ,
    \Tile_X4Y6_SS4BEG[1] ,
    \Tile_X4Y6_SS4BEG[0] }),
    .SS4END({\Tile_X4Y5_SS4BEG[15] ,
    \Tile_X4Y5_SS4BEG[14] ,
    \Tile_X4Y5_SS4BEG[13] ,
    \Tile_X4Y5_SS4BEG[12] ,
    \Tile_X4Y5_SS4BEG[11] ,
    \Tile_X4Y5_SS4BEG[10] ,
    \Tile_X4Y5_SS4BEG[9] ,
    \Tile_X4Y5_SS4BEG[8] ,
    \Tile_X4Y5_SS4BEG[7] ,
    \Tile_X4Y5_SS4BEG[6] ,
    \Tile_X4Y5_SS4BEG[5] ,
    \Tile_X4Y5_SS4BEG[4] ,
    \Tile_X4Y5_SS4BEG[3] ,
    \Tile_X4Y5_SS4BEG[2] ,
    \Tile_X4Y5_SS4BEG[1] ,
    \Tile_X4Y5_SS4BEG[0] }),
    .W1BEG({\Tile_X4Y6_W1BEG[3] ,
    \Tile_X4Y6_W1BEG[2] ,
    \Tile_X4Y6_W1BEG[1] ,
    \Tile_X4Y6_W1BEG[0] }),
    .W1END({\Tile_X5Y6_W1BEG[3] ,
    \Tile_X5Y6_W1BEG[2] ,
    \Tile_X5Y6_W1BEG[1] ,
    \Tile_X5Y6_W1BEG[0] }),
    .W2BEG({\Tile_X4Y6_W2BEG[7] ,
    \Tile_X4Y6_W2BEG[6] ,
    \Tile_X4Y6_W2BEG[5] ,
    \Tile_X4Y6_W2BEG[4] ,
    \Tile_X4Y6_W2BEG[3] ,
    \Tile_X4Y6_W2BEG[2] ,
    \Tile_X4Y6_W2BEG[1] ,
    \Tile_X4Y6_W2BEG[0] }),
    .W2BEGb({\Tile_X4Y6_W2BEGb[7] ,
    \Tile_X4Y6_W2BEGb[6] ,
    \Tile_X4Y6_W2BEGb[5] ,
    \Tile_X4Y6_W2BEGb[4] ,
    \Tile_X4Y6_W2BEGb[3] ,
    \Tile_X4Y6_W2BEGb[2] ,
    \Tile_X4Y6_W2BEGb[1] ,
    \Tile_X4Y6_W2BEGb[0] }),
    .W2END({\Tile_X5Y6_W2BEGb[7] ,
    \Tile_X5Y6_W2BEGb[6] ,
    \Tile_X5Y6_W2BEGb[5] ,
    \Tile_X5Y6_W2BEGb[4] ,
    \Tile_X5Y6_W2BEGb[3] ,
    \Tile_X5Y6_W2BEGb[2] ,
    \Tile_X5Y6_W2BEGb[1] ,
    \Tile_X5Y6_W2BEGb[0] }),
    .W2MID({\Tile_X5Y6_W2BEG[7] ,
    \Tile_X5Y6_W2BEG[6] ,
    \Tile_X5Y6_W2BEG[5] ,
    \Tile_X5Y6_W2BEG[4] ,
    \Tile_X5Y6_W2BEG[3] ,
    \Tile_X5Y6_W2BEG[2] ,
    \Tile_X5Y6_W2BEG[1] ,
    \Tile_X5Y6_W2BEG[0] }),
    .W6BEG({\Tile_X4Y6_W6BEG[11] ,
    \Tile_X4Y6_W6BEG[10] ,
    \Tile_X4Y6_W6BEG[9] ,
    \Tile_X4Y6_W6BEG[8] ,
    \Tile_X4Y6_W6BEG[7] ,
    \Tile_X4Y6_W6BEG[6] ,
    \Tile_X4Y6_W6BEG[5] ,
    \Tile_X4Y6_W6BEG[4] ,
    \Tile_X4Y6_W6BEG[3] ,
    \Tile_X4Y6_W6BEG[2] ,
    \Tile_X4Y6_W6BEG[1] ,
    \Tile_X4Y6_W6BEG[0] }),
    .W6END({\Tile_X5Y6_W6BEG[11] ,
    \Tile_X5Y6_W6BEG[10] ,
    \Tile_X5Y6_W6BEG[9] ,
    \Tile_X5Y6_W6BEG[8] ,
    \Tile_X5Y6_W6BEG[7] ,
    \Tile_X5Y6_W6BEG[6] ,
    \Tile_X5Y6_W6BEG[5] ,
    \Tile_X5Y6_W6BEG[4] ,
    \Tile_X5Y6_W6BEG[3] ,
    \Tile_X5Y6_W6BEG[2] ,
    \Tile_X5Y6_W6BEG[1] ,
    \Tile_X5Y6_W6BEG[0] }),
    .WW4BEG({\Tile_X4Y6_WW4BEG[15] ,
    \Tile_X4Y6_WW4BEG[14] ,
    \Tile_X4Y6_WW4BEG[13] ,
    \Tile_X4Y6_WW4BEG[12] ,
    \Tile_X4Y6_WW4BEG[11] ,
    \Tile_X4Y6_WW4BEG[10] ,
    \Tile_X4Y6_WW4BEG[9] ,
    \Tile_X4Y6_WW4BEG[8] ,
    \Tile_X4Y6_WW4BEG[7] ,
    \Tile_X4Y6_WW4BEG[6] ,
    \Tile_X4Y6_WW4BEG[5] ,
    \Tile_X4Y6_WW4BEG[4] ,
    \Tile_X4Y6_WW4BEG[3] ,
    \Tile_X4Y6_WW4BEG[2] ,
    \Tile_X4Y6_WW4BEG[1] ,
    \Tile_X4Y6_WW4BEG[0] }),
    .WW4END({\Tile_X5Y6_WW4BEG[15] ,
    \Tile_X5Y6_WW4BEG[14] ,
    \Tile_X5Y6_WW4BEG[13] ,
    \Tile_X5Y6_WW4BEG[12] ,
    \Tile_X5Y6_WW4BEG[11] ,
    \Tile_X5Y6_WW4BEG[10] ,
    \Tile_X5Y6_WW4BEG[9] ,
    \Tile_X5Y6_WW4BEG[8] ,
    \Tile_X5Y6_WW4BEG[7] ,
    \Tile_X5Y6_WW4BEG[6] ,
    \Tile_X5Y6_WW4BEG[5] ,
    \Tile_X5Y6_WW4BEG[4] ,
    \Tile_X5Y6_WW4BEG[3] ,
    \Tile_X5Y6_WW4BEG[2] ,
    \Tile_X5Y6_WW4BEG[1] ,
    \Tile_X5Y6_WW4BEG[0] }));
 LUT4AB Tile_X4Y7_LUT4AB (.Ci(Tile_X4Y8_Co),
    .Co(Tile_X4Y7_Co),
    .UserCLK(Tile_X4Y8_UserCLKo),
    .UserCLKo(Tile_X4Y7_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X4Y7_E1BEG[3] ,
    \Tile_X4Y7_E1BEG[2] ,
    \Tile_X4Y7_E1BEG[1] ,
    \Tile_X4Y7_E1BEG[0] }),
    .E1END({\Tile_X3Y7_E1BEG[3] ,
    \Tile_X3Y7_E1BEG[2] ,
    \Tile_X3Y7_E1BEG[1] ,
    \Tile_X3Y7_E1BEG[0] }),
    .E2BEG({\Tile_X4Y7_E2BEG[7] ,
    \Tile_X4Y7_E2BEG[6] ,
    \Tile_X4Y7_E2BEG[5] ,
    \Tile_X4Y7_E2BEG[4] ,
    \Tile_X4Y7_E2BEG[3] ,
    \Tile_X4Y7_E2BEG[2] ,
    \Tile_X4Y7_E2BEG[1] ,
    \Tile_X4Y7_E2BEG[0] }),
    .E2BEGb({\Tile_X4Y7_E2BEGb[7] ,
    \Tile_X4Y7_E2BEGb[6] ,
    \Tile_X4Y7_E2BEGb[5] ,
    \Tile_X4Y7_E2BEGb[4] ,
    \Tile_X4Y7_E2BEGb[3] ,
    \Tile_X4Y7_E2BEGb[2] ,
    \Tile_X4Y7_E2BEGb[1] ,
    \Tile_X4Y7_E2BEGb[0] }),
    .E2END({\Tile_X3Y7_E2BEGb[7] ,
    \Tile_X3Y7_E2BEGb[6] ,
    \Tile_X3Y7_E2BEGb[5] ,
    \Tile_X3Y7_E2BEGb[4] ,
    \Tile_X3Y7_E2BEGb[3] ,
    \Tile_X3Y7_E2BEGb[2] ,
    \Tile_X3Y7_E2BEGb[1] ,
    \Tile_X3Y7_E2BEGb[0] }),
    .E2MID({\Tile_X3Y7_E2BEG[7] ,
    \Tile_X3Y7_E2BEG[6] ,
    \Tile_X3Y7_E2BEG[5] ,
    \Tile_X3Y7_E2BEG[4] ,
    \Tile_X3Y7_E2BEG[3] ,
    \Tile_X3Y7_E2BEG[2] ,
    \Tile_X3Y7_E2BEG[1] ,
    \Tile_X3Y7_E2BEG[0] }),
    .E6BEG({\Tile_X4Y7_E6BEG[11] ,
    \Tile_X4Y7_E6BEG[10] ,
    \Tile_X4Y7_E6BEG[9] ,
    \Tile_X4Y7_E6BEG[8] ,
    \Tile_X4Y7_E6BEG[7] ,
    \Tile_X4Y7_E6BEG[6] ,
    \Tile_X4Y7_E6BEG[5] ,
    \Tile_X4Y7_E6BEG[4] ,
    \Tile_X4Y7_E6BEG[3] ,
    \Tile_X4Y7_E6BEG[2] ,
    \Tile_X4Y7_E6BEG[1] ,
    \Tile_X4Y7_E6BEG[0] }),
    .E6END({\Tile_X3Y7_E6BEG[11] ,
    \Tile_X3Y7_E6BEG[10] ,
    \Tile_X3Y7_E6BEG[9] ,
    \Tile_X3Y7_E6BEG[8] ,
    \Tile_X3Y7_E6BEG[7] ,
    \Tile_X3Y7_E6BEG[6] ,
    \Tile_X3Y7_E6BEG[5] ,
    \Tile_X3Y7_E6BEG[4] ,
    \Tile_X3Y7_E6BEG[3] ,
    \Tile_X3Y7_E6BEG[2] ,
    \Tile_X3Y7_E6BEG[1] ,
    \Tile_X3Y7_E6BEG[0] }),
    .EE4BEG({\Tile_X4Y7_EE4BEG[15] ,
    \Tile_X4Y7_EE4BEG[14] ,
    \Tile_X4Y7_EE4BEG[13] ,
    \Tile_X4Y7_EE4BEG[12] ,
    \Tile_X4Y7_EE4BEG[11] ,
    \Tile_X4Y7_EE4BEG[10] ,
    \Tile_X4Y7_EE4BEG[9] ,
    \Tile_X4Y7_EE4BEG[8] ,
    \Tile_X4Y7_EE4BEG[7] ,
    \Tile_X4Y7_EE4BEG[6] ,
    \Tile_X4Y7_EE4BEG[5] ,
    \Tile_X4Y7_EE4BEG[4] ,
    \Tile_X4Y7_EE4BEG[3] ,
    \Tile_X4Y7_EE4BEG[2] ,
    \Tile_X4Y7_EE4BEG[1] ,
    \Tile_X4Y7_EE4BEG[0] }),
    .EE4END({\Tile_X3Y7_EE4BEG[15] ,
    \Tile_X3Y7_EE4BEG[14] ,
    \Tile_X3Y7_EE4BEG[13] ,
    \Tile_X3Y7_EE4BEG[12] ,
    \Tile_X3Y7_EE4BEG[11] ,
    \Tile_X3Y7_EE4BEG[10] ,
    \Tile_X3Y7_EE4BEG[9] ,
    \Tile_X3Y7_EE4BEG[8] ,
    \Tile_X3Y7_EE4BEG[7] ,
    \Tile_X3Y7_EE4BEG[6] ,
    \Tile_X3Y7_EE4BEG[5] ,
    \Tile_X3Y7_EE4BEG[4] ,
    \Tile_X3Y7_EE4BEG[3] ,
    \Tile_X3Y7_EE4BEG[2] ,
    \Tile_X3Y7_EE4BEG[1] ,
    \Tile_X3Y7_EE4BEG[0] }),
    .FrameData({\Tile_X3Y7_FrameData_O[31] ,
    \Tile_X3Y7_FrameData_O[30] ,
    \Tile_X3Y7_FrameData_O[29] ,
    \Tile_X3Y7_FrameData_O[28] ,
    \Tile_X3Y7_FrameData_O[27] ,
    \Tile_X3Y7_FrameData_O[26] ,
    \Tile_X3Y7_FrameData_O[25] ,
    \Tile_X3Y7_FrameData_O[24] ,
    \Tile_X3Y7_FrameData_O[23] ,
    \Tile_X3Y7_FrameData_O[22] ,
    \Tile_X3Y7_FrameData_O[21] ,
    \Tile_X3Y7_FrameData_O[20] ,
    \Tile_X3Y7_FrameData_O[19] ,
    \Tile_X3Y7_FrameData_O[18] ,
    \Tile_X3Y7_FrameData_O[17] ,
    \Tile_X3Y7_FrameData_O[16] ,
    \Tile_X3Y7_FrameData_O[15] ,
    \Tile_X3Y7_FrameData_O[14] ,
    \Tile_X3Y7_FrameData_O[13] ,
    \Tile_X3Y7_FrameData_O[12] ,
    \Tile_X3Y7_FrameData_O[11] ,
    \Tile_X3Y7_FrameData_O[10] ,
    \Tile_X3Y7_FrameData_O[9] ,
    \Tile_X3Y7_FrameData_O[8] ,
    \Tile_X3Y7_FrameData_O[7] ,
    \Tile_X3Y7_FrameData_O[6] ,
    \Tile_X3Y7_FrameData_O[5] ,
    \Tile_X3Y7_FrameData_O[4] ,
    \Tile_X3Y7_FrameData_O[3] ,
    \Tile_X3Y7_FrameData_O[2] ,
    \Tile_X3Y7_FrameData_O[1] ,
    \Tile_X3Y7_FrameData_O[0] }),
    .FrameData_O({\Tile_X4Y7_FrameData_O[31] ,
    \Tile_X4Y7_FrameData_O[30] ,
    \Tile_X4Y7_FrameData_O[29] ,
    \Tile_X4Y7_FrameData_O[28] ,
    \Tile_X4Y7_FrameData_O[27] ,
    \Tile_X4Y7_FrameData_O[26] ,
    \Tile_X4Y7_FrameData_O[25] ,
    \Tile_X4Y7_FrameData_O[24] ,
    \Tile_X4Y7_FrameData_O[23] ,
    \Tile_X4Y7_FrameData_O[22] ,
    \Tile_X4Y7_FrameData_O[21] ,
    \Tile_X4Y7_FrameData_O[20] ,
    \Tile_X4Y7_FrameData_O[19] ,
    \Tile_X4Y7_FrameData_O[18] ,
    \Tile_X4Y7_FrameData_O[17] ,
    \Tile_X4Y7_FrameData_O[16] ,
    \Tile_X4Y7_FrameData_O[15] ,
    \Tile_X4Y7_FrameData_O[14] ,
    \Tile_X4Y7_FrameData_O[13] ,
    \Tile_X4Y7_FrameData_O[12] ,
    \Tile_X4Y7_FrameData_O[11] ,
    \Tile_X4Y7_FrameData_O[10] ,
    \Tile_X4Y7_FrameData_O[9] ,
    \Tile_X4Y7_FrameData_O[8] ,
    \Tile_X4Y7_FrameData_O[7] ,
    \Tile_X4Y7_FrameData_O[6] ,
    \Tile_X4Y7_FrameData_O[5] ,
    \Tile_X4Y7_FrameData_O[4] ,
    \Tile_X4Y7_FrameData_O[3] ,
    \Tile_X4Y7_FrameData_O[2] ,
    \Tile_X4Y7_FrameData_O[1] ,
    \Tile_X4Y7_FrameData_O[0] }),
    .FrameStrobe({\Tile_X4Y8_FrameStrobe_O[19] ,
    \Tile_X4Y8_FrameStrobe_O[18] ,
    \Tile_X4Y8_FrameStrobe_O[17] ,
    \Tile_X4Y8_FrameStrobe_O[16] ,
    \Tile_X4Y8_FrameStrobe_O[15] ,
    \Tile_X4Y8_FrameStrobe_O[14] ,
    \Tile_X4Y8_FrameStrobe_O[13] ,
    \Tile_X4Y8_FrameStrobe_O[12] ,
    \Tile_X4Y8_FrameStrobe_O[11] ,
    \Tile_X4Y8_FrameStrobe_O[10] ,
    \Tile_X4Y8_FrameStrobe_O[9] ,
    \Tile_X4Y8_FrameStrobe_O[8] ,
    \Tile_X4Y8_FrameStrobe_O[7] ,
    \Tile_X4Y8_FrameStrobe_O[6] ,
    \Tile_X4Y8_FrameStrobe_O[5] ,
    \Tile_X4Y8_FrameStrobe_O[4] ,
    \Tile_X4Y8_FrameStrobe_O[3] ,
    \Tile_X4Y8_FrameStrobe_O[2] ,
    \Tile_X4Y8_FrameStrobe_O[1] ,
    \Tile_X4Y8_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X4Y7_FrameStrobe_O[19] ,
    \Tile_X4Y7_FrameStrobe_O[18] ,
    \Tile_X4Y7_FrameStrobe_O[17] ,
    \Tile_X4Y7_FrameStrobe_O[16] ,
    \Tile_X4Y7_FrameStrobe_O[15] ,
    \Tile_X4Y7_FrameStrobe_O[14] ,
    \Tile_X4Y7_FrameStrobe_O[13] ,
    \Tile_X4Y7_FrameStrobe_O[12] ,
    \Tile_X4Y7_FrameStrobe_O[11] ,
    \Tile_X4Y7_FrameStrobe_O[10] ,
    \Tile_X4Y7_FrameStrobe_O[9] ,
    \Tile_X4Y7_FrameStrobe_O[8] ,
    \Tile_X4Y7_FrameStrobe_O[7] ,
    \Tile_X4Y7_FrameStrobe_O[6] ,
    \Tile_X4Y7_FrameStrobe_O[5] ,
    \Tile_X4Y7_FrameStrobe_O[4] ,
    \Tile_X4Y7_FrameStrobe_O[3] ,
    \Tile_X4Y7_FrameStrobe_O[2] ,
    \Tile_X4Y7_FrameStrobe_O[1] ,
    \Tile_X4Y7_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X4Y7_N1BEG[3] ,
    \Tile_X4Y7_N1BEG[2] ,
    \Tile_X4Y7_N1BEG[1] ,
    \Tile_X4Y7_N1BEG[0] }),
    .N1END({\Tile_X4Y8_N1BEG[3] ,
    \Tile_X4Y8_N1BEG[2] ,
    \Tile_X4Y8_N1BEG[1] ,
    \Tile_X4Y8_N1BEG[0] }),
    .N2BEG({\Tile_X4Y7_N2BEG[7] ,
    \Tile_X4Y7_N2BEG[6] ,
    \Tile_X4Y7_N2BEG[5] ,
    \Tile_X4Y7_N2BEG[4] ,
    \Tile_X4Y7_N2BEG[3] ,
    \Tile_X4Y7_N2BEG[2] ,
    \Tile_X4Y7_N2BEG[1] ,
    \Tile_X4Y7_N2BEG[0] }),
    .N2BEGb({\Tile_X4Y7_N2BEGb[7] ,
    \Tile_X4Y7_N2BEGb[6] ,
    \Tile_X4Y7_N2BEGb[5] ,
    \Tile_X4Y7_N2BEGb[4] ,
    \Tile_X4Y7_N2BEGb[3] ,
    \Tile_X4Y7_N2BEGb[2] ,
    \Tile_X4Y7_N2BEGb[1] ,
    \Tile_X4Y7_N2BEGb[0] }),
    .N2END({\Tile_X4Y8_N2BEGb[7] ,
    \Tile_X4Y8_N2BEGb[6] ,
    \Tile_X4Y8_N2BEGb[5] ,
    \Tile_X4Y8_N2BEGb[4] ,
    \Tile_X4Y8_N2BEGb[3] ,
    \Tile_X4Y8_N2BEGb[2] ,
    \Tile_X4Y8_N2BEGb[1] ,
    \Tile_X4Y8_N2BEGb[0] }),
    .N2MID({\Tile_X4Y8_N2BEG[7] ,
    \Tile_X4Y8_N2BEG[6] ,
    \Tile_X4Y8_N2BEG[5] ,
    \Tile_X4Y8_N2BEG[4] ,
    \Tile_X4Y8_N2BEG[3] ,
    \Tile_X4Y8_N2BEG[2] ,
    \Tile_X4Y8_N2BEG[1] ,
    \Tile_X4Y8_N2BEG[0] }),
    .N4BEG({\Tile_X4Y7_N4BEG[15] ,
    \Tile_X4Y7_N4BEG[14] ,
    \Tile_X4Y7_N4BEG[13] ,
    \Tile_X4Y7_N4BEG[12] ,
    \Tile_X4Y7_N4BEG[11] ,
    \Tile_X4Y7_N4BEG[10] ,
    \Tile_X4Y7_N4BEG[9] ,
    \Tile_X4Y7_N4BEG[8] ,
    \Tile_X4Y7_N4BEG[7] ,
    \Tile_X4Y7_N4BEG[6] ,
    \Tile_X4Y7_N4BEG[5] ,
    \Tile_X4Y7_N4BEG[4] ,
    \Tile_X4Y7_N4BEG[3] ,
    \Tile_X4Y7_N4BEG[2] ,
    \Tile_X4Y7_N4BEG[1] ,
    \Tile_X4Y7_N4BEG[0] }),
    .N4END({\Tile_X4Y8_N4BEG[15] ,
    \Tile_X4Y8_N4BEG[14] ,
    \Tile_X4Y8_N4BEG[13] ,
    \Tile_X4Y8_N4BEG[12] ,
    \Tile_X4Y8_N4BEG[11] ,
    \Tile_X4Y8_N4BEG[10] ,
    \Tile_X4Y8_N4BEG[9] ,
    \Tile_X4Y8_N4BEG[8] ,
    \Tile_X4Y8_N4BEG[7] ,
    \Tile_X4Y8_N4BEG[6] ,
    \Tile_X4Y8_N4BEG[5] ,
    \Tile_X4Y8_N4BEG[4] ,
    \Tile_X4Y8_N4BEG[3] ,
    \Tile_X4Y8_N4BEG[2] ,
    \Tile_X4Y8_N4BEG[1] ,
    \Tile_X4Y8_N4BEG[0] }),
    .NN4BEG({\Tile_X4Y7_NN4BEG[15] ,
    \Tile_X4Y7_NN4BEG[14] ,
    \Tile_X4Y7_NN4BEG[13] ,
    \Tile_X4Y7_NN4BEG[12] ,
    \Tile_X4Y7_NN4BEG[11] ,
    \Tile_X4Y7_NN4BEG[10] ,
    \Tile_X4Y7_NN4BEG[9] ,
    \Tile_X4Y7_NN4BEG[8] ,
    \Tile_X4Y7_NN4BEG[7] ,
    \Tile_X4Y7_NN4BEG[6] ,
    \Tile_X4Y7_NN4BEG[5] ,
    \Tile_X4Y7_NN4BEG[4] ,
    \Tile_X4Y7_NN4BEG[3] ,
    \Tile_X4Y7_NN4BEG[2] ,
    \Tile_X4Y7_NN4BEG[1] ,
    \Tile_X4Y7_NN4BEG[0] }),
    .NN4END({\Tile_X4Y8_NN4BEG[15] ,
    \Tile_X4Y8_NN4BEG[14] ,
    \Tile_X4Y8_NN4BEG[13] ,
    \Tile_X4Y8_NN4BEG[12] ,
    \Tile_X4Y8_NN4BEG[11] ,
    \Tile_X4Y8_NN4BEG[10] ,
    \Tile_X4Y8_NN4BEG[9] ,
    \Tile_X4Y8_NN4BEG[8] ,
    \Tile_X4Y8_NN4BEG[7] ,
    \Tile_X4Y8_NN4BEG[6] ,
    \Tile_X4Y8_NN4BEG[5] ,
    \Tile_X4Y8_NN4BEG[4] ,
    \Tile_X4Y8_NN4BEG[3] ,
    \Tile_X4Y8_NN4BEG[2] ,
    \Tile_X4Y8_NN4BEG[1] ,
    \Tile_X4Y8_NN4BEG[0] }),
    .S1BEG({\Tile_X4Y7_S1BEG[3] ,
    \Tile_X4Y7_S1BEG[2] ,
    \Tile_X4Y7_S1BEG[1] ,
    \Tile_X4Y7_S1BEG[0] }),
    .S1END({\Tile_X4Y6_S1BEG[3] ,
    \Tile_X4Y6_S1BEG[2] ,
    \Tile_X4Y6_S1BEG[1] ,
    \Tile_X4Y6_S1BEG[0] }),
    .S2BEG({\Tile_X4Y7_S2BEG[7] ,
    \Tile_X4Y7_S2BEG[6] ,
    \Tile_X4Y7_S2BEG[5] ,
    \Tile_X4Y7_S2BEG[4] ,
    \Tile_X4Y7_S2BEG[3] ,
    \Tile_X4Y7_S2BEG[2] ,
    \Tile_X4Y7_S2BEG[1] ,
    \Tile_X4Y7_S2BEG[0] }),
    .S2BEGb({\Tile_X4Y7_S2BEGb[7] ,
    \Tile_X4Y7_S2BEGb[6] ,
    \Tile_X4Y7_S2BEGb[5] ,
    \Tile_X4Y7_S2BEGb[4] ,
    \Tile_X4Y7_S2BEGb[3] ,
    \Tile_X4Y7_S2BEGb[2] ,
    \Tile_X4Y7_S2BEGb[1] ,
    \Tile_X4Y7_S2BEGb[0] }),
    .S2END({\Tile_X4Y6_S2BEGb[7] ,
    \Tile_X4Y6_S2BEGb[6] ,
    \Tile_X4Y6_S2BEGb[5] ,
    \Tile_X4Y6_S2BEGb[4] ,
    \Tile_X4Y6_S2BEGb[3] ,
    \Tile_X4Y6_S2BEGb[2] ,
    \Tile_X4Y6_S2BEGb[1] ,
    \Tile_X4Y6_S2BEGb[0] }),
    .S2MID({\Tile_X4Y6_S2BEG[7] ,
    \Tile_X4Y6_S2BEG[6] ,
    \Tile_X4Y6_S2BEG[5] ,
    \Tile_X4Y6_S2BEG[4] ,
    \Tile_X4Y6_S2BEG[3] ,
    \Tile_X4Y6_S2BEG[2] ,
    \Tile_X4Y6_S2BEG[1] ,
    \Tile_X4Y6_S2BEG[0] }),
    .S4BEG({\Tile_X4Y7_S4BEG[15] ,
    \Tile_X4Y7_S4BEG[14] ,
    \Tile_X4Y7_S4BEG[13] ,
    \Tile_X4Y7_S4BEG[12] ,
    \Tile_X4Y7_S4BEG[11] ,
    \Tile_X4Y7_S4BEG[10] ,
    \Tile_X4Y7_S4BEG[9] ,
    \Tile_X4Y7_S4BEG[8] ,
    \Tile_X4Y7_S4BEG[7] ,
    \Tile_X4Y7_S4BEG[6] ,
    \Tile_X4Y7_S4BEG[5] ,
    \Tile_X4Y7_S4BEG[4] ,
    \Tile_X4Y7_S4BEG[3] ,
    \Tile_X4Y7_S4BEG[2] ,
    \Tile_X4Y7_S4BEG[1] ,
    \Tile_X4Y7_S4BEG[0] }),
    .S4END({\Tile_X4Y6_S4BEG[15] ,
    \Tile_X4Y6_S4BEG[14] ,
    \Tile_X4Y6_S4BEG[13] ,
    \Tile_X4Y6_S4BEG[12] ,
    \Tile_X4Y6_S4BEG[11] ,
    \Tile_X4Y6_S4BEG[10] ,
    \Tile_X4Y6_S4BEG[9] ,
    \Tile_X4Y6_S4BEG[8] ,
    \Tile_X4Y6_S4BEG[7] ,
    \Tile_X4Y6_S4BEG[6] ,
    \Tile_X4Y6_S4BEG[5] ,
    \Tile_X4Y6_S4BEG[4] ,
    \Tile_X4Y6_S4BEG[3] ,
    \Tile_X4Y6_S4BEG[2] ,
    \Tile_X4Y6_S4BEG[1] ,
    \Tile_X4Y6_S4BEG[0] }),
    .SS4BEG({\Tile_X4Y7_SS4BEG[15] ,
    \Tile_X4Y7_SS4BEG[14] ,
    \Tile_X4Y7_SS4BEG[13] ,
    \Tile_X4Y7_SS4BEG[12] ,
    \Tile_X4Y7_SS4BEG[11] ,
    \Tile_X4Y7_SS4BEG[10] ,
    \Tile_X4Y7_SS4BEG[9] ,
    \Tile_X4Y7_SS4BEG[8] ,
    \Tile_X4Y7_SS4BEG[7] ,
    \Tile_X4Y7_SS4BEG[6] ,
    \Tile_X4Y7_SS4BEG[5] ,
    \Tile_X4Y7_SS4BEG[4] ,
    \Tile_X4Y7_SS4BEG[3] ,
    \Tile_X4Y7_SS4BEG[2] ,
    \Tile_X4Y7_SS4BEG[1] ,
    \Tile_X4Y7_SS4BEG[0] }),
    .SS4END({\Tile_X4Y6_SS4BEG[15] ,
    \Tile_X4Y6_SS4BEG[14] ,
    \Tile_X4Y6_SS4BEG[13] ,
    \Tile_X4Y6_SS4BEG[12] ,
    \Tile_X4Y6_SS4BEG[11] ,
    \Tile_X4Y6_SS4BEG[10] ,
    \Tile_X4Y6_SS4BEG[9] ,
    \Tile_X4Y6_SS4BEG[8] ,
    \Tile_X4Y6_SS4BEG[7] ,
    \Tile_X4Y6_SS4BEG[6] ,
    \Tile_X4Y6_SS4BEG[5] ,
    \Tile_X4Y6_SS4BEG[4] ,
    \Tile_X4Y6_SS4BEG[3] ,
    \Tile_X4Y6_SS4BEG[2] ,
    \Tile_X4Y6_SS4BEG[1] ,
    \Tile_X4Y6_SS4BEG[0] }),
    .W1BEG({\Tile_X4Y7_W1BEG[3] ,
    \Tile_X4Y7_W1BEG[2] ,
    \Tile_X4Y7_W1BEG[1] ,
    \Tile_X4Y7_W1BEG[0] }),
    .W1END({\Tile_X5Y7_W1BEG[3] ,
    \Tile_X5Y7_W1BEG[2] ,
    \Tile_X5Y7_W1BEG[1] ,
    \Tile_X5Y7_W1BEG[0] }),
    .W2BEG({\Tile_X4Y7_W2BEG[7] ,
    \Tile_X4Y7_W2BEG[6] ,
    \Tile_X4Y7_W2BEG[5] ,
    \Tile_X4Y7_W2BEG[4] ,
    \Tile_X4Y7_W2BEG[3] ,
    \Tile_X4Y7_W2BEG[2] ,
    \Tile_X4Y7_W2BEG[1] ,
    \Tile_X4Y7_W2BEG[0] }),
    .W2BEGb({\Tile_X4Y7_W2BEGb[7] ,
    \Tile_X4Y7_W2BEGb[6] ,
    \Tile_X4Y7_W2BEGb[5] ,
    \Tile_X4Y7_W2BEGb[4] ,
    \Tile_X4Y7_W2BEGb[3] ,
    \Tile_X4Y7_W2BEGb[2] ,
    \Tile_X4Y7_W2BEGb[1] ,
    \Tile_X4Y7_W2BEGb[0] }),
    .W2END({\Tile_X5Y7_W2BEGb[7] ,
    \Tile_X5Y7_W2BEGb[6] ,
    \Tile_X5Y7_W2BEGb[5] ,
    \Tile_X5Y7_W2BEGb[4] ,
    \Tile_X5Y7_W2BEGb[3] ,
    \Tile_X5Y7_W2BEGb[2] ,
    \Tile_X5Y7_W2BEGb[1] ,
    \Tile_X5Y7_W2BEGb[0] }),
    .W2MID({\Tile_X5Y7_W2BEG[7] ,
    \Tile_X5Y7_W2BEG[6] ,
    \Tile_X5Y7_W2BEG[5] ,
    \Tile_X5Y7_W2BEG[4] ,
    \Tile_X5Y7_W2BEG[3] ,
    \Tile_X5Y7_W2BEG[2] ,
    \Tile_X5Y7_W2BEG[1] ,
    \Tile_X5Y7_W2BEG[0] }),
    .W6BEG({\Tile_X4Y7_W6BEG[11] ,
    \Tile_X4Y7_W6BEG[10] ,
    \Tile_X4Y7_W6BEG[9] ,
    \Tile_X4Y7_W6BEG[8] ,
    \Tile_X4Y7_W6BEG[7] ,
    \Tile_X4Y7_W6BEG[6] ,
    \Tile_X4Y7_W6BEG[5] ,
    \Tile_X4Y7_W6BEG[4] ,
    \Tile_X4Y7_W6BEG[3] ,
    \Tile_X4Y7_W6BEG[2] ,
    \Tile_X4Y7_W6BEG[1] ,
    \Tile_X4Y7_W6BEG[0] }),
    .W6END({\Tile_X5Y7_W6BEG[11] ,
    \Tile_X5Y7_W6BEG[10] ,
    \Tile_X5Y7_W6BEG[9] ,
    \Tile_X5Y7_W6BEG[8] ,
    \Tile_X5Y7_W6BEG[7] ,
    \Tile_X5Y7_W6BEG[6] ,
    \Tile_X5Y7_W6BEG[5] ,
    \Tile_X5Y7_W6BEG[4] ,
    \Tile_X5Y7_W6BEG[3] ,
    \Tile_X5Y7_W6BEG[2] ,
    \Tile_X5Y7_W6BEG[1] ,
    \Tile_X5Y7_W6BEG[0] }),
    .WW4BEG({\Tile_X4Y7_WW4BEG[15] ,
    \Tile_X4Y7_WW4BEG[14] ,
    \Tile_X4Y7_WW4BEG[13] ,
    \Tile_X4Y7_WW4BEG[12] ,
    \Tile_X4Y7_WW4BEG[11] ,
    \Tile_X4Y7_WW4BEG[10] ,
    \Tile_X4Y7_WW4BEG[9] ,
    \Tile_X4Y7_WW4BEG[8] ,
    \Tile_X4Y7_WW4BEG[7] ,
    \Tile_X4Y7_WW4BEG[6] ,
    \Tile_X4Y7_WW4BEG[5] ,
    \Tile_X4Y7_WW4BEG[4] ,
    \Tile_X4Y7_WW4BEG[3] ,
    \Tile_X4Y7_WW4BEG[2] ,
    \Tile_X4Y7_WW4BEG[1] ,
    \Tile_X4Y7_WW4BEG[0] }),
    .WW4END({\Tile_X5Y7_WW4BEG[15] ,
    \Tile_X5Y7_WW4BEG[14] ,
    \Tile_X5Y7_WW4BEG[13] ,
    \Tile_X5Y7_WW4BEG[12] ,
    \Tile_X5Y7_WW4BEG[11] ,
    \Tile_X5Y7_WW4BEG[10] ,
    \Tile_X5Y7_WW4BEG[9] ,
    \Tile_X5Y7_WW4BEG[8] ,
    \Tile_X5Y7_WW4BEG[7] ,
    \Tile_X5Y7_WW4BEG[6] ,
    \Tile_X5Y7_WW4BEG[5] ,
    \Tile_X5Y7_WW4BEG[4] ,
    \Tile_X5Y7_WW4BEG[3] ,
    \Tile_X5Y7_WW4BEG[2] ,
    \Tile_X5Y7_WW4BEG[1] ,
    \Tile_X5Y7_WW4BEG[0] }));
 LUT4AB Tile_X4Y8_LUT4AB (.Ci(Tile_X4Y9_Co),
    .Co(Tile_X4Y8_Co),
    .UserCLK(Tile_X4Y9_UserCLKo),
    .UserCLKo(Tile_X4Y8_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X4Y8_E1BEG[3] ,
    \Tile_X4Y8_E1BEG[2] ,
    \Tile_X4Y8_E1BEG[1] ,
    \Tile_X4Y8_E1BEG[0] }),
    .E1END({\Tile_X3Y8_E1BEG[3] ,
    \Tile_X3Y8_E1BEG[2] ,
    \Tile_X3Y8_E1BEG[1] ,
    \Tile_X3Y8_E1BEG[0] }),
    .E2BEG({\Tile_X4Y8_E2BEG[7] ,
    \Tile_X4Y8_E2BEG[6] ,
    \Tile_X4Y8_E2BEG[5] ,
    \Tile_X4Y8_E2BEG[4] ,
    \Tile_X4Y8_E2BEG[3] ,
    \Tile_X4Y8_E2BEG[2] ,
    \Tile_X4Y8_E2BEG[1] ,
    \Tile_X4Y8_E2BEG[0] }),
    .E2BEGb({\Tile_X4Y8_E2BEGb[7] ,
    \Tile_X4Y8_E2BEGb[6] ,
    \Tile_X4Y8_E2BEGb[5] ,
    \Tile_X4Y8_E2BEGb[4] ,
    \Tile_X4Y8_E2BEGb[3] ,
    \Tile_X4Y8_E2BEGb[2] ,
    \Tile_X4Y8_E2BEGb[1] ,
    \Tile_X4Y8_E2BEGb[0] }),
    .E2END({\Tile_X3Y8_E2BEGb[7] ,
    \Tile_X3Y8_E2BEGb[6] ,
    \Tile_X3Y8_E2BEGb[5] ,
    \Tile_X3Y8_E2BEGb[4] ,
    \Tile_X3Y8_E2BEGb[3] ,
    \Tile_X3Y8_E2BEGb[2] ,
    \Tile_X3Y8_E2BEGb[1] ,
    \Tile_X3Y8_E2BEGb[0] }),
    .E2MID({\Tile_X3Y8_E2BEG[7] ,
    \Tile_X3Y8_E2BEG[6] ,
    \Tile_X3Y8_E2BEG[5] ,
    \Tile_X3Y8_E2BEG[4] ,
    \Tile_X3Y8_E2BEG[3] ,
    \Tile_X3Y8_E2BEG[2] ,
    \Tile_X3Y8_E2BEG[1] ,
    \Tile_X3Y8_E2BEG[0] }),
    .E6BEG({\Tile_X4Y8_E6BEG[11] ,
    \Tile_X4Y8_E6BEG[10] ,
    \Tile_X4Y8_E6BEG[9] ,
    \Tile_X4Y8_E6BEG[8] ,
    \Tile_X4Y8_E6BEG[7] ,
    \Tile_X4Y8_E6BEG[6] ,
    \Tile_X4Y8_E6BEG[5] ,
    \Tile_X4Y8_E6BEG[4] ,
    \Tile_X4Y8_E6BEG[3] ,
    \Tile_X4Y8_E6BEG[2] ,
    \Tile_X4Y8_E6BEG[1] ,
    \Tile_X4Y8_E6BEG[0] }),
    .E6END({\Tile_X3Y8_E6BEG[11] ,
    \Tile_X3Y8_E6BEG[10] ,
    \Tile_X3Y8_E6BEG[9] ,
    \Tile_X3Y8_E6BEG[8] ,
    \Tile_X3Y8_E6BEG[7] ,
    \Tile_X3Y8_E6BEG[6] ,
    \Tile_X3Y8_E6BEG[5] ,
    \Tile_X3Y8_E6BEG[4] ,
    \Tile_X3Y8_E6BEG[3] ,
    \Tile_X3Y8_E6BEG[2] ,
    \Tile_X3Y8_E6BEG[1] ,
    \Tile_X3Y8_E6BEG[0] }),
    .EE4BEG({\Tile_X4Y8_EE4BEG[15] ,
    \Tile_X4Y8_EE4BEG[14] ,
    \Tile_X4Y8_EE4BEG[13] ,
    \Tile_X4Y8_EE4BEG[12] ,
    \Tile_X4Y8_EE4BEG[11] ,
    \Tile_X4Y8_EE4BEG[10] ,
    \Tile_X4Y8_EE4BEG[9] ,
    \Tile_X4Y8_EE4BEG[8] ,
    \Tile_X4Y8_EE4BEG[7] ,
    \Tile_X4Y8_EE4BEG[6] ,
    \Tile_X4Y8_EE4BEG[5] ,
    \Tile_X4Y8_EE4BEG[4] ,
    \Tile_X4Y8_EE4BEG[3] ,
    \Tile_X4Y8_EE4BEG[2] ,
    \Tile_X4Y8_EE4BEG[1] ,
    \Tile_X4Y8_EE4BEG[0] }),
    .EE4END({\Tile_X3Y8_EE4BEG[15] ,
    \Tile_X3Y8_EE4BEG[14] ,
    \Tile_X3Y8_EE4BEG[13] ,
    \Tile_X3Y8_EE4BEG[12] ,
    \Tile_X3Y8_EE4BEG[11] ,
    \Tile_X3Y8_EE4BEG[10] ,
    \Tile_X3Y8_EE4BEG[9] ,
    \Tile_X3Y8_EE4BEG[8] ,
    \Tile_X3Y8_EE4BEG[7] ,
    \Tile_X3Y8_EE4BEG[6] ,
    \Tile_X3Y8_EE4BEG[5] ,
    \Tile_X3Y8_EE4BEG[4] ,
    \Tile_X3Y8_EE4BEG[3] ,
    \Tile_X3Y8_EE4BEG[2] ,
    \Tile_X3Y8_EE4BEG[1] ,
    \Tile_X3Y8_EE4BEG[0] }),
    .FrameData({\Tile_X3Y8_FrameData_O[31] ,
    \Tile_X3Y8_FrameData_O[30] ,
    \Tile_X3Y8_FrameData_O[29] ,
    \Tile_X3Y8_FrameData_O[28] ,
    \Tile_X3Y8_FrameData_O[27] ,
    \Tile_X3Y8_FrameData_O[26] ,
    \Tile_X3Y8_FrameData_O[25] ,
    \Tile_X3Y8_FrameData_O[24] ,
    \Tile_X3Y8_FrameData_O[23] ,
    \Tile_X3Y8_FrameData_O[22] ,
    \Tile_X3Y8_FrameData_O[21] ,
    \Tile_X3Y8_FrameData_O[20] ,
    \Tile_X3Y8_FrameData_O[19] ,
    \Tile_X3Y8_FrameData_O[18] ,
    \Tile_X3Y8_FrameData_O[17] ,
    \Tile_X3Y8_FrameData_O[16] ,
    \Tile_X3Y8_FrameData_O[15] ,
    \Tile_X3Y8_FrameData_O[14] ,
    \Tile_X3Y8_FrameData_O[13] ,
    \Tile_X3Y8_FrameData_O[12] ,
    \Tile_X3Y8_FrameData_O[11] ,
    \Tile_X3Y8_FrameData_O[10] ,
    \Tile_X3Y8_FrameData_O[9] ,
    \Tile_X3Y8_FrameData_O[8] ,
    \Tile_X3Y8_FrameData_O[7] ,
    \Tile_X3Y8_FrameData_O[6] ,
    \Tile_X3Y8_FrameData_O[5] ,
    \Tile_X3Y8_FrameData_O[4] ,
    \Tile_X3Y8_FrameData_O[3] ,
    \Tile_X3Y8_FrameData_O[2] ,
    \Tile_X3Y8_FrameData_O[1] ,
    \Tile_X3Y8_FrameData_O[0] }),
    .FrameData_O({\Tile_X4Y8_FrameData_O[31] ,
    \Tile_X4Y8_FrameData_O[30] ,
    \Tile_X4Y8_FrameData_O[29] ,
    \Tile_X4Y8_FrameData_O[28] ,
    \Tile_X4Y8_FrameData_O[27] ,
    \Tile_X4Y8_FrameData_O[26] ,
    \Tile_X4Y8_FrameData_O[25] ,
    \Tile_X4Y8_FrameData_O[24] ,
    \Tile_X4Y8_FrameData_O[23] ,
    \Tile_X4Y8_FrameData_O[22] ,
    \Tile_X4Y8_FrameData_O[21] ,
    \Tile_X4Y8_FrameData_O[20] ,
    \Tile_X4Y8_FrameData_O[19] ,
    \Tile_X4Y8_FrameData_O[18] ,
    \Tile_X4Y8_FrameData_O[17] ,
    \Tile_X4Y8_FrameData_O[16] ,
    \Tile_X4Y8_FrameData_O[15] ,
    \Tile_X4Y8_FrameData_O[14] ,
    \Tile_X4Y8_FrameData_O[13] ,
    \Tile_X4Y8_FrameData_O[12] ,
    \Tile_X4Y8_FrameData_O[11] ,
    \Tile_X4Y8_FrameData_O[10] ,
    \Tile_X4Y8_FrameData_O[9] ,
    \Tile_X4Y8_FrameData_O[8] ,
    \Tile_X4Y8_FrameData_O[7] ,
    \Tile_X4Y8_FrameData_O[6] ,
    \Tile_X4Y8_FrameData_O[5] ,
    \Tile_X4Y8_FrameData_O[4] ,
    \Tile_X4Y8_FrameData_O[3] ,
    \Tile_X4Y8_FrameData_O[2] ,
    \Tile_X4Y8_FrameData_O[1] ,
    \Tile_X4Y8_FrameData_O[0] }),
    .FrameStrobe({\Tile_X4Y9_FrameStrobe_O[19] ,
    \Tile_X4Y9_FrameStrobe_O[18] ,
    \Tile_X4Y9_FrameStrobe_O[17] ,
    \Tile_X4Y9_FrameStrobe_O[16] ,
    \Tile_X4Y9_FrameStrobe_O[15] ,
    \Tile_X4Y9_FrameStrobe_O[14] ,
    \Tile_X4Y9_FrameStrobe_O[13] ,
    \Tile_X4Y9_FrameStrobe_O[12] ,
    \Tile_X4Y9_FrameStrobe_O[11] ,
    \Tile_X4Y9_FrameStrobe_O[10] ,
    \Tile_X4Y9_FrameStrobe_O[9] ,
    \Tile_X4Y9_FrameStrobe_O[8] ,
    \Tile_X4Y9_FrameStrobe_O[7] ,
    \Tile_X4Y9_FrameStrobe_O[6] ,
    \Tile_X4Y9_FrameStrobe_O[5] ,
    \Tile_X4Y9_FrameStrobe_O[4] ,
    \Tile_X4Y9_FrameStrobe_O[3] ,
    \Tile_X4Y9_FrameStrobe_O[2] ,
    \Tile_X4Y9_FrameStrobe_O[1] ,
    \Tile_X4Y9_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X4Y8_FrameStrobe_O[19] ,
    \Tile_X4Y8_FrameStrobe_O[18] ,
    \Tile_X4Y8_FrameStrobe_O[17] ,
    \Tile_X4Y8_FrameStrobe_O[16] ,
    \Tile_X4Y8_FrameStrobe_O[15] ,
    \Tile_X4Y8_FrameStrobe_O[14] ,
    \Tile_X4Y8_FrameStrobe_O[13] ,
    \Tile_X4Y8_FrameStrobe_O[12] ,
    \Tile_X4Y8_FrameStrobe_O[11] ,
    \Tile_X4Y8_FrameStrobe_O[10] ,
    \Tile_X4Y8_FrameStrobe_O[9] ,
    \Tile_X4Y8_FrameStrobe_O[8] ,
    \Tile_X4Y8_FrameStrobe_O[7] ,
    \Tile_X4Y8_FrameStrobe_O[6] ,
    \Tile_X4Y8_FrameStrobe_O[5] ,
    \Tile_X4Y8_FrameStrobe_O[4] ,
    \Tile_X4Y8_FrameStrobe_O[3] ,
    \Tile_X4Y8_FrameStrobe_O[2] ,
    \Tile_X4Y8_FrameStrobe_O[1] ,
    \Tile_X4Y8_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X4Y8_N1BEG[3] ,
    \Tile_X4Y8_N1BEG[2] ,
    \Tile_X4Y8_N1BEG[1] ,
    \Tile_X4Y8_N1BEG[0] }),
    .N1END({\Tile_X4Y9_N1BEG[3] ,
    \Tile_X4Y9_N1BEG[2] ,
    \Tile_X4Y9_N1BEG[1] ,
    \Tile_X4Y9_N1BEG[0] }),
    .N2BEG({\Tile_X4Y8_N2BEG[7] ,
    \Tile_X4Y8_N2BEG[6] ,
    \Tile_X4Y8_N2BEG[5] ,
    \Tile_X4Y8_N2BEG[4] ,
    \Tile_X4Y8_N2BEG[3] ,
    \Tile_X4Y8_N2BEG[2] ,
    \Tile_X4Y8_N2BEG[1] ,
    \Tile_X4Y8_N2BEG[0] }),
    .N2BEGb({\Tile_X4Y8_N2BEGb[7] ,
    \Tile_X4Y8_N2BEGb[6] ,
    \Tile_X4Y8_N2BEGb[5] ,
    \Tile_X4Y8_N2BEGb[4] ,
    \Tile_X4Y8_N2BEGb[3] ,
    \Tile_X4Y8_N2BEGb[2] ,
    \Tile_X4Y8_N2BEGb[1] ,
    \Tile_X4Y8_N2BEGb[0] }),
    .N2END({\Tile_X4Y9_N2BEGb[7] ,
    \Tile_X4Y9_N2BEGb[6] ,
    \Tile_X4Y9_N2BEGb[5] ,
    \Tile_X4Y9_N2BEGb[4] ,
    \Tile_X4Y9_N2BEGb[3] ,
    \Tile_X4Y9_N2BEGb[2] ,
    \Tile_X4Y9_N2BEGb[1] ,
    \Tile_X4Y9_N2BEGb[0] }),
    .N2MID({\Tile_X4Y9_N2BEG[7] ,
    \Tile_X4Y9_N2BEG[6] ,
    \Tile_X4Y9_N2BEG[5] ,
    \Tile_X4Y9_N2BEG[4] ,
    \Tile_X4Y9_N2BEG[3] ,
    \Tile_X4Y9_N2BEG[2] ,
    \Tile_X4Y9_N2BEG[1] ,
    \Tile_X4Y9_N2BEG[0] }),
    .N4BEG({\Tile_X4Y8_N4BEG[15] ,
    \Tile_X4Y8_N4BEG[14] ,
    \Tile_X4Y8_N4BEG[13] ,
    \Tile_X4Y8_N4BEG[12] ,
    \Tile_X4Y8_N4BEG[11] ,
    \Tile_X4Y8_N4BEG[10] ,
    \Tile_X4Y8_N4BEG[9] ,
    \Tile_X4Y8_N4BEG[8] ,
    \Tile_X4Y8_N4BEG[7] ,
    \Tile_X4Y8_N4BEG[6] ,
    \Tile_X4Y8_N4BEG[5] ,
    \Tile_X4Y8_N4BEG[4] ,
    \Tile_X4Y8_N4BEG[3] ,
    \Tile_X4Y8_N4BEG[2] ,
    \Tile_X4Y8_N4BEG[1] ,
    \Tile_X4Y8_N4BEG[0] }),
    .N4END({\Tile_X4Y9_N4BEG[15] ,
    \Tile_X4Y9_N4BEG[14] ,
    \Tile_X4Y9_N4BEG[13] ,
    \Tile_X4Y9_N4BEG[12] ,
    \Tile_X4Y9_N4BEG[11] ,
    \Tile_X4Y9_N4BEG[10] ,
    \Tile_X4Y9_N4BEG[9] ,
    \Tile_X4Y9_N4BEG[8] ,
    \Tile_X4Y9_N4BEG[7] ,
    \Tile_X4Y9_N4BEG[6] ,
    \Tile_X4Y9_N4BEG[5] ,
    \Tile_X4Y9_N4BEG[4] ,
    \Tile_X4Y9_N4BEG[3] ,
    \Tile_X4Y9_N4BEG[2] ,
    \Tile_X4Y9_N4BEG[1] ,
    \Tile_X4Y9_N4BEG[0] }),
    .NN4BEG({\Tile_X4Y8_NN4BEG[15] ,
    \Tile_X4Y8_NN4BEG[14] ,
    \Tile_X4Y8_NN4BEG[13] ,
    \Tile_X4Y8_NN4BEG[12] ,
    \Tile_X4Y8_NN4BEG[11] ,
    \Tile_X4Y8_NN4BEG[10] ,
    \Tile_X4Y8_NN4BEG[9] ,
    \Tile_X4Y8_NN4BEG[8] ,
    \Tile_X4Y8_NN4BEG[7] ,
    \Tile_X4Y8_NN4BEG[6] ,
    \Tile_X4Y8_NN4BEG[5] ,
    \Tile_X4Y8_NN4BEG[4] ,
    \Tile_X4Y8_NN4BEG[3] ,
    \Tile_X4Y8_NN4BEG[2] ,
    \Tile_X4Y8_NN4BEG[1] ,
    \Tile_X4Y8_NN4BEG[0] }),
    .NN4END({\Tile_X4Y9_NN4BEG[15] ,
    \Tile_X4Y9_NN4BEG[14] ,
    \Tile_X4Y9_NN4BEG[13] ,
    \Tile_X4Y9_NN4BEG[12] ,
    \Tile_X4Y9_NN4BEG[11] ,
    \Tile_X4Y9_NN4BEG[10] ,
    \Tile_X4Y9_NN4BEG[9] ,
    \Tile_X4Y9_NN4BEG[8] ,
    \Tile_X4Y9_NN4BEG[7] ,
    \Tile_X4Y9_NN4BEG[6] ,
    \Tile_X4Y9_NN4BEG[5] ,
    \Tile_X4Y9_NN4BEG[4] ,
    \Tile_X4Y9_NN4BEG[3] ,
    \Tile_X4Y9_NN4BEG[2] ,
    \Tile_X4Y9_NN4BEG[1] ,
    \Tile_X4Y9_NN4BEG[0] }),
    .S1BEG({\Tile_X4Y8_S1BEG[3] ,
    \Tile_X4Y8_S1BEG[2] ,
    \Tile_X4Y8_S1BEG[1] ,
    \Tile_X4Y8_S1BEG[0] }),
    .S1END({\Tile_X4Y7_S1BEG[3] ,
    \Tile_X4Y7_S1BEG[2] ,
    \Tile_X4Y7_S1BEG[1] ,
    \Tile_X4Y7_S1BEG[0] }),
    .S2BEG({\Tile_X4Y8_S2BEG[7] ,
    \Tile_X4Y8_S2BEG[6] ,
    \Tile_X4Y8_S2BEG[5] ,
    \Tile_X4Y8_S2BEG[4] ,
    \Tile_X4Y8_S2BEG[3] ,
    \Tile_X4Y8_S2BEG[2] ,
    \Tile_X4Y8_S2BEG[1] ,
    \Tile_X4Y8_S2BEG[0] }),
    .S2BEGb({\Tile_X4Y8_S2BEGb[7] ,
    \Tile_X4Y8_S2BEGb[6] ,
    \Tile_X4Y8_S2BEGb[5] ,
    \Tile_X4Y8_S2BEGb[4] ,
    \Tile_X4Y8_S2BEGb[3] ,
    \Tile_X4Y8_S2BEGb[2] ,
    \Tile_X4Y8_S2BEGb[1] ,
    \Tile_X4Y8_S2BEGb[0] }),
    .S2END({\Tile_X4Y7_S2BEGb[7] ,
    \Tile_X4Y7_S2BEGb[6] ,
    \Tile_X4Y7_S2BEGb[5] ,
    \Tile_X4Y7_S2BEGb[4] ,
    \Tile_X4Y7_S2BEGb[3] ,
    \Tile_X4Y7_S2BEGb[2] ,
    \Tile_X4Y7_S2BEGb[1] ,
    \Tile_X4Y7_S2BEGb[0] }),
    .S2MID({\Tile_X4Y7_S2BEG[7] ,
    \Tile_X4Y7_S2BEG[6] ,
    \Tile_X4Y7_S2BEG[5] ,
    \Tile_X4Y7_S2BEG[4] ,
    \Tile_X4Y7_S2BEG[3] ,
    \Tile_X4Y7_S2BEG[2] ,
    \Tile_X4Y7_S2BEG[1] ,
    \Tile_X4Y7_S2BEG[0] }),
    .S4BEG({\Tile_X4Y8_S4BEG[15] ,
    \Tile_X4Y8_S4BEG[14] ,
    \Tile_X4Y8_S4BEG[13] ,
    \Tile_X4Y8_S4BEG[12] ,
    \Tile_X4Y8_S4BEG[11] ,
    \Tile_X4Y8_S4BEG[10] ,
    \Tile_X4Y8_S4BEG[9] ,
    \Tile_X4Y8_S4BEG[8] ,
    \Tile_X4Y8_S4BEG[7] ,
    \Tile_X4Y8_S4BEG[6] ,
    \Tile_X4Y8_S4BEG[5] ,
    \Tile_X4Y8_S4BEG[4] ,
    \Tile_X4Y8_S4BEG[3] ,
    \Tile_X4Y8_S4BEG[2] ,
    \Tile_X4Y8_S4BEG[1] ,
    \Tile_X4Y8_S4BEG[0] }),
    .S4END({\Tile_X4Y7_S4BEG[15] ,
    \Tile_X4Y7_S4BEG[14] ,
    \Tile_X4Y7_S4BEG[13] ,
    \Tile_X4Y7_S4BEG[12] ,
    \Tile_X4Y7_S4BEG[11] ,
    \Tile_X4Y7_S4BEG[10] ,
    \Tile_X4Y7_S4BEG[9] ,
    \Tile_X4Y7_S4BEG[8] ,
    \Tile_X4Y7_S4BEG[7] ,
    \Tile_X4Y7_S4BEG[6] ,
    \Tile_X4Y7_S4BEG[5] ,
    \Tile_X4Y7_S4BEG[4] ,
    \Tile_X4Y7_S4BEG[3] ,
    \Tile_X4Y7_S4BEG[2] ,
    \Tile_X4Y7_S4BEG[1] ,
    \Tile_X4Y7_S4BEG[0] }),
    .SS4BEG({\Tile_X4Y8_SS4BEG[15] ,
    \Tile_X4Y8_SS4BEG[14] ,
    \Tile_X4Y8_SS4BEG[13] ,
    \Tile_X4Y8_SS4BEG[12] ,
    \Tile_X4Y8_SS4BEG[11] ,
    \Tile_X4Y8_SS4BEG[10] ,
    \Tile_X4Y8_SS4BEG[9] ,
    \Tile_X4Y8_SS4BEG[8] ,
    \Tile_X4Y8_SS4BEG[7] ,
    \Tile_X4Y8_SS4BEG[6] ,
    \Tile_X4Y8_SS4BEG[5] ,
    \Tile_X4Y8_SS4BEG[4] ,
    \Tile_X4Y8_SS4BEG[3] ,
    \Tile_X4Y8_SS4BEG[2] ,
    \Tile_X4Y8_SS4BEG[1] ,
    \Tile_X4Y8_SS4BEG[0] }),
    .SS4END({\Tile_X4Y7_SS4BEG[15] ,
    \Tile_X4Y7_SS4BEG[14] ,
    \Tile_X4Y7_SS4BEG[13] ,
    \Tile_X4Y7_SS4BEG[12] ,
    \Tile_X4Y7_SS4BEG[11] ,
    \Tile_X4Y7_SS4BEG[10] ,
    \Tile_X4Y7_SS4BEG[9] ,
    \Tile_X4Y7_SS4BEG[8] ,
    \Tile_X4Y7_SS4BEG[7] ,
    \Tile_X4Y7_SS4BEG[6] ,
    \Tile_X4Y7_SS4BEG[5] ,
    \Tile_X4Y7_SS4BEG[4] ,
    \Tile_X4Y7_SS4BEG[3] ,
    \Tile_X4Y7_SS4BEG[2] ,
    \Tile_X4Y7_SS4BEG[1] ,
    \Tile_X4Y7_SS4BEG[0] }),
    .W1BEG({\Tile_X4Y8_W1BEG[3] ,
    \Tile_X4Y8_W1BEG[2] ,
    \Tile_X4Y8_W1BEG[1] ,
    \Tile_X4Y8_W1BEG[0] }),
    .W1END({\Tile_X5Y8_W1BEG[3] ,
    \Tile_X5Y8_W1BEG[2] ,
    \Tile_X5Y8_W1BEG[1] ,
    \Tile_X5Y8_W1BEG[0] }),
    .W2BEG({\Tile_X4Y8_W2BEG[7] ,
    \Tile_X4Y8_W2BEG[6] ,
    \Tile_X4Y8_W2BEG[5] ,
    \Tile_X4Y8_W2BEG[4] ,
    \Tile_X4Y8_W2BEG[3] ,
    \Tile_X4Y8_W2BEG[2] ,
    \Tile_X4Y8_W2BEG[1] ,
    \Tile_X4Y8_W2BEG[0] }),
    .W2BEGb({\Tile_X4Y8_W2BEGb[7] ,
    \Tile_X4Y8_W2BEGb[6] ,
    \Tile_X4Y8_W2BEGb[5] ,
    \Tile_X4Y8_W2BEGb[4] ,
    \Tile_X4Y8_W2BEGb[3] ,
    \Tile_X4Y8_W2BEGb[2] ,
    \Tile_X4Y8_W2BEGb[1] ,
    \Tile_X4Y8_W2BEGb[0] }),
    .W2END({\Tile_X5Y8_W2BEGb[7] ,
    \Tile_X5Y8_W2BEGb[6] ,
    \Tile_X5Y8_W2BEGb[5] ,
    \Tile_X5Y8_W2BEGb[4] ,
    \Tile_X5Y8_W2BEGb[3] ,
    \Tile_X5Y8_W2BEGb[2] ,
    \Tile_X5Y8_W2BEGb[1] ,
    \Tile_X5Y8_W2BEGb[0] }),
    .W2MID({\Tile_X5Y8_W2BEG[7] ,
    \Tile_X5Y8_W2BEG[6] ,
    \Tile_X5Y8_W2BEG[5] ,
    \Tile_X5Y8_W2BEG[4] ,
    \Tile_X5Y8_W2BEG[3] ,
    \Tile_X5Y8_W2BEG[2] ,
    \Tile_X5Y8_W2BEG[1] ,
    \Tile_X5Y8_W2BEG[0] }),
    .W6BEG({\Tile_X4Y8_W6BEG[11] ,
    \Tile_X4Y8_W6BEG[10] ,
    \Tile_X4Y8_W6BEG[9] ,
    \Tile_X4Y8_W6BEG[8] ,
    \Tile_X4Y8_W6BEG[7] ,
    \Tile_X4Y8_W6BEG[6] ,
    \Tile_X4Y8_W6BEG[5] ,
    \Tile_X4Y8_W6BEG[4] ,
    \Tile_X4Y8_W6BEG[3] ,
    \Tile_X4Y8_W6BEG[2] ,
    \Tile_X4Y8_W6BEG[1] ,
    \Tile_X4Y8_W6BEG[0] }),
    .W6END({\Tile_X5Y8_W6BEG[11] ,
    \Tile_X5Y8_W6BEG[10] ,
    \Tile_X5Y8_W6BEG[9] ,
    \Tile_X5Y8_W6BEG[8] ,
    \Tile_X5Y8_W6BEG[7] ,
    \Tile_X5Y8_W6BEG[6] ,
    \Tile_X5Y8_W6BEG[5] ,
    \Tile_X5Y8_W6BEG[4] ,
    \Tile_X5Y8_W6BEG[3] ,
    \Tile_X5Y8_W6BEG[2] ,
    \Tile_X5Y8_W6BEG[1] ,
    \Tile_X5Y8_W6BEG[0] }),
    .WW4BEG({\Tile_X4Y8_WW4BEG[15] ,
    \Tile_X4Y8_WW4BEG[14] ,
    \Tile_X4Y8_WW4BEG[13] ,
    \Tile_X4Y8_WW4BEG[12] ,
    \Tile_X4Y8_WW4BEG[11] ,
    \Tile_X4Y8_WW4BEG[10] ,
    \Tile_X4Y8_WW4BEG[9] ,
    \Tile_X4Y8_WW4BEG[8] ,
    \Tile_X4Y8_WW4BEG[7] ,
    \Tile_X4Y8_WW4BEG[6] ,
    \Tile_X4Y8_WW4BEG[5] ,
    \Tile_X4Y8_WW4BEG[4] ,
    \Tile_X4Y8_WW4BEG[3] ,
    \Tile_X4Y8_WW4BEG[2] ,
    \Tile_X4Y8_WW4BEG[1] ,
    \Tile_X4Y8_WW4BEG[0] }),
    .WW4END({\Tile_X5Y8_WW4BEG[15] ,
    \Tile_X5Y8_WW4BEG[14] ,
    \Tile_X5Y8_WW4BEG[13] ,
    \Tile_X5Y8_WW4BEG[12] ,
    \Tile_X5Y8_WW4BEG[11] ,
    \Tile_X5Y8_WW4BEG[10] ,
    \Tile_X5Y8_WW4BEG[9] ,
    \Tile_X5Y8_WW4BEG[8] ,
    \Tile_X5Y8_WW4BEG[7] ,
    \Tile_X5Y8_WW4BEG[6] ,
    \Tile_X5Y8_WW4BEG[5] ,
    \Tile_X5Y8_WW4BEG[4] ,
    \Tile_X5Y8_WW4BEG[3] ,
    \Tile_X5Y8_WW4BEG[2] ,
    \Tile_X5Y8_WW4BEG[1] ,
    \Tile_X5Y8_WW4BEG[0] }));
 S_IO4 Tile_X4Y9_S_IO4 (.A_I_top(Tile_X4Y9_A_I_top),
    .A_O_top(Tile_X4Y9_A_O_top),
    .A_T_top(Tile_X4Y9_A_T_top),
    .B_I_top(Tile_X4Y9_B_I_top),
    .B_O_top(Tile_X4Y9_B_O_top),
    .B_T_top(Tile_X4Y9_B_T_top),
    .C_I_top(Tile_X4Y9_C_I_top),
    .C_O_top(Tile_X4Y9_C_O_top),
    .C_T_top(Tile_X4Y9_C_T_top),
    .Co(Tile_X4Y9_Co),
    .D_I_top(Tile_X4Y9_D_I_top),
    .D_O_top(Tile_X4Y9_D_O_top),
    .D_T_top(Tile_X4Y9_D_T_top),
    .UserCLK(UserCLK),
    .UserCLKo(Tile_X4Y9_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .FrameData({\Tile_X3Y9_FrameData_O[31] ,
    \Tile_X3Y9_FrameData_O[30] ,
    \Tile_X3Y9_FrameData_O[29] ,
    \Tile_X3Y9_FrameData_O[28] ,
    \Tile_X3Y9_FrameData_O[27] ,
    \Tile_X3Y9_FrameData_O[26] ,
    \Tile_X3Y9_FrameData_O[25] ,
    \Tile_X3Y9_FrameData_O[24] ,
    \Tile_X3Y9_FrameData_O[23] ,
    \Tile_X3Y9_FrameData_O[22] ,
    \Tile_X3Y9_FrameData_O[21] ,
    \Tile_X3Y9_FrameData_O[20] ,
    \Tile_X3Y9_FrameData_O[19] ,
    \Tile_X3Y9_FrameData_O[18] ,
    \Tile_X3Y9_FrameData_O[17] ,
    \Tile_X3Y9_FrameData_O[16] ,
    \Tile_X3Y9_FrameData_O[15] ,
    \Tile_X3Y9_FrameData_O[14] ,
    \Tile_X3Y9_FrameData_O[13] ,
    \Tile_X3Y9_FrameData_O[12] ,
    \Tile_X3Y9_FrameData_O[11] ,
    \Tile_X3Y9_FrameData_O[10] ,
    \Tile_X3Y9_FrameData_O[9] ,
    \Tile_X3Y9_FrameData_O[8] ,
    \Tile_X3Y9_FrameData_O[7] ,
    \Tile_X3Y9_FrameData_O[6] ,
    \Tile_X3Y9_FrameData_O[5] ,
    \Tile_X3Y9_FrameData_O[4] ,
    \Tile_X3Y9_FrameData_O[3] ,
    \Tile_X3Y9_FrameData_O[2] ,
    \Tile_X3Y9_FrameData_O[1] ,
    \Tile_X3Y9_FrameData_O[0] }),
    .FrameData_O({\Tile_X4Y9_FrameData_O[31] ,
    \Tile_X4Y9_FrameData_O[30] ,
    \Tile_X4Y9_FrameData_O[29] ,
    \Tile_X4Y9_FrameData_O[28] ,
    \Tile_X4Y9_FrameData_O[27] ,
    \Tile_X4Y9_FrameData_O[26] ,
    \Tile_X4Y9_FrameData_O[25] ,
    \Tile_X4Y9_FrameData_O[24] ,
    \Tile_X4Y9_FrameData_O[23] ,
    \Tile_X4Y9_FrameData_O[22] ,
    \Tile_X4Y9_FrameData_O[21] ,
    \Tile_X4Y9_FrameData_O[20] ,
    \Tile_X4Y9_FrameData_O[19] ,
    \Tile_X4Y9_FrameData_O[18] ,
    \Tile_X4Y9_FrameData_O[17] ,
    \Tile_X4Y9_FrameData_O[16] ,
    \Tile_X4Y9_FrameData_O[15] ,
    \Tile_X4Y9_FrameData_O[14] ,
    \Tile_X4Y9_FrameData_O[13] ,
    \Tile_X4Y9_FrameData_O[12] ,
    \Tile_X4Y9_FrameData_O[11] ,
    \Tile_X4Y9_FrameData_O[10] ,
    \Tile_X4Y9_FrameData_O[9] ,
    \Tile_X4Y9_FrameData_O[8] ,
    \Tile_X4Y9_FrameData_O[7] ,
    \Tile_X4Y9_FrameData_O[6] ,
    \Tile_X4Y9_FrameData_O[5] ,
    \Tile_X4Y9_FrameData_O[4] ,
    \Tile_X4Y9_FrameData_O[3] ,
    \Tile_X4Y9_FrameData_O[2] ,
    \Tile_X4Y9_FrameData_O[1] ,
    \Tile_X4Y9_FrameData_O[0] }),
    .FrameStrobe({FrameStrobe[99],
    FrameStrobe[98],
    FrameStrobe[97],
    FrameStrobe[96],
    FrameStrobe[95],
    FrameStrobe[94],
    FrameStrobe[93],
    FrameStrobe[92],
    FrameStrobe[91],
    FrameStrobe[90],
    FrameStrobe[89],
    FrameStrobe[88],
    FrameStrobe[87],
    FrameStrobe[86],
    FrameStrobe[85],
    FrameStrobe[84],
    FrameStrobe[83],
    FrameStrobe[82],
    FrameStrobe[81],
    FrameStrobe[80]}),
    .FrameStrobe_O({\Tile_X4Y9_FrameStrobe_O[19] ,
    \Tile_X4Y9_FrameStrobe_O[18] ,
    \Tile_X4Y9_FrameStrobe_O[17] ,
    \Tile_X4Y9_FrameStrobe_O[16] ,
    \Tile_X4Y9_FrameStrobe_O[15] ,
    \Tile_X4Y9_FrameStrobe_O[14] ,
    \Tile_X4Y9_FrameStrobe_O[13] ,
    \Tile_X4Y9_FrameStrobe_O[12] ,
    \Tile_X4Y9_FrameStrobe_O[11] ,
    \Tile_X4Y9_FrameStrobe_O[10] ,
    \Tile_X4Y9_FrameStrobe_O[9] ,
    \Tile_X4Y9_FrameStrobe_O[8] ,
    \Tile_X4Y9_FrameStrobe_O[7] ,
    \Tile_X4Y9_FrameStrobe_O[6] ,
    \Tile_X4Y9_FrameStrobe_O[5] ,
    \Tile_X4Y9_FrameStrobe_O[4] ,
    \Tile_X4Y9_FrameStrobe_O[3] ,
    \Tile_X4Y9_FrameStrobe_O[2] ,
    \Tile_X4Y9_FrameStrobe_O[1] ,
    \Tile_X4Y9_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X4Y9_N1BEG[3] ,
    \Tile_X4Y9_N1BEG[2] ,
    \Tile_X4Y9_N1BEG[1] ,
    \Tile_X4Y9_N1BEG[0] }),
    .N2BEG({\Tile_X4Y9_N2BEG[7] ,
    \Tile_X4Y9_N2BEG[6] ,
    \Tile_X4Y9_N2BEG[5] ,
    \Tile_X4Y9_N2BEG[4] ,
    \Tile_X4Y9_N2BEG[3] ,
    \Tile_X4Y9_N2BEG[2] ,
    \Tile_X4Y9_N2BEG[1] ,
    \Tile_X4Y9_N2BEG[0] }),
    .N2BEGb({\Tile_X4Y9_N2BEGb[7] ,
    \Tile_X4Y9_N2BEGb[6] ,
    \Tile_X4Y9_N2BEGb[5] ,
    \Tile_X4Y9_N2BEGb[4] ,
    \Tile_X4Y9_N2BEGb[3] ,
    \Tile_X4Y9_N2BEGb[2] ,
    \Tile_X4Y9_N2BEGb[1] ,
    \Tile_X4Y9_N2BEGb[0] }),
    .N4BEG({\Tile_X4Y9_N4BEG[15] ,
    \Tile_X4Y9_N4BEG[14] ,
    \Tile_X4Y9_N4BEG[13] ,
    \Tile_X4Y9_N4BEG[12] ,
    \Tile_X4Y9_N4BEG[11] ,
    \Tile_X4Y9_N4BEG[10] ,
    \Tile_X4Y9_N4BEG[9] ,
    \Tile_X4Y9_N4BEG[8] ,
    \Tile_X4Y9_N4BEG[7] ,
    \Tile_X4Y9_N4BEG[6] ,
    \Tile_X4Y9_N4BEG[5] ,
    \Tile_X4Y9_N4BEG[4] ,
    \Tile_X4Y9_N4BEG[3] ,
    \Tile_X4Y9_N4BEG[2] ,
    \Tile_X4Y9_N4BEG[1] ,
    \Tile_X4Y9_N4BEG[0] }),
    .NN4BEG({\Tile_X4Y9_NN4BEG[15] ,
    \Tile_X4Y9_NN4BEG[14] ,
    \Tile_X4Y9_NN4BEG[13] ,
    \Tile_X4Y9_NN4BEG[12] ,
    \Tile_X4Y9_NN4BEG[11] ,
    \Tile_X4Y9_NN4BEG[10] ,
    \Tile_X4Y9_NN4BEG[9] ,
    \Tile_X4Y9_NN4BEG[8] ,
    \Tile_X4Y9_NN4BEG[7] ,
    \Tile_X4Y9_NN4BEG[6] ,
    \Tile_X4Y9_NN4BEG[5] ,
    \Tile_X4Y9_NN4BEG[4] ,
    \Tile_X4Y9_NN4BEG[3] ,
    \Tile_X4Y9_NN4BEG[2] ,
    \Tile_X4Y9_NN4BEG[1] ,
    \Tile_X4Y9_NN4BEG[0] }),
    .S1END({\Tile_X4Y8_S1BEG[3] ,
    \Tile_X4Y8_S1BEG[2] ,
    \Tile_X4Y8_S1BEG[1] ,
    \Tile_X4Y8_S1BEG[0] }),
    .S2END({\Tile_X4Y8_S2BEGb[7] ,
    \Tile_X4Y8_S2BEGb[6] ,
    \Tile_X4Y8_S2BEGb[5] ,
    \Tile_X4Y8_S2BEGb[4] ,
    \Tile_X4Y8_S2BEGb[3] ,
    \Tile_X4Y8_S2BEGb[2] ,
    \Tile_X4Y8_S2BEGb[1] ,
    \Tile_X4Y8_S2BEGb[0] }),
    .S2MID({\Tile_X4Y8_S2BEG[7] ,
    \Tile_X4Y8_S2BEG[6] ,
    \Tile_X4Y8_S2BEG[5] ,
    \Tile_X4Y8_S2BEG[4] ,
    \Tile_X4Y8_S2BEG[3] ,
    \Tile_X4Y8_S2BEG[2] ,
    \Tile_X4Y8_S2BEG[1] ,
    \Tile_X4Y8_S2BEG[0] }),
    .S4END({\Tile_X4Y8_S4BEG[15] ,
    \Tile_X4Y8_S4BEG[14] ,
    \Tile_X4Y8_S4BEG[13] ,
    \Tile_X4Y8_S4BEG[12] ,
    \Tile_X4Y8_S4BEG[11] ,
    \Tile_X4Y8_S4BEG[10] ,
    \Tile_X4Y8_S4BEG[9] ,
    \Tile_X4Y8_S4BEG[8] ,
    \Tile_X4Y8_S4BEG[7] ,
    \Tile_X4Y8_S4BEG[6] ,
    \Tile_X4Y8_S4BEG[5] ,
    \Tile_X4Y8_S4BEG[4] ,
    \Tile_X4Y8_S4BEG[3] ,
    \Tile_X4Y8_S4BEG[2] ,
    \Tile_X4Y8_S4BEG[1] ,
    \Tile_X4Y8_S4BEG[0] }),
    .SS4END({\Tile_X4Y8_SS4BEG[15] ,
    \Tile_X4Y8_SS4BEG[14] ,
    \Tile_X4Y8_SS4BEG[13] ,
    \Tile_X4Y8_SS4BEG[12] ,
    \Tile_X4Y8_SS4BEG[11] ,
    \Tile_X4Y8_SS4BEG[10] ,
    \Tile_X4Y8_SS4BEG[9] ,
    \Tile_X4Y8_SS4BEG[8] ,
    \Tile_X4Y8_SS4BEG[7] ,
    \Tile_X4Y8_SS4BEG[6] ,
    \Tile_X4Y8_SS4BEG[5] ,
    \Tile_X4Y8_SS4BEG[4] ,
    \Tile_X4Y8_SS4BEG[3] ,
    \Tile_X4Y8_SS4BEG[2] ,
    \Tile_X4Y8_SS4BEG[1] ,
    \Tile_X4Y8_SS4BEG[0] }));
 NE_term Tile_X5Y0_NE_term (.UserCLK(Tile_X5Y1_UserCLKo),
    .UserCLKo(Tile_X5Y0_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .FrameData({\Tile_X4Y0_FrameData_O[31] ,
    \Tile_X4Y0_FrameData_O[30] ,
    \Tile_X4Y0_FrameData_O[29] ,
    \Tile_X4Y0_FrameData_O[28] ,
    \Tile_X4Y0_FrameData_O[27] ,
    \Tile_X4Y0_FrameData_O[26] ,
    \Tile_X4Y0_FrameData_O[25] ,
    \Tile_X4Y0_FrameData_O[24] ,
    \Tile_X4Y0_FrameData_O[23] ,
    \Tile_X4Y0_FrameData_O[22] ,
    \Tile_X4Y0_FrameData_O[21] ,
    \Tile_X4Y0_FrameData_O[20] ,
    \Tile_X4Y0_FrameData_O[19] ,
    \Tile_X4Y0_FrameData_O[18] ,
    \Tile_X4Y0_FrameData_O[17] ,
    \Tile_X4Y0_FrameData_O[16] ,
    \Tile_X4Y0_FrameData_O[15] ,
    \Tile_X4Y0_FrameData_O[14] ,
    \Tile_X4Y0_FrameData_O[13] ,
    \Tile_X4Y0_FrameData_O[12] ,
    \Tile_X4Y0_FrameData_O[11] ,
    \Tile_X4Y0_FrameData_O[10] ,
    \Tile_X4Y0_FrameData_O[9] ,
    \Tile_X4Y0_FrameData_O[8] ,
    \Tile_X4Y0_FrameData_O[7] ,
    \Tile_X4Y0_FrameData_O[6] ,
    \Tile_X4Y0_FrameData_O[5] ,
    \Tile_X4Y0_FrameData_O[4] ,
    \Tile_X4Y0_FrameData_O[3] ,
    \Tile_X4Y0_FrameData_O[2] ,
    \Tile_X4Y0_FrameData_O[1] ,
    \Tile_X4Y0_FrameData_O[0] }),
    .FrameData_O({\Tile_X5Y0_FrameData_O[31] ,
    \Tile_X5Y0_FrameData_O[30] ,
    \Tile_X5Y0_FrameData_O[29] ,
    \Tile_X5Y0_FrameData_O[28] ,
    \Tile_X5Y0_FrameData_O[27] ,
    \Tile_X5Y0_FrameData_O[26] ,
    \Tile_X5Y0_FrameData_O[25] ,
    \Tile_X5Y0_FrameData_O[24] ,
    \Tile_X5Y0_FrameData_O[23] ,
    \Tile_X5Y0_FrameData_O[22] ,
    \Tile_X5Y0_FrameData_O[21] ,
    \Tile_X5Y0_FrameData_O[20] ,
    \Tile_X5Y0_FrameData_O[19] ,
    \Tile_X5Y0_FrameData_O[18] ,
    \Tile_X5Y0_FrameData_O[17] ,
    \Tile_X5Y0_FrameData_O[16] ,
    \Tile_X5Y0_FrameData_O[15] ,
    \Tile_X5Y0_FrameData_O[14] ,
    \Tile_X5Y0_FrameData_O[13] ,
    \Tile_X5Y0_FrameData_O[12] ,
    \Tile_X5Y0_FrameData_O[11] ,
    \Tile_X5Y0_FrameData_O[10] ,
    \Tile_X5Y0_FrameData_O[9] ,
    \Tile_X5Y0_FrameData_O[8] ,
    \Tile_X5Y0_FrameData_O[7] ,
    \Tile_X5Y0_FrameData_O[6] ,
    \Tile_X5Y0_FrameData_O[5] ,
    \Tile_X5Y0_FrameData_O[4] ,
    \Tile_X5Y0_FrameData_O[3] ,
    \Tile_X5Y0_FrameData_O[2] ,
    \Tile_X5Y0_FrameData_O[1] ,
    \Tile_X5Y0_FrameData_O[0] }),
    .FrameStrobe({\Tile_X5Y1_FrameStrobe_O[19] ,
    \Tile_X5Y1_FrameStrobe_O[18] ,
    \Tile_X5Y1_FrameStrobe_O[17] ,
    \Tile_X5Y1_FrameStrobe_O[16] ,
    \Tile_X5Y1_FrameStrobe_O[15] ,
    \Tile_X5Y1_FrameStrobe_O[14] ,
    \Tile_X5Y1_FrameStrobe_O[13] ,
    \Tile_X5Y1_FrameStrobe_O[12] ,
    \Tile_X5Y1_FrameStrobe_O[11] ,
    \Tile_X5Y1_FrameStrobe_O[10] ,
    \Tile_X5Y1_FrameStrobe_O[9] ,
    \Tile_X5Y1_FrameStrobe_O[8] ,
    \Tile_X5Y1_FrameStrobe_O[7] ,
    \Tile_X5Y1_FrameStrobe_O[6] ,
    \Tile_X5Y1_FrameStrobe_O[5] ,
    \Tile_X5Y1_FrameStrobe_O[4] ,
    \Tile_X5Y1_FrameStrobe_O[3] ,
    \Tile_X5Y1_FrameStrobe_O[2] ,
    \Tile_X5Y1_FrameStrobe_O[1] ,
    \Tile_X5Y1_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X5Y0_FrameStrobe_O[19] ,
    \Tile_X5Y0_FrameStrobe_O[18] ,
    \Tile_X5Y0_FrameStrobe_O[17] ,
    \Tile_X5Y0_FrameStrobe_O[16] ,
    \Tile_X5Y0_FrameStrobe_O[15] ,
    \Tile_X5Y0_FrameStrobe_O[14] ,
    \Tile_X5Y0_FrameStrobe_O[13] ,
    \Tile_X5Y0_FrameStrobe_O[12] ,
    \Tile_X5Y0_FrameStrobe_O[11] ,
    \Tile_X5Y0_FrameStrobe_O[10] ,
    \Tile_X5Y0_FrameStrobe_O[9] ,
    \Tile_X5Y0_FrameStrobe_O[8] ,
    \Tile_X5Y0_FrameStrobe_O[7] ,
    \Tile_X5Y0_FrameStrobe_O[6] ,
    \Tile_X5Y0_FrameStrobe_O[5] ,
    \Tile_X5Y0_FrameStrobe_O[4] ,
    \Tile_X5Y0_FrameStrobe_O[3] ,
    \Tile_X5Y0_FrameStrobe_O[2] ,
    \Tile_X5Y0_FrameStrobe_O[1] ,
    \Tile_X5Y0_FrameStrobe_O[0] }),
    .N1END({\Tile_X5Y1_N1BEG[3] ,
    \Tile_X5Y1_N1BEG[2] ,
    \Tile_X5Y1_N1BEG[1] ,
    \Tile_X5Y1_N1BEG[0] }),
    .N2END({\Tile_X5Y1_N2BEGb[7] ,
    \Tile_X5Y1_N2BEGb[6] ,
    \Tile_X5Y1_N2BEGb[5] ,
    \Tile_X5Y1_N2BEGb[4] ,
    \Tile_X5Y1_N2BEGb[3] ,
    \Tile_X5Y1_N2BEGb[2] ,
    \Tile_X5Y1_N2BEGb[1] ,
    \Tile_X5Y1_N2BEGb[0] }),
    .N2MID({\Tile_X5Y1_N2BEG[7] ,
    \Tile_X5Y1_N2BEG[6] ,
    \Tile_X5Y1_N2BEG[5] ,
    \Tile_X5Y1_N2BEG[4] ,
    \Tile_X5Y1_N2BEG[3] ,
    \Tile_X5Y1_N2BEG[2] ,
    \Tile_X5Y1_N2BEG[1] ,
    \Tile_X5Y1_N2BEG[0] }),
    .N4END({\Tile_X5Y1_N4BEG[15] ,
    \Tile_X5Y1_N4BEG[14] ,
    \Tile_X5Y1_N4BEG[13] ,
    \Tile_X5Y1_N4BEG[12] ,
    \Tile_X5Y1_N4BEG[11] ,
    \Tile_X5Y1_N4BEG[10] ,
    \Tile_X5Y1_N4BEG[9] ,
    \Tile_X5Y1_N4BEG[8] ,
    \Tile_X5Y1_N4BEG[7] ,
    \Tile_X5Y1_N4BEG[6] ,
    \Tile_X5Y1_N4BEG[5] ,
    \Tile_X5Y1_N4BEG[4] ,
    \Tile_X5Y1_N4BEG[3] ,
    \Tile_X5Y1_N4BEG[2] ,
    \Tile_X5Y1_N4BEG[1] ,
    \Tile_X5Y1_N4BEG[0] }),
    .S1BEG({\Tile_X5Y0_S1BEG[3] ,
    \Tile_X5Y0_S1BEG[2] ,
    \Tile_X5Y0_S1BEG[1] ,
    \Tile_X5Y0_S1BEG[0] }),
    .S2BEG({\Tile_X5Y0_S2BEG[7] ,
    \Tile_X5Y0_S2BEG[6] ,
    \Tile_X5Y0_S2BEG[5] ,
    \Tile_X5Y0_S2BEG[4] ,
    \Tile_X5Y0_S2BEG[3] ,
    \Tile_X5Y0_S2BEG[2] ,
    \Tile_X5Y0_S2BEG[1] ,
    \Tile_X5Y0_S2BEG[0] }),
    .S2BEGb({\Tile_X5Y0_S2BEGb[7] ,
    \Tile_X5Y0_S2BEGb[6] ,
    \Tile_X5Y0_S2BEGb[5] ,
    \Tile_X5Y0_S2BEGb[4] ,
    \Tile_X5Y0_S2BEGb[3] ,
    \Tile_X5Y0_S2BEGb[2] ,
    \Tile_X5Y0_S2BEGb[1] ,
    \Tile_X5Y0_S2BEGb[0] }),
    .S4BEG({\Tile_X5Y0_S4BEG[15] ,
    \Tile_X5Y0_S4BEG[14] ,
    \Tile_X5Y0_S4BEG[13] ,
    \Tile_X5Y0_S4BEG[12] ,
    \Tile_X5Y0_S4BEG[11] ,
    \Tile_X5Y0_S4BEG[10] ,
    \Tile_X5Y0_S4BEG[9] ,
    \Tile_X5Y0_S4BEG[8] ,
    \Tile_X5Y0_S4BEG[7] ,
    \Tile_X5Y0_S4BEG[6] ,
    \Tile_X5Y0_S4BEG[5] ,
    \Tile_X5Y0_S4BEG[4] ,
    \Tile_X5Y0_S4BEG[3] ,
    \Tile_X5Y0_S4BEG[2] ,
    \Tile_X5Y0_S4BEG[1] ,
    \Tile_X5Y0_S4BEG[0] }));
 IHP_SRAM Tile_X5Y1_IHP_SRAM (.ADDR_SRAM0(Tile_X5Y2_ADDR_SRAM0),
    .ADDR_SRAM1(Tile_X5Y2_ADDR_SRAM1),
    .ADDR_SRAM2(Tile_X5Y2_ADDR_SRAM2),
    .ADDR_SRAM3(Tile_X5Y2_ADDR_SRAM3),
    .ADDR_SRAM4(Tile_X5Y2_ADDR_SRAM4),
    .ADDR_SRAM5(Tile_X5Y2_ADDR_SRAM5),
    .ADDR_SRAM6(Tile_X5Y2_ADDR_SRAM6),
    .ADDR_SRAM7(Tile_X5Y2_ADDR_SRAM7),
    .ADDR_SRAM8(Tile_X5Y2_ADDR_SRAM8),
    .ADDR_SRAM9(Tile_X5Y2_ADDR_SRAM9),
    .BM_SRAM0(Tile_X5Y2_BM_SRAM0),
    .BM_SRAM1(Tile_X5Y2_BM_SRAM1),
    .BM_SRAM10(Tile_X5Y2_BM_SRAM10),
    .BM_SRAM11(Tile_X5Y2_BM_SRAM11),
    .BM_SRAM12(Tile_X5Y2_BM_SRAM12),
    .BM_SRAM13(Tile_X5Y2_BM_SRAM13),
    .BM_SRAM14(Tile_X5Y2_BM_SRAM14),
    .BM_SRAM15(Tile_X5Y2_BM_SRAM15),
    .BM_SRAM16(Tile_X5Y2_BM_SRAM16),
    .BM_SRAM17(Tile_X5Y2_BM_SRAM17),
    .BM_SRAM18(Tile_X5Y2_BM_SRAM18),
    .BM_SRAM19(Tile_X5Y2_BM_SRAM19),
    .BM_SRAM2(Tile_X5Y2_BM_SRAM2),
    .BM_SRAM20(Tile_X5Y2_BM_SRAM20),
    .BM_SRAM21(Tile_X5Y2_BM_SRAM21),
    .BM_SRAM22(Tile_X5Y2_BM_SRAM22),
    .BM_SRAM23(Tile_X5Y2_BM_SRAM23),
    .BM_SRAM24(Tile_X5Y2_BM_SRAM24),
    .BM_SRAM25(Tile_X5Y2_BM_SRAM25),
    .BM_SRAM26(Tile_X5Y2_BM_SRAM26),
    .BM_SRAM27(Tile_X5Y2_BM_SRAM27),
    .BM_SRAM28(Tile_X5Y2_BM_SRAM28),
    .BM_SRAM29(Tile_X5Y2_BM_SRAM29),
    .BM_SRAM3(Tile_X5Y2_BM_SRAM3),
    .BM_SRAM30(Tile_X5Y2_BM_SRAM30),
    .BM_SRAM31(Tile_X5Y2_BM_SRAM31),
    .BM_SRAM4(Tile_X5Y2_BM_SRAM4),
    .BM_SRAM5(Tile_X5Y2_BM_SRAM5),
    .BM_SRAM6(Tile_X5Y2_BM_SRAM6),
    .BM_SRAM7(Tile_X5Y2_BM_SRAM7),
    .BM_SRAM8(Tile_X5Y2_BM_SRAM8),
    .BM_SRAM9(Tile_X5Y2_BM_SRAM9),
    .CLK_SRAM(Tile_X5Y2_CLK_SRAM),
    .CONFIGURED_top(Tile_X5Y2_CONFIGURED_top),
    .DIN_SRAM0(Tile_X5Y2_DIN_SRAM0),
    .DIN_SRAM1(Tile_X5Y2_DIN_SRAM1),
    .DIN_SRAM10(Tile_X5Y2_DIN_SRAM10),
    .DIN_SRAM11(Tile_X5Y2_DIN_SRAM11),
    .DIN_SRAM12(Tile_X5Y2_DIN_SRAM12),
    .DIN_SRAM13(Tile_X5Y2_DIN_SRAM13),
    .DIN_SRAM14(Tile_X5Y2_DIN_SRAM14),
    .DIN_SRAM15(Tile_X5Y2_DIN_SRAM15),
    .DIN_SRAM16(Tile_X5Y2_DIN_SRAM16),
    .DIN_SRAM17(Tile_X5Y2_DIN_SRAM17),
    .DIN_SRAM18(Tile_X5Y2_DIN_SRAM18),
    .DIN_SRAM19(Tile_X5Y2_DIN_SRAM19),
    .DIN_SRAM2(Tile_X5Y2_DIN_SRAM2),
    .DIN_SRAM20(Tile_X5Y2_DIN_SRAM20),
    .DIN_SRAM21(Tile_X5Y2_DIN_SRAM21),
    .DIN_SRAM22(Tile_X5Y2_DIN_SRAM22),
    .DIN_SRAM23(Tile_X5Y2_DIN_SRAM23),
    .DIN_SRAM24(Tile_X5Y2_DIN_SRAM24),
    .DIN_SRAM25(Tile_X5Y2_DIN_SRAM25),
    .DIN_SRAM26(Tile_X5Y2_DIN_SRAM26),
    .DIN_SRAM27(Tile_X5Y2_DIN_SRAM27),
    .DIN_SRAM28(Tile_X5Y2_DIN_SRAM28),
    .DIN_SRAM29(Tile_X5Y2_DIN_SRAM29),
    .DIN_SRAM3(Tile_X5Y2_DIN_SRAM3),
    .DIN_SRAM30(Tile_X5Y2_DIN_SRAM30),
    .DIN_SRAM31(Tile_X5Y2_DIN_SRAM31),
    .DIN_SRAM4(Tile_X5Y2_DIN_SRAM4),
    .DIN_SRAM5(Tile_X5Y2_DIN_SRAM5),
    .DIN_SRAM6(Tile_X5Y2_DIN_SRAM6),
    .DIN_SRAM7(Tile_X5Y2_DIN_SRAM7),
    .DIN_SRAM8(Tile_X5Y2_DIN_SRAM8),
    .DIN_SRAM9(Tile_X5Y2_DIN_SRAM9),
    .DOUT_SRAM0(Tile_X5Y2_DOUT_SRAM0),
    .DOUT_SRAM1(Tile_X5Y2_DOUT_SRAM1),
    .DOUT_SRAM10(Tile_X5Y2_DOUT_SRAM10),
    .DOUT_SRAM11(Tile_X5Y2_DOUT_SRAM11),
    .DOUT_SRAM12(Tile_X5Y2_DOUT_SRAM12),
    .DOUT_SRAM13(Tile_X5Y2_DOUT_SRAM13),
    .DOUT_SRAM14(Tile_X5Y2_DOUT_SRAM14),
    .DOUT_SRAM15(Tile_X5Y2_DOUT_SRAM15),
    .DOUT_SRAM16(Tile_X5Y2_DOUT_SRAM16),
    .DOUT_SRAM17(Tile_X5Y2_DOUT_SRAM17),
    .DOUT_SRAM18(Tile_X5Y2_DOUT_SRAM18),
    .DOUT_SRAM19(Tile_X5Y2_DOUT_SRAM19),
    .DOUT_SRAM2(Tile_X5Y2_DOUT_SRAM2),
    .DOUT_SRAM20(Tile_X5Y2_DOUT_SRAM20),
    .DOUT_SRAM21(Tile_X5Y2_DOUT_SRAM21),
    .DOUT_SRAM22(Tile_X5Y2_DOUT_SRAM22),
    .DOUT_SRAM23(Tile_X5Y2_DOUT_SRAM23),
    .DOUT_SRAM24(Tile_X5Y2_DOUT_SRAM24),
    .DOUT_SRAM25(Tile_X5Y2_DOUT_SRAM25),
    .DOUT_SRAM26(Tile_X5Y2_DOUT_SRAM26),
    .DOUT_SRAM27(Tile_X5Y2_DOUT_SRAM27),
    .DOUT_SRAM28(Tile_X5Y2_DOUT_SRAM28),
    .DOUT_SRAM29(Tile_X5Y2_DOUT_SRAM29),
    .DOUT_SRAM3(Tile_X5Y2_DOUT_SRAM3),
    .DOUT_SRAM30(Tile_X5Y2_DOUT_SRAM30),
    .DOUT_SRAM31(Tile_X5Y2_DOUT_SRAM31),
    .DOUT_SRAM4(Tile_X5Y2_DOUT_SRAM4),
    .DOUT_SRAM5(Tile_X5Y2_DOUT_SRAM5),
    .DOUT_SRAM6(Tile_X5Y2_DOUT_SRAM6),
    .DOUT_SRAM7(Tile_X5Y2_DOUT_SRAM7),
    .DOUT_SRAM8(Tile_X5Y2_DOUT_SRAM8),
    .DOUT_SRAM9(Tile_X5Y2_DOUT_SRAM9),
    .MEN_SRAM(Tile_X5Y2_MEN_SRAM),
    .REN_SRAM(Tile_X5Y2_REN_SRAM),
    .TIE_HIGH_SRAM(Tile_X5Y2_TIE_HIGH_SRAM),
    .TIE_LOW_SRAM(Tile_X5Y2_TIE_LOW_SRAM),
    .Tile_X0Y0_UserCLKo(Tile_X5Y1_UserCLKo),
    .Tile_X0Y1_UserCLK(Tile_X5Y3_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .WEN_SRAM(Tile_X5Y2_WEN_SRAM),
    .Tile_X0Y0_E1END({\Tile_X4Y1_E1BEG[3] ,
    \Tile_X4Y1_E1BEG[2] ,
    \Tile_X4Y1_E1BEG[1] ,
    \Tile_X4Y1_E1BEG[0] }),
    .Tile_X0Y0_E2END({\Tile_X4Y1_E2BEGb[7] ,
    \Tile_X4Y1_E2BEGb[6] ,
    \Tile_X4Y1_E2BEGb[5] ,
    \Tile_X4Y1_E2BEGb[4] ,
    \Tile_X4Y1_E2BEGb[3] ,
    \Tile_X4Y1_E2BEGb[2] ,
    \Tile_X4Y1_E2BEGb[1] ,
    \Tile_X4Y1_E2BEGb[0] }),
    .Tile_X0Y0_E2MID({\Tile_X4Y1_E2BEG[7] ,
    \Tile_X4Y1_E2BEG[6] ,
    \Tile_X4Y1_E2BEG[5] ,
    \Tile_X4Y1_E2BEG[4] ,
    \Tile_X4Y1_E2BEG[3] ,
    \Tile_X4Y1_E2BEG[2] ,
    \Tile_X4Y1_E2BEG[1] ,
    \Tile_X4Y1_E2BEG[0] }),
    .Tile_X0Y0_E6END({\Tile_X4Y1_E6BEG[11] ,
    \Tile_X4Y1_E6BEG[10] ,
    \Tile_X4Y1_E6BEG[9] ,
    \Tile_X4Y1_E6BEG[8] ,
    \Tile_X4Y1_E6BEG[7] ,
    \Tile_X4Y1_E6BEG[6] ,
    \Tile_X4Y1_E6BEG[5] ,
    \Tile_X4Y1_E6BEG[4] ,
    \Tile_X4Y1_E6BEG[3] ,
    \Tile_X4Y1_E6BEG[2] ,
    \Tile_X4Y1_E6BEG[1] ,
    \Tile_X4Y1_E6BEG[0] }),
    .Tile_X0Y0_EE4END({\Tile_X4Y1_EE4BEG[15] ,
    \Tile_X4Y1_EE4BEG[14] ,
    \Tile_X4Y1_EE4BEG[13] ,
    \Tile_X4Y1_EE4BEG[12] ,
    \Tile_X4Y1_EE4BEG[11] ,
    \Tile_X4Y1_EE4BEG[10] ,
    \Tile_X4Y1_EE4BEG[9] ,
    \Tile_X4Y1_EE4BEG[8] ,
    \Tile_X4Y1_EE4BEG[7] ,
    \Tile_X4Y1_EE4BEG[6] ,
    \Tile_X4Y1_EE4BEG[5] ,
    \Tile_X4Y1_EE4BEG[4] ,
    \Tile_X4Y1_EE4BEG[3] ,
    \Tile_X4Y1_EE4BEG[2] ,
    \Tile_X4Y1_EE4BEG[1] ,
    \Tile_X4Y1_EE4BEG[0] }),
    .Tile_X0Y0_FrameData({\Tile_X4Y1_FrameData_O[31] ,
    \Tile_X4Y1_FrameData_O[30] ,
    \Tile_X4Y1_FrameData_O[29] ,
    \Tile_X4Y1_FrameData_O[28] ,
    \Tile_X4Y1_FrameData_O[27] ,
    \Tile_X4Y1_FrameData_O[26] ,
    \Tile_X4Y1_FrameData_O[25] ,
    \Tile_X4Y1_FrameData_O[24] ,
    \Tile_X4Y1_FrameData_O[23] ,
    \Tile_X4Y1_FrameData_O[22] ,
    \Tile_X4Y1_FrameData_O[21] ,
    \Tile_X4Y1_FrameData_O[20] ,
    \Tile_X4Y1_FrameData_O[19] ,
    \Tile_X4Y1_FrameData_O[18] ,
    \Tile_X4Y1_FrameData_O[17] ,
    \Tile_X4Y1_FrameData_O[16] ,
    \Tile_X4Y1_FrameData_O[15] ,
    \Tile_X4Y1_FrameData_O[14] ,
    \Tile_X4Y1_FrameData_O[13] ,
    \Tile_X4Y1_FrameData_O[12] ,
    \Tile_X4Y1_FrameData_O[11] ,
    \Tile_X4Y1_FrameData_O[10] ,
    \Tile_X4Y1_FrameData_O[9] ,
    \Tile_X4Y1_FrameData_O[8] ,
    \Tile_X4Y1_FrameData_O[7] ,
    \Tile_X4Y1_FrameData_O[6] ,
    \Tile_X4Y1_FrameData_O[5] ,
    \Tile_X4Y1_FrameData_O[4] ,
    \Tile_X4Y1_FrameData_O[3] ,
    \Tile_X4Y1_FrameData_O[2] ,
    \Tile_X4Y1_FrameData_O[1] ,
    \Tile_X4Y1_FrameData_O[0] }),
    .Tile_X0Y0_FrameData_O({\Tile_X5Y1_FrameData_O[31] ,
    \Tile_X5Y1_FrameData_O[30] ,
    \Tile_X5Y1_FrameData_O[29] ,
    \Tile_X5Y1_FrameData_O[28] ,
    \Tile_X5Y1_FrameData_O[27] ,
    \Tile_X5Y1_FrameData_O[26] ,
    \Tile_X5Y1_FrameData_O[25] ,
    \Tile_X5Y1_FrameData_O[24] ,
    \Tile_X5Y1_FrameData_O[23] ,
    \Tile_X5Y1_FrameData_O[22] ,
    \Tile_X5Y1_FrameData_O[21] ,
    \Tile_X5Y1_FrameData_O[20] ,
    \Tile_X5Y1_FrameData_O[19] ,
    \Tile_X5Y1_FrameData_O[18] ,
    \Tile_X5Y1_FrameData_O[17] ,
    \Tile_X5Y1_FrameData_O[16] ,
    \Tile_X5Y1_FrameData_O[15] ,
    \Tile_X5Y1_FrameData_O[14] ,
    \Tile_X5Y1_FrameData_O[13] ,
    \Tile_X5Y1_FrameData_O[12] ,
    \Tile_X5Y1_FrameData_O[11] ,
    \Tile_X5Y1_FrameData_O[10] ,
    \Tile_X5Y1_FrameData_O[9] ,
    \Tile_X5Y1_FrameData_O[8] ,
    \Tile_X5Y1_FrameData_O[7] ,
    \Tile_X5Y1_FrameData_O[6] ,
    \Tile_X5Y1_FrameData_O[5] ,
    \Tile_X5Y1_FrameData_O[4] ,
    \Tile_X5Y1_FrameData_O[3] ,
    \Tile_X5Y1_FrameData_O[2] ,
    \Tile_X5Y1_FrameData_O[1] ,
    \Tile_X5Y1_FrameData_O[0] }),
    .Tile_X0Y0_FrameStrobe_O({\Tile_X5Y1_FrameStrobe_O[19] ,
    \Tile_X5Y1_FrameStrobe_O[18] ,
    \Tile_X5Y1_FrameStrobe_O[17] ,
    \Tile_X5Y1_FrameStrobe_O[16] ,
    \Tile_X5Y1_FrameStrobe_O[15] ,
    \Tile_X5Y1_FrameStrobe_O[14] ,
    \Tile_X5Y1_FrameStrobe_O[13] ,
    \Tile_X5Y1_FrameStrobe_O[12] ,
    \Tile_X5Y1_FrameStrobe_O[11] ,
    \Tile_X5Y1_FrameStrobe_O[10] ,
    \Tile_X5Y1_FrameStrobe_O[9] ,
    \Tile_X5Y1_FrameStrobe_O[8] ,
    \Tile_X5Y1_FrameStrobe_O[7] ,
    \Tile_X5Y1_FrameStrobe_O[6] ,
    \Tile_X5Y1_FrameStrobe_O[5] ,
    \Tile_X5Y1_FrameStrobe_O[4] ,
    \Tile_X5Y1_FrameStrobe_O[3] ,
    \Tile_X5Y1_FrameStrobe_O[2] ,
    \Tile_X5Y1_FrameStrobe_O[1] ,
    \Tile_X5Y1_FrameStrobe_O[0] }),
    .Tile_X0Y0_N1BEG({\Tile_X5Y1_N1BEG[3] ,
    \Tile_X5Y1_N1BEG[2] ,
    \Tile_X5Y1_N1BEG[1] ,
    \Tile_X5Y1_N1BEG[0] }),
    .Tile_X0Y0_N2BEG({\Tile_X5Y1_N2BEG[7] ,
    \Tile_X5Y1_N2BEG[6] ,
    \Tile_X5Y1_N2BEG[5] ,
    \Tile_X5Y1_N2BEG[4] ,
    \Tile_X5Y1_N2BEG[3] ,
    \Tile_X5Y1_N2BEG[2] ,
    \Tile_X5Y1_N2BEG[1] ,
    \Tile_X5Y1_N2BEG[0] }),
    .Tile_X0Y0_N2BEGb({\Tile_X5Y1_N2BEGb[7] ,
    \Tile_X5Y1_N2BEGb[6] ,
    \Tile_X5Y1_N2BEGb[5] ,
    \Tile_X5Y1_N2BEGb[4] ,
    \Tile_X5Y1_N2BEGb[3] ,
    \Tile_X5Y1_N2BEGb[2] ,
    \Tile_X5Y1_N2BEGb[1] ,
    \Tile_X5Y1_N2BEGb[0] }),
    .Tile_X0Y0_N4BEG({\Tile_X5Y1_N4BEG[15] ,
    \Tile_X5Y1_N4BEG[14] ,
    \Tile_X5Y1_N4BEG[13] ,
    \Tile_X5Y1_N4BEG[12] ,
    \Tile_X5Y1_N4BEG[11] ,
    \Tile_X5Y1_N4BEG[10] ,
    \Tile_X5Y1_N4BEG[9] ,
    \Tile_X5Y1_N4BEG[8] ,
    \Tile_X5Y1_N4BEG[7] ,
    \Tile_X5Y1_N4BEG[6] ,
    \Tile_X5Y1_N4BEG[5] ,
    \Tile_X5Y1_N4BEG[4] ,
    \Tile_X5Y1_N4BEG[3] ,
    \Tile_X5Y1_N4BEG[2] ,
    \Tile_X5Y1_N4BEG[1] ,
    \Tile_X5Y1_N4BEG[0] }),
    .Tile_X0Y0_S1END({\Tile_X5Y0_S1BEG[3] ,
    \Tile_X5Y0_S1BEG[2] ,
    \Tile_X5Y0_S1BEG[1] ,
    \Tile_X5Y0_S1BEG[0] }),
    .Tile_X0Y0_S2END({\Tile_X5Y0_S2BEGb[7] ,
    \Tile_X5Y0_S2BEGb[6] ,
    \Tile_X5Y0_S2BEGb[5] ,
    \Tile_X5Y0_S2BEGb[4] ,
    \Tile_X5Y0_S2BEGb[3] ,
    \Tile_X5Y0_S2BEGb[2] ,
    \Tile_X5Y0_S2BEGb[1] ,
    \Tile_X5Y0_S2BEGb[0] }),
    .Tile_X0Y0_S2MID({\Tile_X5Y0_S2BEG[7] ,
    \Tile_X5Y0_S2BEG[6] ,
    \Tile_X5Y0_S2BEG[5] ,
    \Tile_X5Y0_S2BEG[4] ,
    \Tile_X5Y0_S2BEG[3] ,
    \Tile_X5Y0_S2BEG[2] ,
    \Tile_X5Y0_S2BEG[1] ,
    \Tile_X5Y0_S2BEG[0] }),
    .Tile_X0Y0_S4END({\Tile_X5Y0_S4BEG[15] ,
    \Tile_X5Y0_S4BEG[14] ,
    \Tile_X5Y0_S4BEG[13] ,
    \Tile_X5Y0_S4BEG[12] ,
    \Tile_X5Y0_S4BEG[11] ,
    \Tile_X5Y0_S4BEG[10] ,
    \Tile_X5Y0_S4BEG[9] ,
    \Tile_X5Y0_S4BEG[8] ,
    \Tile_X5Y0_S4BEG[7] ,
    \Tile_X5Y0_S4BEG[6] ,
    \Tile_X5Y0_S4BEG[5] ,
    \Tile_X5Y0_S4BEG[4] ,
    \Tile_X5Y0_S4BEG[3] ,
    \Tile_X5Y0_S4BEG[2] ,
    \Tile_X5Y0_S4BEG[1] ,
    \Tile_X5Y0_S4BEG[0] }),
    .Tile_X0Y0_W1BEG({\Tile_X5Y1_W1BEG[3] ,
    \Tile_X5Y1_W1BEG[2] ,
    \Tile_X5Y1_W1BEG[1] ,
    \Tile_X5Y1_W1BEG[0] }),
    .Tile_X0Y0_W2BEG({\Tile_X5Y1_W2BEG[7] ,
    \Tile_X5Y1_W2BEG[6] ,
    \Tile_X5Y1_W2BEG[5] ,
    \Tile_X5Y1_W2BEG[4] ,
    \Tile_X5Y1_W2BEG[3] ,
    \Tile_X5Y1_W2BEG[2] ,
    \Tile_X5Y1_W2BEG[1] ,
    \Tile_X5Y1_W2BEG[0] }),
    .Tile_X0Y0_W2BEGb({\Tile_X5Y1_W2BEGb[7] ,
    \Tile_X5Y1_W2BEGb[6] ,
    \Tile_X5Y1_W2BEGb[5] ,
    \Tile_X5Y1_W2BEGb[4] ,
    \Tile_X5Y1_W2BEGb[3] ,
    \Tile_X5Y1_W2BEGb[2] ,
    \Tile_X5Y1_W2BEGb[1] ,
    \Tile_X5Y1_W2BEGb[0] }),
    .Tile_X0Y0_W6BEG({\Tile_X5Y1_W6BEG[11] ,
    \Tile_X5Y1_W6BEG[10] ,
    \Tile_X5Y1_W6BEG[9] ,
    \Tile_X5Y1_W6BEG[8] ,
    \Tile_X5Y1_W6BEG[7] ,
    \Tile_X5Y1_W6BEG[6] ,
    \Tile_X5Y1_W6BEG[5] ,
    \Tile_X5Y1_W6BEG[4] ,
    \Tile_X5Y1_W6BEG[3] ,
    \Tile_X5Y1_W6BEG[2] ,
    \Tile_X5Y1_W6BEG[1] ,
    \Tile_X5Y1_W6BEG[0] }),
    .Tile_X0Y0_WW4BEG({\Tile_X5Y1_WW4BEG[15] ,
    \Tile_X5Y1_WW4BEG[14] ,
    \Tile_X5Y1_WW4BEG[13] ,
    \Tile_X5Y1_WW4BEG[12] ,
    \Tile_X5Y1_WW4BEG[11] ,
    \Tile_X5Y1_WW4BEG[10] ,
    \Tile_X5Y1_WW4BEG[9] ,
    \Tile_X5Y1_WW4BEG[8] ,
    \Tile_X5Y1_WW4BEG[7] ,
    \Tile_X5Y1_WW4BEG[6] ,
    \Tile_X5Y1_WW4BEG[5] ,
    \Tile_X5Y1_WW4BEG[4] ,
    \Tile_X5Y1_WW4BEG[3] ,
    \Tile_X5Y1_WW4BEG[2] ,
    \Tile_X5Y1_WW4BEG[1] ,
    \Tile_X5Y1_WW4BEG[0] }),
    .Tile_X0Y1_E1END({\Tile_X4Y2_E1BEG[3] ,
    \Tile_X4Y2_E1BEG[2] ,
    \Tile_X4Y2_E1BEG[1] ,
    \Tile_X4Y2_E1BEG[0] }),
    .Tile_X0Y1_E2END({\Tile_X4Y2_E2BEGb[7] ,
    \Tile_X4Y2_E2BEGb[6] ,
    \Tile_X4Y2_E2BEGb[5] ,
    \Tile_X4Y2_E2BEGb[4] ,
    \Tile_X4Y2_E2BEGb[3] ,
    \Tile_X4Y2_E2BEGb[2] ,
    \Tile_X4Y2_E2BEGb[1] ,
    \Tile_X4Y2_E2BEGb[0] }),
    .Tile_X0Y1_E2MID({\Tile_X4Y2_E2BEG[7] ,
    \Tile_X4Y2_E2BEG[6] ,
    \Tile_X4Y2_E2BEG[5] ,
    \Tile_X4Y2_E2BEG[4] ,
    \Tile_X4Y2_E2BEG[3] ,
    \Tile_X4Y2_E2BEG[2] ,
    \Tile_X4Y2_E2BEG[1] ,
    \Tile_X4Y2_E2BEG[0] }),
    .Tile_X0Y1_E6END({\Tile_X4Y2_E6BEG[11] ,
    \Tile_X4Y2_E6BEG[10] ,
    \Tile_X4Y2_E6BEG[9] ,
    \Tile_X4Y2_E6BEG[8] ,
    \Tile_X4Y2_E6BEG[7] ,
    \Tile_X4Y2_E6BEG[6] ,
    \Tile_X4Y2_E6BEG[5] ,
    \Tile_X4Y2_E6BEG[4] ,
    \Tile_X4Y2_E6BEG[3] ,
    \Tile_X4Y2_E6BEG[2] ,
    \Tile_X4Y2_E6BEG[1] ,
    \Tile_X4Y2_E6BEG[0] }),
    .Tile_X0Y1_EE4END({\Tile_X4Y2_EE4BEG[15] ,
    \Tile_X4Y2_EE4BEG[14] ,
    \Tile_X4Y2_EE4BEG[13] ,
    \Tile_X4Y2_EE4BEG[12] ,
    \Tile_X4Y2_EE4BEG[11] ,
    \Tile_X4Y2_EE4BEG[10] ,
    \Tile_X4Y2_EE4BEG[9] ,
    \Tile_X4Y2_EE4BEG[8] ,
    \Tile_X4Y2_EE4BEG[7] ,
    \Tile_X4Y2_EE4BEG[6] ,
    \Tile_X4Y2_EE4BEG[5] ,
    \Tile_X4Y2_EE4BEG[4] ,
    \Tile_X4Y2_EE4BEG[3] ,
    \Tile_X4Y2_EE4BEG[2] ,
    \Tile_X4Y2_EE4BEG[1] ,
    \Tile_X4Y2_EE4BEG[0] }),
    .Tile_X0Y1_FrameData({\Tile_X4Y2_FrameData_O[31] ,
    \Tile_X4Y2_FrameData_O[30] ,
    \Tile_X4Y2_FrameData_O[29] ,
    \Tile_X4Y2_FrameData_O[28] ,
    \Tile_X4Y2_FrameData_O[27] ,
    \Tile_X4Y2_FrameData_O[26] ,
    \Tile_X4Y2_FrameData_O[25] ,
    \Tile_X4Y2_FrameData_O[24] ,
    \Tile_X4Y2_FrameData_O[23] ,
    \Tile_X4Y2_FrameData_O[22] ,
    \Tile_X4Y2_FrameData_O[21] ,
    \Tile_X4Y2_FrameData_O[20] ,
    \Tile_X4Y2_FrameData_O[19] ,
    \Tile_X4Y2_FrameData_O[18] ,
    \Tile_X4Y2_FrameData_O[17] ,
    \Tile_X4Y2_FrameData_O[16] ,
    \Tile_X4Y2_FrameData_O[15] ,
    \Tile_X4Y2_FrameData_O[14] ,
    \Tile_X4Y2_FrameData_O[13] ,
    \Tile_X4Y2_FrameData_O[12] ,
    \Tile_X4Y2_FrameData_O[11] ,
    \Tile_X4Y2_FrameData_O[10] ,
    \Tile_X4Y2_FrameData_O[9] ,
    \Tile_X4Y2_FrameData_O[8] ,
    \Tile_X4Y2_FrameData_O[7] ,
    \Tile_X4Y2_FrameData_O[6] ,
    \Tile_X4Y2_FrameData_O[5] ,
    \Tile_X4Y2_FrameData_O[4] ,
    \Tile_X4Y2_FrameData_O[3] ,
    \Tile_X4Y2_FrameData_O[2] ,
    \Tile_X4Y2_FrameData_O[1] ,
    \Tile_X4Y2_FrameData_O[0] }),
    .Tile_X0Y1_FrameData_O({\Tile_X5Y2_FrameData_O[31] ,
    \Tile_X5Y2_FrameData_O[30] ,
    \Tile_X5Y2_FrameData_O[29] ,
    \Tile_X5Y2_FrameData_O[28] ,
    \Tile_X5Y2_FrameData_O[27] ,
    \Tile_X5Y2_FrameData_O[26] ,
    \Tile_X5Y2_FrameData_O[25] ,
    \Tile_X5Y2_FrameData_O[24] ,
    \Tile_X5Y2_FrameData_O[23] ,
    \Tile_X5Y2_FrameData_O[22] ,
    \Tile_X5Y2_FrameData_O[21] ,
    \Tile_X5Y2_FrameData_O[20] ,
    \Tile_X5Y2_FrameData_O[19] ,
    \Tile_X5Y2_FrameData_O[18] ,
    \Tile_X5Y2_FrameData_O[17] ,
    \Tile_X5Y2_FrameData_O[16] ,
    \Tile_X5Y2_FrameData_O[15] ,
    \Tile_X5Y2_FrameData_O[14] ,
    \Tile_X5Y2_FrameData_O[13] ,
    \Tile_X5Y2_FrameData_O[12] ,
    \Tile_X5Y2_FrameData_O[11] ,
    \Tile_X5Y2_FrameData_O[10] ,
    \Tile_X5Y2_FrameData_O[9] ,
    \Tile_X5Y2_FrameData_O[8] ,
    \Tile_X5Y2_FrameData_O[7] ,
    \Tile_X5Y2_FrameData_O[6] ,
    \Tile_X5Y2_FrameData_O[5] ,
    \Tile_X5Y2_FrameData_O[4] ,
    \Tile_X5Y2_FrameData_O[3] ,
    \Tile_X5Y2_FrameData_O[2] ,
    \Tile_X5Y2_FrameData_O[1] ,
    \Tile_X5Y2_FrameData_O[0] }),
    .Tile_X0Y1_FrameStrobe({\Tile_X5Y3_FrameStrobe_O[19] ,
    \Tile_X5Y3_FrameStrobe_O[18] ,
    \Tile_X5Y3_FrameStrobe_O[17] ,
    \Tile_X5Y3_FrameStrobe_O[16] ,
    \Tile_X5Y3_FrameStrobe_O[15] ,
    \Tile_X5Y3_FrameStrobe_O[14] ,
    \Tile_X5Y3_FrameStrobe_O[13] ,
    \Tile_X5Y3_FrameStrobe_O[12] ,
    \Tile_X5Y3_FrameStrobe_O[11] ,
    \Tile_X5Y3_FrameStrobe_O[10] ,
    \Tile_X5Y3_FrameStrobe_O[9] ,
    \Tile_X5Y3_FrameStrobe_O[8] ,
    \Tile_X5Y3_FrameStrobe_O[7] ,
    \Tile_X5Y3_FrameStrobe_O[6] ,
    \Tile_X5Y3_FrameStrobe_O[5] ,
    \Tile_X5Y3_FrameStrobe_O[4] ,
    \Tile_X5Y3_FrameStrobe_O[3] ,
    \Tile_X5Y3_FrameStrobe_O[2] ,
    \Tile_X5Y3_FrameStrobe_O[1] ,
    \Tile_X5Y3_FrameStrobe_O[0] }),
    .Tile_X0Y1_N1END({\Tile_X5Y3_N1BEG[3] ,
    \Tile_X5Y3_N1BEG[2] ,
    \Tile_X5Y3_N1BEG[1] ,
    \Tile_X5Y3_N1BEG[0] }),
    .Tile_X0Y1_N2END({\Tile_X5Y3_N2BEGb[7] ,
    \Tile_X5Y3_N2BEGb[6] ,
    \Tile_X5Y3_N2BEGb[5] ,
    \Tile_X5Y3_N2BEGb[4] ,
    \Tile_X5Y3_N2BEGb[3] ,
    \Tile_X5Y3_N2BEGb[2] ,
    \Tile_X5Y3_N2BEGb[1] ,
    \Tile_X5Y3_N2BEGb[0] }),
    .Tile_X0Y1_N2MID({\Tile_X5Y3_N2BEG[7] ,
    \Tile_X5Y3_N2BEG[6] ,
    \Tile_X5Y3_N2BEG[5] ,
    \Tile_X5Y3_N2BEG[4] ,
    \Tile_X5Y3_N2BEG[3] ,
    \Tile_X5Y3_N2BEG[2] ,
    \Tile_X5Y3_N2BEG[1] ,
    \Tile_X5Y3_N2BEG[0] }),
    .Tile_X0Y1_N4END({\Tile_X5Y3_N4BEG[15] ,
    \Tile_X5Y3_N4BEG[14] ,
    \Tile_X5Y3_N4BEG[13] ,
    \Tile_X5Y3_N4BEG[12] ,
    \Tile_X5Y3_N4BEG[11] ,
    \Tile_X5Y3_N4BEG[10] ,
    \Tile_X5Y3_N4BEG[9] ,
    \Tile_X5Y3_N4BEG[8] ,
    \Tile_X5Y3_N4BEG[7] ,
    \Tile_X5Y3_N4BEG[6] ,
    \Tile_X5Y3_N4BEG[5] ,
    \Tile_X5Y3_N4BEG[4] ,
    \Tile_X5Y3_N4BEG[3] ,
    \Tile_X5Y3_N4BEG[2] ,
    \Tile_X5Y3_N4BEG[1] ,
    \Tile_X5Y3_N4BEG[0] }),
    .Tile_X0Y1_S1BEG({\Tile_X5Y2_S1BEG[3] ,
    \Tile_X5Y2_S1BEG[2] ,
    \Tile_X5Y2_S1BEG[1] ,
    \Tile_X5Y2_S1BEG[0] }),
    .Tile_X0Y1_S2BEG({\Tile_X5Y2_S2BEG[7] ,
    \Tile_X5Y2_S2BEG[6] ,
    \Tile_X5Y2_S2BEG[5] ,
    \Tile_X5Y2_S2BEG[4] ,
    \Tile_X5Y2_S2BEG[3] ,
    \Tile_X5Y2_S2BEG[2] ,
    \Tile_X5Y2_S2BEG[1] ,
    \Tile_X5Y2_S2BEG[0] }),
    .Tile_X0Y1_S2BEGb({\Tile_X5Y2_S2BEGb[7] ,
    \Tile_X5Y2_S2BEGb[6] ,
    \Tile_X5Y2_S2BEGb[5] ,
    \Tile_X5Y2_S2BEGb[4] ,
    \Tile_X5Y2_S2BEGb[3] ,
    \Tile_X5Y2_S2BEGb[2] ,
    \Tile_X5Y2_S2BEGb[1] ,
    \Tile_X5Y2_S2BEGb[0] }),
    .Tile_X0Y1_S4BEG({\Tile_X5Y2_S4BEG[15] ,
    \Tile_X5Y2_S4BEG[14] ,
    \Tile_X5Y2_S4BEG[13] ,
    \Tile_X5Y2_S4BEG[12] ,
    \Tile_X5Y2_S4BEG[11] ,
    \Tile_X5Y2_S4BEG[10] ,
    \Tile_X5Y2_S4BEG[9] ,
    \Tile_X5Y2_S4BEG[8] ,
    \Tile_X5Y2_S4BEG[7] ,
    \Tile_X5Y2_S4BEG[6] ,
    \Tile_X5Y2_S4BEG[5] ,
    \Tile_X5Y2_S4BEG[4] ,
    \Tile_X5Y2_S4BEG[3] ,
    \Tile_X5Y2_S4BEG[2] ,
    \Tile_X5Y2_S4BEG[1] ,
    \Tile_X5Y2_S4BEG[0] }),
    .Tile_X0Y1_W1BEG({\Tile_X5Y2_W1BEG[3] ,
    \Tile_X5Y2_W1BEG[2] ,
    \Tile_X5Y2_W1BEG[1] ,
    \Tile_X5Y2_W1BEG[0] }),
    .Tile_X0Y1_W2BEG({\Tile_X5Y2_W2BEG[7] ,
    \Tile_X5Y2_W2BEG[6] ,
    \Tile_X5Y2_W2BEG[5] ,
    \Tile_X5Y2_W2BEG[4] ,
    \Tile_X5Y2_W2BEG[3] ,
    \Tile_X5Y2_W2BEG[2] ,
    \Tile_X5Y2_W2BEG[1] ,
    \Tile_X5Y2_W2BEG[0] }),
    .Tile_X0Y1_W2BEGb({\Tile_X5Y2_W2BEGb[7] ,
    \Tile_X5Y2_W2BEGb[6] ,
    \Tile_X5Y2_W2BEGb[5] ,
    \Tile_X5Y2_W2BEGb[4] ,
    \Tile_X5Y2_W2BEGb[3] ,
    \Tile_X5Y2_W2BEGb[2] ,
    \Tile_X5Y2_W2BEGb[1] ,
    \Tile_X5Y2_W2BEGb[0] }),
    .Tile_X0Y1_W6BEG({\Tile_X5Y2_W6BEG[11] ,
    \Tile_X5Y2_W6BEG[10] ,
    \Tile_X5Y2_W6BEG[9] ,
    \Tile_X5Y2_W6BEG[8] ,
    \Tile_X5Y2_W6BEG[7] ,
    \Tile_X5Y2_W6BEG[6] ,
    \Tile_X5Y2_W6BEG[5] ,
    \Tile_X5Y2_W6BEG[4] ,
    \Tile_X5Y2_W6BEG[3] ,
    \Tile_X5Y2_W6BEG[2] ,
    \Tile_X5Y2_W6BEG[1] ,
    \Tile_X5Y2_W6BEG[0] }),
    .Tile_X0Y1_WW4BEG({\Tile_X5Y2_WW4BEG[15] ,
    \Tile_X5Y2_WW4BEG[14] ,
    \Tile_X5Y2_WW4BEG[13] ,
    \Tile_X5Y2_WW4BEG[12] ,
    \Tile_X5Y2_WW4BEG[11] ,
    \Tile_X5Y2_WW4BEG[10] ,
    \Tile_X5Y2_WW4BEG[9] ,
    \Tile_X5Y2_WW4BEG[8] ,
    \Tile_X5Y2_WW4BEG[7] ,
    \Tile_X5Y2_WW4BEG[6] ,
    \Tile_X5Y2_WW4BEG[5] ,
    \Tile_X5Y2_WW4BEG[4] ,
    \Tile_X5Y2_WW4BEG[3] ,
    \Tile_X5Y2_WW4BEG[2] ,
    \Tile_X5Y2_WW4BEG[1] ,
    \Tile_X5Y2_WW4BEG[0] }));
 E_TT_IF2 Tile_X5Y3_E_TT_IF2 (.CLK_TT_PROJECT(Tile_X5Y4_CLK_TT_PROJECT),
    .ENA_TT_PROJECT(Tile_X5Y4_ENA_TT_PROJECT),
    .RST_N_TT_PROJECT(Tile_X5Y4_RST_N_TT_PROJECT),
    .Tile_X0Y0_UserCLKo(Tile_X5Y3_UserCLKo),
    .Tile_X0Y1_UserCLK(Tile_X5Y5_UserCLKo),
    .UIO_IN_TT_PROJECT0(Tile_X5Y4_UIO_IN_TT_PROJECT0),
    .UIO_IN_TT_PROJECT1(Tile_X5Y4_UIO_IN_TT_PROJECT1),
    .UIO_IN_TT_PROJECT2(Tile_X5Y4_UIO_IN_TT_PROJECT2),
    .UIO_IN_TT_PROJECT3(Tile_X5Y4_UIO_IN_TT_PROJECT3),
    .UIO_IN_TT_PROJECT4(Tile_X5Y4_UIO_IN_TT_PROJECT4),
    .UIO_IN_TT_PROJECT5(Tile_X5Y4_UIO_IN_TT_PROJECT5),
    .UIO_IN_TT_PROJECT6(Tile_X5Y4_UIO_IN_TT_PROJECT6),
    .UIO_IN_TT_PROJECT7(Tile_X5Y4_UIO_IN_TT_PROJECT7),
    .UIO_OE_TT_PROJECT0(Tile_X5Y4_UIO_OE_TT_PROJECT0),
    .UIO_OE_TT_PROJECT1(Tile_X5Y4_UIO_OE_TT_PROJECT1),
    .UIO_OE_TT_PROJECT2(Tile_X5Y4_UIO_OE_TT_PROJECT2),
    .UIO_OE_TT_PROJECT3(Tile_X5Y4_UIO_OE_TT_PROJECT3),
    .UIO_OE_TT_PROJECT4(Tile_X5Y4_UIO_OE_TT_PROJECT4),
    .UIO_OE_TT_PROJECT5(Tile_X5Y4_UIO_OE_TT_PROJECT5),
    .UIO_OE_TT_PROJECT6(Tile_X5Y4_UIO_OE_TT_PROJECT6),
    .UIO_OE_TT_PROJECT7(Tile_X5Y4_UIO_OE_TT_PROJECT7),
    .UIO_OUT_TT_PROJECT0(Tile_X5Y4_UIO_OUT_TT_PROJECT0),
    .UIO_OUT_TT_PROJECT1(Tile_X5Y4_UIO_OUT_TT_PROJECT1),
    .UIO_OUT_TT_PROJECT2(Tile_X5Y4_UIO_OUT_TT_PROJECT2),
    .UIO_OUT_TT_PROJECT3(Tile_X5Y4_UIO_OUT_TT_PROJECT3),
    .UIO_OUT_TT_PROJECT4(Tile_X5Y4_UIO_OUT_TT_PROJECT4),
    .UIO_OUT_TT_PROJECT5(Tile_X5Y4_UIO_OUT_TT_PROJECT5),
    .UIO_OUT_TT_PROJECT6(Tile_X5Y4_UIO_OUT_TT_PROJECT6),
    .UIO_OUT_TT_PROJECT7(Tile_X5Y4_UIO_OUT_TT_PROJECT7),
    .UI_IN_TT_PROJECT0(Tile_X5Y4_UI_IN_TT_PROJECT0),
    .UI_IN_TT_PROJECT1(Tile_X5Y4_UI_IN_TT_PROJECT1),
    .UI_IN_TT_PROJECT2(Tile_X5Y4_UI_IN_TT_PROJECT2),
    .UI_IN_TT_PROJECT3(Tile_X5Y4_UI_IN_TT_PROJECT3),
    .UI_IN_TT_PROJECT4(Tile_X5Y4_UI_IN_TT_PROJECT4),
    .UI_IN_TT_PROJECT5(Tile_X5Y4_UI_IN_TT_PROJECT5),
    .UI_IN_TT_PROJECT6(Tile_X5Y4_UI_IN_TT_PROJECT6),
    .UI_IN_TT_PROJECT7(Tile_X5Y4_UI_IN_TT_PROJECT7),
    .UO_OUT_TT_PROJECT0(Tile_X5Y4_UO_OUT_TT_PROJECT0),
    .UO_OUT_TT_PROJECT1(Tile_X5Y4_UO_OUT_TT_PROJECT1),
    .UO_OUT_TT_PROJECT2(Tile_X5Y4_UO_OUT_TT_PROJECT2),
    .UO_OUT_TT_PROJECT3(Tile_X5Y4_UO_OUT_TT_PROJECT3),
    .UO_OUT_TT_PROJECT4(Tile_X5Y4_UO_OUT_TT_PROJECT4),
    .UO_OUT_TT_PROJECT5(Tile_X5Y4_UO_OUT_TT_PROJECT5),
    .UO_OUT_TT_PROJECT6(Tile_X5Y4_UO_OUT_TT_PROJECT6),
    .UO_OUT_TT_PROJECT7(Tile_X5Y4_UO_OUT_TT_PROJECT7),
    .VGND(VGND),
    .VPWR(VPWR),
    .Tile_X0Y0_E1END({\Tile_X4Y3_E1BEG[3] ,
    \Tile_X4Y3_E1BEG[2] ,
    \Tile_X4Y3_E1BEG[1] ,
    \Tile_X4Y3_E1BEG[0] }),
    .Tile_X0Y0_E2END({\Tile_X4Y3_E2BEGb[7] ,
    \Tile_X4Y3_E2BEGb[6] ,
    \Tile_X4Y3_E2BEGb[5] ,
    \Tile_X4Y3_E2BEGb[4] ,
    \Tile_X4Y3_E2BEGb[3] ,
    \Tile_X4Y3_E2BEGb[2] ,
    \Tile_X4Y3_E2BEGb[1] ,
    \Tile_X4Y3_E2BEGb[0] }),
    .Tile_X0Y0_E2MID({\Tile_X4Y3_E2BEG[7] ,
    \Tile_X4Y3_E2BEG[6] ,
    \Tile_X4Y3_E2BEG[5] ,
    \Tile_X4Y3_E2BEG[4] ,
    \Tile_X4Y3_E2BEG[3] ,
    \Tile_X4Y3_E2BEG[2] ,
    \Tile_X4Y3_E2BEG[1] ,
    \Tile_X4Y3_E2BEG[0] }),
    .Tile_X0Y0_E6END({\Tile_X4Y3_E6BEG[11] ,
    \Tile_X4Y3_E6BEG[10] ,
    \Tile_X4Y3_E6BEG[9] ,
    \Tile_X4Y3_E6BEG[8] ,
    \Tile_X4Y3_E6BEG[7] ,
    \Tile_X4Y3_E6BEG[6] ,
    \Tile_X4Y3_E6BEG[5] ,
    \Tile_X4Y3_E6BEG[4] ,
    \Tile_X4Y3_E6BEG[3] ,
    \Tile_X4Y3_E6BEG[2] ,
    \Tile_X4Y3_E6BEG[1] ,
    \Tile_X4Y3_E6BEG[0] }),
    .Tile_X0Y0_EE4END({\Tile_X4Y3_EE4BEG[15] ,
    \Tile_X4Y3_EE4BEG[14] ,
    \Tile_X4Y3_EE4BEG[13] ,
    \Tile_X4Y3_EE4BEG[12] ,
    \Tile_X4Y3_EE4BEG[11] ,
    \Tile_X4Y3_EE4BEG[10] ,
    \Tile_X4Y3_EE4BEG[9] ,
    \Tile_X4Y3_EE4BEG[8] ,
    \Tile_X4Y3_EE4BEG[7] ,
    \Tile_X4Y3_EE4BEG[6] ,
    \Tile_X4Y3_EE4BEG[5] ,
    \Tile_X4Y3_EE4BEG[4] ,
    \Tile_X4Y3_EE4BEG[3] ,
    \Tile_X4Y3_EE4BEG[2] ,
    \Tile_X4Y3_EE4BEG[1] ,
    \Tile_X4Y3_EE4BEG[0] }),
    .Tile_X0Y0_FrameData({\Tile_X4Y3_FrameData_O[31] ,
    \Tile_X4Y3_FrameData_O[30] ,
    \Tile_X4Y3_FrameData_O[29] ,
    \Tile_X4Y3_FrameData_O[28] ,
    \Tile_X4Y3_FrameData_O[27] ,
    \Tile_X4Y3_FrameData_O[26] ,
    \Tile_X4Y3_FrameData_O[25] ,
    \Tile_X4Y3_FrameData_O[24] ,
    \Tile_X4Y3_FrameData_O[23] ,
    \Tile_X4Y3_FrameData_O[22] ,
    \Tile_X4Y3_FrameData_O[21] ,
    \Tile_X4Y3_FrameData_O[20] ,
    \Tile_X4Y3_FrameData_O[19] ,
    \Tile_X4Y3_FrameData_O[18] ,
    \Tile_X4Y3_FrameData_O[17] ,
    \Tile_X4Y3_FrameData_O[16] ,
    \Tile_X4Y3_FrameData_O[15] ,
    \Tile_X4Y3_FrameData_O[14] ,
    \Tile_X4Y3_FrameData_O[13] ,
    \Tile_X4Y3_FrameData_O[12] ,
    \Tile_X4Y3_FrameData_O[11] ,
    \Tile_X4Y3_FrameData_O[10] ,
    \Tile_X4Y3_FrameData_O[9] ,
    \Tile_X4Y3_FrameData_O[8] ,
    \Tile_X4Y3_FrameData_O[7] ,
    \Tile_X4Y3_FrameData_O[6] ,
    \Tile_X4Y3_FrameData_O[5] ,
    \Tile_X4Y3_FrameData_O[4] ,
    \Tile_X4Y3_FrameData_O[3] ,
    \Tile_X4Y3_FrameData_O[2] ,
    \Tile_X4Y3_FrameData_O[1] ,
    \Tile_X4Y3_FrameData_O[0] }),
    .Tile_X0Y0_FrameData_O({\Tile_X5Y3_FrameData_O[31] ,
    \Tile_X5Y3_FrameData_O[30] ,
    \Tile_X5Y3_FrameData_O[29] ,
    \Tile_X5Y3_FrameData_O[28] ,
    \Tile_X5Y3_FrameData_O[27] ,
    \Tile_X5Y3_FrameData_O[26] ,
    \Tile_X5Y3_FrameData_O[25] ,
    \Tile_X5Y3_FrameData_O[24] ,
    \Tile_X5Y3_FrameData_O[23] ,
    \Tile_X5Y3_FrameData_O[22] ,
    \Tile_X5Y3_FrameData_O[21] ,
    \Tile_X5Y3_FrameData_O[20] ,
    \Tile_X5Y3_FrameData_O[19] ,
    \Tile_X5Y3_FrameData_O[18] ,
    \Tile_X5Y3_FrameData_O[17] ,
    \Tile_X5Y3_FrameData_O[16] ,
    \Tile_X5Y3_FrameData_O[15] ,
    \Tile_X5Y3_FrameData_O[14] ,
    \Tile_X5Y3_FrameData_O[13] ,
    \Tile_X5Y3_FrameData_O[12] ,
    \Tile_X5Y3_FrameData_O[11] ,
    \Tile_X5Y3_FrameData_O[10] ,
    \Tile_X5Y3_FrameData_O[9] ,
    \Tile_X5Y3_FrameData_O[8] ,
    \Tile_X5Y3_FrameData_O[7] ,
    \Tile_X5Y3_FrameData_O[6] ,
    \Tile_X5Y3_FrameData_O[5] ,
    \Tile_X5Y3_FrameData_O[4] ,
    \Tile_X5Y3_FrameData_O[3] ,
    \Tile_X5Y3_FrameData_O[2] ,
    \Tile_X5Y3_FrameData_O[1] ,
    \Tile_X5Y3_FrameData_O[0] }),
    .Tile_X0Y0_FrameStrobe_O({\Tile_X5Y3_FrameStrobe_O[19] ,
    \Tile_X5Y3_FrameStrobe_O[18] ,
    \Tile_X5Y3_FrameStrobe_O[17] ,
    \Tile_X5Y3_FrameStrobe_O[16] ,
    \Tile_X5Y3_FrameStrobe_O[15] ,
    \Tile_X5Y3_FrameStrobe_O[14] ,
    \Tile_X5Y3_FrameStrobe_O[13] ,
    \Tile_X5Y3_FrameStrobe_O[12] ,
    \Tile_X5Y3_FrameStrobe_O[11] ,
    \Tile_X5Y3_FrameStrobe_O[10] ,
    \Tile_X5Y3_FrameStrobe_O[9] ,
    \Tile_X5Y3_FrameStrobe_O[8] ,
    \Tile_X5Y3_FrameStrobe_O[7] ,
    \Tile_X5Y3_FrameStrobe_O[6] ,
    \Tile_X5Y3_FrameStrobe_O[5] ,
    \Tile_X5Y3_FrameStrobe_O[4] ,
    \Tile_X5Y3_FrameStrobe_O[3] ,
    \Tile_X5Y3_FrameStrobe_O[2] ,
    \Tile_X5Y3_FrameStrobe_O[1] ,
    \Tile_X5Y3_FrameStrobe_O[0] }),
    .Tile_X0Y0_N1BEG({\Tile_X5Y3_N1BEG[3] ,
    \Tile_X5Y3_N1BEG[2] ,
    \Tile_X5Y3_N1BEG[1] ,
    \Tile_X5Y3_N1BEG[0] }),
    .Tile_X0Y0_N2BEG({\Tile_X5Y3_N2BEG[7] ,
    \Tile_X5Y3_N2BEG[6] ,
    \Tile_X5Y3_N2BEG[5] ,
    \Tile_X5Y3_N2BEG[4] ,
    \Tile_X5Y3_N2BEG[3] ,
    \Tile_X5Y3_N2BEG[2] ,
    \Tile_X5Y3_N2BEG[1] ,
    \Tile_X5Y3_N2BEG[0] }),
    .Tile_X0Y0_N2BEGb({\Tile_X5Y3_N2BEGb[7] ,
    \Tile_X5Y3_N2BEGb[6] ,
    \Tile_X5Y3_N2BEGb[5] ,
    \Tile_X5Y3_N2BEGb[4] ,
    \Tile_X5Y3_N2BEGb[3] ,
    \Tile_X5Y3_N2BEGb[2] ,
    \Tile_X5Y3_N2BEGb[1] ,
    \Tile_X5Y3_N2BEGb[0] }),
    .Tile_X0Y0_N4BEG({\Tile_X5Y3_N4BEG[15] ,
    \Tile_X5Y3_N4BEG[14] ,
    \Tile_X5Y3_N4BEG[13] ,
    \Tile_X5Y3_N4BEG[12] ,
    \Tile_X5Y3_N4BEG[11] ,
    \Tile_X5Y3_N4BEG[10] ,
    \Tile_X5Y3_N4BEG[9] ,
    \Tile_X5Y3_N4BEG[8] ,
    \Tile_X5Y3_N4BEG[7] ,
    \Tile_X5Y3_N4BEG[6] ,
    \Tile_X5Y3_N4BEG[5] ,
    \Tile_X5Y3_N4BEG[4] ,
    \Tile_X5Y3_N4BEG[3] ,
    \Tile_X5Y3_N4BEG[2] ,
    \Tile_X5Y3_N4BEG[1] ,
    \Tile_X5Y3_N4BEG[0] }),
    .Tile_X0Y0_S1END({\Tile_X5Y2_S1BEG[3] ,
    \Tile_X5Y2_S1BEG[2] ,
    \Tile_X5Y2_S1BEG[1] ,
    \Tile_X5Y2_S1BEG[0] }),
    .Tile_X0Y0_S2END({\Tile_X5Y2_S2BEGb[7] ,
    \Tile_X5Y2_S2BEGb[6] ,
    \Tile_X5Y2_S2BEGb[5] ,
    \Tile_X5Y2_S2BEGb[4] ,
    \Tile_X5Y2_S2BEGb[3] ,
    \Tile_X5Y2_S2BEGb[2] ,
    \Tile_X5Y2_S2BEGb[1] ,
    \Tile_X5Y2_S2BEGb[0] }),
    .Tile_X0Y0_S2MID({\Tile_X5Y2_S2BEG[7] ,
    \Tile_X5Y2_S2BEG[6] ,
    \Tile_X5Y2_S2BEG[5] ,
    \Tile_X5Y2_S2BEG[4] ,
    \Tile_X5Y2_S2BEG[3] ,
    \Tile_X5Y2_S2BEG[2] ,
    \Tile_X5Y2_S2BEG[1] ,
    \Tile_X5Y2_S2BEG[0] }),
    .Tile_X0Y0_S4END({\Tile_X5Y2_S4BEG[15] ,
    \Tile_X5Y2_S4BEG[14] ,
    \Tile_X5Y2_S4BEG[13] ,
    \Tile_X5Y2_S4BEG[12] ,
    \Tile_X5Y2_S4BEG[11] ,
    \Tile_X5Y2_S4BEG[10] ,
    \Tile_X5Y2_S4BEG[9] ,
    \Tile_X5Y2_S4BEG[8] ,
    \Tile_X5Y2_S4BEG[7] ,
    \Tile_X5Y2_S4BEG[6] ,
    \Tile_X5Y2_S4BEG[5] ,
    \Tile_X5Y2_S4BEG[4] ,
    \Tile_X5Y2_S4BEG[3] ,
    \Tile_X5Y2_S4BEG[2] ,
    \Tile_X5Y2_S4BEG[1] ,
    \Tile_X5Y2_S4BEG[0] }),
    .Tile_X0Y0_W1BEG({\Tile_X5Y3_W1BEG[3] ,
    \Tile_X5Y3_W1BEG[2] ,
    \Tile_X5Y3_W1BEG[1] ,
    \Tile_X5Y3_W1BEG[0] }),
    .Tile_X0Y0_W2BEG({\Tile_X5Y3_W2BEG[7] ,
    \Tile_X5Y3_W2BEG[6] ,
    \Tile_X5Y3_W2BEG[5] ,
    \Tile_X5Y3_W2BEG[4] ,
    \Tile_X5Y3_W2BEG[3] ,
    \Tile_X5Y3_W2BEG[2] ,
    \Tile_X5Y3_W2BEG[1] ,
    \Tile_X5Y3_W2BEG[0] }),
    .Tile_X0Y0_W2BEGb({\Tile_X5Y3_W2BEGb[7] ,
    \Tile_X5Y3_W2BEGb[6] ,
    \Tile_X5Y3_W2BEGb[5] ,
    \Tile_X5Y3_W2BEGb[4] ,
    \Tile_X5Y3_W2BEGb[3] ,
    \Tile_X5Y3_W2BEGb[2] ,
    \Tile_X5Y3_W2BEGb[1] ,
    \Tile_X5Y3_W2BEGb[0] }),
    .Tile_X0Y0_W6BEG({\Tile_X5Y3_W6BEG[11] ,
    \Tile_X5Y3_W6BEG[10] ,
    \Tile_X5Y3_W6BEG[9] ,
    \Tile_X5Y3_W6BEG[8] ,
    \Tile_X5Y3_W6BEG[7] ,
    \Tile_X5Y3_W6BEG[6] ,
    \Tile_X5Y3_W6BEG[5] ,
    \Tile_X5Y3_W6BEG[4] ,
    \Tile_X5Y3_W6BEG[3] ,
    \Tile_X5Y3_W6BEG[2] ,
    \Tile_X5Y3_W6BEG[1] ,
    \Tile_X5Y3_W6BEG[0] }),
    .Tile_X0Y0_WW4BEG({\Tile_X5Y3_WW4BEG[15] ,
    \Tile_X5Y3_WW4BEG[14] ,
    \Tile_X5Y3_WW4BEG[13] ,
    \Tile_X5Y3_WW4BEG[12] ,
    \Tile_X5Y3_WW4BEG[11] ,
    \Tile_X5Y3_WW4BEG[10] ,
    \Tile_X5Y3_WW4BEG[9] ,
    \Tile_X5Y3_WW4BEG[8] ,
    \Tile_X5Y3_WW4BEG[7] ,
    \Tile_X5Y3_WW4BEG[6] ,
    \Tile_X5Y3_WW4BEG[5] ,
    \Tile_X5Y3_WW4BEG[4] ,
    \Tile_X5Y3_WW4BEG[3] ,
    \Tile_X5Y3_WW4BEG[2] ,
    \Tile_X5Y3_WW4BEG[1] ,
    \Tile_X5Y3_WW4BEG[0] }),
    .Tile_X0Y1_E1END({\Tile_X4Y4_E1BEG[3] ,
    \Tile_X4Y4_E1BEG[2] ,
    \Tile_X4Y4_E1BEG[1] ,
    \Tile_X4Y4_E1BEG[0] }),
    .Tile_X0Y1_E2END({\Tile_X4Y4_E2BEGb[7] ,
    \Tile_X4Y4_E2BEGb[6] ,
    \Tile_X4Y4_E2BEGb[5] ,
    \Tile_X4Y4_E2BEGb[4] ,
    \Tile_X4Y4_E2BEGb[3] ,
    \Tile_X4Y4_E2BEGb[2] ,
    \Tile_X4Y4_E2BEGb[1] ,
    \Tile_X4Y4_E2BEGb[0] }),
    .Tile_X0Y1_E2MID({\Tile_X4Y4_E2BEG[7] ,
    \Tile_X4Y4_E2BEG[6] ,
    \Tile_X4Y4_E2BEG[5] ,
    \Tile_X4Y4_E2BEG[4] ,
    \Tile_X4Y4_E2BEG[3] ,
    \Tile_X4Y4_E2BEG[2] ,
    \Tile_X4Y4_E2BEG[1] ,
    \Tile_X4Y4_E2BEG[0] }),
    .Tile_X0Y1_E6END({\Tile_X4Y4_E6BEG[11] ,
    \Tile_X4Y4_E6BEG[10] ,
    \Tile_X4Y4_E6BEG[9] ,
    \Tile_X4Y4_E6BEG[8] ,
    \Tile_X4Y4_E6BEG[7] ,
    \Tile_X4Y4_E6BEG[6] ,
    \Tile_X4Y4_E6BEG[5] ,
    \Tile_X4Y4_E6BEG[4] ,
    \Tile_X4Y4_E6BEG[3] ,
    \Tile_X4Y4_E6BEG[2] ,
    \Tile_X4Y4_E6BEG[1] ,
    \Tile_X4Y4_E6BEG[0] }),
    .Tile_X0Y1_EE4END({\Tile_X4Y4_EE4BEG[15] ,
    \Tile_X4Y4_EE4BEG[14] ,
    \Tile_X4Y4_EE4BEG[13] ,
    \Tile_X4Y4_EE4BEG[12] ,
    \Tile_X4Y4_EE4BEG[11] ,
    \Tile_X4Y4_EE4BEG[10] ,
    \Tile_X4Y4_EE4BEG[9] ,
    \Tile_X4Y4_EE4BEG[8] ,
    \Tile_X4Y4_EE4BEG[7] ,
    \Tile_X4Y4_EE4BEG[6] ,
    \Tile_X4Y4_EE4BEG[5] ,
    \Tile_X4Y4_EE4BEG[4] ,
    \Tile_X4Y4_EE4BEG[3] ,
    \Tile_X4Y4_EE4BEG[2] ,
    \Tile_X4Y4_EE4BEG[1] ,
    \Tile_X4Y4_EE4BEG[0] }),
    .Tile_X0Y1_FrameData({\Tile_X4Y4_FrameData_O[31] ,
    \Tile_X4Y4_FrameData_O[30] ,
    \Tile_X4Y4_FrameData_O[29] ,
    \Tile_X4Y4_FrameData_O[28] ,
    \Tile_X4Y4_FrameData_O[27] ,
    \Tile_X4Y4_FrameData_O[26] ,
    \Tile_X4Y4_FrameData_O[25] ,
    \Tile_X4Y4_FrameData_O[24] ,
    \Tile_X4Y4_FrameData_O[23] ,
    \Tile_X4Y4_FrameData_O[22] ,
    \Tile_X4Y4_FrameData_O[21] ,
    \Tile_X4Y4_FrameData_O[20] ,
    \Tile_X4Y4_FrameData_O[19] ,
    \Tile_X4Y4_FrameData_O[18] ,
    \Tile_X4Y4_FrameData_O[17] ,
    \Tile_X4Y4_FrameData_O[16] ,
    \Tile_X4Y4_FrameData_O[15] ,
    \Tile_X4Y4_FrameData_O[14] ,
    \Tile_X4Y4_FrameData_O[13] ,
    \Tile_X4Y4_FrameData_O[12] ,
    \Tile_X4Y4_FrameData_O[11] ,
    \Tile_X4Y4_FrameData_O[10] ,
    \Tile_X4Y4_FrameData_O[9] ,
    \Tile_X4Y4_FrameData_O[8] ,
    \Tile_X4Y4_FrameData_O[7] ,
    \Tile_X4Y4_FrameData_O[6] ,
    \Tile_X4Y4_FrameData_O[5] ,
    \Tile_X4Y4_FrameData_O[4] ,
    \Tile_X4Y4_FrameData_O[3] ,
    \Tile_X4Y4_FrameData_O[2] ,
    \Tile_X4Y4_FrameData_O[1] ,
    \Tile_X4Y4_FrameData_O[0] }),
    .Tile_X0Y1_FrameData_O({\Tile_X5Y4_FrameData_O[31] ,
    \Tile_X5Y4_FrameData_O[30] ,
    \Tile_X5Y4_FrameData_O[29] ,
    \Tile_X5Y4_FrameData_O[28] ,
    \Tile_X5Y4_FrameData_O[27] ,
    \Tile_X5Y4_FrameData_O[26] ,
    \Tile_X5Y4_FrameData_O[25] ,
    \Tile_X5Y4_FrameData_O[24] ,
    \Tile_X5Y4_FrameData_O[23] ,
    \Tile_X5Y4_FrameData_O[22] ,
    \Tile_X5Y4_FrameData_O[21] ,
    \Tile_X5Y4_FrameData_O[20] ,
    \Tile_X5Y4_FrameData_O[19] ,
    \Tile_X5Y4_FrameData_O[18] ,
    \Tile_X5Y4_FrameData_O[17] ,
    \Tile_X5Y4_FrameData_O[16] ,
    \Tile_X5Y4_FrameData_O[15] ,
    \Tile_X5Y4_FrameData_O[14] ,
    \Tile_X5Y4_FrameData_O[13] ,
    \Tile_X5Y4_FrameData_O[12] ,
    \Tile_X5Y4_FrameData_O[11] ,
    \Tile_X5Y4_FrameData_O[10] ,
    \Tile_X5Y4_FrameData_O[9] ,
    \Tile_X5Y4_FrameData_O[8] ,
    \Tile_X5Y4_FrameData_O[7] ,
    \Tile_X5Y4_FrameData_O[6] ,
    \Tile_X5Y4_FrameData_O[5] ,
    \Tile_X5Y4_FrameData_O[4] ,
    \Tile_X5Y4_FrameData_O[3] ,
    \Tile_X5Y4_FrameData_O[2] ,
    \Tile_X5Y4_FrameData_O[1] ,
    \Tile_X5Y4_FrameData_O[0] }),
    .Tile_X0Y1_FrameStrobe({\Tile_X5Y5_FrameStrobe_O[19] ,
    \Tile_X5Y5_FrameStrobe_O[18] ,
    \Tile_X5Y5_FrameStrobe_O[17] ,
    \Tile_X5Y5_FrameStrobe_O[16] ,
    \Tile_X5Y5_FrameStrobe_O[15] ,
    \Tile_X5Y5_FrameStrobe_O[14] ,
    \Tile_X5Y5_FrameStrobe_O[13] ,
    \Tile_X5Y5_FrameStrobe_O[12] ,
    \Tile_X5Y5_FrameStrobe_O[11] ,
    \Tile_X5Y5_FrameStrobe_O[10] ,
    \Tile_X5Y5_FrameStrobe_O[9] ,
    \Tile_X5Y5_FrameStrobe_O[8] ,
    \Tile_X5Y5_FrameStrobe_O[7] ,
    \Tile_X5Y5_FrameStrobe_O[6] ,
    \Tile_X5Y5_FrameStrobe_O[5] ,
    \Tile_X5Y5_FrameStrobe_O[4] ,
    \Tile_X5Y5_FrameStrobe_O[3] ,
    \Tile_X5Y5_FrameStrobe_O[2] ,
    \Tile_X5Y5_FrameStrobe_O[1] ,
    \Tile_X5Y5_FrameStrobe_O[0] }),
    .Tile_X0Y1_N1END({\Tile_X5Y5_N1BEG[3] ,
    \Tile_X5Y5_N1BEG[2] ,
    \Tile_X5Y5_N1BEG[1] ,
    \Tile_X5Y5_N1BEG[0] }),
    .Tile_X0Y1_N2END({\Tile_X5Y5_N2BEGb[7] ,
    \Tile_X5Y5_N2BEGb[6] ,
    \Tile_X5Y5_N2BEGb[5] ,
    \Tile_X5Y5_N2BEGb[4] ,
    \Tile_X5Y5_N2BEGb[3] ,
    \Tile_X5Y5_N2BEGb[2] ,
    \Tile_X5Y5_N2BEGb[1] ,
    \Tile_X5Y5_N2BEGb[0] }),
    .Tile_X0Y1_N2MID({\Tile_X5Y5_N2BEG[7] ,
    \Tile_X5Y5_N2BEG[6] ,
    \Tile_X5Y5_N2BEG[5] ,
    \Tile_X5Y5_N2BEG[4] ,
    \Tile_X5Y5_N2BEG[3] ,
    \Tile_X5Y5_N2BEG[2] ,
    \Tile_X5Y5_N2BEG[1] ,
    \Tile_X5Y5_N2BEG[0] }),
    .Tile_X0Y1_N4END({\Tile_X5Y5_N4BEG[15] ,
    \Tile_X5Y5_N4BEG[14] ,
    \Tile_X5Y5_N4BEG[13] ,
    \Tile_X5Y5_N4BEG[12] ,
    \Tile_X5Y5_N4BEG[11] ,
    \Tile_X5Y5_N4BEG[10] ,
    \Tile_X5Y5_N4BEG[9] ,
    \Tile_X5Y5_N4BEG[8] ,
    \Tile_X5Y5_N4BEG[7] ,
    \Tile_X5Y5_N4BEG[6] ,
    \Tile_X5Y5_N4BEG[5] ,
    \Tile_X5Y5_N4BEG[4] ,
    \Tile_X5Y5_N4BEG[3] ,
    \Tile_X5Y5_N4BEG[2] ,
    \Tile_X5Y5_N4BEG[1] ,
    \Tile_X5Y5_N4BEG[0] }),
    .Tile_X0Y1_S1BEG({\Tile_X5Y4_S1BEG[3] ,
    \Tile_X5Y4_S1BEG[2] ,
    \Tile_X5Y4_S1BEG[1] ,
    \Tile_X5Y4_S1BEG[0] }),
    .Tile_X0Y1_S2BEG({\Tile_X5Y4_S2BEG[7] ,
    \Tile_X5Y4_S2BEG[6] ,
    \Tile_X5Y4_S2BEG[5] ,
    \Tile_X5Y4_S2BEG[4] ,
    \Tile_X5Y4_S2BEG[3] ,
    \Tile_X5Y4_S2BEG[2] ,
    \Tile_X5Y4_S2BEG[1] ,
    \Tile_X5Y4_S2BEG[0] }),
    .Tile_X0Y1_S2BEGb({\Tile_X5Y4_S2BEGb[7] ,
    \Tile_X5Y4_S2BEGb[6] ,
    \Tile_X5Y4_S2BEGb[5] ,
    \Tile_X5Y4_S2BEGb[4] ,
    \Tile_X5Y4_S2BEGb[3] ,
    \Tile_X5Y4_S2BEGb[2] ,
    \Tile_X5Y4_S2BEGb[1] ,
    \Tile_X5Y4_S2BEGb[0] }),
    .Tile_X0Y1_S4BEG({\Tile_X5Y4_S4BEG[15] ,
    \Tile_X5Y4_S4BEG[14] ,
    \Tile_X5Y4_S4BEG[13] ,
    \Tile_X5Y4_S4BEG[12] ,
    \Tile_X5Y4_S4BEG[11] ,
    \Tile_X5Y4_S4BEG[10] ,
    \Tile_X5Y4_S4BEG[9] ,
    \Tile_X5Y4_S4BEG[8] ,
    \Tile_X5Y4_S4BEG[7] ,
    \Tile_X5Y4_S4BEG[6] ,
    \Tile_X5Y4_S4BEG[5] ,
    \Tile_X5Y4_S4BEG[4] ,
    \Tile_X5Y4_S4BEG[3] ,
    \Tile_X5Y4_S4BEG[2] ,
    \Tile_X5Y4_S4BEG[1] ,
    \Tile_X5Y4_S4BEG[0] }),
    .Tile_X0Y1_W1BEG({\Tile_X5Y4_W1BEG[3] ,
    \Tile_X5Y4_W1BEG[2] ,
    \Tile_X5Y4_W1BEG[1] ,
    \Tile_X5Y4_W1BEG[0] }),
    .Tile_X0Y1_W2BEG({\Tile_X5Y4_W2BEG[7] ,
    \Tile_X5Y4_W2BEG[6] ,
    \Tile_X5Y4_W2BEG[5] ,
    \Tile_X5Y4_W2BEG[4] ,
    \Tile_X5Y4_W2BEG[3] ,
    \Tile_X5Y4_W2BEG[2] ,
    \Tile_X5Y4_W2BEG[1] ,
    \Tile_X5Y4_W2BEG[0] }),
    .Tile_X0Y1_W2BEGb({\Tile_X5Y4_W2BEGb[7] ,
    \Tile_X5Y4_W2BEGb[6] ,
    \Tile_X5Y4_W2BEGb[5] ,
    \Tile_X5Y4_W2BEGb[4] ,
    \Tile_X5Y4_W2BEGb[3] ,
    \Tile_X5Y4_W2BEGb[2] ,
    \Tile_X5Y4_W2BEGb[1] ,
    \Tile_X5Y4_W2BEGb[0] }),
    .Tile_X0Y1_W6BEG({\Tile_X5Y4_W6BEG[11] ,
    \Tile_X5Y4_W6BEG[10] ,
    \Tile_X5Y4_W6BEG[9] ,
    \Tile_X5Y4_W6BEG[8] ,
    \Tile_X5Y4_W6BEG[7] ,
    \Tile_X5Y4_W6BEG[6] ,
    \Tile_X5Y4_W6BEG[5] ,
    \Tile_X5Y4_W6BEG[4] ,
    \Tile_X5Y4_W6BEG[3] ,
    \Tile_X5Y4_W6BEG[2] ,
    \Tile_X5Y4_W6BEG[1] ,
    \Tile_X5Y4_W6BEG[0] }),
    .Tile_X0Y1_WW4BEG({\Tile_X5Y4_WW4BEG[15] ,
    \Tile_X5Y4_WW4BEG[14] ,
    \Tile_X5Y4_WW4BEG[13] ,
    \Tile_X5Y4_WW4BEG[12] ,
    \Tile_X5Y4_WW4BEG[11] ,
    \Tile_X5Y4_WW4BEG[10] ,
    \Tile_X5Y4_WW4BEG[9] ,
    \Tile_X5Y4_WW4BEG[8] ,
    \Tile_X5Y4_WW4BEG[7] ,
    \Tile_X5Y4_WW4BEG[6] ,
    \Tile_X5Y4_WW4BEG[5] ,
    \Tile_X5Y4_WW4BEG[4] ,
    \Tile_X5Y4_WW4BEG[3] ,
    \Tile_X5Y4_WW4BEG[2] ,
    \Tile_X5Y4_WW4BEG[1] ,
    \Tile_X5Y4_WW4BEG[0] }));
 E_TT_IF Tile_X5Y5_E_TT_IF (.CLK_TT_PROJECT(Tile_X5Y5_CLK_TT_PROJECT),
    .ENA_TT_PROJECT(Tile_X5Y5_ENA_TT_PROJECT),
    .RST_N_TT_PROJECT(Tile_X5Y5_RST_N_TT_PROJECT),
    .UIO_IN_TT_PROJECT0(Tile_X5Y5_UIO_IN_TT_PROJECT0),
    .UIO_IN_TT_PROJECT1(Tile_X5Y5_UIO_IN_TT_PROJECT1),
    .UIO_IN_TT_PROJECT2(Tile_X5Y5_UIO_IN_TT_PROJECT2),
    .UIO_IN_TT_PROJECT3(Tile_X5Y5_UIO_IN_TT_PROJECT3),
    .UIO_IN_TT_PROJECT4(Tile_X5Y5_UIO_IN_TT_PROJECT4),
    .UIO_IN_TT_PROJECT5(Tile_X5Y5_UIO_IN_TT_PROJECT5),
    .UIO_IN_TT_PROJECT6(Tile_X5Y5_UIO_IN_TT_PROJECT6),
    .UIO_IN_TT_PROJECT7(Tile_X5Y5_UIO_IN_TT_PROJECT7),
    .UIO_OE_TT_PROJECT0(Tile_X5Y5_UIO_OE_TT_PROJECT0),
    .UIO_OE_TT_PROJECT1(Tile_X5Y5_UIO_OE_TT_PROJECT1),
    .UIO_OE_TT_PROJECT2(Tile_X5Y5_UIO_OE_TT_PROJECT2),
    .UIO_OE_TT_PROJECT3(Tile_X5Y5_UIO_OE_TT_PROJECT3),
    .UIO_OE_TT_PROJECT4(Tile_X5Y5_UIO_OE_TT_PROJECT4),
    .UIO_OE_TT_PROJECT5(Tile_X5Y5_UIO_OE_TT_PROJECT5),
    .UIO_OE_TT_PROJECT6(Tile_X5Y5_UIO_OE_TT_PROJECT6),
    .UIO_OE_TT_PROJECT7(Tile_X5Y5_UIO_OE_TT_PROJECT7),
    .UIO_OUT_TT_PROJECT0(Tile_X5Y5_UIO_OUT_TT_PROJECT0),
    .UIO_OUT_TT_PROJECT1(Tile_X5Y5_UIO_OUT_TT_PROJECT1),
    .UIO_OUT_TT_PROJECT2(Tile_X5Y5_UIO_OUT_TT_PROJECT2),
    .UIO_OUT_TT_PROJECT3(Tile_X5Y5_UIO_OUT_TT_PROJECT3),
    .UIO_OUT_TT_PROJECT4(Tile_X5Y5_UIO_OUT_TT_PROJECT4),
    .UIO_OUT_TT_PROJECT5(Tile_X5Y5_UIO_OUT_TT_PROJECT5),
    .UIO_OUT_TT_PROJECT6(Tile_X5Y5_UIO_OUT_TT_PROJECT6),
    .UIO_OUT_TT_PROJECT7(Tile_X5Y5_UIO_OUT_TT_PROJECT7),
    .UI_IN_TT_PROJECT0(Tile_X5Y5_UI_IN_TT_PROJECT0),
    .UI_IN_TT_PROJECT1(Tile_X5Y5_UI_IN_TT_PROJECT1),
    .UI_IN_TT_PROJECT2(Tile_X5Y5_UI_IN_TT_PROJECT2),
    .UI_IN_TT_PROJECT3(Tile_X5Y5_UI_IN_TT_PROJECT3),
    .UI_IN_TT_PROJECT4(Tile_X5Y5_UI_IN_TT_PROJECT4),
    .UI_IN_TT_PROJECT5(Tile_X5Y5_UI_IN_TT_PROJECT5),
    .UI_IN_TT_PROJECT6(Tile_X5Y5_UI_IN_TT_PROJECT6),
    .UI_IN_TT_PROJECT7(Tile_X5Y5_UI_IN_TT_PROJECT7),
    .UO_OUT_TT_PROJECT0(Tile_X5Y5_UO_OUT_TT_PROJECT0),
    .UO_OUT_TT_PROJECT1(Tile_X5Y5_UO_OUT_TT_PROJECT1),
    .UO_OUT_TT_PROJECT2(Tile_X5Y5_UO_OUT_TT_PROJECT2),
    .UO_OUT_TT_PROJECT3(Tile_X5Y5_UO_OUT_TT_PROJECT3),
    .UO_OUT_TT_PROJECT4(Tile_X5Y5_UO_OUT_TT_PROJECT4),
    .UO_OUT_TT_PROJECT5(Tile_X5Y5_UO_OUT_TT_PROJECT5),
    .UO_OUT_TT_PROJECT6(Tile_X5Y5_UO_OUT_TT_PROJECT6),
    .UO_OUT_TT_PROJECT7(Tile_X5Y5_UO_OUT_TT_PROJECT7),
    .UserCLK(Tile_X5Y6_UserCLKo),
    .UserCLKo(Tile_X5Y5_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1END({\Tile_X4Y5_E1BEG[3] ,
    \Tile_X4Y5_E1BEG[2] ,
    \Tile_X4Y5_E1BEG[1] ,
    \Tile_X4Y5_E1BEG[0] }),
    .E2END({\Tile_X4Y5_E2BEGb[7] ,
    \Tile_X4Y5_E2BEGb[6] ,
    \Tile_X4Y5_E2BEGb[5] ,
    \Tile_X4Y5_E2BEGb[4] ,
    \Tile_X4Y5_E2BEGb[3] ,
    \Tile_X4Y5_E2BEGb[2] ,
    \Tile_X4Y5_E2BEGb[1] ,
    \Tile_X4Y5_E2BEGb[0] }),
    .E2MID({\Tile_X4Y5_E2BEG[7] ,
    \Tile_X4Y5_E2BEG[6] ,
    \Tile_X4Y5_E2BEG[5] ,
    \Tile_X4Y5_E2BEG[4] ,
    \Tile_X4Y5_E2BEG[3] ,
    \Tile_X4Y5_E2BEG[2] ,
    \Tile_X4Y5_E2BEG[1] ,
    \Tile_X4Y5_E2BEG[0] }),
    .E6END({\Tile_X4Y5_E6BEG[11] ,
    \Tile_X4Y5_E6BEG[10] ,
    \Tile_X4Y5_E6BEG[9] ,
    \Tile_X4Y5_E6BEG[8] ,
    \Tile_X4Y5_E6BEG[7] ,
    \Tile_X4Y5_E6BEG[6] ,
    \Tile_X4Y5_E6BEG[5] ,
    \Tile_X4Y5_E6BEG[4] ,
    \Tile_X4Y5_E6BEG[3] ,
    \Tile_X4Y5_E6BEG[2] ,
    \Tile_X4Y5_E6BEG[1] ,
    \Tile_X4Y5_E6BEG[0] }),
    .EE4END({\Tile_X4Y5_EE4BEG[15] ,
    \Tile_X4Y5_EE4BEG[14] ,
    \Tile_X4Y5_EE4BEG[13] ,
    \Tile_X4Y5_EE4BEG[12] ,
    \Tile_X4Y5_EE4BEG[11] ,
    \Tile_X4Y5_EE4BEG[10] ,
    \Tile_X4Y5_EE4BEG[9] ,
    \Tile_X4Y5_EE4BEG[8] ,
    \Tile_X4Y5_EE4BEG[7] ,
    \Tile_X4Y5_EE4BEG[6] ,
    \Tile_X4Y5_EE4BEG[5] ,
    \Tile_X4Y5_EE4BEG[4] ,
    \Tile_X4Y5_EE4BEG[3] ,
    \Tile_X4Y5_EE4BEG[2] ,
    \Tile_X4Y5_EE4BEG[1] ,
    \Tile_X4Y5_EE4BEG[0] }),
    .FrameData({\Tile_X4Y5_FrameData_O[31] ,
    \Tile_X4Y5_FrameData_O[30] ,
    \Tile_X4Y5_FrameData_O[29] ,
    \Tile_X4Y5_FrameData_O[28] ,
    \Tile_X4Y5_FrameData_O[27] ,
    \Tile_X4Y5_FrameData_O[26] ,
    \Tile_X4Y5_FrameData_O[25] ,
    \Tile_X4Y5_FrameData_O[24] ,
    \Tile_X4Y5_FrameData_O[23] ,
    \Tile_X4Y5_FrameData_O[22] ,
    \Tile_X4Y5_FrameData_O[21] ,
    \Tile_X4Y5_FrameData_O[20] ,
    \Tile_X4Y5_FrameData_O[19] ,
    \Tile_X4Y5_FrameData_O[18] ,
    \Tile_X4Y5_FrameData_O[17] ,
    \Tile_X4Y5_FrameData_O[16] ,
    \Tile_X4Y5_FrameData_O[15] ,
    \Tile_X4Y5_FrameData_O[14] ,
    \Tile_X4Y5_FrameData_O[13] ,
    \Tile_X4Y5_FrameData_O[12] ,
    \Tile_X4Y5_FrameData_O[11] ,
    \Tile_X4Y5_FrameData_O[10] ,
    \Tile_X4Y5_FrameData_O[9] ,
    \Tile_X4Y5_FrameData_O[8] ,
    \Tile_X4Y5_FrameData_O[7] ,
    \Tile_X4Y5_FrameData_O[6] ,
    \Tile_X4Y5_FrameData_O[5] ,
    \Tile_X4Y5_FrameData_O[4] ,
    \Tile_X4Y5_FrameData_O[3] ,
    \Tile_X4Y5_FrameData_O[2] ,
    \Tile_X4Y5_FrameData_O[1] ,
    \Tile_X4Y5_FrameData_O[0] }),
    .FrameData_O({\Tile_X5Y5_FrameData_O[31] ,
    \Tile_X5Y5_FrameData_O[30] ,
    \Tile_X5Y5_FrameData_O[29] ,
    \Tile_X5Y5_FrameData_O[28] ,
    \Tile_X5Y5_FrameData_O[27] ,
    \Tile_X5Y5_FrameData_O[26] ,
    \Tile_X5Y5_FrameData_O[25] ,
    \Tile_X5Y5_FrameData_O[24] ,
    \Tile_X5Y5_FrameData_O[23] ,
    \Tile_X5Y5_FrameData_O[22] ,
    \Tile_X5Y5_FrameData_O[21] ,
    \Tile_X5Y5_FrameData_O[20] ,
    \Tile_X5Y5_FrameData_O[19] ,
    \Tile_X5Y5_FrameData_O[18] ,
    \Tile_X5Y5_FrameData_O[17] ,
    \Tile_X5Y5_FrameData_O[16] ,
    \Tile_X5Y5_FrameData_O[15] ,
    \Tile_X5Y5_FrameData_O[14] ,
    \Tile_X5Y5_FrameData_O[13] ,
    \Tile_X5Y5_FrameData_O[12] ,
    \Tile_X5Y5_FrameData_O[11] ,
    \Tile_X5Y5_FrameData_O[10] ,
    \Tile_X5Y5_FrameData_O[9] ,
    \Tile_X5Y5_FrameData_O[8] ,
    \Tile_X5Y5_FrameData_O[7] ,
    \Tile_X5Y5_FrameData_O[6] ,
    \Tile_X5Y5_FrameData_O[5] ,
    \Tile_X5Y5_FrameData_O[4] ,
    \Tile_X5Y5_FrameData_O[3] ,
    \Tile_X5Y5_FrameData_O[2] ,
    \Tile_X5Y5_FrameData_O[1] ,
    \Tile_X5Y5_FrameData_O[0] }),
    .FrameStrobe({\Tile_X5Y6_FrameStrobe_O[19] ,
    \Tile_X5Y6_FrameStrobe_O[18] ,
    \Tile_X5Y6_FrameStrobe_O[17] ,
    \Tile_X5Y6_FrameStrobe_O[16] ,
    \Tile_X5Y6_FrameStrobe_O[15] ,
    \Tile_X5Y6_FrameStrobe_O[14] ,
    \Tile_X5Y6_FrameStrobe_O[13] ,
    \Tile_X5Y6_FrameStrobe_O[12] ,
    \Tile_X5Y6_FrameStrobe_O[11] ,
    \Tile_X5Y6_FrameStrobe_O[10] ,
    \Tile_X5Y6_FrameStrobe_O[9] ,
    \Tile_X5Y6_FrameStrobe_O[8] ,
    \Tile_X5Y6_FrameStrobe_O[7] ,
    \Tile_X5Y6_FrameStrobe_O[6] ,
    \Tile_X5Y6_FrameStrobe_O[5] ,
    \Tile_X5Y6_FrameStrobe_O[4] ,
    \Tile_X5Y6_FrameStrobe_O[3] ,
    \Tile_X5Y6_FrameStrobe_O[2] ,
    \Tile_X5Y6_FrameStrobe_O[1] ,
    \Tile_X5Y6_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X5Y5_FrameStrobe_O[19] ,
    \Tile_X5Y5_FrameStrobe_O[18] ,
    \Tile_X5Y5_FrameStrobe_O[17] ,
    \Tile_X5Y5_FrameStrobe_O[16] ,
    \Tile_X5Y5_FrameStrobe_O[15] ,
    \Tile_X5Y5_FrameStrobe_O[14] ,
    \Tile_X5Y5_FrameStrobe_O[13] ,
    \Tile_X5Y5_FrameStrobe_O[12] ,
    \Tile_X5Y5_FrameStrobe_O[11] ,
    \Tile_X5Y5_FrameStrobe_O[10] ,
    \Tile_X5Y5_FrameStrobe_O[9] ,
    \Tile_X5Y5_FrameStrobe_O[8] ,
    \Tile_X5Y5_FrameStrobe_O[7] ,
    \Tile_X5Y5_FrameStrobe_O[6] ,
    \Tile_X5Y5_FrameStrobe_O[5] ,
    \Tile_X5Y5_FrameStrobe_O[4] ,
    \Tile_X5Y5_FrameStrobe_O[3] ,
    \Tile_X5Y5_FrameStrobe_O[2] ,
    \Tile_X5Y5_FrameStrobe_O[1] ,
    \Tile_X5Y5_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X5Y5_N1BEG[3] ,
    \Tile_X5Y5_N1BEG[2] ,
    \Tile_X5Y5_N1BEG[1] ,
    \Tile_X5Y5_N1BEG[0] }),
    .N1END({\Tile_X5Y6_N1BEG[3] ,
    \Tile_X5Y6_N1BEG[2] ,
    \Tile_X5Y6_N1BEG[1] ,
    \Tile_X5Y6_N1BEG[0] }),
    .N2BEG({\Tile_X5Y5_N2BEG[7] ,
    \Tile_X5Y5_N2BEG[6] ,
    \Tile_X5Y5_N2BEG[5] ,
    \Tile_X5Y5_N2BEG[4] ,
    \Tile_X5Y5_N2BEG[3] ,
    \Tile_X5Y5_N2BEG[2] ,
    \Tile_X5Y5_N2BEG[1] ,
    \Tile_X5Y5_N2BEG[0] }),
    .N2BEGb({\Tile_X5Y5_N2BEGb[7] ,
    \Tile_X5Y5_N2BEGb[6] ,
    \Tile_X5Y5_N2BEGb[5] ,
    \Tile_X5Y5_N2BEGb[4] ,
    \Tile_X5Y5_N2BEGb[3] ,
    \Tile_X5Y5_N2BEGb[2] ,
    \Tile_X5Y5_N2BEGb[1] ,
    \Tile_X5Y5_N2BEGb[0] }),
    .N2END({\Tile_X5Y6_N2BEGb[7] ,
    \Tile_X5Y6_N2BEGb[6] ,
    \Tile_X5Y6_N2BEGb[5] ,
    \Tile_X5Y6_N2BEGb[4] ,
    \Tile_X5Y6_N2BEGb[3] ,
    \Tile_X5Y6_N2BEGb[2] ,
    \Tile_X5Y6_N2BEGb[1] ,
    \Tile_X5Y6_N2BEGb[0] }),
    .N2MID({\Tile_X5Y6_N2BEG[7] ,
    \Tile_X5Y6_N2BEG[6] ,
    \Tile_X5Y6_N2BEG[5] ,
    \Tile_X5Y6_N2BEG[4] ,
    \Tile_X5Y6_N2BEG[3] ,
    \Tile_X5Y6_N2BEG[2] ,
    \Tile_X5Y6_N2BEG[1] ,
    \Tile_X5Y6_N2BEG[0] }),
    .N4BEG({\Tile_X5Y5_N4BEG[15] ,
    \Tile_X5Y5_N4BEG[14] ,
    \Tile_X5Y5_N4BEG[13] ,
    \Tile_X5Y5_N4BEG[12] ,
    \Tile_X5Y5_N4BEG[11] ,
    \Tile_X5Y5_N4BEG[10] ,
    \Tile_X5Y5_N4BEG[9] ,
    \Tile_X5Y5_N4BEG[8] ,
    \Tile_X5Y5_N4BEG[7] ,
    \Tile_X5Y5_N4BEG[6] ,
    \Tile_X5Y5_N4BEG[5] ,
    \Tile_X5Y5_N4BEG[4] ,
    \Tile_X5Y5_N4BEG[3] ,
    \Tile_X5Y5_N4BEG[2] ,
    \Tile_X5Y5_N4BEG[1] ,
    \Tile_X5Y5_N4BEG[0] }),
    .N4END({\Tile_X5Y6_N4BEG[15] ,
    \Tile_X5Y6_N4BEG[14] ,
    \Tile_X5Y6_N4BEG[13] ,
    \Tile_X5Y6_N4BEG[12] ,
    \Tile_X5Y6_N4BEG[11] ,
    \Tile_X5Y6_N4BEG[10] ,
    \Tile_X5Y6_N4BEG[9] ,
    \Tile_X5Y6_N4BEG[8] ,
    \Tile_X5Y6_N4BEG[7] ,
    \Tile_X5Y6_N4BEG[6] ,
    \Tile_X5Y6_N4BEG[5] ,
    \Tile_X5Y6_N4BEG[4] ,
    \Tile_X5Y6_N4BEG[3] ,
    \Tile_X5Y6_N4BEG[2] ,
    \Tile_X5Y6_N4BEG[1] ,
    \Tile_X5Y6_N4BEG[0] }),
    .S1BEG({\Tile_X5Y5_S1BEG[3] ,
    \Tile_X5Y5_S1BEG[2] ,
    \Tile_X5Y5_S1BEG[1] ,
    \Tile_X5Y5_S1BEG[0] }),
    .S1END({\Tile_X5Y4_S1BEG[3] ,
    \Tile_X5Y4_S1BEG[2] ,
    \Tile_X5Y4_S1BEG[1] ,
    \Tile_X5Y4_S1BEG[0] }),
    .S2BEG({\Tile_X5Y5_S2BEG[7] ,
    \Tile_X5Y5_S2BEG[6] ,
    \Tile_X5Y5_S2BEG[5] ,
    \Tile_X5Y5_S2BEG[4] ,
    \Tile_X5Y5_S2BEG[3] ,
    \Tile_X5Y5_S2BEG[2] ,
    \Tile_X5Y5_S2BEG[1] ,
    \Tile_X5Y5_S2BEG[0] }),
    .S2BEGb({\Tile_X5Y5_S2BEGb[7] ,
    \Tile_X5Y5_S2BEGb[6] ,
    \Tile_X5Y5_S2BEGb[5] ,
    \Tile_X5Y5_S2BEGb[4] ,
    \Tile_X5Y5_S2BEGb[3] ,
    \Tile_X5Y5_S2BEGb[2] ,
    \Tile_X5Y5_S2BEGb[1] ,
    \Tile_X5Y5_S2BEGb[0] }),
    .S2END({\Tile_X5Y4_S2BEGb[7] ,
    \Tile_X5Y4_S2BEGb[6] ,
    \Tile_X5Y4_S2BEGb[5] ,
    \Tile_X5Y4_S2BEGb[4] ,
    \Tile_X5Y4_S2BEGb[3] ,
    \Tile_X5Y4_S2BEGb[2] ,
    \Tile_X5Y4_S2BEGb[1] ,
    \Tile_X5Y4_S2BEGb[0] }),
    .S2MID({\Tile_X5Y4_S2BEG[7] ,
    \Tile_X5Y4_S2BEG[6] ,
    \Tile_X5Y4_S2BEG[5] ,
    \Tile_X5Y4_S2BEG[4] ,
    \Tile_X5Y4_S2BEG[3] ,
    \Tile_X5Y4_S2BEG[2] ,
    \Tile_X5Y4_S2BEG[1] ,
    \Tile_X5Y4_S2BEG[0] }),
    .S4BEG({\Tile_X5Y5_S4BEG[15] ,
    \Tile_X5Y5_S4BEG[14] ,
    \Tile_X5Y5_S4BEG[13] ,
    \Tile_X5Y5_S4BEG[12] ,
    \Tile_X5Y5_S4BEG[11] ,
    \Tile_X5Y5_S4BEG[10] ,
    \Tile_X5Y5_S4BEG[9] ,
    \Tile_X5Y5_S4BEG[8] ,
    \Tile_X5Y5_S4BEG[7] ,
    \Tile_X5Y5_S4BEG[6] ,
    \Tile_X5Y5_S4BEG[5] ,
    \Tile_X5Y5_S4BEG[4] ,
    \Tile_X5Y5_S4BEG[3] ,
    \Tile_X5Y5_S4BEG[2] ,
    \Tile_X5Y5_S4BEG[1] ,
    \Tile_X5Y5_S4BEG[0] }),
    .S4END({\Tile_X5Y4_S4BEG[15] ,
    \Tile_X5Y4_S4BEG[14] ,
    \Tile_X5Y4_S4BEG[13] ,
    \Tile_X5Y4_S4BEG[12] ,
    \Tile_X5Y4_S4BEG[11] ,
    \Tile_X5Y4_S4BEG[10] ,
    \Tile_X5Y4_S4BEG[9] ,
    \Tile_X5Y4_S4BEG[8] ,
    \Tile_X5Y4_S4BEG[7] ,
    \Tile_X5Y4_S4BEG[6] ,
    \Tile_X5Y4_S4BEG[5] ,
    \Tile_X5Y4_S4BEG[4] ,
    \Tile_X5Y4_S4BEG[3] ,
    \Tile_X5Y4_S4BEG[2] ,
    \Tile_X5Y4_S4BEG[1] ,
    \Tile_X5Y4_S4BEG[0] }),
    .W1BEG({\Tile_X5Y5_W1BEG[3] ,
    \Tile_X5Y5_W1BEG[2] ,
    \Tile_X5Y5_W1BEG[1] ,
    \Tile_X5Y5_W1BEG[0] }),
    .W2BEG({\Tile_X5Y5_W2BEG[7] ,
    \Tile_X5Y5_W2BEG[6] ,
    \Tile_X5Y5_W2BEG[5] ,
    \Tile_X5Y5_W2BEG[4] ,
    \Tile_X5Y5_W2BEG[3] ,
    \Tile_X5Y5_W2BEG[2] ,
    \Tile_X5Y5_W2BEG[1] ,
    \Tile_X5Y5_W2BEG[0] }),
    .W2BEGb({\Tile_X5Y5_W2BEGb[7] ,
    \Tile_X5Y5_W2BEGb[6] ,
    \Tile_X5Y5_W2BEGb[5] ,
    \Tile_X5Y5_W2BEGb[4] ,
    \Tile_X5Y5_W2BEGb[3] ,
    \Tile_X5Y5_W2BEGb[2] ,
    \Tile_X5Y5_W2BEGb[1] ,
    \Tile_X5Y5_W2BEGb[0] }),
    .W6BEG({\Tile_X5Y5_W6BEG[11] ,
    \Tile_X5Y5_W6BEG[10] ,
    \Tile_X5Y5_W6BEG[9] ,
    \Tile_X5Y5_W6BEG[8] ,
    \Tile_X5Y5_W6BEG[7] ,
    \Tile_X5Y5_W6BEG[6] ,
    \Tile_X5Y5_W6BEG[5] ,
    \Tile_X5Y5_W6BEG[4] ,
    \Tile_X5Y5_W6BEG[3] ,
    \Tile_X5Y5_W6BEG[2] ,
    \Tile_X5Y5_W6BEG[1] ,
    \Tile_X5Y5_W6BEG[0] }),
    .WW4BEG({\Tile_X5Y5_WW4BEG[15] ,
    \Tile_X5Y5_WW4BEG[14] ,
    \Tile_X5Y5_WW4BEG[13] ,
    \Tile_X5Y5_WW4BEG[12] ,
    \Tile_X5Y5_WW4BEG[11] ,
    \Tile_X5Y5_WW4BEG[10] ,
    \Tile_X5Y5_WW4BEG[9] ,
    \Tile_X5Y5_WW4BEG[8] ,
    \Tile_X5Y5_WW4BEG[7] ,
    \Tile_X5Y5_WW4BEG[6] ,
    \Tile_X5Y5_WW4BEG[5] ,
    \Tile_X5Y5_WW4BEG[4] ,
    \Tile_X5Y5_WW4BEG[3] ,
    \Tile_X5Y5_WW4BEG[2] ,
    \Tile_X5Y5_WW4BEG[1] ,
    \Tile_X5Y5_WW4BEG[0] }));
 E_TT_IF Tile_X5Y6_E_TT_IF (.CLK_TT_PROJECT(Tile_X5Y6_CLK_TT_PROJECT),
    .ENA_TT_PROJECT(Tile_X5Y6_ENA_TT_PROJECT),
    .RST_N_TT_PROJECT(Tile_X5Y6_RST_N_TT_PROJECT),
    .UIO_IN_TT_PROJECT0(Tile_X5Y6_UIO_IN_TT_PROJECT0),
    .UIO_IN_TT_PROJECT1(Tile_X5Y6_UIO_IN_TT_PROJECT1),
    .UIO_IN_TT_PROJECT2(Tile_X5Y6_UIO_IN_TT_PROJECT2),
    .UIO_IN_TT_PROJECT3(Tile_X5Y6_UIO_IN_TT_PROJECT3),
    .UIO_IN_TT_PROJECT4(Tile_X5Y6_UIO_IN_TT_PROJECT4),
    .UIO_IN_TT_PROJECT5(Tile_X5Y6_UIO_IN_TT_PROJECT5),
    .UIO_IN_TT_PROJECT6(Tile_X5Y6_UIO_IN_TT_PROJECT6),
    .UIO_IN_TT_PROJECT7(Tile_X5Y6_UIO_IN_TT_PROJECT7),
    .UIO_OE_TT_PROJECT0(Tile_X5Y6_UIO_OE_TT_PROJECT0),
    .UIO_OE_TT_PROJECT1(Tile_X5Y6_UIO_OE_TT_PROJECT1),
    .UIO_OE_TT_PROJECT2(Tile_X5Y6_UIO_OE_TT_PROJECT2),
    .UIO_OE_TT_PROJECT3(Tile_X5Y6_UIO_OE_TT_PROJECT3),
    .UIO_OE_TT_PROJECT4(Tile_X5Y6_UIO_OE_TT_PROJECT4),
    .UIO_OE_TT_PROJECT5(Tile_X5Y6_UIO_OE_TT_PROJECT5),
    .UIO_OE_TT_PROJECT6(Tile_X5Y6_UIO_OE_TT_PROJECT6),
    .UIO_OE_TT_PROJECT7(Tile_X5Y6_UIO_OE_TT_PROJECT7),
    .UIO_OUT_TT_PROJECT0(Tile_X5Y6_UIO_OUT_TT_PROJECT0),
    .UIO_OUT_TT_PROJECT1(Tile_X5Y6_UIO_OUT_TT_PROJECT1),
    .UIO_OUT_TT_PROJECT2(Tile_X5Y6_UIO_OUT_TT_PROJECT2),
    .UIO_OUT_TT_PROJECT3(Tile_X5Y6_UIO_OUT_TT_PROJECT3),
    .UIO_OUT_TT_PROJECT4(Tile_X5Y6_UIO_OUT_TT_PROJECT4),
    .UIO_OUT_TT_PROJECT5(Tile_X5Y6_UIO_OUT_TT_PROJECT5),
    .UIO_OUT_TT_PROJECT6(Tile_X5Y6_UIO_OUT_TT_PROJECT6),
    .UIO_OUT_TT_PROJECT7(Tile_X5Y6_UIO_OUT_TT_PROJECT7),
    .UI_IN_TT_PROJECT0(Tile_X5Y6_UI_IN_TT_PROJECT0),
    .UI_IN_TT_PROJECT1(Tile_X5Y6_UI_IN_TT_PROJECT1),
    .UI_IN_TT_PROJECT2(Tile_X5Y6_UI_IN_TT_PROJECT2),
    .UI_IN_TT_PROJECT3(Tile_X5Y6_UI_IN_TT_PROJECT3),
    .UI_IN_TT_PROJECT4(Tile_X5Y6_UI_IN_TT_PROJECT4),
    .UI_IN_TT_PROJECT5(Tile_X5Y6_UI_IN_TT_PROJECT5),
    .UI_IN_TT_PROJECT6(Tile_X5Y6_UI_IN_TT_PROJECT6),
    .UI_IN_TT_PROJECT7(Tile_X5Y6_UI_IN_TT_PROJECT7),
    .UO_OUT_TT_PROJECT0(Tile_X5Y6_UO_OUT_TT_PROJECT0),
    .UO_OUT_TT_PROJECT1(Tile_X5Y6_UO_OUT_TT_PROJECT1),
    .UO_OUT_TT_PROJECT2(Tile_X5Y6_UO_OUT_TT_PROJECT2),
    .UO_OUT_TT_PROJECT3(Tile_X5Y6_UO_OUT_TT_PROJECT3),
    .UO_OUT_TT_PROJECT4(Tile_X5Y6_UO_OUT_TT_PROJECT4),
    .UO_OUT_TT_PROJECT5(Tile_X5Y6_UO_OUT_TT_PROJECT5),
    .UO_OUT_TT_PROJECT6(Tile_X5Y6_UO_OUT_TT_PROJECT6),
    .UO_OUT_TT_PROJECT7(Tile_X5Y6_UO_OUT_TT_PROJECT7),
    .UserCLK(Tile_X5Y7_UserCLKo),
    .UserCLKo(Tile_X5Y6_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1END({\Tile_X4Y6_E1BEG[3] ,
    \Tile_X4Y6_E1BEG[2] ,
    \Tile_X4Y6_E1BEG[1] ,
    \Tile_X4Y6_E1BEG[0] }),
    .E2END({\Tile_X4Y6_E2BEGb[7] ,
    \Tile_X4Y6_E2BEGb[6] ,
    \Tile_X4Y6_E2BEGb[5] ,
    \Tile_X4Y6_E2BEGb[4] ,
    \Tile_X4Y6_E2BEGb[3] ,
    \Tile_X4Y6_E2BEGb[2] ,
    \Tile_X4Y6_E2BEGb[1] ,
    \Tile_X4Y6_E2BEGb[0] }),
    .E2MID({\Tile_X4Y6_E2BEG[7] ,
    \Tile_X4Y6_E2BEG[6] ,
    \Tile_X4Y6_E2BEG[5] ,
    \Tile_X4Y6_E2BEG[4] ,
    \Tile_X4Y6_E2BEG[3] ,
    \Tile_X4Y6_E2BEG[2] ,
    \Tile_X4Y6_E2BEG[1] ,
    \Tile_X4Y6_E2BEG[0] }),
    .E6END({\Tile_X4Y6_E6BEG[11] ,
    \Tile_X4Y6_E6BEG[10] ,
    \Tile_X4Y6_E6BEG[9] ,
    \Tile_X4Y6_E6BEG[8] ,
    \Tile_X4Y6_E6BEG[7] ,
    \Tile_X4Y6_E6BEG[6] ,
    \Tile_X4Y6_E6BEG[5] ,
    \Tile_X4Y6_E6BEG[4] ,
    \Tile_X4Y6_E6BEG[3] ,
    \Tile_X4Y6_E6BEG[2] ,
    \Tile_X4Y6_E6BEG[1] ,
    \Tile_X4Y6_E6BEG[0] }),
    .EE4END({\Tile_X4Y6_EE4BEG[15] ,
    \Tile_X4Y6_EE4BEG[14] ,
    \Tile_X4Y6_EE4BEG[13] ,
    \Tile_X4Y6_EE4BEG[12] ,
    \Tile_X4Y6_EE4BEG[11] ,
    \Tile_X4Y6_EE4BEG[10] ,
    \Tile_X4Y6_EE4BEG[9] ,
    \Tile_X4Y6_EE4BEG[8] ,
    \Tile_X4Y6_EE4BEG[7] ,
    \Tile_X4Y6_EE4BEG[6] ,
    \Tile_X4Y6_EE4BEG[5] ,
    \Tile_X4Y6_EE4BEG[4] ,
    \Tile_X4Y6_EE4BEG[3] ,
    \Tile_X4Y6_EE4BEG[2] ,
    \Tile_X4Y6_EE4BEG[1] ,
    \Tile_X4Y6_EE4BEG[0] }),
    .FrameData({\Tile_X4Y6_FrameData_O[31] ,
    \Tile_X4Y6_FrameData_O[30] ,
    \Tile_X4Y6_FrameData_O[29] ,
    \Tile_X4Y6_FrameData_O[28] ,
    \Tile_X4Y6_FrameData_O[27] ,
    \Tile_X4Y6_FrameData_O[26] ,
    \Tile_X4Y6_FrameData_O[25] ,
    \Tile_X4Y6_FrameData_O[24] ,
    \Tile_X4Y6_FrameData_O[23] ,
    \Tile_X4Y6_FrameData_O[22] ,
    \Tile_X4Y6_FrameData_O[21] ,
    \Tile_X4Y6_FrameData_O[20] ,
    \Tile_X4Y6_FrameData_O[19] ,
    \Tile_X4Y6_FrameData_O[18] ,
    \Tile_X4Y6_FrameData_O[17] ,
    \Tile_X4Y6_FrameData_O[16] ,
    \Tile_X4Y6_FrameData_O[15] ,
    \Tile_X4Y6_FrameData_O[14] ,
    \Tile_X4Y6_FrameData_O[13] ,
    \Tile_X4Y6_FrameData_O[12] ,
    \Tile_X4Y6_FrameData_O[11] ,
    \Tile_X4Y6_FrameData_O[10] ,
    \Tile_X4Y6_FrameData_O[9] ,
    \Tile_X4Y6_FrameData_O[8] ,
    \Tile_X4Y6_FrameData_O[7] ,
    \Tile_X4Y6_FrameData_O[6] ,
    \Tile_X4Y6_FrameData_O[5] ,
    \Tile_X4Y6_FrameData_O[4] ,
    \Tile_X4Y6_FrameData_O[3] ,
    \Tile_X4Y6_FrameData_O[2] ,
    \Tile_X4Y6_FrameData_O[1] ,
    \Tile_X4Y6_FrameData_O[0] }),
    .FrameData_O({\Tile_X5Y6_FrameData_O[31] ,
    \Tile_X5Y6_FrameData_O[30] ,
    \Tile_X5Y6_FrameData_O[29] ,
    \Tile_X5Y6_FrameData_O[28] ,
    \Tile_X5Y6_FrameData_O[27] ,
    \Tile_X5Y6_FrameData_O[26] ,
    \Tile_X5Y6_FrameData_O[25] ,
    \Tile_X5Y6_FrameData_O[24] ,
    \Tile_X5Y6_FrameData_O[23] ,
    \Tile_X5Y6_FrameData_O[22] ,
    \Tile_X5Y6_FrameData_O[21] ,
    \Tile_X5Y6_FrameData_O[20] ,
    \Tile_X5Y6_FrameData_O[19] ,
    \Tile_X5Y6_FrameData_O[18] ,
    \Tile_X5Y6_FrameData_O[17] ,
    \Tile_X5Y6_FrameData_O[16] ,
    \Tile_X5Y6_FrameData_O[15] ,
    \Tile_X5Y6_FrameData_O[14] ,
    \Tile_X5Y6_FrameData_O[13] ,
    \Tile_X5Y6_FrameData_O[12] ,
    \Tile_X5Y6_FrameData_O[11] ,
    \Tile_X5Y6_FrameData_O[10] ,
    \Tile_X5Y6_FrameData_O[9] ,
    \Tile_X5Y6_FrameData_O[8] ,
    \Tile_X5Y6_FrameData_O[7] ,
    \Tile_X5Y6_FrameData_O[6] ,
    \Tile_X5Y6_FrameData_O[5] ,
    \Tile_X5Y6_FrameData_O[4] ,
    \Tile_X5Y6_FrameData_O[3] ,
    \Tile_X5Y6_FrameData_O[2] ,
    \Tile_X5Y6_FrameData_O[1] ,
    \Tile_X5Y6_FrameData_O[0] }),
    .FrameStrobe({\Tile_X5Y7_FrameStrobe_O[19] ,
    \Tile_X5Y7_FrameStrobe_O[18] ,
    \Tile_X5Y7_FrameStrobe_O[17] ,
    \Tile_X5Y7_FrameStrobe_O[16] ,
    \Tile_X5Y7_FrameStrobe_O[15] ,
    \Tile_X5Y7_FrameStrobe_O[14] ,
    \Tile_X5Y7_FrameStrobe_O[13] ,
    \Tile_X5Y7_FrameStrobe_O[12] ,
    \Tile_X5Y7_FrameStrobe_O[11] ,
    \Tile_X5Y7_FrameStrobe_O[10] ,
    \Tile_X5Y7_FrameStrobe_O[9] ,
    \Tile_X5Y7_FrameStrobe_O[8] ,
    \Tile_X5Y7_FrameStrobe_O[7] ,
    \Tile_X5Y7_FrameStrobe_O[6] ,
    \Tile_X5Y7_FrameStrobe_O[5] ,
    \Tile_X5Y7_FrameStrobe_O[4] ,
    \Tile_X5Y7_FrameStrobe_O[3] ,
    \Tile_X5Y7_FrameStrobe_O[2] ,
    \Tile_X5Y7_FrameStrobe_O[1] ,
    \Tile_X5Y7_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X5Y6_FrameStrobe_O[19] ,
    \Tile_X5Y6_FrameStrobe_O[18] ,
    \Tile_X5Y6_FrameStrobe_O[17] ,
    \Tile_X5Y6_FrameStrobe_O[16] ,
    \Tile_X5Y6_FrameStrobe_O[15] ,
    \Tile_X5Y6_FrameStrobe_O[14] ,
    \Tile_X5Y6_FrameStrobe_O[13] ,
    \Tile_X5Y6_FrameStrobe_O[12] ,
    \Tile_X5Y6_FrameStrobe_O[11] ,
    \Tile_X5Y6_FrameStrobe_O[10] ,
    \Tile_X5Y6_FrameStrobe_O[9] ,
    \Tile_X5Y6_FrameStrobe_O[8] ,
    \Tile_X5Y6_FrameStrobe_O[7] ,
    \Tile_X5Y6_FrameStrobe_O[6] ,
    \Tile_X5Y6_FrameStrobe_O[5] ,
    \Tile_X5Y6_FrameStrobe_O[4] ,
    \Tile_X5Y6_FrameStrobe_O[3] ,
    \Tile_X5Y6_FrameStrobe_O[2] ,
    \Tile_X5Y6_FrameStrobe_O[1] ,
    \Tile_X5Y6_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X5Y6_N1BEG[3] ,
    \Tile_X5Y6_N1BEG[2] ,
    \Tile_X5Y6_N1BEG[1] ,
    \Tile_X5Y6_N1BEG[0] }),
    .N1END({\Tile_X5Y7_N1BEG[3] ,
    \Tile_X5Y7_N1BEG[2] ,
    \Tile_X5Y7_N1BEG[1] ,
    \Tile_X5Y7_N1BEG[0] }),
    .N2BEG({\Tile_X5Y6_N2BEG[7] ,
    \Tile_X5Y6_N2BEG[6] ,
    \Tile_X5Y6_N2BEG[5] ,
    \Tile_X5Y6_N2BEG[4] ,
    \Tile_X5Y6_N2BEG[3] ,
    \Tile_X5Y6_N2BEG[2] ,
    \Tile_X5Y6_N2BEG[1] ,
    \Tile_X5Y6_N2BEG[0] }),
    .N2BEGb({\Tile_X5Y6_N2BEGb[7] ,
    \Tile_X5Y6_N2BEGb[6] ,
    \Tile_X5Y6_N2BEGb[5] ,
    \Tile_X5Y6_N2BEGb[4] ,
    \Tile_X5Y6_N2BEGb[3] ,
    \Tile_X5Y6_N2BEGb[2] ,
    \Tile_X5Y6_N2BEGb[1] ,
    \Tile_X5Y6_N2BEGb[0] }),
    .N2END({\Tile_X5Y7_N2BEGb[7] ,
    \Tile_X5Y7_N2BEGb[6] ,
    \Tile_X5Y7_N2BEGb[5] ,
    \Tile_X5Y7_N2BEGb[4] ,
    \Tile_X5Y7_N2BEGb[3] ,
    \Tile_X5Y7_N2BEGb[2] ,
    \Tile_X5Y7_N2BEGb[1] ,
    \Tile_X5Y7_N2BEGb[0] }),
    .N2MID({\Tile_X5Y7_N2BEG[7] ,
    \Tile_X5Y7_N2BEG[6] ,
    \Tile_X5Y7_N2BEG[5] ,
    \Tile_X5Y7_N2BEG[4] ,
    \Tile_X5Y7_N2BEG[3] ,
    \Tile_X5Y7_N2BEG[2] ,
    \Tile_X5Y7_N2BEG[1] ,
    \Tile_X5Y7_N2BEG[0] }),
    .N4BEG({\Tile_X5Y6_N4BEG[15] ,
    \Tile_X5Y6_N4BEG[14] ,
    \Tile_X5Y6_N4BEG[13] ,
    \Tile_X5Y6_N4BEG[12] ,
    \Tile_X5Y6_N4BEG[11] ,
    \Tile_X5Y6_N4BEG[10] ,
    \Tile_X5Y6_N4BEG[9] ,
    \Tile_X5Y6_N4BEG[8] ,
    \Tile_X5Y6_N4BEG[7] ,
    \Tile_X5Y6_N4BEG[6] ,
    \Tile_X5Y6_N4BEG[5] ,
    \Tile_X5Y6_N4BEG[4] ,
    \Tile_X5Y6_N4BEG[3] ,
    \Tile_X5Y6_N4BEG[2] ,
    \Tile_X5Y6_N4BEG[1] ,
    \Tile_X5Y6_N4BEG[0] }),
    .N4END({\Tile_X5Y7_N4BEG[15] ,
    \Tile_X5Y7_N4BEG[14] ,
    \Tile_X5Y7_N4BEG[13] ,
    \Tile_X5Y7_N4BEG[12] ,
    \Tile_X5Y7_N4BEG[11] ,
    \Tile_X5Y7_N4BEG[10] ,
    \Tile_X5Y7_N4BEG[9] ,
    \Tile_X5Y7_N4BEG[8] ,
    \Tile_X5Y7_N4BEG[7] ,
    \Tile_X5Y7_N4BEG[6] ,
    \Tile_X5Y7_N4BEG[5] ,
    \Tile_X5Y7_N4BEG[4] ,
    \Tile_X5Y7_N4BEG[3] ,
    \Tile_X5Y7_N4BEG[2] ,
    \Tile_X5Y7_N4BEG[1] ,
    \Tile_X5Y7_N4BEG[0] }),
    .S1BEG({\Tile_X5Y6_S1BEG[3] ,
    \Tile_X5Y6_S1BEG[2] ,
    \Tile_X5Y6_S1BEG[1] ,
    \Tile_X5Y6_S1BEG[0] }),
    .S1END({\Tile_X5Y5_S1BEG[3] ,
    \Tile_X5Y5_S1BEG[2] ,
    \Tile_X5Y5_S1BEG[1] ,
    \Tile_X5Y5_S1BEG[0] }),
    .S2BEG({\Tile_X5Y6_S2BEG[7] ,
    \Tile_X5Y6_S2BEG[6] ,
    \Tile_X5Y6_S2BEG[5] ,
    \Tile_X5Y6_S2BEG[4] ,
    \Tile_X5Y6_S2BEG[3] ,
    \Tile_X5Y6_S2BEG[2] ,
    \Tile_X5Y6_S2BEG[1] ,
    \Tile_X5Y6_S2BEG[0] }),
    .S2BEGb({\Tile_X5Y6_S2BEGb[7] ,
    \Tile_X5Y6_S2BEGb[6] ,
    \Tile_X5Y6_S2BEGb[5] ,
    \Tile_X5Y6_S2BEGb[4] ,
    \Tile_X5Y6_S2BEGb[3] ,
    \Tile_X5Y6_S2BEGb[2] ,
    \Tile_X5Y6_S2BEGb[1] ,
    \Tile_X5Y6_S2BEGb[0] }),
    .S2END({\Tile_X5Y5_S2BEGb[7] ,
    \Tile_X5Y5_S2BEGb[6] ,
    \Tile_X5Y5_S2BEGb[5] ,
    \Tile_X5Y5_S2BEGb[4] ,
    \Tile_X5Y5_S2BEGb[3] ,
    \Tile_X5Y5_S2BEGb[2] ,
    \Tile_X5Y5_S2BEGb[1] ,
    \Tile_X5Y5_S2BEGb[0] }),
    .S2MID({\Tile_X5Y5_S2BEG[7] ,
    \Tile_X5Y5_S2BEG[6] ,
    \Tile_X5Y5_S2BEG[5] ,
    \Tile_X5Y5_S2BEG[4] ,
    \Tile_X5Y5_S2BEG[3] ,
    \Tile_X5Y5_S2BEG[2] ,
    \Tile_X5Y5_S2BEG[1] ,
    \Tile_X5Y5_S2BEG[0] }),
    .S4BEG({\Tile_X5Y6_S4BEG[15] ,
    \Tile_X5Y6_S4BEG[14] ,
    \Tile_X5Y6_S4BEG[13] ,
    \Tile_X5Y6_S4BEG[12] ,
    \Tile_X5Y6_S4BEG[11] ,
    \Tile_X5Y6_S4BEG[10] ,
    \Tile_X5Y6_S4BEG[9] ,
    \Tile_X5Y6_S4BEG[8] ,
    \Tile_X5Y6_S4BEG[7] ,
    \Tile_X5Y6_S4BEG[6] ,
    \Tile_X5Y6_S4BEG[5] ,
    \Tile_X5Y6_S4BEG[4] ,
    \Tile_X5Y6_S4BEG[3] ,
    \Tile_X5Y6_S4BEG[2] ,
    \Tile_X5Y6_S4BEG[1] ,
    \Tile_X5Y6_S4BEG[0] }),
    .S4END({\Tile_X5Y5_S4BEG[15] ,
    \Tile_X5Y5_S4BEG[14] ,
    \Tile_X5Y5_S4BEG[13] ,
    \Tile_X5Y5_S4BEG[12] ,
    \Tile_X5Y5_S4BEG[11] ,
    \Tile_X5Y5_S4BEG[10] ,
    \Tile_X5Y5_S4BEG[9] ,
    \Tile_X5Y5_S4BEG[8] ,
    \Tile_X5Y5_S4BEG[7] ,
    \Tile_X5Y5_S4BEG[6] ,
    \Tile_X5Y5_S4BEG[5] ,
    \Tile_X5Y5_S4BEG[4] ,
    \Tile_X5Y5_S4BEG[3] ,
    \Tile_X5Y5_S4BEG[2] ,
    \Tile_X5Y5_S4BEG[1] ,
    \Tile_X5Y5_S4BEG[0] }),
    .W1BEG({\Tile_X5Y6_W1BEG[3] ,
    \Tile_X5Y6_W1BEG[2] ,
    \Tile_X5Y6_W1BEG[1] ,
    \Tile_X5Y6_W1BEG[0] }),
    .W2BEG({\Tile_X5Y6_W2BEG[7] ,
    \Tile_X5Y6_W2BEG[6] ,
    \Tile_X5Y6_W2BEG[5] ,
    \Tile_X5Y6_W2BEG[4] ,
    \Tile_X5Y6_W2BEG[3] ,
    \Tile_X5Y6_W2BEG[2] ,
    \Tile_X5Y6_W2BEG[1] ,
    \Tile_X5Y6_W2BEG[0] }),
    .W2BEGb({\Tile_X5Y6_W2BEGb[7] ,
    \Tile_X5Y6_W2BEGb[6] ,
    \Tile_X5Y6_W2BEGb[5] ,
    \Tile_X5Y6_W2BEGb[4] ,
    \Tile_X5Y6_W2BEGb[3] ,
    \Tile_X5Y6_W2BEGb[2] ,
    \Tile_X5Y6_W2BEGb[1] ,
    \Tile_X5Y6_W2BEGb[0] }),
    .W6BEG({\Tile_X5Y6_W6BEG[11] ,
    \Tile_X5Y6_W6BEG[10] ,
    \Tile_X5Y6_W6BEG[9] ,
    \Tile_X5Y6_W6BEG[8] ,
    \Tile_X5Y6_W6BEG[7] ,
    \Tile_X5Y6_W6BEG[6] ,
    \Tile_X5Y6_W6BEG[5] ,
    \Tile_X5Y6_W6BEG[4] ,
    \Tile_X5Y6_W6BEG[3] ,
    \Tile_X5Y6_W6BEG[2] ,
    \Tile_X5Y6_W6BEG[1] ,
    \Tile_X5Y6_W6BEG[0] }),
    .WW4BEG({\Tile_X5Y6_WW4BEG[15] ,
    \Tile_X5Y6_WW4BEG[14] ,
    \Tile_X5Y6_WW4BEG[13] ,
    \Tile_X5Y6_WW4BEG[12] ,
    \Tile_X5Y6_WW4BEG[11] ,
    \Tile_X5Y6_WW4BEG[10] ,
    \Tile_X5Y6_WW4BEG[9] ,
    \Tile_X5Y6_WW4BEG[8] ,
    \Tile_X5Y6_WW4BEG[7] ,
    \Tile_X5Y6_WW4BEG[6] ,
    \Tile_X5Y6_WW4BEG[5] ,
    \Tile_X5Y6_WW4BEG[4] ,
    \Tile_X5Y6_WW4BEG[3] ,
    \Tile_X5Y6_WW4BEG[2] ,
    \Tile_X5Y6_WW4BEG[1] ,
    \Tile_X5Y6_WW4BEG[0] }));
 E_TT_IF Tile_X5Y7_E_TT_IF (.CLK_TT_PROJECT(Tile_X5Y7_CLK_TT_PROJECT),
    .ENA_TT_PROJECT(Tile_X5Y7_ENA_TT_PROJECT),
    .RST_N_TT_PROJECT(Tile_X5Y7_RST_N_TT_PROJECT),
    .UIO_IN_TT_PROJECT0(Tile_X5Y7_UIO_IN_TT_PROJECT0),
    .UIO_IN_TT_PROJECT1(Tile_X5Y7_UIO_IN_TT_PROJECT1),
    .UIO_IN_TT_PROJECT2(Tile_X5Y7_UIO_IN_TT_PROJECT2),
    .UIO_IN_TT_PROJECT3(Tile_X5Y7_UIO_IN_TT_PROJECT3),
    .UIO_IN_TT_PROJECT4(Tile_X5Y7_UIO_IN_TT_PROJECT4),
    .UIO_IN_TT_PROJECT5(Tile_X5Y7_UIO_IN_TT_PROJECT5),
    .UIO_IN_TT_PROJECT6(Tile_X5Y7_UIO_IN_TT_PROJECT6),
    .UIO_IN_TT_PROJECT7(Tile_X5Y7_UIO_IN_TT_PROJECT7),
    .UIO_OE_TT_PROJECT0(Tile_X5Y7_UIO_OE_TT_PROJECT0),
    .UIO_OE_TT_PROJECT1(Tile_X5Y7_UIO_OE_TT_PROJECT1),
    .UIO_OE_TT_PROJECT2(Tile_X5Y7_UIO_OE_TT_PROJECT2),
    .UIO_OE_TT_PROJECT3(Tile_X5Y7_UIO_OE_TT_PROJECT3),
    .UIO_OE_TT_PROJECT4(Tile_X5Y7_UIO_OE_TT_PROJECT4),
    .UIO_OE_TT_PROJECT5(Tile_X5Y7_UIO_OE_TT_PROJECT5),
    .UIO_OE_TT_PROJECT6(Tile_X5Y7_UIO_OE_TT_PROJECT6),
    .UIO_OE_TT_PROJECT7(Tile_X5Y7_UIO_OE_TT_PROJECT7),
    .UIO_OUT_TT_PROJECT0(Tile_X5Y7_UIO_OUT_TT_PROJECT0),
    .UIO_OUT_TT_PROJECT1(Tile_X5Y7_UIO_OUT_TT_PROJECT1),
    .UIO_OUT_TT_PROJECT2(Tile_X5Y7_UIO_OUT_TT_PROJECT2),
    .UIO_OUT_TT_PROJECT3(Tile_X5Y7_UIO_OUT_TT_PROJECT3),
    .UIO_OUT_TT_PROJECT4(Tile_X5Y7_UIO_OUT_TT_PROJECT4),
    .UIO_OUT_TT_PROJECT5(Tile_X5Y7_UIO_OUT_TT_PROJECT5),
    .UIO_OUT_TT_PROJECT6(Tile_X5Y7_UIO_OUT_TT_PROJECT6),
    .UIO_OUT_TT_PROJECT7(Tile_X5Y7_UIO_OUT_TT_PROJECT7),
    .UI_IN_TT_PROJECT0(Tile_X5Y7_UI_IN_TT_PROJECT0),
    .UI_IN_TT_PROJECT1(Tile_X5Y7_UI_IN_TT_PROJECT1),
    .UI_IN_TT_PROJECT2(Tile_X5Y7_UI_IN_TT_PROJECT2),
    .UI_IN_TT_PROJECT3(Tile_X5Y7_UI_IN_TT_PROJECT3),
    .UI_IN_TT_PROJECT4(Tile_X5Y7_UI_IN_TT_PROJECT4),
    .UI_IN_TT_PROJECT5(Tile_X5Y7_UI_IN_TT_PROJECT5),
    .UI_IN_TT_PROJECT6(Tile_X5Y7_UI_IN_TT_PROJECT6),
    .UI_IN_TT_PROJECT7(Tile_X5Y7_UI_IN_TT_PROJECT7),
    .UO_OUT_TT_PROJECT0(Tile_X5Y7_UO_OUT_TT_PROJECT0),
    .UO_OUT_TT_PROJECT1(Tile_X5Y7_UO_OUT_TT_PROJECT1),
    .UO_OUT_TT_PROJECT2(Tile_X5Y7_UO_OUT_TT_PROJECT2),
    .UO_OUT_TT_PROJECT3(Tile_X5Y7_UO_OUT_TT_PROJECT3),
    .UO_OUT_TT_PROJECT4(Tile_X5Y7_UO_OUT_TT_PROJECT4),
    .UO_OUT_TT_PROJECT5(Tile_X5Y7_UO_OUT_TT_PROJECT5),
    .UO_OUT_TT_PROJECT6(Tile_X5Y7_UO_OUT_TT_PROJECT6),
    .UO_OUT_TT_PROJECT7(Tile_X5Y7_UO_OUT_TT_PROJECT7),
    .UserCLK(Tile_X5Y8_UserCLKo),
    .UserCLKo(Tile_X5Y7_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1END({\Tile_X4Y7_E1BEG[3] ,
    \Tile_X4Y7_E1BEG[2] ,
    \Tile_X4Y7_E1BEG[1] ,
    \Tile_X4Y7_E1BEG[0] }),
    .E2END({\Tile_X4Y7_E2BEGb[7] ,
    \Tile_X4Y7_E2BEGb[6] ,
    \Tile_X4Y7_E2BEGb[5] ,
    \Tile_X4Y7_E2BEGb[4] ,
    \Tile_X4Y7_E2BEGb[3] ,
    \Tile_X4Y7_E2BEGb[2] ,
    \Tile_X4Y7_E2BEGb[1] ,
    \Tile_X4Y7_E2BEGb[0] }),
    .E2MID({\Tile_X4Y7_E2BEG[7] ,
    \Tile_X4Y7_E2BEG[6] ,
    \Tile_X4Y7_E2BEG[5] ,
    \Tile_X4Y7_E2BEG[4] ,
    \Tile_X4Y7_E2BEG[3] ,
    \Tile_X4Y7_E2BEG[2] ,
    \Tile_X4Y7_E2BEG[1] ,
    \Tile_X4Y7_E2BEG[0] }),
    .E6END({\Tile_X4Y7_E6BEG[11] ,
    \Tile_X4Y7_E6BEG[10] ,
    \Tile_X4Y7_E6BEG[9] ,
    \Tile_X4Y7_E6BEG[8] ,
    \Tile_X4Y7_E6BEG[7] ,
    \Tile_X4Y7_E6BEG[6] ,
    \Tile_X4Y7_E6BEG[5] ,
    \Tile_X4Y7_E6BEG[4] ,
    \Tile_X4Y7_E6BEG[3] ,
    \Tile_X4Y7_E6BEG[2] ,
    \Tile_X4Y7_E6BEG[1] ,
    \Tile_X4Y7_E6BEG[0] }),
    .EE4END({\Tile_X4Y7_EE4BEG[15] ,
    \Tile_X4Y7_EE4BEG[14] ,
    \Tile_X4Y7_EE4BEG[13] ,
    \Tile_X4Y7_EE4BEG[12] ,
    \Tile_X4Y7_EE4BEG[11] ,
    \Tile_X4Y7_EE4BEG[10] ,
    \Tile_X4Y7_EE4BEG[9] ,
    \Tile_X4Y7_EE4BEG[8] ,
    \Tile_X4Y7_EE4BEG[7] ,
    \Tile_X4Y7_EE4BEG[6] ,
    \Tile_X4Y7_EE4BEG[5] ,
    \Tile_X4Y7_EE4BEG[4] ,
    \Tile_X4Y7_EE4BEG[3] ,
    \Tile_X4Y7_EE4BEG[2] ,
    \Tile_X4Y7_EE4BEG[1] ,
    \Tile_X4Y7_EE4BEG[0] }),
    .FrameData({\Tile_X4Y7_FrameData_O[31] ,
    \Tile_X4Y7_FrameData_O[30] ,
    \Tile_X4Y7_FrameData_O[29] ,
    \Tile_X4Y7_FrameData_O[28] ,
    \Tile_X4Y7_FrameData_O[27] ,
    \Tile_X4Y7_FrameData_O[26] ,
    \Tile_X4Y7_FrameData_O[25] ,
    \Tile_X4Y7_FrameData_O[24] ,
    \Tile_X4Y7_FrameData_O[23] ,
    \Tile_X4Y7_FrameData_O[22] ,
    \Tile_X4Y7_FrameData_O[21] ,
    \Tile_X4Y7_FrameData_O[20] ,
    \Tile_X4Y7_FrameData_O[19] ,
    \Tile_X4Y7_FrameData_O[18] ,
    \Tile_X4Y7_FrameData_O[17] ,
    \Tile_X4Y7_FrameData_O[16] ,
    \Tile_X4Y7_FrameData_O[15] ,
    \Tile_X4Y7_FrameData_O[14] ,
    \Tile_X4Y7_FrameData_O[13] ,
    \Tile_X4Y7_FrameData_O[12] ,
    \Tile_X4Y7_FrameData_O[11] ,
    \Tile_X4Y7_FrameData_O[10] ,
    \Tile_X4Y7_FrameData_O[9] ,
    \Tile_X4Y7_FrameData_O[8] ,
    \Tile_X4Y7_FrameData_O[7] ,
    \Tile_X4Y7_FrameData_O[6] ,
    \Tile_X4Y7_FrameData_O[5] ,
    \Tile_X4Y7_FrameData_O[4] ,
    \Tile_X4Y7_FrameData_O[3] ,
    \Tile_X4Y7_FrameData_O[2] ,
    \Tile_X4Y7_FrameData_O[1] ,
    \Tile_X4Y7_FrameData_O[0] }),
    .FrameData_O({\Tile_X5Y7_FrameData_O[31] ,
    \Tile_X5Y7_FrameData_O[30] ,
    \Tile_X5Y7_FrameData_O[29] ,
    \Tile_X5Y7_FrameData_O[28] ,
    \Tile_X5Y7_FrameData_O[27] ,
    \Tile_X5Y7_FrameData_O[26] ,
    \Tile_X5Y7_FrameData_O[25] ,
    \Tile_X5Y7_FrameData_O[24] ,
    \Tile_X5Y7_FrameData_O[23] ,
    \Tile_X5Y7_FrameData_O[22] ,
    \Tile_X5Y7_FrameData_O[21] ,
    \Tile_X5Y7_FrameData_O[20] ,
    \Tile_X5Y7_FrameData_O[19] ,
    \Tile_X5Y7_FrameData_O[18] ,
    \Tile_X5Y7_FrameData_O[17] ,
    \Tile_X5Y7_FrameData_O[16] ,
    \Tile_X5Y7_FrameData_O[15] ,
    \Tile_X5Y7_FrameData_O[14] ,
    \Tile_X5Y7_FrameData_O[13] ,
    \Tile_X5Y7_FrameData_O[12] ,
    \Tile_X5Y7_FrameData_O[11] ,
    \Tile_X5Y7_FrameData_O[10] ,
    \Tile_X5Y7_FrameData_O[9] ,
    \Tile_X5Y7_FrameData_O[8] ,
    \Tile_X5Y7_FrameData_O[7] ,
    \Tile_X5Y7_FrameData_O[6] ,
    \Tile_X5Y7_FrameData_O[5] ,
    \Tile_X5Y7_FrameData_O[4] ,
    \Tile_X5Y7_FrameData_O[3] ,
    \Tile_X5Y7_FrameData_O[2] ,
    \Tile_X5Y7_FrameData_O[1] ,
    \Tile_X5Y7_FrameData_O[0] }),
    .FrameStrobe({\Tile_X5Y8_FrameStrobe_O[19] ,
    \Tile_X5Y8_FrameStrobe_O[18] ,
    \Tile_X5Y8_FrameStrobe_O[17] ,
    \Tile_X5Y8_FrameStrobe_O[16] ,
    \Tile_X5Y8_FrameStrobe_O[15] ,
    \Tile_X5Y8_FrameStrobe_O[14] ,
    \Tile_X5Y8_FrameStrobe_O[13] ,
    \Tile_X5Y8_FrameStrobe_O[12] ,
    \Tile_X5Y8_FrameStrobe_O[11] ,
    \Tile_X5Y8_FrameStrobe_O[10] ,
    \Tile_X5Y8_FrameStrobe_O[9] ,
    \Tile_X5Y8_FrameStrobe_O[8] ,
    \Tile_X5Y8_FrameStrobe_O[7] ,
    \Tile_X5Y8_FrameStrobe_O[6] ,
    \Tile_X5Y8_FrameStrobe_O[5] ,
    \Tile_X5Y8_FrameStrobe_O[4] ,
    \Tile_X5Y8_FrameStrobe_O[3] ,
    \Tile_X5Y8_FrameStrobe_O[2] ,
    \Tile_X5Y8_FrameStrobe_O[1] ,
    \Tile_X5Y8_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X5Y7_FrameStrobe_O[19] ,
    \Tile_X5Y7_FrameStrobe_O[18] ,
    \Tile_X5Y7_FrameStrobe_O[17] ,
    \Tile_X5Y7_FrameStrobe_O[16] ,
    \Tile_X5Y7_FrameStrobe_O[15] ,
    \Tile_X5Y7_FrameStrobe_O[14] ,
    \Tile_X5Y7_FrameStrobe_O[13] ,
    \Tile_X5Y7_FrameStrobe_O[12] ,
    \Tile_X5Y7_FrameStrobe_O[11] ,
    \Tile_X5Y7_FrameStrobe_O[10] ,
    \Tile_X5Y7_FrameStrobe_O[9] ,
    \Tile_X5Y7_FrameStrobe_O[8] ,
    \Tile_X5Y7_FrameStrobe_O[7] ,
    \Tile_X5Y7_FrameStrobe_O[6] ,
    \Tile_X5Y7_FrameStrobe_O[5] ,
    \Tile_X5Y7_FrameStrobe_O[4] ,
    \Tile_X5Y7_FrameStrobe_O[3] ,
    \Tile_X5Y7_FrameStrobe_O[2] ,
    \Tile_X5Y7_FrameStrobe_O[1] ,
    \Tile_X5Y7_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X5Y7_N1BEG[3] ,
    \Tile_X5Y7_N1BEG[2] ,
    \Tile_X5Y7_N1BEG[1] ,
    \Tile_X5Y7_N1BEG[0] }),
    .N1END({\Tile_X5Y8_N1BEG[3] ,
    \Tile_X5Y8_N1BEG[2] ,
    \Tile_X5Y8_N1BEG[1] ,
    \Tile_X5Y8_N1BEG[0] }),
    .N2BEG({\Tile_X5Y7_N2BEG[7] ,
    \Tile_X5Y7_N2BEG[6] ,
    \Tile_X5Y7_N2BEG[5] ,
    \Tile_X5Y7_N2BEG[4] ,
    \Tile_X5Y7_N2BEG[3] ,
    \Tile_X5Y7_N2BEG[2] ,
    \Tile_X5Y7_N2BEG[1] ,
    \Tile_X5Y7_N2BEG[0] }),
    .N2BEGb({\Tile_X5Y7_N2BEGb[7] ,
    \Tile_X5Y7_N2BEGb[6] ,
    \Tile_X5Y7_N2BEGb[5] ,
    \Tile_X5Y7_N2BEGb[4] ,
    \Tile_X5Y7_N2BEGb[3] ,
    \Tile_X5Y7_N2BEGb[2] ,
    \Tile_X5Y7_N2BEGb[1] ,
    \Tile_X5Y7_N2BEGb[0] }),
    .N2END({\Tile_X5Y8_N2BEGb[7] ,
    \Tile_X5Y8_N2BEGb[6] ,
    \Tile_X5Y8_N2BEGb[5] ,
    \Tile_X5Y8_N2BEGb[4] ,
    \Tile_X5Y8_N2BEGb[3] ,
    \Tile_X5Y8_N2BEGb[2] ,
    \Tile_X5Y8_N2BEGb[1] ,
    \Tile_X5Y8_N2BEGb[0] }),
    .N2MID({\Tile_X5Y8_N2BEG[7] ,
    \Tile_X5Y8_N2BEG[6] ,
    \Tile_X5Y8_N2BEG[5] ,
    \Tile_X5Y8_N2BEG[4] ,
    \Tile_X5Y8_N2BEG[3] ,
    \Tile_X5Y8_N2BEG[2] ,
    \Tile_X5Y8_N2BEG[1] ,
    \Tile_X5Y8_N2BEG[0] }),
    .N4BEG({\Tile_X5Y7_N4BEG[15] ,
    \Tile_X5Y7_N4BEG[14] ,
    \Tile_X5Y7_N4BEG[13] ,
    \Tile_X5Y7_N4BEG[12] ,
    \Tile_X5Y7_N4BEG[11] ,
    \Tile_X5Y7_N4BEG[10] ,
    \Tile_X5Y7_N4BEG[9] ,
    \Tile_X5Y7_N4BEG[8] ,
    \Tile_X5Y7_N4BEG[7] ,
    \Tile_X5Y7_N4BEG[6] ,
    \Tile_X5Y7_N4BEG[5] ,
    \Tile_X5Y7_N4BEG[4] ,
    \Tile_X5Y7_N4BEG[3] ,
    \Tile_X5Y7_N4BEG[2] ,
    \Tile_X5Y7_N4BEG[1] ,
    \Tile_X5Y7_N4BEG[0] }),
    .N4END({\Tile_X5Y8_N4BEG[15] ,
    \Tile_X5Y8_N4BEG[14] ,
    \Tile_X5Y8_N4BEG[13] ,
    \Tile_X5Y8_N4BEG[12] ,
    \Tile_X5Y8_N4BEG[11] ,
    \Tile_X5Y8_N4BEG[10] ,
    \Tile_X5Y8_N4BEG[9] ,
    \Tile_X5Y8_N4BEG[8] ,
    \Tile_X5Y8_N4BEG[7] ,
    \Tile_X5Y8_N4BEG[6] ,
    \Tile_X5Y8_N4BEG[5] ,
    \Tile_X5Y8_N4BEG[4] ,
    \Tile_X5Y8_N4BEG[3] ,
    \Tile_X5Y8_N4BEG[2] ,
    \Tile_X5Y8_N4BEG[1] ,
    \Tile_X5Y8_N4BEG[0] }),
    .S1BEG({\Tile_X5Y7_S1BEG[3] ,
    \Tile_X5Y7_S1BEG[2] ,
    \Tile_X5Y7_S1BEG[1] ,
    \Tile_X5Y7_S1BEG[0] }),
    .S1END({\Tile_X5Y6_S1BEG[3] ,
    \Tile_X5Y6_S1BEG[2] ,
    \Tile_X5Y6_S1BEG[1] ,
    \Tile_X5Y6_S1BEG[0] }),
    .S2BEG({\Tile_X5Y7_S2BEG[7] ,
    \Tile_X5Y7_S2BEG[6] ,
    \Tile_X5Y7_S2BEG[5] ,
    \Tile_X5Y7_S2BEG[4] ,
    \Tile_X5Y7_S2BEG[3] ,
    \Tile_X5Y7_S2BEG[2] ,
    \Tile_X5Y7_S2BEG[1] ,
    \Tile_X5Y7_S2BEG[0] }),
    .S2BEGb({\Tile_X5Y7_S2BEGb[7] ,
    \Tile_X5Y7_S2BEGb[6] ,
    \Tile_X5Y7_S2BEGb[5] ,
    \Tile_X5Y7_S2BEGb[4] ,
    \Tile_X5Y7_S2BEGb[3] ,
    \Tile_X5Y7_S2BEGb[2] ,
    \Tile_X5Y7_S2BEGb[1] ,
    \Tile_X5Y7_S2BEGb[0] }),
    .S2END({\Tile_X5Y6_S2BEGb[7] ,
    \Tile_X5Y6_S2BEGb[6] ,
    \Tile_X5Y6_S2BEGb[5] ,
    \Tile_X5Y6_S2BEGb[4] ,
    \Tile_X5Y6_S2BEGb[3] ,
    \Tile_X5Y6_S2BEGb[2] ,
    \Tile_X5Y6_S2BEGb[1] ,
    \Tile_X5Y6_S2BEGb[0] }),
    .S2MID({\Tile_X5Y6_S2BEG[7] ,
    \Tile_X5Y6_S2BEG[6] ,
    \Tile_X5Y6_S2BEG[5] ,
    \Tile_X5Y6_S2BEG[4] ,
    \Tile_X5Y6_S2BEG[3] ,
    \Tile_X5Y6_S2BEG[2] ,
    \Tile_X5Y6_S2BEG[1] ,
    \Tile_X5Y6_S2BEG[0] }),
    .S4BEG({\Tile_X5Y7_S4BEG[15] ,
    \Tile_X5Y7_S4BEG[14] ,
    \Tile_X5Y7_S4BEG[13] ,
    \Tile_X5Y7_S4BEG[12] ,
    \Tile_X5Y7_S4BEG[11] ,
    \Tile_X5Y7_S4BEG[10] ,
    \Tile_X5Y7_S4BEG[9] ,
    \Tile_X5Y7_S4BEG[8] ,
    \Tile_X5Y7_S4BEG[7] ,
    \Tile_X5Y7_S4BEG[6] ,
    \Tile_X5Y7_S4BEG[5] ,
    \Tile_X5Y7_S4BEG[4] ,
    \Tile_X5Y7_S4BEG[3] ,
    \Tile_X5Y7_S4BEG[2] ,
    \Tile_X5Y7_S4BEG[1] ,
    \Tile_X5Y7_S4BEG[0] }),
    .S4END({\Tile_X5Y6_S4BEG[15] ,
    \Tile_X5Y6_S4BEG[14] ,
    \Tile_X5Y6_S4BEG[13] ,
    \Tile_X5Y6_S4BEG[12] ,
    \Tile_X5Y6_S4BEG[11] ,
    \Tile_X5Y6_S4BEG[10] ,
    \Tile_X5Y6_S4BEG[9] ,
    \Tile_X5Y6_S4BEG[8] ,
    \Tile_X5Y6_S4BEG[7] ,
    \Tile_X5Y6_S4BEG[6] ,
    \Tile_X5Y6_S4BEG[5] ,
    \Tile_X5Y6_S4BEG[4] ,
    \Tile_X5Y6_S4BEG[3] ,
    \Tile_X5Y6_S4BEG[2] ,
    \Tile_X5Y6_S4BEG[1] ,
    \Tile_X5Y6_S4BEG[0] }),
    .W1BEG({\Tile_X5Y7_W1BEG[3] ,
    \Tile_X5Y7_W1BEG[2] ,
    \Tile_X5Y7_W1BEG[1] ,
    \Tile_X5Y7_W1BEG[0] }),
    .W2BEG({\Tile_X5Y7_W2BEG[7] ,
    \Tile_X5Y7_W2BEG[6] ,
    \Tile_X5Y7_W2BEG[5] ,
    \Tile_X5Y7_W2BEG[4] ,
    \Tile_X5Y7_W2BEG[3] ,
    \Tile_X5Y7_W2BEG[2] ,
    \Tile_X5Y7_W2BEG[1] ,
    \Tile_X5Y7_W2BEG[0] }),
    .W2BEGb({\Tile_X5Y7_W2BEGb[7] ,
    \Tile_X5Y7_W2BEGb[6] ,
    \Tile_X5Y7_W2BEGb[5] ,
    \Tile_X5Y7_W2BEGb[4] ,
    \Tile_X5Y7_W2BEGb[3] ,
    \Tile_X5Y7_W2BEGb[2] ,
    \Tile_X5Y7_W2BEGb[1] ,
    \Tile_X5Y7_W2BEGb[0] }),
    .W6BEG({\Tile_X5Y7_W6BEG[11] ,
    \Tile_X5Y7_W6BEG[10] ,
    \Tile_X5Y7_W6BEG[9] ,
    \Tile_X5Y7_W6BEG[8] ,
    \Tile_X5Y7_W6BEG[7] ,
    \Tile_X5Y7_W6BEG[6] ,
    \Tile_X5Y7_W6BEG[5] ,
    \Tile_X5Y7_W6BEG[4] ,
    \Tile_X5Y7_W6BEG[3] ,
    \Tile_X5Y7_W6BEG[2] ,
    \Tile_X5Y7_W6BEG[1] ,
    \Tile_X5Y7_W6BEG[0] }),
    .WW4BEG({\Tile_X5Y7_WW4BEG[15] ,
    \Tile_X5Y7_WW4BEG[14] ,
    \Tile_X5Y7_WW4BEG[13] ,
    \Tile_X5Y7_WW4BEG[12] ,
    \Tile_X5Y7_WW4BEG[11] ,
    \Tile_X5Y7_WW4BEG[10] ,
    \Tile_X5Y7_WW4BEG[9] ,
    \Tile_X5Y7_WW4BEG[8] ,
    \Tile_X5Y7_WW4BEG[7] ,
    \Tile_X5Y7_WW4BEG[6] ,
    \Tile_X5Y7_WW4BEG[5] ,
    \Tile_X5Y7_WW4BEG[4] ,
    \Tile_X5Y7_WW4BEG[3] ,
    \Tile_X5Y7_WW4BEG[2] ,
    \Tile_X5Y7_WW4BEG[1] ,
    \Tile_X5Y7_WW4BEG[0] }));
 E_TT_IF Tile_X5Y8_E_TT_IF (.CLK_TT_PROJECT(Tile_X5Y8_CLK_TT_PROJECT),
    .ENA_TT_PROJECT(Tile_X5Y8_ENA_TT_PROJECT),
    .RST_N_TT_PROJECT(Tile_X5Y8_RST_N_TT_PROJECT),
    .UIO_IN_TT_PROJECT0(Tile_X5Y8_UIO_IN_TT_PROJECT0),
    .UIO_IN_TT_PROJECT1(Tile_X5Y8_UIO_IN_TT_PROJECT1),
    .UIO_IN_TT_PROJECT2(Tile_X5Y8_UIO_IN_TT_PROJECT2),
    .UIO_IN_TT_PROJECT3(Tile_X5Y8_UIO_IN_TT_PROJECT3),
    .UIO_IN_TT_PROJECT4(Tile_X5Y8_UIO_IN_TT_PROJECT4),
    .UIO_IN_TT_PROJECT5(Tile_X5Y8_UIO_IN_TT_PROJECT5),
    .UIO_IN_TT_PROJECT6(Tile_X5Y8_UIO_IN_TT_PROJECT6),
    .UIO_IN_TT_PROJECT7(Tile_X5Y8_UIO_IN_TT_PROJECT7),
    .UIO_OE_TT_PROJECT0(Tile_X5Y8_UIO_OE_TT_PROJECT0),
    .UIO_OE_TT_PROJECT1(Tile_X5Y8_UIO_OE_TT_PROJECT1),
    .UIO_OE_TT_PROJECT2(Tile_X5Y8_UIO_OE_TT_PROJECT2),
    .UIO_OE_TT_PROJECT3(Tile_X5Y8_UIO_OE_TT_PROJECT3),
    .UIO_OE_TT_PROJECT4(Tile_X5Y8_UIO_OE_TT_PROJECT4),
    .UIO_OE_TT_PROJECT5(Tile_X5Y8_UIO_OE_TT_PROJECT5),
    .UIO_OE_TT_PROJECT6(Tile_X5Y8_UIO_OE_TT_PROJECT6),
    .UIO_OE_TT_PROJECT7(Tile_X5Y8_UIO_OE_TT_PROJECT7),
    .UIO_OUT_TT_PROJECT0(Tile_X5Y8_UIO_OUT_TT_PROJECT0),
    .UIO_OUT_TT_PROJECT1(Tile_X5Y8_UIO_OUT_TT_PROJECT1),
    .UIO_OUT_TT_PROJECT2(Tile_X5Y8_UIO_OUT_TT_PROJECT2),
    .UIO_OUT_TT_PROJECT3(Tile_X5Y8_UIO_OUT_TT_PROJECT3),
    .UIO_OUT_TT_PROJECT4(Tile_X5Y8_UIO_OUT_TT_PROJECT4),
    .UIO_OUT_TT_PROJECT5(Tile_X5Y8_UIO_OUT_TT_PROJECT5),
    .UIO_OUT_TT_PROJECT6(Tile_X5Y8_UIO_OUT_TT_PROJECT6),
    .UIO_OUT_TT_PROJECT7(Tile_X5Y8_UIO_OUT_TT_PROJECT7),
    .UI_IN_TT_PROJECT0(Tile_X5Y8_UI_IN_TT_PROJECT0),
    .UI_IN_TT_PROJECT1(Tile_X5Y8_UI_IN_TT_PROJECT1),
    .UI_IN_TT_PROJECT2(Tile_X5Y8_UI_IN_TT_PROJECT2),
    .UI_IN_TT_PROJECT3(Tile_X5Y8_UI_IN_TT_PROJECT3),
    .UI_IN_TT_PROJECT4(Tile_X5Y8_UI_IN_TT_PROJECT4),
    .UI_IN_TT_PROJECT5(Tile_X5Y8_UI_IN_TT_PROJECT5),
    .UI_IN_TT_PROJECT6(Tile_X5Y8_UI_IN_TT_PROJECT6),
    .UI_IN_TT_PROJECT7(Tile_X5Y8_UI_IN_TT_PROJECT7),
    .UO_OUT_TT_PROJECT0(Tile_X5Y8_UO_OUT_TT_PROJECT0),
    .UO_OUT_TT_PROJECT1(Tile_X5Y8_UO_OUT_TT_PROJECT1),
    .UO_OUT_TT_PROJECT2(Tile_X5Y8_UO_OUT_TT_PROJECT2),
    .UO_OUT_TT_PROJECT3(Tile_X5Y8_UO_OUT_TT_PROJECT3),
    .UO_OUT_TT_PROJECT4(Tile_X5Y8_UO_OUT_TT_PROJECT4),
    .UO_OUT_TT_PROJECT5(Tile_X5Y8_UO_OUT_TT_PROJECT5),
    .UO_OUT_TT_PROJECT6(Tile_X5Y8_UO_OUT_TT_PROJECT6),
    .UO_OUT_TT_PROJECT7(Tile_X5Y8_UO_OUT_TT_PROJECT7),
    .UserCLK(Tile_X5Y9_UserCLKo),
    .UserCLKo(Tile_X5Y8_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1END({\Tile_X4Y8_E1BEG[3] ,
    \Tile_X4Y8_E1BEG[2] ,
    \Tile_X4Y8_E1BEG[1] ,
    \Tile_X4Y8_E1BEG[0] }),
    .E2END({\Tile_X4Y8_E2BEGb[7] ,
    \Tile_X4Y8_E2BEGb[6] ,
    \Tile_X4Y8_E2BEGb[5] ,
    \Tile_X4Y8_E2BEGb[4] ,
    \Tile_X4Y8_E2BEGb[3] ,
    \Tile_X4Y8_E2BEGb[2] ,
    \Tile_X4Y8_E2BEGb[1] ,
    \Tile_X4Y8_E2BEGb[0] }),
    .E2MID({\Tile_X4Y8_E2BEG[7] ,
    \Tile_X4Y8_E2BEG[6] ,
    \Tile_X4Y8_E2BEG[5] ,
    \Tile_X4Y8_E2BEG[4] ,
    \Tile_X4Y8_E2BEG[3] ,
    \Tile_X4Y8_E2BEG[2] ,
    \Tile_X4Y8_E2BEG[1] ,
    \Tile_X4Y8_E2BEG[0] }),
    .E6END({\Tile_X4Y8_E6BEG[11] ,
    \Tile_X4Y8_E6BEG[10] ,
    \Tile_X4Y8_E6BEG[9] ,
    \Tile_X4Y8_E6BEG[8] ,
    \Tile_X4Y8_E6BEG[7] ,
    \Tile_X4Y8_E6BEG[6] ,
    \Tile_X4Y8_E6BEG[5] ,
    \Tile_X4Y8_E6BEG[4] ,
    \Tile_X4Y8_E6BEG[3] ,
    \Tile_X4Y8_E6BEG[2] ,
    \Tile_X4Y8_E6BEG[1] ,
    \Tile_X4Y8_E6BEG[0] }),
    .EE4END({\Tile_X4Y8_EE4BEG[15] ,
    \Tile_X4Y8_EE4BEG[14] ,
    \Tile_X4Y8_EE4BEG[13] ,
    \Tile_X4Y8_EE4BEG[12] ,
    \Tile_X4Y8_EE4BEG[11] ,
    \Tile_X4Y8_EE4BEG[10] ,
    \Tile_X4Y8_EE4BEG[9] ,
    \Tile_X4Y8_EE4BEG[8] ,
    \Tile_X4Y8_EE4BEG[7] ,
    \Tile_X4Y8_EE4BEG[6] ,
    \Tile_X4Y8_EE4BEG[5] ,
    \Tile_X4Y8_EE4BEG[4] ,
    \Tile_X4Y8_EE4BEG[3] ,
    \Tile_X4Y8_EE4BEG[2] ,
    \Tile_X4Y8_EE4BEG[1] ,
    \Tile_X4Y8_EE4BEG[0] }),
    .FrameData({\Tile_X4Y8_FrameData_O[31] ,
    \Tile_X4Y8_FrameData_O[30] ,
    \Tile_X4Y8_FrameData_O[29] ,
    \Tile_X4Y8_FrameData_O[28] ,
    \Tile_X4Y8_FrameData_O[27] ,
    \Tile_X4Y8_FrameData_O[26] ,
    \Tile_X4Y8_FrameData_O[25] ,
    \Tile_X4Y8_FrameData_O[24] ,
    \Tile_X4Y8_FrameData_O[23] ,
    \Tile_X4Y8_FrameData_O[22] ,
    \Tile_X4Y8_FrameData_O[21] ,
    \Tile_X4Y8_FrameData_O[20] ,
    \Tile_X4Y8_FrameData_O[19] ,
    \Tile_X4Y8_FrameData_O[18] ,
    \Tile_X4Y8_FrameData_O[17] ,
    \Tile_X4Y8_FrameData_O[16] ,
    \Tile_X4Y8_FrameData_O[15] ,
    \Tile_X4Y8_FrameData_O[14] ,
    \Tile_X4Y8_FrameData_O[13] ,
    \Tile_X4Y8_FrameData_O[12] ,
    \Tile_X4Y8_FrameData_O[11] ,
    \Tile_X4Y8_FrameData_O[10] ,
    \Tile_X4Y8_FrameData_O[9] ,
    \Tile_X4Y8_FrameData_O[8] ,
    \Tile_X4Y8_FrameData_O[7] ,
    \Tile_X4Y8_FrameData_O[6] ,
    \Tile_X4Y8_FrameData_O[5] ,
    \Tile_X4Y8_FrameData_O[4] ,
    \Tile_X4Y8_FrameData_O[3] ,
    \Tile_X4Y8_FrameData_O[2] ,
    \Tile_X4Y8_FrameData_O[1] ,
    \Tile_X4Y8_FrameData_O[0] }),
    .FrameData_O({\Tile_X5Y8_FrameData_O[31] ,
    \Tile_X5Y8_FrameData_O[30] ,
    \Tile_X5Y8_FrameData_O[29] ,
    \Tile_X5Y8_FrameData_O[28] ,
    \Tile_X5Y8_FrameData_O[27] ,
    \Tile_X5Y8_FrameData_O[26] ,
    \Tile_X5Y8_FrameData_O[25] ,
    \Tile_X5Y8_FrameData_O[24] ,
    \Tile_X5Y8_FrameData_O[23] ,
    \Tile_X5Y8_FrameData_O[22] ,
    \Tile_X5Y8_FrameData_O[21] ,
    \Tile_X5Y8_FrameData_O[20] ,
    \Tile_X5Y8_FrameData_O[19] ,
    \Tile_X5Y8_FrameData_O[18] ,
    \Tile_X5Y8_FrameData_O[17] ,
    \Tile_X5Y8_FrameData_O[16] ,
    \Tile_X5Y8_FrameData_O[15] ,
    \Tile_X5Y8_FrameData_O[14] ,
    \Tile_X5Y8_FrameData_O[13] ,
    \Tile_X5Y8_FrameData_O[12] ,
    \Tile_X5Y8_FrameData_O[11] ,
    \Tile_X5Y8_FrameData_O[10] ,
    \Tile_X5Y8_FrameData_O[9] ,
    \Tile_X5Y8_FrameData_O[8] ,
    \Tile_X5Y8_FrameData_O[7] ,
    \Tile_X5Y8_FrameData_O[6] ,
    \Tile_X5Y8_FrameData_O[5] ,
    \Tile_X5Y8_FrameData_O[4] ,
    \Tile_X5Y8_FrameData_O[3] ,
    \Tile_X5Y8_FrameData_O[2] ,
    \Tile_X5Y8_FrameData_O[1] ,
    \Tile_X5Y8_FrameData_O[0] }),
    .FrameStrobe({\Tile_X5Y9_FrameStrobe_O[19] ,
    \Tile_X5Y9_FrameStrobe_O[18] ,
    \Tile_X5Y9_FrameStrobe_O[17] ,
    \Tile_X5Y9_FrameStrobe_O[16] ,
    \Tile_X5Y9_FrameStrobe_O[15] ,
    \Tile_X5Y9_FrameStrobe_O[14] ,
    \Tile_X5Y9_FrameStrobe_O[13] ,
    \Tile_X5Y9_FrameStrobe_O[12] ,
    \Tile_X5Y9_FrameStrobe_O[11] ,
    \Tile_X5Y9_FrameStrobe_O[10] ,
    \Tile_X5Y9_FrameStrobe_O[9] ,
    \Tile_X5Y9_FrameStrobe_O[8] ,
    \Tile_X5Y9_FrameStrobe_O[7] ,
    \Tile_X5Y9_FrameStrobe_O[6] ,
    \Tile_X5Y9_FrameStrobe_O[5] ,
    \Tile_X5Y9_FrameStrobe_O[4] ,
    \Tile_X5Y9_FrameStrobe_O[3] ,
    \Tile_X5Y9_FrameStrobe_O[2] ,
    \Tile_X5Y9_FrameStrobe_O[1] ,
    \Tile_X5Y9_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X5Y8_FrameStrobe_O[19] ,
    \Tile_X5Y8_FrameStrobe_O[18] ,
    \Tile_X5Y8_FrameStrobe_O[17] ,
    \Tile_X5Y8_FrameStrobe_O[16] ,
    \Tile_X5Y8_FrameStrobe_O[15] ,
    \Tile_X5Y8_FrameStrobe_O[14] ,
    \Tile_X5Y8_FrameStrobe_O[13] ,
    \Tile_X5Y8_FrameStrobe_O[12] ,
    \Tile_X5Y8_FrameStrobe_O[11] ,
    \Tile_X5Y8_FrameStrobe_O[10] ,
    \Tile_X5Y8_FrameStrobe_O[9] ,
    \Tile_X5Y8_FrameStrobe_O[8] ,
    \Tile_X5Y8_FrameStrobe_O[7] ,
    \Tile_X5Y8_FrameStrobe_O[6] ,
    \Tile_X5Y8_FrameStrobe_O[5] ,
    \Tile_X5Y8_FrameStrobe_O[4] ,
    \Tile_X5Y8_FrameStrobe_O[3] ,
    \Tile_X5Y8_FrameStrobe_O[2] ,
    \Tile_X5Y8_FrameStrobe_O[1] ,
    \Tile_X5Y8_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X5Y8_N1BEG[3] ,
    \Tile_X5Y8_N1BEG[2] ,
    \Tile_X5Y8_N1BEG[1] ,
    \Tile_X5Y8_N1BEG[0] }),
    .N1END({\Tile_X5Y9_N1BEG[3] ,
    \Tile_X5Y9_N1BEG[2] ,
    \Tile_X5Y9_N1BEG[1] ,
    \Tile_X5Y9_N1BEG[0] }),
    .N2BEG({\Tile_X5Y8_N2BEG[7] ,
    \Tile_X5Y8_N2BEG[6] ,
    \Tile_X5Y8_N2BEG[5] ,
    \Tile_X5Y8_N2BEG[4] ,
    \Tile_X5Y8_N2BEG[3] ,
    \Tile_X5Y8_N2BEG[2] ,
    \Tile_X5Y8_N2BEG[1] ,
    \Tile_X5Y8_N2BEG[0] }),
    .N2BEGb({\Tile_X5Y8_N2BEGb[7] ,
    \Tile_X5Y8_N2BEGb[6] ,
    \Tile_X5Y8_N2BEGb[5] ,
    \Tile_X5Y8_N2BEGb[4] ,
    \Tile_X5Y8_N2BEGb[3] ,
    \Tile_X5Y8_N2BEGb[2] ,
    \Tile_X5Y8_N2BEGb[1] ,
    \Tile_X5Y8_N2BEGb[0] }),
    .N2END({\Tile_X5Y9_N2BEGb[7] ,
    \Tile_X5Y9_N2BEGb[6] ,
    \Tile_X5Y9_N2BEGb[5] ,
    \Tile_X5Y9_N2BEGb[4] ,
    \Tile_X5Y9_N2BEGb[3] ,
    \Tile_X5Y9_N2BEGb[2] ,
    \Tile_X5Y9_N2BEGb[1] ,
    \Tile_X5Y9_N2BEGb[0] }),
    .N2MID({\Tile_X5Y9_N2BEG[7] ,
    \Tile_X5Y9_N2BEG[6] ,
    \Tile_X5Y9_N2BEG[5] ,
    \Tile_X5Y9_N2BEG[4] ,
    \Tile_X5Y9_N2BEG[3] ,
    \Tile_X5Y9_N2BEG[2] ,
    \Tile_X5Y9_N2BEG[1] ,
    \Tile_X5Y9_N2BEG[0] }),
    .N4BEG({\Tile_X5Y8_N4BEG[15] ,
    \Tile_X5Y8_N4BEG[14] ,
    \Tile_X5Y8_N4BEG[13] ,
    \Tile_X5Y8_N4BEG[12] ,
    \Tile_X5Y8_N4BEG[11] ,
    \Tile_X5Y8_N4BEG[10] ,
    \Tile_X5Y8_N4BEG[9] ,
    \Tile_X5Y8_N4BEG[8] ,
    \Tile_X5Y8_N4BEG[7] ,
    \Tile_X5Y8_N4BEG[6] ,
    \Tile_X5Y8_N4BEG[5] ,
    \Tile_X5Y8_N4BEG[4] ,
    \Tile_X5Y8_N4BEG[3] ,
    \Tile_X5Y8_N4BEG[2] ,
    \Tile_X5Y8_N4BEG[1] ,
    \Tile_X5Y8_N4BEG[0] }),
    .N4END({\Tile_X5Y9_N4BEG[15] ,
    \Tile_X5Y9_N4BEG[14] ,
    \Tile_X5Y9_N4BEG[13] ,
    \Tile_X5Y9_N4BEG[12] ,
    \Tile_X5Y9_N4BEG[11] ,
    \Tile_X5Y9_N4BEG[10] ,
    \Tile_X5Y9_N4BEG[9] ,
    \Tile_X5Y9_N4BEG[8] ,
    \Tile_X5Y9_N4BEG[7] ,
    \Tile_X5Y9_N4BEG[6] ,
    \Tile_X5Y9_N4BEG[5] ,
    \Tile_X5Y9_N4BEG[4] ,
    \Tile_X5Y9_N4BEG[3] ,
    \Tile_X5Y9_N4BEG[2] ,
    \Tile_X5Y9_N4BEG[1] ,
    \Tile_X5Y9_N4BEG[0] }),
    .S1BEG({\Tile_X5Y8_S1BEG[3] ,
    \Tile_X5Y8_S1BEG[2] ,
    \Tile_X5Y8_S1BEG[1] ,
    \Tile_X5Y8_S1BEG[0] }),
    .S1END({\Tile_X5Y7_S1BEG[3] ,
    \Tile_X5Y7_S1BEG[2] ,
    \Tile_X5Y7_S1BEG[1] ,
    \Tile_X5Y7_S1BEG[0] }),
    .S2BEG({\Tile_X5Y8_S2BEG[7] ,
    \Tile_X5Y8_S2BEG[6] ,
    \Tile_X5Y8_S2BEG[5] ,
    \Tile_X5Y8_S2BEG[4] ,
    \Tile_X5Y8_S2BEG[3] ,
    \Tile_X5Y8_S2BEG[2] ,
    \Tile_X5Y8_S2BEG[1] ,
    \Tile_X5Y8_S2BEG[0] }),
    .S2BEGb({\Tile_X5Y8_S2BEGb[7] ,
    \Tile_X5Y8_S2BEGb[6] ,
    \Tile_X5Y8_S2BEGb[5] ,
    \Tile_X5Y8_S2BEGb[4] ,
    \Tile_X5Y8_S2BEGb[3] ,
    \Tile_X5Y8_S2BEGb[2] ,
    \Tile_X5Y8_S2BEGb[1] ,
    \Tile_X5Y8_S2BEGb[0] }),
    .S2END({\Tile_X5Y7_S2BEGb[7] ,
    \Tile_X5Y7_S2BEGb[6] ,
    \Tile_X5Y7_S2BEGb[5] ,
    \Tile_X5Y7_S2BEGb[4] ,
    \Tile_X5Y7_S2BEGb[3] ,
    \Tile_X5Y7_S2BEGb[2] ,
    \Tile_X5Y7_S2BEGb[1] ,
    \Tile_X5Y7_S2BEGb[0] }),
    .S2MID({\Tile_X5Y7_S2BEG[7] ,
    \Tile_X5Y7_S2BEG[6] ,
    \Tile_X5Y7_S2BEG[5] ,
    \Tile_X5Y7_S2BEG[4] ,
    \Tile_X5Y7_S2BEG[3] ,
    \Tile_X5Y7_S2BEG[2] ,
    \Tile_X5Y7_S2BEG[1] ,
    \Tile_X5Y7_S2BEG[0] }),
    .S4BEG({\Tile_X5Y8_S4BEG[15] ,
    \Tile_X5Y8_S4BEG[14] ,
    \Tile_X5Y8_S4BEG[13] ,
    \Tile_X5Y8_S4BEG[12] ,
    \Tile_X5Y8_S4BEG[11] ,
    \Tile_X5Y8_S4BEG[10] ,
    \Tile_X5Y8_S4BEG[9] ,
    \Tile_X5Y8_S4BEG[8] ,
    \Tile_X5Y8_S4BEG[7] ,
    \Tile_X5Y8_S4BEG[6] ,
    \Tile_X5Y8_S4BEG[5] ,
    \Tile_X5Y8_S4BEG[4] ,
    \Tile_X5Y8_S4BEG[3] ,
    \Tile_X5Y8_S4BEG[2] ,
    \Tile_X5Y8_S4BEG[1] ,
    \Tile_X5Y8_S4BEG[0] }),
    .S4END({\Tile_X5Y7_S4BEG[15] ,
    \Tile_X5Y7_S4BEG[14] ,
    \Tile_X5Y7_S4BEG[13] ,
    \Tile_X5Y7_S4BEG[12] ,
    \Tile_X5Y7_S4BEG[11] ,
    \Tile_X5Y7_S4BEG[10] ,
    \Tile_X5Y7_S4BEG[9] ,
    \Tile_X5Y7_S4BEG[8] ,
    \Tile_X5Y7_S4BEG[7] ,
    \Tile_X5Y7_S4BEG[6] ,
    \Tile_X5Y7_S4BEG[5] ,
    \Tile_X5Y7_S4BEG[4] ,
    \Tile_X5Y7_S4BEG[3] ,
    \Tile_X5Y7_S4BEG[2] ,
    \Tile_X5Y7_S4BEG[1] ,
    \Tile_X5Y7_S4BEG[0] }),
    .W1BEG({\Tile_X5Y8_W1BEG[3] ,
    \Tile_X5Y8_W1BEG[2] ,
    \Tile_X5Y8_W1BEG[1] ,
    \Tile_X5Y8_W1BEG[0] }),
    .W2BEG({\Tile_X5Y8_W2BEG[7] ,
    \Tile_X5Y8_W2BEG[6] ,
    \Tile_X5Y8_W2BEG[5] ,
    \Tile_X5Y8_W2BEG[4] ,
    \Tile_X5Y8_W2BEG[3] ,
    \Tile_X5Y8_W2BEG[2] ,
    \Tile_X5Y8_W2BEG[1] ,
    \Tile_X5Y8_W2BEG[0] }),
    .W2BEGb({\Tile_X5Y8_W2BEGb[7] ,
    \Tile_X5Y8_W2BEGb[6] ,
    \Tile_X5Y8_W2BEGb[5] ,
    \Tile_X5Y8_W2BEGb[4] ,
    \Tile_X5Y8_W2BEGb[3] ,
    \Tile_X5Y8_W2BEGb[2] ,
    \Tile_X5Y8_W2BEGb[1] ,
    \Tile_X5Y8_W2BEGb[0] }),
    .W6BEG({\Tile_X5Y8_W6BEG[11] ,
    \Tile_X5Y8_W6BEG[10] ,
    \Tile_X5Y8_W6BEG[9] ,
    \Tile_X5Y8_W6BEG[8] ,
    \Tile_X5Y8_W6BEG[7] ,
    \Tile_X5Y8_W6BEG[6] ,
    \Tile_X5Y8_W6BEG[5] ,
    \Tile_X5Y8_W6BEG[4] ,
    \Tile_X5Y8_W6BEG[3] ,
    \Tile_X5Y8_W6BEG[2] ,
    \Tile_X5Y8_W6BEG[1] ,
    \Tile_X5Y8_W6BEG[0] }),
    .WW4BEG({\Tile_X5Y8_WW4BEG[15] ,
    \Tile_X5Y8_WW4BEG[14] ,
    \Tile_X5Y8_WW4BEG[13] ,
    \Tile_X5Y8_WW4BEG[12] ,
    \Tile_X5Y8_WW4BEG[11] ,
    \Tile_X5Y8_WW4BEG[10] ,
    \Tile_X5Y8_WW4BEG[9] ,
    \Tile_X5Y8_WW4BEG[8] ,
    \Tile_X5Y8_WW4BEG[7] ,
    \Tile_X5Y8_WW4BEG[6] ,
    \Tile_X5Y8_WW4BEG[5] ,
    \Tile_X5Y8_WW4BEG[4] ,
    \Tile_X5Y8_WW4BEG[3] ,
    \Tile_X5Y8_WW4BEG[2] ,
    \Tile_X5Y8_WW4BEG[1] ,
    \Tile_X5Y8_WW4BEG[0] }));
 SE_term Tile_X5Y9_SE_term (.UserCLK(UserCLK),
    .UserCLKo(Tile_X5Y9_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .FrameData({\Tile_X4Y9_FrameData_O[31] ,
    \Tile_X4Y9_FrameData_O[30] ,
    \Tile_X4Y9_FrameData_O[29] ,
    \Tile_X4Y9_FrameData_O[28] ,
    \Tile_X4Y9_FrameData_O[27] ,
    \Tile_X4Y9_FrameData_O[26] ,
    \Tile_X4Y9_FrameData_O[25] ,
    \Tile_X4Y9_FrameData_O[24] ,
    \Tile_X4Y9_FrameData_O[23] ,
    \Tile_X4Y9_FrameData_O[22] ,
    \Tile_X4Y9_FrameData_O[21] ,
    \Tile_X4Y9_FrameData_O[20] ,
    \Tile_X4Y9_FrameData_O[19] ,
    \Tile_X4Y9_FrameData_O[18] ,
    \Tile_X4Y9_FrameData_O[17] ,
    \Tile_X4Y9_FrameData_O[16] ,
    \Tile_X4Y9_FrameData_O[15] ,
    \Tile_X4Y9_FrameData_O[14] ,
    \Tile_X4Y9_FrameData_O[13] ,
    \Tile_X4Y9_FrameData_O[12] ,
    \Tile_X4Y9_FrameData_O[11] ,
    \Tile_X4Y9_FrameData_O[10] ,
    \Tile_X4Y9_FrameData_O[9] ,
    \Tile_X4Y9_FrameData_O[8] ,
    \Tile_X4Y9_FrameData_O[7] ,
    \Tile_X4Y9_FrameData_O[6] ,
    \Tile_X4Y9_FrameData_O[5] ,
    \Tile_X4Y9_FrameData_O[4] ,
    \Tile_X4Y9_FrameData_O[3] ,
    \Tile_X4Y9_FrameData_O[2] ,
    \Tile_X4Y9_FrameData_O[1] ,
    \Tile_X4Y9_FrameData_O[0] }),
    .FrameData_O({\Tile_X5Y9_FrameData_O[31] ,
    \Tile_X5Y9_FrameData_O[30] ,
    \Tile_X5Y9_FrameData_O[29] ,
    \Tile_X5Y9_FrameData_O[28] ,
    \Tile_X5Y9_FrameData_O[27] ,
    \Tile_X5Y9_FrameData_O[26] ,
    \Tile_X5Y9_FrameData_O[25] ,
    \Tile_X5Y9_FrameData_O[24] ,
    \Tile_X5Y9_FrameData_O[23] ,
    \Tile_X5Y9_FrameData_O[22] ,
    \Tile_X5Y9_FrameData_O[21] ,
    \Tile_X5Y9_FrameData_O[20] ,
    \Tile_X5Y9_FrameData_O[19] ,
    \Tile_X5Y9_FrameData_O[18] ,
    \Tile_X5Y9_FrameData_O[17] ,
    \Tile_X5Y9_FrameData_O[16] ,
    \Tile_X5Y9_FrameData_O[15] ,
    \Tile_X5Y9_FrameData_O[14] ,
    \Tile_X5Y9_FrameData_O[13] ,
    \Tile_X5Y9_FrameData_O[12] ,
    \Tile_X5Y9_FrameData_O[11] ,
    \Tile_X5Y9_FrameData_O[10] ,
    \Tile_X5Y9_FrameData_O[9] ,
    \Tile_X5Y9_FrameData_O[8] ,
    \Tile_X5Y9_FrameData_O[7] ,
    \Tile_X5Y9_FrameData_O[6] ,
    \Tile_X5Y9_FrameData_O[5] ,
    \Tile_X5Y9_FrameData_O[4] ,
    \Tile_X5Y9_FrameData_O[3] ,
    \Tile_X5Y9_FrameData_O[2] ,
    \Tile_X5Y9_FrameData_O[1] ,
    \Tile_X5Y9_FrameData_O[0] }),
    .FrameStrobe({FrameStrobe[119],
    FrameStrobe[118],
    FrameStrobe[117],
    FrameStrobe[116],
    FrameStrobe[115],
    FrameStrobe[114],
    FrameStrobe[113],
    FrameStrobe[112],
    FrameStrobe[111],
    FrameStrobe[110],
    FrameStrobe[109],
    FrameStrobe[108],
    FrameStrobe[107],
    FrameStrobe[106],
    FrameStrobe[105],
    FrameStrobe[104],
    FrameStrobe[103],
    FrameStrobe[102],
    FrameStrobe[101],
    FrameStrobe[100]}),
    .FrameStrobe_O({\Tile_X5Y9_FrameStrobe_O[19] ,
    \Tile_X5Y9_FrameStrobe_O[18] ,
    \Tile_X5Y9_FrameStrobe_O[17] ,
    \Tile_X5Y9_FrameStrobe_O[16] ,
    \Tile_X5Y9_FrameStrobe_O[15] ,
    \Tile_X5Y9_FrameStrobe_O[14] ,
    \Tile_X5Y9_FrameStrobe_O[13] ,
    \Tile_X5Y9_FrameStrobe_O[12] ,
    \Tile_X5Y9_FrameStrobe_O[11] ,
    \Tile_X5Y9_FrameStrobe_O[10] ,
    \Tile_X5Y9_FrameStrobe_O[9] ,
    \Tile_X5Y9_FrameStrobe_O[8] ,
    \Tile_X5Y9_FrameStrobe_O[7] ,
    \Tile_X5Y9_FrameStrobe_O[6] ,
    \Tile_X5Y9_FrameStrobe_O[5] ,
    \Tile_X5Y9_FrameStrobe_O[4] ,
    \Tile_X5Y9_FrameStrobe_O[3] ,
    \Tile_X5Y9_FrameStrobe_O[2] ,
    \Tile_X5Y9_FrameStrobe_O[1] ,
    \Tile_X5Y9_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X5Y9_N1BEG[3] ,
    \Tile_X5Y9_N1BEG[2] ,
    \Tile_X5Y9_N1BEG[1] ,
    \Tile_X5Y9_N1BEG[0] }),
    .N2BEG({\Tile_X5Y9_N2BEG[7] ,
    \Tile_X5Y9_N2BEG[6] ,
    \Tile_X5Y9_N2BEG[5] ,
    \Tile_X5Y9_N2BEG[4] ,
    \Tile_X5Y9_N2BEG[3] ,
    \Tile_X5Y9_N2BEG[2] ,
    \Tile_X5Y9_N2BEG[1] ,
    \Tile_X5Y9_N2BEG[0] }),
    .N2BEGb({\Tile_X5Y9_N2BEGb[7] ,
    \Tile_X5Y9_N2BEGb[6] ,
    \Tile_X5Y9_N2BEGb[5] ,
    \Tile_X5Y9_N2BEGb[4] ,
    \Tile_X5Y9_N2BEGb[3] ,
    \Tile_X5Y9_N2BEGb[2] ,
    \Tile_X5Y9_N2BEGb[1] ,
    \Tile_X5Y9_N2BEGb[0] }),
    .N4BEG({\Tile_X5Y9_N4BEG[15] ,
    \Tile_X5Y9_N4BEG[14] ,
    \Tile_X5Y9_N4BEG[13] ,
    \Tile_X5Y9_N4BEG[12] ,
    \Tile_X5Y9_N4BEG[11] ,
    \Tile_X5Y9_N4BEG[10] ,
    \Tile_X5Y9_N4BEG[9] ,
    \Tile_X5Y9_N4BEG[8] ,
    \Tile_X5Y9_N4BEG[7] ,
    \Tile_X5Y9_N4BEG[6] ,
    \Tile_X5Y9_N4BEG[5] ,
    \Tile_X5Y9_N4BEG[4] ,
    \Tile_X5Y9_N4BEG[3] ,
    \Tile_X5Y9_N4BEG[2] ,
    \Tile_X5Y9_N4BEG[1] ,
    \Tile_X5Y9_N4BEG[0] }),
    .S1END({\Tile_X5Y8_S1BEG[3] ,
    \Tile_X5Y8_S1BEG[2] ,
    \Tile_X5Y8_S1BEG[1] ,
    \Tile_X5Y8_S1BEG[0] }),
    .S2END({\Tile_X5Y8_S2BEGb[7] ,
    \Tile_X5Y8_S2BEGb[6] ,
    \Tile_X5Y8_S2BEGb[5] ,
    \Tile_X5Y8_S2BEGb[4] ,
    \Tile_X5Y8_S2BEGb[3] ,
    \Tile_X5Y8_S2BEGb[2] ,
    \Tile_X5Y8_S2BEGb[1] ,
    \Tile_X5Y8_S2BEGb[0] }),
    .S2MID({\Tile_X5Y8_S2BEG[7] ,
    \Tile_X5Y8_S2BEG[6] ,
    \Tile_X5Y8_S2BEG[5] ,
    \Tile_X5Y8_S2BEG[4] ,
    \Tile_X5Y8_S2BEG[3] ,
    \Tile_X5Y8_S2BEG[2] ,
    \Tile_X5Y8_S2BEG[1] ,
    \Tile_X5Y8_S2BEG[0] }),
    .S4END({\Tile_X5Y8_S4BEG[15] ,
    \Tile_X5Y8_S4BEG[14] ,
    \Tile_X5Y8_S4BEG[13] ,
    \Tile_X5Y8_S4BEG[12] ,
    \Tile_X5Y8_S4BEG[11] ,
    \Tile_X5Y8_S4BEG[10] ,
    \Tile_X5Y8_S4BEG[9] ,
    \Tile_X5Y8_S4BEG[8] ,
    \Tile_X5Y8_S4BEG[7] ,
    \Tile_X5Y8_S4BEG[6] ,
    \Tile_X5Y8_S4BEG[5] ,
    \Tile_X5Y8_S4BEG[4] ,
    \Tile_X5Y8_S4BEG[3] ,
    \Tile_X5Y8_S4BEG[2] ,
    \Tile_X5Y8_S4BEG[1] ,
    \Tile_X5Y8_S4BEG[0] }));
endmodule
