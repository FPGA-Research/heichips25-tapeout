module N_IO4 (A_I_top,
    A_O_top,
    A_T_top,
    B_I_top,
    B_O_top,
    B_T_top,
    C_I_top,
    C_O_top,
    C_T_top,
    Ci,
    D_I_top,
    D_O_top,
    D_T_top,
    UserCLK,
    UserCLKo,
    FrameData,
    FrameData_O,
    FrameStrobe,
    FrameStrobe_O,
    N1END,
    N2END,
    N2MID,
    N4END,
    NN4END,
    S1BEG,
    S2BEG,
    S2BEGb,
    S4BEG,
    SS4BEG);
 output A_I_top;
 input A_O_top;
 output A_T_top;
 output B_I_top;
 input B_O_top;
 output B_T_top;
 output C_I_top;
 input C_O_top;
 output C_T_top;
 input Ci;
 output D_I_top;
 input D_O_top;
 output D_T_top;
 input UserCLK;
 output UserCLKo;
 input [31:0] FrameData;
 output [31:0] FrameData_O;
 input [19:0] FrameStrobe;
 output [19:0] FrameStrobe_O;
 input [3:0] N1END;
 input [7:0] N2END;
 input [7:0] N2MID;
 input [15:0] N4END;
 input [15:0] NN4END;
 output [3:0] S1BEG;
 output [7:0] S2BEG;
 output [7:0] S2BEGb;
 output [15:0] S4BEG;
 output [15:0] SS4BEG;

 wire \Inst_A_IO_1_bidirectional_frame_config_pass.Q ;
 wire \Inst_B_IO_1_bidirectional_frame_config_pass.Q ;
 wire \Inst_C_IO_1_bidirectional_frame_config_pass.Q ;
 wire \Inst_D_IO_1_bidirectional_frame_config_pass.Q ;
 wire \Inst_N_IO4_ConfigMem.Inst_frame0_bit0.Q ;
 wire \Inst_N_IO4_ConfigMem.Inst_frame0_bit1.Q ;
 wire \Inst_N_IO4_ConfigMem.Inst_frame0_bit10.Q ;
 wire \Inst_N_IO4_ConfigMem.Inst_frame0_bit11.Q ;
 wire \Inst_N_IO4_ConfigMem.Inst_frame0_bit12.Q ;
 wire \Inst_N_IO4_ConfigMem.Inst_frame0_bit13.Q ;
 wire \Inst_N_IO4_ConfigMem.Inst_frame0_bit14.Q ;
 wire \Inst_N_IO4_ConfigMem.Inst_frame0_bit15.Q ;
 wire \Inst_N_IO4_ConfigMem.Inst_frame0_bit16.Q ;
 wire \Inst_N_IO4_ConfigMem.Inst_frame0_bit17.Q ;
 wire \Inst_N_IO4_ConfigMem.Inst_frame0_bit18.Q ;
 wire \Inst_N_IO4_ConfigMem.Inst_frame0_bit19.Q ;
 wire \Inst_N_IO4_ConfigMem.Inst_frame0_bit2.Q ;
 wire \Inst_N_IO4_ConfigMem.Inst_frame0_bit20.Q ;
 wire \Inst_N_IO4_ConfigMem.Inst_frame0_bit21.Q ;
 wire \Inst_N_IO4_ConfigMem.Inst_frame0_bit22.Q ;
 wire \Inst_N_IO4_ConfigMem.Inst_frame0_bit23.Q ;
 wire \Inst_N_IO4_ConfigMem.Inst_frame0_bit24.Q ;
 wire \Inst_N_IO4_ConfigMem.Inst_frame0_bit25.Q ;
 wire \Inst_N_IO4_ConfigMem.Inst_frame0_bit26.Q ;
 wire \Inst_N_IO4_ConfigMem.Inst_frame0_bit27.Q ;
 wire \Inst_N_IO4_ConfigMem.Inst_frame0_bit28.Q ;
 wire \Inst_N_IO4_ConfigMem.Inst_frame0_bit29.Q ;
 wire \Inst_N_IO4_ConfigMem.Inst_frame0_bit3.Q ;
 wire \Inst_N_IO4_ConfigMem.Inst_frame0_bit30.Q ;
 wire \Inst_N_IO4_ConfigMem.Inst_frame0_bit31.Q ;
 wire \Inst_N_IO4_ConfigMem.Inst_frame0_bit4.Q ;
 wire \Inst_N_IO4_ConfigMem.Inst_frame0_bit5.Q ;
 wire \Inst_N_IO4_ConfigMem.Inst_frame0_bit6.Q ;
 wire \Inst_N_IO4_ConfigMem.Inst_frame0_bit7.Q ;
 wire \Inst_N_IO4_ConfigMem.Inst_frame0_bit8.Q ;
 wire \Inst_N_IO4_ConfigMem.Inst_frame0_bit9.Q ;
 wire \Inst_N_IO4_ConfigMem.Inst_frame1_bit0.Q ;
 wire \Inst_N_IO4_ConfigMem.Inst_frame1_bit1.Q ;
 wire \Inst_N_IO4_ConfigMem.Inst_frame1_bit10.Q ;
 wire \Inst_N_IO4_ConfigMem.Inst_frame1_bit11.Q ;
 wire \Inst_N_IO4_ConfigMem.Inst_frame1_bit12.Q ;
 wire \Inst_N_IO4_ConfigMem.Inst_frame1_bit13.Q ;
 wire \Inst_N_IO4_ConfigMem.Inst_frame1_bit14.Q ;
 wire \Inst_N_IO4_ConfigMem.Inst_frame1_bit15.Q ;
 wire \Inst_N_IO4_ConfigMem.Inst_frame1_bit16.Q ;
 wire \Inst_N_IO4_ConfigMem.Inst_frame1_bit17.Q ;
 wire \Inst_N_IO4_ConfigMem.Inst_frame1_bit18.Q ;
 wire \Inst_N_IO4_ConfigMem.Inst_frame1_bit19.Q ;
 wire \Inst_N_IO4_ConfigMem.Inst_frame1_bit2.Q ;
 wire \Inst_N_IO4_ConfigMem.Inst_frame1_bit20.Q ;
 wire \Inst_N_IO4_ConfigMem.Inst_frame1_bit21.Q ;
 wire \Inst_N_IO4_ConfigMem.Inst_frame1_bit22.Q ;
 wire \Inst_N_IO4_ConfigMem.Inst_frame1_bit23.Q ;
 wire \Inst_N_IO4_ConfigMem.Inst_frame1_bit24.Q ;
 wire \Inst_N_IO4_ConfigMem.Inst_frame1_bit25.Q ;
 wire \Inst_N_IO4_ConfigMem.Inst_frame1_bit26.Q ;
 wire \Inst_N_IO4_ConfigMem.Inst_frame1_bit27.Q ;
 wire \Inst_N_IO4_ConfigMem.Inst_frame1_bit28.Q ;
 wire \Inst_N_IO4_ConfigMem.Inst_frame1_bit29.Q ;
 wire \Inst_N_IO4_ConfigMem.Inst_frame1_bit3.Q ;
 wire \Inst_N_IO4_ConfigMem.Inst_frame1_bit30.Q ;
 wire \Inst_N_IO4_ConfigMem.Inst_frame1_bit31.Q ;
 wire \Inst_N_IO4_ConfigMem.Inst_frame1_bit4.Q ;
 wire \Inst_N_IO4_ConfigMem.Inst_frame1_bit5.Q ;
 wire \Inst_N_IO4_ConfigMem.Inst_frame1_bit6.Q ;
 wire \Inst_N_IO4_ConfigMem.Inst_frame1_bit7.Q ;
 wire \Inst_N_IO4_ConfigMem.Inst_frame1_bit8.Q ;
 wire \Inst_N_IO4_ConfigMem.Inst_frame1_bit9.Q ;
 wire \Inst_N_IO4_ConfigMem.Inst_frame2_bit0.Q ;
 wire \Inst_N_IO4_ConfigMem.Inst_frame2_bit1.Q ;
 wire \Inst_N_IO4_ConfigMem.Inst_frame2_bit10.Q ;
 wire \Inst_N_IO4_ConfigMem.Inst_frame2_bit11.Q ;
 wire \Inst_N_IO4_ConfigMem.Inst_frame2_bit12.Q ;
 wire \Inst_N_IO4_ConfigMem.Inst_frame2_bit13.Q ;
 wire \Inst_N_IO4_ConfigMem.Inst_frame2_bit14.Q ;
 wire \Inst_N_IO4_ConfigMem.Inst_frame2_bit15.Q ;
 wire \Inst_N_IO4_ConfigMem.Inst_frame2_bit16.Q ;
 wire \Inst_N_IO4_ConfigMem.Inst_frame2_bit17.Q ;
 wire \Inst_N_IO4_ConfigMem.Inst_frame2_bit18.Q ;
 wire \Inst_N_IO4_ConfigMem.Inst_frame2_bit19.Q ;
 wire \Inst_N_IO4_ConfigMem.Inst_frame2_bit2.Q ;
 wire \Inst_N_IO4_ConfigMem.Inst_frame2_bit20.Q ;
 wire \Inst_N_IO4_ConfigMem.Inst_frame2_bit21.Q ;
 wire \Inst_N_IO4_ConfigMem.Inst_frame2_bit22.Q ;
 wire \Inst_N_IO4_ConfigMem.Inst_frame2_bit23.Q ;
 wire \Inst_N_IO4_ConfigMem.Inst_frame2_bit24.Q ;
 wire \Inst_N_IO4_ConfigMem.Inst_frame2_bit25.Q ;
 wire \Inst_N_IO4_ConfigMem.Inst_frame2_bit26.Q ;
 wire \Inst_N_IO4_ConfigMem.Inst_frame2_bit27.Q ;
 wire \Inst_N_IO4_ConfigMem.Inst_frame2_bit28.Q ;
 wire \Inst_N_IO4_ConfigMem.Inst_frame2_bit29.Q ;
 wire \Inst_N_IO4_ConfigMem.Inst_frame2_bit3.Q ;
 wire \Inst_N_IO4_ConfigMem.Inst_frame2_bit30.Q ;
 wire \Inst_N_IO4_ConfigMem.Inst_frame2_bit31.Q ;
 wire \Inst_N_IO4_ConfigMem.Inst_frame2_bit4.Q ;
 wire \Inst_N_IO4_ConfigMem.Inst_frame2_bit5.Q ;
 wire \Inst_N_IO4_ConfigMem.Inst_frame2_bit6.Q ;
 wire \Inst_N_IO4_ConfigMem.Inst_frame2_bit7.Q ;
 wire \Inst_N_IO4_ConfigMem.Inst_frame2_bit8.Q ;
 wire \Inst_N_IO4_ConfigMem.Inst_frame2_bit9.Q ;
 wire \Inst_N_IO4_ConfigMem.Inst_frame3_bit0.Q ;
 wire \Inst_N_IO4_ConfigMem.Inst_frame3_bit1.Q ;
 wire \Inst_N_IO4_ConfigMem.Inst_frame3_bit10.Q ;
 wire \Inst_N_IO4_ConfigMem.Inst_frame3_bit11.Q ;
 wire \Inst_N_IO4_ConfigMem.Inst_frame3_bit12.Q ;
 wire \Inst_N_IO4_ConfigMem.Inst_frame3_bit13.Q ;
 wire \Inst_N_IO4_ConfigMem.Inst_frame3_bit14.Q ;
 wire \Inst_N_IO4_ConfigMem.Inst_frame3_bit15.Q ;
 wire \Inst_N_IO4_ConfigMem.Inst_frame3_bit16.Q ;
 wire \Inst_N_IO4_ConfigMem.Inst_frame3_bit17.Q ;
 wire \Inst_N_IO4_ConfigMem.Inst_frame3_bit18.Q ;
 wire \Inst_N_IO4_ConfigMem.Inst_frame3_bit19.Q ;
 wire \Inst_N_IO4_ConfigMem.Inst_frame3_bit2.Q ;
 wire \Inst_N_IO4_ConfigMem.Inst_frame3_bit20.Q ;
 wire \Inst_N_IO4_ConfigMem.Inst_frame3_bit21.Q ;
 wire \Inst_N_IO4_ConfigMem.Inst_frame3_bit22.Q ;
 wire \Inst_N_IO4_ConfigMem.Inst_frame3_bit23.Q ;
 wire \Inst_N_IO4_ConfigMem.Inst_frame3_bit24.Q ;
 wire \Inst_N_IO4_ConfigMem.Inst_frame3_bit25.Q ;
 wire \Inst_N_IO4_ConfigMem.Inst_frame3_bit26.Q ;
 wire \Inst_N_IO4_ConfigMem.Inst_frame3_bit27.Q ;
 wire \Inst_N_IO4_ConfigMem.Inst_frame3_bit28.Q ;
 wire \Inst_N_IO4_ConfigMem.Inst_frame3_bit29.Q ;
 wire \Inst_N_IO4_ConfigMem.Inst_frame3_bit3.Q ;
 wire \Inst_N_IO4_ConfigMem.Inst_frame3_bit30.Q ;
 wire \Inst_N_IO4_ConfigMem.Inst_frame3_bit31.Q ;
 wire \Inst_N_IO4_ConfigMem.Inst_frame3_bit4.Q ;
 wire \Inst_N_IO4_ConfigMem.Inst_frame3_bit5.Q ;
 wire \Inst_N_IO4_ConfigMem.Inst_frame3_bit6.Q ;
 wire \Inst_N_IO4_ConfigMem.Inst_frame3_bit7.Q ;
 wire \Inst_N_IO4_ConfigMem.Inst_frame3_bit8.Q ;
 wire \Inst_N_IO4_ConfigMem.Inst_frame3_bit9.Q ;
 wire \Inst_N_IO4_ConfigMem.Inst_frame4_bit28.Q ;
 wire \Inst_N_IO4_ConfigMem.Inst_frame4_bit29.Q ;
 wire \Inst_N_IO4_ConfigMem.Inst_frame4_bit30.Q ;
 wire \Inst_N_IO4_ConfigMem.Inst_frame4_bit31.Q ;
 wire \Inst_N_IO4_switch_matrix.S1BEG0 ;
 wire \Inst_N_IO4_switch_matrix.S1BEG1 ;
 wire \Inst_N_IO4_switch_matrix.S1BEG2 ;
 wire \Inst_N_IO4_switch_matrix.S1BEG3 ;
 wire \Inst_N_IO4_switch_matrix.S2BEG0 ;
 wire \Inst_N_IO4_switch_matrix.S2BEG1 ;
 wire \Inst_N_IO4_switch_matrix.S2BEG2 ;
 wire \Inst_N_IO4_switch_matrix.S2BEG3 ;
 wire \Inst_N_IO4_switch_matrix.S2BEG4 ;
 wire \Inst_N_IO4_switch_matrix.S2BEG5 ;
 wire \Inst_N_IO4_switch_matrix.S2BEG6 ;
 wire \Inst_N_IO4_switch_matrix.S2BEG7 ;
 wire \Inst_N_IO4_switch_matrix.S2BEGb0 ;
 wire \Inst_N_IO4_switch_matrix.S2BEGb1 ;
 wire \Inst_N_IO4_switch_matrix.S2BEGb2 ;
 wire \Inst_N_IO4_switch_matrix.S2BEGb3 ;
 wire \Inst_N_IO4_switch_matrix.S2BEGb4 ;
 wire \Inst_N_IO4_switch_matrix.S2BEGb5 ;
 wire \Inst_N_IO4_switch_matrix.S2BEGb6 ;
 wire \Inst_N_IO4_switch_matrix.S2BEGb7 ;
 wire \Inst_N_IO4_switch_matrix.S4BEG0 ;
 wire \Inst_N_IO4_switch_matrix.S4BEG1 ;
 wire \Inst_N_IO4_switch_matrix.S4BEG10 ;
 wire \Inst_N_IO4_switch_matrix.S4BEG11 ;
 wire \Inst_N_IO4_switch_matrix.S4BEG12 ;
 wire \Inst_N_IO4_switch_matrix.S4BEG13 ;
 wire \Inst_N_IO4_switch_matrix.S4BEG14 ;
 wire \Inst_N_IO4_switch_matrix.S4BEG15 ;
 wire \Inst_N_IO4_switch_matrix.S4BEG2 ;
 wire \Inst_N_IO4_switch_matrix.S4BEG3 ;
 wire \Inst_N_IO4_switch_matrix.S4BEG4 ;
 wire \Inst_N_IO4_switch_matrix.S4BEG5 ;
 wire \Inst_N_IO4_switch_matrix.S4BEG6 ;
 wire \Inst_N_IO4_switch_matrix.S4BEG7 ;
 wire \Inst_N_IO4_switch_matrix.S4BEG8 ;
 wire \Inst_N_IO4_switch_matrix.S4BEG9 ;
 wire \Inst_N_IO4_switch_matrix.SS4BEG0 ;
 wire \Inst_N_IO4_switch_matrix.SS4BEG1 ;
 wire \Inst_N_IO4_switch_matrix.SS4BEG10 ;
 wire \Inst_N_IO4_switch_matrix.SS4BEG11 ;
 wire \Inst_N_IO4_switch_matrix.SS4BEG12 ;
 wire \Inst_N_IO4_switch_matrix.SS4BEG13 ;
 wire \Inst_N_IO4_switch_matrix.SS4BEG14 ;
 wire \Inst_N_IO4_switch_matrix.SS4BEG15 ;
 wire \Inst_N_IO4_switch_matrix.SS4BEG2 ;
 wire \Inst_N_IO4_switch_matrix.SS4BEG3 ;
 wire \Inst_N_IO4_switch_matrix.SS4BEG4 ;
 wire \Inst_N_IO4_switch_matrix.SS4BEG5 ;
 wire \Inst_N_IO4_switch_matrix.SS4BEG6 ;
 wire \Inst_N_IO4_switch_matrix.SS4BEG7 ;
 wire \Inst_N_IO4_switch_matrix.SS4BEG8 ;
 wire \Inst_N_IO4_switch_matrix.SS4BEG9 ;
 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire UserCLK_regs;
 wire clknet_0_UserCLK;
 wire clknet_1_0__leaf_UserCLK;
 wire clknet_0_UserCLK_regs;
 wire clknet_1_0__leaf_UserCLK_regs;
 wire clknet_1_1__leaf_UserCLK_regs;

 sg13g2_inv_1 _083_ (.Y(_000_),
    .A(N2END[1]));
 sg13g2_inv_1 _084_ (.Y(_001_),
    .A(\Inst_N_IO4_ConfigMem.Inst_frame0_bit20.Q ));
 sg13g2_inv_1 _085_ (.Y(_002_),
    .A(\Inst_N_IO4_ConfigMem.Inst_frame0_bit21.Q ));
 sg13g2_inv_1 _086_ (.Y(_003_),
    .A(\Inst_N_IO4_ConfigMem.Inst_frame0_bit12.Q ));
 sg13g2_mux4_1 _087_ (.S0(\Inst_N_IO4_ConfigMem.Inst_frame3_bit14.Q ),
    .A0(N2MID[2]),
    .A1(N4END[2]),
    .A2(NN4END[2]),
    .A3(NN4END[10]),
    .S1(\Inst_N_IO4_ConfigMem.Inst_frame3_bit15.Q ),
    .X(\Inst_N_IO4_switch_matrix.S2BEG5 ));
 sg13g2_mux4_1 _088_ (.S0(\Inst_N_IO4_ConfigMem.Inst_frame3_bit12.Q ),
    .A0(N2MID[3]),
    .A1(N4END[3]),
    .A2(NN4END[3]),
    .A3(NN4END[11]),
    .S1(\Inst_N_IO4_ConfigMem.Inst_frame3_bit13.Q ),
    .X(\Inst_N_IO4_switch_matrix.S2BEG4 ));
 sg13g2_mux4_1 _089_ (.S0(\Inst_N_IO4_ConfigMem.Inst_frame3_bit10.Q ),
    .A0(N2MID[4]),
    .A1(N4END[4]),
    .A2(NN4END[4]),
    .A3(NN4END[12]),
    .S1(\Inst_N_IO4_ConfigMem.Inst_frame3_bit11.Q ),
    .X(\Inst_N_IO4_switch_matrix.S2BEG3 ));
 sg13g2_mux4_1 _090_ (.S0(\Inst_N_IO4_ConfigMem.Inst_frame3_bit8.Q ),
    .A0(N2MID[5]),
    .A1(N4END[5]),
    .A2(NN4END[5]),
    .A3(NN4END[13]),
    .S1(\Inst_N_IO4_ConfigMem.Inst_frame3_bit9.Q ),
    .X(\Inst_N_IO4_switch_matrix.S2BEG2 ));
 sg13g2_mux4_1 _091_ (.S0(\Inst_N_IO4_ConfigMem.Inst_frame3_bit6.Q ),
    .A0(N2MID[6]),
    .A1(N4END[6]),
    .A2(NN4END[6]),
    .A3(NN4END[14]),
    .S1(\Inst_N_IO4_ConfigMem.Inst_frame3_bit7.Q ),
    .X(\Inst_N_IO4_switch_matrix.S2BEG1 ));
 sg13g2_mux4_1 _092_ (.S0(\Inst_N_IO4_ConfigMem.Inst_frame3_bit4.Q ),
    .A0(N2MID[7]),
    .A1(N4END[7]),
    .A2(NN4END[7]),
    .A3(NN4END[15]),
    .S1(\Inst_N_IO4_ConfigMem.Inst_frame3_bit5.Q ),
    .X(\Inst_N_IO4_switch_matrix.S2BEG0 ));
 sg13g2_mux4_1 _093_ (.S0(\Inst_N_IO4_ConfigMem.Inst_frame3_bit2.Q ),
    .A0(N1END[0]),
    .A1(N1END[3]),
    .A2(\Inst_B_IO_1_bidirectional_frame_config_pass.Q ),
    .A3(\Inst_D_IO_1_bidirectional_frame_config_pass.Q ),
    .S1(\Inst_N_IO4_ConfigMem.Inst_frame3_bit3.Q ),
    .X(\Inst_N_IO4_switch_matrix.S1BEG3 ));
 sg13g2_mux4_1 _094_ (.S0(\Inst_N_IO4_ConfigMem.Inst_frame3_bit0.Q ),
    .A0(N1END[0]),
    .A1(N1END[1]),
    .A2(B_O_top),
    .A3(D_O_top),
    .S1(\Inst_N_IO4_ConfigMem.Inst_frame3_bit1.Q ),
    .X(\Inst_N_IO4_switch_matrix.S1BEG2 ));
 sg13g2_mux4_1 _095_ (.S0(\Inst_N_IO4_ConfigMem.Inst_frame4_bit30.Q ),
    .A0(N1END[1]),
    .A1(N1END[2]),
    .A2(\Inst_A_IO_1_bidirectional_frame_config_pass.Q ),
    .A3(\Inst_C_IO_1_bidirectional_frame_config_pass.Q ),
    .S1(\Inst_N_IO4_ConfigMem.Inst_frame4_bit31.Q ),
    .X(\Inst_N_IO4_switch_matrix.S1BEG1 ));
 sg13g2_mux4_1 _096_ (.S0(\Inst_N_IO4_ConfigMem.Inst_frame4_bit29.Q ),
    .A0(N1END[2]),
    .A1(A_O_top),
    .A2(N1END[3]),
    .A3(C_O_top),
    .S1(\Inst_N_IO4_ConfigMem.Inst_frame4_bit28.Q ),
    .X(\Inst_N_IO4_switch_matrix.S1BEG0 ));
 sg13g2_mux4_1 _097_ (.S0(\Inst_N_IO4_ConfigMem.Inst_frame0_bit8.Q ),
    .A0(N2MID[7]),
    .A1(N2END[0]),
    .A2(N2END[1]),
    .A3(N2END[2]),
    .S1(\Inst_N_IO4_ConfigMem.Inst_frame0_bit9.Q ),
    .X(_004_));
 sg13g2_o21ai_1 _098_ (.B1(\Inst_N_IO4_ConfigMem.Inst_frame0_bit8.Q ),
    .Y(_005_),
    .A1(\Inst_N_IO4_ConfigMem.Inst_frame0_bit9.Q ),
    .A2(N2END[4]));
 sg13g2_nor2_1 _099_ (.A(\Inst_N_IO4_ConfigMem.Inst_frame0_bit8.Q ),
    .B(\Inst_N_IO4_ConfigMem.Inst_frame0_bit9.Q ),
    .Y(_006_));
 sg13g2_nand2_1 _100_ (.Y(_007_),
    .A(N2END[3]),
    .B(_006_));
 sg13g2_nand3_1 _101_ (.B(_005_),
    .C(_007_),
    .A(\Inst_N_IO4_ConfigMem.Inst_frame0_bit10.Q ),
    .Y(_008_));
 sg13g2_o21ai_1 _102_ (.B1(_008_),
    .Y(A_T_top),
    .A1(\Inst_N_IO4_ConfigMem.Inst_frame0_bit10.Q ),
    .A2(_004_));
 sg13g2_mux4_1 _103_ (.S0(\Inst_N_IO4_ConfigMem.Inst_frame0_bit15.Q ),
    .A0(N2MID[6]),
    .A1(N2MID[7]),
    .A2(N2END[0]),
    .A3(N2END[4]),
    .S1(\Inst_N_IO4_ConfigMem.Inst_frame0_bit16.Q ),
    .X(_009_));
 sg13g2_o21ai_1 _104_ (.B1(\Inst_N_IO4_ConfigMem.Inst_frame0_bit15.Q ),
    .Y(_010_),
    .A1(\Inst_N_IO4_ConfigMem.Inst_frame0_bit16.Q ),
    .A2(N2END[6]));
 sg13g2_nor2_1 _105_ (.A(\Inst_N_IO4_ConfigMem.Inst_frame0_bit15.Q ),
    .B(\Inst_N_IO4_ConfigMem.Inst_frame0_bit16.Q ),
    .Y(_011_));
 sg13g2_nand2_1 _106_ (.Y(_012_),
    .A(N2END[5]),
    .B(_011_));
 sg13g2_nand3_1 _107_ (.B(_010_),
    .C(_012_),
    .A(\Inst_N_IO4_ConfigMem.Inst_frame0_bit17.Q ),
    .Y(_013_));
 sg13g2_o21ai_1 _108_ (.B1(_013_),
    .Y(B_T_top),
    .A1(\Inst_N_IO4_ConfigMem.Inst_frame0_bit17.Q ),
    .A2(_009_));
 sg13g2_nand2b_1 _109_ (.Y(_014_),
    .B(N2END[5]),
    .A_N(\Inst_N_IO4_ConfigMem.Inst_frame0_bit23.Q ));
 sg13g2_mux4_1 _110_ (.S0(\Inst_N_IO4_ConfigMem.Inst_frame0_bit22.Q ),
    .A0(N2MID[6]),
    .A1(N2MID[7]),
    .A2(N2END[0]),
    .A3(N2END[4]),
    .S1(\Inst_N_IO4_ConfigMem.Inst_frame0_bit23.Q ),
    .X(_015_));
 sg13g2_o21ai_1 _111_ (.B1(\Inst_N_IO4_ConfigMem.Inst_frame0_bit22.Q ),
    .Y(_016_),
    .A1(N2END[6]),
    .A2(\Inst_N_IO4_ConfigMem.Inst_frame0_bit23.Q ));
 sg13g2_o21ai_1 _112_ (.B1(\Inst_N_IO4_ConfigMem.Inst_frame0_bit24.Q ),
    .Y(_017_),
    .A1(\Inst_N_IO4_ConfigMem.Inst_frame0_bit22.Q ),
    .A2(_014_));
 sg13g2_nand2b_1 _113_ (.Y(_018_),
    .B(_016_),
    .A_N(_017_));
 sg13g2_o21ai_1 _114_ (.B1(_018_),
    .Y(C_T_top),
    .A1(\Inst_N_IO4_ConfigMem.Inst_frame0_bit24.Q ),
    .A2(_015_));
 sg13g2_nand2b_1 _115_ (.Y(_019_),
    .B(N2END[5]),
    .A_N(\Inst_N_IO4_ConfigMem.Inst_frame0_bit30.Q ));
 sg13g2_mux4_1 _116_ (.S0(\Inst_N_IO4_ConfigMem.Inst_frame0_bit29.Q ),
    .A0(N2MID[6]),
    .A1(N2MID[7]),
    .A2(N2END[0]),
    .A3(N2END[4]),
    .S1(\Inst_N_IO4_ConfigMem.Inst_frame0_bit30.Q ),
    .X(_020_));
 sg13g2_o21ai_1 _117_ (.B1(\Inst_N_IO4_ConfigMem.Inst_frame0_bit29.Q ),
    .Y(_021_),
    .A1(N2END[6]),
    .A2(\Inst_N_IO4_ConfigMem.Inst_frame0_bit30.Q ));
 sg13g2_o21ai_1 _118_ (.B1(\Inst_N_IO4_ConfigMem.Inst_frame0_bit31.Q ),
    .Y(_022_),
    .A1(\Inst_N_IO4_ConfigMem.Inst_frame0_bit29.Q ),
    .A2(_019_));
 sg13g2_nand2b_1 _119_ (.Y(_023_),
    .B(_021_),
    .A_N(_022_));
 sg13g2_o21ai_1 _120_ (.B1(_023_),
    .Y(D_T_top),
    .A1(\Inst_N_IO4_ConfigMem.Inst_frame0_bit31.Q ),
    .A2(_020_));
 sg13g2_nand2_1 _121_ (.Y(_024_),
    .A(N2END[5]),
    .B(\Inst_N_IO4_ConfigMem.Inst_frame0_bit25.Q ));
 sg13g2_nand2b_1 _122_ (.Y(_025_),
    .B(N2END[4]),
    .A_N(\Inst_N_IO4_ConfigMem.Inst_frame0_bit25.Q ));
 sg13g2_a21oi_1 _123_ (.A1(_024_),
    .A2(_025_),
    .Y(_026_),
    .B1(\Inst_N_IO4_ConfigMem.Inst_frame0_bit26.Q ));
 sg13g2_nor2b_1 _124_ (.A(N2END[7]),
    .B_N(\Inst_N_IO4_ConfigMem.Inst_frame0_bit25.Q ),
    .Y(_027_));
 sg13g2_o21ai_1 _125_ (.B1(\Inst_N_IO4_ConfigMem.Inst_frame0_bit26.Q ),
    .Y(_028_),
    .A1(N2END[6]),
    .A2(\Inst_N_IO4_ConfigMem.Inst_frame0_bit25.Q ));
 sg13g2_o21ai_1 _126_ (.B1(\Inst_N_IO4_ConfigMem.Inst_frame0_bit27.Q ),
    .Y(_029_),
    .A1(_027_),
    .A2(_028_));
 sg13g2_mux2_1 _127_ (.A0(N2END[2]),
    .A1(N2END[3]),
    .S(\Inst_N_IO4_ConfigMem.Inst_frame0_bit25.Q ),
    .X(_030_));
 sg13g2_or2_1 _128_ (.X(_031_),
    .B(\Inst_N_IO4_ConfigMem.Inst_frame0_bit25.Q ),
    .A(N2END[0]));
 sg13g2_a21oi_1 _129_ (.A1(_000_),
    .A2(\Inst_N_IO4_ConfigMem.Inst_frame0_bit25.Q ),
    .Y(_032_),
    .B1(\Inst_N_IO4_ConfigMem.Inst_frame0_bit26.Q ));
 sg13g2_a221oi_1 _130_ (.B2(_032_),
    .C1(\Inst_N_IO4_ConfigMem.Inst_frame0_bit27.Q ),
    .B1(_031_),
    .A1(\Inst_N_IO4_ConfigMem.Inst_frame0_bit26.Q ),
    .Y(_033_),
    .A2(_030_));
 sg13g2_o21ai_1 _131_ (.B1(\Inst_N_IO4_ConfigMem.Inst_frame0_bit28.Q ),
    .Y(_034_),
    .A1(_026_),
    .A2(_029_));
 sg13g2_mux4_1 _132_ (.S0(\Inst_N_IO4_ConfigMem.Inst_frame0_bit25.Q ),
    .A0(N2MID[0]),
    .A1(N2MID[1]),
    .A2(N2MID[2]),
    .A3(N2MID[3]),
    .S1(\Inst_N_IO4_ConfigMem.Inst_frame0_bit26.Q ),
    .X(_035_));
 sg13g2_mux4_1 _133_ (.S0(\Inst_N_IO4_ConfigMem.Inst_frame0_bit25.Q ),
    .A0(N2MID[4]),
    .A1(N2MID[5]),
    .A2(N2MID[6]),
    .A3(N2MID[7]),
    .S1(\Inst_N_IO4_ConfigMem.Inst_frame0_bit26.Q ),
    .X(_036_));
 sg13g2_mux2_1 _134_ (.A0(_035_),
    .A1(_036_),
    .S(\Inst_N_IO4_ConfigMem.Inst_frame0_bit27.Q ),
    .X(_037_));
 sg13g2_nand2b_1 _135_ (.Y(_038_),
    .B(_037_),
    .A_N(\Inst_N_IO4_ConfigMem.Inst_frame0_bit28.Q ));
 sg13g2_o21ai_1 _136_ (.B1(_038_),
    .Y(D_I_top),
    .A1(_033_),
    .A2(_034_));
 sg13g2_mux2_1 _137_ (.A0(N2END[2]),
    .A1(N2END[3]),
    .S(\Inst_N_IO4_ConfigMem.Inst_frame0_bit18.Q ),
    .X(_039_));
 sg13g2_mux2_1 _138_ (.A0(N2END[0]),
    .A1(N2END[1]),
    .S(\Inst_N_IO4_ConfigMem.Inst_frame0_bit18.Q ),
    .X(_040_));
 sg13g2_nand2b_1 _139_ (.Y(_041_),
    .B(_040_),
    .A_N(\Inst_N_IO4_ConfigMem.Inst_frame0_bit19.Q ));
 sg13g2_a21oi_1 _140_ (.A1(\Inst_N_IO4_ConfigMem.Inst_frame0_bit19.Q ),
    .A2(_039_),
    .Y(_042_),
    .B1(\Inst_N_IO4_ConfigMem.Inst_frame0_bit20.Q ));
 sg13g2_mux2_1 _141_ (.A0(N2END[4]),
    .A1(N2END[5]),
    .S(\Inst_N_IO4_ConfigMem.Inst_frame0_bit18.Q ),
    .X(_043_));
 sg13g2_nand2b_1 _142_ (.Y(_044_),
    .B(_043_),
    .A_N(\Inst_N_IO4_ConfigMem.Inst_frame0_bit19.Q ));
 sg13g2_mux2_1 _143_ (.A0(N2END[6]),
    .A1(N2END[7]),
    .S(\Inst_N_IO4_ConfigMem.Inst_frame0_bit18.Q ),
    .X(_045_));
 sg13g2_a21oi_1 _144_ (.A1(\Inst_N_IO4_ConfigMem.Inst_frame0_bit19.Q ),
    .A2(_045_),
    .Y(_046_),
    .B1(_001_));
 sg13g2_a221oi_1 _145_ (.B2(_046_),
    .C1(_002_),
    .B1(_044_),
    .A1(_041_),
    .Y(_047_),
    .A2(_042_));
 sg13g2_mux2_1 _146_ (.A0(N2MID[2]),
    .A1(N2MID[3]),
    .S(\Inst_N_IO4_ConfigMem.Inst_frame0_bit18.Q ),
    .X(_048_));
 sg13g2_mux2_1 _147_ (.A0(N2MID[0]),
    .A1(N2MID[1]),
    .S(\Inst_N_IO4_ConfigMem.Inst_frame0_bit18.Q ),
    .X(_049_));
 sg13g2_mux2_1 _148_ (.A0(N2MID[6]),
    .A1(N2MID[7]),
    .S(\Inst_N_IO4_ConfigMem.Inst_frame0_bit18.Q ),
    .X(_050_));
 sg13g2_mux2_1 _149_ (.A0(N2MID[4]),
    .A1(N2MID[5]),
    .S(\Inst_N_IO4_ConfigMem.Inst_frame0_bit18.Q ),
    .X(_051_));
 sg13g2_mux4_1 _150_ (.S0(\Inst_N_IO4_ConfigMem.Inst_frame0_bit20.Q ),
    .A0(_049_),
    .A1(_051_),
    .A2(_048_),
    .A3(_050_),
    .S1(\Inst_N_IO4_ConfigMem.Inst_frame0_bit19.Q ),
    .X(_052_));
 sg13g2_a21o_1 _151_ (.A2(_052_),
    .A1(_002_),
    .B1(_047_),
    .X(C_I_top));
 sg13g2_mux4_1 _152_ (.S0(\Inst_N_IO4_ConfigMem.Inst_frame0_bit12.Q ),
    .A0(N2END[0]),
    .A1(N2END[2]),
    .A2(N2END[1]),
    .A3(N2END[3]),
    .S1(\Inst_N_IO4_ConfigMem.Inst_frame0_bit11.Q ),
    .X(_053_));
 sg13g2_mux2_1 _153_ (.A0(N2END[4]),
    .A1(N2END[5]),
    .S(\Inst_N_IO4_ConfigMem.Inst_frame0_bit11.Q ),
    .X(_054_));
 sg13g2_nor2b_1 _154_ (.A(N2END[7]),
    .B_N(\Inst_N_IO4_ConfigMem.Inst_frame0_bit11.Q ),
    .Y(_055_));
 sg13g2_o21ai_1 _155_ (.B1(\Inst_N_IO4_ConfigMem.Inst_frame0_bit12.Q ),
    .Y(_056_),
    .A1(N2END[6]),
    .A2(\Inst_N_IO4_ConfigMem.Inst_frame0_bit11.Q ));
 sg13g2_o21ai_1 _156_ (.B1(\Inst_N_IO4_ConfigMem.Inst_frame0_bit13.Q ),
    .Y(_057_),
    .A1(_055_),
    .A2(_056_));
 sg13g2_a21oi_1 _157_ (.A1(_003_),
    .A2(_054_),
    .Y(_058_),
    .B1(_057_));
 sg13g2_o21ai_1 _158_ (.B1(\Inst_N_IO4_ConfigMem.Inst_frame0_bit14.Q ),
    .Y(_059_),
    .A1(\Inst_N_IO4_ConfigMem.Inst_frame0_bit13.Q ),
    .A2(_053_));
 sg13g2_mux4_1 _159_ (.S0(\Inst_N_IO4_ConfigMem.Inst_frame0_bit11.Q ),
    .A0(N2MID[0]),
    .A1(N2MID[1]),
    .A2(N2MID[2]),
    .A3(N2MID[3]),
    .S1(\Inst_N_IO4_ConfigMem.Inst_frame0_bit12.Q ),
    .X(_060_));
 sg13g2_mux4_1 _160_ (.S0(\Inst_N_IO4_ConfigMem.Inst_frame0_bit11.Q ),
    .A0(N2MID[4]),
    .A1(N2MID[5]),
    .A2(N2MID[6]),
    .A3(N2MID[7]),
    .S1(\Inst_N_IO4_ConfigMem.Inst_frame0_bit12.Q ),
    .X(_061_));
 sg13g2_mux2_1 _161_ (.A0(_060_),
    .A1(_061_),
    .S(\Inst_N_IO4_ConfigMem.Inst_frame0_bit13.Q ),
    .X(_062_));
 sg13g2_nand2b_1 _162_ (.Y(_063_),
    .B(_062_),
    .A_N(\Inst_N_IO4_ConfigMem.Inst_frame0_bit14.Q ));
 sg13g2_o21ai_1 _163_ (.B1(_063_),
    .Y(B_I_top),
    .A1(_058_),
    .A2(_059_));
 sg13g2_mux2_1 _164_ (.A0(N2END[2]),
    .A1(N2END[3]),
    .S(\Inst_N_IO4_ConfigMem.Inst_frame0_bit4.Q ),
    .X(_064_));
 sg13g2_or2_1 _165_ (.X(_065_),
    .B(\Inst_N_IO4_ConfigMem.Inst_frame0_bit4.Q ),
    .A(N2END[0]));
 sg13g2_a21oi_1 _166_ (.A1(_000_),
    .A2(\Inst_N_IO4_ConfigMem.Inst_frame0_bit4.Q ),
    .Y(_066_),
    .B1(\Inst_N_IO4_ConfigMem.Inst_frame0_bit5.Q ));
 sg13g2_a221oi_1 _167_ (.B2(_066_),
    .C1(\Inst_N_IO4_ConfigMem.Inst_frame0_bit6.Q ),
    .B1(_065_),
    .A1(\Inst_N_IO4_ConfigMem.Inst_frame0_bit5.Q ),
    .Y(_067_),
    .A2(_064_));
 sg13g2_nor2b_1 _168_ (.A(N2END[7]),
    .B_N(\Inst_N_IO4_ConfigMem.Inst_frame0_bit4.Q ),
    .Y(_068_));
 sg13g2_o21ai_1 _169_ (.B1(\Inst_N_IO4_ConfigMem.Inst_frame0_bit5.Q ),
    .Y(_069_),
    .A1(N2END[6]),
    .A2(\Inst_N_IO4_ConfigMem.Inst_frame0_bit4.Q ));
 sg13g2_nand2_1 _170_ (.Y(_070_),
    .A(N2END[5]),
    .B(\Inst_N_IO4_ConfigMem.Inst_frame0_bit4.Q ));
 sg13g2_nand2b_1 _171_ (.Y(_071_),
    .B(N2END[4]),
    .A_N(\Inst_N_IO4_ConfigMem.Inst_frame0_bit4.Q ));
 sg13g2_a21oi_1 _172_ (.A1(_070_),
    .A2(_071_),
    .Y(_072_),
    .B1(\Inst_N_IO4_ConfigMem.Inst_frame0_bit5.Q ));
 sg13g2_o21ai_1 _173_ (.B1(\Inst_N_IO4_ConfigMem.Inst_frame0_bit6.Q ),
    .Y(_073_),
    .A1(_068_),
    .A2(_069_));
 sg13g2_o21ai_1 _174_ (.B1(\Inst_N_IO4_ConfigMem.Inst_frame0_bit7.Q ),
    .Y(_074_),
    .A1(_072_),
    .A2(_073_));
 sg13g2_mux4_1 _175_ (.S0(\Inst_N_IO4_ConfigMem.Inst_frame0_bit4.Q ),
    .A0(N2MID[0]),
    .A1(N2MID[1]),
    .A2(N2MID[2]),
    .A3(N2MID[3]),
    .S1(\Inst_N_IO4_ConfigMem.Inst_frame0_bit5.Q ),
    .X(_075_));
 sg13g2_mux4_1 _176_ (.S0(\Inst_N_IO4_ConfigMem.Inst_frame0_bit4.Q ),
    .A0(N2MID[4]),
    .A1(N2MID[5]),
    .A2(N2MID[6]),
    .A3(N2MID[7]),
    .S1(\Inst_N_IO4_ConfigMem.Inst_frame0_bit5.Q ),
    .X(_076_));
 sg13g2_mux2_1 _177_ (.A0(_075_),
    .A1(_076_),
    .S(\Inst_N_IO4_ConfigMem.Inst_frame0_bit6.Q ),
    .X(_077_));
 sg13g2_nand2b_1 _178_ (.Y(_078_),
    .B(_077_),
    .A_N(\Inst_N_IO4_ConfigMem.Inst_frame0_bit7.Q ));
 sg13g2_o21ai_1 _179_ (.B1(_078_),
    .Y(A_I_top),
    .A1(_067_),
    .A2(_074_));
 sg13g2_mux4_1 _180_ (.S0(\Inst_N_IO4_ConfigMem.Inst_frame0_bit3.Q ),
    .A0(N2MID[1]),
    .A1(N2MID[5]),
    .A2(N2MID[3]),
    .A3(D_O_top),
    .S1(\Inst_N_IO4_ConfigMem.Inst_frame0_bit2.Q ),
    .X(\Inst_N_IO4_switch_matrix.SS4BEG15 ));
 sg13g2_mux4_1 _181_ (.S0(\Inst_N_IO4_ConfigMem.Inst_frame0_bit0.Q ),
    .A0(N2MID[0]),
    .A1(N2MID[2]),
    .A2(N2MID[4]),
    .A3(C_O_top),
    .S1(\Inst_N_IO4_ConfigMem.Inst_frame0_bit1.Q ),
    .X(\Inst_N_IO4_switch_matrix.SS4BEG14 ));
 sg13g2_mux4_1 _182_ (.S0(\Inst_N_IO4_ConfigMem.Inst_frame1_bit30.Q ),
    .A0(N4END[7]),
    .A1(N4END[9]),
    .A2(N4END[11]),
    .A3(\Inst_B_IO_1_bidirectional_frame_config_pass.Q ),
    .S1(\Inst_N_IO4_ConfigMem.Inst_frame1_bit31.Q ),
    .X(\Inst_N_IO4_switch_matrix.SS4BEG13 ));
 sg13g2_mux4_1 _183_ (.S0(\Inst_N_IO4_ConfigMem.Inst_frame1_bit29.Q ),
    .A0(N4END[1]),
    .A1(N4END[5]),
    .A2(N4END[3]),
    .A3(\Inst_A_IO_1_bidirectional_frame_config_pass.Q ),
    .S1(\Inst_N_IO4_ConfigMem.Inst_frame1_bit28.Q ),
    .X(\Inst_N_IO4_switch_matrix.SS4BEG12 ));
 sg13g2_mux4_1 _184_ (.S0(\Inst_N_IO4_ConfigMem.Inst_frame1_bit26.Q ),
    .A0(N4END[6]),
    .A1(N4END[8]),
    .A2(N4END[10]),
    .A3(B_O_top),
    .S1(\Inst_N_IO4_ConfigMem.Inst_frame1_bit27.Q ),
    .X(\Inst_N_IO4_switch_matrix.SS4BEG11 ));
 sg13g2_mux4_1 _185_ (.S0(\Inst_N_IO4_ConfigMem.Inst_frame1_bit24.Q ),
    .A0(N4END[0]),
    .A1(N4END[2]),
    .A2(N4END[4]),
    .A3(A_O_top),
    .S1(\Inst_N_IO4_ConfigMem.Inst_frame1_bit25.Q ),
    .X(\Inst_N_IO4_switch_matrix.SS4BEG10 ));
 sg13g2_mux4_1 _186_ (.S0(\Inst_N_IO4_ConfigMem.Inst_frame1_bit22.Q ),
    .A0(N4END[3]),
    .A1(N4END[5]),
    .A2(N4END[7]),
    .A3(\Inst_D_IO_1_bidirectional_frame_config_pass.Q ),
    .S1(\Inst_N_IO4_ConfigMem.Inst_frame1_bit23.Q ),
    .X(\Inst_N_IO4_switch_matrix.SS4BEG9 ));
 sg13g2_mux4_1 _187_ (.S0(\Inst_N_IO4_ConfigMem.Inst_frame1_bit20.Q ),
    .A0(N4END[6]),
    .A1(N4END[8]),
    .A2(N4END[10]),
    .A3(\Inst_C_IO_1_bidirectional_frame_config_pass.Q ),
    .S1(\Inst_N_IO4_ConfigMem.Inst_frame1_bit21.Q ),
    .X(\Inst_N_IO4_switch_matrix.SS4BEG8 ));
 sg13g2_mux4_1 _188_ (.S0(\Inst_N_IO4_ConfigMem.Inst_frame1_bit18.Q ),
    .A0(N2MID[3]),
    .A1(N2MID[5]),
    .A2(N2MID[7]),
    .A3(D_O_top),
    .S1(\Inst_N_IO4_ConfigMem.Inst_frame1_bit19.Q ),
    .X(\Inst_N_IO4_switch_matrix.SS4BEG7 ));
 sg13g2_mux4_1 _189_ (.S0(\Inst_N_IO4_ConfigMem.Inst_frame1_bit17.Q ),
    .A0(N2MID[2]),
    .A1(N2MID[6]),
    .A2(N2MID[4]),
    .A3(C_O_top),
    .S1(\Inst_N_IO4_ConfigMem.Inst_frame1_bit16.Q ),
    .X(\Inst_N_IO4_switch_matrix.SS4BEG6 ));
 sg13g2_mux4_1 _190_ (.S0(\Inst_N_IO4_ConfigMem.Inst_frame1_bit14.Q ),
    .A0(N2END[1]),
    .A1(N2END[3]),
    .A2(N2END[5]),
    .A3(\Inst_D_IO_1_bidirectional_frame_config_pass.Q ),
    .S1(\Inst_N_IO4_ConfigMem.Inst_frame1_bit15.Q ),
    .X(\Inst_N_IO4_switch_matrix.SS4BEG5 ));
 sg13g2_mux4_1 _191_ (.S0(\Inst_N_IO4_ConfigMem.Inst_frame1_bit12.Q ),
    .A0(N2END[0]),
    .A1(N2END[2]),
    .A2(N2END[4]),
    .A3(\Inst_C_IO_1_bidirectional_frame_config_pass.Q ),
    .S1(\Inst_N_IO4_ConfigMem.Inst_frame1_bit13.Q ),
    .X(\Inst_N_IO4_switch_matrix.SS4BEG4 ));
 sg13g2_mux4_1 _192_ (.S0(\Inst_N_IO4_ConfigMem.Inst_frame1_bit10.Q ),
    .A0(N4END[7]),
    .A1(N4END[9]),
    .A2(N4END[11]),
    .A3(\Inst_B_IO_1_bidirectional_frame_config_pass.Q ),
    .S1(\Inst_N_IO4_ConfigMem.Inst_frame1_bit11.Q ),
    .X(\Inst_N_IO4_switch_matrix.SS4BEG3 ));
 sg13g2_mux4_1 _193_ (.S0(\Inst_N_IO4_ConfigMem.Inst_frame1_bit8.Q ),
    .A0(N2END[6]),
    .A1(N2END[7]),
    .A2(N4END[1]),
    .A3(\Inst_A_IO_1_bidirectional_frame_config_pass.Q ),
    .S1(\Inst_N_IO4_ConfigMem.Inst_frame1_bit9.Q ),
    .X(\Inst_N_IO4_switch_matrix.SS4BEG2 ));
 sg13g2_mux4_1 _194_ (.S0(\Inst_N_IO4_ConfigMem.Inst_frame1_bit6.Q ),
    .A0(N4END[6]),
    .A1(N4END[8]),
    .A2(N4END[10]),
    .A3(B_O_top),
    .S1(\Inst_N_IO4_ConfigMem.Inst_frame1_bit7.Q ),
    .X(\Inst_N_IO4_switch_matrix.SS4BEG1 ));
 sg13g2_mux4_1 _195_ (.S0(\Inst_N_IO4_ConfigMem.Inst_frame1_bit4.Q ),
    .A0(N4END[0]),
    .A1(N4END[2]),
    .A2(N4END[4]),
    .A3(A_O_top),
    .S1(\Inst_N_IO4_ConfigMem.Inst_frame1_bit5.Q ),
    .X(\Inst_N_IO4_switch_matrix.SS4BEG0 ));
 sg13g2_mux4_1 _196_ (.S0(\Inst_N_IO4_ConfigMem.Inst_frame1_bit2.Q ),
    .A0(N4END[0]),
    .A1(NN4END[0]),
    .A2(\Inst_B_IO_1_bidirectional_frame_config_pass.Q ),
    .A3(\Inst_D_IO_1_bidirectional_frame_config_pass.Q ),
    .S1(\Inst_N_IO4_ConfigMem.Inst_frame1_bit3.Q ),
    .X(\Inst_N_IO4_switch_matrix.S4BEG15 ));
 sg13g2_mux4_1 _197_ (.S0(\Inst_N_IO4_ConfigMem.Inst_frame1_bit0.Q ),
    .A0(N4END[1]),
    .A1(NN4END[1]),
    .A2(\Inst_A_IO_1_bidirectional_frame_config_pass.Q ),
    .A3(\Inst_C_IO_1_bidirectional_frame_config_pass.Q ),
    .S1(\Inst_N_IO4_ConfigMem.Inst_frame1_bit1.Q ),
    .X(\Inst_N_IO4_switch_matrix.S4BEG14 ));
 sg13g2_mux4_1 _198_ (.S0(\Inst_N_IO4_ConfigMem.Inst_frame2_bit30.Q ),
    .A0(N4END[4]),
    .A1(NN4END[4]),
    .A2(\Inst_B_IO_1_bidirectional_frame_config_pass.Q ),
    .A3(\Inst_D_IO_1_bidirectional_frame_config_pass.Q ),
    .S1(\Inst_N_IO4_ConfigMem.Inst_frame2_bit31.Q ),
    .X(\Inst_N_IO4_switch_matrix.S4BEG13 ));
 sg13g2_mux4_1 _199_ (.S0(\Inst_N_IO4_ConfigMem.Inst_frame2_bit28.Q ),
    .A0(N4END[5]),
    .A1(NN4END[5]),
    .A2(\Inst_A_IO_1_bidirectional_frame_config_pass.Q ),
    .A3(\Inst_C_IO_1_bidirectional_frame_config_pass.Q ),
    .S1(\Inst_N_IO4_ConfigMem.Inst_frame2_bit29.Q ),
    .X(\Inst_N_IO4_switch_matrix.S4BEG12 ));
 sg13g2_mux4_1 _200_ (.S0(\Inst_N_IO4_ConfigMem.Inst_frame2_bit26.Q ),
    .A0(N4END[8]),
    .A1(NN4END[8]),
    .A2(\Inst_B_IO_1_bidirectional_frame_config_pass.Q ),
    .A3(\Inst_D_IO_1_bidirectional_frame_config_pass.Q ),
    .S1(\Inst_N_IO4_ConfigMem.Inst_frame2_bit27.Q ),
    .X(\Inst_N_IO4_switch_matrix.S4BEG11 ));
 sg13g2_mux4_1 _201_ (.S0(\Inst_N_IO4_ConfigMem.Inst_frame2_bit24.Q ),
    .A0(N4END[9]),
    .A1(NN4END[9]),
    .A2(\Inst_A_IO_1_bidirectional_frame_config_pass.Q ),
    .A3(\Inst_C_IO_1_bidirectional_frame_config_pass.Q ),
    .S1(\Inst_N_IO4_ConfigMem.Inst_frame2_bit25.Q ),
    .X(\Inst_N_IO4_switch_matrix.S4BEG10 ));
 sg13g2_mux4_1 _202_ (.S0(\Inst_N_IO4_ConfigMem.Inst_frame2_bit23.Q ),
    .A0(N4END[12]),
    .A1(\Inst_B_IO_1_bidirectional_frame_config_pass.Q ),
    .A2(NN4END[12]),
    .A3(\Inst_D_IO_1_bidirectional_frame_config_pass.Q ),
    .S1(\Inst_N_IO4_ConfigMem.Inst_frame2_bit22.Q ),
    .X(\Inst_N_IO4_switch_matrix.S4BEG9 ));
 sg13g2_mux4_1 _203_ (.S0(\Inst_N_IO4_ConfigMem.Inst_frame2_bit21.Q ),
    .A0(N4END[13]),
    .A1(\Inst_A_IO_1_bidirectional_frame_config_pass.Q ),
    .A2(NN4END[13]),
    .A3(\Inst_C_IO_1_bidirectional_frame_config_pass.Q ),
    .S1(\Inst_N_IO4_ConfigMem.Inst_frame2_bit20.Q ),
    .X(\Inst_N_IO4_switch_matrix.S4BEG8 ));
 sg13g2_mux4_1 _204_ (.S0(\Inst_N_IO4_ConfigMem.Inst_frame2_bit19.Q ),
    .A0(N4END[2]),
    .A1(B_O_top),
    .A2(NN4END[2]),
    .A3(D_O_top),
    .S1(\Inst_N_IO4_ConfigMem.Inst_frame2_bit18.Q ),
    .X(\Inst_N_IO4_switch_matrix.S4BEG7 ));
 sg13g2_mux4_1 _205_ (.S0(\Inst_N_IO4_ConfigMem.Inst_frame2_bit16.Q ),
    .A0(N4END[3]),
    .A1(NN4END[3]),
    .A2(A_O_top),
    .A3(C_O_top),
    .S1(\Inst_N_IO4_ConfigMem.Inst_frame2_bit17.Q ),
    .X(\Inst_N_IO4_switch_matrix.S4BEG6 ));
 sg13g2_mux4_1 _206_ (.S0(\Inst_N_IO4_ConfigMem.Inst_frame2_bit14.Q ),
    .A0(N4END[6]),
    .A1(NN4END[6]),
    .A2(B_O_top),
    .A3(D_O_top),
    .S1(\Inst_N_IO4_ConfigMem.Inst_frame2_bit15.Q ),
    .X(\Inst_N_IO4_switch_matrix.S4BEG5 ));
 sg13g2_mux4_1 _207_ (.S0(\Inst_N_IO4_ConfigMem.Inst_frame2_bit12.Q ),
    .A0(N4END[7]),
    .A1(NN4END[7]),
    .A2(A_O_top),
    .A3(C_O_top),
    .S1(\Inst_N_IO4_ConfigMem.Inst_frame2_bit13.Q ),
    .X(\Inst_N_IO4_switch_matrix.S4BEG4 ));
 sg13g2_mux4_1 _208_ (.S0(\Inst_N_IO4_ConfigMem.Inst_frame2_bit11.Q ),
    .A0(N4END[10]),
    .A1(B_O_top),
    .A2(NN4END[10]),
    .A3(D_O_top),
    .S1(\Inst_N_IO4_ConfigMem.Inst_frame2_bit10.Q ),
    .X(\Inst_N_IO4_switch_matrix.S4BEG3 ));
 sg13g2_mux4_1 _209_ (.S0(\Inst_N_IO4_ConfigMem.Inst_frame2_bit9.Q ),
    .A0(N4END[11]),
    .A1(A_O_top),
    .A2(NN4END[11]),
    .A3(C_O_top),
    .S1(\Inst_N_IO4_ConfigMem.Inst_frame2_bit8.Q ),
    .X(\Inst_N_IO4_switch_matrix.S4BEG2 ));
 sg13g2_mux4_1 _210_ (.S0(\Inst_N_IO4_ConfigMem.Inst_frame2_bit7.Q ),
    .A0(N4END[14]),
    .A1(B_O_top),
    .A2(NN4END[14]),
    .A3(D_O_top),
    .S1(\Inst_N_IO4_ConfigMem.Inst_frame2_bit6.Q ),
    .X(\Inst_N_IO4_switch_matrix.S4BEG1 ));
 sg13g2_mux4_1 _211_ (.S0(\Inst_N_IO4_ConfigMem.Inst_frame2_bit5.Q ),
    .A0(N4END[15]),
    .A1(A_O_top),
    .A2(NN4END[15]),
    .A3(C_O_top),
    .S1(\Inst_N_IO4_ConfigMem.Inst_frame2_bit4.Q ),
    .X(\Inst_N_IO4_switch_matrix.S4BEG0 ));
 sg13g2_mux4_1 _212_ (.S0(\Inst_N_IO4_ConfigMem.Inst_frame2_bit2.Q ),
    .A0(N2END[0]),
    .A1(N4END[0]),
    .A2(NN4END[0]),
    .A3(NN4END[8]),
    .S1(\Inst_N_IO4_ConfigMem.Inst_frame2_bit3.Q ),
    .X(\Inst_N_IO4_switch_matrix.S2BEGb7 ));
 sg13g2_mux4_1 _213_ (.S0(\Inst_N_IO4_ConfigMem.Inst_frame2_bit0.Q ),
    .A0(N2END[1]),
    .A1(N4END[1]),
    .A2(NN4END[1]),
    .A3(NN4END[9]),
    .S1(\Inst_N_IO4_ConfigMem.Inst_frame2_bit1.Q ),
    .X(\Inst_N_IO4_switch_matrix.S2BEGb6 ));
 sg13g2_mux4_1 _214_ (.S0(\Inst_N_IO4_ConfigMem.Inst_frame3_bit30.Q ),
    .A0(N2END[2]),
    .A1(N4END[2]),
    .A2(NN4END[2]),
    .A3(NN4END[10]),
    .S1(\Inst_N_IO4_ConfigMem.Inst_frame3_bit31.Q ),
    .X(\Inst_N_IO4_switch_matrix.S2BEGb5 ));
 sg13g2_mux4_1 _215_ (.S0(\Inst_N_IO4_ConfigMem.Inst_frame3_bit29.Q ),
    .A0(N2END[3]),
    .A1(NN4END[3]),
    .A2(N4END[3]),
    .A3(NN4END[11]),
    .S1(\Inst_N_IO4_ConfigMem.Inst_frame3_bit28.Q ),
    .X(\Inst_N_IO4_switch_matrix.S2BEGb4 ));
 sg13g2_mux4_1 _216_ (.S0(\Inst_N_IO4_ConfigMem.Inst_frame3_bit27.Q ),
    .A0(N2END[4]),
    .A1(NN4END[4]),
    .A2(N4END[4]),
    .A3(NN4END[12]),
    .S1(\Inst_N_IO4_ConfigMem.Inst_frame3_bit26.Q ),
    .X(\Inst_N_IO4_switch_matrix.S2BEGb3 ));
 sg13g2_mux4_1 _217_ (.S0(\Inst_N_IO4_ConfigMem.Inst_frame3_bit25.Q ),
    .A0(N2END[5]),
    .A1(NN4END[5]),
    .A2(N4END[5]),
    .A3(NN4END[13]),
    .S1(\Inst_N_IO4_ConfigMem.Inst_frame3_bit24.Q ),
    .X(\Inst_N_IO4_switch_matrix.S2BEGb2 ));
 sg13g2_mux4_1 _218_ (.S0(\Inst_N_IO4_ConfigMem.Inst_frame3_bit23.Q ),
    .A0(N2END[6]),
    .A1(NN4END[6]),
    .A2(N4END[6]),
    .A3(NN4END[14]),
    .S1(\Inst_N_IO4_ConfigMem.Inst_frame3_bit22.Q ),
    .X(\Inst_N_IO4_switch_matrix.S2BEGb1 ));
 sg13g2_mux4_1 _219_ (.S0(\Inst_N_IO4_ConfigMem.Inst_frame3_bit21.Q ),
    .A0(N2END[7]),
    .A1(NN4END[7]),
    .A2(N4END[7]),
    .A3(NN4END[15]),
    .S1(\Inst_N_IO4_ConfigMem.Inst_frame3_bit20.Q ),
    .X(\Inst_N_IO4_switch_matrix.S2BEGb0 ));
 sg13g2_mux4_1 _220_ (.S0(\Inst_N_IO4_ConfigMem.Inst_frame3_bit18.Q ),
    .A0(N2MID[0]),
    .A1(N4END[0]),
    .A2(NN4END[0]),
    .A3(NN4END[8]),
    .S1(\Inst_N_IO4_ConfigMem.Inst_frame3_bit19.Q ),
    .X(\Inst_N_IO4_switch_matrix.S2BEG7 ));
 sg13g2_mux4_1 _221_ (.S0(\Inst_N_IO4_ConfigMem.Inst_frame3_bit16.Q ),
    .A0(N2MID[1]),
    .A1(N4END[1]),
    .A2(NN4END[1]),
    .A3(NN4END[9]),
    .S1(\Inst_N_IO4_ConfigMem.Inst_frame3_bit17.Q ),
    .X(\Inst_N_IO4_switch_matrix.S2BEG6 ));
 sg13g2_dlhq_1 _222_ (.D(FrameData[28]),
    .GATE(FrameStrobe[4]),
    .Q(\Inst_N_IO4_ConfigMem.Inst_frame4_bit28.Q ));
 sg13g2_dlhq_1 _223_ (.D(FrameData[29]),
    .GATE(FrameStrobe[4]),
    .Q(\Inst_N_IO4_ConfigMem.Inst_frame4_bit29.Q ));
 sg13g2_dlhq_1 _224_ (.D(FrameData[30]),
    .GATE(FrameStrobe[4]),
    .Q(\Inst_N_IO4_ConfigMem.Inst_frame4_bit30.Q ));
 sg13g2_dlhq_1 _225_ (.D(FrameData[31]),
    .GATE(FrameStrobe[4]),
    .Q(\Inst_N_IO4_ConfigMem.Inst_frame4_bit31.Q ));
 sg13g2_dlhq_1 _226_ (.D(FrameData[0]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_N_IO4_ConfigMem.Inst_frame3_bit0.Q ));
 sg13g2_dlhq_1 _227_ (.D(FrameData[1]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_N_IO4_ConfigMem.Inst_frame3_bit1.Q ));
 sg13g2_dlhq_1 _228_ (.D(FrameData[2]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_N_IO4_ConfigMem.Inst_frame3_bit2.Q ));
 sg13g2_dlhq_1 _229_ (.D(FrameData[3]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_N_IO4_ConfigMem.Inst_frame3_bit3.Q ));
 sg13g2_dlhq_1 _230_ (.D(FrameData[4]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_N_IO4_ConfigMem.Inst_frame3_bit4.Q ));
 sg13g2_dlhq_1 _231_ (.D(FrameData[5]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_N_IO4_ConfigMem.Inst_frame3_bit5.Q ));
 sg13g2_dlhq_1 _232_ (.D(FrameData[6]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_N_IO4_ConfigMem.Inst_frame3_bit6.Q ));
 sg13g2_dlhq_1 _233_ (.D(FrameData[7]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_N_IO4_ConfigMem.Inst_frame3_bit7.Q ));
 sg13g2_dlhq_1 _234_ (.D(FrameData[8]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_N_IO4_ConfigMem.Inst_frame3_bit8.Q ));
 sg13g2_dlhq_1 _235_ (.D(FrameData[9]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_N_IO4_ConfigMem.Inst_frame3_bit9.Q ));
 sg13g2_dlhq_1 _236_ (.D(FrameData[10]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_N_IO4_ConfigMem.Inst_frame3_bit10.Q ));
 sg13g2_dlhq_1 _237_ (.D(FrameData[11]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_N_IO4_ConfigMem.Inst_frame3_bit11.Q ));
 sg13g2_dlhq_1 _238_ (.D(FrameData[12]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_N_IO4_ConfigMem.Inst_frame3_bit12.Q ));
 sg13g2_dlhq_1 _239_ (.D(FrameData[13]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_N_IO4_ConfigMem.Inst_frame3_bit13.Q ));
 sg13g2_dlhq_1 _240_ (.D(FrameData[14]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_N_IO4_ConfigMem.Inst_frame3_bit14.Q ));
 sg13g2_dlhq_1 _241_ (.D(FrameData[15]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_N_IO4_ConfigMem.Inst_frame3_bit15.Q ));
 sg13g2_dlhq_1 _242_ (.D(FrameData[16]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_N_IO4_ConfigMem.Inst_frame3_bit16.Q ));
 sg13g2_dlhq_1 _243_ (.D(FrameData[17]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_N_IO4_ConfigMem.Inst_frame3_bit17.Q ));
 sg13g2_dlhq_1 _244_ (.D(FrameData[18]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_N_IO4_ConfigMem.Inst_frame3_bit18.Q ));
 sg13g2_dlhq_1 _245_ (.D(FrameData[19]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_N_IO4_ConfigMem.Inst_frame3_bit19.Q ));
 sg13g2_dlhq_1 _246_ (.D(FrameData[20]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_N_IO4_ConfigMem.Inst_frame3_bit20.Q ));
 sg13g2_dlhq_1 _247_ (.D(FrameData[21]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_N_IO4_ConfigMem.Inst_frame3_bit21.Q ));
 sg13g2_dlhq_1 _248_ (.D(FrameData[22]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_N_IO4_ConfigMem.Inst_frame3_bit22.Q ));
 sg13g2_dlhq_1 _249_ (.D(FrameData[23]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_N_IO4_ConfigMem.Inst_frame3_bit23.Q ));
 sg13g2_dlhq_1 _250_ (.D(FrameData[24]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_N_IO4_ConfigMem.Inst_frame3_bit24.Q ));
 sg13g2_dlhq_1 _251_ (.D(FrameData[25]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_N_IO4_ConfigMem.Inst_frame3_bit25.Q ));
 sg13g2_dlhq_1 _252_ (.D(FrameData[26]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_N_IO4_ConfigMem.Inst_frame3_bit26.Q ));
 sg13g2_dlhq_1 _253_ (.D(FrameData[27]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_N_IO4_ConfigMem.Inst_frame3_bit27.Q ));
 sg13g2_dlhq_1 _254_ (.D(FrameData[28]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_N_IO4_ConfigMem.Inst_frame3_bit28.Q ));
 sg13g2_dlhq_1 _255_ (.D(FrameData[29]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_N_IO4_ConfigMem.Inst_frame3_bit29.Q ));
 sg13g2_dlhq_1 _256_ (.D(FrameData[30]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_N_IO4_ConfigMem.Inst_frame3_bit30.Q ));
 sg13g2_dlhq_1 _257_ (.D(FrameData[31]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_N_IO4_ConfigMem.Inst_frame3_bit31.Q ));
 sg13g2_dlhq_1 _258_ (.D(FrameData[0]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_N_IO4_ConfigMem.Inst_frame2_bit0.Q ));
 sg13g2_dlhq_1 _259_ (.D(FrameData[1]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_N_IO4_ConfigMem.Inst_frame2_bit1.Q ));
 sg13g2_dlhq_1 _260_ (.D(FrameData[2]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_N_IO4_ConfigMem.Inst_frame2_bit2.Q ));
 sg13g2_dlhq_1 _261_ (.D(FrameData[3]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_N_IO4_ConfigMem.Inst_frame2_bit3.Q ));
 sg13g2_dlhq_1 _262_ (.D(FrameData[4]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_N_IO4_ConfigMem.Inst_frame2_bit4.Q ));
 sg13g2_dlhq_1 _263_ (.D(FrameData[5]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_N_IO4_ConfigMem.Inst_frame2_bit5.Q ));
 sg13g2_dlhq_1 _264_ (.D(FrameData[6]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_N_IO4_ConfigMem.Inst_frame2_bit6.Q ));
 sg13g2_dlhq_1 _265_ (.D(FrameData[7]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_N_IO4_ConfigMem.Inst_frame2_bit7.Q ));
 sg13g2_dlhq_1 _266_ (.D(FrameData[8]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_N_IO4_ConfigMem.Inst_frame2_bit8.Q ));
 sg13g2_dlhq_1 _267_ (.D(FrameData[9]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_N_IO4_ConfigMem.Inst_frame2_bit9.Q ));
 sg13g2_dlhq_1 _268_ (.D(FrameData[10]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_N_IO4_ConfigMem.Inst_frame2_bit10.Q ));
 sg13g2_dlhq_1 _269_ (.D(FrameData[11]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_N_IO4_ConfigMem.Inst_frame2_bit11.Q ));
 sg13g2_dlhq_1 _270_ (.D(FrameData[12]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_N_IO4_ConfigMem.Inst_frame2_bit12.Q ));
 sg13g2_dlhq_1 _271_ (.D(FrameData[13]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_N_IO4_ConfigMem.Inst_frame2_bit13.Q ));
 sg13g2_dlhq_1 _272_ (.D(FrameData[14]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_N_IO4_ConfigMem.Inst_frame2_bit14.Q ));
 sg13g2_dlhq_1 _273_ (.D(FrameData[15]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_N_IO4_ConfigMem.Inst_frame2_bit15.Q ));
 sg13g2_dlhq_1 _274_ (.D(FrameData[16]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_N_IO4_ConfigMem.Inst_frame2_bit16.Q ));
 sg13g2_dlhq_1 _275_ (.D(FrameData[17]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_N_IO4_ConfigMem.Inst_frame2_bit17.Q ));
 sg13g2_dlhq_1 _276_ (.D(FrameData[18]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_N_IO4_ConfigMem.Inst_frame2_bit18.Q ));
 sg13g2_dlhq_1 _277_ (.D(FrameData[19]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_N_IO4_ConfigMem.Inst_frame2_bit19.Q ));
 sg13g2_dlhq_1 _278_ (.D(FrameData[20]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_N_IO4_ConfigMem.Inst_frame2_bit20.Q ));
 sg13g2_dlhq_1 _279_ (.D(FrameData[21]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_N_IO4_ConfigMem.Inst_frame2_bit21.Q ));
 sg13g2_dlhq_1 _280_ (.D(FrameData[22]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_N_IO4_ConfigMem.Inst_frame2_bit22.Q ));
 sg13g2_dlhq_1 _281_ (.D(FrameData[23]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_N_IO4_ConfigMem.Inst_frame2_bit23.Q ));
 sg13g2_dlhq_1 _282_ (.D(FrameData[24]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_N_IO4_ConfigMem.Inst_frame2_bit24.Q ));
 sg13g2_dlhq_1 _283_ (.D(FrameData[25]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_N_IO4_ConfigMem.Inst_frame2_bit25.Q ));
 sg13g2_dlhq_1 _284_ (.D(FrameData[26]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_N_IO4_ConfigMem.Inst_frame2_bit26.Q ));
 sg13g2_dlhq_1 _285_ (.D(FrameData[27]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_N_IO4_ConfigMem.Inst_frame2_bit27.Q ));
 sg13g2_dlhq_1 _286_ (.D(FrameData[28]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_N_IO4_ConfigMem.Inst_frame2_bit28.Q ));
 sg13g2_dlhq_1 _287_ (.D(FrameData[29]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_N_IO4_ConfigMem.Inst_frame2_bit29.Q ));
 sg13g2_dlhq_1 _288_ (.D(FrameData[30]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_N_IO4_ConfigMem.Inst_frame2_bit30.Q ));
 sg13g2_dlhq_1 _289_ (.D(FrameData[31]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_N_IO4_ConfigMem.Inst_frame2_bit31.Q ));
 sg13g2_dlhq_1 _290_ (.D(FrameData[0]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_N_IO4_ConfigMem.Inst_frame1_bit0.Q ));
 sg13g2_dlhq_1 _291_ (.D(FrameData[1]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_N_IO4_ConfigMem.Inst_frame1_bit1.Q ));
 sg13g2_dlhq_1 _292_ (.D(FrameData[2]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_N_IO4_ConfigMem.Inst_frame1_bit2.Q ));
 sg13g2_dlhq_1 _293_ (.D(FrameData[3]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_N_IO4_ConfigMem.Inst_frame1_bit3.Q ));
 sg13g2_dlhq_1 _294_ (.D(FrameData[4]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_N_IO4_ConfigMem.Inst_frame1_bit4.Q ));
 sg13g2_dlhq_1 _295_ (.D(FrameData[5]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_N_IO4_ConfigMem.Inst_frame1_bit5.Q ));
 sg13g2_dlhq_1 _296_ (.D(FrameData[6]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_N_IO4_ConfigMem.Inst_frame1_bit6.Q ));
 sg13g2_dlhq_1 _297_ (.D(FrameData[7]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_N_IO4_ConfigMem.Inst_frame1_bit7.Q ));
 sg13g2_dlhq_1 _298_ (.D(FrameData[8]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_N_IO4_ConfigMem.Inst_frame1_bit8.Q ));
 sg13g2_dlhq_1 _299_ (.D(FrameData[9]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_N_IO4_ConfigMem.Inst_frame1_bit9.Q ));
 sg13g2_dlhq_1 _300_ (.D(FrameData[10]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_N_IO4_ConfigMem.Inst_frame1_bit10.Q ));
 sg13g2_dlhq_1 _301_ (.D(FrameData[11]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_N_IO4_ConfigMem.Inst_frame1_bit11.Q ));
 sg13g2_dlhq_1 _302_ (.D(FrameData[12]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_N_IO4_ConfigMem.Inst_frame1_bit12.Q ));
 sg13g2_dlhq_1 _303_ (.D(FrameData[13]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_N_IO4_ConfigMem.Inst_frame1_bit13.Q ));
 sg13g2_dlhq_1 _304_ (.D(FrameData[14]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_N_IO4_ConfigMem.Inst_frame1_bit14.Q ));
 sg13g2_dlhq_1 _305_ (.D(FrameData[15]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_N_IO4_ConfigMem.Inst_frame1_bit15.Q ));
 sg13g2_dlhq_1 _306_ (.D(FrameData[16]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_N_IO4_ConfigMem.Inst_frame1_bit16.Q ));
 sg13g2_dlhq_1 _307_ (.D(FrameData[17]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_N_IO4_ConfigMem.Inst_frame1_bit17.Q ));
 sg13g2_dlhq_1 _308_ (.D(FrameData[18]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_N_IO4_ConfigMem.Inst_frame1_bit18.Q ));
 sg13g2_dlhq_1 _309_ (.D(FrameData[19]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_N_IO4_ConfigMem.Inst_frame1_bit19.Q ));
 sg13g2_dlhq_1 _310_ (.D(FrameData[20]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_N_IO4_ConfigMem.Inst_frame1_bit20.Q ));
 sg13g2_dlhq_1 _311_ (.D(FrameData[21]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_N_IO4_ConfigMem.Inst_frame1_bit21.Q ));
 sg13g2_dlhq_1 _312_ (.D(FrameData[22]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_N_IO4_ConfigMem.Inst_frame1_bit22.Q ));
 sg13g2_dlhq_1 _313_ (.D(FrameData[23]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_N_IO4_ConfigMem.Inst_frame1_bit23.Q ));
 sg13g2_dlhq_1 _314_ (.D(FrameData[24]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_N_IO4_ConfigMem.Inst_frame1_bit24.Q ));
 sg13g2_dlhq_1 _315_ (.D(FrameData[25]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_N_IO4_ConfigMem.Inst_frame1_bit25.Q ));
 sg13g2_dlhq_1 _316_ (.D(FrameData[26]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_N_IO4_ConfigMem.Inst_frame1_bit26.Q ));
 sg13g2_dlhq_1 _317_ (.D(FrameData[27]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_N_IO4_ConfigMem.Inst_frame1_bit27.Q ));
 sg13g2_dlhq_1 _318_ (.D(FrameData[28]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_N_IO4_ConfigMem.Inst_frame1_bit28.Q ));
 sg13g2_dlhq_1 _319_ (.D(FrameData[29]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_N_IO4_ConfigMem.Inst_frame1_bit29.Q ));
 sg13g2_dlhq_1 _320_ (.D(FrameData[30]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_N_IO4_ConfigMem.Inst_frame1_bit30.Q ));
 sg13g2_dlhq_1 _321_ (.D(FrameData[31]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_N_IO4_ConfigMem.Inst_frame1_bit31.Q ));
 sg13g2_dlhq_1 _322_ (.D(FrameData[0]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_N_IO4_ConfigMem.Inst_frame0_bit0.Q ));
 sg13g2_dlhq_1 _323_ (.D(FrameData[1]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_N_IO4_ConfigMem.Inst_frame0_bit1.Q ));
 sg13g2_dlhq_1 _324_ (.D(FrameData[2]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_N_IO4_ConfigMem.Inst_frame0_bit2.Q ));
 sg13g2_dlhq_1 _325_ (.D(FrameData[3]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_N_IO4_ConfigMem.Inst_frame0_bit3.Q ));
 sg13g2_dlhq_1 _326_ (.D(FrameData[4]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_N_IO4_ConfigMem.Inst_frame0_bit4.Q ));
 sg13g2_dlhq_1 _327_ (.D(FrameData[5]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_N_IO4_ConfigMem.Inst_frame0_bit5.Q ));
 sg13g2_dlhq_1 _328_ (.D(FrameData[6]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_N_IO4_ConfigMem.Inst_frame0_bit6.Q ));
 sg13g2_dlhq_1 _329_ (.D(FrameData[7]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_N_IO4_ConfigMem.Inst_frame0_bit7.Q ));
 sg13g2_dlhq_1 _330_ (.D(FrameData[8]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_N_IO4_ConfigMem.Inst_frame0_bit8.Q ));
 sg13g2_dlhq_1 _331_ (.D(FrameData[9]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_N_IO4_ConfigMem.Inst_frame0_bit9.Q ));
 sg13g2_dlhq_1 _332_ (.D(FrameData[10]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_N_IO4_ConfigMem.Inst_frame0_bit10.Q ));
 sg13g2_dlhq_1 _333_ (.D(FrameData[11]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_N_IO4_ConfigMem.Inst_frame0_bit11.Q ));
 sg13g2_dlhq_1 _334_ (.D(FrameData[12]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_N_IO4_ConfigMem.Inst_frame0_bit12.Q ));
 sg13g2_dlhq_1 _335_ (.D(FrameData[13]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_N_IO4_ConfigMem.Inst_frame0_bit13.Q ));
 sg13g2_dlhq_1 _336_ (.D(FrameData[14]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_N_IO4_ConfigMem.Inst_frame0_bit14.Q ));
 sg13g2_dlhq_1 _337_ (.D(FrameData[15]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_N_IO4_ConfigMem.Inst_frame0_bit15.Q ));
 sg13g2_dlhq_1 _338_ (.D(FrameData[16]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_N_IO4_ConfigMem.Inst_frame0_bit16.Q ));
 sg13g2_dlhq_1 _339_ (.D(FrameData[17]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_N_IO4_ConfigMem.Inst_frame0_bit17.Q ));
 sg13g2_dlhq_1 _340_ (.D(FrameData[18]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_N_IO4_ConfigMem.Inst_frame0_bit18.Q ));
 sg13g2_dlhq_1 _341_ (.D(FrameData[19]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_N_IO4_ConfigMem.Inst_frame0_bit19.Q ));
 sg13g2_dlhq_1 _342_ (.D(FrameData[20]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_N_IO4_ConfigMem.Inst_frame0_bit20.Q ));
 sg13g2_dlhq_1 _343_ (.D(FrameData[21]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_N_IO4_ConfigMem.Inst_frame0_bit21.Q ));
 sg13g2_dlhq_1 _344_ (.D(FrameData[22]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_N_IO4_ConfigMem.Inst_frame0_bit22.Q ));
 sg13g2_dlhq_1 _345_ (.D(FrameData[23]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_N_IO4_ConfigMem.Inst_frame0_bit23.Q ));
 sg13g2_dlhq_1 _346_ (.D(FrameData[24]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_N_IO4_ConfigMem.Inst_frame0_bit24.Q ));
 sg13g2_dlhq_1 _347_ (.D(FrameData[25]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_N_IO4_ConfigMem.Inst_frame0_bit25.Q ));
 sg13g2_dlhq_1 _348_ (.D(FrameData[26]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_N_IO4_ConfigMem.Inst_frame0_bit26.Q ));
 sg13g2_dlhq_1 _349_ (.D(FrameData[27]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_N_IO4_ConfigMem.Inst_frame0_bit27.Q ));
 sg13g2_dlhq_1 _350_ (.D(FrameData[28]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_N_IO4_ConfigMem.Inst_frame0_bit28.Q ));
 sg13g2_dlhq_1 _351_ (.D(FrameData[29]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_N_IO4_ConfigMem.Inst_frame0_bit29.Q ));
 sg13g2_dlhq_1 _352_ (.D(FrameData[30]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_N_IO4_ConfigMem.Inst_frame0_bit30.Q ));
 sg13g2_dlhq_1 _353_ (.D(FrameData[31]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_N_IO4_ConfigMem.Inst_frame0_bit31.Q ));
 sg13g2_dfrbpq_1 _354_ (.RESET_B(_081_),
    .D(A_O_top),
    .Q(\Inst_A_IO_1_bidirectional_frame_config_pass.Q ),
    .CLK(clknet_1_0__leaf_UserCLK_regs));
 sg13g2_dfrbpq_1 _355_ (.RESET_B(_082_),
    .D(B_O_top),
    .Q(\Inst_B_IO_1_bidirectional_frame_config_pass.Q ),
    .CLK(clknet_1_1__leaf_UserCLK_regs));
 sg13g2_dfrbpq_1 _356_ (.RESET_B(_079_),
    .D(C_O_top),
    .Q(\Inst_C_IO_1_bidirectional_frame_config_pass.Q ),
    .CLK(clknet_1_0__leaf_UserCLK_regs));
 sg13g2_dfrbpq_1 _357_ (.RESET_B(_080_),
    .D(D_O_top),
    .Q(\Inst_D_IO_1_bidirectional_frame_config_pass.Q ),
    .CLK(clknet_1_1__leaf_UserCLK_regs));
 sg13g2_tiehi _358_ (.L_HI(_079_));
 sg13g2_tiehi _359_ (.L_HI(_080_));
 sg13g2_tiehi _360_ (.L_HI(_081_));
 sg13g2_tiehi _361_ (.L_HI(_082_));
 sg13g2_buf_1 _362_ (.A(FrameData[0]),
    .X(FrameData_O[0]));
 sg13g2_buf_1 _363_ (.A(FrameData[1]),
    .X(FrameData_O[1]));
 sg13g2_buf_1 _364_ (.A(FrameData[2]),
    .X(FrameData_O[2]));
 sg13g2_buf_1 _365_ (.A(FrameData[3]),
    .X(FrameData_O[3]));
 sg13g2_buf_1 _366_ (.A(FrameData[4]),
    .X(FrameData_O[4]));
 sg13g2_buf_1 _367_ (.A(FrameData[5]),
    .X(FrameData_O[5]));
 sg13g2_buf_1 _368_ (.A(FrameData[6]),
    .X(FrameData_O[6]));
 sg13g2_buf_1 _369_ (.A(FrameData[7]),
    .X(FrameData_O[7]));
 sg13g2_buf_1 _370_ (.A(FrameData[8]),
    .X(FrameData_O[8]));
 sg13g2_buf_1 _371_ (.A(FrameData[9]),
    .X(FrameData_O[9]));
 sg13g2_buf_1 _372_ (.A(FrameData[10]),
    .X(FrameData_O[10]));
 sg13g2_buf_1 _373_ (.A(FrameData[11]),
    .X(FrameData_O[11]));
 sg13g2_buf_1 _374_ (.A(FrameData[12]),
    .X(FrameData_O[12]));
 sg13g2_buf_1 _375_ (.A(FrameData[13]),
    .X(FrameData_O[13]));
 sg13g2_buf_1 _376_ (.A(FrameData[14]),
    .X(FrameData_O[14]));
 sg13g2_buf_1 _377_ (.A(FrameData[15]),
    .X(FrameData_O[15]));
 sg13g2_buf_1 _378_ (.A(FrameData[16]),
    .X(FrameData_O[16]));
 sg13g2_buf_1 _379_ (.A(FrameData[17]),
    .X(FrameData_O[17]));
 sg13g2_buf_1 _380_ (.A(FrameData[18]),
    .X(FrameData_O[18]));
 sg13g2_buf_1 _381_ (.A(FrameData[19]),
    .X(FrameData_O[19]));
 sg13g2_buf_1 _382_ (.A(FrameData[20]),
    .X(FrameData_O[20]));
 sg13g2_buf_1 _383_ (.A(FrameData[21]),
    .X(FrameData_O[21]));
 sg13g2_buf_1 _384_ (.A(FrameData[22]),
    .X(FrameData_O[22]));
 sg13g2_buf_1 _385_ (.A(FrameData[23]),
    .X(FrameData_O[23]));
 sg13g2_buf_1 _386_ (.A(FrameData[24]),
    .X(FrameData_O[24]));
 sg13g2_buf_1 _387_ (.A(FrameData[25]),
    .X(FrameData_O[25]));
 sg13g2_buf_1 _388_ (.A(FrameData[26]),
    .X(FrameData_O[26]));
 sg13g2_buf_1 _389_ (.A(FrameData[27]),
    .X(FrameData_O[27]));
 sg13g2_buf_1 _390_ (.A(FrameData[28]),
    .X(FrameData_O[28]));
 sg13g2_buf_1 _391_ (.A(FrameData[29]),
    .X(FrameData_O[29]));
 sg13g2_buf_1 _392_ (.A(FrameData[30]),
    .X(FrameData_O[30]));
 sg13g2_buf_1 _393_ (.A(FrameData[31]),
    .X(FrameData_O[31]));
 sg13g2_buf_1 _394_ (.A(FrameStrobe[0]),
    .X(FrameStrobe_O[0]));
 sg13g2_buf_1 _395_ (.A(FrameStrobe[1]),
    .X(FrameStrobe_O[1]));
 sg13g2_buf_1 _396_ (.A(FrameStrobe[2]),
    .X(FrameStrobe_O[2]));
 sg13g2_buf_1 _397_ (.A(FrameStrobe[3]),
    .X(FrameStrobe_O[3]));
 sg13g2_buf_1 _398_ (.A(FrameStrobe[4]),
    .X(FrameStrobe_O[4]));
 sg13g2_buf_1 _399_ (.A(FrameStrobe[5]),
    .X(FrameStrobe_O[5]));
 sg13g2_buf_1 _400_ (.A(FrameStrobe[6]),
    .X(FrameStrobe_O[6]));
 sg13g2_buf_1 _401_ (.A(FrameStrobe[7]),
    .X(FrameStrobe_O[7]));
 sg13g2_buf_1 _402_ (.A(FrameStrobe[8]),
    .X(FrameStrobe_O[8]));
 sg13g2_buf_1 _403_ (.A(FrameStrobe[9]),
    .X(FrameStrobe_O[9]));
 sg13g2_buf_1 _404_ (.A(FrameStrobe[10]),
    .X(FrameStrobe_O[10]));
 sg13g2_buf_1 _405_ (.A(FrameStrobe[11]),
    .X(FrameStrobe_O[11]));
 sg13g2_buf_1 _406_ (.A(FrameStrobe[12]),
    .X(FrameStrobe_O[12]));
 sg13g2_buf_1 _407_ (.A(FrameStrobe[13]),
    .X(FrameStrobe_O[13]));
 sg13g2_buf_1 _408_ (.A(FrameStrobe[14]),
    .X(FrameStrobe_O[14]));
 sg13g2_buf_1 _409_ (.A(FrameStrobe[15]),
    .X(FrameStrobe_O[15]));
 sg13g2_buf_1 _410_ (.A(FrameStrobe[16]),
    .X(FrameStrobe_O[16]));
 sg13g2_buf_1 _411_ (.A(FrameStrobe[17]),
    .X(FrameStrobe_O[17]));
 sg13g2_buf_1 _412_ (.A(FrameStrobe[18]),
    .X(FrameStrobe_O[18]));
 sg13g2_buf_1 _413_ (.A(FrameStrobe[19]),
    .X(FrameStrobe_O[19]));
 sg13g2_buf_1 _414_ (.A(\Inst_N_IO4_switch_matrix.S1BEG0 ),
    .X(S1BEG[0]));
 sg13g2_buf_1 _415_ (.A(\Inst_N_IO4_switch_matrix.S1BEG1 ),
    .X(S1BEG[1]));
 sg13g2_buf_1 _416_ (.A(\Inst_N_IO4_switch_matrix.S1BEG2 ),
    .X(S1BEG[2]));
 sg13g2_buf_1 _417_ (.A(\Inst_N_IO4_switch_matrix.S1BEG3 ),
    .X(S1BEG[3]));
 sg13g2_buf_1 _418_ (.A(\Inst_N_IO4_switch_matrix.S2BEG0 ),
    .X(S2BEG[0]));
 sg13g2_buf_1 _419_ (.A(\Inst_N_IO4_switch_matrix.S2BEG1 ),
    .X(S2BEG[1]));
 sg13g2_buf_1 _420_ (.A(\Inst_N_IO4_switch_matrix.S2BEG2 ),
    .X(S2BEG[2]));
 sg13g2_buf_1 _421_ (.A(\Inst_N_IO4_switch_matrix.S2BEG3 ),
    .X(S2BEG[3]));
 sg13g2_buf_1 _422_ (.A(\Inst_N_IO4_switch_matrix.S2BEG4 ),
    .X(S2BEG[4]));
 sg13g2_buf_1 _423_ (.A(\Inst_N_IO4_switch_matrix.S2BEG5 ),
    .X(S2BEG[5]));
 sg13g2_buf_1 _424_ (.A(\Inst_N_IO4_switch_matrix.S2BEG6 ),
    .X(S2BEG[6]));
 sg13g2_buf_1 _425_ (.A(\Inst_N_IO4_switch_matrix.S2BEG7 ),
    .X(S2BEG[7]));
 sg13g2_buf_1 _426_ (.A(\Inst_N_IO4_switch_matrix.S2BEGb0 ),
    .X(S2BEGb[0]));
 sg13g2_buf_1 _427_ (.A(\Inst_N_IO4_switch_matrix.S2BEGb1 ),
    .X(S2BEGb[1]));
 sg13g2_buf_1 _428_ (.A(\Inst_N_IO4_switch_matrix.S2BEGb2 ),
    .X(S2BEGb[2]));
 sg13g2_buf_1 _429_ (.A(\Inst_N_IO4_switch_matrix.S2BEGb3 ),
    .X(S2BEGb[3]));
 sg13g2_buf_1 _430_ (.A(\Inst_N_IO4_switch_matrix.S2BEGb4 ),
    .X(S2BEGb[4]));
 sg13g2_buf_1 _431_ (.A(\Inst_N_IO4_switch_matrix.S2BEGb5 ),
    .X(S2BEGb[5]));
 sg13g2_buf_1 _432_ (.A(\Inst_N_IO4_switch_matrix.S2BEGb6 ),
    .X(S2BEGb[6]));
 sg13g2_buf_1 _433_ (.A(\Inst_N_IO4_switch_matrix.S2BEGb7 ),
    .X(S2BEGb[7]));
 sg13g2_buf_1 _434_ (.A(\Inst_N_IO4_switch_matrix.S4BEG0 ),
    .X(S4BEG[0]));
 sg13g2_buf_1 _435_ (.A(\Inst_N_IO4_switch_matrix.S4BEG1 ),
    .X(S4BEG[1]));
 sg13g2_buf_1 _436_ (.A(\Inst_N_IO4_switch_matrix.S4BEG2 ),
    .X(S4BEG[2]));
 sg13g2_buf_1 _437_ (.A(\Inst_N_IO4_switch_matrix.S4BEG3 ),
    .X(S4BEG[3]));
 sg13g2_buf_1 _438_ (.A(\Inst_N_IO4_switch_matrix.S4BEG4 ),
    .X(S4BEG[4]));
 sg13g2_buf_1 _439_ (.A(\Inst_N_IO4_switch_matrix.S4BEG5 ),
    .X(S4BEG[5]));
 sg13g2_buf_1 _440_ (.A(\Inst_N_IO4_switch_matrix.S4BEG6 ),
    .X(S4BEG[6]));
 sg13g2_buf_1 _441_ (.A(\Inst_N_IO4_switch_matrix.S4BEG7 ),
    .X(S4BEG[7]));
 sg13g2_buf_1 _442_ (.A(\Inst_N_IO4_switch_matrix.S4BEG8 ),
    .X(S4BEG[8]));
 sg13g2_buf_1 _443_ (.A(\Inst_N_IO4_switch_matrix.S4BEG9 ),
    .X(S4BEG[9]));
 sg13g2_buf_1 _444_ (.A(\Inst_N_IO4_switch_matrix.S4BEG10 ),
    .X(S4BEG[10]));
 sg13g2_buf_1 _445_ (.A(\Inst_N_IO4_switch_matrix.S4BEG11 ),
    .X(S4BEG[11]));
 sg13g2_buf_1 _446_ (.A(\Inst_N_IO4_switch_matrix.S4BEG12 ),
    .X(S4BEG[12]));
 sg13g2_buf_1 _447_ (.A(\Inst_N_IO4_switch_matrix.S4BEG13 ),
    .X(S4BEG[13]));
 sg13g2_buf_1 _448_ (.A(\Inst_N_IO4_switch_matrix.S4BEG14 ),
    .X(S4BEG[14]));
 sg13g2_buf_1 _449_ (.A(\Inst_N_IO4_switch_matrix.S4BEG15 ),
    .X(S4BEG[15]));
 sg13g2_buf_1 _450_ (.A(\Inst_N_IO4_switch_matrix.SS4BEG0 ),
    .X(SS4BEG[0]));
 sg13g2_buf_1 _451_ (.A(\Inst_N_IO4_switch_matrix.SS4BEG1 ),
    .X(SS4BEG[1]));
 sg13g2_buf_1 _452_ (.A(\Inst_N_IO4_switch_matrix.SS4BEG2 ),
    .X(SS4BEG[2]));
 sg13g2_buf_1 _453_ (.A(\Inst_N_IO4_switch_matrix.SS4BEG3 ),
    .X(SS4BEG[3]));
 sg13g2_buf_1 _454_ (.A(\Inst_N_IO4_switch_matrix.SS4BEG4 ),
    .X(SS4BEG[4]));
 sg13g2_buf_1 _455_ (.A(\Inst_N_IO4_switch_matrix.SS4BEG5 ),
    .X(SS4BEG[5]));
 sg13g2_buf_1 _456_ (.A(\Inst_N_IO4_switch_matrix.SS4BEG6 ),
    .X(SS4BEG[6]));
 sg13g2_buf_1 _457_ (.A(\Inst_N_IO4_switch_matrix.SS4BEG7 ),
    .X(SS4BEG[7]));
 sg13g2_buf_1 _458_ (.A(\Inst_N_IO4_switch_matrix.SS4BEG8 ),
    .X(SS4BEG[8]));
 sg13g2_buf_1 _459_ (.A(\Inst_N_IO4_switch_matrix.SS4BEG9 ),
    .X(SS4BEG[9]));
 sg13g2_buf_1 _460_ (.A(\Inst_N_IO4_switch_matrix.SS4BEG10 ),
    .X(SS4BEG[10]));
 sg13g2_buf_1 _461_ (.A(\Inst_N_IO4_switch_matrix.SS4BEG11 ),
    .X(SS4BEG[11]));
 sg13g2_buf_1 _462_ (.A(\Inst_N_IO4_switch_matrix.SS4BEG12 ),
    .X(SS4BEG[12]));
 sg13g2_buf_1 _463_ (.A(\Inst_N_IO4_switch_matrix.SS4BEG13 ),
    .X(SS4BEG[13]));
 sg13g2_buf_1 _464_ (.A(\Inst_N_IO4_switch_matrix.SS4BEG14 ),
    .X(SS4BEG[14]));
 sg13g2_buf_1 _465_ (.A(\Inst_N_IO4_switch_matrix.SS4BEG15 ),
    .X(SS4BEG[15]));
 sg13g2_buf_1 _466_ (.A(clknet_1_0__leaf_UserCLK),
    .X(UserCLKo));
 sg13g2_buf_8 clkbuf_regs_0_UserCLK (.A(UserCLK),
    .X(UserCLK_regs));
 sg13g2_buf_8 clkbuf_0_UserCLK (.A(UserCLK),
    .X(clknet_0_UserCLK));
 sg13g2_buf_8 clkbuf_1_0__f_UserCLK (.A(clknet_0_UserCLK),
    .X(clknet_1_0__leaf_UserCLK));
 sg13g2_buf_8 clkbuf_0_UserCLK_regs (.A(UserCLK_regs),
    .X(clknet_0_UserCLK_regs));
 sg13g2_buf_8 clkbuf_1_0__f_UserCLK_regs (.A(clknet_0_UserCLK_regs),
    .X(clknet_1_0__leaf_UserCLK_regs));
 sg13g2_buf_8 clkbuf_1_1__f_UserCLK_regs (.A(clknet_0_UserCLK_regs),
    .X(clknet_1_1__leaf_UserCLK_regs));
 sg13g2_fill_1 FILLER_0_0 ();
 sg13g2_fill_1 FILLER_0_23 ();
 sg13g2_fill_2 FILLER_0_125 ();
 sg13g2_decap_8 FILLER_0_153 ();
 sg13g2_decap_8 FILLER_0_160 ();
 sg13g2_decap_8 FILLER_0_167 ();
 sg13g2_fill_2 FILLER_0_174 ();
 sg13g2_decap_8 FILLER_0_193 ();
 sg13g2_fill_2 FILLER_0_200 ();
 sg13g2_fill_1 FILLER_0_202 ();
 sg13g2_fill_2 FILLER_0_411 ();
 sg13g2_fill_2 FILLER_0_421 ();
 sg13g2_fill_1 FILLER_0_423 ();
 sg13g2_fill_1 FILLER_1_0 ();
 sg13g2_fill_2 FILLER_1_61 ();
 sg13g2_fill_1 FILLER_1_130 ();
 sg13g2_fill_2 FILLER_1_156 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_fill_2 FILLER_1_203 ();
 sg13g2_fill_1 FILLER_1_238 ();
 sg13g2_fill_2 FILLER_1_285 ();
 sg13g2_fill_1 FILLER_1_287 ();
 sg13g2_fill_1 FILLER_1_317 ();
 sg13g2_fill_1 FILLER_1_343 ();
 sg13g2_fill_1 FILLER_1_423 ();
 sg13g2_fill_1 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_157 ();
 sg13g2_decap_8 FILLER_2_164 ();
 sg13g2_decap_8 FILLER_2_171 ();
 sg13g2_decap_8 FILLER_2_178 ();
 sg13g2_decap_8 FILLER_2_185 ();
 sg13g2_decap_4 FILLER_2_192 ();
 sg13g2_fill_2 FILLER_2_213 ();
 sg13g2_fill_2 FILLER_2_257 ();
 sg13g2_fill_2 FILLER_2_348 ();
 sg13g2_fill_1 FILLER_2_350 ();
 sg13g2_fill_1 FILLER_2_423 ();
 sg13g2_fill_1 FILLER_3_51 ();
 sg13g2_fill_2 FILLER_3_79 ();
 sg13g2_decap_8 FILLER_3_144 ();
 sg13g2_fill_2 FILLER_3_151 ();
 sg13g2_fill_1 FILLER_3_153 ();
 sg13g2_decap_8 FILLER_3_188 ();
 sg13g2_fill_2 FILLER_3_199 ();
 sg13g2_decap_4 FILLER_3_218 ();
 sg13g2_fill_2 FILLER_3_222 ();
 sg13g2_fill_2 FILLER_3_245 ();
 sg13g2_fill_1 FILLER_3_247 ();
 sg13g2_fill_2 FILLER_3_277 ();
 sg13g2_fill_1 FILLER_3_279 ();
 sg13g2_fill_2 FILLER_3_301 ();
 sg13g2_fill_2 FILLER_3_328 ();
 sg13g2_fill_1 FILLER_3_330 ();
 sg13g2_fill_2 FILLER_3_369 ();
 sg13g2_fill_1 FILLER_3_371 ();
 sg13g2_fill_2 FILLER_3_421 ();
 sg13g2_fill_1 FILLER_3_423 ();
 sg13g2_fill_2 FILLER_4_0 ();
 sg13g2_fill_2 FILLER_4_71 ();
 sg13g2_decap_8 FILLER_4_155 ();
 sg13g2_decap_8 FILLER_4_162 ();
 sg13g2_decap_4 FILLER_4_190 ();
 sg13g2_fill_2 FILLER_4_194 ();
 sg13g2_decap_4 FILLER_4_234 ();
 sg13g2_fill_1 FILLER_4_238 ();
 sg13g2_fill_2 FILLER_4_277 ();
 sg13g2_fill_2 FILLER_4_317 ();
 sg13g2_fill_2 FILLER_4_348 ();
 sg13g2_fill_2 FILLER_4_379 ();
 sg13g2_fill_1 FILLER_4_402 ();
 sg13g2_fill_2 FILLER_4_411 ();
 sg13g2_fill_2 FILLER_4_421 ();
 sg13g2_fill_1 FILLER_4_423 ();
 sg13g2_fill_1 FILLER_5_0 ();
 sg13g2_fill_1 FILLER_5_18 ();
 sg13g2_fill_1 FILLER_5_34 ();
 sg13g2_fill_1 FILLER_5_95 ();
 sg13g2_decap_8 FILLER_5_135 ();
 sg13g2_decap_8 FILLER_5_180 ();
 sg13g2_decap_8 FILLER_5_187 ();
 sg13g2_decap_4 FILLER_5_194 ();
 sg13g2_decap_4 FILLER_5_202 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_234 ();
 sg13g2_fill_2 FILLER_5_241 ();
 sg13g2_decap_4 FILLER_5_260 ();
 sg13g2_fill_2 FILLER_5_289 ();
 sg13g2_fill_1 FILLER_5_291 ();
 sg13g2_fill_2 FILLER_5_330 ();
 sg13g2_fill_1 FILLER_5_332 ();
 sg13g2_fill_1 FILLER_5_358 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_fill_2 FILLER_5_421 ();
 sg13g2_fill_1 FILLER_5_423 ();
 sg13g2_fill_1 FILLER_6_71 ();
 sg13g2_fill_1 FILLER_6_100 ();
 sg13g2_decap_8 FILLER_6_139 ();
 sg13g2_decap_8 FILLER_6_146 ();
 sg13g2_fill_2 FILLER_6_153 ();
 sg13g2_fill_1 FILLER_6_155 ();
 sg13g2_decap_8 FILLER_6_194 ();
 sg13g2_fill_1 FILLER_6_222 ();
 sg13g2_decap_4 FILLER_6_231 ();
 sg13g2_fill_1 FILLER_6_235 ();
 sg13g2_decap_4 FILLER_6_265 ();
 sg13g2_fill_1 FILLER_6_269 ();
 sg13g2_fill_1 FILLER_6_274 ();
 sg13g2_fill_2 FILLER_6_321 ();
 sg13g2_fill_1 FILLER_6_348 ();
 sg13g2_fill_2 FILLER_6_370 ();
 sg13g2_fill_1 FILLER_6_372 ();
 sg13g2_decap_4 FILLER_6_398 ();
 sg13g2_fill_1 FILLER_6_402 ();
 sg13g2_fill_2 FILLER_6_407 ();
 sg13g2_fill_2 FILLER_6_421 ();
 sg13g2_fill_1 FILLER_6_423 ();
 sg13g2_fill_2 FILLER_7_22 ();
 sg13g2_fill_1 FILLER_7_54 ();
 sg13g2_fill_1 FILLER_7_86 ();
 sg13g2_fill_2 FILLER_7_104 ();
 sg13g2_fill_2 FILLER_7_149 ();
 sg13g2_fill_2 FILLER_7_172 ();
 sg13g2_fill_1 FILLER_7_174 ();
 sg13g2_decap_8 FILLER_7_200 ();
 sg13g2_fill_2 FILLER_7_245 ();
 sg13g2_decap_4 FILLER_7_264 ();
 sg13g2_fill_1 FILLER_7_306 ();
 sg13g2_fill_2 FILLER_7_374 ();
 sg13g2_fill_2 FILLER_7_393 ();
 sg13g2_fill_1 FILLER_7_412 ();
 sg13g2_fill_2 FILLER_7_421 ();
 sg13g2_fill_1 FILLER_7_423 ();
 sg13g2_fill_1 FILLER_8_59 ();
 sg13g2_decap_4 FILLER_8_107 ();
 sg13g2_decap_4 FILLER_8_206 ();
 sg13g2_fill_1 FILLER_8_256 ();
 sg13g2_fill_2 FILLER_8_328 ();
 sg13g2_fill_2 FILLER_8_385 ();
 sg13g2_fill_1 FILLER_8_387 ();
 sg13g2_fill_2 FILLER_8_421 ();
 sg13g2_fill_1 FILLER_8_423 ();
 sg13g2_fill_2 FILLER_9_0 ();
 sg13g2_fill_2 FILLER_9_36 ();
 sg13g2_fill_2 FILLER_9_65 ();
 sg13g2_fill_2 FILLER_9_112 ();
 sg13g2_fill_1 FILLER_9_158 ();
 sg13g2_fill_2 FILLER_9_197 ();
 sg13g2_fill_1 FILLER_9_199 ();
 sg13g2_decap_8 FILLER_9_225 ();
 sg13g2_fill_2 FILLER_9_287 ();
 sg13g2_fill_1 FILLER_9_340 ();
 sg13g2_fill_1 FILLER_9_389 ();
 sg13g2_fill_1 FILLER_9_423 ();
 sg13g2_fill_1 FILLER_10_0 ();
 sg13g2_fill_2 FILLER_10_39 ();
 sg13g2_fill_2 FILLER_10_48 ();
 sg13g2_fill_1 FILLER_10_50 ();
 sg13g2_fill_1 FILLER_10_85 ();
 sg13g2_fill_2 FILLER_10_153 ();
 sg13g2_fill_1 FILLER_10_155 ();
 sg13g2_fill_2 FILLER_10_194 ();
 sg13g2_fill_1 FILLER_10_200 ();
 sg13g2_fill_1 FILLER_10_247 ();
 sg13g2_fill_2 FILLER_10_273 ();
 sg13g2_fill_1 FILLER_10_315 ();
 sg13g2_fill_2 FILLER_10_343 ();
 sg13g2_fill_2 FILLER_10_393 ();
 sg13g2_fill_1 FILLER_10_412 ();
 sg13g2_fill_2 FILLER_10_421 ();
 sg13g2_fill_1 FILLER_10_423 ();
 sg13g2_fill_2 FILLER_11_0 ();
 sg13g2_fill_2 FILLER_11_29 ();
 sg13g2_fill_2 FILLER_11_87 ();
 sg13g2_fill_1 FILLER_11_89 ();
 sg13g2_fill_1 FILLER_11_175 ();
 sg13g2_fill_2 FILLER_11_227 ();
 sg13g2_fill_2 FILLER_11_327 ();
 sg13g2_fill_1 FILLER_11_329 ();
 sg13g2_fill_2 FILLER_11_421 ();
 sg13g2_fill_1 FILLER_11_423 ();
endmodule
