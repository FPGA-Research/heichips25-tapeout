magic
tech ihp-sg13g2
magscale 1 2
timestamp 1753461245
<< metal1 >>
rect 1152 9848 20452 9872
rect 1152 9808 4928 9848
rect 4968 9808 5010 9848
rect 5050 9808 5092 9848
rect 5132 9808 5174 9848
rect 5214 9808 5256 9848
rect 5296 9808 20048 9848
rect 20088 9808 20130 9848
rect 20170 9808 20212 9848
rect 20252 9808 20294 9848
rect 20334 9808 20376 9848
rect 20416 9808 20452 9848
rect 1152 9784 20452 9808
rect 1152 9092 20352 9116
rect 1152 9052 3688 9092
rect 3728 9052 3770 9092
rect 3810 9052 3852 9092
rect 3892 9052 3934 9092
rect 3974 9052 4016 9092
rect 4056 9052 18808 9092
rect 18848 9052 18890 9092
rect 18930 9052 18972 9092
rect 19012 9052 19054 9092
rect 19094 9052 19136 9092
rect 19176 9052 20352 9092
rect 1152 9028 20352 9052
rect 8811 8924 8853 8933
rect 8811 8884 8812 8924
rect 8852 8884 8853 8924
rect 8811 8875 8853 8884
rect 3435 8840 3477 8849
rect 3435 8800 3436 8840
rect 3476 8800 3477 8840
rect 3435 8791 3477 8800
rect 3819 8840 3861 8849
rect 3819 8800 3820 8840
rect 3860 8800 3861 8840
rect 3819 8791 3861 8800
rect 4779 8840 4821 8849
rect 4779 8800 4780 8840
rect 4820 8800 4821 8840
rect 4779 8791 4821 8800
rect 5739 8840 5781 8849
rect 5739 8800 5740 8840
rect 5780 8800 5781 8840
rect 5739 8791 5781 8800
rect 6603 8840 6645 8849
rect 6603 8800 6604 8840
rect 6644 8800 6645 8840
rect 6603 8791 6645 8800
rect 7851 8840 7893 8849
rect 7851 8800 7852 8840
rect 7892 8800 7893 8840
rect 7851 8791 7893 8800
rect 9387 8840 9429 8849
rect 9387 8800 9388 8840
rect 9428 8800 9429 8840
rect 9387 8791 9429 8800
rect 10443 8840 10485 8849
rect 10443 8800 10444 8840
rect 10484 8800 10485 8840
rect 10443 8791 10485 8800
rect 11403 8840 11445 8849
rect 11403 8800 11404 8840
rect 11444 8800 11445 8840
rect 11403 8791 11445 8800
rect 11595 8840 11637 8849
rect 11595 8800 11596 8840
rect 11636 8800 11637 8840
rect 11595 8791 11637 8800
rect 11979 8840 12021 8849
rect 11979 8800 11980 8840
rect 12020 8800 12021 8840
rect 11979 8791 12021 8800
rect 13035 8840 13077 8849
rect 13035 8800 13036 8840
rect 13076 8800 13077 8840
rect 13035 8791 13077 8800
rect 14091 8840 14133 8849
rect 14091 8800 14092 8840
rect 14132 8800 14133 8840
rect 14091 8791 14133 8800
rect 15435 8840 15477 8849
rect 15435 8800 15436 8840
rect 15476 8800 15477 8840
rect 15435 8791 15477 8800
rect 16107 8840 16149 8849
rect 16107 8800 16108 8840
rect 16148 8800 16149 8840
rect 16107 8791 16149 8800
rect 16491 8840 16533 8849
rect 16491 8800 16492 8840
rect 16532 8800 16533 8840
rect 16491 8791 16533 8800
rect 17067 8840 17109 8849
rect 17067 8800 17068 8840
rect 17108 8800 17109 8840
rect 17067 8791 17109 8800
rect 17835 8840 17877 8849
rect 17835 8800 17836 8840
rect 17876 8800 17877 8840
rect 17835 8791 17877 8800
rect 18411 8840 18453 8849
rect 18411 8800 18412 8840
rect 18452 8800 18453 8840
rect 18411 8791 18453 8800
rect 19563 8840 19605 8849
rect 19563 8800 19564 8840
rect 19604 8800 19605 8840
rect 19563 8791 19605 8800
rect 19755 8840 19797 8849
rect 19755 8800 19756 8840
rect 19796 8800 19797 8840
rect 19755 8791 19797 8800
rect 1507 8756 1565 8757
rect 1507 8716 1516 8756
rect 1556 8716 1565 8756
rect 1507 8715 1565 8716
rect 1891 8756 1949 8757
rect 1891 8716 1900 8756
rect 1940 8716 1949 8756
rect 1891 8715 1949 8716
rect 2275 8756 2333 8757
rect 2275 8716 2284 8756
rect 2324 8716 2333 8756
rect 2275 8715 2333 8716
rect 3619 8756 3677 8757
rect 3619 8716 3628 8756
rect 3668 8716 3677 8756
rect 3619 8715 3677 8716
rect 4003 8756 4061 8757
rect 4003 8716 4012 8756
rect 4052 8716 4061 8756
rect 4003 8715 4061 8716
rect 4963 8756 5021 8757
rect 4963 8716 4972 8756
rect 5012 8716 5021 8756
rect 4963 8715 5021 8716
rect 5923 8756 5981 8757
rect 5923 8716 5932 8756
rect 5972 8716 5981 8756
rect 5923 8715 5981 8716
rect 6787 8756 6845 8757
rect 6787 8716 6796 8756
rect 6836 8716 6845 8756
rect 6787 8715 6845 8716
rect 8035 8756 8093 8757
rect 8035 8716 8044 8756
rect 8084 8716 8093 8756
rect 8035 8715 8093 8716
rect 8995 8756 9053 8757
rect 8995 8716 9004 8756
rect 9044 8716 9053 8756
rect 8995 8715 9053 8716
rect 9571 8756 9629 8757
rect 9571 8716 9580 8756
rect 9620 8716 9629 8756
rect 9571 8715 9629 8716
rect 10627 8756 10685 8757
rect 10627 8716 10636 8756
rect 10676 8716 10685 8756
rect 10627 8715 10685 8716
rect 11203 8756 11261 8757
rect 11203 8716 11212 8756
rect 11252 8716 11261 8756
rect 11203 8715 11261 8716
rect 11779 8756 11837 8757
rect 11779 8716 11788 8756
rect 11828 8716 11837 8756
rect 11779 8715 11837 8716
rect 12163 8756 12221 8757
rect 12163 8716 12172 8756
rect 12212 8716 12221 8756
rect 12163 8715 12221 8716
rect 13219 8756 13277 8757
rect 13219 8716 13228 8756
rect 13268 8716 13277 8756
rect 13219 8715 13277 8716
rect 14275 8756 14333 8757
rect 14275 8716 14284 8756
rect 14324 8716 14333 8756
rect 14275 8715 14333 8716
rect 15619 8756 15677 8757
rect 15619 8716 15628 8756
rect 15668 8716 15677 8756
rect 15619 8715 15677 8716
rect 16291 8756 16349 8757
rect 16291 8716 16300 8756
rect 16340 8716 16349 8756
rect 16291 8715 16349 8716
rect 16675 8756 16733 8757
rect 16675 8716 16684 8756
rect 16724 8716 16733 8756
rect 16675 8715 16733 8716
rect 16867 8756 16925 8757
rect 16867 8716 16876 8756
rect 16916 8716 16925 8756
rect 16867 8715 16925 8716
rect 17635 8756 17693 8757
rect 17635 8716 17644 8756
rect 17684 8716 17693 8756
rect 17635 8715 17693 8716
rect 18211 8756 18269 8757
rect 18211 8716 18220 8756
rect 18260 8716 18269 8756
rect 18211 8715 18269 8716
rect 18979 8756 19037 8757
rect 18979 8716 18988 8756
rect 19028 8716 19037 8756
rect 18979 8715 19037 8716
rect 19363 8756 19421 8757
rect 19363 8716 19372 8756
rect 19412 8716 19421 8756
rect 19363 8715 19421 8716
rect 19939 8756 19997 8757
rect 19939 8716 19948 8756
rect 19988 8716 19997 8756
rect 19939 8715 19997 8716
rect 1707 8504 1749 8513
rect 1707 8464 1708 8504
rect 1748 8464 1749 8504
rect 1707 8455 1749 8464
rect 2091 8504 2133 8513
rect 2091 8464 2092 8504
rect 2132 8464 2133 8504
rect 2091 8455 2133 8464
rect 2475 8504 2517 8513
rect 2475 8464 2476 8504
rect 2516 8464 2517 8504
rect 2475 8455 2517 8464
rect 19179 8504 19221 8513
rect 19179 8464 19180 8504
rect 19220 8464 19221 8504
rect 19179 8455 19221 8464
rect 1152 8336 20452 8360
rect 1152 8296 4928 8336
rect 4968 8296 5010 8336
rect 5050 8296 5092 8336
rect 5132 8296 5174 8336
rect 5214 8296 5256 8336
rect 5296 8296 20048 8336
rect 20088 8296 20130 8336
rect 20170 8296 20212 8336
rect 20252 8296 20294 8336
rect 20334 8296 20376 8336
rect 20416 8296 20452 8336
rect 1152 8272 20452 8296
rect 2179 7916 2237 7917
rect 2179 7876 2188 7916
rect 2228 7876 2237 7916
rect 2179 7875 2237 7876
rect 13603 7916 13661 7917
rect 13603 7876 13612 7916
rect 13652 7876 13661 7916
rect 13603 7875 13661 7876
rect 13803 7832 13845 7841
rect 13803 7792 13804 7832
rect 13844 7792 13845 7832
rect 13803 7783 13845 7792
rect 2379 7748 2421 7757
rect 2379 7708 2380 7748
rect 2420 7708 2421 7748
rect 2379 7699 2421 7708
rect 1152 7580 20352 7604
rect 1152 7540 3688 7580
rect 3728 7540 3770 7580
rect 3810 7540 3852 7580
rect 3892 7540 3934 7580
rect 3974 7540 4016 7580
rect 4056 7540 18808 7580
rect 18848 7540 18890 7580
rect 18930 7540 18972 7580
rect 19012 7540 19054 7580
rect 19094 7540 19136 7580
rect 19176 7540 20352 7580
rect 1152 7516 20352 7540
rect 19267 7244 19325 7245
rect 19267 7204 19276 7244
rect 19316 7204 19325 7244
rect 19267 7203 19325 7204
rect 19467 6992 19509 7001
rect 19467 6952 19468 6992
rect 19508 6952 19509 6992
rect 19467 6943 19509 6952
rect 1152 6824 20452 6848
rect 1152 6784 4928 6824
rect 4968 6784 5010 6824
rect 5050 6784 5092 6824
rect 5132 6784 5174 6824
rect 5214 6784 5256 6824
rect 5296 6784 20048 6824
rect 20088 6784 20130 6824
rect 20170 6784 20212 6824
rect 20252 6784 20294 6824
rect 20334 6784 20376 6824
rect 20416 6784 20452 6824
rect 1152 6760 20452 6784
rect 2379 6656 2421 6665
rect 2379 6616 2380 6656
rect 2420 6616 2421 6656
rect 2379 6607 2421 6616
rect 2763 6656 2805 6665
rect 2763 6616 2764 6656
rect 2804 6616 2805 6656
rect 2763 6607 2805 6616
rect 18123 6656 18165 6665
rect 18123 6616 18124 6656
rect 18164 6616 18165 6656
rect 18123 6607 18165 6616
rect 19851 6656 19893 6665
rect 19851 6616 19852 6656
rect 19892 6616 19893 6656
rect 19851 6607 19893 6616
rect 1795 6404 1853 6405
rect 1795 6364 1804 6404
rect 1844 6364 1853 6404
rect 1795 6363 1853 6364
rect 2179 6404 2237 6405
rect 2179 6364 2188 6404
rect 2228 6364 2237 6404
rect 2179 6363 2237 6364
rect 2563 6404 2621 6405
rect 2563 6364 2572 6404
rect 2612 6364 2621 6404
rect 2563 6363 2621 6364
rect 17923 6404 17981 6405
rect 17923 6364 17932 6404
rect 17972 6364 17981 6404
rect 17923 6363 17981 6364
rect 19267 6404 19325 6405
rect 19267 6364 19276 6404
rect 19316 6364 19325 6404
rect 19267 6363 19325 6364
rect 19651 6404 19709 6405
rect 19651 6364 19660 6404
rect 19700 6364 19709 6404
rect 19651 6363 19709 6364
rect 1995 6236 2037 6245
rect 1995 6196 1996 6236
rect 2036 6196 2037 6236
rect 1995 6187 2037 6196
rect 19467 6236 19509 6245
rect 19467 6196 19468 6236
rect 19508 6196 19509 6236
rect 19467 6187 19509 6196
rect 1152 6068 20352 6092
rect 1152 6028 3688 6068
rect 3728 6028 3770 6068
rect 3810 6028 3852 6068
rect 3892 6028 3934 6068
rect 3974 6028 4016 6068
rect 4056 6028 18808 6068
rect 18848 6028 18890 6068
rect 18930 6028 18972 6068
rect 19012 6028 19054 6068
rect 19094 6028 19136 6068
rect 19176 6028 20352 6068
rect 1152 6004 20352 6028
rect 1891 5732 1949 5733
rect 1891 5692 1900 5732
rect 1940 5692 1949 5732
rect 1891 5691 1949 5692
rect 19171 5732 19229 5733
rect 19171 5692 19180 5732
rect 19220 5692 19229 5732
rect 19171 5691 19229 5692
rect 2091 5480 2133 5489
rect 2091 5440 2092 5480
rect 2132 5440 2133 5480
rect 2091 5431 2133 5440
rect 19371 5480 19413 5489
rect 19371 5440 19372 5480
rect 19412 5440 19413 5480
rect 19371 5431 19413 5440
rect 1152 5312 20452 5336
rect 1152 5272 4928 5312
rect 4968 5272 5010 5312
rect 5050 5272 5092 5312
rect 5132 5272 5174 5312
rect 5214 5272 5256 5312
rect 5296 5272 20048 5312
rect 20088 5272 20130 5312
rect 20170 5272 20212 5312
rect 20252 5272 20294 5312
rect 20334 5272 20376 5312
rect 20416 5272 20452 5312
rect 1152 5248 20452 5272
rect 1891 4892 1949 4893
rect 1891 4852 1900 4892
rect 1940 4852 1949 4892
rect 1891 4851 1949 4852
rect 16675 4892 16733 4893
rect 16675 4852 16684 4892
rect 16724 4852 16733 4892
rect 16675 4851 16733 4852
rect 17251 4892 17309 4893
rect 17251 4852 17260 4892
rect 17300 4852 17309 4892
rect 17251 4851 17309 4852
rect 2091 4724 2133 4733
rect 2091 4684 2092 4724
rect 2132 4684 2133 4724
rect 2091 4675 2133 4684
rect 16875 4724 16917 4733
rect 16875 4684 16876 4724
rect 16916 4684 16917 4724
rect 16875 4675 16917 4684
rect 17451 4724 17493 4733
rect 17451 4684 17452 4724
rect 17492 4684 17493 4724
rect 17451 4675 17493 4684
rect 1152 4556 20352 4580
rect 1152 4516 3688 4556
rect 3728 4516 3770 4556
rect 3810 4516 3852 4556
rect 3892 4516 3934 4556
rect 3974 4516 4016 4556
rect 4056 4516 18808 4556
rect 18848 4516 18890 4556
rect 18930 4516 18972 4556
rect 19012 4516 19054 4556
rect 19094 4516 19136 4556
rect 19176 4516 20352 4556
rect 1152 4492 20352 4516
rect 1899 4388 1941 4397
rect 1899 4348 1900 4388
rect 1940 4348 1941 4388
rect 1899 4339 1941 4348
rect 19371 4388 19413 4397
rect 19371 4348 19372 4388
rect 19412 4348 19413 4388
rect 19371 4339 19413 4348
rect 2083 4220 2141 4221
rect 2083 4180 2092 4220
rect 2132 4180 2141 4220
rect 2083 4179 2141 4180
rect 18787 4220 18845 4221
rect 18787 4180 18796 4220
rect 18836 4180 18845 4220
rect 18787 4179 18845 4180
rect 19171 4220 19229 4221
rect 19171 4180 19180 4220
rect 19220 4180 19229 4220
rect 19171 4179 19229 4180
rect 19555 4220 19613 4221
rect 19555 4180 19564 4220
rect 19604 4180 19613 4220
rect 19555 4179 19613 4180
rect 18987 3968 19029 3977
rect 18987 3928 18988 3968
rect 19028 3928 19029 3968
rect 18987 3919 19029 3928
rect 19755 3968 19797 3977
rect 19755 3928 19756 3968
rect 19796 3928 19797 3968
rect 19755 3919 19797 3928
rect 1152 3800 20452 3824
rect 1152 3760 4928 3800
rect 4968 3760 5010 3800
rect 5050 3760 5092 3800
rect 5132 3760 5174 3800
rect 5214 3760 5256 3800
rect 5296 3760 20048 3800
rect 20088 3760 20130 3800
rect 20170 3760 20212 3800
rect 20252 3760 20294 3800
rect 20334 3760 20376 3800
rect 20416 3760 20452 3800
rect 1152 3736 20452 3760
rect 1891 3380 1949 3381
rect 1891 3340 1900 3380
rect 1940 3340 1949 3380
rect 1891 3339 1949 3340
rect 19267 3380 19325 3381
rect 19267 3340 19276 3380
rect 19316 3340 19325 3380
rect 19267 3339 19325 3340
rect 2091 3212 2133 3221
rect 2091 3172 2092 3212
rect 2132 3172 2133 3212
rect 2091 3163 2133 3172
rect 19467 3212 19509 3221
rect 19467 3172 19468 3212
rect 19508 3172 19509 3212
rect 19467 3163 19509 3172
rect 1152 3044 20352 3068
rect 1152 3004 3688 3044
rect 3728 3004 3770 3044
rect 3810 3004 3852 3044
rect 3892 3004 3934 3044
rect 3974 3004 4016 3044
rect 4056 3004 18808 3044
rect 18848 3004 18890 3044
rect 18930 3004 18972 3044
rect 19012 3004 19054 3044
rect 19094 3004 19136 3044
rect 19176 3004 20352 3044
rect 1152 2980 20352 3004
rect 2955 2876 2997 2885
rect 2955 2836 2956 2876
rect 2996 2836 2997 2876
rect 2955 2827 2997 2836
rect 3723 2876 3765 2885
rect 3723 2836 3724 2876
rect 3764 2836 3765 2876
rect 3723 2827 3765 2836
rect 6891 2792 6933 2801
rect 6891 2752 6892 2792
rect 6932 2752 6933 2792
rect 6891 2743 6933 2752
rect 1891 2708 1949 2709
rect 1891 2668 1900 2708
rect 1940 2668 1949 2708
rect 1891 2667 1949 2668
rect 2755 2708 2813 2709
rect 2755 2668 2764 2708
rect 2804 2668 2813 2708
rect 2755 2667 2813 2668
rect 3523 2708 3581 2709
rect 3523 2668 3532 2708
rect 3572 2668 3581 2708
rect 3523 2667 3581 2668
rect 6691 2708 6749 2709
rect 6691 2668 6700 2708
rect 6740 2668 6749 2708
rect 6691 2667 6749 2668
rect 8707 2708 8765 2709
rect 8707 2668 8716 2708
rect 8756 2668 8765 2708
rect 8707 2667 8765 2668
rect 9667 2708 9725 2709
rect 9667 2668 9676 2708
rect 9716 2668 9725 2708
rect 9667 2667 9725 2668
rect 15139 2708 15197 2709
rect 15139 2668 15148 2708
rect 15188 2668 15197 2708
rect 15139 2667 15197 2668
rect 15523 2708 15581 2709
rect 15523 2668 15532 2708
rect 15572 2668 15581 2708
rect 15523 2667 15581 2668
rect 16099 2708 16157 2709
rect 16099 2668 16108 2708
rect 16148 2668 16157 2708
rect 16099 2667 16157 2668
rect 17347 2708 17405 2709
rect 17347 2668 17356 2708
rect 17396 2668 17405 2708
rect 17347 2667 17405 2668
rect 2091 2456 2133 2465
rect 2091 2416 2092 2456
rect 2132 2416 2133 2456
rect 2091 2407 2133 2416
rect 8907 2456 8949 2465
rect 8907 2416 8908 2456
rect 8948 2416 8949 2456
rect 8907 2407 8949 2416
rect 9867 2456 9909 2465
rect 9867 2416 9868 2456
rect 9908 2416 9909 2456
rect 9867 2407 9909 2416
rect 14955 2456 14997 2465
rect 14955 2416 14956 2456
rect 14996 2416 14997 2456
rect 14955 2407 14997 2416
rect 15339 2456 15381 2465
rect 15339 2416 15340 2456
rect 15380 2416 15381 2456
rect 15339 2407 15381 2416
rect 15915 2456 15957 2465
rect 15915 2416 15916 2456
rect 15956 2416 15957 2456
rect 15915 2407 15957 2416
rect 17547 2456 17589 2465
rect 17547 2416 17548 2456
rect 17588 2416 17589 2456
rect 17547 2407 17589 2416
rect 1152 2288 20452 2312
rect 1152 2248 4928 2288
rect 4968 2248 5010 2288
rect 5050 2248 5092 2288
rect 5132 2248 5174 2288
rect 5214 2248 5256 2288
rect 5296 2248 20048 2288
rect 20088 2248 20130 2288
rect 20170 2248 20212 2288
rect 20252 2248 20294 2288
rect 20334 2248 20376 2288
rect 20416 2248 20452 2288
rect 1152 2224 20452 2248
rect 2091 2120 2133 2129
rect 2091 2080 2092 2120
rect 2132 2080 2133 2120
rect 2091 2071 2133 2080
rect 2475 2120 2517 2129
rect 2475 2080 2476 2120
rect 2516 2080 2517 2120
rect 2475 2071 2517 2080
rect 2859 2120 2901 2129
rect 2859 2080 2860 2120
rect 2900 2080 2901 2120
rect 2859 2071 2901 2080
rect 5355 2120 5397 2129
rect 5355 2080 5356 2120
rect 5396 2080 5397 2120
rect 5355 2071 5397 2080
rect 19563 2120 19605 2129
rect 19563 2080 19564 2120
rect 19604 2080 19605 2120
rect 19563 2071 19605 2080
rect 19947 2120 19989 2129
rect 19947 2080 19948 2120
rect 19988 2080 19989 2120
rect 19947 2071 19989 2080
rect 1891 1868 1949 1869
rect 1891 1828 1900 1868
rect 1940 1828 1949 1868
rect 1891 1827 1949 1828
rect 2275 1868 2333 1869
rect 2275 1828 2284 1868
rect 2324 1828 2333 1868
rect 2275 1827 2333 1828
rect 2659 1868 2717 1869
rect 2659 1828 2668 1868
rect 2708 1828 2717 1868
rect 2659 1827 2717 1828
rect 3715 1868 3773 1869
rect 3715 1828 3724 1868
rect 3764 1828 3773 1868
rect 3715 1827 3773 1828
rect 4099 1868 4157 1869
rect 4099 1828 4108 1868
rect 4148 1828 4157 1868
rect 4099 1827 4157 1828
rect 4483 1868 4541 1869
rect 4483 1828 4492 1868
rect 4532 1828 4541 1868
rect 4483 1827 4541 1828
rect 5155 1868 5213 1869
rect 5155 1828 5164 1868
rect 5204 1828 5213 1868
rect 5155 1827 5213 1828
rect 5635 1868 5693 1869
rect 5635 1828 5644 1868
rect 5684 1828 5693 1868
rect 5635 1827 5693 1828
rect 6115 1868 6173 1869
rect 6115 1828 6124 1868
rect 6164 1828 6173 1868
rect 6115 1827 6173 1828
rect 6883 1868 6941 1869
rect 6883 1828 6892 1868
rect 6932 1828 6941 1868
rect 6883 1827 6941 1828
rect 7267 1868 7325 1869
rect 7267 1828 7276 1868
rect 7316 1828 7325 1868
rect 7267 1827 7325 1828
rect 7651 1868 7709 1869
rect 7651 1828 7660 1868
rect 7700 1828 7709 1868
rect 7651 1827 7709 1828
rect 8035 1868 8093 1869
rect 8035 1828 8044 1868
rect 8084 1828 8093 1868
rect 8035 1827 8093 1828
rect 8419 1868 8477 1869
rect 8419 1828 8428 1868
rect 8468 1828 8477 1868
rect 8419 1827 8477 1828
rect 9955 1868 10013 1869
rect 9955 1828 9964 1868
rect 10004 1828 10013 1868
rect 9955 1827 10013 1828
rect 10339 1868 10397 1869
rect 10339 1828 10348 1868
rect 10388 1828 10397 1868
rect 10339 1827 10397 1828
rect 10819 1868 10877 1869
rect 10819 1828 10828 1868
rect 10868 1828 10877 1868
rect 10819 1827 10877 1828
rect 11203 1868 11261 1869
rect 11203 1828 11212 1868
rect 11252 1828 11261 1868
rect 11203 1827 11261 1828
rect 11587 1868 11645 1869
rect 11587 1828 11596 1868
rect 11636 1828 11645 1868
rect 11587 1827 11645 1828
rect 11971 1868 12029 1869
rect 11971 1828 11980 1868
rect 12020 1828 12029 1868
rect 11971 1827 12029 1828
rect 12835 1868 12893 1869
rect 12835 1828 12844 1868
rect 12884 1828 12893 1868
rect 12835 1827 12893 1828
rect 13219 1868 13277 1869
rect 13219 1828 13228 1868
rect 13268 1828 13277 1868
rect 13219 1827 13277 1828
rect 13603 1868 13661 1869
rect 13603 1828 13612 1868
rect 13652 1828 13661 1868
rect 13603 1827 13661 1828
rect 13987 1868 14045 1869
rect 13987 1828 13996 1868
rect 14036 1828 14045 1868
rect 13987 1827 14045 1828
rect 14563 1868 14621 1869
rect 14563 1828 14572 1868
rect 14612 1828 14621 1868
rect 14563 1827 14621 1828
rect 16099 1868 16157 1869
rect 16099 1828 16108 1868
rect 16148 1828 16157 1868
rect 16099 1827 16157 1828
rect 16963 1868 17021 1869
rect 16963 1828 16972 1868
rect 17012 1828 17021 1868
rect 16963 1827 17021 1828
rect 17347 1868 17405 1869
rect 17347 1828 17356 1868
rect 17396 1828 17405 1868
rect 17347 1827 17405 1828
rect 17731 1868 17789 1869
rect 17731 1828 17740 1868
rect 17780 1828 17789 1868
rect 17731 1827 17789 1828
rect 18979 1868 19037 1869
rect 18979 1828 18988 1868
rect 19028 1828 19037 1868
rect 18979 1827 19037 1828
rect 19363 1868 19421 1869
rect 19363 1828 19372 1868
rect 19412 1828 19421 1868
rect 19363 1827 19421 1828
rect 19747 1868 19805 1869
rect 19747 1828 19756 1868
rect 19796 1828 19805 1868
rect 19747 1827 19805 1828
rect 19179 1784 19221 1793
rect 19179 1744 19180 1784
rect 19220 1744 19221 1784
rect 19179 1735 19221 1744
rect 3915 1700 3957 1709
rect 3915 1660 3916 1700
rect 3956 1660 3957 1700
rect 3915 1651 3957 1660
rect 4299 1700 4341 1709
rect 4299 1660 4300 1700
rect 4340 1660 4341 1700
rect 4299 1651 4341 1660
rect 4683 1700 4725 1709
rect 4683 1660 4684 1700
rect 4724 1660 4725 1700
rect 4683 1651 4725 1660
rect 5835 1700 5877 1709
rect 5835 1660 5836 1700
rect 5876 1660 5877 1700
rect 5835 1651 5877 1660
rect 6315 1700 6357 1709
rect 6315 1660 6316 1700
rect 6356 1660 6357 1700
rect 6315 1651 6357 1660
rect 7083 1700 7125 1709
rect 7083 1660 7084 1700
rect 7124 1660 7125 1700
rect 7083 1651 7125 1660
rect 7467 1700 7509 1709
rect 7467 1660 7468 1700
rect 7508 1660 7509 1700
rect 7467 1651 7509 1660
rect 7851 1700 7893 1709
rect 7851 1660 7852 1700
rect 7892 1660 7893 1700
rect 7851 1651 7893 1660
rect 8235 1700 8277 1709
rect 8235 1660 8236 1700
rect 8276 1660 8277 1700
rect 8235 1651 8277 1660
rect 8619 1700 8661 1709
rect 8619 1660 8620 1700
rect 8660 1660 8661 1700
rect 8619 1651 8661 1660
rect 10155 1700 10197 1709
rect 10155 1660 10156 1700
rect 10196 1660 10197 1700
rect 10155 1651 10197 1660
rect 10539 1700 10581 1709
rect 10539 1660 10540 1700
rect 10580 1660 10581 1700
rect 10539 1651 10581 1660
rect 11019 1700 11061 1709
rect 11019 1660 11020 1700
rect 11060 1660 11061 1700
rect 11019 1651 11061 1660
rect 11403 1700 11445 1709
rect 11403 1660 11404 1700
rect 11444 1660 11445 1700
rect 11403 1651 11445 1660
rect 11787 1700 11829 1709
rect 11787 1660 11788 1700
rect 11828 1660 11829 1700
rect 11787 1651 11829 1660
rect 12171 1700 12213 1709
rect 12171 1660 12172 1700
rect 12212 1660 12213 1700
rect 12171 1651 12213 1660
rect 13035 1700 13077 1709
rect 13035 1660 13036 1700
rect 13076 1660 13077 1700
rect 13035 1651 13077 1660
rect 13419 1700 13461 1709
rect 13419 1660 13420 1700
rect 13460 1660 13461 1700
rect 13419 1651 13461 1660
rect 13803 1700 13845 1709
rect 13803 1660 13804 1700
rect 13844 1660 13845 1700
rect 13803 1651 13845 1660
rect 14187 1700 14229 1709
rect 14187 1660 14188 1700
rect 14228 1660 14229 1700
rect 14187 1651 14229 1660
rect 14763 1700 14805 1709
rect 14763 1660 14764 1700
rect 14804 1660 14805 1700
rect 14763 1651 14805 1660
rect 15915 1700 15957 1709
rect 15915 1660 15916 1700
rect 15956 1660 15957 1700
rect 15915 1651 15957 1660
rect 17163 1700 17205 1709
rect 17163 1660 17164 1700
rect 17204 1660 17205 1700
rect 17163 1651 17205 1660
rect 17547 1700 17589 1709
rect 17547 1660 17548 1700
rect 17588 1660 17589 1700
rect 17547 1651 17589 1660
rect 17931 1700 17973 1709
rect 17931 1660 17932 1700
rect 17972 1660 17973 1700
rect 17931 1651 17973 1660
rect 1152 1532 20352 1556
rect 1152 1492 3688 1532
rect 3728 1492 3770 1532
rect 3810 1492 3852 1532
rect 3892 1492 3934 1532
rect 3974 1492 4016 1532
rect 4056 1492 18808 1532
rect 18848 1492 18890 1532
rect 18930 1492 18972 1532
rect 19012 1492 19054 1532
rect 19094 1492 19136 1532
rect 19176 1492 20352 1532
rect 1152 1468 20352 1492
rect 17347 1196 17405 1197
rect 17347 1156 17356 1196
rect 17396 1156 17405 1196
rect 17347 1155 17405 1156
rect 17547 944 17589 953
rect 17547 904 17548 944
rect 17588 904 17589 944
rect 17547 895 17589 904
rect 1152 776 20452 800
rect 1152 736 4928 776
rect 4968 736 5010 776
rect 5050 736 5092 776
rect 5132 736 5174 776
rect 5214 736 5256 776
rect 5296 736 20048 776
rect 20088 736 20130 776
rect 20170 736 20212 776
rect 20252 736 20294 776
rect 20334 736 20376 776
rect 20416 736 20452 776
rect 1152 712 20452 736
<< via1 >>
rect 4928 9808 4968 9848
rect 5010 9808 5050 9848
rect 5092 9808 5132 9848
rect 5174 9808 5214 9848
rect 5256 9808 5296 9848
rect 20048 9808 20088 9848
rect 20130 9808 20170 9848
rect 20212 9808 20252 9848
rect 20294 9808 20334 9848
rect 20376 9808 20416 9848
rect 3688 9052 3728 9092
rect 3770 9052 3810 9092
rect 3852 9052 3892 9092
rect 3934 9052 3974 9092
rect 4016 9052 4056 9092
rect 18808 9052 18848 9092
rect 18890 9052 18930 9092
rect 18972 9052 19012 9092
rect 19054 9052 19094 9092
rect 19136 9052 19176 9092
rect 8812 8884 8852 8924
rect 3436 8800 3476 8840
rect 3820 8800 3860 8840
rect 4780 8800 4820 8840
rect 5740 8800 5780 8840
rect 6604 8800 6644 8840
rect 7852 8800 7892 8840
rect 9388 8800 9428 8840
rect 10444 8800 10484 8840
rect 11404 8800 11444 8840
rect 11596 8800 11636 8840
rect 11980 8800 12020 8840
rect 13036 8800 13076 8840
rect 14092 8800 14132 8840
rect 15436 8800 15476 8840
rect 16108 8800 16148 8840
rect 16492 8800 16532 8840
rect 17068 8800 17108 8840
rect 17836 8800 17876 8840
rect 18412 8800 18452 8840
rect 19564 8800 19604 8840
rect 19756 8800 19796 8840
rect 1516 8716 1556 8756
rect 1900 8716 1940 8756
rect 2284 8716 2324 8756
rect 3628 8716 3668 8756
rect 4012 8716 4052 8756
rect 4972 8716 5012 8756
rect 5932 8716 5972 8756
rect 6796 8716 6836 8756
rect 8044 8716 8084 8756
rect 9004 8716 9044 8756
rect 9580 8716 9620 8756
rect 10636 8716 10676 8756
rect 11212 8716 11252 8756
rect 11788 8716 11828 8756
rect 12172 8716 12212 8756
rect 13228 8716 13268 8756
rect 14284 8716 14324 8756
rect 15628 8716 15668 8756
rect 16300 8716 16340 8756
rect 16684 8716 16724 8756
rect 16876 8716 16916 8756
rect 17644 8716 17684 8756
rect 18220 8716 18260 8756
rect 18988 8716 19028 8756
rect 19372 8716 19412 8756
rect 19948 8716 19988 8756
rect 1708 8464 1748 8504
rect 2092 8464 2132 8504
rect 2476 8464 2516 8504
rect 19180 8464 19220 8504
rect 4928 8296 4968 8336
rect 5010 8296 5050 8336
rect 5092 8296 5132 8336
rect 5174 8296 5214 8336
rect 5256 8296 5296 8336
rect 20048 8296 20088 8336
rect 20130 8296 20170 8336
rect 20212 8296 20252 8336
rect 20294 8296 20334 8336
rect 20376 8296 20416 8336
rect 2188 7876 2228 7916
rect 13612 7876 13652 7916
rect 13804 7792 13844 7832
rect 2380 7708 2420 7748
rect 3688 7540 3728 7580
rect 3770 7540 3810 7580
rect 3852 7540 3892 7580
rect 3934 7540 3974 7580
rect 4016 7540 4056 7580
rect 18808 7540 18848 7580
rect 18890 7540 18930 7580
rect 18972 7540 19012 7580
rect 19054 7540 19094 7580
rect 19136 7540 19176 7580
rect 19276 7204 19316 7244
rect 19468 6952 19508 6992
rect 4928 6784 4968 6824
rect 5010 6784 5050 6824
rect 5092 6784 5132 6824
rect 5174 6784 5214 6824
rect 5256 6784 5296 6824
rect 20048 6784 20088 6824
rect 20130 6784 20170 6824
rect 20212 6784 20252 6824
rect 20294 6784 20334 6824
rect 20376 6784 20416 6824
rect 2380 6616 2420 6656
rect 2764 6616 2804 6656
rect 18124 6616 18164 6656
rect 19852 6616 19892 6656
rect 1804 6364 1844 6404
rect 2188 6364 2228 6404
rect 2572 6364 2612 6404
rect 17932 6364 17972 6404
rect 19276 6364 19316 6404
rect 19660 6364 19700 6404
rect 1996 6196 2036 6236
rect 19468 6196 19508 6236
rect 3688 6028 3728 6068
rect 3770 6028 3810 6068
rect 3852 6028 3892 6068
rect 3934 6028 3974 6068
rect 4016 6028 4056 6068
rect 18808 6028 18848 6068
rect 18890 6028 18930 6068
rect 18972 6028 19012 6068
rect 19054 6028 19094 6068
rect 19136 6028 19176 6068
rect 1900 5692 1940 5732
rect 19180 5692 19220 5732
rect 2092 5440 2132 5480
rect 19372 5440 19412 5480
rect 4928 5272 4968 5312
rect 5010 5272 5050 5312
rect 5092 5272 5132 5312
rect 5174 5272 5214 5312
rect 5256 5272 5296 5312
rect 20048 5272 20088 5312
rect 20130 5272 20170 5312
rect 20212 5272 20252 5312
rect 20294 5272 20334 5312
rect 20376 5272 20416 5312
rect 1900 4852 1940 4892
rect 16684 4852 16724 4892
rect 17260 4852 17300 4892
rect 2092 4684 2132 4724
rect 16876 4684 16916 4724
rect 17452 4684 17492 4724
rect 3688 4516 3728 4556
rect 3770 4516 3810 4556
rect 3852 4516 3892 4556
rect 3934 4516 3974 4556
rect 4016 4516 4056 4556
rect 18808 4516 18848 4556
rect 18890 4516 18930 4556
rect 18972 4516 19012 4556
rect 19054 4516 19094 4556
rect 19136 4516 19176 4556
rect 1900 4348 1940 4388
rect 19372 4348 19412 4388
rect 2092 4180 2132 4220
rect 18796 4180 18836 4220
rect 19180 4180 19220 4220
rect 19564 4180 19604 4220
rect 18988 3928 19028 3968
rect 19756 3928 19796 3968
rect 4928 3760 4968 3800
rect 5010 3760 5050 3800
rect 5092 3760 5132 3800
rect 5174 3760 5214 3800
rect 5256 3760 5296 3800
rect 20048 3760 20088 3800
rect 20130 3760 20170 3800
rect 20212 3760 20252 3800
rect 20294 3760 20334 3800
rect 20376 3760 20416 3800
rect 1900 3340 1940 3380
rect 19276 3340 19316 3380
rect 2092 3172 2132 3212
rect 19468 3172 19508 3212
rect 3688 3004 3728 3044
rect 3770 3004 3810 3044
rect 3852 3004 3892 3044
rect 3934 3004 3974 3044
rect 4016 3004 4056 3044
rect 18808 3004 18848 3044
rect 18890 3004 18930 3044
rect 18972 3004 19012 3044
rect 19054 3004 19094 3044
rect 19136 3004 19176 3044
rect 2956 2836 2996 2876
rect 3724 2836 3764 2876
rect 6892 2752 6932 2792
rect 1900 2668 1940 2708
rect 2764 2668 2804 2708
rect 3532 2668 3572 2708
rect 6700 2668 6740 2708
rect 8716 2668 8756 2708
rect 9676 2668 9716 2708
rect 15148 2668 15188 2708
rect 15532 2668 15572 2708
rect 16108 2668 16148 2708
rect 17356 2668 17396 2708
rect 2092 2416 2132 2456
rect 8908 2416 8948 2456
rect 9868 2416 9908 2456
rect 14956 2416 14996 2456
rect 15340 2416 15380 2456
rect 15916 2416 15956 2456
rect 17548 2416 17588 2456
rect 4928 2248 4968 2288
rect 5010 2248 5050 2288
rect 5092 2248 5132 2288
rect 5174 2248 5214 2288
rect 5256 2248 5296 2288
rect 20048 2248 20088 2288
rect 20130 2248 20170 2288
rect 20212 2248 20252 2288
rect 20294 2248 20334 2288
rect 20376 2248 20416 2288
rect 2092 2080 2132 2120
rect 2476 2080 2516 2120
rect 2860 2080 2900 2120
rect 5356 2080 5396 2120
rect 19564 2080 19604 2120
rect 19948 2080 19988 2120
rect 1900 1828 1940 1868
rect 2284 1828 2324 1868
rect 2668 1828 2708 1868
rect 3724 1828 3764 1868
rect 4108 1828 4148 1868
rect 4492 1828 4532 1868
rect 5164 1828 5204 1868
rect 5644 1828 5684 1868
rect 6124 1828 6164 1868
rect 6892 1828 6932 1868
rect 7276 1828 7316 1868
rect 7660 1828 7700 1868
rect 8044 1828 8084 1868
rect 8428 1828 8468 1868
rect 9964 1828 10004 1868
rect 10348 1828 10388 1868
rect 10828 1828 10868 1868
rect 11212 1828 11252 1868
rect 11596 1828 11636 1868
rect 11980 1828 12020 1868
rect 12844 1828 12884 1868
rect 13228 1828 13268 1868
rect 13612 1828 13652 1868
rect 13996 1828 14036 1868
rect 14572 1828 14612 1868
rect 16108 1828 16148 1868
rect 16972 1828 17012 1868
rect 17356 1828 17396 1868
rect 17740 1828 17780 1868
rect 18988 1828 19028 1868
rect 19372 1828 19412 1868
rect 19756 1828 19796 1868
rect 19180 1744 19220 1784
rect 3916 1660 3956 1700
rect 4300 1660 4340 1700
rect 4684 1660 4724 1700
rect 5836 1660 5876 1700
rect 6316 1660 6356 1700
rect 7084 1660 7124 1700
rect 7468 1660 7508 1700
rect 7852 1660 7892 1700
rect 8236 1660 8276 1700
rect 8620 1660 8660 1700
rect 10156 1660 10196 1700
rect 10540 1660 10580 1700
rect 11020 1660 11060 1700
rect 11404 1660 11444 1700
rect 11788 1660 11828 1700
rect 12172 1660 12212 1700
rect 13036 1660 13076 1700
rect 13420 1660 13460 1700
rect 13804 1660 13844 1700
rect 14188 1660 14228 1700
rect 14764 1660 14804 1700
rect 15916 1660 15956 1700
rect 17164 1660 17204 1700
rect 17548 1660 17588 1700
rect 17932 1660 17972 1700
rect 3688 1492 3728 1532
rect 3770 1492 3810 1532
rect 3852 1492 3892 1532
rect 3934 1492 3974 1532
rect 4016 1492 4056 1532
rect 18808 1492 18848 1532
rect 18890 1492 18930 1532
rect 18972 1492 19012 1532
rect 19054 1492 19094 1532
rect 19136 1492 19176 1532
rect 17356 1156 17396 1196
rect 17548 904 17588 944
rect 4928 736 4968 776
rect 5010 736 5050 776
rect 5092 736 5132 776
rect 5174 736 5214 776
rect 5256 736 5296 776
rect 20048 736 20088 776
rect 20130 736 20170 776
rect 20212 736 20252 776
rect 20294 736 20334 776
rect 20376 736 20416 776
<< metal2 >>
rect 1016 10672 1096 10752
rect 1976 10672 2056 10752
rect 2936 10672 3016 10752
rect 3896 10672 3976 10752
rect 4108 10692 4724 10732
rect 555 10520 597 10529
rect 555 10480 556 10520
rect 596 10480 597 10520
rect 555 10471 597 10480
rect 556 8009 596 10471
rect 555 8000 597 8009
rect 555 7960 556 8000
rect 596 7960 597 8000
rect 555 7951 597 7960
rect 1036 4397 1076 10672
rect 1515 9848 1557 9857
rect 1515 9808 1516 9848
rect 1556 9808 1557 9848
rect 1515 9799 1557 9808
rect 1516 8756 1556 9799
rect 1899 9512 1941 9521
rect 1899 9472 1900 9512
rect 1940 9472 1941 9512
rect 1899 9463 1941 9472
rect 1516 8707 1556 8716
rect 1900 8756 1940 9463
rect 1900 8707 1940 8716
rect 1996 8681 2036 10672
rect 2283 10184 2325 10193
rect 2283 10144 2284 10184
rect 2324 10144 2325 10184
rect 2283 10135 2325 10144
rect 2284 8756 2324 10135
rect 2956 8765 2996 10672
rect 3916 10604 3956 10672
rect 4108 10604 4148 10692
rect 3916 10564 4148 10604
rect 3688 9092 4056 9101
rect 3728 9052 3770 9092
rect 3810 9052 3852 9092
rect 3892 9052 3934 9092
rect 3974 9052 4016 9092
rect 3688 9043 4056 9052
rect 3436 8840 3476 8849
rect 2284 8707 2324 8716
rect 2955 8756 2997 8765
rect 2955 8716 2956 8756
rect 2996 8716 2997 8756
rect 2955 8707 2997 8716
rect 3436 8681 3476 8800
rect 3820 8840 3860 8851
rect 4684 8840 4724 10692
rect 4856 10672 4936 10752
rect 5816 10672 5896 10752
rect 6776 10672 6856 10752
rect 7736 10672 7816 10752
rect 8696 10672 8776 10752
rect 9656 10672 9736 10752
rect 10616 10672 10696 10752
rect 11576 10672 11656 10752
rect 11788 10692 12020 10732
rect 4876 10016 4916 10672
rect 5836 10604 5876 10672
rect 5836 10564 6068 10604
rect 4780 9976 4916 10016
rect 4780 9008 4820 9976
rect 4928 9848 5296 9857
rect 4968 9808 5010 9848
rect 5050 9808 5092 9848
rect 5132 9808 5174 9848
rect 5214 9808 5256 9848
rect 4928 9799 5296 9808
rect 4780 8968 4916 9008
rect 4780 8840 4820 8849
rect 4684 8800 4780 8840
rect 3820 8765 3860 8800
rect 4780 8791 4820 8800
rect 4876 8765 4916 8968
rect 5740 8840 5780 8851
rect 5740 8765 5780 8800
rect 6028 8765 6068 10564
rect 6796 8924 6836 10672
rect 7756 9689 7796 10672
rect 7755 9680 7797 9689
rect 7755 9640 7756 9680
rect 7796 9640 7797 9680
rect 7755 9631 7797 9640
rect 6796 8884 6932 8924
rect 6603 8840 6645 8849
rect 6603 8800 6604 8840
rect 6644 8800 6645 8840
rect 6603 8791 6645 8800
rect 3628 8756 3668 8765
rect 3532 8716 3628 8756
rect 1995 8672 2037 8681
rect 1995 8632 1996 8672
rect 2036 8632 2037 8672
rect 1995 8623 2037 8632
rect 3435 8672 3477 8681
rect 3435 8632 3436 8672
rect 3476 8632 3477 8672
rect 3435 8623 3477 8632
rect 1708 8504 1748 8513
rect 1708 8345 1748 8464
rect 2091 8504 2133 8513
rect 2091 8464 2092 8504
rect 2132 8464 2133 8504
rect 2091 8455 2133 8464
rect 2475 8504 2517 8513
rect 2475 8464 2476 8504
rect 2516 8464 2517 8504
rect 2475 8455 2517 8464
rect 2092 8370 2132 8455
rect 2476 8370 2516 8455
rect 1707 8336 1749 8345
rect 1707 8296 1708 8336
rect 1748 8296 1749 8336
rect 1707 8287 1749 8296
rect 2187 7916 2229 7925
rect 2187 7876 2188 7916
rect 2228 7876 2229 7916
rect 2187 7867 2229 7876
rect 2188 7782 2228 7867
rect 2379 7748 2421 7757
rect 2379 7708 2380 7748
rect 2420 7708 2421 7748
rect 2379 7699 2421 7708
rect 2380 7614 2420 7699
rect 2571 7160 2613 7169
rect 2571 7120 2572 7160
rect 2612 7120 2613 7160
rect 2571 7111 2613 7120
rect 2187 6824 2229 6833
rect 2187 6784 2188 6824
rect 2228 6784 2229 6824
rect 2187 6775 2229 6784
rect 1804 6404 1844 6413
rect 1804 6161 1844 6364
rect 2188 6404 2228 6775
rect 2379 6740 2421 6749
rect 2379 6700 2380 6740
rect 2420 6700 2421 6740
rect 2379 6691 2421 6700
rect 2380 6656 2420 6691
rect 2380 6605 2420 6616
rect 2188 6355 2228 6364
rect 2572 6404 2612 7111
rect 2763 6656 2805 6665
rect 2763 6616 2764 6656
rect 2804 6616 2805 6656
rect 2763 6607 2805 6616
rect 2764 6522 2804 6607
rect 2572 6355 2612 6364
rect 1995 6236 2037 6245
rect 1995 6196 1996 6236
rect 2036 6196 2037 6236
rect 1995 6187 2037 6196
rect 1803 6152 1845 6161
rect 1803 6112 1804 6152
rect 1844 6112 1845 6152
rect 1803 6103 1845 6112
rect 1996 6102 2036 6187
rect 1900 5732 1940 5741
rect 1900 5153 1940 5692
rect 3532 5657 3572 8716
rect 3628 8707 3668 8716
rect 3819 8756 3861 8765
rect 3819 8716 3820 8756
rect 3860 8716 3861 8756
rect 3819 8707 3861 8716
rect 4012 8756 4052 8765
rect 3915 8672 3957 8681
rect 3915 8632 3916 8672
rect 3956 8632 3957 8672
rect 3915 8623 3957 8632
rect 3916 8345 3956 8623
rect 3915 8336 3957 8345
rect 3915 8296 3916 8336
rect 3956 8296 3957 8336
rect 3915 8287 3957 8296
rect 4012 7925 4052 8716
rect 4875 8756 4917 8765
rect 4875 8716 4876 8756
rect 4916 8716 4917 8756
rect 4875 8707 4917 8716
rect 4972 8756 5012 8765
rect 4972 8504 5012 8716
rect 5739 8756 5781 8765
rect 5739 8716 5740 8756
rect 5780 8716 5781 8756
rect 5739 8707 5781 8716
rect 5932 8756 5972 8765
rect 4780 8464 5012 8504
rect 4011 7916 4053 7925
rect 4011 7876 4012 7916
rect 4052 7876 4053 7916
rect 4011 7867 4053 7876
rect 3688 7580 4056 7589
rect 3728 7540 3770 7580
rect 3810 7540 3852 7580
rect 3892 7540 3934 7580
rect 3974 7540 4016 7580
rect 3688 7531 4056 7540
rect 4780 6917 4820 8464
rect 4928 8336 5296 8345
rect 4968 8296 5010 8336
rect 5050 8296 5092 8336
rect 5132 8296 5174 8336
rect 5214 8296 5256 8336
rect 4928 8287 5296 8296
rect 5163 7916 5205 7925
rect 5163 7876 5164 7916
rect 5204 7876 5205 7916
rect 5163 7867 5205 7876
rect 5164 7001 5204 7867
rect 5932 7589 5972 8716
rect 6027 8756 6069 8765
rect 6027 8716 6028 8756
rect 6068 8716 6069 8756
rect 6027 8707 6069 8716
rect 6604 8706 6644 8791
rect 6892 8765 6932 8884
rect 7852 8840 7892 8851
rect 8716 8849 8756 10672
rect 8811 9680 8853 9689
rect 8811 9640 8812 9680
rect 8852 9640 8853 9680
rect 8811 9631 8853 9640
rect 8812 8924 8852 9631
rect 8812 8875 8852 8884
rect 9676 8849 9716 10672
rect 10636 8924 10676 10672
rect 11596 10604 11636 10672
rect 11788 10604 11828 10692
rect 11596 10564 11828 10604
rect 11211 9176 11253 9185
rect 11211 9136 11212 9176
rect 11252 9136 11253 9176
rect 11211 9127 11253 9136
rect 11403 9176 11445 9185
rect 11403 9136 11404 9176
rect 11444 9136 11445 9176
rect 11403 9127 11445 9136
rect 10636 8884 10772 8924
rect 7852 8765 7892 8800
rect 8715 8840 8757 8849
rect 8715 8800 8716 8840
rect 8756 8800 8757 8840
rect 8715 8791 8757 8800
rect 9387 8840 9429 8849
rect 9387 8800 9388 8840
rect 9428 8800 9429 8840
rect 9387 8791 9429 8800
rect 9675 8840 9717 8849
rect 9675 8800 9676 8840
rect 9716 8800 9717 8840
rect 9675 8791 9717 8800
rect 10443 8840 10485 8849
rect 10443 8800 10444 8840
rect 10484 8800 10485 8840
rect 10443 8791 10485 8800
rect 6796 8756 6836 8765
rect 5931 7580 5973 7589
rect 5931 7540 5932 7580
rect 5972 7540 5973 7580
rect 5931 7531 5973 7540
rect 5163 6992 5205 7001
rect 5163 6952 5164 6992
rect 5204 6952 5205 6992
rect 5163 6943 5205 6952
rect 4779 6908 4821 6917
rect 4779 6868 4780 6908
rect 4820 6868 4821 6908
rect 4779 6859 4821 6868
rect 4928 6824 5296 6833
rect 4968 6784 5010 6824
rect 5050 6784 5092 6824
rect 5132 6784 5174 6824
rect 5214 6784 5256 6824
rect 4928 6775 5296 6784
rect 3688 6068 4056 6077
rect 3728 6028 3770 6068
rect 3810 6028 3852 6068
rect 3892 6028 3934 6068
rect 3974 6028 4016 6068
rect 3688 6019 4056 6028
rect 6796 5741 6836 8716
rect 6891 8756 6933 8765
rect 6891 8716 6892 8756
rect 6932 8716 6933 8756
rect 6891 8707 6933 8716
rect 7851 8756 7893 8765
rect 7851 8716 7852 8756
rect 7892 8716 7893 8756
rect 7851 8707 7893 8716
rect 8044 8756 8084 8765
rect 7371 7580 7413 7589
rect 7371 7540 7372 7580
rect 7412 7540 7413 7580
rect 7371 7531 7413 7540
rect 7372 5909 7412 7531
rect 7371 5900 7413 5909
rect 7371 5860 7372 5900
rect 7412 5860 7413 5900
rect 7371 5851 7413 5860
rect 6795 5732 6837 5741
rect 6795 5692 6796 5732
rect 6836 5692 6837 5732
rect 6795 5683 6837 5692
rect 3531 5648 3573 5657
rect 3531 5608 3532 5648
rect 3572 5608 3573 5648
rect 3531 5599 3573 5608
rect 2187 5564 2229 5573
rect 2092 5524 2188 5564
rect 2228 5524 2229 5564
rect 2092 5480 2132 5524
rect 2187 5515 2229 5524
rect 2092 5431 2132 5440
rect 4928 5312 5296 5321
rect 4968 5272 5010 5312
rect 5050 5272 5092 5312
rect 5132 5272 5174 5312
rect 5214 5272 5256 5312
rect 4928 5263 5296 5272
rect 1899 5144 1941 5153
rect 1899 5104 1900 5144
rect 1940 5104 1941 5144
rect 1899 5095 1941 5104
rect 1227 4976 1269 4985
rect 1227 4936 1228 4976
rect 1268 4936 1269 4976
rect 1227 4927 1269 4936
rect 1035 4388 1077 4397
rect 1035 4348 1036 4388
rect 1076 4348 1077 4388
rect 1035 4339 1077 4348
rect 1228 3137 1268 4927
rect 1899 4892 1941 4901
rect 1899 4852 1900 4892
rect 1940 4852 1941 4892
rect 1899 4843 1941 4852
rect 6411 4892 6453 4901
rect 6411 4852 6412 4892
rect 6452 4852 6453 4892
rect 6411 4843 6453 4852
rect 1900 4758 1940 4843
rect 2091 4724 2133 4733
rect 2091 4684 2092 4724
rect 2132 4684 2133 4724
rect 2091 4675 2133 4684
rect 2092 4590 2132 4675
rect 3688 4556 4056 4565
rect 3728 4516 3770 4556
rect 3810 4516 3852 4556
rect 3892 4516 3934 4556
rect 3974 4516 4016 4556
rect 3688 4507 4056 4516
rect 1899 4388 1941 4397
rect 1899 4348 1900 4388
rect 1940 4348 1941 4388
rect 1899 4339 1941 4348
rect 1900 4254 1940 4339
rect 3147 4304 3189 4313
rect 3147 4264 3148 4304
rect 3188 4264 3189 4304
rect 3147 4255 3189 4264
rect 2091 4220 2133 4229
rect 2091 4180 2092 4220
rect 2132 4180 2133 4220
rect 2091 4171 2133 4180
rect 2092 4086 2132 4171
rect 2475 3968 2517 3977
rect 2475 3928 2476 3968
rect 2516 3928 2517 3968
rect 2475 3919 2517 3928
rect 1900 3380 1940 3389
rect 1804 3340 1900 3380
rect 1227 3128 1269 3137
rect 1227 3088 1228 3128
rect 1268 3088 1269 3128
rect 1227 3079 1269 3088
rect 1804 2045 1844 3340
rect 1900 3331 1940 3340
rect 2091 3212 2133 3221
rect 2091 3172 2092 3212
rect 2132 3172 2133 3212
rect 2091 3163 2133 3172
rect 2092 3078 2132 3163
rect 1900 2708 1940 2717
rect 1940 2668 2420 2708
rect 1900 2659 1940 2668
rect 2092 2456 2132 2465
rect 2132 2416 2228 2456
rect 2092 2407 2132 2416
rect 2091 2288 2133 2297
rect 2091 2248 2092 2288
rect 2132 2248 2133 2288
rect 2091 2239 2133 2248
rect 2092 2120 2132 2239
rect 2092 2071 2132 2080
rect 1803 2036 1845 2045
rect 1803 1996 1804 2036
rect 1844 1996 1845 2036
rect 1803 1987 1845 1996
rect 1803 1868 1845 1877
rect 1803 1828 1804 1868
rect 1844 1828 1845 1868
rect 1803 1819 1845 1828
rect 1900 1868 1940 1877
rect 1804 80 1844 1819
rect 1900 785 1940 1828
rect 2188 1205 2228 2416
rect 2284 1868 2324 1877
rect 2187 1196 2229 1205
rect 2187 1156 2188 1196
rect 2228 1156 2229 1196
rect 2187 1147 2229 1156
rect 2284 944 2324 1828
rect 1996 904 2324 944
rect 1899 776 1941 785
rect 1899 736 1900 776
rect 1940 736 1941 776
rect 1899 727 1941 736
rect 1996 80 2036 904
rect 2187 776 2229 785
rect 2187 736 2188 776
rect 2228 736 2229 776
rect 2187 727 2229 736
rect 2188 80 2228 727
rect 2380 80 2420 2668
rect 2476 2120 2516 3919
rect 3148 3809 3188 4255
rect 3147 3800 3189 3809
rect 3147 3760 3148 3800
rect 3188 3760 3189 3800
rect 3147 3751 3189 3760
rect 4928 3800 5296 3809
rect 4968 3760 5010 3800
rect 5050 3760 5092 3800
rect 5132 3760 5174 3800
rect 5214 3760 5256 3800
rect 4928 3751 5296 3760
rect 6412 3473 6452 4843
rect 6987 3800 7029 3809
rect 6987 3760 6988 3800
rect 7028 3760 7029 3800
rect 6987 3751 7029 3760
rect 6411 3464 6453 3473
rect 6411 3424 6412 3464
rect 6452 3424 6453 3464
rect 6411 3415 6453 3424
rect 3531 3296 3573 3305
rect 3531 3256 3532 3296
rect 3572 3256 3573 3296
rect 3531 3247 3573 3256
rect 2955 2960 2997 2969
rect 2955 2920 2956 2960
rect 2996 2920 2997 2960
rect 2955 2911 2997 2920
rect 2956 2876 2996 2911
rect 3532 2876 3572 3247
rect 3688 3044 4056 3053
rect 3728 3004 3770 3044
rect 3810 3004 3852 3044
rect 3892 3004 3934 3044
rect 3974 3004 4016 3044
rect 3688 2995 4056 3004
rect 6219 3044 6261 3053
rect 6219 3004 6220 3044
rect 6260 3004 6261 3044
rect 6219 2995 6261 3004
rect 3724 2876 3764 2885
rect 3532 2836 3724 2876
rect 2956 2825 2996 2836
rect 3724 2827 3764 2836
rect 6027 2876 6069 2885
rect 6027 2836 6028 2876
rect 6068 2836 6069 2876
rect 6027 2827 6069 2836
rect 2476 2071 2516 2080
rect 2764 2708 2804 2717
rect 3532 2708 3572 2717
rect 2571 2036 2613 2045
rect 2571 1996 2572 2036
rect 2612 1996 2613 2036
rect 2571 1987 2613 1996
rect 2572 80 2612 1987
rect 2667 1868 2709 1877
rect 2667 1828 2668 1868
rect 2708 1828 2709 1868
rect 2667 1819 2709 1828
rect 2668 1734 2708 1819
rect 2764 80 2804 2668
rect 3052 2668 3532 2708
rect 2859 2120 2901 2129
rect 2859 2080 2860 2120
rect 2900 2080 2901 2120
rect 2859 2071 2901 2080
rect 2860 1986 2900 2071
rect 3052 1364 3092 2668
rect 3532 2659 3572 2668
rect 5931 2708 5973 2717
rect 5931 2668 5932 2708
rect 5972 2668 5973 2708
rect 5931 2659 5973 2668
rect 4928 2288 5296 2297
rect 4968 2248 5010 2288
rect 5050 2248 5092 2288
rect 5132 2248 5174 2288
rect 5214 2248 5256 2288
rect 4928 2239 5296 2248
rect 5355 2120 5397 2129
rect 5355 2080 5356 2120
rect 5396 2080 5397 2120
rect 5355 2071 5397 2080
rect 5356 1986 5396 2071
rect 3724 1868 3764 1877
rect 2956 1324 3092 1364
rect 3148 1828 3724 1868
rect 2956 80 2996 1324
rect 3148 80 3188 1828
rect 3724 1819 3764 1828
rect 4108 1868 4148 1877
rect 3916 1709 3956 1794
rect 3915 1700 3957 1709
rect 3915 1660 3916 1700
rect 3956 1660 3957 1700
rect 3915 1651 3957 1660
rect 3688 1532 4056 1541
rect 3728 1492 3770 1532
rect 3810 1492 3852 1532
rect 3892 1492 3934 1532
rect 3974 1492 4016 1532
rect 3688 1483 4056 1492
rect 3339 1364 3381 1373
rect 3339 1324 3340 1364
rect 3380 1324 3381 1364
rect 3339 1315 3381 1324
rect 3340 80 3380 1315
rect 4108 1289 4148 1828
rect 4203 1868 4245 1877
rect 4203 1828 4204 1868
rect 4244 1828 4245 1868
rect 4203 1819 4245 1828
rect 4492 1868 4532 1877
rect 3531 1280 3573 1289
rect 3531 1240 3532 1280
rect 3572 1240 3573 1280
rect 3531 1231 3573 1240
rect 4107 1280 4149 1289
rect 4107 1240 4108 1280
rect 4148 1240 4149 1280
rect 4107 1231 4149 1240
rect 3532 80 3572 1231
rect 3723 944 3765 953
rect 4204 944 4244 1819
rect 4300 1700 4340 1709
rect 4340 1660 4436 1700
rect 4300 1651 4340 1660
rect 4299 1280 4341 1289
rect 4299 1240 4300 1280
rect 4340 1240 4341 1280
rect 4299 1231 4341 1240
rect 3723 904 3724 944
rect 3764 904 3765 944
rect 3723 895 3765 904
rect 4108 904 4244 944
rect 3724 80 3764 895
rect 3915 860 3957 869
rect 3915 820 3916 860
rect 3956 820 3957 860
rect 3915 811 3957 820
rect 3916 80 3956 811
rect 4108 80 4148 904
rect 4300 80 4340 1231
rect 4396 281 4436 1660
rect 4492 1373 4532 1828
rect 5163 1868 5205 1877
rect 5163 1828 5164 1868
rect 5204 1828 5205 1868
rect 5163 1819 5205 1828
rect 5451 1868 5493 1877
rect 5451 1828 5452 1868
rect 5492 1828 5493 1868
rect 5451 1819 5493 1828
rect 5644 1868 5684 1877
rect 5164 1734 5204 1819
rect 4684 1700 4724 1709
rect 4684 1541 4724 1660
rect 4779 1700 4821 1709
rect 4779 1660 4780 1700
rect 4820 1660 4821 1700
rect 4779 1651 4821 1660
rect 4683 1532 4725 1541
rect 4683 1492 4684 1532
rect 4724 1492 4725 1532
rect 4683 1483 4725 1492
rect 4587 1448 4629 1457
rect 4587 1408 4588 1448
rect 4628 1408 4629 1448
rect 4587 1399 4629 1408
rect 4491 1364 4533 1373
rect 4491 1324 4492 1364
rect 4532 1324 4533 1364
rect 4491 1315 4533 1324
rect 4588 944 4628 1399
rect 4683 1364 4725 1373
rect 4683 1324 4684 1364
rect 4724 1324 4725 1364
rect 4683 1315 4725 1324
rect 4492 904 4628 944
rect 4395 272 4437 281
rect 4395 232 4396 272
rect 4436 232 4437 272
rect 4395 223 4437 232
rect 4492 80 4532 904
rect 4684 80 4724 1315
rect 4780 197 4820 1651
rect 4928 776 5296 785
rect 4968 736 5010 776
rect 5050 736 5092 776
rect 5132 736 5174 776
rect 5214 736 5256 776
rect 4928 727 5296 736
rect 4875 608 4917 617
rect 4875 568 4876 608
rect 4916 568 4917 608
rect 4875 559 4917 568
rect 4779 188 4821 197
rect 4779 148 4780 188
rect 4820 148 4821 188
rect 4779 139 4821 148
rect 4876 80 4916 559
rect 5067 524 5109 533
rect 5067 484 5068 524
rect 5108 484 5109 524
rect 5067 475 5109 484
rect 5068 80 5108 475
rect 5259 356 5301 365
rect 5259 316 5260 356
rect 5300 316 5301 356
rect 5259 307 5301 316
rect 5260 80 5300 307
rect 5452 80 5492 1819
rect 5644 1289 5684 1828
rect 5835 1700 5877 1709
rect 5835 1660 5836 1700
rect 5876 1660 5877 1700
rect 5835 1651 5877 1660
rect 5836 1566 5876 1651
rect 5643 1280 5685 1289
rect 5835 1280 5877 1289
rect 5643 1240 5644 1280
rect 5684 1240 5685 1280
rect 5643 1231 5685 1240
rect 5740 1240 5836 1280
rect 5876 1240 5877 1280
rect 5740 692 5780 1240
rect 5835 1231 5877 1240
rect 5644 652 5780 692
rect 5644 80 5684 652
rect 5932 524 5972 2659
rect 5836 484 5972 524
rect 5836 80 5876 484
rect 6028 80 6068 2827
rect 6124 1868 6164 1877
rect 6124 1457 6164 1828
rect 6123 1448 6165 1457
rect 6123 1408 6124 1448
rect 6164 1408 6165 1448
rect 6123 1399 6165 1408
rect 6220 80 6260 2995
rect 6891 2792 6933 2801
rect 6891 2752 6892 2792
rect 6932 2752 6933 2792
rect 6891 2743 6933 2752
rect 6700 2708 6740 2717
rect 6316 1700 6356 1709
rect 6316 1457 6356 1660
rect 6315 1448 6357 1457
rect 6315 1408 6316 1448
rect 6356 1408 6357 1448
rect 6315 1399 6357 1408
rect 6700 1373 6740 2668
rect 6892 2658 6932 2743
rect 6892 1868 6932 1877
rect 6795 1616 6837 1625
rect 6795 1576 6796 1616
rect 6836 1576 6837 1616
rect 6795 1567 6837 1576
rect 6699 1364 6741 1373
rect 6699 1324 6700 1364
rect 6740 1324 6741 1364
rect 6699 1315 6741 1324
rect 6603 944 6645 953
rect 6603 904 6604 944
rect 6644 904 6645 944
rect 6603 895 6645 904
rect 6411 440 6453 449
rect 6411 400 6412 440
rect 6452 400 6453 440
rect 6411 391 6453 400
rect 6412 80 6452 391
rect 6604 80 6644 895
rect 6796 80 6836 1567
rect 6892 617 6932 1828
rect 6891 608 6933 617
rect 6891 568 6892 608
rect 6932 568 6933 608
rect 6891 559 6933 568
rect 6988 80 7028 3751
rect 8044 3137 8084 8716
rect 9004 8756 9044 8765
rect 9004 5153 9044 8716
rect 9388 8706 9428 8791
rect 9580 8756 9620 8765
rect 9003 5144 9045 5153
rect 9003 5104 9004 5144
rect 9044 5104 9045 5144
rect 9003 5095 9045 5104
rect 9580 5069 9620 8716
rect 10444 8706 10484 8791
rect 10732 8765 10772 8884
rect 10636 8756 10676 8765
rect 9579 5060 9621 5069
rect 9579 5020 9580 5060
rect 9620 5020 9621 5060
rect 9579 5011 9621 5020
rect 9099 3968 9141 3977
rect 9099 3928 9100 3968
rect 9140 3928 9141 3968
rect 9099 3919 9141 3928
rect 8043 3128 8085 3137
rect 8043 3088 8044 3128
rect 8084 3088 8085 3128
rect 8043 3079 8085 3088
rect 8716 2708 8756 2717
rect 7756 2668 8716 2708
rect 7371 2624 7413 2633
rect 7371 2584 7372 2624
rect 7412 2584 7413 2624
rect 7371 2575 7413 2584
rect 7275 1868 7317 1877
rect 7275 1828 7276 1868
rect 7316 1828 7317 1868
rect 7275 1819 7317 1828
rect 7276 1734 7316 1819
rect 7372 1709 7412 2575
rect 7660 1868 7700 1877
rect 7084 1700 7124 1709
rect 7084 785 7124 1660
rect 7371 1700 7413 1709
rect 7371 1660 7372 1700
rect 7412 1660 7413 1700
rect 7371 1651 7413 1660
rect 7468 1700 7508 1709
rect 7179 1364 7221 1373
rect 7179 1324 7180 1364
rect 7220 1324 7221 1364
rect 7179 1315 7221 1324
rect 7083 776 7125 785
rect 7083 736 7084 776
rect 7124 736 7125 776
rect 7083 727 7125 736
rect 7180 80 7220 1315
rect 7468 701 7508 1660
rect 7660 869 7700 1828
rect 7659 860 7701 869
rect 7659 820 7660 860
rect 7700 820 7701 860
rect 7659 811 7701 820
rect 7467 692 7509 701
rect 7467 652 7468 692
rect 7508 652 7509 692
rect 7467 643 7509 652
rect 7563 608 7605 617
rect 7563 568 7564 608
rect 7604 568 7605 608
rect 7563 559 7605 568
rect 7371 104 7413 113
rect 7371 80 7372 104
rect 1784 0 1864 80
rect 1976 0 2056 80
rect 2168 0 2248 80
rect 2360 0 2440 80
rect 2552 0 2632 80
rect 2744 0 2824 80
rect 2936 0 3016 80
rect 3128 0 3208 80
rect 3320 0 3400 80
rect 3512 0 3592 80
rect 3704 0 3784 80
rect 3896 0 3976 80
rect 4088 0 4168 80
rect 4280 0 4360 80
rect 4472 0 4552 80
rect 4664 0 4744 80
rect 4856 0 4936 80
rect 5048 0 5128 80
rect 5240 0 5320 80
rect 5432 0 5512 80
rect 5624 0 5704 80
rect 5816 0 5896 80
rect 6008 0 6088 80
rect 6200 0 6280 80
rect 6392 0 6472 80
rect 6584 0 6664 80
rect 6776 0 6856 80
rect 6968 0 7048 80
rect 7160 0 7240 80
rect 7352 64 7372 80
rect 7412 80 7413 104
rect 7564 80 7604 559
rect 7756 80 7796 2668
rect 8716 2659 8756 2668
rect 8331 2540 8373 2549
rect 8331 2500 8332 2540
rect 8372 2500 8373 2540
rect 8331 2491 8373 2500
rect 8044 1868 8084 1877
rect 7852 1700 7892 1709
rect 7852 953 7892 1660
rect 8044 1037 8084 1828
rect 8139 1868 8181 1877
rect 8139 1828 8140 1868
rect 8180 1828 8181 1868
rect 8139 1819 8181 1828
rect 8043 1028 8085 1037
rect 8043 988 8044 1028
rect 8084 988 8085 1028
rect 8043 979 8085 988
rect 7851 944 7893 953
rect 7851 904 7852 944
rect 7892 904 7893 944
rect 7851 895 7893 904
rect 8140 440 8180 1819
rect 8235 1700 8277 1709
rect 8235 1660 8236 1700
rect 8276 1660 8277 1700
rect 8235 1651 8277 1660
rect 8236 1566 8276 1651
rect 8235 1280 8277 1289
rect 8235 1240 8236 1280
rect 8276 1240 8277 1280
rect 8235 1231 8277 1240
rect 8044 400 8180 440
rect 8044 356 8084 400
rect 8236 356 8276 1231
rect 8044 316 8095 356
rect 8055 272 8095 316
rect 8044 232 8095 272
rect 8140 316 8276 356
rect 8044 188 8084 232
rect 8026 148 8084 188
rect 8026 104 8066 148
rect 7948 80 8066 104
rect 8140 80 8180 316
rect 8332 80 8372 2491
rect 8908 2456 8948 2465
rect 8811 2372 8853 2381
rect 8811 2332 8812 2372
rect 8852 2332 8853 2372
rect 8811 2323 8853 2332
rect 8428 1868 8468 1877
rect 8428 617 8468 1828
rect 8620 1700 8660 1709
rect 8523 860 8565 869
rect 8523 820 8524 860
rect 8564 820 8565 860
rect 8523 811 8565 820
rect 8427 608 8469 617
rect 8427 568 8428 608
rect 8468 568 8469 608
rect 8427 559 8469 568
rect 8524 80 8564 811
rect 8620 617 8660 1660
rect 8715 1196 8757 1205
rect 8715 1156 8716 1196
rect 8756 1156 8757 1196
rect 8715 1147 8757 1156
rect 8619 608 8661 617
rect 8619 568 8620 608
rect 8660 568 8661 608
rect 8619 559 8661 568
rect 8716 80 8756 1147
rect 8812 272 8852 2323
rect 8908 449 8948 2416
rect 8907 440 8949 449
rect 8907 400 8908 440
rect 8948 400 8949 440
rect 8907 391 8949 400
rect 8812 232 8948 272
rect 8908 80 8948 232
rect 9100 80 9140 3919
rect 10443 3296 10485 3305
rect 10443 3256 10444 3296
rect 10484 3256 10485 3296
rect 10443 3247 10485 3256
rect 9676 2708 9716 2717
rect 9676 2549 9716 2668
rect 9675 2540 9717 2549
rect 9675 2500 9676 2540
rect 9716 2500 9717 2540
rect 9675 2491 9717 2500
rect 9868 2456 9908 2465
rect 9291 2036 9333 2045
rect 9291 1996 9292 2036
rect 9332 1996 9333 2036
rect 9291 1987 9333 1996
rect 9292 80 9332 1987
rect 9675 1700 9717 1709
rect 9675 1660 9676 1700
rect 9716 1660 9717 1700
rect 9675 1651 9717 1660
rect 9483 944 9525 953
rect 9483 904 9484 944
rect 9524 904 9525 944
rect 9483 895 9525 904
rect 9484 80 9524 895
rect 9676 80 9716 1651
rect 9868 1205 9908 2416
rect 9964 1868 10004 1877
rect 9867 1196 9909 1205
rect 9867 1156 9868 1196
rect 9908 1156 9909 1196
rect 9867 1147 9909 1156
rect 9964 533 10004 1828
rect 10348 1868 10388 1877
rect 10156 1700 10196 1709
rect 10059 1532 10101 1541
rect 10059 1492 10060 1532
rect 10100 1492 10101 1532
rect 10059 1483 10101 1492
rect 9963 524 10005 533
rect 9963 484 9964 524
rect 10004 484 10005 524
rect 9963 475 10005 484
rect 9867 272 9909 281
rect 9867 232 9868 272
rect 9908 232 9909 272
rect 9867 223 9909 232
rect 9868 80 9908 223
rect 10060 80 10100 1483
rect 10156 953 10196 1660
rect 10155 944 10197 953
rect 10155 904 10156 944
rect 10196 904 10197 944
rect 10155 895 10197 904
rect 10348 365 10388 1828
rect 10347 356 10389 365
rect 10347 316 10348 356
rect 10388 316 10389 356
rect 10347 307 10389 316
rect 10251 188 10293 197
rect 10251 148 10252 188
rect 10292 148 10293 188
rect 10251 139 10293 148
rect 10252 80 10292 139
rect 10444 80 10484 3247
rect 10539 2960 10581 2969
rect 10539 2920 10540 2960
rect 10580 2920 10581 2960
rect 10539 2911 10581 2920
rect 10540 1868 10580 2911
rect 10636 2297 10676 8716
rect 10731 8756 10773 8765
rect 10731 8716 10732 8756
rect 10772 8716 10773 8756
rect 10731 8707 10773 8716
rect 11212 8756 11252 9127
rect 11404 8840 11444 9127
rect 11404 8791 11444 8800
rect 11596 8840 11636 8851
rect 11596 8765 11636 8800
rect 11980 8840 12020 10692
rect 12536 10672 12616 10752
rect 13496 10672 13576 10752
rect 14456 10672 14536 10752
rect 15416 10672 15496 10752
rect 15628 10692 16148 10732
rect 12556 8849 12596 10672
rect 13516 8849 13556 10672
rect 14476 8849 14516 10672
rect 15436 10604 15476 10672
rect 15628 10604 15668 10692
rect 15436 10564 15668 10604
rect 11980 8791 12020 8800
rect 12555 8840 12597 8849
rect 12555 8800 12556 8840
rect 12596 8800 12597 8840
rect 12555 8791 12597 8800
rect 13035 8840 13077 8849
rect 13035 8800 13036 8840
rect 13076 8800 13077 8840
rect 13035 8791 13077 8800
rect 13515 8840 13557 8849
rect 13515 8800 13516 8840
rect 13556 8800 13557 8840
rect 13515 8791 13557 8800
rect 14091 8840 14133 8849
rect 14091 8800 14092 8840
rect 14132 8800 14133 8840
rect 14091 8791 14133 8800
rect 14475 8840 14517 8849
rect 14475 8800 14476 8840
rect 14516 8800 14517 8840
rect 14475 8791 14517 8800
rect 15435 8840 15477 8849
rect 15435 8800 15436 8840
rect 15476 8800 15477 8840
rect 15435 8791 15477 8800
rect 16108 8840 16148 10692
rect 16376 10672 16456 10752
rect 17336 10672 17416 10752
rect 17836 10692 18164 10732
rect 16203 9512 16245 9521
rect 16203 9472 16204 9512
rect 16244 9472 16245 9512
rect 16203 9463 16245 9472
rect 16108 8791 16148 8800
rect 11212 8707 11252 8716
rect 11595 8756 11637 8765
rect 11595 8716 11596 8756
rect 11636 8716 11637 8756
rect 11595 8707 11637 8716
rect 11788 8756 11828 8765
rect 10731 3212 10773 3221
rect 10731 3172 10732 3212
rect 10772 3172 10773 3212
rect 10731 3163 10773 3172
rect 10635 2288 10677 2297
rect 10635 2248 10636 2288
rect 10676 2248 10677 2288
rect 10635 2239 10677 2248
rect 10540 1828 10676 1868
rect 10540 1700 10580 1709
rect 10540 1037 10580 1660
rect 10539 1028 10581 1037
rect 10539 988 10540 1028
rect 10580 988 10581 1028
rect 10539 979 10581 988
rect 10636 80 10676 1828
rect 10732 272 10772 3163
rect 11691 2792 11733 2801
rect 11691 2752 11692 2792
rect 11732 2752 11733 2792
rect 11691 2743 11733 2752
rect 10828 1868 10868 1877
rect 10828 869 10868 1828
rect 11211 1868 11253 1877
rect 11211 1828 11212 1868
rect 11252 1828 11253 1868
rect 11211 1819 11253 1828
rect 11596 1868 11636 1877
rect 11212 1734 11252 1819
rect 11020 1700 11060 1709
rect 11020 869 11060 1660
rect 11404 1700 11444 1709
rect 11404 1121 11444 1660
rect 11596 1289 11636 1828
rect 11595 1280 11637 1289
rect 11595 1240 11596 1280
rect 11636 1240 11637 1280
rect 11595 1231 11637 1240
rect 11403 1112 11445 1121
rect 11403 1072 11404 1112
rect 11444 1072 11445 1112
rect 11403 1063 11445 1072
rect 11211 1028 11253 1037
rect 11211 988 11212 1028
rect 11252 988 11253 1028
rect 11211 979 11253 988
rect 10827 860 10869 869
rect 10827 820 10828 860
rect 10868 820 10869 860
rect 10827 811 10869 820
rect 11019 860 11061 869
rect 11019 820 11020 860
rect 11060 820 11061 860
rect 11019 811 11061 820
rect 11019 692 11061 701
rect 11019 652 11020 692
rect 11060 652 11061 692
rect 11019 643 11061 652
rect 10732 232 10868 272
rect 10828 80 10868 232
rect 11020 80 11060 643
rect 11212 80 11252 979
rect 11403 944 11445 953
rect 11403 904 11404 944
rect 11444 904 11445 944
rect 11403 895 11445 904
rect 11404 80 11444 895
rect 11595 776 11637 785
rect 11595 736 11596 776
rect 11636 736 11637 776
rect 11692 776 11732 2743
rect 11788 2465 11828 8716
rect 12172 8756 12212 8765
rect 12172 6320 12212 8716
rect 13036 8706 13076 8791
rect 13228 8756 13268 8765
rect 13228 6320 13268 8716
rect 14092 8706 14132 8791
rect 14284 8756 14324 8765
rect 13611 8420 13653 8429
rect 13611 8380 13612 8420
rect 13652 8380 13653 8420
rect 13611 8371 13653 8380
rect 13612 7916 13652 8371
rect 13612 7867 13652 7876
rect 13803 7832 13845 7841
rect 13803 7792 13804 7832
rect 13844 7792 13845 7832
rect 13803 7783 13845 7792
rect 13804 7698 13844 7783
rect 12172 6280 12308 6320
rect 13228 6280 13364 6320
rect 11787 2456 11829 2465
rect 11787 2416 11788 2456
rect 11828 2416 11829 2456
rect 11787 2407 11829 2416
rect 11980 1868 12020 1877
rect 11884 1828 11980 1868
rect 11788 1700 11828 1709
rect 11788 953 11828 1660
rect 11787 944 11829 953
rect 11787 904 11788 944
rect 11828 904 11829 944
rect 11787 895 11829 904
rect 11692 736 11828 776
rect 11595 727 11637 736
rect 11596 80 11636 727
rect 11788 80 11828 736
rect 11884 197 11924 1828
rect 11980 1819 12020 1828
rect 12075 1700 12117 1709
rect 12075 1660 12076 1700
rect 12116 1660 12117 1700
rect 12075 1651 12117 1660
rect 12172 1700 12212 1709
rect 11979 1448 12021 1457
rect 11979 1408 11980 1448
rect 12020 1408 12021 1448
rect 11979 1399 12021 1408
rect 11883 188 11925 197
rect 11883 148 11884 188
rect 11924 148 11925 188
rect 11883 139 11925 148
rect 11980 80 12020 1399
rect 12076 860 12116 1651
rect 12172 1037 12212 1660
rect 12171 1028 12213 1037
rect 12171 988 12172 1028
rect 12212 988 12213 1028
rect 12171 979 12213 988
rect 12076 820 12212 860
rect 12172 80 12212 820
rect 12268 701 12308 6280
rect 13227 3800 13269 3809
rect 13227 3760 13228 3800
rect 13268 3760 13269 3800
rect 13227 3751 13269 3760
rect 12363 2120 12405 2129
rect 12363 2080 12364 2120
rect 12404 2080 12405 2120
rect 12363 2071 12405 2080
rect 12267 692 12309 701
rect 12267 652 12268 692
rect 12308 652 12309 692
rect 12267 643 12309 652
rect 12364 80 12404 2071
rect 12844 1868 12884 1877
rect 12844 1373 12884 1828
rect 13228 1868 13268 3751
rect 13324 2129 13364 6280
rect 14284 3389 14324 8716
rect 15436 8706 15476 8791
rect 15628 8756 15668 8765
rect 15628 6320 15668 8716
rect 16204 8597 16244 9463
rect 16396 8840 16436 10672
rect 17356 9596 17396 10672
rect 17068 9556 17396 9596
rect 16492 8840 16532 8849
rect 16396 8800 16492 8840
rect 16492 8791 16532 8800
rect 17068 8840 17108 9556
rect 17068 8791 17108 8800
rect 17836 8840 17876 10692
rect 18124 10604 18164 10692
rect 18296 10672 18376 10752
rect 19256 10672 19336 10752
rect 19468 10692 19796 10732
rect 18316 10604 18356 10672
rect 18124 10564 18356 10604
rect 19276 10604 19316 10672
rect 19468 10604 19508 10692
rect 19276 10564 19508 10604
rect 19563 10520 19605 10529
rect 19563 10480 19564 10520
rect 19604 10480 19605 10520
rect 19563 10471 19605 10480
rect 18808 9092 19176 9101
rect 18848 9052 18890 9092
rect 18930 9052 18972 9092
rect 19012 9052 19054 9092
rect 19094 9052 19136 9092
rect 18808 9043 19176 9052
rect 18219 8924 18261 8933
rect 18219 8884 18220 8924
rect 18260 8884 18261 8924
rect 18219 8875 18261 8884
rect 17836 8791 17876 8800
rect 16300 8756 16340 8765
rect 16203 8588 16245 8597
rect 16203 8548 16204 8588
rect 16244 8548 16245 8588
rect 16203 8539 16245 8548
rect 16011 6992 16053 7001
rect 16011 6952 16012 6992
rect 16052 6952 16053 6992
rect 16011 6943 16053 6952
rect 15628 6280 15764 6320
rect 15627 4220 15669 4229
rect 15627 4180 15628 4220
rect 15668 4180 15669 4220
rect 15627 4171 15669 4180
rect 14283 3380 14325 3389
rect 14283 3340 14284 3380
rect 14324 3340 14325 3380
rect 14283 3331 14325 3340
rect 15147 3044 15189 3053
rect 15147 3004 15148 3044
rect 15188 3004 15189 3044
rect 15147 2995 15189 3004
rect 15148 2708 15188 2995
rect 15531 2876 15573 2885
rect 15531 2836 15532 2876
rect 15572 2836 15573 2876
rect 15531 2827 15573 2836
rect 15148 2659 15188 2668
rect 15532 2708 15572 2827
rect 15532 2659 15572 2668
rect 14956 2456 14996 2465
rect 15340 2456 15380 2465
rect 14860 2416 14956 2456
rect 13323 2120 13365 2129
rect 13323 2080 13324 2120
rect 13364 2080 13365 2120
rect 13323 2071 13365 2080
rect 13228 1819 13268 1828
rect 13612 1868 13652 1877
rect 13036 1700 13076 1709
rect 12843 1364 12885 1373
rect 12843 1324 12844 1364
rect 12884 1324 12885 1364
rect 12843 1315 12885 1324
rect 12747 1196 12789 1205
rect 12747 1156 12748 1196
rect 12788 1156 12789 1196
rect 12747 1147 12789 1156
rect 12555 860 12597 869
rect 12555 820 12556 860
rect 12596 820 12597 860
rect 12555 811 12597 820
rect 12556 80 12596 811
rect 12748 80 12788 1147
rect 12939 944 12981 953
rect 12939 904 12940 944
rect 12980 904 12981 944
rect 12939 895 12981 904
rect 12940 80 12980 895
rect 13036 785 13076 1660
rect 13420 1700 13460 1709
rect 13131 1112 13173 1121
rect 13131 1072 13132 1112
rect 13172 1072 13173 1112
rect 13131 1063 13173 1072
rect 13035 776 13077 785
rect 13035 736 13036 776
rect 13076 736 13077 776
rect 13035 727 13077 736
rect 13132 80 13172 1063
rect 13420 953 13460 1660
rect 13612 1625 13652 1828
rect 13996 1868 14036 1877
rect 13804 1700 13844 1709
rect 13611 1616 13653 1625
rect 13611 1576 13612 1616
rect 13652 1576 13653 1616
rect 13611 1567 13653 1576
rect 13707 1028 13749 1037
rect 13707 988 13708 1028
rect 13748 988 13749 1028
rect 13707 979 13749 988
rect 13419 944 13461 953
rect 13419 904 13420 944
rect 13460 904 13461 944
rect 13419 895 13461 904
rect 13515 608 13557 617
rect 13515 568 13516 608
rect 13556 568 13557 608
rect 13515 559 13557 568
rect 13323 440 13365 449
rect 13323 400 13324 440
rect 13364 400 13365 440
rect 13323 391 13365 400
rect 13324 80 13364 391
rect 13516 80 13556 559
rect 13708 80 13748 979
rect 13804 869 13844 1660
rect 13996 1121 14036 1828
rect 14572 1868 14612 1877
rect 14188 1700 14228 1709
rect 14228 1660 14516 1700
rect 14188 1651 14228 1660
rect 13995 1112 14037 1121
rect 13995 1072 13996 1112
rect 14036 1072 14037 1112
rect 13995 1063 14037 1072
rect 14091 944 14133 953
rect 14091 904 14092 944
rect 14132 904 14133 944
rect 14091 895 14133 904
rect 13803 860 13845 869
rect 13803 820 13804 860
rect 13844 820 13845 860
rect 13803 811 13845 820
rect 13899 776 13941 785
rect 13899 736 13900 776
rect 13940 736 13941 776
rect 13899 727 13941 736
rect 13900 80 13940 727
rect 14092 80 14132 895
rect 14283 860 14325 869
rect 14283 820 14284 860
rect 14324 820 14325 860
rect 14283 811 14325 820
rect 14284 80 14324 811
rect 14476 80 14516 1660
rect 14572 449 14612 1828
rect 14764 1700 14804 1709
rect 14668 1660 14764 1700
rect 14571 440 14613 449
rect 14571 400 14572 440
rect 14612 400 14613 440
rect 14571 391 14613 400
rect 14668 80 14708 1660
rect 14764 1651 14804 1660
rect 14860 80 14900 2416
rect 14956 2407 14996 2416
rect 15052 2416 15340 2456
rect 15052 80 15092 2416
rect 15340 2407 15380 2416
rect 15243 1868 15285 1877
rect 15243 1828 15244 1868
rect 15284 1828 15285 1868
rect 15243 1819 15285 1828
rect 15244 80 15284 1819
rect 15435 1700 15477 1709
rect 15435 1660 15436 1700
rect 15476 1660 15477 1700
rect 15435 1651 15477 1660
rect 15436 80 15476 1651
rect 15628 80 15668 4171
rect 15724 3305 15764 6280
rect 15819 5648 15861 5657
rect 15819 5608 15820 5648
rect 15860 5608 15861 5648
rect 15819 5599 15861 5608
rect 15723 3296 15765 3305
rect 15723 3256 15724 3296
rect 15764 3256 15765 3296
rect 15723 3247 15765 3256
rect 15820 80 15860 5599
rect 15916 2456 15956 2465
rect 15916 1877 15956 2416
rect 15915 1868 15957 1877
rect 15915 1828 15916 1868
rect 15956 1828 15957 1868
rect 15915 1819 15957 1828
rect 15915 1700 15957 1709
rect 15915 1660 15916 1700
rect 15956 1660 15957 1700
rect 15915 1651 15957 1660
rect 15916 1566 15956 1651
rect 16012 80 16052 6943
rect 16203 6908 16245 6917
rect 16203 6868 16204 6908
rect 16244 6868 16245 6908
rect 16203 6859 16245 6868
rect 16107 2708 16149 2717
rect 16107 2668 16108 2708
rect 16148 2668 16149 2708
rect 16107 2659 16149 2668
rect 16108 2574 16148 2659
rect 16107 1868 16149 1877
rect 16107 1828 16108 1868
rect 16148 1828 16149 1868
rect 16107 1819 16149 1828
rect 16108 1734 16148 1819
rect 16204 80 16244 6859
rect 16300 3221 16340 8716
rect 16684 8756 16724 8765
rect 16395 6404 16437 6413
rect 16395 6364 16396 6404
rect 16436 6364 16437 6404
rect 16395 6355 16437 6364
rect 16396 5825 16436 6355
rect 16684 6320 16724 8716
rect 16876 8756 16916 8765
rect 16876 6320 16916 8716
rect 17644 8756 17684 8765
rect 17644 6320 17684 8716
rect 18220 8756 18260 8875
rect 18411 8840 18453 8849
rect 18411 8800 18412 8840
rect 18452 8800 18453 8840
rect 18411 8791 18453 8800
rect 19564 8840 19604 10471
rect 19564 8791 19604 8800
rect 19756 8840 19796 10692
rect 20216 10672 20296 10752
rect 20236 10016 20276 10672
rect 20236 9976 20564 10016
rect 20048 9848 20416 9857
rect 20088 9808 20130 9848
rect 20170 9808 20212 9848
rect 20252 9808 20294 9848
rect 20334 9808 20376 9848
rect 20048 9799 20416 9808
rect 19756 8791 19796 8800
rect 18220 8707 18260 8716
rect 18412 8706 18452 8791
rect 18988 8756 19028 8765
rect 19372 8756 19412 8765
rect 19028 8716 19316 8756
rect 18988 8707 19028 8716
rect 19179 8504 19221 8513
rect 19179 8464 19180 8504
rect 19220 8464 19221 8504
rect 19179 8455 19221 8464
rect 19180 8370 19220 8455
rect 17931 8168 17973 8177
rect 17931 8128 17932 8168
rect 17972 8128 17973 8168
rect 17931 8119 17973 8128
rect 18123 8168 18165 8177
rect 18123 8128 18124 8168
rect 18164 8128 18165 8168
rect 18123 8119 18165 8128
rect 17932 6404 17972 8119
rect 18124 6656 18164 8119
rect 18808 7580 19176 7589
rect 18848 7540 18890 7580
rect 18930 7540 18972 7580
rect 19012 7540 19054 7580
rect 19094 7540 19136 7580
rect 18808 7531 19176 7540
rect 19276 7496 19316 8716
rect 19372 8009 19412 8716
rect 19948 8756 19988 8765
rect 19371 8000 19413 8009
rect 19371 7960 19372 8000
rect 19412 7960 19413 8000
rect 19371 7951 19413 7960
rect 19659 7496 19701 7505
rect 19276 7456 19412 7496
rect 19276 7244 19316 7253
rect 19180 7204 19276 7244
rect 18315 7160 18357 7169
rect 18315 7120 18316 7160
rect 18356 7120 18357 7160
rect 18315 7111 18357 7120
rect 18124 6607 18164 6616
rect 18316 6581 18356 7111
rect 18315 6572 18357 6581
rect 18315 6532 18316 6572
rect 18356 6532 18357 6572
rect 18315 6523 18357 6532
rect 19180 6497 19220 7204
rect 19276 7195 19316 7204
rect 19179 6488 19221 6497
rect 19179 6448 19180 6488
rect 19220 6448 19221 6488
rect 19179 6439 19221 6448
rect 19276 6413 19316 6498
rect 17932 6355 17972 6364
rect 19275 6404 19317 6413
rect 19275 6364 19276 6404
rect 19316 6364 19317 6404
rect 19275 6355 19317 6364
rect 16684 6280 16820 6320
rect 16876 6280 17012 6320
rect 17644 6280 17876 6320
rect 16491 5900 16533 5909
rect 16491 5860 16492 5900
rect 16532 5860 16533 5900
rect 16491 5851 16533 5860
rect 16395 5816 16437 5825
rect 16395 5776 16396 5816
rect 16436 5776 16437 5816
rect 16395 5767 16437 5776
rect 16395 5060 16437 5069
rect 16395 5020 16396 5060
rect 16436 5020 16437 5060
rect 16395 5011 16437 5020
rect 16299 3212 16341 3221
rect 16299 3172 16300 3212
rect 16340 3172 16341 3212
rect 16299 3163 16341 3172
rect 16396 2549 16436 5011
rect 16395 2540 16437 2549
rect 16395 2500 16396 2540
rect 16436 2500 16437 2540
rect 16395 2491 16437 2500
rect 16492 1280 16532 5851
rect 16587 5732 16629 5741
rect 16587 5692 16588 5732
rect 16628 5692 16629 5732
rect 16587 5683 16629 5692
rect 16396 1240 16532 1280
rect 16396 80 16436 1240
rect 16588 80 16628 5683
rect 16683 4892 16725 4901
rect 16683 4852 16684 4892
rect 16724 4852 16725 4892
rect 16683 4843 16725 4852
rect 16684 4758 16724 4843
rect 16780 3137 16820 6280
rect 16876 4724 16916 4733
rect 16876 3473 16916 4684
rect 16875 3464 16917 3473
rect 16875 3424 16876 3464
rect 16916 3424 16917 3464
rect 16875 3415 16917 3424
rect 16779 3128 16821 3137
rect 16779 3088 16780 3128
rect 16820 3088 16821 3128
rect 16779 3079 16821 3088
rect 16779 2960 16821 2969
rect 16779 2920 16780 2960
rect 16820 2920 16821 2960
rect 16779 2911 16821 2920
rect 16683 2540 16725 2549
rect 16683 2500 16684 2540
rect 16724 2500 16725 2540
rect 16683 2491 16725 2500
rect 16684 281 16724 2491
rect 16683 272 16725 281
rect 16683 232 16684 272
rect 16724 232 16725 272
rect 16683 223 16725 232
rect 16780 80 16820 2911
rect 16972 2885 17012 6280
rect 17067 5144 17109 5153
rect 17067 5104 17068 5144
rect 17108 5104 17109 5144
rect 17067 5095 17109 5104
rect 16971 2876 17013 2885
rect 16971 2836 16972 2876
rect 17012 2836 17013 2876
rect 16971 2827 17013 2836
rect 17068 2624 17108 5095
rect 17260 4892 17300 4901
rect 17260 4313 17300 4852
rect 17452 4724 17492 4733
rect 17259 4304 17301 4313
rect 17259 4264 17260 4304
rect 17300 4264 17301 4304
rect 17259 4255 17301 4264
rect 17452 3893 17492 4684
rect 17451 3884 17493 3893
rect 17451 3844 17452 3884
rect 17492 3844 17493 3884
rect 17451 3835 17493 3844
rect 17355 2708 17397 2717
rect 17355 2668 17356 2708
rect 17396 2668 17397 2708
rect 17355 2659 17397 2668
rect 16876 2584 17108 2624
rect 16876 1112 16916 2584
rect 17356 2574 17396 2659
rect 17067 2456 17109 2465
rect 17067 2416 17068 2456
rect 17108 2416 17109 2456
rect 17067 2407 17109 2416
rect 17548 2456 17588 2465
rect 16972 1868 17012 1877
rect 16972 1289 17012 1828
rect 16971 1280 17013 1289
rect 16971 1240 16972 1280
rect 17012 1240 17013 1280
rect 16971 1231 17013 1240
rect 16876 1072 17012 1112
rect 16972 80 17012 1072
rect 17068 785 17108 2407
rect 17259 2288 17301 2297
rect 17259 2248 17260 2288
rect 17300 2248 17301 2288
rect 17259 2239 17301 2248
rect 17164 1700 17204 1709
rect 17067 776 17109 785
rect 17067 736 17068 776
rect 17108 736 17109 776
rect 17067 727 17109 736
rect 17164 449 17204 1660
rect 17163 440 17205 449
rect 17163 400 17164 440
rect 17204 400 17205 440
rect 17260 440 17300 2239
rect 17356 1868 17396 1877
rect 17548 1868 17588 2416
rect 17739 1868 17781 1877
rect 17548 1828 17684 1868
rect 17356 1541 17396 1828
rect 17548 1700 17588 1709
rect 17452 1660 17548 1700
rect 17355 1532 17397 1541
rect 17355 1492 17356 1532
rect 17396 1492 17397 1532
rect 17355 1483 17397 1492
rect 17356 1196 17396 1205
rect 17356 617 17396 1156
rect 17355 608 17397 617
rect 17355 568 17356 608
rect 17396 568 17397 608
rect 17355 559 17397 568
rect 17260 400 17396 440
rect 17163 391 17205 400
rect 17163 272 17205 281
rect 17163 232 17164 272
rect 17204 232 17205 272
rect 17163 223 17205 232
rect 17164 80 17204 223
rect 17356 80 17396 400
rect 17452 197 17492 1660
rect 17548 1651 17588 1660
rect 17644 1457 17684 1828
rect 17739 1828 17740 1868
rect 17780 1828 17781 1868
rect 17739 1819 17781 1828
rect 17740 1734 17780 1819
rect 17643 1448 17685 1457
rect 17643 1408 17644 1448
rect 17684 1408 17685 1448
rect 17643 1399 17685 1408
rect 17836 1373 17876 6280
rect 18808 6068 19176 6077
rect 18848 6028 18890 6068
rect 18930 6028 18972 6068
rect 19012 6028 19054 6068
rect 19094 6028 19136 6068
rect 18808 6019 19176 6028
rect 19180 5732 19220 5741
rect 19180 5405 19220 5692
rect 19372 5648 19412 7456
rect 19659 7456 19660 7496
rect 19700 7456 19701 7496
rect 19659 7447 19701 7456
rect 19851 7496 19893 7505
rect 19851 7456 19852 7496
rect 19892 7456 19893 7496
rect 19851 7447 19893 7456
rect 19468 6992 19508 7001
rect 19468 6497 19508 6952
rect 19467 6488 19509 6497
rect 19467 6448 19468 6488
rect 19508 6448 19509 6488
rect 19467 6439 19509 6448
rect 19660 6404 19700 7447
rect 19852 6656 19892 7447
rect 19852 6607 19892 6616
rect 19660 6355 19700 6364
rect 19468 6236 19508 6245
rect 19468 5825 19508 6196
rect 19467 5816 19509 5825
rect 19467 5776 19468 5816
rect 19508 5776 19509 5816
rect 19467 5767 19509 5776
rect 19372 5608 19508 5648
rect 19371 5480 19413 5489
rect 19371 5440 19372 5480
rect 19412 5440 19413 5480
rect 19371 5431 19413 5440
rect 19179 5396 19221 5405
rect 19179 5356 19180 5396
rect 19220 5356 19221 5396
rect 19179 5347 19221 5356
rect 19372 5346 19412 5431
rect 18699 4976 18741 4985
rect 18699 4936 18700 4976
rect 18740 4936 18741 4976
rect 18699 4927 18741 4936
rect 18700 4220 18740 4927
rect 18808 4556 19176 4565
rect 18848 4516 18890 4556
rect 18930 4516 18972 4556
rect 19012 4516 19054 4556
rect 19094 4516 19136 4556
rect 18808 4507 19176 4516
rect 19371 4472 19413 4481
rect 19371 4432 19372 4472
rect 19412 4432 19413 4472
rect 19371 4423 19413 4432
rect 19179 4388 19221 4397
rect 19179 4348 19180 4388
rect 19220 4348 19221 4388
rect 19179 4339 19221 4348
rect 19372 4388 19412 4423
rect 18796 4220 18836 4229
rect 18700 4180 18796 4220
rect 18796 4171 18836 4180
rect 19180 4220 19220 4339
rect 19372 4337 19412 4348
rect 19180 4171 19220 4180
rect 18988 3968 19028 3977
rect 18123 3380 18165 3389
rect 18123 3340 18124 3380
rect 18164 3340 18165 3380
rect 18123 3331 18165 3340
rect 18027 2120 18069 2129
rect 18027 2080 18028 2120
rect 18068 2080 18069 2120
rect 18027 2071 18069 2080
rect 17932 1700 17972 1709
rect 17835 1364 17877 1373
rect 17835 1324 17836 1364
rect 17876 1324 17877 1364
rect 17835 1315 17877 1324
rect 17547 1112 17589 1121
rect 17547 1072 17548 1112
rect 17588 1072 17589 1112
rect 17547 1063 17589 1072
rect 17548 944 17588 1063
rect 17548 895 17588 904
rect 17932 869 17972 1660
rect 17931 860 17973 869
rect 17931 820 17932 860
rect 17972 820 17973 860
rect 17931 811 17973 820
rect 17547 776 17589 785
rect 17547 736 17548 776
rect 17588 736 17589 776
rect 17547 727 17589 736
rect 17451 188 17493 197
rect 17451 148 17452 188
rect 17492 148 17493 188
rect 17451 139 17493 148
rect 17548 80 17588 727
rect 17739 692 17781 701
rect 18028 692 18068 2071
rect 17739 652 17740 692
rect 17780 652 17781 692
rect 17739 643 17781 652
rect 17932 652 18068 692
rect 17740 80 17780 643
rect 17932 80 17972 652
rect 18124 80 18164 3331
rect 18315 3296 18357 3305
rect 18315 3256 18316 3296
rect 18356 3256 18357 3296
rect 18315 3247 18357 3256
rect 18316 80 18356 3247
rect 18988 3221 19028 3928
rect 19275 3380 19317 3389
rect 19275 3340 19276 3380
rect 19316 3340 19317 3380
rect 19468 3380 19508 5608
rect 19563 4220 19605 4229
rect 19563 4180 19564 4220
rect 19604 4180 19605 4220
rect 19563 4171 19605 4180
rect 19564 4086 19604 4171
rect 19755 4136 19797 4145
rect 19755 4096 19756 4136
rect 19796 4096 19797 4136
rect 19755 4087 19797 4096
rect 19756 3968 19796 4087
rect 19756 3919 19796 3928
rect 19468 3340 19604 3380
rect 19275 3331 19317 3340
rect 19276 3246 19316 3331
rect 18507 3212 18549 3221
rect 18507 3172 18508 3212
rect 18548 3172 18549 3212
rect 18507 3163 18549 3172
rect 18987 3212 19029 3221
rect 18987 3172 18988 3212
rect 19028 3172 19029 3212
rect 18987 3163 19029 3172
rect 19468 3212 19508 3221
rect 18508 80 18548 3163
rect 18603 3128 18645 3137
rect 18603 3088 18604 3128
rect 18644 3088 18645 3128
rect 18603 3079 18645 3088
rect 18604 1280 18644 3079
rect 18808 3044 19176 3053
rect 18848 3004 18890 3044
rect 18930 3004 18972 3044
rect 19012 3004 19054 3044
rect 19094 3004 19136 3044
rect 18808 2995 19176 3004
rect 19275 3044 19317 3053
rect 19275 3004 19276 3044
rect 19316 3004 19317 3044
rect 19275 2995 19317 3004
rect 18891 2876 18933 2885
rect 18891 2836 18892 2876
rect 18932 2836 18933 2876
rect 18891 2827 18933 2836
rect 18892 1700 18932 2827
rect 18987 1868 19029 1877
rect 18987 1828 18988 1868
rect 19028 1828 19029 1868
rect 18987 1819 19029 1828
rect 18988 1734 19028 1819
rect 19180 1793 19220 1878
rect 19179 1784 19221 1793
rect 19179 1744 19180 1784
rect 19220 1744 19221 1784
rect 19179 1735 19221 1744
rect 18700 1660 18932 1700
rect 18700 1364 18740 1660
rect 18808 1532 19176 1541
rect 18848 1492 18890 1532
rect 18930 1492 18972 1532
rect 19012 1492 19054 1532
rect 19094 1492 19136 1532
rect 18808 1483 19176 1492
rect 19083 1364 19125 1373
rect 18700 1324 18932 1364
rect 18604 1240 18740 1280
rect 18700 80 18740 1240
rect 18892 80 18932 1324
rect 19083 1324 19084 1364
rect 19124 1324 19125 1364
rect 19083 1315 19125 1324
rect 19084 80 19124 1315
rect 19276 80 19316 2995
rect 19468 2801 19508 3172
rect 19467 2792 19509 2801
rect 19467 2752 19468 2792
rect 19508 2752 19509 2792
rect 19467 2743 19509 2752
rect 19564 2624 19604 3340
rect 19948 3053 19988 8716
rect 20524 8513 20564 9976
rect 20619 9848 20661 9857
rect 20619 9808 20620 9848
rect 20660 9808 20661 9848
rect 20619 9799 20661 9808
rect 20620 8681 20660 9799
rect 20619 8672 20661 8681
rect 20619 8632 20620 8672
rect 20660 8632 20661 8672
rect 20619 8623 20661 8632
rect 20523 8504 20565 8513
rect 20523 8464 20524 8504
rect 20564 8464 20565 8504
rect 20523 8455 20565 8464
rect 21387 8504 21429 8513
rect 21387 8464 21388 8504
rect 21428 8464 21429 8504
rect 21387 8455 21429 8464
rect 20048 8336 20416 8345
rect 20088 8296 20130 8336
rect 20170 8296 20212 8336
rect 20252 8296 20294 8336
rect 20334 8296 20376 8336
rect 20048 8287 20416 8296
rect 21388 8009 21428 8455
rect 21387 8000 21429 8009
rect 21387 7960 21388 8000
rect 21428 7960 21429 8000
rect 21387 7951 21429 7960
rect 20048 6824 20416 6833
rect 20088 6784 20130 6824
rect 20170 6784 20212 6824
rect 20252 6784 20294 6824
rect 20334 6784 20376 6824
rect 20048 6775 20416 6784
rect 20048 5312 20416 5321
rect 20088 5272 20130 5312
rect 20170 5272 20212 5312
rect 20252 5272 20294 5312
rect 20334 5272 20376 5312
rect 20048 5263 20416 5272
rect 20048 3800 20416 3809
rect 20088 3760 20130 3800
rect 20170 3760 20212 3800
rect 20252 3760 20294 3800
rect 20334 3760 20376 3800
rect 20048 3751 20416 3760
rect 19947 3044 19989 3053
rect 19947 3004 19948 3044
rect 19988 3004 19989 3044
rect 19947 2995 19989 3004
rect 19468 2584 19604 2624
rect 19371 1868 19413 1877
rect 19371 1828 19372 1868
rect 19412 1828 19413 1868
rect 19371 1819 19413 1828
rect 19372 1734 19412 1819
rect 19468 80 19508 2584
rect 19563 2456 19605 2465
rect 19563 2416 19564 2456
rect 19604 2416 19605 2456
rect 19563 2407 19605 2416
rect 19564 2120 19604 2407
rect 20048 2288 20416 2297
rect 20088 2248 20130 2288
rect 20170 2248 20212 2288
rect 20252 2248 20294 2288
rect 20334 2248 20376 2288
rect 20048 2239 20416 2248
rect 19564 2071 19604 2080
rect 19947 2120 19989 2129
rect 19947 2080 19948 2120
rect 19988 2080 19989 2120
rect 19947 2071 19989 2080
rect 19948 1986 19988 2071
rect 19755 1868 19797 1877
rect 19755 1828 19756 1868
rect 19796 1828 19797 1868
rect 19755 1819 19797 1828
rect 19756 1734 19796 1819
rect 20048 776 20416 785
rect 20088 736 20130 776
rect 20170 736 20212 776
rect 20252 736 20294 776
rect 20334 736 20376 776
rect 20048 727 20416 736
rect 7412 64 7432 80
rect 7352 0 7432 64
rect 7544 0 7624 80
rect 7736 0 7816 80
rect 7928 64 8066 80
rect 7928 0 8008 64
rect 8120 0 8200 80
rect 8312 0 8392 80
rect 8504 0 8584 80
rect 8696 0 8776 80
rect 8888 0 8968 80
rect 9080 0 9160 80
rect 9272 0 9352 80
rect 9464 0 9544 80
rect 9656 0 9736 80
rect 9848 0 9928 80
rect 10040 0 10120 80
rect 10232 0 10312 80
rect 10424 0 10504 80
rect 10616 0 10696 80
rect 10808 0 10888 80
rect 11000 0 11080 80
rect 11192 0 11272 80
rect 11384 0 11464 80
rect 11576 0 11656 80
rect 11768 0 11848 80
rect 11960 0 12040 80
rect 12152 0 12232 80
rect 12344 0 12424 80
rect 12536 0 12616 80
rect 12728 0 12808 80
rect 12920 0 13000 80
rect 13112 0 13192 80
rect 13304 0 13384 80
rect 13496 0 13576 80
rect 13688 0 13768 80
rect 13880 0 13960 80
rect 14072 0 14152 80
rect 14264 0 14344 80
rect 14456 0 14536 80
rect 14648 0 14728 80
rect 14840 0 14920 80
rect 15032 0 15112 80
rect 15224 0 15304 80
rect 15416 0 15496 80
rect 15608 0 15688 80
rect 15800 0 15880 80
rect 15992 0 16072 80
rect 16184 0 16264 80
rect 16376 0 16456 80
rect 16568 0 16648 80
rect 16760 0 16840 80
rect 16952 0 17032 80
rect 17144 0 17224 80
rect 17336 0 17416 80
rect 17528 0 17608 80
rect 17720 0 17800 80
rect 17912 0 17992 80
rect 18104 0 18184 80
rect 18296 0 18376 80
rect 18488 0 18568 80
rect 18680 0 18760 80
rect 18872 0 18952 80
rect 19064 0 19144 80
rect 19256 0 19336 80
rect 19448 0 19528 80
<< via2 >>
rect 556 10480 596 10520
rect 556 7960 596 8000
rect 1516 9808 1556 9848
rect 1900 9472 1940 9512
rect 2284 10144 2324 10184
rect 3688 9052 3728 9092
rect 3770 9052 3810 9092
rect 3852 9052 3892 9092
rect 3934 9052 3974 9092
rect 4016 9052 4056 9092
rect 2956 8716 2996 8756
rect 4928 9808 4968 9848
rect 5010 9808 5050 9848
rect 5092 9808 5132 9848
rect 5174 9808 5214 9848
rect 5256 9808 5296 9848
rect 7756 9640 7796 9680
rect 6604 8800 6644 8840
rect 1996 8632 2036 8672
rect 3436 8632 3476 8672
rect 2092 8464 2132 8504
rect 2476 8464 2516 8504
rect 1708 8296 1748 8336
rect 2188 7876 2228 7916
rect 2380 7708 2420 7748
rect 2572 7120 2612 7160
rect 2188 6784 2228 6824
rect 2380 6700 2420 6740
rect 2764 6616 2804 6656
rect 1996 6196 2036 6236
rect 1804 6112 1844 6152
rect 3820 8716 3860 8756
rect 3916 8632 3956 8672
rect 3916 8296 3956 8336
rect 4876 8716 4916 8756
rect 5740 8716 5780 8756
rect 4012 7876 4052 7916
rect 3688 7540 3728 7580
rect 3770 7540 3810 7580
rect 3852 7540 3892 7580
rect 3934 7540 3974 7580
rect 4016 7540 4056 7580
rect 4928 8296 4968 8336
rect 5010 8296 5050 8336
rect 5092 8296 5132 8336
rect 5174 8296 5214 8336
rect 5256 8296 5296 8336
rect 5164 7876 5204 7916
rect 6028 8716 6068 8756
rect 8812 9640 8852 9680
rect 11212 9136 11252 9176
rect 11404 9136 11444 9176
rect 8716 8800 8756 8840
rect 9388 8800 9428 8840
rect 9676 8800 9716 8840
rect 10444 8800 10484 8840
rect 5932 7540 5972 7580
rect 5164 6952 5204 6992
rect 4780 6868 4820 6908
rect 4928 6784 4968 6824
rect 5010 6784 5050 6824
rect 5092 6784 5132 6824
rect 5174 6784 5214 6824
rect 5256 6784 5296 6824
rect 3688 6028 3728 6068
rect 3770 6028 3810 6068
rect 3852 6028 3892 6068
rect 3934 6028 3974 6068
rect 4016 6028 4056 6068
rect 6892 8716 6932 8756
rect 7852 8716 7892 8756
rect 7372 7540 7412 7580
rect 7372 5860 7412 5900
rect 6796 5692 6836 5732
rect 3532 5608 3572 5648
rect 2188 5524 2228 5564
rect 4928 5272 4968 5312
rect 5010 5272 5050 5312
rect 5092 5272 5132 5312
rect 5174 5272 5214 5312
rect 5256 5272 5296 5312
rect 1900 5104 1940 5144
rect 1228 4936 1268 4976
rect 1036 4348 1076 4388
rect 1900 4852 1940 4892
rect 6412 4852 6452 4892
rect 2092 4684 2132 4724
rect 3688 4516 3728 4556
rect 3770 4516 3810 4556
rect 3852 4516 3892 4556
rect 3934 4516 3974 4556
rect 4016 4516 4056 4556
rect 1900 4348 1940 4388
rect 3148 4264 3188 4304
rect 2092 4180 2132 4220
rect 2476 3928 2516 3968
rect 1228 3088 1268 3128
rect 2092 3172 2132 3212
rect 2092 2248 2132 2288
rect 1804 1996 1844 2036
rect 1804 1828 1844 1868
rect 2188 1156 2228 1196
rect 1900 736 1940 776
rect 2188 736 2228 776
rect 3148 3760 3188 3800
rect 4928 3760 4968 3800
rect 5010 3760 5050 3800
rect 5092 3760 5132 3800
rect 5174 3760 5214 3800
rect 5256 3760 5296 3800
rect 6988 3760 7028 3800
rect 6412 3424 6452 3464
rect 3532 3256 3572 3296
rect 2956 2920 2996 2960
rect 3688 3004 3728 3044
rect 3770 3004 3810 3044
rect 3852 3004 3892 3044
rect 3934 3004 3974 3044
rect 4016 3004 4056 3044
rect 6220 3004 6260 3044
rect 6028 2836 6068 2876
rect 2572 1996 2612 2036
rect 2668 1828 2708 1868
rect 2860 2080 2900 2120
rect 5932 2668 5972 2708
rect 4928 2248 4968 2288
rect 5010 2248 5050 2288
rect 5092 2248 5132 2288
rect 5174 2248 5214 2288
rect 5256 2248 5296 2288
rect 5356 2080 5396 2120
rect 3916 1660 3956 1700
rect 3688 1492 3728 1532
rect 3770 1492 3810 1532
rect 3852 1492 3892 1532
rect 3934 1492 3974 1532
rect 4016 1492 4056 1532
rect 3340 1324 3380 1364
rect 4204 1828 4244 1868
rect 3532 1240 3572 1280
rect 4108 1240 4148 1280
rect 4300 1240 4340 1280
rect 3724 904 3764 944
rect 3916 820 3956 860
rect 5164 1828 5204 1868
rect 5452 1828 5492 1868
rect 4780 1660 4820 1700
rect 4684 1492 4724 1532
rect 4588 1408 4628 1448
rect 4492 1324 4532 1364
rect 4684 1324 4724 1364
rect 4396 232 4436 272
rect 4928 736 4968 776
rect 5010 736 5050 776
rect 5092 736 5132 776
rect 5174 736 5214 776
rect 5256 736 5296 776
rect 4876 568 4916 608
rect 4780 148 4820 188
rect 5068 484 5108 524
rect 5260 316 5300 356
rect 5836 1660 5876 1700
rect 5644 1240 5684 1280
rect 5836 1240 5876 1280
rect 6124 1408 6164 1448
rect 6892 2752 6932 2792
rect 6316 1408 6356 1448
rect 6796 1576 6836 1616
rect 6700 1324 6740 1364
rect 6604 904 6644 944
rect 6412 400 6452 440
rect 6892 568 6932 608
rect 9004 5104 9044 5144
rect 9580 5020 9620 5060
rect 9100 3928 9140 3968
rect 8044 3088 8084 3128
rect 7372 2584 7412 2624
rect 7276 1828 7316 1868
rect 7372 1660 7412 1700
rect 7180 1324 7220 1364
rect 7084 736 7124 776
rect 7660 820 7700 860
rect 7468 652 7508 692
rect 7564 568 7604 608
rect 7372 64 7412 104
rect 8332 2500 8372 2540
rect 8140 1828 8180 1868
rect 8044 988 8084 1028
rect 7852 904 7892 944
rect 8236 1660 8276 1700
rect 8236 1240 8276 1280
rect 8812 2332 8852 2372
rect 8524 820 8564 860
rect 8428 568 8468 608
rect 8716 1156 8756 1196
rect 8620 568 8660 608
rect 8908 400 8948 440
rect 10444 3256 10484 3296
rect 9676 2500 9716 2540
rect 9292 1996 9332 2036
rect 9676 1660 9716 1700
rect 9484 904 9524 944
rect 9868 1156 9908 1196
rect 10060 1492 10100 1532
rect 9964 484 10004 524
rect 9868 232 9908 272
rect 10156 904 10196 944
rect 10348 316 10388 356
rect 10252 148 10292 188
rect 10540 2920 10580 2960
rect 10732 8716 10772 8756
rect 12556 8800 12596 8840
rect 13036 8800 13076 8840
rect 13516 8800 13556 8840
rect 14092 8800 14132 8840
rect 14476 8800 14516 8840
rect 15436 8800 15476 8840
rect 16204 9472 16244 9512
rect 11596 8716 11636 8756
rect 10732 3172 10772 3212
rect 10636 2248 10676 2288
rect 10540 988 10580 1028
rect 11692 2752 11732 2792
rect 11212 1828 11252 1868
rect 11596 1240 11636 1280
rect 11404 1072 11444 1112
rect 11212 988 11252 1028
rect 10828 820 10868 860
rect 11020 820 11060 860
rect 11020 652 11060 692
rect 11404 904 11444 944
rect 11596 736 11636 776
rect 13612 8380 13652 8420
rect 13804 7792 13844 7832
rect 11788 2416 11828 2456
rect 11788 904 11828 944
rect 12076 1660 12116 1700
rect 11980 1408 12020 1448
rect 11884 148 11924 188
rect 12172 988 12212 1028
rect 13228 3760 13268 3800
rect 12364 2080 12404 2120
rect 12268 652 12308 692
rect 19564 10480 19604 10520
rect 18808 9052 18848 9092
rect 18890 9052 18930 9092
rect 18972 9052 19012 9092
rect 19054 9052 19094 9092
rect 19136 9052 19176 9092
rect 18220 8884 18260 8924
rect 16204 8548 16244 8588
rect 16012 6952 16052 6992
rect 15628 4180 15668 4220
rect 14284 3340 14324 3380
rect 15148 3004 15188 3044
rect 15532 2836 15572 2876
rect 13324 2080 13364 2120
rect 12844 1324 12884 1364
rect 12748 1156 12788 1196
rect 12556 820 12596 860
rect 12940 904 12980 944
rect 13132 1072 13172 1112
rect 13036 736 13076 776
rect 13612 1576 13652 1616
rect 13708 988 13748 1028
rect 13420 904 13460 944
rect 13516 568 13556 608
rect 13324 400 13364 440
rect 13996 1072 14036 1112
rect 14092 904 14132 944
rect 13804 820 13844 860
rect 13900 736 13940 776
rect 14284 820 14324 860
rect 14572 400 14612 440
rect 15244 1828 15284 1868
rect 15436 1660 15476 1700
rect 15820 5608 15860 5648
rect 15724 3256 15764 3296
rect 15916 1828 15956 1868
rect 15916 1660 15956 1700
rect 16204 6868 16244 6908
rect 16108 2668 16148 2708
rect 16108 1828 16148 1868
rect 16396 6364 16436 6404
rect 18412 8800 18452 8840
rect 20048 9808 20088 9848
rect 20130 9808 20170 9848
rect 20212 9808 20252 9848
rect 20294 9808 20334 9848
rect 20376 9808 20416 9848
rect 19180 8464 19220 8504
rect 17932 8128 17972 8168
rect 18124 8128 18164 8168
rect 18808 7540 18848 7580
rect 18890 7540 18930 7580
rect 18972 7540 19012 7580
rect 19054 7540 19094 7580
rect 19136 7540 19176 7580
rect 19372 7960 19412 8000
rect 18316 7120 18356 7160
rect 18316 6532 18356 6572
rect 19180 6448 19220 6488
rect 19276 6364 19316 6404
rect 16492 5860 16532 5900
rect 16396 5776 16436 5816
rect 16396 5020 16436 5060
rect 16300 3172 16340 3212
rect 16396 2500 16436 2540
rect 16588 5692 16628 5732
rect 16684 4852 16724 4892
rect 16876 3424 16916 3464
rect 16780 3088 16820 3128
rect 16780 2920 16820 2960
rect 16684 2500 16724 2540
rect 16684 232 16724 272
rect 17068 5104 17108 5144
rect 16972 2836 17012 2876
rect 17260 4264 17300 4304
rect 17452 3844 17492 3884
rect 17356 2668 17396 2708
rect 17068 2416 17108 2456
rect 16972 1240 17012 1280
rect 17260 2248 17300 2288
rect 17068 736 17108 776
rect 17164 400 17204 440
rect 17356 1492 17396 1532
rect 17356 568 17396 608
rect 17164 232 17204 272
rect 17740 1828 17780 1868
rect 17644 1408 17684 1448
rect 18808 6028 18848 6068
rect 18890 6028 18930 6068
rect 18972 6028 19012 6068
rect 19054 6028 19094 6068
rect 19136 6028 19176 6068
rect 19660 7456 19700 7496
rect 19852 7456 19892 7496
rect 19468 6448 19508 6488
rect 19468 5776 19508 5816
rect 19372 5440 19412 5480
rect 19180 5356 19220 5396
rect 18700 4936 18740 4976
rect 18808 4516 18848 4556
rect 18890 4516 18930 4556
rect 18972 4516 19012 4556
rect 19054 4516 19094 4556
rect 19136 4516 19176 4556
rect 19372 4432 19412 4472
rect 19180 4348 19220 4388
rect 18124 3340 18164 3380
rect 18028 2080 18068 2120
rect 17836 1324 17876 1364
rect 17548 1072 17588 1112
rect 17932 820 17972 860
rect 17548 736 17588 776
rect 17452 148 17492 188
rect 17740 652 17780 692
rect 18316 3256 18356 3296
rect 19276 3340 19316 3380
rect 19564 4180 19604 4220
rect 19756 4096 19796 4136
rect 18508 3172 18548 3212
rect 18988 3172 19028 3212
rect 18604 3088 18644 3128
rect 18808 3004 18848 3044
rect 18890 3004 18930 3044
rect 18972 3004 19012 3044
rect 19054 3004 19094 3044
rect 19136 3004 19176 3044
rect 19276 3004 19316 3044
rect 18892 2836 18932 2876
rect 18988 1828 19028 1868
rect 19180 1744 19220 1784
rect 18808 1492 18848 1532
rect 18890 1492 18930 1532
rect 18972 1492 19012 1532
rect 19054 1492 19094 1532
rect 19136 1492 19176 1532
rect 19084 1324 19124 1364
rect 19468 2752 19508 2792
rect 20620 9808 20660 9848
rect 20620 8632 20660 8672
rect 20524 8464 20564 8504
rect 21388 8464 21428 8504
rect 20048 8296 20088 8336
rect 20130 8296 20170 8336
rect 20212 8296 20252 8336
rect 20294 8296 20334 8336
rect 20376 8296 20416 8336
rect 21388 7960 21428 8000
rect 20048 6784 20088 6824
rect 20130 6784 20170 6824
rect 20212 6784 20252 6824
rect 20294 6784 20334 6824
rect 20376 6784 20416 6824
rect 20048 5272 20088 5312
rect 20130 5272 20170 5312
rect 20212 5272 20252 5312
rect 20294 5272 20334 5312
rect 20376 5272 20416 5312
rect 20048 3760 20088 3800
rect 20130 3760 20170 3800
rect 20212 3760 20252 3800
rect 20294 3760 20334 3800
rect 20376 3760 20416 3800
rect 19948 3004 19988 3044
rect 19372 1828 19412 1868
rect 19564 2416 19604 2456
rect 20048 2248 20088 2288
rect 20130 2248 20170 2288
rect 20212 2248 20252 2288
rect 20294 2248 20334 2288
rect 20376 2248 20416 2288
rect 19948 2080 19988 2120
rect 19756 1828 19796 1868
rect 20048 736 20088 776
rect 20130 736 20170 776
rect 20212 736 20252 776
rect 20294 736 20334 776
rect 20376 736 20416 776
<< metal3 >>
rect 0 10520 80 10540
rect 21424 10520 21504 10540
rect 0 10480 556 10520
rect 596 10480 605 10520
rect 19555 10480 19564 10520
rect 19604 10480 21504 10520
rect 0 10460 80 10480
rect 21424 10460 21504 10480
rect 0 10184 80 10204
rect 21283 10184 21341 10185
rect 21424 10184 21504 10204
rect 0 10144 2284 10184
rect 2324 10144 2333 10184
rect 21283 10144 21292 10184
rect 21332 10144 21504 10184
rect 0 10124 80 10144
rect 21283 10143 21341 10144
rect 21424 10124 21504 10144
rect 0 9848 80 9868
rect 21424 9848 21504 9868
rect 0 9808 1516 9848
rect 1556 9808 1565 9848
rect 4919 9808 4928 9848
rect 4968 9808 5010 9848
rect 5050 9808 5092 9848
rect 5132 9808 5174 9848
rect 5214 9808 5256 9848
rect 5296 9808 5305 9848
rect 20039 9808 20048 9848
rect 20088 9808 20130 9848
rect 20170 9808 20212 9848
rect 20252 9808 20294 9848
rect 20334 9808 20376 9848
rect 20416 9808 20425 9848
rect 20611 9808 20620 9848
rect 20660 9808 21504 9848
rect 0 9788 80 9808
rect 21424 9788 21504 9808
rect 7747 9640 7756 9680
rect 7796 9640 8812 9680
rect 8852 9640 8861 9680
rect 0 9512 80 9532
rect 21424 9512 21504 9532
rect 0 9472 1900 9512
rect 1940 9472 1949 9512
rect 16195 9472 16204 9512
rect 16244 9472 21504 9512
rect 0 9452 80 9472
rect 21424 9452 21504 9472
rect 0 9176 80 9196
rect 21424 9176 21504 9196
rect 0 9136 11212 9176
rect 11252 9136 11261 9176
rect 11395 9136 11404 9176
rect 11444 9136 21504 9176
rect 0 9116 80 9136
rect 21424 9116 21504 9136
rect 3679 9052 3688 9092
rect 3728 9052 3770 9092
rect 3810 9052 3852 9092
rect 3892 9052 3934 9092
rect 3974 9052 4016 9092
rect 4056 9052 4065 9092
rect 18799 9052 18808 9092
rect 18848 9052 18890 9092
rect 18930 9052 18972 9092
rect 19012 9052 19054 9092
rect 19094 9052 19136 9092
rect 19176 9052 19185 9092
rect 6280 8884 18220 8924
rect 18260 8884 18269 8924
rect 0 8840 80 8860
rect 6280 8840 6320 8884
rect 21424 8840 21504 8860
rect 0 8800 6320 8840
rect 6595 8800 6604 8840
rect 6644 8800 6653 8840
rect 8707 8800 8716 8840
rect 8756 8800 9388 8840
rect 9428 8800 9437 8840
rect 9667 8800 9676 8840
rect 9716 8800 10444 8840
rect 10484 8800 10493 8840
rect 12547 8800 12556 8840
rect 12596 8800 13036 8840
rect 13076 8800 13085 8840
rect 13507 8800 13516 8840
rect 13556 8800 14092 8840
rect 14132 8800 14141 8840
rect 14467 8800 14476 8840
rect 14516 8800 15436 8840
rect 15476 8800 15485 8840
rect 18403 8800 18412 8840
rect 18452 8800 21504 8840
rect 0 8780 80 8800
rect 6604 8756 6644 8800
rect 21424 8780 21504 8800
rect 2947 8716 2956 8756
rect 2996 8716 3820 8756
rect 3860 8716 3869 8756
rect 4867 8716 4876 8756
rect 4916 8716 5740 8756
rect 5780 8716 5789 8756
rect 6019 8716 6028 8756
rect 6068 8716 6644 8756
rect 6883 8716 6892 8756
rect 6932 8716 7852 8756
rect 7892 8716 7901 8756
rect 10723 8716 10732 8756
rect 10772 8716 11596 8756
rect 11636 8716 11645 8756
rect 1987 8632 1996 8672
rect 2036 8632 3436 8672
rect 3476 8632 3485 8672
rect 3907 8632 3916 8672
rect 3956 8632 20620 8672
rect 20660 8632 20669 8672
rect 2092 8548 16204 8588
rect 16244 8548 16253 8588
rect 0 8504 80 8524
rect 2092 8504 2132 8548
rect 2467 8504 2525 8505
rect 21424 8504 21504 8524
rect 0 8464 2036 8504
rect 2083 8464 2092 8504
rect 2132 8464 2141 8504
rect 2382 8464 2476 8504
rect 2516 8464 2525 8504
rect 19171 8464 19180 8504
rect 19220 8464 20524 8504
rect 20564 8464 20573 8504
rect 21379 8464 21388 8504
rect 21428 8464 21504 8504
rect 0 8444 80 8464
rect 1996 8420 2036 8464
rect 2467 8463 2525 8464
rect 21424 8444 21504 8464
rect 1996 8380 13612 8420
rect 13652 8380 13661 8420
rect 1699 8296 1708 8336
rect 1748 8296 3916 8336
rect 3956 8296 3965 8336
rect 4919 8296 4928 8336
rect 4968 8296 5010 8336
rect 5050 8296 5092 8336
rect 5132 8296 5174 8336
rect 5214 8296 5256 8336
rect 5296 8296 5305 8336
rect 20039 8296 20048 8336
rect 20088 8296 20130 8336
rect 20170 8296 20212 8336
rect 20252 8296 20294 8336
rect 20334 8296 20376 8336
rect 20416 8296 20425 8336
rect 0 8168 80 8188
rect 21424 8168 21504 8188
rect 0 8128 17932 8168
rect 17972 8128 17981 8168
rect 18115 8128 18124 8168
rect 18164 8128 21504 8168
rect 0 8108 80 8128
rect 21424 8108 21504 8128
rect 547 7960 556 8000
rect 596 7960 19372 8000
rect 19412 7960 19421 8000
rect 21292 7960 21388 8000
rect 21428 7960 21437 8000
rect 21292 7916 21332 7960
rect 2179 7876 2188 7916
rect 2228 7876 2237 7916
rect 4003 7876 4012 7916
rect 4052 7876 5164 7916
rect 5204 7876 5213 7916
rect 15100 7876 21332 7916
rect 0 7832 80 7852
rect 2188 7832 2228 7876
rect 15100 7832 15140 7876
rect 21424 7832 21504 7852
rect 0 7792 2228 7832
rect 13795 7792 13804 7832
rect 13844 7792 15140 7832
rect 18316 7792 21504 7832
rect 0 7772 80 7792
rect 2371 7708 2380 7748
rect 2420 7708 6320 7748
rect 6280 7664 6320 7708
rect 18316 7664 18356 7792
rect 21424 7772 21504 7792
rect 6280 7624 18356 7664
rect 3679 7540 3688 7580
rect 3728 7540 3770 7580
rect 3810 7540 3852 7580
rect 3892 7540 3934 7580
rect 3974 7540 4016 7580
rect 4056 7540 4065 7580
rect 5923 7540 5932 7580
rect 5972 7540 7372 7580
rect 7412 7540 7421 7580
rect 18799 7540 18808 7580
rect 18848 7540 18890 7580
rect 18930 7540 18972 7580
rect 19012 7540 19054 7580
rect 19094 7540 19136 7580
rect 19176 7540 19185 7580
rect 0 7496 80 7516
rect 21424 7496 21504 7516
rect 0 7456 19660 7496
rect 19700 7456 19709 7496
rect 19843 7456 19852 7496
rect 19892 7456 21504 7496
rect 0 7436 80 7456
rect 21424 7436 21504 7456
rect 0 7160 80 7180
rect 21424 7160 21504 7180
rect 0 7120 2572 7160
rect 2612 7120 2621 7160
rect 18307 7120 18316 7160
rect 18356 7120 21504 7160
rect 0 7100 80 7120
rect 21424 7100 21504 7120
rect 5155 6952 5164 6992
rect 5204 6952 16012 6992
rect 16052 6952 16061 6992
rect 4771 6868 4780 6908
rect 4820 6868 16204 6908
rect 16244 6868 16253 6908
rect 0 6824 80 6844
rect 21424 6824 21504 6844
rect 0 6784 2188 6824
rect 2228 6784 2237 6824
rect 4919 6784 4928 6824
rect 4968 6784 5010 6824
rect 5050 6784 5092 6824
rect 5132 6784 5174 6824
rect 5214 6784 5256 6824
rect 5296 6784 5305 6824
rect 20039 6784 20048 6824
rect 20088 6784 20130 6824
rect 20170 6784 20212 6824
rect 20252 6784 20294 6824
rect 20334 6784 20376 6824
rect 20416 6784 20425 6824
rect 21292 6784 21504 6824
rect 0 6764 80 6784
rect 2371 6700 2380 6740
rect 2420 6700 6320 6740
rect 6280 6656 6320 6700
rect 21292 6656 21332 6784
rect 21424 6764 21504 6784
rect 2755 6616 2764 6656
rect 2804 6616 2813 6656
rect 6280 6616 21332 6656
rect 2764 6572 2804 6616
rect 2764 6532 18316 6572
rect 18356 6532 18365 6572
rect 0 6488 80 6508
rect 21424 6488 21504 6508
rect 0 6448 19180 6488
rect 19220 6448 19229 6488
rect 19459 6448 19468 6488
rect 19508 6448 21504 6488
rect 0 6428 80 6448
rect 21424 6428 21504 6448
rect 16387 6364 16396 6404
rect 16436 6364 19276 6404
rect 19316 6364 19325 6404
rect 1987 6196 1996 6236
rect 2036 6196 6320 6236
rect 0 6152 80 6172
rect 6280 6152 6320 6196
rect 21424 6152 21504 6172
rect 0 6112 1804 6152
rect 1844 6112 1853 6152
rect 6280 6112 21504 6152
rect 0 6092 80 6112
rect 21424 6092 21504 6112
rect 3679 6028 3688 6068
rect 3728 6028 3770 6068
rect 3810 6028 3852 6068
rect 3892 6028 3934 6068
rect 3974 6028 4016 6068
rect 4056 6028 4065 6068
rect 18799 6028 18808 6068
rect 18848 6028 18890 6068
rect 18930 6028 18972 6068
rect 19012 6028 19054 6068
rect 19094 6028 19136 6068
rect 19176 6028 19185 6068
rect 7363 5860 7372 5900
rect 7412 5860 16492 5900
rect 16532 5860 16541 5900
rect 0 5816 80 5836
rect 21424 5816 21504 5836
rect 0 5776 16396 5816
rect 16436 5776 16445 5816
rect 19459 5776 19468 5816
rect 19508 5776 21504 5816
rect 0 5756 80 5776
rect 21424 5756 21504 5776
rect 6787 5692 6796 5732
rect 6836 5692 16588 5732
rect 16628 5692 16637 5732
rect 3523 5608 3532 5648
rect 3572 5608 15820 5648
rect 15860 5608 15869 5648
rect 2179 5524 2188 5564
rect 2228 5524 15140 5564
rect 0 5480 80 5500
rect 15100 5480 15140 5524
rect 21424 5480 21504 5500
rect 0 5440 6320 5480
rect 15100 5440 19316 5480
rect 19363 5440 19372 5480
rect 19412 5440 21504 5480
rect 0 5420 80 5440
rect 6280 5396 6320 5440
rect 6280 5356 19180 5396
rect 19220 5356 19229 5396
rect 4919 5272 4928 5312
rect 4968 5272 5010 5312
rect 5050 5272 5092 5312
rect 5132 5272 5174 5312
rect 5214 5272 5256 5312
rect 5296 5272 5305 5312
rect 0 5144 80 5164
rect 19276 5144 19316 5440
rect 21424 5420 21504 5440
rect 20039 5272 20048 5312
rect 20088 5272 20130 5312
rect 20170 5272 20212 5312
rect 20252 5272 20294 5312
rect 20334 5272 20376 5312
rect 20416 5272 20425 5312
rect 21424 5144 21504 5164
rect 0 5104 1900 5144
rect 1940 5104 1949 5144
rect 8995 5104 9004 5144
rect 9044 5104 17068 5144
rect 17108 5104 17117 5144
rect 19276 5104 21504 5144
rect 0 5084 80 5104
rect 21424 5084 21504 5104
rect 9571 5020 9580 5060
rect 9620 5020 16396 5060
rect 16436 5020 16445 5060
rect 1219 4936 1228 4976
rect 1268 4936 18700 4976
rect 18740 4936 18749 4976
rect 1891 4852 1900 4892
rect 1940 4852 1949 4892
rect 6403 4852 6412 4892
rect 6452 4852 16684 4892
rect 16724 4852 16733 4892
rect 0 4808 80 4828
rect 1900 4808 1940 4852
rect 21424 4808 21504 4828
rect 0 4768 1940 4808
rect 21292 4768 21504 4808
rect 0 4748 80 4768
rect 2083 4684 2092 4724
rect 2132 4684 6320 4724
rect 6280 4640 6320 4684
rect 21292 4640 21332 4768
rect 21424 4748 21504 4768
rect 6280 4600 21332 4640
rect 3679 4516 3688 4556
rect 3728 4516 3770 4556
rect 3810 4516 3852 4556
rect 3892 4516 3934 4556
rect 3974 4516 4016 4556
rect 4056 4516 4065 4556
rect 18799 4516 18808 4556
rect 18848 4516 18890 4556
rect 18930 4516 18972 4556
rect 19012 4516 19054 4556
rect 19094 4516 19136 4556
rect 19176 4516 19185 4556
rect 0 4472 80 4492
rect 21424 4472 21504 4492
rect 0 4432 6320 4472
rect 19363 4432 19372 4472
rect 19412 4432 21504 4472
rect 0 4412 80 4432
rect 6280 4388 6320 4432
rect 21424 4412 21504 4432
rect 1027 4348 1036 4388
rect 1076 4348 1900 4388
rect 1940 4348 1949 4388
rect 6280 4348 19180 4388
rect 19220 4348 19229 4388
rect 3139 4264 3148 4304
rect 3188 4264 17260 4304
rect 17300 4264 17309 4304
rect 2083 4180 2092 4220
rect 2132 4180 15628 4220
rect 15668 4180 15677 4220
rect 19555 4180 19564 4220
rect 19604 4180 19613 4220
rect 0 4136 80 4156
rect 19564 4136 19604 4180
rect 21424 4136 21504 4156
rect 0 4096 19604 4136
rect 19747 4096 19756 4136
rect 19796 4096 21504 4136
rect 0 4076 80 4096
rect 21424 4076 21504 4096
rect 2467 3928 2476 3968
rect 2516 3928 9100 3968
rect 9140 3928 9149 3968
rect 17443 3844 17452 3884
rect 17492 3844 20564 3884
rect 0 3800 80 3820
rect 20524 3800 20564 3844
rect 21424 3800 21504 3820
rect 0 3760 3148 3800
rect 3188 3760 3197 3800
rect 4919 3760 4928 3800
rect 4968 3760 5010 3800
rect 5050 3760 5092 3800
rect 5132 3760 5174 3800
rect 5214 3760 5256 3800
rect 5296 3760 5305 3800
rect 6979 3760 6988 3800
rect 7028 3760 13228 3800
rect 13268 3760 13277 3800
rect 20039 3760 20048 3800
rect 20088 3760 20130 3800
rect 20170 3760 20212 3800
rect 20252 3760 20294 3800
rect 20334 3760 20376 3800
rect 20416 3760 20425 3800
rect 20524 3760 21504 3800
rect 0 3740 80 3760
rect 21424 3740 21504 3760
rect 0 3464 80 3484
rect 21424 3464 21504 3484
rect 0 3424 6412 3464
rect 6452 3424 6461 3464
rect 16867 3424 16876 3464
rect 16916 3424 21504 3464
rect 0 3404 80 3424
rect 21424 3404 21504 3424
rect 19267 3380 19325 3381
rect 14275 3340 14284 3380
rect 14324 3340 18124 3380
rect 18164 3340 18173 3380
rect 19182 3340 19276 3380
rect 19316 3340 19325 3380
rect 19267 3339 19325 3340
rect 3523 3256 3532 3296
rect 3572 3256 10444 3296
rect 10484 3256 10493 3296
rect 15715 3256 15724 3296
rect 15764 3256 18316 3296
rect 18356 3256 18365 3296
rect 2083 3172 2092 3212
rect 2132 3172 10732 3212
rect 10772 3172 10781 3212
rect 16291 3172 16300 3212
rect 16340 3172 18508 3212
rect 18548 3172 18557 3212
rect 18979 3172 18988 3212
rect 19028 3172 19037 3212
rect 0 3128 80 3148
rect 18988 3128 19028 3172
rect 21424 3128 21504 3148
rect 0 3088 1228 3128
rect 1268 3088 1277 3128
rect 8035 3088 8044 3128
rect 8084 3088 16724 3128
rect 16771 3088 16780 3128
rect 16820 3088 18604 3128
rect 18644 3088 18653 3128
rect 18988 3088 21504 3128
rect 0 3068 80 3088
rect 3679 3004 3688 3044
rect 3728 3004 3770 3044
rect 3810 3004 3852 3044
rect 3892 3004 3934 3044
rect 3974 3004 4016 3044
rect 4056 3004 4065 3044
rect 6211 3004 6220 3044
rect 6260 3004 15148 3044
rect 15188 3004 15197 3044
rect 16684 2960 16724 3088
rect 21424 3068 21504 3088
rect 18799 3004 18808 3044
rect 18848 3004 18890 3044
rect 18930 3004 18972 3044
rect 19012 3004 19054 3044
rect 19094 3004 19136 3044
rect 19176 3004 19185 3044
rect 19267 3004 19276 3044
rect 19316 3004 19948 3044
rect 19988 3004 19997 3044
rect 2947 2920 2956 2960
rect 2996 2920 10540 2960
rect 10580 2920 10589 2960
rect 16684 2920 16780 2960
rect 16820 2920 16829 2960
rect 6019 2836 6028 2876
rect 6068 2836 15532 2876
rect 15572 2836 15581 2876
rect 16963 2836 16972 2876
rect 17012 2836 18892 2876
rect 18932 2836 18941 2876
rect 0 2792 80 2812
rect 1219 2792 1277 2793
rect 21424 2792 21504 2812
rect 0 2752 1228 2792
rect 1268 2752 1277 2792
rect 6883 2752 6892 2792
rect 6932 2752 11692 2792
rect 11732 2752 11741 2792
rect 19459 2752 19468 2792
rect 19508 2752 21504 2792
rect 0 2732 80 2752
rect 1219 2751 1277 2752
rect 21424 2732 21504 2752
rect 5923 2668 5932 2708
rect 5972 2668 16108 2708
rect 16148 2668 16157 2708
rect 17347 2668 17356 2708
rect 17396 2668 17405 2708
rect 17356 2624 17396 2668
rect 7363 2584 7372 2624
rect 7412 2584 17396 2624
rect 8323 2500 8332 2540
rect 8372 2500 9676 2540
rect 9716 2500 9725 2540
rect 16387 2500 16396 2540
rect 16436 2500 16684 2540
rect 16724 2500 16733 2540
rect 0 2456 80 2476
rect 1219 2456 1277 2457
rect 21424 2456 21504 2476
rect 0 2416 1228 2456
rect 1268 2416 1277 2456
rect 11779 2416 11788 2456
rect 11828 2416 17068 2456
rect 17108 2416 17117 2456
rect 19555 2416 19564 2456
rect 19604 2416 21504 2456
rect 0 2396 80 2416
rect 1219 2415 1277 2416
rect 21424 2396 21504 2416
rect 2092 2332 8812 2372
rect 8852 2332 8861 2372
rect 2092 2288 2132 2332
rect 2083 2248 2092 2288
rect 2132 2248 2141 2288
rect 4919 2248 4928 2288
rect 4968 2248 5010 2288
rect 5050 2248 5092 2288
rect 5132 2248 5174 2288
rect 5214 2248 5256 2288
rect 5296 2248 5305 2288
rect 10627 2248 10636 2288
rect 10676 2248 17260 2288
rect 17300 2248 17309 2288
rect 20039 2248 20048 2288
rect 20088 2248 20130 2288
rect 20170 2248 20212 2288
rect 20252 2248 20294 2288
rect 20334 2248 20376 2288
rect 20416 2248 20425 2288
rect 0 2120 80 2140
rect 1219 2120 1277 2121
rect 21424 2120 21504 2140
rect 0 2080 1228 2120
rect 1268 2080 1277 2120
rect 2851 2080 2860 2120
rect 2900 2080 2909 2120
rect 5347 2080 5356 2120
rect 5396 2080 12364 2120
rect 12404 2080 12413 2120
rect 13315 2080 13324 2120
rect 13364 2080 18028 2120
rect 18068 2080 18077 2120
rect 19939 2080 19948 2120
rect 19988 2080 21504 2120
rect 0 2060 80 2080
rect 1219 2079 1277 2080
rect 2860 2036 2900 2080
rect 21424 2060 21504 2080
rect 1795 1996 1804 2036
rect 1844 1996 2572 2036
rect 2612 1996 2621 2036
rect 2860 1996 9292 2036
rect 9332 1996 9341 2036
rect 17635 1952 17693 1953
rect 17635 1912 17644 1952
rect 17684 1912 19028 1952
rect 17635 1911 17693 1912
rect 16099 1868 16157 1869
rect 17731 1868 17789 1869
rect 18988 1868 19028 1912
rect 19363 1868 19421 1869
rect 19747 1868 19805 1869
rect 1795 1828 1804 1868
rect 1844 1828 2668 1868
rect 2708 1828 2717 1868
rect 4195 1828 4204 1868
rect 4244 1828 5164 1868
rect 5204 1828 5213 1868
rect 5443 1828 5452 1868
rect 5492 1828 7276 1868
rect 7316 1828 7325 1868
rect 8131 1828 8140 1868
rect 8180 1828 11212 1868
rect 11252 1828 11261 1868
rect 15235 1828 15244 1868
rect 15284 1828 15916 1868
rect 15956 1828 15965 1868
rect 16014 1828 16108 1868
rect 16148 1828 16157 1868
rect 17646 1828 17740 1868
rect 17780 1828 17789 1868
rect 18979 1828 18988 1868
rect 19028 1828 19037 1868
rect 19278 1828 19372 1868
rect 19412 1828 19421 1868
rect 19662 1828 19756 1868
rect 19796 1828 19805 1868
rect 16099 1827 16157 1828
rect 17731 1827 17789 1828
rect 19363 1827 19421 1828
rect 19747 1827 19805 1828
rect 0 1784 80 1804
rect 8707 1784 8765 1785
rect 21424 1784 21504 1804
rect 0 1744 8716 1784
rect 8756 1744 8765 1784
rect 19171 1744 19180 1784
rect 19220 1744 21504 1784
rect 0 1724 80 1744
rect 8707 1743 8765 1744
rect 21424 1724 21504 1744
rect 5827 1700 5885 1701
rect 11299 1700 11357 1701
rect 3907 1660 3916 1700
rect 3956 1660 4780 1700
rect 4820 1660 4829 1700
rect 5742 1660 5836 1700
rect 5876 1660 5885 1700
rect 5827 1659 5885 1660
rect 5932 1660 7372 1700
rect 7412 1660 7421 1700
rect 8227 1660 8236 1700
rect 8276 1660 9676 1700
rect 9716 1660 9725 1700
rect 11299 1660 11308 1700
rect 11348 1660 12076 1700
rect 12116 1660 12125 1700
rect 15427 1660 15436 1700
rect 15476 1660 15916 1700
rect 15956 1660 15965 1700
rect 5932 1616 5972 1660
rect 11299 1659 11357 1660
rect 3244 1576 5972 1616
rect 6787 1576 6796 1616
rect 6836 1576 13612 1616
rect 13652 1576 13661 1616
rect 0 1448 80 1468
rect 3244 1448 3284 1576
rect 13987 1532 14045 1533
rect 3679 1492 3688 1532
rect 3728 1492 3770 1532
rect 3810 1492 3852 1532
rect 3892 1492 3934 1532
rect 3974 1492 4016 1532
rect 4056 1492 4065 1532
rect 4675 1492 4684 1532
rect 4724 1492 10060 1532
rect 10100 1492 10109 1532
rect 13987 1492 13996 1532
rect 14036 1492 17356 1532
rect 17396 1492 17405 1532
rect 18799 1492 18808 1532
rect 18848 1492 18890 1532
rect 18930 1492 18972 1532
rect 19012 1492 19054 1532
rect 19094 1492 19136 1532
rect 19176 1492 19185 1532
rect 13987 1491 14045 1492
rect 21424 1448 21504 1468
rect 0 1408 3284 1448
rect 4579 1408 4588 1448
rect 4628 1408 6124 1448
rect 6164 1408 6173 1448
rect 6307 1408 6316 1448
rect 6356 1408 11980 1448
rect 12020 1408 12029 1448
rect 17635 1408 17644 1448
rect 17684 1408 21504 1448
rect 0 1388 80 1408
rect 21424 1388 21504 1408
rect 3331 1324 3340 1364
rect 3380 1324 4492 1364
rect 4532 1324 4541 1364
rect 4675 1324 4684 1364
rect 4724 1324 6700 1364
rect 6740 1324 6749 1364
rect 7171 1324 7180 1364
rect 7220 1324 12844 1364
rect 12884 1324 12893 1364
rect 17827 1324 17836 1364
rect 17876 1324 19084 1364
rect 19124 1324 19133 1364
rect 8035 1280 8093 1281
rect 13891 1280 13949 1281
rect 3523 1240 3532 1280
rect 3572 1240 4108 1280
rect 4148 1240 4157 1280
rect 4291 1240 4300 1280
rect 4340 1240 5644 1280
rect 5684 1240 5693 1280
rect 5827 1240 5836 1280
rect 5876 1240 8044 1280
rect 8084 1240 8093 1280
rect 8227 1240 8236 1280
rect 8276 1240 11596 1280
rect 11636 1240 11645 1280
rect 13891 1240 13900 1280
rect 13940 1240 16972 1280
rect 17012 1240 17021 1280
rect 8035 1239 8093 1240
rect 13891 1239 13949 1240
rect 2179 1156 2188 1196
rect 2228 1156 8716 1196
rect 8756 1156 8765 1196
rect 9859 1156 9868 1196
rect 9908 1156 12748 1196
rect 12788 1156 12797 1196
rect 0 1112 80 1132
rect 7459 1112 7517 1113
rect 13315 1112 13373 1113
rect 21424 1112 21504 1132
rect 0 1072 7468 1112
rect 7508 1072 7517 1112
rect 11395 1072 11404 1112
rect 11444 1072 13132 1112
rect 13172 1072 13181 1112
rect 13315 1072 13324 1112
rect 13364 1072 13996 1112
rect 14036 1072 14045 1112
rect 17539 1072 17548 1112
rect 17588 1072 21504 1112
rect 0 1052 80 1072
rect 7459 1071 7517 1072
rect 13315 1071 13373 1072
rect 21424 1052 21504 1072
rect 6280 988 8044 1028
rect 8084 988 8093 1028
rect 10531 988 10540 1028
rect 10580 988 11212 1028
rect 11252 988 11261 1028
rect 12163 988 12172 1028
rect 12212 988 13708 1028
rect 13748 988 13757 1028
rect 6280 944 6320 988
rect 6595 944 6653 945
rect 3715 904 3724 944
rect 3764 904 6320 944
rect 6510 904 6604 944
rect 6644 904 6653 944
rect 7843 904 7852 944
rect 7892 904 9484 944
rect 9524 904 9533 944
rect 10147 904 10156 944
rect 10196 904 11404 944
rect 11444 904 11453 944
rect 11779 904 11788 944
rect 11828 904 12940 944
rect 12980 904 12989 944
rect 13411 904 13420 944
rect 13460 904 14092 944
rect 14132 904 14141 944
rect 6595 903 6653 904
rect 3907 820 3916 860
rect 3956 820 7660 860
rect 7700 820 7709 860
rect 8515 820 8524 860
rect 8564 820 10828 860
rect 10868 820 10877 860
rect 11011 820 11020 860
rect 11060 820 12556 860
rect 12596 820 12605 860
rect 13795 820 13804 860
rect 13844 820 14284 860
rect 14324 820 14333 860
rect 17923 820 17932 860
rect 17972 820 20564 860
rect 0 776 80 796
rect 1699 776 1757 777
rect 20524 776 20564 820
rect 21424 776 21504 796
rect 0 736 1708 776
rect 1748 736 1757 776
rect 1891 736 1900 776
rect 1940 736 2188 776
rect 2228 736 2237 776
rect 4919 736 4928 776
rect 4968 736 5010 776
rect 5050 736 5092 776
rect 5132 736 5174 776
rect 5214 736 5256 776
rect 5296 736 5305 776
rect 7075 736 7084 776
rect 7124 736 11596 776
rect 11636 736 11645 776
rect 13027 736 13036 776
rect 13076 736 13900 776
rect 13940 736 13949 776
rect 17059 736 17068 776
rect 17108 736 17548 776
rect 17588 736 17597 776
rect 20039 736 20048 776
rect 20088 736 20130 776
rect 20170 736 20212 776
rect 20252 736 20294 776
rect 20334 736 20376 776
rect 20416 736 20425 776
rect 20524 736 21504 776
rect 0 716 80 736
rect 1699 735 1757 736
rect 21424 716 21504 736
rect 7459 652 7468 692
rect 7508 652 11020 692
rect 11060 652 11069 692
rect 12259 652 12268 692
rect 12308 652 17740 692
rect 17780 652 17789 692
rect 15331 608 15389 609
rect 4867 568 4876 608
rect 4916 568 6892 608
rect 6932 568 6941 608
rect 7555 568 7564 608
rect 7604 568 8428 608
rect 8468 568 8477 608
rect 8611 568 8620 608
rect 8660 568 13516 608
rect 13556 568 13565 608
rect 15331 568 15340 608
rect 15380 568 17356 608
rect 17396 568 17405 608
rect 15331 567 15389 568
rect 5059 484 5068 524
rect 5108 484 9964 524
rect 10004 484 10013 524
rect 0 440 80 460
rect 5347 440 5405 441
rect 6403 440 6461 441
rect 13795 440 13853 441
rect 21424 440 21504 460
rect 0 400 5356 440
rect 5396 400 5405 440
rect 6318 400 6412 440
rect 6452 400 6461 440
rect 8899 400 8908 440
rect 8948 400 13324 440
rect 13364 400 13373 440
rect 13795 400 13804 440
rect 13844 400 14572 440
rect 14612 400 14621 440
rect 17155 400 17164 440
rect 17204 400 21504 440
rect 0 380 80 400
rect 5347 399 5405 400
rect 6403 399 6461 400
rect 13795 399 13853 400
rect 21424 380 21504 400
rect 5251 316 5260 356
rect 5300 316 10348 356
rect 10388 316 10397 356
rect 4387 232 4396 272
rect 4436 232 9868 272
rect 9908 232 9917 272
rect 16675 232 16684 272
rect 16724 232 17164 272
rect 17204 232 17213 272
rect 4771 148 4780 188
rect 4820 148 10252 188
rect 10292 148 10301 188
rect 11875 148 11884 188
rect 11924 148 11933 188
rect 17443 148 17452 188
rect 17492 148 17501 188
rect 0 104 80 124
rect 3235 104 3293 105
rect 11884 104 11924 148
rect 0 64 3244 104
rect 3284 64 3293 104
rect 7363 64 7372 104
rect 7412 64 11924 104
rect 17452 104 17492 148
rect 21424 104 21504 124
rect 17452 64 21504 104
rect 0 44 80 64
rect 3235 63 3293 64
rect 21424 44 21504 64
<< via3 >>
rect 21292 10144 21332 10184
rect 4928 9808 4968 9848
rect 5010 9808 5050 9848
rect 5092 9808 5132 9848
rect 5174 9808 5214 9848
rect 5256 9808 5296 9848
rect 20048 9808 20088 9848
rect 20130 9808 20170 9848
rect 20212 9808 20252 9848
rect 20294 9808 20334 9848
rect 20376 9808 20416 9848
rect 3688 9052 3728 9092
rect 3770 9052 3810 9092
rect 3852 9052 3892 9092
rect 3934 9052 3974 9092
rect 4016 9052 4056 9092
rect 18808 9052 18848 9092
rect 18890 9052 18930 9092
rect 18972 9052 19012 9092
rect 19054 9052 19094 9092
rect 19136 9052 19176 9092
rect 2476 8464 2516 8504
rect 4928 8296 4968 8336
rect 5010 8296 5050 8336
rect 5092 8296 5132 8336
rect 5174 8296 5214 8336
rect 5256 8296 5296 8336
rect 20048 8296 20088 8336
rect 20130 8296 20170 8336
rect 20212 8296 20252 8336
rect 20294 8296 20334 8336
rect 20376 8296 20416 8336
rect 3688 7540 3728 7580
rect 3770 7540 3810 7580
rect 3852 7540 3892 7580
rect 3934 7540 3974 7580
rect 4016 7540 4056 7580
rect 18808 7540 18848 7580
rect 18890 7540 18930 7580
rect 18972 7540 19012 7580
rect 19054 7540 19094 7580
rect 19136 7540 19176 7580
rect 4928 6784 4968 6824
rect 5010 6784 5050 6824
rect 5092 6784 5132 6824
rect 5174 6784 5214 6824
rect 5256 6784 5296 6824
rect 20048 6784 20088 6824
rect 20130 6784 20170 6824
rect 20212 6784 20252 6824
rect 20294 6784 20334 6824
rect 20376 6784 20416 6824
rect 3688 6028 3728 6068
rect 3770 6028 3810 6068
rect 3852 6028 3892 6068
rect 3934 6028 3974 6068
rect 4016 6028 4056 6068
rect 18808 6028 18848 6068
rect 18890 6028 18930 6068
rect 18972 6028 19012 6068
rect 19054 6028 19094 6068
rect 19136 6028 19176 6068
rect 4928 5272 4968 5312
rect 5010 5272 5050 5312
rect 5092 5272 5132 5312
rect 5174 5272 5214 5312
rect 5256 5272 5296 5312
rect 20048 5272 20088 5312
rect 20130 5272 20170 5312
rect 20212 5272 20252 5312
rect 20294 5272 20334 5312
rect 20376 5272 20416 5312
rect 3688 4516 3728 4556
rect 3770 4516 3810 4556
rect 3852 4516 3892 4556
rect 3934 4516 3974 4556
rect 4016 4516 4056 4556
rect 18808 4516 18848 4556
rect 18890 4516 18930 4556
rect 18972 4516 19012 4556
rect 19054 4516 19094 4556
rect 19136 4516 19176 4556
rect 4928 3760 4968 3800
rect 5010 3760 5050 3800
rect 5092 3760 5132 3800
rect 5174 3760 5214 3800
rect 5256 3760 5296 3800
rect 20048 3760 20088 3800
rect 20130 3760 20170 3800
rect 20212 3760 20252 3800
rect 20294 3760 20334 3800
rect 20376 3760 20416 3800
rect 19276 3340 19316 3380
rect 3688 3004 3728 3044
rect 3770 3004 3810 3044
rect 3852 3004 3892 3044
rect 3934 3004 3974 3044
rect 4016 3004 4056 3044
rect 18808 3004 18848 3044
rect 18890 3004 18930 3044
rect 18972 3004 19012 3044
rect 19054 3004 19094 3044
rect 19136 3004 19176 3044
rect 1228 2752 1268 2792
rect 1228 2416 1268 2456
rect 4928 2248 4968 2288
rect 5010 2248 5050 2288
rect 5092 2248 5132 2288
rect 5174 2248 5214 2288
rect 5256 2248 5296 2288
rect 20048 2248 20088 2288
rect 20130 2248 20170 2288
rect 20212 2248 20252 2288
rect 20294 2248 20334 2288
rect 20376 2248 20416 2288
rect 1228 2080 1268 2120
rect 17644 1912 17684 1952
rect 16108 1828 16148 1868
rect 17740 1828 17780 1868
rect 19372 1828 19412 1868
rect 19756 1828 19796 1868
rect 8716 1744 8756 1784
rect 5836 1660 5876 1700
rect 11308 1660 11348 1700
rect 3688 1492 3728 1532
rect 3770 1492 3810 1532
rect 3852 1492 3892 1532
rect 3934 1492 3974 1532
rect 4016 1492 4056 1532
rect 13996 1492 14036 1532
rect 18808 1492 18848 1532
rect 18890 1492 18930 1532
rect 18972 1492 19012 1532
rect 19054 1492 19094 1532
rect 19136 1492 19176 1532
rect 8044 1240 8084 1280
rect 13900 1240 13940 1280
rect 7468 1072 7508 1112
rect 13324 1072 13364 1112
rect 6604 904 6644 944
rect 1708 736 1748 776
rect 4928 736 4968 776
rect 5010 736 5050 776
rect 5092 736 5132 776
rect 5174 736 5214 776
rect 5256 736 5296 776
rect 20048 736 20088 776
rect 20130 736 20170 776
rect 20212 736 20252 776
rect 20294 736 20334 776
rect 20376 736 20416 776
rect 15340 568 15380 608
rect 5356 400 5396 440
rect 6412 400 6452 440
rect 13804 400 13844 440
rect 3244 64 3284 104
<< metal4 >>
rect 21292 10184 21332 10193
rect 4928 9848 5296 9857
rect 4968 9808 5010 9848
rect 5050 9808 5092 9848
rect 5132 9808 5174 9848
rect 5214 9808 5256 9848
rect 4928 9799 5296 9808
rect 20048 9848 20416 9857
rect 20088 9808 20130 9848
rect 20170 9808 20212 9848
rect 20252 9808 20294 9848
rect 20334 9808 20376 9848
rect 20048 9799 20416 9808
rect 3688 9092 4056 9101
rect 3728 9052 3770 9092
rect 3810 9052 3852 9092
rect 3892 9052 3934 9092
rect 3974 9052 4016 9092
rect 3688 9043 4056 9052
rect 18808 9092 19176 9101
rect 18848 9052 18890 9092
rect 18930 9052 18972 9092
rect 19012 9052 19054 9092
rect 19094 9052 19136 9092
rect 18808 9043 19176 9052
rect 21292 8513 21332 10144
rect 2475 8504 2517 8513
rect 2475 8464 2476 8504
rect 2516 8464 2517 8504
rect 2475 8455 2517 8464
rect 21291 8504 21333 8513
rect 21291 8464 21292 8504
rect 21332 8464 21333 8504
rect 21291 8455 21333 8464
rect 2476 8370 2516 8455
rect 4928 8336 5296 8345
rect 4968 8296 5010 8336
rect 5050 8296 5092 8336
rect 5132 8296 5174 8336
rect 5214 8296 5256 8336
rect 4928 8287 5296 8296
rect 20048 8336 20416 8345
rect 20088 8296 20130 8336
rect 20170 8296 20212 8336
rect 20252 8296 20294 8336
rect 20334 8296 20376 8336
rect 20048 8287 20416 8296
rect 3688 7580 4056 7589
rect 3728 7540 3770 7580
rect 3810 7540 3852 7580
rect 3892 7540 3934 7580
rect 3974 7540 4016 7580
rect 3688 7531 4056 7540
rect 18808 7580 19176 7589
rect 18848 7540 18890 7580
rect 18930 7540 18972 7580
rect 19012 7540 19054 7580
rect 19094 7540 19136 7580
rect 18808 7531 19176 7540
rect 4928 6824 5296 6833
rect 4968 6784 5010 6824
rect 5050 6784 5092 6824
rect 5132 6784 5174 6824
rect 5214 6784 5256 6824
rect 4928 6775 5296 6784
rect 20048 6824 20416 6833
rect 20088 6784 20130 6824
rect 20170 6784 20212 6824
rect 20252 6784 20294 6824
rect 20334 6784 20376 6824
rect 20048 6775 20416 6784
rect 3688 6068 4056 6077
rect 3728 6028 3770 6068
rect 3810 6028 3852 6068
rect 3892 6028 3934 6068
rect 3974 6028 4016 6068
rect 3688 6019 4056 6028
rect 18808 6068 19176 6077
rect 18848 6028 18890 6068
rect 18930 6028 18972 6068
rect 19012 6028 19054 6068
rect 19094 6028 19136 6068
rect 18808 6019 19176 6028
rect 4928 5312 5296 5321
rect 4968 5272 5010 5312
rect 5050 5272 5092 5312
rect 5132 5272 5174 5312
rect 5214 5272 5256 5312
rect 4928 5263 5296 5272
rect 20048 5312 20416 5321
rect 20088 5272 20130 5312
rect 20170 5272 20212 5312
rect 20252 5272 20294 5312
rect 20334 5272 20376 5312
rect 20048 5263 20416 5272
rect 3688 4556 4056 4565
rect 3728 4516 3770 4556
rect 3810 4516 3852 4556
rect 3892 4516 3934 4556
rect 3974 4516 4016 4556
rect 3688 4507 4056 4516
rect 18808 4556 19176 4565
rect 18848 4516 18890 4556
rect 18930 4516 18972 4556
rect 19012 4516 19054 4556
rect 19094 4516 19136 4556
rect 18808 4507 19176 4516
rect 4928 3800 5296 3809
rect 4968 3760 5010 3800
rect 5050 3760 5092 3800
rect 5132 3760 5174 3800
rect 5214 3760 5256 3800
rect 4928 3751 5296 3760
rect 20048 3800 20416 3809
rect 20088 3760 20130 3800
rect 20170 3760 20212 3800
rect 20252 3760 20294 3800
rect 20334 3760 20376 3800
rect 20048 3751 20416 3760
rect 19276 3380 19316 3389
rect 3688 3044 4056 3053
rect 3728 3004 3770 3044
rect 3810 3004 3852 3044
rect 3892 3004 3934 3044
rect 3974 3004 4016 3044
rect 3688 2995 4056 3004
rect 18808 3044 19176 3053
rect 18848 3004 18890 3044
rect 18930 3004 18972 3044
rect 19012 3004 19054 3044
rect 19094 3004 19136 3044
rect 18808 2995 19176 3004
rect 19276 2801 19316 3340
rect 1227 2792 1269 2801
rect 1227 2752 1228 2792
rect 1268 2752 1269 2792
rect 1227 2743 1269 2752
rect 19275 2792 19317 2801
rect 19275 2752 19276 2792
rect 19316 2752 19317 2792
rect 19275 2743 19317 2752
rect 1228 2658 1268 2743
rect 1227 2456 1269 2465
rect 1227 2416 1228 2456
rect 1268 2416 1269 2456
rect 1227 2407 1269 2416
rect 19371 2456 19413 2465
rect 19371 2416 19372 2456
rect 19412 2416 19413 2456
rect 19371 2407 19413 2416
rect 1228 2322 1268 2407
rect 4928 2288 5296 2297
rect 4968 2248 5010 2288
rect 5050 2248 5092 2288
rect 5132 2248 5174 2288
rect 5214 2248 5256 2288
rect 4928 2239 5296 2248
rect 1227 2120 1269 2129
rect 1227 2080 1228 2120
rect 1268 2080 1269 2120
rect 1227 2071 1269 2080
rect 1228 1986 1268 2071
rect 8715 1952 8757 1961
rect 8715 1912 8716 1952
rect 8756 1912 8757 1952
rect 8715 1903 8757 1912
rect 17643 1952 17685 1961
rect 17643 1912 17644 1952
rect 17684 1912 17685 1952
rect 17643 1903 17685 1912
rect 8043 1868 8085 1877
rect 8043 1828 8044 1868
rect 8084 1828 8085 1868
rect 8043 1819 8085 1828
rect 1707 1784 1749 1793
rect 1707 1744 1708 1784
rect 1748 1744 1749 1784
rect 1707 1735 1749 1744
rect 1708 776 1748 1735
rect 5835 1700 5877 1709
rect 5835 1660 5836 1700
rect 5876 1660 5877 1700
rect 5835 1651 5877 1660
rect 5836 1566 5876 1651
rect 3688 1532 4056 1541
rect 3728 1492 3770 1532
rect 3810 1492 3852 1532
rect 3892 1492 3934 1532
rect 3974 1492 4016 1532
rect 3688 1483 4056 1492
rect 5355 1280 5397 1289
rect 5355 1240 5356 1280
rect 5396 1240 5397 1280
rect 5355 1231 5397 1240
rect 8044 1280 8084 1819
rect 8716 1784 8756 1903
rect 16107 1868 16149 1877
rect 16107 1828 16108 1868
rect 16148 1828 16149 1868
rect 16107 1819 16149 1828
rect 8716 1735 8756 1744
rect 16108 1734 16148 1819
rect 17644 1818 17684 1903
rect 17739 1868 17781 1877
rect 17739 1828 17740 1868
rect 17780 1828 17781 1868
rect 17739 1819 17781 1828
rect 19372 1868 19412 2407
rect 20048 2288 20416 2297
rect 20088 2248 20130 2288
rect 20170 2248 20212 2288
rect 20252 2248 20294 2288
rect 20334 2248 20376 2288
rect 20048 2239 20416 2248
rect 19755 2120 19797 2129
rect 19755 2080 19756 2120
rect 19796 2080 19797 2120
rect 19755 2071 19797 2080
rect 19372 1819 19412 1828
rect 19756 1868 19796 2071
rect 19756 1819 19796 1828
rect 17740 1734 17780 1819
rect 11307 1700 11349 1709
rect 11307 1660 11308 1700
rect 11348 1660 11349 1700
rect 11307 1651 11349 1660
rect 11308 1566 11348 1651
rect 13996 1532 14036 1541
rect 8044 1231 8084 1240
rect 13899 1280 13941 1289
rect 13899 1240 13900 1280
rect 13940 1240 13941 1280
rect 13899 1231 13941 1240
rect 3243 1196 3285 1205
rect 3243 1156 3244 1196
rect 3284 1156 3285 1196
rect 3243 1147 3285 1156
rect 1708 727 1748 736
rect 3244 104 3284 1147
rect 4928 776 5296 785
rect 4968 736 5010 776
rect 5050 736 5092 776
rect 5132 736 5174 776
rect 5214 736 5256 776
rect 4928 727 5296 736
rect 5356 440 5396 1231
rect 13900 1146 13940 1231
rect 13996 1205 14036 1492
rect 18808 1532 19176 1541
rect 18848 1492 18890 1532
rect 18930 1492 18972 1532
rect 19012 1492 19054 1532
rect 19094 1492 19136 1532
rect 18808 1483 19176 1492
rect 13995 1196 14037 1205
rect 13995 1156 13996 1196
rect 14036 1156 14037 1196
rect 13995 1147 14037 1156
rect 6603 1112 6645 1121
rect 6603 1072 6604 1112
rect 6644 1072 6645 1112
rect 6603 1063 6645 1072
rect 7468 1112 7508 1121
rect 6604 944 6644 1063
rect 6604 895 6644 904
rect 7468 617 7508 1072
rect 13323 1112 13365 1121
rect 13323 1072 13324 1112
rect 13364 1072 13365 1112
rect 13323 1063 13365 1072
rect 13324 978 13364 1063
rect 20048 776 20416 785
rect 20088 736 20130 776
rect 20170 736 20212 776
rect 20252 736 20294 776
rect 20334 736 20376 776
rect 20048 727 20416 736
rect 7467 608 7509 617
rect 7467 568 7468 608
rect 7508 568 7509 608
rect 7467 559 7509 568
rect 15339 608 15381 617
rect 15339 568 15340 608
rect 15380 568 15381 608
rect 15339 559 15381 568
rect 15340 474 15380 559
rect 5356 391 5396 400
rect 6411 440 6453 449
rect 6411 400 6412 440
rect 6452 400 6453 440
rect 6411 391 6453 400
rect 13803 440 13845 449
rect 13803 400 13804 440
rect 13844 400 13845 440
rect 13803 391 13845 400
rect 6412 306 6452 391
rect 13804 306 13844 391
rect 3244 55 3284 64
<< via4 >>
rect 4928 9808 4968 9848
rect 5010 9808 5050 9848
rect 5092 9808 5132 9848
rect 5174 9808 5214 9848
rect 5256 9808 5296 9848
rect 20048 9808 20088 9848
rect 20130 9808 20170 9848
rect 20212 9808 20252 9848
rect 20294 9808 20334 9848
rect 20376 9808 20416 9848
rect 3688 9052 3728 9092
rect 3770 9052 3810 9092
rect 3852 9052 3892 9092
rect 3934 9052 3974 9092
rect 4016 9052 4056 9092
rect 18808 9052 18848 9092
rect 18890 9052 18930 9092
rect 18972 9052 19012 9092
rect 19054 9052 19094 9092
rect 19136 9052 19176 9092
rect 2476 8464 2516 8504
rect 21292 8464 21332 8504
rect 4928 8296 4968 8336
rect 5010 8296 5050 8336
rect 5092 8296 5132 8336
rect 5174 8296 5214 8336
rect 5256 8296 5296 8336
rect 20048 8296 20088 8336
rect 20130 8296 20170 8336
rect 20212 8296 20252 8336
rect 20294 8296 20334 8336
rect 20376 8296 20416 8336
rect 3688 7540 3728 7580
rect 3770 7540 3810 7580
rect 3852 7540 3892 7580
rect 3934 7540 3974 7580
rect 4016 7540 4056 7580
rect 18808 7540 18848 7580
rect 18890 7540 18930 7580
rect 18972 7540 19012 7580
rect 19054 7540 19094 7580
rect 19136 7540 19176 7580
rect 4928 6784 4968 6824
rect 5010 6784 5050 6824
rect 5092 6784 5132 6824
rect 5174 6784 5214 6824
rect 5256 6784 5296 6824
rect 20048 6784 20088 6824
rect 20130 6784 20170 6824
rect 20212 6784 20252 6824
rect 20294 6784 20334 6824
rect 20376 6784 20416 6824
rect 3688 6028 3728 6068
rect 3770 6028 3810 6068
rect 3852 6028 3892 6068
rect 3934 6028 3974 6068
rect 4016 6028 4056 6068
rect 18808 6028 18848 6068
rect 18890 6028 18930 6068
rect 18972 6028 19012 6068
rect 19054 6028 19094 6068
rect 19136 6028 19176 6068
rect 4928 5272 4968 5312
rect 5010 5272 5050 5312
rect 5092 5272 5132 5312
rect 5174 5272 5214 5312
rect 5256 5272 5296 5312
rect 20048 5272 20088 5312
rect 20130 5272 20170 5312
rect 20212 5272 20252 5312
rect 20294 5272 20334 5312
rect 20376 5272 20416 5312
rect 3688 4516 3728 4556
rect 3770 4516 3810 4556
rect 3852 4516 3892 4556
rect 3934 4516 3974 4556
rect 4016 4516 4056 4556
rect 18808 4516 18848 4556
rect 18890 4516 18930 4556
rect 18972 4516 19012 4556
rect 19054 4516 19094 4556
rect 19136 4516 19176 4556
rect 4928 3760 4968 3800
rect 5010 3760 5050 3800
rect 5092 3760 5132 3800
rect 5174 3760 5214 3800
rect 5256 3760 5296 3800
rect 20048 3760 20088 3800
rect 20130 3760 20170 3800
rect 20212 3760 20252 3800
rect 20294 3760 20334 3800
rect 20376 3760 20416 3800
rect 3688 3004 3728 3044
rect 3770 3004 3810 3044
rect 3852 3004 3892 3044
rect 3934 3004 3974 3044
rect 4016 3004 4056 3044
rect 18808 3004 18848 3044
rect 18890 3004 18930 3044
rect 18972 3004 19012 3044
rect 19054 3004 19094 3044
rect 19136 3004 19176 3044
rect 1228 2752 1268 2792
rect 19276 2752 19316 2792
rect 1228 2416 1268 2456
rect 19372 2416 19412 2456
rect 4928 2248 4968 2288
rect 5010 2248 5050 2288
rect 5092 2248 5132 2288
rect 5174 2248 5214 2288
rect 5256 2248 5296 2288
rect 1228 2080 1268 2120
rect 8716 1912 8756 1952
rect 17644 1912 17684 1952
rect 8044 1828 8084 1868
rect 1708 1744 1748 1784
rect 5836 1660 5876 1700
rect 3688 1492 3728 1532
rect 3770 1492 3810 1532
rect 3852 1492 3892 1532
rect 3934 1492 3974 1532
rect 4016 1492 4056 1532
rect 5356 1240 5396 1280
rect 16108 1828 16148 1868
rect 17740 1828 17780 1868
rect 20048 2248 20088 2288
rect 20130 2248 20170 2288
rect 20212 2248 20252 2288
rect 20294 2248 20334 2288
rect 20376 2248 20416 2288
rect 19756 2080 19796 2120
rect 11308 1660 11348 1700
rect 13900 1240 13940 1280
rect 3244 1156 3284 1196
rect 4928 736 4968 776
rect 5010 736 5050 776
rect 5092 736 5132 776
rect 5174 736 5214 776
rect 5256 736 5296 776
rect 18808 1492 18848 1532
rect 18890 1492 18930 1532
rect 18972 1492 19012 1532
rect 19054 1492 19094 1532
rect 19136 1492 19176 1532
rect 13996 1156 14036 1196
rect 6604 1072 6644 1112
rect 13324 1072 13364 1112
rect 20048 736 20088 776
rect 20130 736 20170 776
rect 20212 736 20252 776
rect 20294 736 20334 776
rect 20376 736 20416 776
rect 7468 568 7508 608
rect 15340 568 15380 608
rect 6412 400 6452 440
rect 13804 400 13844 440
<< metal5 >>
rect 4919 9871 5305 9890
rect 4919 9848 4985 9871
rect 5071 9848 5153 9871
rect 5239 9848 5305 9871
rect 4919 9808 4928 9848
rect 4968 9808 4985 9848
rect 5071 9808 5092 9848
rect 5132 9808 5153 9848
rect 5239 9808 5256 9848
rect 5296 9808 5305 9848
rect 4919 9785 4985 9808
rect 5071 9785 5153 9808
rect 5239 9785 5305 9808
rect 4919 9766 5305 9785
rect 20039 9871 20425 9890
rect 20039 9848 20105 9871
rect 20191 9848 20273 9871
rect 20359 9848 20425 9871
rect 20039 9808 20048 9848
rect 20088 9808 20105 9848
rect 20191 9808 20212 9848
rect 20252 9808 20273 9848
rect 20359 9808 20376 9848
rect 20416 9808 20425 9848
rect 20039 9785 20105 9808
rect 20191 9785 20273 9808
rect 20359 9785 20425 9808
rect 20039 9766 20425 9785
rect 3679 9115 4065 9134
rect 3679 9092 3745 9115
rect 3831 9092 3913 9115
rect 3999 9092 4065 9115
rect 3679 9052 3688 9092
rect 3728 9052 3745 9092
rect 3831 9052 3852 9092
rect 3892 9052 3913 9092
rect 3999 9052 4016 9092
rect 4056 9052 4065 9092
rect 3679 9029 3745 9052
rect 3831 9029 3913 9052
rect 3999 9029 4065 9052
rect 3679 9010 4065 9029
rect 18799 9115 19185 9134
rect 18799 9092 18865 9115
rect 18951 9092 19033 9115
rect 19119 9092 19185 9115
rect 18799 9052 18808 9092
rect 18848 9052 18865 9092
rect 18951 9052 18972 9092
rect 19012 9052 19033 9092
rect 19119 9052 19136 9092
rect 19176 9052 19185 9092
rect 18799 9029 18865 9052
rect 18951 9029 19033 9052
rect 19119 9029 19185 9052
rect 18799 9010 19185 9029
rect 2467 8464 2476 8504
rect 2516 8464 21292 8504
rect 21332 8464 21341 8504
rect 4919 8359 5305 8378
rect 4919 8336 4985 8359
rect 5071 8336 5153 8359
rect 5239 8336 5305 8359
rect 4919 8296 4928 8336
rect 4968 8296 4985 8336
rect 5071 8296 5092 8336
rect 5132 8296 5153 8336
rect 5239 8296 5256 8336
rect 5296 8296 5305 8336
rect 4919 8273 4985 8296
rect 5071 8273 5153 8296
rect 5239 8273 5305 8296
rect 4919 8254 5305 8273
rect 20039 8359 20425 8378
rect 20039 8336 20105 8359
rect 20191 8336 20273 8359
rect 20359 8336 20425 8359
rect 20039 8296 20048 8336
rect 20088 8296 20105 8336
rect 20191 8296 20212 8336
rect 20252 8296 20273 8336
rect 20359 8296 20376 8336
rect 20416 8296 20425 8336
rect 20039 8273 20105 8296
rect 20191 8273 20273 8296
rect 20359 8273 20425 8296
rect 20039 8254 20425 8273
rect 3679 7603 4065 7622
rect 3679 7580 3745 7603
rect 3831 7580 3913 7603
rect 3999 7580 4065 7603
rect 3679 7540 3688 7580
rect 3728 7540 3745 7580
rect 3831 7540 3852 7580
rect 3892 7540 3913 7580
rect 3999 7540 4016 7580
rect 4056 7540 4065 7580
rect 3679 7517 3745 7540
rect 3831 7517 3913 7540
rect 3999 7517 4065 7540
rect 3679 7498 4065 7517
rect 18799 7603 19185 7622
rect 18799 7580 18865 7603
rect 18951 7580 19033 7603
rect 19119 7580 19185 7603
rect 18799 7540 18808 7580
rect 18848 7540 18865 7580
rect 18951 7540 18972 7580
rect 19012 7540 19033 7580
rect 19119 7540 19136 7580
rect 19176 7540 19185 7580
rect 18799 7517 18865 7540
rect 18951 7517 19033 7540
rect 19119 7517 19185 7540
rect 18799 7498 19185 7517
rect 4919 6847 5305 6866
rect 4919 6824 4985 6847
rect 5071 6824 5153 6847
rect 5239 6824 5305 6847
rect 4919 6784 4928 6824
rect 4968 6784 4985 6824
rect 5071 6784 5092 6824
rect 5132 6784 5153 6824
rect 5239 6784 5256 6824
rect 5296 6784 5305 6824
rect 4919 6761 4985 6784
rect 5071 6761 5153 6784
rect 5239 6761 5305 6784
rect 4919 6742 5305 6761
rect 20039 6847 20425 6866
rect 20039 6824 20105 6847
rect 20191 6824 20273 6847
rect 20359 6824 20425 6847
rect 20039 6784 20048 6824
rect 20088 6784 20105 6824
rect 20191 6784 20212 6824
rect 20252 6784 20273 6824
rect 20359 6784 20376 6824
rect 20416 6784 20425 6824
rect 20039 6761 20105 6784
rect 20191 6761 20273 6784
rect 20359 6761 20425 6784
rect 20039 6742 20425 6761
rect 3679 6091 4065 6110
rect 3679 6068 3745 6091
rect 3831 6068 3913 6091
rect 3999 6068 4065 6091
rect 3679 6028 3688 6068
rect 3728 6028 3745 6068
rect 3831 6028 3852 6068
rect 3892 6028 3913 6068
rect 3999 6028 4016 6068
rect 4056 6028 4065 6068
rect 3679 6005 3745 6028
rect 3831 6005 3913 6028
rect 3999 6005 4065 6028
rect 3679 5986 4065 6005
rect 18799 6091 19185 6110
rect 18799 6068 18865 6091
rect 18951 6068 19033 6091
rect 19119 6068 19185 6091
rect 18799 6028 18808 6068
rect 18848 6028 18865 6068
rect 18951 6028 18972 6068
rect 19012 6028 19033 6068
rect 19119 6028 19136 6068
rect 19176 6028 19185 6068
rect 18799 6005 18865 6028
rect 18951 6005 19033 6028
rect 19119 6005 19185 6028
rect 18799 5986 19185 6005
rect 4919 5335 5305 5354
rect 4919 5312 4985 5335
rect 5071 5312 5153 5335
rect 5239 5312 5305 5335
rect 4919 5272 4928 5312
rect 4968 5272 4985 5312
rect 5071 5272 5092 5312
rect 5132 5272 5153 5312
rect 5239 5272 5256 5312
rect 5296 5272 5305 5312
rect 4919 5249 4985 5272
rect 5071 5249 5153 5272
rect 5239 5249 5305 5272
rect 4919 5230 5305 5249
rect 20039 5335 20425 5354
rect 20039 5312 20105 5335
rect 20191 5312 20273 5335
rect 20359 5312 20425 5335
rect 20039 5272 20048 5312
rect 20088 5272 20105 5312
rect 20191 5272 20212 5312
rect 20252 5272 20273 5312
rect 20359 5272 20376 5312
rect 20416 5272 20425 5312
rect 20039 5249 20105 5272
rect 20191 5249 20273 5272
rect 20359 5249 20425 5272
rect 20039 5230 20425 5249
rect 3679 4579 4065 4598
rect 3679 4556 3745 4579
rect 3831 4556 3913 4579
rect 3999 4556 4065 4579
rect 3679 4516 3688 4556
rect 3728 4516 3745 4556
rect 3831 4516 3852 4556
rect 3892 4516 3913 4556
rect 3999 4516 4016 4556
rect 4056 4516 4065 4556
rect 3679 4493 3745 4516
rect 3831 4493 3913 4516
rect 3999 4493 4065 4516
rect 3679 4474 4065 4493
rect 18799 4579 19185 4598
rect 18799 4556 18865 4579
rect 18951 4556 19033 4579
rect 19119 4556 19185 4579
rect 18799 4516 18808 4556
rect 18848 4516 18865 4556
rect 18951 4516 18972 4556
rect 19012 4516 19033 4556
rect 19119 4516 19136 4556
rect 19176 4516 19185 4556
rect 18799 4493 18865 4516
rect 18951 4493 19033 4516
rect 19119 4493 19185 4516
rect 18799 4474 19185 4493
rect 4919 3823 5305 3842
rect 4919 3800 4985 3823
rect 5071 3800 5153 3823
rect 5239 3800 5305 3823
rect 4919 3760 4928 3800
rect 4968 3760 4985 3800
rect 5071 3760 5092 3800
rect 5132 3760 5153 3800
rect 5239 3760 5256 3800
rect 5296 3760 5305 3800
rect 4919 3737 4985 3760
rect 5071 3737 5153 3760
rect 5239 3737 5305 3760
rect 4919 3718 5305 3737
rect 20039 3823 20425 3842
rect 20039 3800 20105 3823
rect 20191 3800 20273 3823
rect 20359 3800 20425 3823
rect 20039 3760 20048 3800
rect 20088 3760 20105 3800
rect 20191 3760 20212 3800
rect 20252 3760 20273 3800
rect 20359 3760 20376 3800
rect 20416 3760 20425 3800
rect 20039 3737 20105 3760
rect 20191 3737 20273 3760
rect 20359 3737 20425 3760
rect 20039 3718 20425 3737
rect 3679 3067 4065 3086
rect 3679 3044 3745 3067
rect 3831 3044 3913 3067
rect 3999 3044 4065 3067
rect 3679 3004 3688 3044
rect 3728 3004 3745 3044
rect 3831 3004 3852 3044
rect 3892 3004 3913 3044
rect 3999 3004 4016 3044
rect 4056 3004 4065 3044
rect 3679 2981 3745 3004
rect 3831 2981 3913 3004
rect 3999 2981 4065 3004
rect 3679 2962 4065 2981
rect 18799 3067 19185 3086
rect 18799 3044 18865 3067
rect 18951 3044 19033 3067
rect 19119 3044 19185 3067
rect 18799 3004 18808 3044
rect 18848 3004 18865 3044
rect 18951 3004 18972 3044
rect 19012 3004 19033 3044
rect 19119 3004 19136 3044
rect 19176 3004 19185 3044
rect 18799 2981 18865 3004
rect 18951 2981 19033 3004
rect 19119 2981 19185 3004
rect 18799 2962 19185 2981
rect 1219 2752 1228 2792
rect 1268 2752 19276 2792
rect 19316 2752 19325 2792
rect 1219 2416 1228 2456
rect 1268 2416 19372 2456
rect 19412 2416 19421 2456
rect 4919 2311 5305 2330
rect 4919 2288 4985 2311
rect 5071 2288 5153 2311
rect 5239 2288 5305 2311
rect 4919 2248 4928 2288
rect 4968 2248 4985 2288
rect 5071 2248 5092 2288
rect 5132 2248 5153 2288
rect 5239 2248 5256 2288
rect 5296 2248 5305 2288
rect 4919 2225 4985 2248
rect 5071 2225 5153 2248
rect 5239 2225 5305 2248
rect 4919 2206 5305 2225
rect 20039 2311 20425 2330
rect 20039 2288 20105 2311
rect 20191 2288 20273 2311
rect 20359 2288 20425 2311
rect 20039 2248 20048 2288
rect 20088 2248 20105 2288
rect 20191 2248 20212 2288
rect 20252 2248 20273 2288
rect 20359 2248 20376 2288
rect 20416 2248 20425 2288
rect 20039 2225 20105 2248
rect 20191 2225 20273 2248
rect 20359 2225 20425 2248
rect 20039 2206 20425 2225
rect 1219 2080 1228 2120
rect 1268 2080 19756 2120
rect 19796 2080 19805 2120
rect 8707 1912 8716 1952
rect 8756 1912 17644 1952
rect 17684 1912 17693 1952
rect 8035 1828 8044 1868
rect 8084 1828 16108 1868
rect 16148 1828 16157 1868
rect 16268 1828 17740 1868
rect 17780 1828 17789 1868
rect 16268 1784 16308 1828
rect 1699 1744 1708 1784
rect 1748 1744 16308 1784
rect 5827 1660 5836 1700
rect 5876 1660 11308 1700
rect 11348 1660 11357 1700
rect 3679 1555 4065 1574
rect 3679 1532 3745 1555
rect 3831 1532 3913 1555
rect 3999 1532 4065 1555
rect 3679 1492 3688 1532
rect 3728 1492 3745 1532
rect 3831 1492 3852 1532
rect 3892 1492 3913 1532
rect 3999 1492 4016 1532
rect 4056 1492 4065 1532
rect 3679 1469 3745 1492
rect 3831 1469 3913 1492
rect 3999 1469 4065 1492
rect 3679 1450 4065 1469
rect 18799 1555 19185 1574
rect 18799 1532 18865 1555
rect 18951 1532 19033 1555
rect 19119 1532 19185 1555
rect 18799 1492 18808 1532
rect 18848 1492 18865 1532
rect 18951 1492 18972 1532
rect 19012 1492 19033 1532
rect 19119 1492 19136 1532
rect 19176 1492 19185 1532
rect 18799 1469 18865 1492
rect 18951 1469 19033 1492
rect 19119 1469 19185 1492
rect 18799 1450 19185 1469
rect 5347 1240 5356 1280
rect 5396 1240 13900 1280
rect 13940 1240 13949 1280
rect 3235 1156 3244 1196
rect 3284 1156 13996 1196
rect 14036 1156 14045 1196
rect 6595 1072 6604 1112
rect 6644 1072 13324 1112
rect 13364 1072 13373 1112
rect 4919 799 5305 818
rect 4919 776 4985 799
rect 5071 776 5153 799
rect 5239 776 5305 799
rect 4919 736 4928 776
rect 4968 736 4985 776
rect 5071 736 5092 776
rect 5132 736 5153 776
rect 5239 736 5256 776
rect 5296 736 5305 776
rect 4919 713 4985 736
rect 5071 713 5153 736
rect 5239 713 5305 736
rect 4919 694 5305 713
rect 20039 799 20425 818
rect 20039 776 20105 799
rect 20191 776 20273 799
rect 20359 776 20425 799
rect 20039 736 20048 776
rect 20088 736 20105 776
rect 20191 736 20212 776
rect 20252 736 20273 776
rect 20359 736 20376 776
rect 20416 736 20425 776
rect 20039 713 20105 736
rect 20191 713 20273 736
rect 20359 713 20425 736
rect 20039 694 20425 713
rect 7459 568 7468 608
rect 7508 568 15340 608
rect 15380 568 15389 608
rect 6403 400 6412 440
rect 6452 400 13804 440
rect 13844 400 13853 440
<< via5 >>
rect 4985 9848 5071 9871
rect 5153 9848 5239 9871
rect 4985 9808 5010 9848
rect 5010 9808 5050 9848
rect 5050 9808 5071 9848
rect 5153 9808 5174 9848
rect 5174 9808 5214 9848
rect 5214 9808 5239 9848
rect 4985 9785 5071 9808
rect 5153 9785 5239 9808
rect 20105 9848 20191 9871
rect 20273 9848 20359 9871
rect 20105 9808 20130 9848
rect 20130 9808 20170 9848
rect 20170 9808 20191 9848
rect 20273 9808 20294 9848
rect 20294 9808 20334 9848
rect 20334 9808 20359 9848
rect 20105 9785 20191 9808
rect 20273 9785 20359 9808
rect 3745 9092 3831 9115
rect 3913 9092 3999 9115
rect 3745 9052 3770 9092
rect 3770 9052 3810 9092
rect 3810 9052 3831 9092
rect 3913 9052 3934 9092
rect 3934 9052 3974 9092
rect 3974 9052 3999 9092
rect 3745 9029 3831 9052
rect 3913 9029 3999 9052
rect 18865 9092 18951 9115
rect 19033 9092 19119 9115
rect 18865 9052 18890 9092
rect 18890 9052 18930 9092
rect 18930 9052 18951 9092
rect 19033 9052 19054 9092
rect 19054 9052 19094 9092
rect 19094 9052 19119 9092
rect 18865 9029 18951 9052
rect 19033 9029 19119 9052
rect 4985 8336 5071 8359
rect 5153 8336 5239 8359
rect 4985 8296 5010 8336
rect 5010 8296 5050 8336
rect 5050 8296 5071 8336
rect 5153 8296 5174 8336
rect 5174 8296 5214 8336
rect 5214 8296 5239 8336
rect 4985 8273 5071 8296
rect 5153 8273 5239 8296
rect 20105 8336 20191 8359
rect 20273 8336 20359 8359
rect 20105 8296 20130 8336
rect 20130 8296 20170 8336
rect 20170 8296 20191 8336
rect 20273 8296 20294 8336
rect 20294 8296 20334 8336
rect 20334 8296 20359 8336
rect 20105 8273 20191 8296
rect 20273 8273 20359 8296
rect 3745 7580 3831 7603
rect 3913 7580 3999 7603
rect 3745 7540 3770 7580
rect 3770 7540 3810 7580
rect 3810 7540 3831 7580
rect 3913 7540 3934 7580
rect 3934 7540 3974 7580
rect 3974 7540 3999 7580
rect 3745 7517 3831 7540
rect 3913 7517 3999 7540
rect 18865 7580 18951 7603
rect 19033 7580 19119 7603
rect 18865 7540 18890 7580
rect 18890 7540 18930 7580
rect 18930 7540 18951 7580
rect 19033 7540 19054 7580
rect 19054 7540 19094 7580
rect 19094 7540 19119 7580
rect 18865 7517 18951 7540
rect 19033 7517 19119 7540
rect 4985 6824 5071 6847
rect 5153 6824 5239 6847
rect 4985 6784 5010 6824
rect 5010 6784 5050 6824
rect 5050 6784 5071 6824
rect 5153 6784 5174 6824
rect 5174 6784 5214 6824
rect 5214 6784 5239 6824
rect 4985 6761 5071 6784
rect 5153 6761 5239 6784
rect 20105 6824 20191 6847
rect 20273 6824 20359 6847
rect 20105 6784 20130 6824
rect 20130 6784 20170 6824
rect 20170 6784 20191 6824
rect 20273 6784 20294 6824
rect 20294 6784 20334 6824
rect 20334 6784 20359 6824
rect 20105 6761 20191 6784
rect 20273 6761 20359 6784
rect 3745 6068 3831 6091
rect 3913 6068 3999 6091
rect 3745 6028 3770 6068
rect 3770 6028 3810 6068
rect 3810 6028 3831 6068
rect 3913 6028 3934 6068
rect 3934 6028 3974 6068
rect 3974 6028 3999 6068
rect 3745 6005 3831 6028
rect 3913 6005 3999 6028
rect 18865 6068 18951 6091
rect 19033 6068 19119 6091
rect 18865 6028 18890 6068
rect 18890 6028 18930 6068
rect 18930 6028 18951 6068
rect 19033 6028 19054 6068
rect 19054 6028 19094 6068
rect 19094 6028 19119 6068
rect 18865 6005 18951 6028
rect 19033 6005 19119 6028
rect 4985 5312 5071 5335
rect 5153 5312 5239 5335
rect 4985 5272 5010 5312
rect 5010 5272 5050 5312
rect 5050 5272 5071 5312
rect 5153 5272 5174 5312
rect 5174 5272 5214 5312
rect 5214 5272 5239 5312
rect 4985 5249 5071 5272
rect 5153 5249 5239 5272
rect 20105 5312 20191 5335
rect 20273 5312 20359 5335
rect 20105 5272 20130 5312
rect 20130 5272 20170 5312
rect 20170 5272 20191 5312
rect 20273 5272 20294 5312
rect 20294 5272 20334 5312
rect 20334 5272 20359 5312
rect 20105 5249 20191 5272
rect 20273 5249 20359 5272
rect 3745 4556 3831 4579
rect 3913 4556 3999 4579
rect 3745 4516 3770 4556
rect 3770 4516 3810 4556
rect 3810 4516 3831 4556
rect 3913 4516 3934 4556
rect 3934 4516 3974 4556
rect 3974 4516 3999 4556
rect 3745 4493 3831 4516
rect 3913 4493 3999 4516
rect 18865 4556 18951 4579
rect 19033 4556 19119 4579
rect 18865 4516 18890 4556
rect 18890 4516 18930 4556
rect 18930 4516 18951 4556
rect 19033 4516 19054 4556
rect 19054 4516 19094 4556
rect 19094 4516 19119 4556
rect 18865 4493 18951 4516
rect 19033 4493 19119 4516
rect 4985 3800 5071 3823
rect 5153 3800 5239 3823
rect 4985 3760 5010 3800
rect 5010 3760 5050 3800
rect 5050 3760 5071 3800
rect 5153 3760 5174 3800
rect 5174 3760 5214 3800
rect 5214 3760 5239 3800
rect 4985 3737 5071 3760
rect 5153 3737 5239 3760
rect 20105 3800 20191 3823
rect 20273 3800 20359 3823
rect 20105 3760 20130 3800
rect 20130 3760 20170 3800
rect 20170 3760 20191 3800
rect 20273 3760 20294 3800
rect 20294 3760 20334 3800
rect 20334 3760 20359 3800
rect 20105 3737 20191 3760
rect 20273 3737 20359 3760
rect 3745 3044 3831 3067
rect 3913 3044 3999 3067
rect 3745 3004 3770 3044
rect 3770 3004 3810 3044
rect 3810 3004 3831 3044
rect 3913 3004 3934 3044
rect 3934 3004 3974 3044
rect 3974 3004 3999 3044
rect 3745 2981 3831 3004
rect 3913 2981 3999 3004
rect 18865 3044 18951 3067
rect 19033 3044 19119 3067
rect 18865 3004 18890 3044
rect 18890 3004 18930 3044
rect 18930 3004 18951 3044
rect 19033 3004 19054 3044
rect 19054 3004 19094 3044
rect 19094 3004 19119 3044
rect 18865 2981 18951 3004
rect 19033 2981 19119 3004
rect 4985 2288 5071 2311
rect 5153 2288 5239 2311
rect 4985 2248 5010 2288
rect 5010 2248 5050 2288
rect 5050 2248 5071 2288
rect 5153 2248 5174 2288
rect 5174 2248 5214 2288
rect 5214 2248 5239 2288
rect 4985 2225 5071 2248
rect 5153 2225 5239 2248
rect 20105 2288 20191 2311
rect 20273 2288 20359 2311
rect 20105 2248 20130 2288
rect 20130 2248 20170 2288
rect 20170 2248 20191 2288
rect 20273 2248 20294 2288
rect 20294 2248 20334 2288
rect 20334 2248 20359 2288
rect 20105 2225 20191 2248
rect 20273 2225 20359 2248
rect 3745 1532 3831 1555
rect 3913 1532 3999 1555
rect 3745 1492 3770 1532
rect 3770 1492 3810 1532
rect 3810 1492 3831 1532
rect 3913 1492 3934 1532
rect 3934 1492 3974 1532
rect 3974 1492 3999 1532
rect 3745 1469 3831 1492
rect 3913 1469 3999 1492
rect 18865 1532 18951 1555
rect 19033 1532 19119 1555
rect 18865 1492 18890 1532
rect 18890 1492 18930 1532
rect 18930 1492 18951 1532
rect 19033 1492 19054 1532
rect 19054 1492 19094 1532
rect 19094 1492 19119 1532
rect 18865 1469 18951 1492
rect 19033 1469 19119 1492
rect 4985 776 5071 799
rect 5153 776 5239 799
rect 4985 736 5010 776
rect 5010 736 5050 776
rect 5050 736 5071 776
rect 5153 736 5174 776
rect 5174 736 5214 776
rect 5214 736 5239 776
rect 4985 713 5071 736
rect 5153 713 5239 736
rect 20105 776 20191 799
rect 20273 776 20359 799
rect 20105 736 20130 776
rect 20130 736 20170 776
rect 20170 736 20191 776
rect 20273 736 20294 776
rect 20294 736 20334 776
rect 20334 736 20359 776
rect 20105 713 20191 736
rect 20273 713 20359 736
<< metal6 >>
rect 3652 9115 4092 10752
rect 3652 9029 3745 9115
rect 3831 9029 3913 9115
rect 3999 9029 4092 9115
rect 3652 7603 4092 9029
rect 3652 7517 3745 7603
rect 3831 7517 3913 7603
rect 3999 7517 4092 7603
rect 3652 6091 4092 7517
rect 3652 6005 3745 6091
rect 3831 6005 3913 6091
rect 3999 6005 4092 6091
rect 3652 4579 4092 6005
rect 3652 4493 3745 4579
rect 3831 4493 3913 4579
rect 3999 4493 4092 4579
rect 3652 3067 4092 4493
rect 3652 2981 3745 3067
rect 3831 2981 3913 3067
rect 3999 2981 4092 3067
rect 3652 1555 4092 2981
rect 3652 1469 3745 1555
rect 3831 1469 3913 1555
rect 3999 1469 4092 1555
rect 3652 0 4092 1469
rect 4892 9871 5332 10752
rect 4892 9785 4985 9871
rect 5071 9785 5153 9871
rect 5239 9785 5332 9871
rect 4892 8359 5332 9785
rect 4892 8273 4985 8359
rect 5071 8273 5153 8359
rect 5239 8273 5332 8359
rect 4892 6847 5332 8273
rect 4892 6761 4985 6847
rect 5071 6761 5153 6847
rect 5239 6761 5332 6847
rect 4892 5335 5332 6761
rect 4892 5249 4985 5335
rect 5071 5249 5153 5335
rect 5239 5249 5332 5335
rect 4892 3823 5332 5249
rect 4892 3737 4985 3823
rect 5071 3737 5153 3823
rect 5239 3737 5332 3823
rect 4892 2311 5332 3737
rect 4892 2225 4985 2311
rect 5071 2225 5153 2311
rect 5239 2225 5332 2311
rect 4892 799 5332 2225
rect 4892 713 4985 799
rect 5071 713 5153 799
rect 5239 713 5332 799
rect 4892 0 5332 713
rect 18772 9115 19212 10752
rect 18772 9029 18865 9115
rect 18951 9029 19033 9115
rect 19119 9029 19212 9115
rect 18772 7603 19212 9029
rect 18772 7517 18865 7603
rect 18951 7517 19033 7603
rect 19119 7517 19212 7603
rect 18772 6091 19212 7517
rect 18772 6005 18865 6091
rect 18951 6005 19033 6091
rect 19119 6005 19212 6091
rect 18772 4579 19212 6005
rect 18772 4493 18865 4579
rect 18951 4493 19033 4579
rect 19119 4493 19212 4579
rect 18772 3067 19212 4493
rect 18772 2981 18865 3067
rect 18951 2981 19033 3067
rect 19119 2981 19212 3067
rect 18772 1555 19212 2981
rect 18772 1469 18865 1555
rect 18951 1469 19033 1555
rect 19119 1469 19212 1555
rect 18772 0 19212 1469
rect 20012 9871 20452 10752
rect 20012 9785 20105 9871
rect 20191 9785 20273 9871
rect 20359 9785 20452 9871
rect 20012 8359 20452 9785
rect 20012 8273 20105 8359
rect 20191 8273 20273 8359
rect 20359 8273 20452 8359
rect 20012 6847 20452 8273
rect 20012 6761 20105 6847
rect 20191 6761 20273 6847
rect 20359 6761 20452 6847
rect 20012 5335 20452 6761
rect 20012 5249 20105 5335
rect 20191 5249 20273 5335
rect 20359 5249 20452 5335
rect 20012 3823 20452 5249
rect 20012 3737 20105 3823
rect 20191 3737 20273 3823
rect 20359 3737 20452 3823
rect 20012 2311 20452 3737
rect 20012 2225 20105 2311
rect 20191 2225 20273 2311
rect 20359 2225 20452 2311
rect 20012 799 20452 2225
rect 20012 713 20105 799
rect 20191 713 20273 799
rect 20359 713 20452 799
rect 20012 0 20452 713
use sg13g2_buf_1  _00_
timestamp 1676381911
transform 1 0 17280 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _01_
timestamp 1676381911
transform 1 0 16896 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _02_
timestamp 1676381911
transform 1 0 17664 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _03_
timestamp 1676381911
transform 1 0 17280 0 1 756
box -48 -56 432 834
use sg13g2_buf_1  _04_
timestamp 1676381911
transform 1 0 17280 0 1 2268
box -48 -56 432 834
use sg13g2_buf_1  _05_
timestamp 1676381911
transform 1 0 18912 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _06_
timestamp 1676381911
transform 1 0 19680 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _07_
timestamp 1676381911
transform 1 0 19296 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _08_
timestamp 1676381911
transform 1 0 19200 0 -1 3780
box -48 -56 432 834
use sg13g2_buf_1  _09_
timestamp 1676381911
transform 1 0 18720 0 1 3780
box -48 -56 432 834
use sg13g2_buf_1  _10_
timestamp 1676381911
transform 1 0 16608 0 -1 5292
box -48 -56 432 834
use sg13g2_buf_1  _11_
timestamp 1676381911
transform 1 0 17184 0 -1 5292
box -48 -56 432 834
use sg13g2_buf_1  _12_
timestamp 1676381911
transform 1 0 19488 0 1 3780
box -48 -56 432 834
use sg13g2_buf_1  _13_
timestamp 1676381911
transform 1 0 19104 0 1 3780
box -48 -56 432 834
use sg13g2_buf_1  _14_
timestamp 1676381911
transform 1 0 1824 0 -1 5292
box -48 -56 432 834
use sg13g2_buf_1  _15_
timestamp 1676381911
transform 1 0 1824 0 1 5292
box -48 -56 432 834
use sg13g2_buf_1  _16_
timestamp 1676381911
transform 1 0 19104 0 1 5292
box -48 -56 432 834
use sg13g2_buf_1  _17_
timestamp 1676381911
transform 1 0 19200 0 -1 6804
box -48 -56 432 834
use sg13g2_buf_1  _18_
timestamp 1676381911
transform 1 0 1728 0 -1 6804
box -48 -56 432 834
use sg13g2_buf_1  _19_
timestamp 1676381911
transform 1 0 19200 0 1 6804
box -48 -56 432 834
use sg13g2_buf_1  _20_
timestamp 1676381911
transform 1 0 2112 0 -1 6804
box -48 -56 432 834
use sg13g2_buf_1  _21_
timestamp 1676381911
transform 1 0 2496 0 -1 6804
box -48 -56 432 834
use sg13g2_buf_1  _22_
timestamp 1676381911
transform 1 0 19584 0 -1 6804
box -48 -56 432 834
use sg13g2_buf_1  _23_
timestamp 1676381911
transform 1 0 2112 0 -1 8316
box -48 -56 432 834
use sg13g2_buf_1  _24_
timestamp 1676381911
transform 1 0 17856 0 -1 6804
box -48 -56 432 834
use sg13g2_buf_1  _25_
timestamp 1676381911
transform 1 0 13536 0 -1 8316
box -48 -56 432 834
use sg13g2_buf_1  _26_
timestamp 1676381911
transform 1 0 18144 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  _27_
timestamp 1676381911
transform 1 0 11136 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  _28_
timestamp 1676381911
transform 1 0 1824 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  _29_
timestamp 1676381911
transform 1 0 1440 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  _30_
timestamp 1676381911
transform 1 0 2208 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  _31_
timestamp 1676381911
transform 1 0 19296 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  _32_
timestamp 1676381911
transform -1 0 3744 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  _33_
timestamp 1676381911
transform -1 0 4128 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  _34_
timestamp 1676381911
transform -1 0 5088 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  _35_
timestamp 1676381911
transform -1 0 6048 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  _36_
timestamp 1676381911
transform -1 0 6912 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  _37_
timestamp 1676381911
transform -1 0 8160 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  _38_
timestamp 1676381911
transform -1 0 9120 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  _39_
timestamp 1676381911
transform -1 0 9696 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  _40_
timestamp 1676381911
transform -1 0 10752 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  _41_
timestamp 1676381911
transform -1 0 11904 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  _42_
timestamp 1676381911
transform -1 0 12288 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  _43_
timestamp 1676381911
transform -1 0 13344 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  _44_
timestamp 1676381911
transform -1 0 14400 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  _45_
timestamp 1676381911
transform -1 0 15744 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  _46_
timestamp 1676381911
transform -1 0 16416 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  _47_
timestamp 1676381911
transform -1 0 16800 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  _48_
timestamp 1676381911
transform 1 0 16800 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  _49_
timestamp 1676381911
transform 1 0 17568 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  _50_
timestamp 1676381911
transform -1 0 20064 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  _51_
timestamp 1676381911
transform 1 0 18912 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  _52_
timestamp 1676381911
transform 1 0 1824 0 1 2268
box -48 -56 432 834
use sg13g2_buf_1  _53_
timestamp 1676381911
transform 1 0 1824 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _54_
timestamp 1676381911
transform 1 0 2208 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _55_
timestamp 1676381911
transform 1 0 2592 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _56_
timestamp 1676381911
transform 1 0 7584 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _57_
timestamp 1676381911
transform 1 0 7968 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _58_
timestamp 1676381911
transform 1 0 4032 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _59_
timestamp 1676381911
transform 1 0 4416 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _60_
timestamp 1676381911
transform 1 0 3648 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _61_
timestamp 1676381911
transform 1 0 3456 0 1 2268
box -48 -56 432 834
use sg13g2_buf_1  _62_
timestamp 1676381911
transform 1 0 2688 0 1 2268
box -48 -56 432 834
use sg13g2_buf_1  _63_
timestamp 1676381911
transform 1 0 1824 0 -1 3780
box -48 -56 432 834
use sg13g2_buf_1  _64_
timestamp 1676381911
transform 1 0 7200 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _65_
timestamp 1676381911
transform 1 0 10272 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _66_
timestamp 1676381911
transform 1 0 9888 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _67_
timestamp 1676381911
transform 1 0 6816 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _68_
timestamp 1676381911
transform 1 0 6624 0 1 2268
box -48 -56 432 834
use sg13g2_buf_1  _69_
timestamp 1676381911
transform 1 0 6048 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _70_
timestamp 1676381911
transform 1 0 5568 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _71_
timestamp 1676381911
transform 1 0 5088 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _72_
timestamp 1676381911
transform 1 0 10752 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _73_
timestamp 1676381911
transform 1 0 9600 0 1 2268
box -48 -56 432 834
use sg13g2_buf_1  _74_
timestamp 1676381911
transform 1 0 11520 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _75_
timestamp 1676381911
transform 1 0 11136 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _76_
timestamp 1676381911
transform 1 0 8640 0 1 2268
box -48 -56 432 834
use sg13g2_buf_1  _77_
timestamp 1676381911
transform 1 0 8352 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _78_
timestamp 1676381911
transform 1 0 11904 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _79_
timestamp 1676381911
transform 1 0 12768 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _80_
timestamp 1676381911
transform 1 0 13152 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _81_
timestamp 1676381911
transform 1 0 13536 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _82_
timestamp 1676381911
transform 1 0 13920 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _83_
timestamp 1676381911
transform 1 0 14496 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _84_
timestamp 1676381911
transform -1 0 15264 0 1 2268
box -48 -56 432 834
use sg13g2_buf_1  _85_
timestamp 1676381911
transform -1 0 15648 0 1 2268
box -48 -56 432 834
use sg13g2_buf_1  _86_
timestamp 1676381911
transform -1 0 16224 0 1 2268
box -48 -56 432 834
use sg13g2_buf_1  _87_
timestamp 1676381911
transform -1 0 16224 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _88_
timestamp 1676381911
transform -1 0 2208 0 1 3780
box -48 -56 432 834
use sg13g2_decap_8  FILLER_0_0
timestamp 1679581782
transform 1 0 1152 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_7
timestamp 1679581782
transform 1 0 1824 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_14
timestamp 1679581782
transform 1 0 2496 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_21
timestamp 1679581782
transform 1 0 3168 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_28
timestamp 1679581782
transform 1 0 3840 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_35
timestamp 1679581782
transform 1 0 4512 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_42
timestamp 1679581782
transform 1 0 5184 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_49
timestamp 1679581782
transform 1 0 5856 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_56
timestamp 1679581782
transform 1 0 6528 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_63
timestamp 1679581782
transform 1 0 7200 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_70
timestamp 1679581782
transform 1 0 7872 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_77
timestamp 1679581782
transform 1 0 8544 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_84
timestamp 1679581782
transform 1 0 9216 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_91
timestamp 1679581782
transform 1 0 9888 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_98
timestamp 1679581782
transform 1 0 10560 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_105
timestamp 1679581782
transform 1 0 11232 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_112
timestamp 1679581782
transform 1 0 11904 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_119
timestamp 1679581782
transform 1 0 12576 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_126
timestamp 1679581782
transform 1 0 13248 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_133
timestamp 1679581782
transform 1 0 13920 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_140
timestamp 1679581782
transform 1 0 14592 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_147
timestamp 1679581782
transform 1 0 15264 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_154
timestamp 1679581782
transform 1 0 15936 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_161
timestamp 1679581782
transform 1 0 16608 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_172
timestamp 1679581782
transform 1 0 17664 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_179
timestamp 1679581782
transform 1 0 18336 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_186
timestamp 1679581782
transform 1 0 19008 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_193
timestamp 1679581782
transform 1 0 19680 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_0
timestamp 1679581782
transform 1 0 1152 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_19
timestamp 1679581782
transform 1 0 2976 0 -1 2268
box -48 -56 720 834
use sg13g2_fill_2  FILLER_1_38
timestamp 1677580104
transform 1 0 4800 0 -1 2268
box -48 -56 240 834
use sg13g2_fill_1  FILLER_1_40
timestamp 1677579658
transform 1 0 4992 0 -1 2268
box -48 -56 144 834
use sg13g2_fill_1  FILLER_1_45
timestamp 1677579658
transform 1 0 5472 0 -1 2268
box -48 -56 144 834
use sg13g2_fill_1  FILLER_1_50
timestamp 1677579658
transform 1 0 5952 0 -1 2268
box -48 -56 144 834
use sg13g2_decap_4  FILLER_1_55
timestamp 1679577901
transform 1 0 6432 0 -1 2268
box -48 -56 432 834
use sg13g2_decap_8  FILLER_1_79
timestamp 1679581782
transform 1 0 8736 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_4  FILLER_1_86
timestamp 1679577901
transform 1 0 9408 0 -1 2268
box -48 -56 432 834
use sg13g2_fill_1  FILLER_1_90
timestamp 1677579658
transform 1 0 9792 0 -1 2268
box -48 -56 144 834
use sg13g2_fill_1  FILLER_1_99
timestamp 1677579658
transform 1 0 10656 0 -1 2268
box -48 -56 144 834
use sg13g2_decap_4  FILLER_1_116
timestamp 1679577901
transform 1 0 12288 0 -1 2268
box -48 -56 432 834
use sg13g2_fill_1  FILLER_1_120
timestamp 1677579658
transform 1 0 12672 0 -1 2268
box -48 -56 144 834
use sg13g2_fill_2  FILLER_1_137
timestamp 1677580104
transform 1 0 14304 0 -1 2268
box -48 -56 240 834
use sg13g2_decap_8  FILLER_1_143
timestamp 1679581782
transform 1 0 14880 0 -1 2268
box -48 -56 720 834
use sg13g2_fill_2  FILLER_1_150
timestamp 1677580104
transform 1 0 15552 0 -1 2268
box -48 -56 240 834
use sg13g2_fill_1  FILLER_1_152
timestamp 1677579658
transform 1 0 15744 0 -1 2268
box -48 -56 144 834
use sg13g2_decap_8  FILLER_1_157
timestamp 1679581782
transform 1 0 16224 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_176
timestamp 1679581782
transform 1 0 18048 0 -1 2268
box -48 -56 720 834
use sg13g2_fill_2  FILLER_1_183
timestamp 1677580104
transform 1 0 18720 0 -1 2268
box -48 -56 240 834
use sg13g2_fill_2  FILLER_1_197
timestamp 1677580104
transform 1 0 20064 0 -1 2268
box -48 -56 240 834
use sg13g2_fill_1  FILLER_1_199
timestamp 1677579658
transform 1 0 20256 0 -1 2268
box -48 -56 144 834
use sg13g2_decap_8  FILLER_2_0
timestamp 1679581782
transform 1 0 1152 0 1 2268
box -48 -56 720 834
use sg13g2_decap_4  FILLER_2_11
timestamp 1679577901
transform 1 0 2208 0 1 2268
box -48 -56 432 834
use sg13g2_fill_1  FILLER_2_15
timestamp 1677579658
transform 1 0 2592 0 1 2268
box -48 -56 144 834
use sg13g2_decap_4  FILLER_2_20
timestamp 1679577901
transform 1 0 3072 0 1 2268
box -48 -56 432 834
use sg13g2_decap_8  FILLER_2_28
timestamp 1679581782
transform 1 0 3840 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_35
timestamp 1679581782
transform 1 0 4512 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_42
timestamp 1679581782
transform 1 0 5184 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_49
timestamp 1679581782
transform 1 0 5856 0 1 2268
box -48 -56 720 834
use sg13g2_fill_1  FILLER_2_56
timestamp 1677579658
transform 1 0 6528 0 1 2268
box -48 -56 144 834
use sg13g2_decap_8  FILLER_2_61
timestamp 1679581782
transform 1 0 7008 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_68
timestamp 1679581782
transform 1 0 7680 0 1 2268
box -48 -56 720 834
use sg13g2_fill_2  FILLER_2_75
timestamp 1677580104
transform 1 0 8352 0 1 2268
box -48 -56 240 834
use sg13g2_fill_1  FILLER_2_77
timestamp 1677579658
transform 1 0 8544 0 1 2268
box -48 -56 144 834
use sg13g2_decap_4  FILLER_2_82
timestamp 1679577901
transform 1 0 9024 0 1 2268
box -48 -56 432 834
use sg13g2_fill_2  FILLER_2_86
timestamp 1677580104
transform 1 0 9408 0 1 2268
box -48 -56 240 834
use sg13g2_decap_8  FILLER_2_92
timestamp 1679581782
transform 1 0 9984 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_99
timestamp 1679581782
transform 1 0 10656 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_106
timestamp 1679581782
transform 1 0 11328 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_113
timestamp 1679581782
transform 1 0 12000 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_120
timestamp 1679581782
transform 1 0 12672 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_127
timestamp 1679581782
transform 1 0 13344 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_134
timestamp 1679581782
transform 1 0 14016 0 1 2268
box -48 -56 720 834
use sg13g2_fill_2  FILLER_2_141
timestamp 1677580104
transform 1 0 14688 0 1 2268
box -48 -56 240 834
use sg13g2_fill_2  FILLER_2_151
timestamp 1677580104
transform 1 0 15648 0 1 2268
box -48 -56 240 834
use sg13g2_decap_8  FILLER_2_157
timestamp 1679581782
transform 1 0 16224 0 1 2268
box -48 -56 720 834
use sg13g2_decap_4  FILLER_2_164
timestamp 1679577901
transform 1 0 16896 0 1 2268
box -48 -56 432 834
use sg13g2_decap_8  FILLER_2_172
timestamp 1679581782
transform 1 0 17664 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_179
timestamp 1679581782
transform 1 0 18336 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_186
timestamp 1679581782
transform 1 0 19008 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_193
timestamp 1679581782
transform 1 0 19680 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_0
timestamp 1679581782
transform 1 0 1152 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_11
timestamp 1679581782
transform 1 0 2208 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_18
timestamp 1679581782
transform 1 0 2880 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_25
timestamp 1679581782
transform 1 0 3552 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_32
timestamp 1679581782
transform 1 0 4224 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_39
timestamp 1679581782
transform 1 0 4896 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_46
timestamp 1679581782
transform 1 0 5568 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_53
timestamp 1679581782
transform 1 0 6240 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_60
timestamp 1679581782
transform 1 0 6912 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_67
timestamp 1679581782
transform 1 0 7584 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_74
timestamp 1679581782
transform 1 0 8256 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_81
timestamp 1679581782
transform 1 0 8928 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_88
timestamp 1679581782
transform 1 0 9600 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_95
timestamp 1679581782
transform 1 0 10272 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_102
timestamp 1679581782
transform 1 0 10944 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_109
timestamp 1679581782
transform 1 0 11616 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_116
timestamp 1679581782
transform 1 0 12288 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_123
timestamp 1679581782
transform 1 0 12960 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_130
timestamp 1679581782
transform 1 0 13632 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_137
timestamp 1679581782
transform 1 0 14304 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_144
timestamp 1679581782
transform 1 0 14976 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_151
timestamp 1679581782
transform 1 0 15648 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_158
timestamp 1679581782
transform 1 0 16320 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_165
timestamp 1679581782
transform 1 0 16992 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_172
timestamp 1679581782
transform 1 0 17664 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_179
timestamp 1679581782
transform 1 0 18336 0 -1 3780
box -48 -56 720 834
use sg13g2_fill_2  FILLER_3_186
timestamp 1677580104
transform 1 0 19008 0 -1 3780
box -48 -56 240 834
use sg13g2_decap_8  FILLER_3_192
timestamp 1679581782
transform 1 0 19584 0 -1 3780
box -48 -56 720 834
use sg13g2_fill_1  FILLER_3_199
timestamp 1677579658
transform 1 0 20256 0 -1 3780
box -48 -56 144 834
use sg13g2_decap_8  FILLER_4_0
timestamp 1679581782
transform 1 0 1152 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_11
timestamp 1679581782
transform 1 0 2208 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_18
timestamp 1679581782
transform 1 0 2880 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_25
timestamp 1679581782
transform 1 0 3552 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_32
timestamp 1679581782
transform 1 0 4224 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_39
timestamp 1679581782
transform 1 0 4896 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_46
timestamp 1679581782
transform 1 0 5568 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_53
timestamp 1679581782
transform 1 0 6240 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_60
timestamp 1679581782
transform 1 0 6912 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_67
timestamp 1679581782
transform 1 0 7584 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_74
timestamp 1679581782
transform 1 0 8256 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_81
timestamp 1679581782
transform 1 0 8928 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_88
timestamp 1679581782
transform 1 0 9600 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_95
timestamp 1679581782
transform 1 0 10272 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_102
timestamp 1679581782
transform 1 0 10944 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_109
timestamp 1679581782
transform 1 0 11616 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_116
timestamp 1679581782
transform 1 0 12288 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_123
timestamp 1679581782
transform 1 0 12960 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_130
timestamp 1679581782
transform 1 0 13632 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_137
timestamp 1679581782
transform 1 0 14304 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_144
timestamp 1679581782
transform 1 0 14976 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_151
timestamp 1679581782
transform 1 0 15648 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_158
timestamp 1679581782
transform 1 0 16320 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_165
timestamp 1679581782
transform 1 0 16992 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_172
timestamp 1679581782
transform 1 0 17664 0 1 3780
box -48 -56 720 834
use sg13g2_decap_4  FILLER_4_179
timestamp 1679577901
transform 1 0 18336 0 1 3780
box -48 -56 432 834
use sg13g2_decap_4  FILLER_4_195
timestamp 1679577901
transform 1 0 19872 0 1 3780
box -48 -56 432 834
use sg13g2_fill_1  FILLER_4_199
timestamp 1677579658
transform 1 0 20256 0 1 3780
box -48 -56 144 834
use sg13g2_decap_8  FILLER_5_0
timestamp 1679581782
transform 1 0 1152 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_11
timestamp 1679581782
transform 1 0 2208 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_18
timestamp 1679581782
transform 1 0 2880 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_25
timestamp 1679581782
transform 1 0 3552 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_32
timestamp 1679581782
transform 1 0 4224 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_39
timestamp 1679581782
transform 1 0 4896 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_46
timestamp 1679581782
transform 1 0 5568 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_53
timestamp 1679581782
transform 1 0 6240 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_60
timestamp 1679581782
transform 1 0 6912 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_67
timestamp 1679581782
transform 1 0 7584 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_74
timestamp 1679581782
transform 1 0 8256 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_81
timestamp 1679581782
transform 1 0 8928 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_88
timestamp 1679581782
transform 1 0 9600 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_95
timestamp 1679581782
transform 1 0 10272 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_102
timestamp 1679581782
transform 1 0 10944 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_109
timestamp 1679581782
transform 1 0 11616 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_116
timestamp 1679581782
transform 1 0 12288 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_123
timestamp 1679581782
transform 1 0 12960 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_130
timestamp 1679581782
transform 1 0 13632 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_137
timestamp 1679581782
transform 1 0 14304 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_144
timestamp 1679581782
transform 1 0 14976 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_151
timestamp 1679581782
transform 1 0 15648 0 -1 5292
box -48 -56 720 834
use sg13g2_fill_2  FILLER_5_158
timestamp 1677580104
transform 1 0 16320 0 -1 5292
box -48 -56 240 834
use sg13g2_fill_1  FILLER_5_160
timestamp 1677579658
transform 1 0 16512 0 -1 5292
box -48 -56 144 834
use sg13g2_fill_2  FILLER_5_165
timestamp 1677580104
transform 1 0 16992 0 -1 5292
box -48 -56 240 834
use sg13g2_decap_8  FILLER_5_171
timestamp 1679581782
transform 1 0 17568 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_178
timestamp 1679581782
transform 1 0 18240 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_185
timestamp 1679581782
transform 1 0 18912 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_192
timestamp 1679581782
transform 1 0 19584 0 -1 5292
box -48 -56 720 834
use sg13g2_fill_1  FILLER_5_199
timestamp 1677579658
transform 1 0 20256 0 -1 5292
box -48 -56 144 834
use sg13g2_decap_8  FILLER_6_0
timestamp 1679581782
transform 1 0 1152 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_11
timestamp 1679581782
transform 1 0 2208 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_18
timestamp 1679581782
transform 1 0 2880 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_25
timestamp 1679581782
transform 1 0 3552 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_32
timestamp 1679581782
transform 1 0 4224 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_39
timestamp 1679581782
transform 1 0 4896 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_46
timestamp 1679581782
transform 1 0 5568 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_53
timestamp 1679581782
transform 1 0 6240 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_60
timestamp 1679581782
transform 1 0 6912 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_67
timestamp 1679581782
transform 1 0 7584 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_74
timestamp 1679581782
transform 1 0 8256 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_81
timestamp 1679581782
transform 1 0 8928 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_88
timestamp 1679581782
transform 1 0 9600 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_95
timestamp 1679581782
transform 1 0 10272 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_102
timestamp 1679581782
transform 1 0 10944 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_109
timestamp 1679581782
transform 1 0 11616 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_116
timestamp 1679581782
transform 1 0 12288 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_123
timestamp 1679581782
transform 1 0 12960 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_130
timestamp 1679581782
transform 1 0 13632 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_137
timestamp 1679581782
transform 1 0 14304 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_144
timestamp 1679581782
transform 1 0 14976 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_151
timestamp 1679581782
transform 1 0 15648 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_158
timestamp 1679581782
transform 1 0 16320 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_165
timestamp 1679581782
transform 1 0 16992 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_172
timestamp 1679581782
transform 1 0 17664 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_179
timestamp 1679581782
transform 1 0 18336 0 1 5292
box -48 -56 720 834
use sg13g2_fill_1  FILLER_6_186
timestamp 1677579658
transform 1 0 19008 0 1 5292
box -48 -56 144 834
use sg13g2_decap_8  FILLER_6_191
timestamp 1679581782
transform 1 0 19488 0 1 5292
box -48 -56 720 834
use sg13g2_fill_2  FILLER_6_198
timestamp 1677580104
transform 1 0 20160 0 1 5292
box -48 -56 240 834
use sg13g2_decap_4  FILLER_7_0
timestamp 1679577901
transform 1 0 1152 0 -1 6804
box -48 -56 432 834
use sg13g2_fill_2  FILLER_7_4
timestamp 1677580104
transform 1 0 1536 0 -1 6804
box -48 -56 240 834
use sg13g2_decap_8  FILLER_7_18
timestamp 1679581782
transform 1 0 2880 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_25
timestamp 1679581782
transform 1 0 3552 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_32
timestamp 1679581782
transform 1 0 4224 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_39
timestamp 1679581782
transform 1 0 4896 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_46
timestamp 1679581782
transform 1 0 5568 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_53
timestamp 1679581782
transform 1 0 6240 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_60
timestamp 1679581782
transform 1 0 6912 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_67
timestamp 1679581782
transform 1 0 7584 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_74
timestamp 1679581782
transform 1 0 8256 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_81
timestamp 1679581782
transform 1 0 8928 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_88
timestamp 1679581782
transform 1 0 9600 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_95
timestamp 1679581782
transform 1 0 10272 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_102
timestamp 1679581782
transform 1 0 10944 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_109
timestamp 1679581782
transform 1 0 11616 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_116
timestamp 1679581782
transform 1 0 12288 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_123
timestamp 1679581782
transform 1 0 12960 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_130
timestamp 1679581782
transform 1 0 13632 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_137
timestamp 1679581782
transform 1 0 14304 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_144
timestamp 1679581782
transform 1 0 14976 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_151
timestamp 1679581782
transform 1 0 15648 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_158
timestamp 1679581782
transform 1 0 16320 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_165
timestamp 1679581782
transform 1 0 16992 0 -1 6804
box -48 -56 720 834
use sg13g2_fill_2  FILLER_7_172
timestamp 1677580104
transform 1 0 17664 0 -1 6804
box -48 -56 240 834
use sg13g2_decap_8  FILLER_7_178
timestamp 1679581782
transform 1 0 18240 0 -1 6804
box -48 -56 720 834
use sg13g2_fill_2  FILLER_7_185
timestamp 1677580104
transform 1 0 18912 0 -1 6804
box -48 -56 240 834
use sg13g2_fill_1  FILLER_7_187
timestamp 1677579658
transform 1 0 19104 0 -1 6804
box -48 -56 144 834
use sg13g2_decap_4  FILLER_7_196
timestamp 1679577901
transform 1 0 19968 0 -1 6804
box -48 -56 432 834
use sg13g2_decap_8  FILLER_8_0
timestamp 1679581782
transform 1 0 1152 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_7
timestamp 1679581782
transform 1 0 1824 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_14
timestamp 1679581782
transform 1 0 2496 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_21
timestamp 1679581782
transform 1 0 3168 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_28
timestamp 1679581782
transform 1 0 3840 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_35
timestamp 1679581782
transform 1 0 4512 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_42
timestamp 1679581782
transform 1 0 5184 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_49
timestamp 1679581782
transform 1 0 5856 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_56
timestamp 1679581782
transform 1 0 6528 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_63
timestamp 1679581782
transform 1 0 7200 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_70
timestamp 1679581782
transform 1 0 7872 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_77
timestamp 1679581782
transform 1 0 8544 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_84
timestamp 1679581782
transform 1 0 9216 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_91
timestamp 1679581782
transform 1 0 9888 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_98
timestamp 1679581782
transform 1 0 10560 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_105
timestamp 1679581782
transform 1 0 11232 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_112
timestamp 1679581782
transform 1 0 11904 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_119
timestamp 1679581782
transform 1 0 12576 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_126
timestamp 1679581782
transform 1 0 13248 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_133
timestamp 1679581782
transform 1 0 13920 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_140
timestamp 1679581782
transform 1 0 14592 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_147
timestamp 1679581782
transform 1 0 15264 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_154
timestamp 1679581782
transform 1 0 15936 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_161
timestamp 1679581782
transform 1 0 16608 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_168
timestamp 1679581782
transform 1 0 17280 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_175
timestamp 1679581782
transform 1 0 17952 0 1 6804
box -48 -56 720 834
use sg13g2_decap_4  FILLER_8_182
timestamp 1679577901
transform 1 0 18624 0 1 6804
box -48 -56 432 834
use sg13g2_fill_2  FILLER_8_186
timestamp 1677580104
transform 1 0 19008 0 1 6804
box -48 -56 240 834
use sg13g2_decap_8  FILLER_8_192
timestamp 1679581782
transform 1 0 19584 0 1 6804
box -48 -56 720 834
use sg13g2_fill_1  FILLER_8_199
timestamp 1677579658
transform 1 0 20256 0 1 6804
box -48 -56 144 834
use sg13g2_decap_8  FILLER_9_0
timestamp 1679581782
transform 1 0 1152 0 -1 8316
box -48 -56 720 834
use sg13g2_fill_2  FILLER_9_7
timestamp 1677580104
transform 1 0 1824 0 -1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_9_9
timestamp 1677579658
transform 1 0 2016 0 -1 8316
box -48 -56 144 834
use sg13g2_decap_8  FILLER_9_14
timestamp 1679581782
transform 1 0 2496 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_21
timestamp 1679581782
transform 1 0 3168 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_28
timestamp 1679581782
transform 1 0 3840 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_35
timestamp 1679581782
transform 1 0 4512 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_42
timestamp 1679581782
transform 1 0 5184 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_49
timestamp 1679581782
transform 1 0 5856 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_56
timestamp 1679581782
transform 1 0 6528 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_63
timestamp 1679581782
transform 1 0 7200 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_70
timestamp 1679581782
transform 1 0 7872 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_77
timestamp 1679581782
transform 1 0 8544 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_84
timestamp 1679581782
transform 1 0 9216 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_91
timestamp 1679581782
transform 1 0 9888 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_98
timestamp 1679581782
transform 1 0 10560 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_105
timestamp 1679581782
transform 1 0 11232 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_112
timestamp 1679581782
transform 1 0 11904 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_119
timestamp 1679581782
transform 1 0 12576 0 -1 8316
box -48 -56 720 834
use sg13g2_fill_2  FILLER_9_126
timestamp 1677580104
transform 1 0 13248 0 -1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_9_128
timestamp 1677579658
transform 1 0 13440 0 -1 8316
box -48 -56 144 834
use sg13g2_decap_8  FILLER_9_133
timestamp 1679581782
transform 1 0 13920 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_140
timestamp 1679581782
transform 1 0 14592 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_147
timestamp 1679581782
transform 1 0 15264 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_154
timestamp 1679581782
transform 1 0 15936 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_161
timestamp 1679581782
transform 1 0 16608 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_168
timestamp 1679581782
transform 1 0 17280 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_175
timestamp 1679581782
transform 1 0 17952 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_182
timestamp 1679581782
transform 1 0 18624 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_189
timestamp 1679581782
transform 1 0 19296 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_4  FILLER_9_196
timestamp 1679577901
transform 1 0 19968 0 -1 8316
box -48 -56 432 834
use sg13g2_fill_2  FILLER_10_0
timestamp 1677580104
transform 1 0 1152 0 1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_10_2
timestamp 1677579658
transform 1 0 1344 0 1 8316
box -48 -56 144 834
use sg13g2_decap_8  FILLER_10_15
timestamp 1679581782
transform 1 0 2592 0 1 8316
box -48 -56 720 834
use sg13g2_fill_1  FILLER_10_22
timestamp 1677579658
transform 1 0 3264 0 1 8316
box -48 -56 144 834
use sg13g2_decap_4  FILLER_10_31
timestamp 1679577901
transform 1 0 4128 0 1 8316
box -48 -56 432 834
use sg13g2_fill_2  FILLER_10_35
timestamp 1677580104
transform 1 0 4512 0 1 8316
box -48 -56 240 834
use sg13g2_decap_4  FILLER_10_41
timestamp 1679577901
transform 1 0 5088 0 1 8316
box -48 -56 432 834
use sg13g2_fill_2  FILLER_10_45
timestamp 1677580104
transform 1 0 5472 0 1 8316
box -48 -56 240 834
use sg13g2_decap_4  FILLER_10_51
timestamp 1679577901
transform 1 0 6048 0 1 8316
box -48 -56 432 834
use sg13g2_fill_1  FILLER_10_55
timestamp 1677579658
transform 1 0 6432 0 1 8316
box -48 -56 144 834
use sg13g2_decap_8  FILLER_10_60
timestamp 1679581782
transform 1 0 6912 0 1 8316
box -48 -56 720 834
use sg13g2_fill_2  FILLER_10_67
timestamp 1677580104
transform 1 0 7584 0 1 8316
box -48 -56 240 834
use sg13g2_decap_4  FILLER_10_73
timestamp 1679577901
transform 1 0 8160 0 1 8316
box -48 -56 432 834
use sg13g2_fill_2  FILLER_10_77
timestamp 1677580104
transform 1 0 8544 0 1 8316
box -48 -56 240 834
use sg13g2_fill_2  FILLER_10_83
timestamp 1677580104
transform 1 0 9120 0 1 8316
box -48 -56 240 834
use sg13g2_decap_8  FILLER_10_89
timestamp 1679581782
transform 1 0 9696 0 1 8316
box -48 -56 720 834
use sg13g2_decap_4  FILLER_10_100
timestamp 1679577901
transform 1 0 10752 0 1 8316
box -48 -56 432 834
use sg13g2_decap_8  FILLER_10_116
timestamp 1679581782
transform 1 0 12288 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_127
timestamp 1679581782
transform 1 0 13344 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_138
timestamp 1679581782
transform 1 0 14400 0 1 8316
box -48 -56 720 834
use sg13g2_fill_2  FILLER_10_145
timestamp 1677580104
transform 1 0 15072 0 1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_10_147
timestamp 1677579658
transform 1 0 15264 0 1 8316
box -48 -56 144 834
use sg13g2_fill_2  FILLER_10_152
timestamp 1677580104
transform 1 0 15744 0 1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_10_154
timestamp 1677579658
transform 1 0 15936 0 1 8316
box -48 -56 144 834
use sg13g2_decap_4  FILLER_10_167
timestamp 1679577901
transform 1 0 17184 0 1 8316
box -48 -56 432 834
use sg13g2_fill_2  FILLER_10_175
timestamp 1677580104
transform 1 0 17952 0 1 8316
box -48 -56 240 834
use sg13g2_decap_4  FILLER_10_181
timestamp 1679577901
transform 1 0 18528 0 1 8316
box -48 -56 432 834
use sg13g2_fill_2  FILLER_10_197
timestamp 1677580104
transform 1 0 20064 0 1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_10_199
timestamp 1677579658
transform 1 0 20256 0 1 8316
box -48 -56 144 834
use sg13g2_decap_8  FILLER_11_0
timestamp 1679581782
transform 1 0 1152 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_7
timestamp 1679581782
transform 1 0 1824 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_14
timestamp 1679581782
transform 1 0 2496 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_21
timestamp 1679581782
transform 1 0 3168 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_28
timestamp 1679581782
transform 1 0 3840 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_35
timestamp 1679581782
transform 1 0 4512 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_42
timestamp 1679581782
transform 1 0 5184 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_49
timestamp 1679581782
transform 1 0 5856 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_56
timestamp 1679581782
transform 1 0 6528 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_63
timestamp 1679581782
transform 1 0 7200 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_70
timestamp 1679581782
transform 1 0 7872 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_77
timestamp 1679581782
transform 1 0 8544 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_84
timestamp 1679581782
transform 1 0 9216 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_91
timestamp 1679581782
transform 1 0 9888 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_98
timestamp 1679581782
transform 1 0 10560 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_105
timestamp 1679581782
transform 1 0 11232 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_112
timestamp 1679581782
transform 1 0 11904 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_119
timestamp 1679581782
transform 1 0 12576 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_126
timestamp 1679581782
transform 1 0 13248 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_133
timestamp 1679581782
transform 1 0 13920 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_140
timestamp 1679581782
transform 1 0 14592 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_147
timestamp 1679581782
transform 1 0 15264 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_154
timestamp 1679581782
transform 1 0 15936 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_161
timestamp 1679581782
transform 1 0 16608 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_168
timestamp 1679581782
transform 1 0 17280 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_175
timestamp 1679581782
transform 1 0 17952 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_182
timestamp 1679581782
transform 1 0 18624 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_189
timestamp 1679581782
transform 1 0 19296 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_4  FILLER_11_196
timestamp 1679577901
transform 1 0 19968 0 -1 9828
box -48 -56 432 834
<< labels >>
flabel metal3 s 0 44 80 124 0 FreeSans 320 0 0 0 FrameData[0]
port 0 nsew signal input
flabel metal3 s 0 3404 80 3484 0 FreeSans 320 0 0 0 FrameData[10]
port 1 nsew signal input
flabel metal3 s 0 3740 80 3820 0 FreeSans 320 0 0 0 FrameData[11]
port 2 nsew signal input
flabel metal3 s 0 4076 80 4156 0 FreeSans 320 0 0 0 FrameData[12]
port 3 nsew signal input
flabel metal3 s 0 4412 80 4492 0 FreeSans 320 0 0 0 FrameData[13]
port 4 nsew signal input
flabel metal3 s 0 4748 80 4828 0 FreeSans 320 0 0 0 FrameData[14]
port 5 nsew signal input
flabel metal3 s 0 5084 80 5164 0 FreeSans 320 0 0 0 FrameData[15]
port 6 nsew signal input
flabel metal3 s 0 5420 80 5500 0 FreeSans 320 0 0 0 FrameData[16]
port 7 nsew signal input
flabel metal3 s 0 5756 80 5836 0 FreeSans 320 0 0 0 FrameData[17]
port 8 nsew signal input
flabel metal3 s 0 6092 80 6172 0 FreeSans 320 0 0 0 FrameData[18]
port 9 nsew signal input
flabel metal3 s 0 6428 80 6508 0 FreeSans 320 0 0 0 FrameData[19]
port 10 nsew signal input
flabel metal3 s 0 380 80 460 0 FreeSans 320 0 0 0 FrameData[1]
port 11 nsew signal input
flabel metal3 s 0 6764 80 6844 0 FreeSans 320 0 0 0 FrameData[20]
port 12 nsew signal input
flabel metal3 s 0 7100 80 7180 0 FreeSans 320 0 0 0 FrameData[21]
port 13 nsew signal input
flabel metal3 s 0 7436 80 7516 0 FreeSans 320 0 0 0 FrameData[22]
port 14 nsew signal input
flabel metal3 s 0 7772 80 7852 0 FreeSans 320 0 0 0 FrameData[23]
port 15 nsew signal input
flabel metal3 s 0 8108 80 8188 0 FreeSans 320 0 0 0 FrameData[24]
port 16 nsew signal input
flabel metal3 s 0 8444 80 8524 0 FreeSans 320 0 0 0 FrameData[25]
port 17 nsew signal input
flabel metal3 s 0 8780 80 8860 0 FreeSans 320 0 0 0 FrameData[26]
port 18 nsew signal input
flabel metal3 s 0 9116 80 9196 0 FreeSans 320 0 0 0 FrameData[27]
port 19 nsew signal input
flabel metal3 s 0 9452 80 9532 0 FreeSans 320 0 0 0 FrameData[28]
port 20 nsew signal input
flabel metal3 s 0 9788 80 9868 0 FreeSans 320 0 0 0 FrameData[29]
port 21 nsew signal input
flabel metal3 s 0 716 80 796 0 FreeSans 320 0 0 0 FrameData[2]
port 22 nsew signal input
flabel metal3 s 0 10124 80 10204 0 FreeSans 320 0 0 0 FrameData[30]
port 23 nsew signal input
flabel metal3 s 0 10460 80 10540 0 FreeSans 320 0 0 0 FrameData[31]
port 24 nsew signal input
flabel metal3 s 0 1052 80 1132 0 FreeSans 320 0 0 0 FrameData[3]
port 25 nsew signal input
flabel metal3 s 0 1388 80 1468 0 FreeSans 320 0 0 0 FrameData[4]
port 26 nsew signal input
flabel metal3 s 0 1724 80 1804 0 FreeSans 320 0 0 0 FrameData[5]
port 27 nsew signal input
flabel metal3 s 0 2060 80 2140 0 FreeSans 320 0 0 0 FrameData[6]
port 28 nsew signal input
flabel metal3 s 0 2396 80 2476 0 FreeSans 320 0 0 0 FrameData[7]
port 29 nsew signal input
flabel metal3 s 0 2732 80 2812 0 FreeSans 320 0 0 0 FrameData[8]
port 30 nsew signal input
flabel metal3 s 0 3068 80 3148 0 FreeSans 320 0 0 0 FrameData[9]
port 31 nsew signal input
flabel metal3 s 21424 44 21504 124 0 FreeSans 320 0 0 0 FrameData_O[0]
port 32 nsew signal output
flabel metal3 s 21424 3404 21504 3484 0 FreeSans 320 0 0 0 FrameData_O[10]
port 33 nsew signal output
flabel metal3 s 21424 3740 21504 3820 0 FreeSans 320 0 0 0 FrameData_O[11]
port 34 nsew signal output
flabel metal3 s 21424 4076 21504 4156 0 FreeSans 320 0 0 0 FrameData_O[12]
port 35 nsew signal output
flabel metal3 s 21424 4412 21504 4492 0 FreeSans 320 0 0 0 FrameData_O[13]
port 36 nsew signal output
flabel metal3 s 21424 4748 21504 4828 0 FreeSans 320 0 0 0 FrameData_O[14]
port 37 nsew signal output
flabel metal3 s 21424 5084 21504 5164 0 FreeSans 320 0 0 0 FrameData_O[15]
port 38 nsew signal output
flabel metal3 s 21424 5420 21504 5500 0 FreeSans 320 0 0 0 FrameData_O[16]
port 39 nsew signal output
flabel metal3 s 21424 5756 21504 5836 0 FreeSans 320 0 0 0 FrameData_O[17]
port 40 nsew signal output
flabel metal3 s 21424 6092 21504 6172 0 FreeSans 320 0 0 0 FrameData_O[18]
port 41 nsew signal output
flabel metal3 s 21424 6428 21504 6508 0 FreeSans 320 0 0 0 FrameData_O[19]
port 42 nsew signal output
flabel metal3 s 21424 380 21504 460 0 FreeSans 320 0 0 0 FrameData_O[1]
port 43 nsew signal output
flabel metal3 s 21424 6764 21504 6844 0 FreeSans 320 0 0 0 FrameData_O[20]
port 44 nsew signal output
flabel metal3 s 21424 7100 21504 7180 0 FreeSans 320 0 0 0 FrameData_O[21]
port 45 nsew signal output
flabel metal3 s 21424 7436 21504 7516 0 FreeSans 320 0 0 0 FrameData_O[22]
port 46 nsew signal output
flabel metal3 s 21424 7772 21504 7852 0 FreeSans 320 0 0 0 FrameData_O[23]
port 47 nsew signal output
flabel metal3 s 21424 8108 21504 8188 0 FreeSans 320 0 0 0 FrameData_O[24]
port 48 nsew signal output
flabel metal3 s 21424 8444 21504 8524 0 FreeSans 320 0 0 0 FrameData_O[25]
port 49 nsew signal output
flabel metal3 s 21424 8780 21504 8860 0 FreeSans 320 0 0 0 FrameData_O[26]
port 50 nsew signal output
flabel metal3 s 21424 9116 21504 9196 0 FreeSans 320 0 0 0 FrameData_O[27]
port 51 nsew signal output
flabel metal3 s 21424 9452 21504 9532 0 FreeSans 320 0 0 0 FrameData_O[28]
port 52 nsew signal output
flabel metal3 s 21424 9788 21504 9868 0 FreeSans 320 0 0 0 FrameData_O[29]
port 53 nsew signal output
flabel metal3 s 21424 716 21504 796 0 FreeSans 320 0 0 0 FrameData_O[2]
port 54 nsew signal output
flabel metal3 s 21424 10124 21504 10204 0 FreeSans 320 0 0 0 FrameData_O[30]
port 55 nsew signal output
flabel metal3 s 21424 10460 21504 10540 0 FreeSans 320 0 0 0 FrameData_O[31]
port 56 nsew signal output
flabel metal3 s 21424 1052 21504 1132 0 FreeSans 320 0 0 0 FrameData_O[3]
port 57 nsew signal output
flabel metal3 s 21424 1388 21504 1468 0 FreeSans 320 0 0 0 FrameData_O[4]
port 58 nsew signal output
flabel metal3 s 21424 1724 21504 1804 0 FreeSans 320 0 0 0 FrameData_O[5]
port 59 nsew signal output
flabel metal3 s 21424 2060 21504 2140 0 FreeSans 320 0 0 0 FrameData_O[6]
port 60 nsew signal output
flabel metal3 s 21424 2396 21504 2476 0 FreeSans 320 0 0 0 FrameData_O[7]
port 61 nsew signal output
flabel metal3 s 21424 2732 21504 2812 0 FreeSans 320 0 0 0 FrameData_O[8]
port 62 nsew signal output
flabel metal3 s 21424 3068 21504 3148 0 FreeSans 320 0 0 0 FrameData_O[9]
port 63 nsew signal output
flabel metal2 s 15800 0 15880 80 0 FreeSans 320 0 0 0 FrameStrobe[0]
port 64 nsew signal input
flabel metal2 s 17720 0 17800 80 0 FreeSans 320 0 0 0 FrameStrobe[10]
port 65 nsew signal input
flabel metal2 s 17912 0 17992 80 0 FreeSans 320 0 0 0 FrameStrobe[11]
port 66 nsew signal input
flabel metal2 s 18104 0 18184 80 0 FreeSans 320 0 0 0 FrameStrobe[12]
port 67 nsew signal input
flabel metal2 s 18296 0 18376 80 0 FreeSans 320 0 0 0 FrameStrobe[13]
port 68 nsew signal input
flabel metal2 s 18488 0 18568 80 0 FreeSans 320 0 0 0 FrameStrobe[14]
port 69 nsew signal input
flabel metal2 s 18680 0 18760 80 0 FreeSans 320 0 0 0 FrameStrobe[15]
port 70 nsew signal input
flabel metal2 s 18872 0 18952 80 0 FreeSans 320 0 0 0 FrameStrobe[16]
port 71 nsew signal input
flabel metal2 s 19064 0 19144 80 0 FreeSans 320 0 0 0 FrameStrobe[17]
port 72 nsew signal input
flabel metal2 s 19256 0 19336 80 0 FreeSans 320 0 0 0 FrameStrobe[18]
port 73 nsew signal input
flabel metal2 s 19448 0 19528 80 0 FreeSans 320 0 0 0 FrameStrobe[19]
port 74 nsew signal input
flabel metal2 s 15992 0 16072 80 0 FreeSans 320 0 0 0 FrameStrobe[1]
port 75 nsew signal input
flabel metal2 s 16184 0 16264 80 0 FreeSans 320 0 0 0 FrameStrobe[2]
port 76 nsew signal input
flabel metal2 s 16376 0 16456 80 0 FreeSans 320 0 0 0 FrameStrobe[3]
port 77 nsew signal input
flabel metal2 s 16568 0 16648 80 0 FreeSans 320 0 0 0 FrameStrobe[4]
port 78 nsew signal input
flabel metal2 s 16760 0 16840 80 0 FreeSans 320 0 0 0 FrameStrobe[5]
port 79 nsew signal input
flabel metal2 s 16952 0 17032 80 0 FreeSans 320 0 0 0 FrameStrobe[6]
port 80 nsew signal input
flabel metal2 s 17144 0 17224 80 0 FreeSans 320 0 0 0 FrameStrobe[7]
port 81 nsew signal input
flabel metal2 s 17336 0 17416 80 0 FreeSans 320 0 0 0 FrameStrobe[8]
port 82 nsew signal input
flabel metal2 s 17528 0 17608 80 0 FreeSans 320 0 0 0 FrameStrobe[9]
port 83 nsew signal input
flabel metal2 s 1976 10672 2056 10752 0 FreeSans 320 0 0 0 FrameStrobe_O[0]
port 84 nsew signal output
flabel metal2 s 11576 10672 11656 10752 0 FreeSans 320 0 0 0 FrameStrobe_O[10]
port 85 nsew signal output
flabel metal2 s 12536 10672 12616 10752 0 FreeSans 320 0 0 0 FrameStrobe_O[11]
port 86 nsew signal output
flabel metal2 s 13496 10672 13576 10752 0 FreeSans 320 0 0 0 FrameStrobe_O[12]
port 87 nsew signal output
flabel metal2 s 14456 10672 14536 10752 0 FreeSans 320 0 0 0 FrameStrobe_O[13]
port 88 nsew signal output
flabel metal2 s 15416 10672 15496 10752 0 FreeSans 320 0 0 0 FrameStrobe_O[14]
port 89 nsew signal output
flabel metal2 s 16376 10672 16456 10752 0 FreeSans 320 0 0 0 FrameStrobe_O[15]
port 90 nsew signal output
flabel metal2 s 17336 10672 17416 10752 0 FreeSans 320 0 0 0 FrameStrobe_O[16]
port 91 nsew signal output
flabel metal2 s 18296 10672 18376 10752 0 FreeSans 320 0 0 0 FrameStrobe_O[17]
port 92 nsew signal output
flabel metal2 s 19256 10672 19336 10752 0 FreeSans 320 0 0 0 FrameStrobe_O[18]
port 93 nsew signal output
flabel metal2 s 20216 10672 20296 10752 0 FreeSans 320 0 0 0 FrameStrobe_O[19]
port 94 nsew signal output
flabel metal2 s 2936 10672 3016 10752 0 FreeSans 320 0 0 0 FrameStrobe_O[1]
port 95 nsew signal output
flabel metal2 s 3896 10672 3976 10752 0 FreeSans 320 0 0 0 FrameStrobe_O[2]
port 96 nsew signal output
flabel metal2 s 4856 10672 4936 10752 0 FreeSans 320 0 0 0 FrameStrobe_O[3]
port 97 nsew signal output
flabel metal2 s 5816 10672 5896 10752 0 FreeSans 320 0 0 0 FrameStrobe_O[4]
port 98 nsew signal output
flabel metal2 s 6776 10672 6856 10752 0 FreeSans 320 0 0 0 FrameStrobe_O[5]
port 99 nsew signal output
flabel metal2 s 7736 10672 7816 10752 0 FreeSans 320 0 0 0 FrameStrobe_O[6]
port 100 nsew signal output
flabel metal2 s 8696 10672 8776 10752 0 FreeSans 320 0 0 0 FrameStrobe_O[7]
port 101 nsew signal output
flabel metal2 s 9656 10672 9736 10752 0 FreeSans 320 0 0 0 FrameStrobe_O[8]
port 102 nsew signal output
flabel metal2 s 10616 10672 10696 10752 0 FreeSans 320 0 0 0 FrameStrobe_O[9]
port 103 nsew signal output
flabel metal2 s 1784 0 1864 80 0 FreeSans 320 0 0 0 N1END[0]
port 104 nsew signal input
flabel metal2 s 1976 0 2056 80 0 FreeSans 320 0 0 0 N1END[1]
port 105 nsew signal input
flabel metal2 s 2168 0 2248 80 0 FreeSans 320 0 0 0 N1END[2]
port 106 nsew signal input
flabel metal2 s 2360 0 2440 80 0 FreeSans 320 0 0 0 N1END[3]
port 107 nsew signal input
flabel metal2 s 4088 0 4168 80 0 FreeSans 320 0 0 0 N2END[0]
port 108 nsew signal input
flabel metal2 s 4280 0 4360 80 0 FreeSans 320 0 0 0 N2END[1]
port 109 nsew signal input
flabel metal2 s 4472 0 4552 80 0 FreeSans 320 0 0 0 N2END[2]
port 110 nsew signal input
flabel metal2 s 4664 0 4744 80 0 FreeSans 320 0 0 0 N2END[3]
port 111 nsew signal input
flabel metal2 s 4856 0 4936 80 0 FreeSans 320 0 0 0 N2END[4]
port 112 nsew signal input
flabel metal2 s 5048 0 5128 80 0 FreeSans 320 0 0 0 N2END[5]
port 113 nsew signal input
flabel metal2 s 5240 0 5320 80 0 FreeSans 320 0 0 0 N2END[6]
port 114 nsew signal input
flabel metal2 s 5432 0 5512 80 0 FreeSans 320 0 0 0 N2END[7]
port 115 nsew signal input
flabel metal2 s 2552 0 2632 80 0 FreeSans 320 0 0 0 N2MID[0]
port 116 nsew signal input
flabel metal2 s 2744 0 2824 80 0 FreeSans 320 0 0 0 N2MID[1]
port 117 nsew signal input
flabel metal2 s 2936 0 3016 80 0 FreeSans 320 0 0 0 N2MID[2]
port 118 nsew signal input
flabel metal2 s 3128 0 3208 80 0 FreeSans 320 0 0 0 N2MID[3]
port 119 nsew signal input
flabel metal2 s 3320 0 3400 80 0 FreeSans 320 0 0 0 N2MID[4]
port 120 nsew signal input
flabel metal2 s 3512 0 3592 80 0 FreeSans 320 0 0 0 N2MID[5]
port 121 nsew signal input
flabel metal2 s 3704 0 3784 80 0 FreeSans 320 0 0 0 N2MID[6]
port 122 nsew signal input
flabel metal2 s 3896 0 3976 80 0 FreeSans 320 0 0 0 N2MID[7]
port 123 nsew signal input
flabel metal2 s 5624 0 5704 80 0 FreeSans 320 0 0 0 N4END[0]
port 124 nsew signal input
flabel metal2 s 7544 0 7624 80 0 FreeSans 320 0 0 0 N4END[10]
port 125 nsew signal input
flabel metal2 s 7736 0 7816 80 0 FreeSans 320 0 0 0 N4END[11]
port 126 nsew signal input
flabel metal2 s 7928 0 8008 80 0 FreeSans 320 0 0 0 N4END[12]
port 127 nsew signal input
flabel metal2 s 8120 0 8200 80 0 FreeSans 320 0 0 0 N4END[13]
port 128 nsew signal input
flabel metal2 s 8312 0 8392 80 0 FreeSans 320 0 0 0 N4END[14]
port 129 nsew signal input
flabel metal2 s 8504 0 8584 80 0 FreeSans 320 0 0 0 N4END[15]
port 130 nsew signal input
flabel metal2 s 5816 0 5896 80 0 FreeSans 320 0 0 0 N4END[1]
port 131 nsew signal input
flabel metal2 s 6008 0 6088 80 0 FreeSans 320 0 0 0 N4END[2]
port 132 nsew signal input
flabel metal2 s 6200 0 6280 80 0 FreeSans 320 0 0 0 N4END[3]
port 133 nsew signal input
flabel metal2 s 6392 0 6472 80 0 FreeSans 320 0 0 0 N4END[4]
port 134 nsew signal input
flabel metal2 s 6584 0 6664 80 0 FreeSans 320 0 0 0 N4END[5]
port 135 nsew signal input
flabel metal2 s 6776 0 6856 80 0 FreeSans 320 0 0 0 N4END[6]
port 136 nsew signal input
flabel metal2 s 6968 0 7048 80 0 FreeSans 320 0 0 0 N4END[7]
port 137 nsew signal input
flabel metal2 s 7160 0 7240 80 0 FreeSans 320 0 0 0 N4END[8]
port 138 nsew signal input
flabel metal2 s 7352 0 7432 80 0 FreeSans 320 0 0 0 N4END[9]
port 139 nsew signal input
flabel metal2 s 8696 0 8776 80 0 FreeSans 320 0 0 0 S1BEG[0]
port 140 nsew signal output
flabel metal2 s 8888 0 8968 80 0 FreeSans 320 0 0 0 S1BEG[1]
port 141 nsew signal output
flabel metal2 s 9080 0 9160 80 0 FreeSans 320 0 0 0 S1BEG[2]
port 142 nsew signal output
flabel metal2 s 9272 0 9352 80 0 FreeSans 320 0 0 0 S1BEG[3]
port 143 nsew signal output
flabel metal2 s 9464 0 9544 80 0 FreeSans 320 0 0 0 S2BEG[0]
port 144 nsew signal output
flabel metal2 s 9656 0 9736 80 0 FreeSans 320 0 0 0 S2BEG[1]
port 145 nsew signal output
flabel metal2 s 9848 0 9928 80 0 FreeSans 320 0 0 0 S2BEG[2]
port 146 nsew signal output
flabel metal2 s 10040 0 10120 80 0 FreeSans 320 0 0 0 S2BEG[3]
port 147 nsew signal output
flabel metal2 s 10232 0 10312 80 0 FreeSans 320 0 0 0 S2BEG[4]
port 148 nsew signal output
flabel metal2 s 10424 0 10504 80 0 FreeSans 320 0 0 0 S2BEG[5]
port 149 nsew signal output
flabel metal2 s 10616 0 10696 80 0 FreeSans 320 0 0 0 S2BEG[6]
port 150 nsew signal output
flabel metal2 s 10808 0 10888 80 0 FreeSans 320 0 0 0 S2BEG[7]
port 151 nsew signal output
flabel metal2 s 11000 0 11080 80 0 FreeSans 320 0 0 0 S2BEGb[0]
port 152 nsew signal output
flabel metal2 s 11192 0 11272 80 0 FreeSans 320 0 0 0 S2BEGb[1]
port 153 nsew signal output
flabel metal2 s 11384 0 11464 80 0 FreeSans 320 0 0 0 S2BEGb[2]
port 154 nsew signal output
flabel metal2 s 11576 0 11656 80 0 FreeSans 320 0 0 0 S2BEGb[3]
port 155 nsew signal output
flabel metal2 s 11768 0 11848 80 0 FreeSans 320 0 0 0 S2BEGb[4]
port 156 nsew signal output
flabel metal2 s 11960 0 12040 80 0 FreeSans 320 0 0 0 S2BEGb[5]
port 157 nsew signal output
flabel metal2 s 12152 0 12232 80 0 FreeSans 320 0 0 0 S2BEGb[6]
port 158 nsew signal output
flabel metal2 s 12344 0 12424 80 0 FreeSans 320 0 0 0 S2BEGb[7]
port 159 nsew signal output
flabel metal2 s 12536 0 12616 80 0 FreeSans 320 0 0 0 S4BEG[0]
port 160 nsew signal output
flabel metal2 s 14456 0 14536 80 0 FreeSans 320 0 0 0 S4BEG[10]
port 161 nsew signal output
flabel metal2 s 14648 0 14728 80 0 FreeSans 320 0 0 0 S4BEG[11]
port 162 nsew signal output
flabel metal2 s 14840 0 14920 80 0 FreeSans 320 0 0 0 S4BEG[12]
port 163 nsew signal output
flabel metal2 s 15032 0 15112 80 0 FreeSans 320 0 0 0 S4BEG[13]
port 164 nsew signal output
flabel metal2 s 15224 0 15304 80 0 FreeSans 320 0 0 0 S4BEG[14]
port 165 nsew signal output
flabel metal2 s 15416 0 15496 80 0 FreeSans 320 0 0 0 S4BEG[15]
port 166 nsew signal output
flabel metal2 s 12728 0 12808 80 0 FreeSans 320 0 0 0 S4BEG[1]
port 167 nsew signal output
flabel metal2 s 12920 0 13000 80 0 FreeSans 320 0 0 0 S4BEG[2]
port 168 nsew signal output
flabel metal2 s 13112 0 13192 80 0 FreeSans 320 0 0 0 S4BEG[3]
port 169 nsew signal output
flabel metal2 s 13304 0 13384 80 0 FreeSans 320 0 0 0 S4BEG[4]
port 170 nsew signal output
flabel metal2 s 13496 0 13576 80 0 FreeSans 320 0 0 0 S4BEG[5]
port 171 nsew signal output
flabel metal2 s 13688 0 13768 80 0 FreeSans 320 0 0 0 S4BEG[6]
port 172 nsew signal output
flabel metal2 s 13880 0 13960 80 0 FreeSans 320 0 0 0 S4BEG[7]
port 173 nsew signal output
flabel metal2 s 14072 0 14152 80 0 FreeSans 320 0 0 0 S4BEG[8]
port 174 nsew signal output
flabel metal2 s 14264 0 14344 80 0 FreeSans 320 0 0 0 S4BEG[9]
port 175 nsew signal output
flabel metal2 s 15608 0 15688 80 0 FreeSans 320 0 0 0 UserCLK
port 176 nsew signal input
flabel metal2 s 1016 10672 1096 10752 0 FreeSans 320 0 0 0 UserCLKo
port 177 nsew signal output
flabel metal6 s 4892 0 5332 10752 0 FreeSans 2624 90 0 0 VGND
port 178 nsew ground bidirectional
flabel metal6 s 4892 0 5332 328 0 FreeSans 2624 0 0 0 VGND
port 178 nsew ground bidirectional
flabel metal6 s 4892 10424 5332 10752 0 FreeSans 2624 0 0 0 VGND
port 178 nsew ground bidirectional
flabel metal6 s 20012 0 20452 10752 0 FreeSans 2624 90 0 0 VGND
port 178 nsew ground bidirectional
flabel metal6 s 20012 0 20452 328 0 FreeSans 2624 0 0 0 VGND
port 178 nsew ground bidirectional
flabel metal6 s 20012 10424 20452 10752 0 FreeSans 2624 0 0 0 VGND
port 178 nsew ground bidirectional
flabel metal6 s 3652 0 4092 10752 0 FreeSans 2624 90 0 0 VPWR
port 179 nsew power bidirectional
flabel metal6 s 3652 0 4092 328 0 FreeSans 2624 0 0 0 VPWR
port 179 nsew power bidirectional
flabel metal6 s 3652 10424 4092 10752 0 FreeSans 2624 0 0 0 VPWR
port 179 nsew power bidirectional
flabel metal6 s 18772 0 19212 10752 0 FreeSans 2624 90 0 0 VPWR
port 179 nsew power bidirectional
flabel metal6 s 18772 0 19212 328 0 FreeSans 2624 0 0 0 VPWR
port 179 nsew power bidirectional
flabel metal6 s 18772 10424 19212 10752 0 FreeSans 2624 0 0 0 VPWR
port 179 nsew power bidirectional
rlabel metal1 10802 9828 10802 9828 0 VGND
rlabel metal1 10752 9072 10752 9072 0 VPWR
rlabel metal3 1662 84 1662 84 0 FrameData[0]
rlabel metal2 6432 4158 6432 4158 0 FrameData[10]
rlabel metal3 1614 3780 1614 3780 0 FrameData[11]
rlabel metal3 19584 4158 19584 4158 0 FrameData[12]
rlabel metal2 19200 4284 19200 4284 0 FrameData[13]
rlabel metal3 990 4788 990 4788 0 FrameData[14]
rlabel metal3 990 5124 990 5124 0 FrameData[15]
rlabel metal2 19200 5544 19200 5544 0 FrameData[16]
rlabel metal3 17856 6384 17856 6384 0 FrameData[17]
rlabel metal3 942 6132 942 6132 0 FrameData[18]
rlabel metal2 19200 6846 19200 6846 0 FrameData[19]
rlabel metal3 2718 420 2718 420 0 FrameData[1]
rlabel metal3 1134 6804 1134 6804 0 FrameData[20]
rlabel metal3 1326 7140 1326 7140 0 FrameData[21]
rlabel metal2 19680 6930 19680 6930 0 FrameData[22]
rlabel metal3 1134 7812 1134 7812 0 FrameData[23]
rlabel metal2 17952 7266 17952 7266 0 FrameData[24]
rlabel metal3 1038 8484 1038 8484 0 FrameData[25]
rlabel metal2 18240 8820 18240 8820 0 FrameData[26]
rlabel metal2 11232 8946 11232 8946 0 FrameData[27]
rlabel metal3 990 9492 990 9492 0 FrameData[28]
rlabel metal3 798 9828 798 9828 0 FrameData[29]
rlabel metal3 894 756 894 756 0 FrameData[2]
rlabel metal3 1182 10164 1182 10164 0 FrameData[30]
rlabel metal3 318 10500 318 10500 0 FrameData[31]
rlabel metal3 16368 588 16368 588 0 FrameData[3]
rlabel metal3 1662 1428 1662 1428 0 FrameData[4]
rlabel metal3 18336 1932 18336 1932 0 FrameData[5]
rlabel metal3 654 2100 654 2100 0 FrameData[6]
rlabel metal3 654 2436 654 2436 0 FrameData[7]
rlabel metal3 654 2772 654 2772 0 FrameData[8]
rlabel metal3 654 3108 654 3108 0 FrameData[9]
rlabel metal3 19458 84 19458 84 0 FrameData_O[0]
rlabel metal3 19170 3444 19170 3444 0 FrameData_O[10]
rlabel metal3 20994 3780 20994 3780 0 FrameData_O[11]
rlabel metal3 20610 4116 20610 4116 0 FrameData_O[12]
rlabel metal2 19392 4410 19392 4410 0 FrameData_O[13]
rlabel metal3 21378 4788 21378 4788 0 FrameData_O[14]
rlabel metal2 2160 5544 2160 5544 0 FrameData_O[15]
rlabel metal3 20418 5460 20418 5460 0 FrameData_O[16]
rlabel metal3 20466 5796 20466 5796 0 FrameData_O[17]
rlabel metal3 4158 6216 4158 6216 0 FrameData_O[18]
rlabel metal3 20466 6468 20466 6468 0 FrameData_O[19]
rlabel metal3 19314 420 19314 420 0 FrameData_O[1]
rlabel metal2 2400 6678 2400 6678 0 FrameData_O[20]
rlabel metal3 2784 6594 2784 6594 0 FrameData_O[21]
rlabel metal2 19872 7056 19872 7056 0 FrameData_O[22]
rlabel metal3 19890 7812 19890 7812 0 FrameData_O[23]
rlabel metal2 18144 7392 18144 7392 0 FrameData_O[24]
rlabel via2 21426 8484 21426 8484 0 FrameData_O[25]
rlabel metal3 19938 8820 19938 8820 0 FrameData_O[26]
rlabel metal2 11424 8988 11424 8988 0 FrameData_O[27]
rlabel metal3 2112 8526 2112 8526 0 FrameData_O[28]
rlabel metal2 3936 8484 3936 8484 0 FrameData_O[29]
rlabel metal3 20994 756 20994 756 0 FrameData_O[2]
rlabel metal3 21378 10164 21378 10164 0 FrameData_O[30]
rlabel metal2 19584 9660 19584 9660 0 FrameData_O[31]
rlabel metal3 19506 1092 19506 1092 0 FrameData_O[3]
rlabel metal3 19554 1428 19554 1428 0 FrameData_O[4]
rlabel metal3 20322 1764 20322 1764 0 FrameData_O[5]
rlabel metal3 20706 2100 20706 2100 0 FrameData_O[6]
rlabel metal2 19584 2268 19584 2268 0 FrameData_O[7]
rlabel metal3 20466 2772 20466 2772 0 FrameData_O[8]
rlabel metal3 20226 3108 20226 3108 0 FrameData_O[9]
rlabel metal2 15840 2844 15840 2844 0 FrameStrobe[0]
rlabel metal2 17760 366 17760 366 0 FrameStrobe[10]
rlabel metal2 17952 366 17952 366 0 FrameStrobe[11]
rlabel metal2 18144 1710 18144 1710 0 FrameStrobe[12]
rlabel metal2 18336 1668 18336 1668 0 FrameStrobe[13]
rlabel metal2 18528 1626 18528 1626 0 FrameStrobe[14]
rlabel metal2 18720 660 18720 660 0 FrameStrobe[15]
rlabel metal2 18912 702 18912 702 0 FrameStrobe[16]
rlabel metal2 19104 702 19104 702 0 FrameStrobe[17]
rlabel metal2 19296 1542 19296 1542 0 FrameStrobe[18]
rlabel metal2 19488 1332 19488 1332 0 FrameStrobe[19]
rlabel metal2 5184 7434 5184 7434 0 FrameStrobe[1]
rlabel metal2 4800 7686 4800 7686 0 FrameStrobe[2]
rlabel metal2 16416 660 16416 660 0 FrameStrobe[3]
rlabel metal2 16608 2886 16608 2886 0 FrameStrobe[4]
rlabel metal2 16800 1500 16800 1500 0 FrameStrobe[5]
rlabel metal2 16992 576 16992 576 0 FrameStrobe[6]
rlabel metal2 17184 156 17184 156 0 FrameStrobe[7]
rlabel metal2 17376 240 17376 240 0 FrameStrobe[8]
rlabel metal2 17568 408 17568 408 0 FrameStrobe[9]
rlabel metal2 3456 8736 3456 8736 0 FrameStrobe_O[0]
rlabel metal2 12000 9766 12000 9766 0 FrameStrobe_O[10]
rlabel metal3 12816 8820 12816 8820 0 FrameStrobe_O[11]
rlabel metal3 13824 8820 13824 8820 0 FrameStrobe_O[12]
rlabel metal2 14496 9756 14496 9756 0 FrameStrobe_O[13]
rlabel metal2 16128 9766 16128 9766 0 FrameStrobe_O[14]
rlabel metal2 16464 8820 16464 8820 0 FrameStrobe_O[15]
rlabel metal2 17088 9198 17088 9198 0 FrameStrobe_O[16]
rlabel metal2 17856 9766 17856 9766 0 FrameStrobe_O[17]
rlabel metal2 19776 9766 19776 9766 0 FrameStrobe_O[18]
rlabel metal3 19872 8484 19872 8484 0 FrameStrobe_O[19]
rlabel metal2 3840 8778 3840 8778 0 FrameStrobe_O[1]
rlabel metal2 4752 8820 4752 8820 0 FrameStrobe_O[2]
rlabel metal2 5760 8778 5760 8778 0 FrameStrobe_O[3]
rlabel metal2 5856 10638 5856 10638 0 FrameStrobe_O[4]
rlabel metal2 7872 8778 7872 8778 0 FrameStrobe_O[5]
rlabel metal2 8832 9282 8832 9282 0 FrameStrobe_O[6]
rlabel metal3 9072 8820 9072 8820 0 FrameStrobe_O[7]
rlabel metal3 10080 8820 10080 8820 0 FrameStrobe_O[8]
rlabel metal2 11616 8778 11616 8778 0 FrameStrobe_O[9]
rlabel metal2 1824 954 1824 954 0 N1END[0]
rlabel metal2 2016 492 2016 492 0 N1END[1]
rlabel metal2 2208 408 2208 408 0 N1END[2]
rlabel metal2 2400 1374 2400 1374 0 N1END[3]
rlabel metal2 4128 492 4128 492 0 N2END[0]
rlabel metal2 4320 660 4320 660 0 N2END[1]
rlabel metal2 4512 492 4512 492 0 N2END[2]
rlabel metal2 4704 702 4704 702 0 N2END[3]
rlabel metal2 4896 324 4896 324 0 N2END[4]
rlabel metal2 5088 282 5088 282 0 N2END[5]
rlabel metal2 5280 198 5280 198 0 N2END[6]
rlabel metal2 5472 954 5472 954 0 N2END[7]
rlabel metal2 2592 1038 2592 1038 0 N2MID[0]
rlabel metal2 2784 1374 2784 1374 0 N2MID[1]
rlabel metal2 2976 702 2976 702 0 N2MID[2]
rlabel metal2 3168 954 3168 954 0 N2MID[3]
rlabel metal2 3360 702 3360 702 0 N2MID[4]
rlabel metal2 3552 660 3552 660 0 N2MID[5]
rlabel metal2 3744 492 3744 492 0 N2MID[6]
rlabel metal2 3936 450 3936 450 0 N2MID[7]
rlabel metal2 5664 366 5664 366 0 N4END[0]
rlabel metal2 7584 324 7584 324 0 N4END[10]
rlabel metal2 7776 1374 7776 1374 0 N4END[11]
rlabel metal2 7968 72 7968 72 0 N4END[12]
rlabel metal2 8160 198 8160 198 0 N4END[13]
rlabel metal2 8352 1290 8352 1290 0 N4END[14]
rlabel metal2 8544 450 8544 450 0 N4END[15]
rlabel metal2 5856 282 5856 282 0 N4END[1]
rlabel metal2 6048 1458 6048 1458 0 N4END[2]
rlabel metal2 6240 1542 6240 1542 0 N4END[3]
rlabel metal2 6432 240 6432 240 0 N4END[4]
rlabel metal2 6624 492 6624 492 0 N4END[5]
rlabel metal2 6816 828 6816 828 0 N4END[6]
rlabel metal2 7008 1920 7008 1920 0 N4END[7]
rlabel metal2 7200 702 7200 702 0 N4END[8]
rlabel via2 7392 72 7392 72 0 N4END[9]
rlabel metal2 2208 1806 2208 1806 0 S1BEG[0]
rlabel metal2 2112 2184 2112 2184 0 S1BEG[1]
rlabel metal2 2496 3024 2496 3024 0 S1BEG[2]
rlabel metal3 2880 2058 2880 2058 0 S1BEG[3]
rlabel metal2 9504 492 9504 492 0 S2BEG[0]
rlabel metal2 9696 870 9696 870 0 S2BEG[1]
rlabel metal2 4416 966 4416 966 0 S2BEG[2]
rlabel metal2 4704 1596 4704 1596 0 S2BEG[3]
rlabel metal2 4800 924 4800 924 0 S2BEG[4]
rlabel metal2 3648 2856 3648 2856 0 S2BEG[5]
rlabel metal2 2976 2898 2976 2898 0 S2BEG[6]
rlabel metal2 10848 156 10848 156 0 S2BEG[7]
rlabel metal2 11040 366 11040 366 0 S2BEGb[0]
rlabel metal2 11232 534 11232 534 0 S2BEGb[1]
rlabel metal2 11424 492 11424 492 0 S2BEGb[2]
rlabel metal2 11616 408 11616 408 0 S2BEGb[3]
rlabel metal2 11808 408 11808 408 0 S2BEGb[4]
rlabel metal2 12000 744 12000 744 0 S2BEGb[5]
rlabel metal2 12192 450 12192 450 0 S2BEGb[6]
rlabel metal2 12384 1080 12384 1080 0 S2BEGb[7]
rlabel metal2 12576 450 12576 450 0 S4BEG[0]
rlabel metal2 14496 870 14496 870 0 S4BEG[10]
rlabel metal2 14688 870 14688 870 0 S4BEG[11]
rlabel metal2 14880 1248 14880 1248 0 S4BEG[12]
rlabel metal2 15072 1248 15072 1248 0 S4BEG[13]
rlabel metal2 15264 954 15264 954 0 S4BEG[14]
rlabel metal2 15456 870 15456 870 0 S4BEG[15]
rlabel metal2 12768 618 12768 618 0 S4BEG[1]
rlabel metal2 12960 492 12960 492 0 S4BEG[2]
rlabel metal2 13152 576 13152 576 0 S4BEG[3]
rlabel metal2 13344 240 13344 240 0 S4BEG[4]
rlabel metal2 13536 324 13536 324 0 S4BEG[5]
rlabel metal2 13728 534 13728 534 0 S4BEG[6]
rlabel metal2 13920 408 13920 408 0 S4BEG[7]
rlabel metal2 14112 492 14112 492 0 S4BEG[8]
rlabel metal2 14304 450 14304 450 0 S4BEG[9]
rlabel metal2 15648 2130 15648 2130 0 UserCLK
rlabel metal3 1488 4368 1488 4368 0 UserCLKo
<< properties >>
string FIXED_BBOX 0 0 21504 10752
<< end >>
