module E_TT_IF2 (CLK_TT_PROJECT,
    ENA_TT_PROJECT,
    RST_N_TT_PROJECT,
    Tile_X0Y0_UserCLKo,
    Tile_X0Y1_UserCLK,
    UIO_IN_TT_PROJECT0,
    UIO_IN_TT_PROJECT1,
    UIO_IN_TT_PROJECT2,
    UIO_IN_TT_PROJECT3,
    UIO_IN_TT_PROJECT4,
    UIO_IN_TT_PROJECT5,
    UIO_IN_TT_PROJECT6,
    UIO_IN_TT_PROJECT7,
    UIO_OE_TT_PROJECT0,
    UIO_OE_TT_PROJECT1,
    UIO_OE_TT_PROJECT2,
    UIO_OE_TT_PROJECT3,
    UIO_OE_TT_PROJECT4,
    UIO_OE_TT_PROJECT5,
    UIO_OE_TT_PROJECT6,
    UIO_OE_TT_PROJECT7,
    UIO_OUT_TT_PROJECT0,
    UIO_OUT_TT_PROJECT1,
    UIO_OUT_TT_PROJECT2,
    UIO_OUT_TT_PROJECT3,
    UIO_OUT_TT_PROJECT4,
    UIO_OUT_TT_PROJECT5,
    UIO_OUT_TT_PROJECT6,
    UIO_OUT_TT_PROJECT7,
    UI_IN_TT_PROJECT0,
    UI_IN_TT_PROJECT1,
    UI_IN_TT_PROJECT2,
    UI_IN_TT_PROJECT3,
    UI_IN_TT_PROJECT4,
    UI_IN_TT_PROJECT5,
    UI_IN_TT_PROJECT6,
    UI_IN_TT_PROJECT7,
    UO_OUT_TT_PROJECT0,
    UO_OUT_TT_PROJECT1,
    UO_OUT_TT_PROJECT2,
    UO_OUT_TT_PROJECT3,
    UO_OUT_TT_PROJECT4,
    UO_OUT_TT_PROJECT5,
    UO_OUT_TT_PROJECT6,
    UO_OUT_TT_PROJECT7,
    VPWR,
    VGND,
    Tile_X0Y0_E1END,
    Tile_X0Y0_E2END,
    Tile_X0Y0_E2MID,
    Tile_X0Y0_E6END,
    Tile_X0Y0_EE4END,
    Tile_X0Y0_FrameData,
    Tile_X0Y0_FrameData_O,
    Tile_X0Y0_FrameStrobe_O,
    Tile_X0Y0_N1BEG,
    Tile_X0Y0_N2BEG,
    Tile_X0Y0_N2BEGb,
    Tile_X0Y0_N4BEG,
    Tile_X0Y0_S1END,
    Tile_X0Y0_S2END,
    Tile_X0Y0_S2MID,
    Tile_X0Y0_S4END,
    Tile_X0Y0_W1BEG,
    Tile_X0Y0_W2BEG,
    Tile_X0Y0_W2BEGb,
    Tile_X0Y0_W6BEG,
    Tile_X0Y0_WW4BEG,
    Tile_X0Y1_E1END,
    Tile_X0Y1_E2END,
    Tile_X0Y1_E2MID,
    Tile_X0Y1_E6END,
    Tile_X0Y1_EE4END,
    Tile_X0Y1_FrameData,
    Tile_X0Y1_FrameData_O,
    Tile_X0Y1_FrameStrobe,
    Tile_X0Y1_N1END,
    Tile_X0Y1_N2END,
    Tile_X0Y1_N2MID,
    Tile_X0Y1_N4END,
    Tile_X0Y1_S1BEG,
    Tile_X0Y1_S2BEG,
    Tile_X0Y1_S2BEGb,
    Tile_X0Y1_S4BEG,
    Tile_X0Y1_W1BEG,
    Tile_X0Y1_W2BEG,
    Tile_X0Y1_W2BEGb,
    Tile_X0Y1_W6BEG,
    Tile_X0Y1_WW4BEG);
 output CLK_TT_PROJECT;
 output ENA_TT_PROJECT;
 output RST_N_TT_PROJECT;
 output Tile_X0Y0_UserCLKo;
 input Tile_X0Y1_UserCLK;
 output UIO_IN_TT_PROJECT0;
 output UIO_IN_TT_PROJECT1;
 output UIO_IN_TT_PROJECT2;
 output UIO_IN_TT_PROJECT3;
 output UIO_IN_TT_PROJECT4;
 output UIO_IN_TT_PROJECT5;
 output UIO_IN_TT_PROJECT6;
 output UIO_IN_TT_PROJECT7;
 input UIO_OE_TT_PROJECT0;
 input UIO_OE_TT_PROJECT1;
 input UIO_OE_TT_PROJECT2;
 input UIO_OE_TT_PROJECT3;
 input UIO_OE_TT_PROJECT4;
 input UIO_OE_TT_PROJECT5;
 input UIO_OE_TT_PROJECT6;
 input UIO_OE_TT_PROJECT7;
 input UIO_OUT_TT_PROJECT0;
 input UIO_OUT_TT_PROJECT1;
 input UIO_OUT_TT_PROJECT2;
 input UIO_OUT_TT_PROJECT3;
 input UIO_OUT_TT_PROJECT4;
 input UIO_OUT_TT_PROJECT5;
 input UIO_OUT_TT_PROJECT6;
 input UIO_OUT_TT_PROJECT7;
 output UI_IN_TT_PROJECT0;
 output UI_IN_TT_PROJECT1;
 output UI_IN_TT_PROJECT2;
 output UI_IN_TT_PROJECT3;
 output UI_IN_TT_PROJECT4;
 output UI_IN_TT_PROJECT5;
 output UI_IN_TT_PROJECT6;
 output UI_IN_TT_PROJECT7;
 input UO_OUT_TT_PROJECT0;
 input UO_OUT_TT_PROJECT1;
 input UO_OUT_TT_PROJECT2;
 input UO_OUT_TT_PROJECT3;
 input UO_OUT_TT_PROJECT4;
 input UO_OUT_TT_PROJECT5;
 input UO_OUT_TT_PROJECT6;
 input UO_OUT_TT_PROJECT7;
 inout VPWR;
 inout VGND;
 input [3:0] Tile_X0Y0_E1END;
 input [7:0] Tile_X0Y0_E2END;
 input [7:0] Tile_X0Y0_E2MID;
 input [11:0] Tile_X0Y0_E6END;
 input [15:0] Tile_X0Y0_EE4END;
 input [31:0] Tile_X0Y0_FrameData;
 output [31:0] Tile_X0Y0_FrameData_O;
 output [19:0] Tile_X0Y0_FrameStrobe_O;
 output [3:0] Tile_X0Y0_N1BEG;
 output [7:0] Tile_X0Y0_N2BEG;
 output [7:0] Tile_X0Y0_N2BEGb;
 output [15:0] Tile_X0Y0_N4BEG;
 input [3:0] Tile_X0Y0_S1END;
 input [7:0] Tile_X0Y0_S2END;
 input [7:0] Tile_X0Y0_S2MID;
 input [15:0] Tile_X0Y0_S4END;
 output [3:0] Tile_X0Y0_W1BEG;
 output [7:0] Tile_X0Y0_W2BEG;
 output [7:0] Tile_X0Y0_W2BEGb;
 output [11:0] Tile_X0Y0_W6BEG;
 output [15:0] Tile_X0Y0_WW4BEG;
 input [3:0] Tile_X0Y1_E1END;
 input [7:0] Tile_X0Y1_E2END;
 input [7:0] Tile_X0Y1_E2MID;
 input [11:0] Tile_X0Y1_E6END;
 input [15:0] Tile_X0Y1_EE4END;
 input [31:0] Tile_X0Y1_FrameData;
 output [31:0] Tile_X0Y1_FrameData_O;
 input [19:0] Tile_X0Y1_FrameStrobe;
 input [3:0] Tile_X0Y1_N1END;
 input [7:0] Tile_X0Y1_N2END;
 input [7:0] Tile_X0Y1_N2MID;
 input [15:0] Tile_X0Y1_N4END;
 output [3:0] Tile_X0Y1_S1BEG;
 output [7:0] Tile_X0Y1_S2BEG;
 output [7:0] Tile_X0Y1_S2BEGb;
 output [15:0] Tile_X0Y1_S4BEG;
 output [3:0] Tile_X0Y1_W1BEG;
 output [7:0] Tile_X0Y1_W2BEG;
 output [7:0] Tile_X0Y1_W2BEGb;
 output [11:0] Tile_X0Y1_W6BEG;
 output [15:0] Tile_X0Y1_WW4BEG;

 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit0.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit1.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit10.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit11.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit12.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit13.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit14.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit15.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit16.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit17.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit18.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit19.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit2.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit20.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit21.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit22.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit23.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit24.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit25.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit26.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit27.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit28.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit29.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit3.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit30.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit31.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit4.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit5.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit6.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit7.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit8.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit9.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit0.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit1.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit10.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit11.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit12.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit13.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit14.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit15.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit16.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit17.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit18.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit19.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit2.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit20.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit21.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit22.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit23.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit24.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit25.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit26.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit27.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit28.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit29.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit3.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit30.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit31.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit4.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit5.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit6.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit7.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit8.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit9.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit0.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit1.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit10.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit11.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit12.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit13.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit14.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit15.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit16.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit17.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit18.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit19.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit2.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit20.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit21.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit22.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit23.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit24.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit25.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit26.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit27.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit28.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit29.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit3.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit30.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit31.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit4.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit5.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit6.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit7.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit8.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit9.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit0.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit1.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit10.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit11.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit12.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit13.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit14.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit15.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit16.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit17.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit18.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit19.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit2.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit20.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit21.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit22.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit23.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit24.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit25.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit26.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit27.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit28.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit29.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit3.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit30.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit31.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit4.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit5.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit6.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit7.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit8.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit9.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit0.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit1.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit10.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit11.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit12.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit13.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit14.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit15.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit16.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit17.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit18.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit19.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit2.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit20.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit21.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit22.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit23.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit24.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit25.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit26.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit27.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit28.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit29.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit3.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit30.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit31.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit4.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit5.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit6.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit7.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit8.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit9.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit0.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit1.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit10.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit11.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit12.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit13.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit14.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit15.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit16.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit17.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit18.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit19.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit2.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit20.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit21.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit22.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit23.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit24.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit25.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit26.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit27.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit28.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit29.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit3.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit30.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit31.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit4.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit5.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit6.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit7.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit8.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit9.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit0.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit1.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit10.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit11.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit12.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit13.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit14.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit15.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit16.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit17.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit18.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit19.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit2.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit20.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit21.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit22.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit23.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit24.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit25.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit26.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit27.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit28.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit29.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit3.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit30.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit31.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit4.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit5.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit6.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit7.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit8.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit9.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit10.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit11.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit12.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit13.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit14.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit15.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit16.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit17.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit18.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit19.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit20.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit21.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit22.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit23.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit24.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit25.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit26.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit27.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit28.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit29.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit30.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit31.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit8.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit9.Q ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG0 ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG1 ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG2 ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG3 ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG4 ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG5 ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG6 ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG7 ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG10 ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG11 ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG12 ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG13 ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG14 ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG15 ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG4 ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG5 ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG6 ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG7 ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG8 ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG9 ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N1BEG0 ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N1BEG1 ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N1BEG2 ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N1BEG3 ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N1END0 ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N1END1 ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N1END2 ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N1END3 ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N2BEG0 ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N2BEG1 ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N2BEG2 ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N2BEG3 ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N2BEG4 ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N2BEG5 ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N2BEG6 ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N2BEG7 ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N2BEGb0 ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N2BEGb1 ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N2BEGb2 ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N2BEGb3 ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N2BEGb4 ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N2BEGb5 ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N2BEGb6 ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N2BEGb7 ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N4BEG0 ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N4BEG1 ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N4BEG2 ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N4BEG3 ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.S2BEG0 ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.S2BEG1 ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.S2BEG2 ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.S2BEG3 ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.S2BEG4 ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.S2BEG5 ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.S2BEG6 ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.S2BEG7 ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.S4BEG0 ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.S4BEG1 ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.S4BEG2 ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.S4BEG3 ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W1BEG0 ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W1BEG1 ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W1BEG2 ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W1BEG3 ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W2BEG0 ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W2BEG1 ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W2BEG2 ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W2BEG3 ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W2BEG4 ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W2BEG5 ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W2BEG6 ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W2BEG7 ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W2BEGb0 ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W2BEGb1 ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W2BEGb2 ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W2BEGb3 ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W2BEGb4 ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W2BEGb5 ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W2BEGb6 ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W2BEGb7 ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W6BEG0 ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W6BEG1 ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W6BEG10 ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W6BEG11 ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W6BEG2 ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W6BEG3 ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W6BEG4 ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W6BEG5 ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W6BEG6 ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W6BEG7 ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W6BEG8 ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W6BEG9 ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.WW4BEG0 ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.WW4BEG1 ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.WW4BEG10 ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.WW4BEG11 ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.WW4BEG12 ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.WW4BEG13 ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.WW4BEG14 ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.WW4BEG15 ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.WW4BEG2 ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.WW4BEG3 ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.WW4BEG4 ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.WW4BEG5 ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.WW4BEG6 ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.WW4BEG7 ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.WW4BEG8 ;
 wire \Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.WW4BEG9 ;
 wire \Tile_X0Y0_E_TT_IF2_top.N4BEG_outbuf_10.A ;
 wire \Tile_X0Y0_E_TT_IF2_top.N4BEG_outbuf_11.A ;
 wire \Tile_X0Y0_E_TT_IF2_top.N4BEG_outbuf_8.A ;
 wire \Tile_X0Y0_E_TT_IF2_top.N4BEG_outbuf_9.A ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit0.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit1.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit10.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit11.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit12.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit13.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit14.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit15.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit16.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit17.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit18.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit19.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit2.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit20.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit21.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit22.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit23.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit24.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit25.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit26.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit27.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit28.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit29.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit3.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit30.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit31.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit4.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit5.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit6.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit7.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit8.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit9.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit0.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit1.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit10.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit11.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit12.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit13.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit14.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit15.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit16.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit17.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit18.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit19.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit2.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit20.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit21.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit22.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit23.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit24.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit25.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit26.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit27.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit28.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit29.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit3.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit30.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit31.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit4.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit5.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit6.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit7.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit8.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit9.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit0.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit1.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit10.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit11.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit12.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit13.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit14.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit15.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit16.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit17.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit18.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit19.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit2.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit20.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit21.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit22.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit23.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit24.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit25.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit26.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit27.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit28.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit29.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit3.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit30.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit31.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit4.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit5.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit6.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit7.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit8.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit9.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit0.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit1.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit10.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit11.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit12.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit13.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit14.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit15.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit16.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit17.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit18.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit19.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit2.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit20.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit21.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit22.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit23.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit24.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit25.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit26.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit27.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit28.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit29.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit3.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit30.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit31.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit4.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit5.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit6.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit7.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit8.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit9.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit0.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit1.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit10.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit11.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit12.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit13.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit14.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit15.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit16.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit17.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit18.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit19.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit2.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit20.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit21.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit22.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit23.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit24.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit25.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit26.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit27.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit28.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit29.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit3.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit30.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit31.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit4.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit5.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit6.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit7.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit8.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit9.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit0.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit1.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit10.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit11.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit12.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit13.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit14.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit15.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit16.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit17.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit18.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit19.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit2.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit20.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit21.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit22.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit23.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit24.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit25.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit26.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit27.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit28.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit29.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit3.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit30.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit31.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit4.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit5.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit6.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit7.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit8.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit9.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit0.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit1.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit10.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit11.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit12.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit13.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit14.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit15.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit16.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit17.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit18.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit19.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit2.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit20.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit21.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit22.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit23.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit24.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit25.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit26.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit27.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit28.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit29.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit3.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit30.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit31.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit4.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit5.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit6.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit7.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit8.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit9.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit0.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit1.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit10.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit11.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit12.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit13.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit14.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit15.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit16.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit17.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit18.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit19.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit2.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit20.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit21.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit22.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit23.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit24.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit25.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit26.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit27.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit28.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit29.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit3.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit30.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit31.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit4.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit5.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit6.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit7.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit8.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit9.Q ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.J_NS4_BEG12 ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.J_NS4_BEG13 ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.J_NS4_BEG14 ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.J_NS4_BEG15 ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.S1BEG0 ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.S1BEG1 ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.S1BEG2 ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.S1BEG3 ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.S2BEG0 ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.S2BEG1 ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.S2BEG2 ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.S2BEG3 ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.S2BEG4 ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.S2BEG5 ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.S2BEG6 ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.S2BEG7 ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.S4BEG0 ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.S4BEG1 ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.S4BEG2 ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.S4BEG3 ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W1BEG0 ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W1BEG1 ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W1BEG2 ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W1BEG3 ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W2BEG0 ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W2BEG1 ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W2BEG2 ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W2BEG3 ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W2BEG4 ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W2BEG5 ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W2BEG6 ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W2BEG7 ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W2BEGb0 ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W2BEGb1 ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W2BEGb2 ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W2BEGb3 ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W2BEGb4 ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W2BEGb5 ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W2BEGb6 ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W2BEGb7 ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W6BEG0 ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W6BEG1 ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W6BEG10 ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W6BEG11 ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W6BEG2 ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W6BEG3 ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W6BEG4 ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W6BEG5 ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W6BEG6 ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W6BEG7 ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W6BEG8 ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W6BEG9 ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.WW4BEG0 ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.WW4BEG1 ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.WW4BEG10 ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.WW4BEG11 ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.WW4BEG12 ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.WW4BEG13 ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.WW4BEG14 ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.WW4BEG15 ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.WW4BEG2 ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.WW4BEG3 ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.WW4BEG4 ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.WW4BEG5 ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.WW4BEG6 ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.WW4BEG7 ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.WW4BEG8 ;
 wire \Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.WW4BEG9 ;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire clknet_0_Tile_X0Y1_UserCLK;
 wire clknet_1_0__leaf_Tile_X0Y1_UserCLK;
 wire clknet_1_1__leaf_Tile_X0Y1_UserCLK;

 sg13g2_inv_1 _0357_ (.VDD(VPWR),
    .Y(_0287_),
    .A(Tile_X0Y0_E6END[1]),
    .VSS(VGND));
 sg13g2_inv_1 _0358_ (.VDD(VPWR),
    .Y(_0288_),
    .A(Tile_X0Y0_E6END[2]),
    .VSS(VGND));
 sg13g2_inv_1 _0359_ (.VDD(VPWR),
    .Y(_0289_),
    .A(Tile_X0Y0_E6END[3]),
    .VSS(VGND));
 sg13g2_inv_1 _0360_ (.VDD(VPWR),
    .Y(_0290_),
    .A(Tile_X0Y0_E6END[0]),
    .VSS(VGND));
 sg13g2_inv_1 _0361_ (.VDD(VPWR),
    .Y(_0291_),
    .A(Tile_X0Y0_E6END[8]),
    .VSS(VGND));
 sg13g2_inv_1 _0362_ (.VDD(VPWR),
    .Y(_0292_),
    .A(Tile_X0Y0_E6END[9]),
    .VSS(VGND));
 sg13g2_inv_1 _0363_ (.VDD(VPWR),
    .Y(_0293_),
    .A(Tile_X0Y0_E6END[10]),
    .VSS(VGND));
 sg13g2_inv_1 _0364_ (.VDD(VPWR),
    .Y(_0294_),
    .A(Tile_X0Y0_E6END[11]),
    .VSS(VGND));
 sg13g2_inv_1 _0365_ (.VDD(VPWR),
    .Y(_0295_),
    .A(Tile_X0Y1_E2END[5]),
    .VSS(VGND));
 sg13g2_inv_1 _0366_ (.VDD(VPWR),
    .Y(_0296_),
    .A(Tile_X0Y0_S2MID[3]),
    .VSS(VGND));
 sg13g2_inv_1 _0367_ (.VDD(VPWR),
    .Y(_0297_),
    .A(Tile_X0Y1_E6END[3]),
    .VSS(VGND));
 sg13g2_inv_1 _0368_ (.VDD(VPWR),
    .Y(_0298_),
    .A(Tile_X0Y1_E6END[2]),
    .VSS(VGND));
 sg13g2_inv_1 _0369_ (.VDD(VPWR),
    .Y(_0299_),
    .A(Tile_X0Y1_E6END[1]),
    .VSS(VGND));
 sg13g2_inv_1 _0370_ (.VDD(VPWR),
    .Y(_0300_),
    .A(Tile_X0Y1_E6END[0]),
    .VSS(VGND));
 sg13g2_inv_1 _0371_ (.VDD(VPWR),
    .Y(_0301_),
    .A(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit30.Q ),
    .VSS(VGND));
 sg13g2_inv_1 _0372_ (.VDD(VPWR),
    .Y(_0302_),
    .A(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit1.Q ),
    .VSS(VGND));
 sg13g2_inv_1 _0373_ (.VDD(VPWR),
    .Y(_0303_),
    .A(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit4.Q ),
    .VSS(VGND));
 sg13g2_inv_1 _0374_ (.VDD(VPWR),
    .Y(_0304_),
    .A(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit7.Q ),
    .VSS(VGND));
 sg13g2_inv_1 _0375_ (.VDD(VPWR),
    .Y(_0305_),
    .A(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit1.Q ),
    .VSS(VGND));
 sg13g2_inv_1 _0376_ (.VDD(VPWR),
    .Y(_0306_),
    .A(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit2.Q ),
    .VSS(VGND));
 sg13g2_inv_1 _0377_ (.VDD(VPWR),
    .Y(_0307_),
    .A(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit7.Q ),
    .VSS(VGND));
 sg13g2_nand2b_1 _0378_ (.Y(_0308_),
    .B(Tile_X0Y0_S1END[1]),
    .A_N(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit26.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _0379_ (.A(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit26.Q ),
    .B(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit27.Q ),
    .C(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N1END1 ),
    .Y(_0309_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _0380_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_0308_),
    .C1(_0309_),
    .B1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit27.Q ),
    .A1(_0287_),
    .Y(_0310_),
    .A2(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit26.Q ));
 sg13g2_mux4_1 _0381_ (.S0(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit14.Q ),
    .A0(Tile_X0Y0_E1END[1]),
    .A1(Tile_X0Y0_E6END[9]),
    .A2(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG13 ),
    .A3(_0310_),
    .S1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit15.Q ),
    .X(_0311_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _0382_ (.Y(_0312_),
    .B(_0311_),
    .A_N(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit26.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _0383_ (.A(Tile_X0Y1_N1END[1]),
    .B(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit26.Q ),
    .C(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit27.Q ),
    .Y(_0313_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _0384_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_0312_),
    .C1(_0313_),
    .B1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit27.Q ),
    .A1(_0299_),
    .Y(_0314_),
    .A2(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit26.Q ));
 sg13g2_mux4_1 _0385_ (.S0(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit3.Q ),
    .A0(Tile_X0Y1_E1END[1]),
    .A1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.J_NS4_BEG13 ),
    .A2(Tile_X0Y1_E6END[5]),
    .A3(_0314_),
    .S1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit2.Q ),
    .X(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N1END1 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0386_ (.S0(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit2.Q ),
    .A0(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N1END1 ),
    .A1(Tile_X0Y1_N4END[5]),
    .A2(Tile_X0Y0_S1END[1]),
    .A3(Tile_X0Y0_S4END[1]),
    .S1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit3.Q ),
    .X(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG13 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0387_ (.S0(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit10.Q ),
    .A0(Tile_X0Y0_E1END[1]),
    .A1(Tile_X0Y0_E6END[5]),
    .A2(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG13 ),
    .A3(_0310_),
    .S1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit11.Q ),
    .X(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N1BEG1 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _0388_ (.Y(_0315_),
    .B(Tile_X0Y0_S1END[2]),
    .A_N(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit28.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _0389_ (.A(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit28.Q ),
    .B(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit29.Q ),
    .C(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N1END2 ),
    .Y(_0316_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _0390_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_0315_),
    .C1(_0316_),
    .B1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit29.Q ),
    .A1(_0288_),
    .Y(_0317_),
    .A2(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit28.Q ));
 sg13g2_mux4_1 _0391_ (.S0(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit16.Q ),
    .A0(Tile_X0Y0_E1END[2]),
    .A1(Tile_X0Y0_E6END[10]),
    .A2(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG14 ),
    .A3(_0317_),
    .S1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit17.Q ),
    .X(_0318_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _0392_ (.Y(_0319_),
    .B(_0318_),
    .A_N(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit28.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _0393_ (.A(Tile_X0Y1_N1END[2]),
    .B(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit28.Q ),
    .C(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit29.Q ),
    .Y(_0320_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _0394_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_0319_),
    .C1(_0320_),
    .B1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit29.Q ),
    .A1(_0298_),
    .Y(_0321_),
    .A2(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit28.Q ));
 sg13g2_mux4_1 _0395_ (.S0(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit5.Q ),
    .A0(Tile_X0Y1_E1END[2]),
    .A1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.J_NS4_BEG14 ),
    .A2(Tile_X0Y1_E6END[6]),
    .A3(_0321_),
    .S1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit4.Q ),
    .X(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N1END2 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0396_ (.S0(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit4.Q ),
    .A0(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N1END2 ),
    .A1(Tile_X0Y1_N4END[6]),
    .A2(Tile_X0Y0_S1END[2]),
    .A3(Tile_X0Y0_S4END[2]),
    .S1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit5.Q ),
    .X(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG14 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0397_ (.S0(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit12.Q ),
    .A0(Tile_X0Y0_E1END[2]),
    .A1(Tile_X0Y0_E6END[6]),
    .A2(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG14 ),
    .A3(_0317_),
    .S1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit13.Q ),
    .X(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N1BEG2 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _0398_ (.Y(_0322_),
    .B(Tile_X0Y0_S1END[3]),
    .A_N(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit30.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _0399_ (.A(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit30.Q ),
    .B(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit31.Q ),
    .C(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N1END3 ),
    .Y(_0323_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _0400_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_0322_),
    .C1(_0323_),
    .B1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit31.Q ),
    .A1(_0289_),
    .Y(_0324_),
    .A2(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit30.Q ));
 sg13g2_mux4_1 _0401_ (.S0(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit18.Q ),
    .A0(Tile_X0Y0_E1END[3]),
    .A1(Tile_X0Y0_E6END[11]),
    .A2(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG15 ),
    .A3(_0324_),
    .S1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit19.Q ),
    .X(_0325_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _0402_ (.Y(_0326_),
    .B(_0325_),
    .A_N(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit30.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _0403_ (.A(Tile_X0Y1_N1END[3]),
    .B(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit30.Q ),
    .C(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit31.Q ),
    .Y(_0327_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _0404_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_0326_),
    .C1(_0327_),
    .B1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit31.Q ),
    .A1(_0297_),
    .Y(_0328_),
    .A2(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit30.Q ));
 sg13g2_mux4_1 _0405_ (.S0(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit7.Q ),
    .A0(Tile_X0Y1_E1END[3]),
    .A1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.J_NS4_BEG15 ),
    .A2(Tile_X0Y1_E6END[7]),
    .A3(_0328_),
    .S1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit6.Q ),
    .X(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N1END3 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0406_ (.S0(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit6.Q ),
    .A0(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N1END3 ),
    .A1(Tile_X0Y1_N4END[7]),
    .A2(Tile_X0Y0_S1END[3]),
    .A3(Tile_X0Y0_S4END[3]),
    .S1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit7.Q ),
    .X(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG15 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0407_ (.S0(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit14.Q ),
    .A0(Tile_X0Y0_E1END[3]),
    .A1(Tile_X0Y0_E6END[7]),
    .A2(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG15 ),
    .A3(_0324_),
    .S1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit15.Q ),
    .X(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N1BEG3 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0408_ (.S0(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit20.Q ),
    .A0(Tile_X0Y0_E2MID[7]),
    .A1(Tile_X0Y0_E2END[7]),
    .A2(Tile_X0Y0_E6END[8]),
    .A3(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG0 ),
    .S1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit21.Q ),
    .X(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.S2BEG0 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _0409_ (.A0(Tile_X0Y1_N2MID[0]),
    .A1(Tile_X0Y1_N2END[0]),
    .S(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit8.Q ),
    .X(_0329_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _0410_ (.A(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit9.Q ),
    .B(_0329_),
    .Y(_0330_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _0411_ (.Y(_0331_),
    .B(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.S2BEG0 ),
    .A_N(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit8.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _0412_ (.Y(_0332_),
    .A(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit8.Q ),
    .B(Tile_X0Y0_S2MID[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _0413_ (.B(_0331_),
    .C(_0332_),
    .A(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit9.Q ),
    .Y(_0333_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _0414_ (.Y(_0334_),
    .B(_0333_),
    .A_N(_0330_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _0415_ (.A(_0330_),
    .B_N(_0333_),
    .Y(_0335_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0416_ (.S0(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit8.Q ),
    .A0(Tile_X0Y1_E2MID[7]),
    .A1(Tile_X0Y1_E2END[7]),
    .A2(Tile_X0Y1_E6END[7]),
    .A3(_0335_),
    .S1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit9.Q ),
    .X(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N2BEGb0 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0417_ (.S0(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit9.Q ),
    .A0(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N2BEGb0 ),
    .A1(Tile_X0Y0_S2MID[0]),
    .A2(Tile_X0Y1_N2MID[0]),
    .A3(Tile_X0Y0_S2END[0]),
    .S1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit8.Q ),
    .X(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG0 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0418_ (.S0(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit16.Q ),
    .A0(Tile_X0Y0_E2MID[7]),
    .A1(Tile_X0Y0_E2END[7]),
    .A2(Tile_X0Y0_E6END[7]),
    .A3(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG0 ),
    .S1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit17.Q ),
    .X(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N2BEG0 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0419_ (.S0(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit22.Q ),
    .A0(Tile_X0Y0_E2MID[6]),
    .A1(Tile_X0Y0_E2END[6]),
    .A2(Tile_X0Y0_E6END[9]),
    .A3(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG1 ),
    .S1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit23.Q ),
    .X(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.S2BEG1 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _0420_ (.A0(Tile_X0Y1_N2MID[1]),
    .A1(Tile_X0Y1_N2END[1]),
    .S(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit10.Q ),
    .X(_0336_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _0421_ (.A(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit11.Q ),
    .B(_0336_),
    .Y(_0337_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _0422_ (.Y(_0338_),
    .B(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.S2BEG1 ),
    .A_N(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit10.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _0423_ (.Y(_0339_),
    .A(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit10.Q ),
    .B(Tile_X0Y0_S2MID[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _0424_ (.B(_0338_),
    .C(_0339_),
    .A(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit11.Q ),
    .Y(_0340_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _0425_ (.Y(_0341_),
    .B(_0340_),
    .A_N(_0337_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _0426_ (.A(_0337_),
    .B_N(_0340_),
    .Y(_0342_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0427_ (.S0(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit10.Q ),
    .A0(Tile_X0Y1_E2MID[6]),
    .A1(Tile_X0Y1_E2END[6]),
    .A2(Tile_X0Y1_E6END[6]),
    .A3(_0342_),
    .S1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit11.Q ),
    .X(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N2BEGb1 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0428_ (.S0(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit11.Q ),
    .A0(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N2BEGb1 ),
    .A1(Tile_X0Y0_S2MID[1]),
    .A2(Tile_X0Y1_N2MID[1]),
    .A3(Tile_X0Y0_S2END[1]),
    .S1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit10.Q ),
    .X(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG1 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0429_ (.S0(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit18.Q ),
    .A0(Tile_X0Y0_E2MID[6]),
    .A1(Tile_X0Y0_E2END[6]),
    .A2(Tile_X0Y0_E6END[6]),
    .A3(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG1 ),
    .S1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit19.Q ),
    .X(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N2BEG1 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0430_ (.S0(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit24.Q ),
    .A0(Tile_X0Y0_E2MID[5]),
    .A1(Tile_X0Y0_E2END[5]),
    .A2(Tile_X0Y0_E6END[10]),
    .A3(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG2 ),
    .S1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit25.Q ),
    .X(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.S2BEG2 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _0431_ (.A0(Tile_X0Y1_N2MID[2]),
    .A1(Tile_X0Y1_N2END[2]),
    .S(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit12.Q ),
    .X(_0343_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _0432_ (.A(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit13.Q ),
    .B(_0343_),
    .Y(_0344_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _0433_ (.Y(_0345_),
    .B(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.S2BEG2 ),
    .A_N(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit12.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _0434_ (.Y(_0346_),
    .A(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit12.Q ),
    .B(Tile_X0Y0_S2MID[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _0435_ (.B(_0345_),
    .C(_0346_),
    .A(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit13.Q ),
    .Y(_0347_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _0436_ (.Y(_0348_),
    .B(_0347_),
    .A_N(_0344_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _0437_ (.A(_0344_),
    .B_N(_0347_),
    .Y(_0349_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0438_ (.S0(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit12.Q ),
    .A0(Tile_X0Y1_E2MID[5]),
    .A1(Tile_X0Y1_E2END[5]),
    .A2(Tile_X0Y1_E6END[5]),
    .A3(_0349_),
    .S1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit13.Q ),
    .X(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N2BEGb2 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0439_ (.S0(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit13.Q ),
    .A0(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N2BEGb2 ),
    .A1(Tile_X0Y0_S2MID[2]),
    .A2(Tile_X0Y1_N2MID[2]),
    .A3(Tile_X0Y0_S2END[2]),
    .S1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit12.Q ),
    .X(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG2 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0440_ (.S0(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit20.Q ),
    .A0(Tile_X0Y0_E2MID[5]),
    .A1(Tile_X0Y0_E2END[5]),
    .A2(Tile_X0Y0_E6END[5]),
    .A3(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG2 ),
    .S1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit21.Q ),
    .X(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N2BEG2 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0441_ (.S0(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit26.Q ),
    .A0(Tile_X0Y0_E2MID[4]),
    .A1(Tile_X0Y0_E2END[4]),
    .A2(Tile_X0Y0_E6END[11]),
    .A3(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG3 ),
    .S1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit27.Q ),
    .X(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.S2BEG3 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _0442_ (.A0(Tile_X0Y1_N2MID[3]),
    .A1(Tile_X0Y1_N2END[3]),
    .S(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit14.Q ),
    .X(_0350_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _0443_ (.A(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit15.Q ),
    .B(_0350_),
    .Y(_0351_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _0444_ (.Y(_0352_),
    .B(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.S2BEG3 ),
    .A_N(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit14.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _0445_ (.Y(_0353_),
    .A(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit14.Q ),
    .B(Tile_X0Y0_S2MID[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _0446_ (.B(_0352_),
    .C(_0353_),
    .A(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit15.Q ),
    .Y(_0354_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _0447_ (.Y(_0355_),
    .B(_0354_),
    .A_N(_0351_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _0448_ (.A(_0351_),
    .B_N(_0354_),
    .Y(_0356_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0449_ (.S0(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit14.Q ),
    .A0(Tile_X0Y1_E2MID[4]),
    .A1(Tile_X0Y1_E2END[4]),
    .A2(Tile_X0Y1_E6END[4]),
    .A3(_0356_),
    .S1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit15.Q ),
    .X(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N2BEGb3 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0450_ (.S0(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit15.Q ),
    .A0(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N2BEGb3 ),
    .A1(Tile_X0Y0_S2MID[3]),
    .A2(Tile_X0Y1_N2MID[3]),
    .A3(Tile_X0Y0_S2END[3]),
    .S1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit14.Q ),
    .X(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG3 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0451_ (.S0(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit22.Q ),
    .A0(Tile_X0Y0_E2MID[4]),
    .A1(Tile_X0Y0_E2END[4]),
    .A2(Tile_X0Y0_E6END[4]),
    .A3(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG3 ),
    .S1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit23.Q ),
    .X(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N2BEG3 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0452_ (.S0(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit29.Q ),
    .A0(Tile_X0Y0_E1END[0]),
    .A1(Tile_X0Y0_E2END[3]),
    .A2(Tile_X0Y0_E2MID[3]),
    .A3(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG4 ),
    .S1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit28.Q ),
    .X(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.S2BEG4 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0453_ (.S0(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit16.Q ),
    .A0(Tile_X0Y1_N2MID[4]),
    .A1(Tile_X0Y1_N2END[4]),
    .A2(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.S2BEG4 ),
    .A3(Tile_X0Y0_S2MID[4]),
    .S1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit17.Q ),
    .X(_0000_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0454_ (.S0(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit16.Q ),
    .A0(Tile_X0Y1_E2MID[3]),
    .A1(Tile_X0Y1_E2END[3]),
    .A2(Tile_X0Y1_E6END[3]),
    .A3(_0000_),
    .S1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit17.Q ),
    .X(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N2BEGb4 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0455_ (.S0(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit17.Q ),
    .A0(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N2BEGb4 ),
    .A1(Tile_X0Y0_S2MID[4]),
    .A2(Tile_X0Y1_N2MID[4]),
    .A3(Tile_X0Y0_S2END[4]),
    .S1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit16.Q ),
    .X(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG4 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0456_ (.S0(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit24.Q ),
    .A0(Tile_X0Y0_E2MID[3]),
    .A1(Tile_X0Y0_E2END[3]),
    .A2(Tile_X0Y0_E6END[3]),
    .A3(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG4 ),
    .S1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit25.Q ),
    .X(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N2BEG4 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0457_ (.S0(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit30.Q ),
    .A0(Tile_X0Y0_E1END[1]),
    .A1(Tile_X0Y0_E2MID[2]),
    .A2(Tile_X0Y0_E2END[2]),
    .A3(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG5 ),
    .S1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit31.Q ),
    .X(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.S2BEG5 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0458_ (.S0(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit18.Q ),
    .A0(Tile_X0Y1_N2MID[5]),
    .A1(Tile_X0Y1_N2END[5]),
    .A2(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.S2BEG5 ),
    .A3(Tile_X0Y0_S2MID[5]),
    .S1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit19.Q ),
    .X(_0001_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0459_ (.S0(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit18.Q ),
    .A0(Tile_X0Y1_E2MID[2]),
    .A1(Tile_X0Y1_E2END[2]),
    .A2(Tile_X0Y1_E6END[2]),
    .A3(_0001_),
    .S1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit19.Q ),
    .X(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N2BEGb5 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0460_ (.S0(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit19.Q ),
    .A0(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N2BEGb5 ),
    .A1(Tile_X0Y0_S2MID[5]),
    .A2(Tile_X0Y1_N2MID[5]),
    .A3(Tile_X0Y0_S2END[5]),
    .S1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit18.Q ),
    .X(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG5 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0461_ (.S0(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit26.Q ),
    .A0(Tile_X0Y0_E2MID[2]),
    .A1(Tile_X0Y0_E2END[2]),
    .A2(Tile_X0Y0_E6END[2]),
    .A3(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG5 ),
    .S1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit27.Q ),
    .X(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N2BEG5 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0462_ (.S0(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit0.Q ),
    .A0(Tile_X0Y0_E1END[2]),
    .A1(Tile_X0Y0_E2MID[1]),
    .A2(Tile_X0Y0_E2END[1]),
    .A3(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG6 ),
    .S1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit1.Q ),
    .X(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.S2BEG6 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0463_ (.S0(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit20.Q ),
    .A0(Tile_X0Y1_N2MID[6]),
    .A1(Tile_X0Y1_N2END[6]),
    .A2(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.S2BEG6 ),
    .A3(Tile_X0Y0_S2MID[6]),
    .S1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit21.Q ),
    .X(_0002_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0464_ (.S0(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit20.Q ),
    .A0(Tile_X0Y1_E2MID[1]),
    .A1(Tile_X0Y1_E2END[1]),
    .A2(Tile_X0Y1_E6END[1]),
    .A3(_0002_),
    .S1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit21.Q ),
    .X(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N2BEGb6 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0465_ (.S0(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit21.Q ),
    .A0(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N2BEGb6 ),
    .A1(Tile_X0Y0_S2MID[6]),
    .A2(Tile_X0Y1_N2MID[6]),
    .A3(Tile_X0Y0_S2END[6]),
    .S1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit20.Q ),
    .X(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG6 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0466_ (.S0(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit28.Q ),
    .A0(Tile_X0Y0_E2MID[1]),
    .A1(Tile_X0Y0_E2END[1]),
    .A2(Tile_X0Y0_E6END[1]),
    .A3(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG6 ),
    .S1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit29.Q ),
    .X(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N2BEG6 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0467_ (.S0(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit2.Q ),
    .A0(Tile_X0Y0_E1END[3]),
    .A1(Tile_X0Y0_E2MID[0]),
    .A2(Tile_X0Y0_E2END[0]),
    .A3(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG7 ),
    .S1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit3.Q ),
    .X(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.S2BEG7 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0468_ (.S0(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit22.Q ),
    .A0(Tile_X0Y1_N2MID[7]),
    .A1(Tile_X0Y1_N2END[7]),
    .A2(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.S2BEG7 ),
    .A3(Tile_X0Y0_S2MID[7]),
    .S1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit23.Q ),
    .X(_0003_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0469_ (.S0(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit22.Q ),
    .A0(Tile_X0Y1_E2MID[0]),
    .A1(Tile_X0Y1_E2END[0]),
    .A2(Tile_X0Y1_E6END[0]),
    .A3(_0003_),
    .S1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit23.Q ),
    .X(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N2BEGb7 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0470_ (.S0(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit23.Q ),
    .A0(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N2BEGb7 ),
    .A1(Tile_X0Y0_S2MID[7]),
    .A2(Tile_X0Y1_N2MID[7]),
    .A3(Tile_X0Y0_S2END[7]),
    .S1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit22.Q ),
    .X(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG7 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0471_ (.S0(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit30.Q ),
    .A0(Tile_X0Y0_E2MID[0]),
    .A1(Tile_X0Y0_E2END[0]),
    .A2(Tile_X0Y0_E6END[0]),
    .A3(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG7 ),
    .S1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit31.Q ),
    .X(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N2BEG7 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _0472_ (.Y(_0004_),
    .B(Tile_X0Y0_S1END[0]),
    .A_N(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit24.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _0473_ (.A(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit24.Q ),
    .B(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit25.Q ),
    .C(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N1END0 ),
    .Y(_0005_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _0474_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_0004_),
    .C1(_0005_),
    .B1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit25.Q ),
    .A1(_0290_),
    .Y(_0006_),
    .A2(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit24.Q ));
 sg13g2_mux4_1 _0475_ (.S0(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit13.Q ),
    .A0(Tile_X0Y0_E1END[0]),
    .A1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG12 ),
    .A2(Tile_X0Y0_E6END[8]),
    .A3(_0006_),
    .S1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit12.Q ),
    .X(_0007_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _0476_ (.Y(_0008_),
    .B(_0007_),
    .A_N(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit24.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _0477_ (.A(Tile_X0Y1_N1END[0]),
    .B(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit24.Q ),
    .C(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit25.Q ),
    .Y(_0009_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _0478_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_0008_),
    .C1(_0009_),
    .B1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit25.Q ),
    .A1(_0300_),
    .Y(_0010_),
    .A2(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit24.Q ));
 sg13g2_mux4_1 _0479_ (.S0(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit1.Q ),
    .A0(Tile_X0Y1_E1END[0]),
    .A1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.J_NS4_BEG12 ),
    .A2(Tile_X0Y1_E6END[4]),
    .A3(_0010_),
    .S1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit0.Q ),
    .X(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N1END0 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0480_ (.S0(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit17.Q ),
    .A0(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N1END0 ),
    .A1(UIO_OUT_TT_PROJECT2),
    .A2(Tile_X0Y0_S1END[0]),
    .A3(UIO_OUT_TT_PROJECT7),
    .S1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit16.Q ),
    .X(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W1BEG0 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0481_ (.S0(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit19.Q ),
    .A0(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N1END1 ),
    .A1(UIO_OUT_TT_PROJECT3),
    .A2(Tile_X0Y0_S1END[1]),
    .A3(UIO_OUT_TT_PROJECT6),
    .S1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit18.Q ),
    .X(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W1BEG1 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0482_ (.S0(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit21.Q ),
    .A0(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N1END2 ),
    .A1(UIO_OUT_TT_PROJECT0),
    .A2(Tile_X0Y0_S1END[2]),
    .A3(UIO_OUT_TT_PROJECT5),
    .S1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit20.Q ),
    .X(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W1BEG2 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0483_ (.S0(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit23.Q ),
    .A0(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N1END3 ),
    .A1(UIO_OUT_TT_PROJECT1),
    .A2(Tile_X0Y0_S1END[3]),
    .A3(UIO_OUT_TT_PROJECT4),
    .S1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit22.Q ),
    .X(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W1BEG3 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0484_ (.S0(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit24.Q ),
    .A0(UIO_OUT_TT_PROJECT0),
    .A1(UIO_OE_TT_PROJECT0),
    .A2(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG0 ),
    .A3(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG7 ),
    .S1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit25.Q ),
    .X(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W2BEG0 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0485_ (.S0(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit26.Q ),
    .A0(UIO_OUT_TT_PROJECT1),
    .A1(UIO_OE_TT_PROJECT1),
    .A2(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG1 ),
    .A3(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG6 ),
    .S1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit27.Q ),
    .X(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W2BEG1 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0486_ (.S0(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit28.Q ),
    .A0(UIO_OUT_TT_PROJECT2),
    .A1(UIO_OE_TT_PROJECT2),
    .A2(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG2 ),
    .A3(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG5 ),
    .S1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit29.Q ),
    .X(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W2BEG2 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0487_ (.S0(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit30.Q ),
    .A0(UIO_OUT_TT_PROJECT3),
    .A1(UIO_OE_TT_PROJECT3),
    .A2(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG3 ),
    .A3(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG4 ),
    .S1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit31.Q ),
    .X(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W2BEG3 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0488_ (.S0(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit0.Q ),
    .A0(UIO_OUT_TT_PROJECT4),
    .A1(UIO_OE_TT_PROJECT4),
    .A2(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG3 ),
    .A3(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG4 ),
    .S1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit1.Q ),
    .X(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W2BEG4 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0489_ (.S0(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit2.Q ),
    .A0(UIO_OUT_TT_PROJECT5),
    .A1(UIO_OE_TT_PROJECT5),
    .A2(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG2 ),
    .A3(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG5 ),
    .S1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit3.Q ),
    .X(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W2BEG5 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0490_ (.S0(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit4.Q ),
    .A0(UIO_OUT_TT_PROJECT6),
    .A1(UIO_OE_TT_PROJECT6),
    .A2(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG1 ),
    .A3(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG6 ),
    .S1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit5.Q ),
    .X(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W2BEG6 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0491_ (.S0(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit6.Q ),
    .A0(UIO_OUT_TT_PROJECT7),
    .A1(UIO_OE_TT_PROJECT7),
    .A2(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG0 ),
    .A3(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG7 ),
    .S1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit7.Q ),
    .X(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W2BEG7 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0492_ (.S0(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit8.Q ),
    .A0(UIO_OUT_TT_PROJECT0),
    .A1(UIO_OE_TT_PROJECT0),
    .A2(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG0 ),
    .A3(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG7 ),
    .S1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit9.Q ),
    .X(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W2BEGb0 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0493_ (.S0(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit10.Q ),
    .A0(UIO_OUT_TT_PROJECT1),
    .A1(UIO_OE_TT_PROJECT1),
    .A2(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG1 ),
    .A3(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG6 ),
    .S1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit11.Q ),
    .X(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W2BEGb1 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0494_ (.S0(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit12.Q ),
    .A0(UIO_OUT_TT_PROJECT2),
    .A1(UIO_OE_TT_PROJECT2),
    .A2(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG2 ),
    .A3(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG5 ),
    .S1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit13.Q ),
    .X(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W2BEGb2 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0495_ (.S0(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit14.Q ),
    .A0(UIO_OUT_TT_PROJECT3),
    .A1(UIO_OE_TT_PROJECT3),
    .A2(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG3 ),
    .A3(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG4 ),
    .S1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit15.Q ),
    .X(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W2BEGb3 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0496_ (.S0(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit16.Q ),
    .A0(UIO_OUT_TT_PROJECT4),
    .A1(UIO_OE_TT_PROJECT4),
    .A2(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG3 ),
    .A3(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG4 ),
    .S1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit17.Q ),
    .X(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W2BEGb4 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0497_ (.S0(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit18.Q ),
    .A0(UIO_OUT_TT_PROJECT5),
    .A1(UIO_OE_TT_PROJECT5),
    .A2(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG2 ),
    .A3(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG5 ),
    .S1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit19.Q ),
    .X(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W2BEGb5 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0498_ (.S0(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit20.Q ),
    .A0(UIO_OUT_TT_PROJECT6),
    .A1(UIO_OE_TT_PROJECT6),
    .A2(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG1 ),
    .A3(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG6 ),
    .S1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit21.Q ),
    .X(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W2BEGb6 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0499_ (.S0(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit22.Q ),
    .A0(UIO_OUT_TT_PROJECT7),
    .A1(UIO_OE_TT_PROJECT7),
    .A2(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG0 ),
    .A3(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG7 ),
    .S1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit23.Q ),
    .X(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W2BEGb7 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0500_ (.S0(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit24.Q ),
    .A0(UIO_OUT_TT_PROJECT0),
    .A1(UIO_OE_TT_PROJECT4),
    .A2(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG15 ),
    .A3(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG7 ),
    .S1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit25.Q ),
    .X(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.WW4BEG0 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0501_ (.S0(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit26.Q ),
    .A0(UIO_OUT_TT_PROJECT1),
    .A1(UIO_OE_TT_PROJECT5),
    .A2(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG14 ),
    .A3(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG6 ),
    .S1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit27.Q ),
    .X(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.WW4BEG1 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0502_ (.S0(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit28.Q ),
    .A0(UIO_OUT_TT_PROJECT2),
    .A1(UIO_OE_TT_PROJECT6),
    .A2(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG13 ),
    .A3(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG5 ),
    .S1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit29.Q ),
    .X(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.WW4BEG2 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0503_ (.S0(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit0.Q ),
    .A0(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N1END0 ),
    .A1(Tile_X0Y1_N4END[4]),
    .A2(Tile_X0Y0_S1END[0]),
    .A3(Tile_X0Y0_S4END[0]),
    .S1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit1.Q ),
    .X(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG12 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0504_ (.S0(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit30.Q ),
    .A0(UIO_OUT_TT_PROJECT3),
    .A1(UIO_OE_TT_PROJECT7),
    .A2(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG12 ),
    .A3(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG4 ),
    .S1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit31.Q ),
    .X(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.WW4BEG3 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0505_ (.S0(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit30.Q ),
    .A0(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N1END3 ),
    .A1(Tile_X0Y1_N4END[7]),
    .A2(Tile_X0Y0_S1END[3]),
    .A3(Tile_X0Y0_S4END[3]),
    .S1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit31.Q ),
    .X(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG11 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0506_ (.S0(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit0.Q ),
    .A0(UIO_OUT_TT_PROJECT4),
    .A1(UIO_OE_TT_PROJECT0),
    .A2(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG11 ),
    .A3(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG3 ),
    .S1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit1.Q ),
    .X(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.WW4BEG4 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0507_ (.S0(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit28.Q ),
    .A0(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N1END2 ),
    .A1(Tile_X0Y1_N4END[6]),
    .A2(Tile_X0Y0_S1END[2]),
    .A3(Tile_X0Y0_S4END[2]),
    .S1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit29.Q ),
    .X(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG10 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0508_ (.S0(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit2.Q ),
    .A0(UIO_OUT_TT_PROJECT5),
    .A1(UIO_OE_TT_PROJECT0),
    .A2(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG10 ),
    .A3(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG2 ),
    .S1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit3.Q ),
    .X(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.WW4BEG5 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0509_ (.S0(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit26.Q ),
    .A0(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N1END1 ),
    .A1(Tile_X0Y1_N4END[5]),
    .A2(Tile_X0Y0_S1END[1]),
    .A3(Tile_X0Y0_S4END[1]),
    .S1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit27.Q ),
    .X(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG9 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0510_ (.S0(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit4.Q ),
    .A0(UIO_OUT_TT_PROJECT6),
    .A1(UIO_OE_TT_PROJECT2),
    .A2(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG9 ),
    .A3(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG1 ),
    .S1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit5.Q ),
    .X(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.WW4BEG6 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0511_ (.S0(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit24.Q ),
    .A0(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N1END0 ),
    .A1(Tile_X0Y1_N4END[4]),
    .A2(Tile_X0Y0_S1END[0]),
    .A3(Tile_X0Y0_S4END[0]),
    .S1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit25.Q ),
    .X(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG8 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0512_ (.S0(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit6.Q ),
    .A0(UIO_OUT_TT_PROJECT7),
    .A1(UIO_OE_TT_PROJECT3),
    .A2(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG8 ),
    .A3(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG0 ),
    .S1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit7.Q ),
    .X(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.WW4BEG7 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0513_ (.S0(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit22.Q ),
    .A0(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N1END3 ),
    .A1(Tile_X0Y1_N4END[7]),
    .A2(Tile_X0Y0_S1END[3]),
    .A3(Tile_X0Y0_S4END[3]),
    .S1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit23.Q ),
    .X(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG7 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0514_ (.S0(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit8.Q ),
    .A0(UIO_OUT_TT_PROJECT4),
    .A1(UIO_OE_TT_PROJECT0),
    .A2(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG7 ),
    .A3(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG7 ),
    .S1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit9.Q ),
    .X(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.WW4BEG8 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0515_ (.S0(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit20.Q ),
    .A0(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N1END2 ),
    .A1(Tile_X0Y1_N4END[6]),
    .A2(Tile_X0Y0_S1END[2]),
    .A3(Tile_X0Y0_S4END[2]),
    .S1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit21.Q ),
    .X(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG6 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0516_ (.S0(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit10.Q ),
    .A0(UIO_OUT_TT_PROJECT5),
    .A1(UIO_OE_TT_PROJECT1),
    .A2(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG6 ),
    .A3(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG6 ),
    .S1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit11.Q ),
    .X(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.WW4BEG9 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0517_ (.S0(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit18.Q ),
    .A0(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N1END1 ),
    .A1(Tile_X0Y1_N4END[5]),
    .A2(Tile_X0Y0_S1END[1]),
    .A3(Tile_X0Y0_S4END[1]),
    .S1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit19.Q ),
    .X(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG5 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0518_ (.S0(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit12.Q ),
    .A0(UIO_OUT_TT_PROJECT6),
    .A1(UIO_OE_TT_PROJECT2),
    .A2(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG5 ),
    .A3(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG5 ),
    .S1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit13.Q ),
    .X(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.WW4BEG10 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0519_ (.S0(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit16.Q ),
    .A0(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N1END0 ),
    .A1(Tile_X0Y1_N4END[4]),
    .A2(Tile_X0Y0_S1END[0]),
    .A3(Tile_X0Y0_S4END[0]),
    .S1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit17.Q ),
    .X(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG4 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0520_ (.S0(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit14.Q ),
    .A0(UIO_OUT_TT_PROJECT7),
    .A1(UIO_OE_TT_PROJECT3),
    .A2(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG4 ),
    .A3(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG4 ),
    .S1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit15.Q ),
    .X(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.WW4BEG11 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0521_ (.S0(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit14.Q ),
    .A0(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N1END3 ),
    .A1(Tile_X0Y1_N4END[7]),
    .A2(Tile_X0Y0_S1END[3]),
    .A3(Tile_X0Y0_S4END[3]),
    .S1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit15.Q ),
    .X(_0011_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0522_ (.S0(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit16.Q ),
    .A0(UIO_OUT_TT_PROJECT0),
    .A1(UIO_OE_TT_PROJECT4),
    .A2(_0011_),
    .A3(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG3 ),
    .S1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit17.Q ),
    .X(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.WW4BEG12 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0523_ (.S0(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit12.Q ),
    .A0(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N1END2 ),
    .A1(Tile_X0Y1_N4END[6]),
    .A2(Tile_X0Y0_S1END[2]),
    .A3(Tile_X0Y0_S4END[2]),
    .S1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit13.Q ),
    .X(_0012_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0524_ (.S0(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit18.Q ),
    .A0(UIO_OUT_TT_PROJECT1),
    .A1(UIO_OE_TT_PROJECT5),
    .A2(_0012_),
    .A3(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG2 ),
    .S1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit19.Q ),
    .X(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.WW4BEG13 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0525_ (.S0(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit10.Q ),
    .A0(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N1END1 ),
    .A1(Tile_X0Y1_N4END[5]),
    .A2(Tile_X0Y0_S1END[1]),
    .A3(Tile_X0Y0_S4END[1]),
    .S1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit11.Q ),
    .X(_0013_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0526_ (.S0(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit20.Q ),
    .A0(UIO_OUT_TT_PROJECT2),
    .A1(UIO_OE_TT_PROJECT6),
    .A2(_0013_),
    .A3(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG1 ),
    .S1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit21.Q ),
    .X(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.WW4BEG14 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0527_ (.S0(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit8.Q ),
    .A0(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N1END0 ),
    .A1(Tile_X0Y1_N4END[4]),
    .A2(Tile_X0Y0_S1END[0]),
    .A3(Tile_X0Y0_S4END[0]),
    .S1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit9.Q ),
    .X(_0014_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0528_ (.S0(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit22.Q ),
    .A0(UIO_OUT_TT_PROJECT3),
    .A1(UIO_OE_TT_PROJECT7),
    .A2(_0014_),
    .A3(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG0 ),
    .S1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit23.Q ),
    .X(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.WW4BEG15 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0529_ (.S0(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit24.Q ),
    .A0(Tile_X0Y1_N4END[4]),
    .A1(Tile_X0Y0_S4END[0]),
    .A2(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG11 ),
    .A3(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG15 ),
    .S1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit25.Q ),
    .X(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W6BEG0 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0530_ (.S0(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit26.Q ),
    .A0(Tile_X0Y1_N4END[5]),
    .A1(Tile_X0Y0_S4END[1]),
    .A2(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG10 ),
    .A3(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG14 ),
    .S1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit27.Q ),
    .X(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W6BEG1 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0531_ (.S0(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit28.Q ),
    .A0(Tile_X0Y1_N4END[6]),
    .A1(Tile_X0Y0_S4END[2]),
    .A2(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG9 ),
    .A3(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG13 ),
    .S1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit29.Q ),
    .X(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W6BEG2 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0532_ (.S0(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit30.Q ),
    .A0(Tile_X0Y1_N4END[7]),
    .A1(Tile_X0Y0_S4END[3]),
    .A2(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG8 ),
    .A3(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG12 ),
    .S1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit31.Q ),
    .X(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W6BEG3 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0533_ (.S0(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit1.Q ),
    .A0(UIO_OUT_TT_PROJECT4),
    .A1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG11 ),
    .A2(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG7 ),
    .A3(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG0 ),
    .S1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit0.Q ),
    .X(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W6BEG4 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0534_ (.S0(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit3.Q ),
    .A0(UIO_OUT_TT_PROJECT5),
    .A1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG10 ),
    .A2(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG6 ),
    .A3(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG1 ),
    .S1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit2.Q ),
    .X(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W6BEG5 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0535_ (.S0(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit4.Q ),
    .A0(UIO_OUT_TT_PROJECT6),
    .A1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG5 ),
    .A2(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG9 ),
    .A3(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG2 ),
    .S1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit5.Q ),
    .X(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W6BEG6 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0536_ (.S0(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit6.Q ),
    .A0(UIO_OUT_TT_PROJECT7),
    .A1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG4 ),
    .A2(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG8 ),
    .A3(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG3 ),
    .S1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit7.Q ),
    .X(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W6BEG7 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0537_ (.S0(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit9.Q ),
    .A0(UIO_OUT_TT_PROJECT0),
    .A1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG7 ),
    .A2(_0011_),
    .A3(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG4 ),
    .S1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit8.Q ),
    .X(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W6BEG8 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0538_ (.S0(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit11.Q ),
    .A0(UIO_OUT_TT_PROJECT1),
    .A1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG6 ),
    .A2(_0012_),
    .A3(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG5 ),
    .S1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit10.Q ),
    .X(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W6BEG9 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0539_ (.S0(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit13.Q ),
    .A0(UIO_OUT_TT_PROJECT2),
    .A1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG5 ),
    .A2(_0013_),
    .A3(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG6 ),
    .S1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit12.Q ),
    .X(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W6BEG10 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0540_ (.S0(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit15.Q ),
    .A0(UIO_OUT_TT_PROJECT3),
    .A1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG4 ),
    .A2(_0014_),
    .A3(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG7 ),
    .S1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit14.Q ),
    .X(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W6BEG11 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _0541_ (.Y(_0015_),
    .B(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit2.Q ),
    .A_N(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG12 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _0542_ (.B1(_0015_),
    .VDD(VPWR),
    .Y(_0016_),
    .VSS(VGND),
    .A1(Tile_X0Y0_E6END[8]),
    .A2(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit2.Q ));
 sg13g2_o21ai_1 _0543_ (.B1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit1.Q ),
    .VDD(VPWR),
    .Y(_0017_),
    .VSS(VGND),
    .A1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit0.Q ),
    .A2(_0016_));
 sg13g2_mux2_1 _0544_ (.A0(_0014_),
    .A1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG0 ),
    .S(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit2.Q ),
    .X(_0018_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _0545_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit0.Q ),
    .A2(_0018_),
    .Y(_0019_),
    .B1(_0017_));
 sg13g2_mux4_1 _0546_ (.S0(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit0.Q ),
    .A0(Tile_X0Y0_E1END[0]),
    .A1(Tile_X0Y0_EE4END[0]),
    .A2(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG4 ),
    .A3(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG8 ),
    .S1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit2.Q ),
    .X(_0020_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _0547_ (.A(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit1.Q ),
    .B(_0020_),
    .Y(_0021_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _0548_ (.A(_0019_),
    .B(_0021_),
    .Y(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N4BEG0 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _0549_ (.Y(_0022_),
    .B(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit5.Q ),
    .A_N(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG13 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _0550_ (.B1(_0022_),
    .VDD(VPWR),
    .Y(_0023_),
    .VSS(VGND),
    .A1(Tile_X0Y0_E6END[9]),
    .A2(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit5.Q ));
 sg13g2_o21ai_1 _0551_ (.B1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit4.Q ),
    .VDD(VPWR),
    .Y(_0024_),
    .VSS(VGND),
    .A1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit3.Q ),
    .A2(_0023_));
 sg13g2_mux2_1 _0552_ (.A0(_0013_),
    .A1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG1 ),
    .S(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit5.Q ),
    .X(_0025_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _0553_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit3.Q ),
    .A2(_0025_),
    .Y(_0026_),
    .B1(_0024_));
 sg13g2_mux4_1 _0554_ (.S0(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit3.Q ),
    .A0(Tile_X0Y0_E1END[1]),
    .A1(Tile_X0Y0_EE4END[1]),
    .A2(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG5 ),
    .A3(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG9 ),
    .S1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit5.Q ),
    .X(_0027_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _0555_ (.A(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit4.Q ),
    .B(_0027_),
    .Y(_0028_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _0556_ (.A(_0026_),
    .B(_0028_),
    .Y(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N4BEG1 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _0557_ (.Y(_0029_),
    .B(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit8.Q ),
    .A_N(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG14 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _0558_ (.B1(_0029_),
    .VDD(VPWR),
    .Y(_0030_),
    .VSS(VGND),
    .A1(Tile_X0Y0_E6END[10]),
    .A2(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit8.Q ));
 sg13g2_o21ai_1 _0559_ (.B1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit7.Q ),
    .VDD(VPWR),
    .Y(_0031_),
    .VSS(VGND),
    .A1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit6.Q ),
    .A2(_0030_));
 sg13g2_mux2_1 _0560_ (.A0(_0012_),
    .A1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG2 ),
    .S(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit8.Q ),
    .X(_0032_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _0561_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit6.Q ),
    .A2(_0032_),
    .Y(_0033_),
    .B1(_0031_));
 sg13g2_mux4_1 _0562_ (.S0(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit6.Q ),
    .A0(Tile_X0Y0_E1END[2]),
    .A1(Tile_X0Y0_EE4END[2]),
    .A2(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG6 ),
    .A3(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG10 ),
    .S1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit8.Q ),
    .X(_0034_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _0563_ (.A(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit7.Q ),
    .B(_0034_),
    .Y(_0035_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _0564_ (.A(_0033_),
    .B(_0035_),
    .Y(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N4BEG2 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _0565_ (.Y(_0036_),
    .B(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit11.Q ),
    .A_N(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG15 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _0566_ (.B1(_0036_),
    .VDD(VPWR),
    .Y(_0037_),
    .VSS(VGND),
    .A1(Tile_X0Y0_E6END[11]),
    .A2(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit11.Q ));
 sg13g2_o21ai_1 _0567_ (.B1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit10.Q ),
    .VDD(VPWR),
    .Y(_0038_),
    .VSS(VGND),
    .A1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit9.Q ),
    .A2(_0037_));
 sg13g2_mux2_1 _0568_ (.A0(_0011_),
    .A1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG3 ),
    .S(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit11.Q ),
    .X(_0039_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _0569_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit9.Q ),
    .A2(_0039_),
    .Y(_0040_),
    .B1(_0038_));
 sg13g2_mux4_1 _0570_ (.S0(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit9.Q ),
    .A0(Tile_X0Y0_E1END[3]),
    .A1(Tile_X0Y0_EE4END[3]),
    .A2(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG7 ),
    .A3(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG11 ),
    .S1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit11.Q ),
    .X(_0041_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _0571_ (.A(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit10.Q ),
    .B(_0041_),
    .Y(_0042_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _0572_ (.A(_0040_),
    .B(_0042_),
    .Y(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N4BEG3 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _0573_ (.Y(_0043_),
    .B(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit6.Q ),
    .A_N(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG12 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _0574_ (.B1(_0043_),
    .VDD(VPWR),
    .Y(_0044_),
    .VSS(VGND),
    .A1(Tile_X0Y0_E6END[4]),
    .A2(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit6.Q ));
 sg13g2_o21ai_1 _0575_ (.B1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit5.Q ),
    .VDD(VPWR),
    .Y(_0045_),
    .VSS(VGND),
    .A1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit4.Q ),
    .A2(_0044_));
 sg13g2_inv_1 _0576_ (.VDD(VPWR),
    .Y(_0046_),
    .A(_0045_),
    .VSS(VGND));
 sg13g2_nand2b_1 _0577_ (.Y(_0047_),
    .B(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit6.Q ),
    .A_N(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG4 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _0578_ (.A(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit4.Q ),
    .B(_0047_),
    .X(_0048_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _0579_ (.B1(_0048_),
    .VDD(VPWR),
    .Y(_0049_),
    .VSS(VGND),
    .A1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit6.Q ),
    .A2(_0014_));
 sg13g2_mux4_1 _0580_ (.S0(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit4.Q ),
    .A0(Tile_X0Y0_E1END[0]),
    .A1(Tile_X0Y0_EE4END[12]),
    .A2(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG4 ),
    .A3(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG8 ),
    .S1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit6.Q ),
    .X(_0050_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _0581_ (.A(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit5.Q ),
    .B(_0050_),
    .Y(_0051_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _0582_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0046_),
    .A2(_0049_),
    .Y(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.S4BEG0 ),
    .B1(_0051_));
 sg13g2_nand2b_1 _0583_ (.Y(_0052_),
    .B(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit9.Q ),
    .A_N(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG13 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _0584_ (.B1(_0052_),
    .VDD(VPWR),
    .Y(_0053_),
    .VSS(VGND),
    .A1(Tile_X0Y0_E6END[5]),
    .A2(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit9.Q ));
 sg13g2_o21ai_1 _0585_ (.B1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit8.Q ),
    .VDD(VPWR),
    .Y(_0054_),
    .VSS(VGND),
    .A1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit7.Q ),
    .A2(_0053_));
 sg13g2_inv_1 _0586_ (.VDD(VPWR),
    .Y(_0055_),
    .A(_0054_),
    .VSS(VGND));
 sg13g2_nand2b_1 _0587_ (.Y(_0056_),
    .B(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit9.Q ),
    .A_N(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG5 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _0588_ (.A(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit7.Q ),
    .B(_0056_),
    .X(_0057_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _0589_ (.B1(_0057_),
    .VDD(VPWR),
    .Y(_0058_),
    .VSS(VGND),
    .A1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit9.Q ),
    .A2(_0013_));
 sg13g2_mux4_1 _0590_ (.S0(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit7.Q ),
    .A0(Tile_X0Y0_E1END[1]),
    .A1(Tile_X0Y0_EE4END[13]),
    .A2(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG5 ),
    .A3(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG9 ),
    .S1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit9.Q ),
    .X(_0059_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _0591_ (.A(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit8.Q ),
    .B(_0059_),
    .Y(_0060_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _0592_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0055_),
    .A2(_0058_),
    .Y(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.S4BEG1 ),
    .B1(_0060_));
 sg13g2_nand2b_1 _0593_ (.Y(_0061_),
    .B(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit12.Q ),
    .A_N(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG14 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _0594_ (.B1(_0061_),
    .VDD(VPWR),
    .Y(_0062_),
    .VSS(VGND),
    .A1(Tile_X0Y0_E6END[6]),
    .A2(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit12.Q ));
 sg13g2_o21ai_1 _0595_ (.B1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit11.Q ),
    .VDD(VPWR),
    .Y(_0063_),
    .VSS(VGND),
    .A1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit10.Q ),
    .A2(_0062_));
 sg13g2_inv_1 _0596_ (.VDD(VPWR),
    .Y(_0064_),
    .A(_0063_),
    .VSS(VGND));
 sg13g2_nand2b_1 _0597_ (.Y(_0065_),
    .B(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit12.Q ),
    .A_N(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG6 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _0598_ (.A(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit10.Q ),
    .B(_0065_),
    .X(_0066_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _0599_ (.B1(_0066_),
    .VDD(VPWR),
    .Y(_0067_),
    .VSS(VGND),
    .A1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit12.Q ),
    .A2(_0012_));
 sg13g2_mux4_1 _0600_ (.S0(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit10.Q ),
    .A0(Tile_X0Y0_E1END[2]),
    .A1(Tile_X0Y0_EE4END[14]),
    .A2(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG6 ),
    .A3(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG10 ),
    .S1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit12.Q ),
    .X(_0068_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _0601_ (.A(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit11.Q ),
    .B(_0068_),
    .Y(_0069_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _0602_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0064_),
    .A2(_0067_),
    .Y(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.S4BEG2 ),
    .B1(_0069_));
 sg13g2_nand2b_1 _0603_ (.Y(_0070_),
    .B(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit15.Q ),
    .A_N(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG15 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _0604_ (.B1(_0070_),
    .VDD(VPWR),
    .Y(_0071_),
    .VSS(VGND),
    .A1(Tile_X0Y0_E6END[7]),
    .A2(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit15.Q ));
 sg13g2_o21ai_1 _0605_ (.B1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit14.Q ),
    .VDD(VPWR),
    .Y(_0072_),
    .VSS(VGND),
    .A1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit13.Q ),
    .A2(_0071_));
 sg13g2_inv_1 _0606_ (.VDD(VPWR),
    .Y(_0073_),
    .A(_0072_),
    .VSS(VGND));
 sg13g2_nand2b_1 _0607_ (.Y(_0074_),
    .B(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit15.Q ),
    .A_N(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG7 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _0608_ (.A(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit13.Q ),
    .B(_0074_),
    .X(_0075_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _0609_ (.B1(_0075_),
    .VDD(VPWR),
    .Y(_0076_),
    .VSS(VGND),
    .A1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit15.Q ),
    .A2(_0011_));
 sg13g2_mux4_1 _0610_ (.S0(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit13.Q ),
    .A0(Tile_X0Y0_E1END[3]),
    .A1(Tile_X0Y0_EE4END[15]),
    .A2(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG7 ),
    .A3(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG11 ),
    .S1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit15.Q ),
    .X(_0077_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _0611_ (.A(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit14.Q ),
    .B(_0077_),
    .Y(_0078_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _0612_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0073_),
    .A2(_0076_),
    .Y(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.S4BEG3 ),
    .B1(_0078_));
 sg13g2_mux4_1 _0613_ (.S0(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit0.Q ),
    .A0(Tile_X0Y1_N1END[0]),
    .A1(Tile_X0Y1_N4END[0]),
    .A2(_0007_),
    .A3(Tile_X0Y0_S4END[4]),
    .S1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit1.Q ),
    .X(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.J_NS4_BEG12 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0614_ (.S0(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit2.Q ),
    .A0(Tile_X0Y1_N1END[1]),
    .A1(Tile_X0Y1_N4END[1]),
    .A2(_0311_),
    .A3(Tile_X0Y0_S4END[5]),
    .S1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit3.Q ),
    .X(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.J_NS4_BEG13 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0615_ (.S0(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit4.Q ),
    .A0(Tile_X0Y1_N1END[2]),
    .A1(Tile_X0Y1_N4END[2]),
    .A2(_0318_),
    .A3(Tile_X0Y0_S4END[6]),
    .S1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit5.Q ),
    .X(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.J_NS4_BEG14 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0616_ (.S0(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit6.Q ),
    .A0(Tile_X0Y1_N1END[3]),
    .A1(Tile_X0Y1_N4END[3]),
    .A2(_0325_),
    .A3(Tile_X0Y0_S4END[7]),
    .S1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit7.Q ),
    .X(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.J_NS4_BEG15 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _0617_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0291_),
    .A2(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit16.Q ),
    .Y(_0079_),
    .B1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit18.Q ));
 sg13g2_o21ai_1 _0618_ (.B1(_0079_),
    .VDD(VPWR),
    .Y(_0080_),
    .VSS(VGND),
    .A1(Tile_X0Y0_E6END[0]),
    .A2(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit16.Q ));
 sg13g2_mux4_1 _0619_ (.S0(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit16.Q ),
    .A0(Tile_X0Y0_EE4END[0]),
    .A1(Tile_X0Y0_EE4END[8]),
    .A2(_0014_),
    .A3(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG8 ),
    .S1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit18.Q ),
    .X(_0081_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _0620_ (.A(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit17.Q ),
    .B(_0081_),
    .Y(_0082_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _0621_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit17.Q ),
    .A2(_0080_),
    .Y(UIO_IN_TT_PROJECT0),
    .B1(_0082_));
 sg13g2_a21oi_1 _0622_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0292_),
    .A2(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit19.Q ),
    .Y(_0083_),
    .B1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit21.Q ));
 sg13g2_o21ai_1 _0623_ (.B1(_0083_),
    .VDD(VPWR),
    .Y(_0084_),
    .VSS(VGND),
    .A1(Tile_X0Y0_E6END[1]),
    .A2(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit19.Q ));
 sg13g2_mux4_1 _0624_ (.S0(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit19.Q ),
    .A0(Tile_X0Y0_EE4END[1]),
    .A1(Tile_X0Y0_EE4END[9]),
    .A2(_0013_),
    .A3(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG9 ),
    .S1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit21.Q ),
    .X(_0085_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _0625_ (.A(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit20.Q ),
    .B(_0085_),
    .Y(_0086_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _0626_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit20.Q ),
    .A2(_0084_),
    .Y(UIO_IN_TT_PROJECT1),
    .B1(_0086_));
 sg13g2_a21oi_1 _0627_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0293_),
    .A2(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit22.Q ),
    .Y(_0087_),
    .B1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit24.Q ));
 sg13g2_o21ai_1 _0628_ (.B1(_0087_),
    .VDD(VPWR),
    .Y(_0088_),
    .VSS(VGND),
    .A1(Tile_X0Y0_E6END[2]),
    .A2(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit22.Q ));
 sg13g2_mux4_1 _0629_ (.S0(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit22.Q ),
    .A0(Tile_X0Y0_EE4END[2]),
    .A1(Tile_X0Y0_EE4END[10]),
    .A2(_0012_),
    .A3(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG10 ),
    .S1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit24.Q ),
    .X(_0089_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _0630_ (.A(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit23.Q ),
    .B(_0089_),
    .Y(_0090_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _0631_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit23.Q ),
    .A2(_0088_),
    .Y(UIO_IN_TT_PROJECT2),
    .B1(_0090_));
 sg13g2_a21oi_1 _0632_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0294_),
    .A2(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit25.Q ),
    .Y(_0091_),
    .B1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit27.Q ));
 sg13g2_o21ai_1 _0633_ (.B1(_0091_),
    .VDD(VPWR),
    .Y(_0092_),
    .VSS(VGND),
    .A1(Tile_X0Y0_E6END[3]),
    .A2(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit25.Q ));
 sg13g2_mux4_1 _0634_ (.S0(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit25.Q ),
    .A0(Tile_X0Y0_EE4END[3]),
    .A1(Tile_X0Y0_EE4END[11]),
    .A2(_0011_),
    .A3(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG11 ),
    .S1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit27.Q ),
    .X(_0093_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _0635_ (.A(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit26.Q ),
    .B(_0093_),
    .Y(_0094_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _0636_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit26.Q ),
    .A2(_0092_),
    .Y(UIO_IN_TT_PROJECT3),
    .B1(_0094_));
 sg13g2_nor2b_1 _0637_ (.A(Tile_X0Y0_E6END[4]),
    .B_N(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit28.Q ),
    .Y(_0095_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _0638_ (.B1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit29.Q ),
    .VDD(VPWR),
    .Y(_0096_),
    .VSS(VGND),
    .A1(Tile_X0Y0_EE4END[12]),
    .A2(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit28.Q ));
 sg13g2_mux4_1 _0639_ (.S0(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit28.Q ),
    .A0(Tile_X0Y0_E1END[0]),
    .A1(Tile_X0Y0_EE4END[4]),
    .A2(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG4 ),
    .A3(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG12 ),
    .S1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit30.Q ),
    .X(_0097_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _0640_ (.A(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit29.Q ),
    .B_N(_0097_),
    .Y(_0098_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _0641_ (.A(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit30.Q ),
    .B(_0095_),
    .C(_0096_),
    .Y(_0099_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _0642_ (.VSS(VGND),
    .VDD(VPWR),
    .X(UIO_IN_TT_PROJECT4),
    .B(_0099_),
    .A(_0098_));
 sg13g2_nor2b_1 _0643_ (.A(Tile_X0Y0_E6END[5]),
    .B_N(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit31.Q ),
    .Y(_0100_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _0644_ (.B1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit0.Q ),
    .VDD(VPWR),
    .Y(_0101_),
    .VSS(VGND),
    .A1(Tile_X0Y0_EE4END[13]),
    .A2(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit31.Q ));
 sg13g2_mux4_1 _0645_ (.S0(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit31.Q ),
    .A0(Tile_X0Y0_E1END[1]),
    .A1(Tile_X0Y0_EE4END[5]),
    .A2(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG5 ),
    .A3(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG13 ),
    .S1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit1.Q ),
    .X(_0102_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _0646_ (.A(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit0.Q ),
    .B_N(_0102_),
    .Y(_0103_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _0647_ (.A(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit1.Q ),
    .B(_0100_),
    .C(_0101_),
    .Y(_0104_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _0648_ (.VSS(VGND),
    .VDD(VPWR),
    .X(UIO_IN_TT_PROJECT5),
    .B(_0104_),
    .A(_0103_));
 sg13g2_nor2b_1 _0649_ (.A(Tile_X0Y0_E6END[6]),
    .B_N(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit2.Q ),
    .Y(_0105_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _0650_ (.B1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit3.Q ),
    .VDD(VPWR),
    .Y(_0106_),
    .VSS(VGND),
    .A1(Tile_X0Y0_EE4END[14]),
    .A2(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit2.Q ));
 sg13g2_mux4_1 _0651_ (.S0(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit2.Q ),
    .A0(Tile_X0Y0_E1END[2]),
    .A1(Tile_X0Y0_EE4END[6]),
    .A2(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG6 ),
    .A3(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG14 ),
    .S1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit4.Q ),
    .X(_0107_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _0652_ (.A(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit3.Q ),
    .B_N(_0107_),
    .Y(_0108_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _0653_ (.A(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit4.Q ),
    .B(_0105_),
    .C(_0106_),
    .Y(_0109_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _0654_ (.VSS(VGND),
    .VDD(VPWR),
    .X(UIO_IN_TT_PROJECT6),
    .B(_0109_),
    .A(_0108_));
 sg13g2_nor2b_1 _0655_ (.A(Tile_X0Y0_E6END[7]),
    .B_N(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit5.Q ),
    .Y(_0110_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _0656_ (.B1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit6.Q ),
    .VDD(VPWR),
    .Y(_0111_),
    .VSS(VGND),
    .A1(Tile_X0Y0_EE4END[15]),
    .A2(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit5.Q ));
 sg13g2_mux4_1 _0657_ (.S0(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit5.Q ),
    .A0(Tile_X0Y0_E1END[3]),
    .A1(Tile_X0Y0_EE4END[7]),
    .A2(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG7 ),
    .A3(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG15 ),
    .S1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit7.Q ),
    .X(_0112_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _0658_ (.A(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit6.Q ),
    .B_N(_0112_),
    .Y(_0113_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _0659_ (.A(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit7.Q ),
    .B(_0110_),
    .C(_0111_),
    .Y(_0114_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _0660_ (.VSS(VGND),
    .VDD(VPWR),
    .X(UIO_IN_TT_PROJECT7),
    .B(_0114_),
    .A(_0113_));
 sg13g2_mux4_1 _0661_ (.S0(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit9.Q ),
    .A0(Tile_X0Y0_E1END[0]),
    .A1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG12 ),
    .A2(Tile_X0Y0_E6END[4]),
    .A3(_0006_),
    .S1(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit8.Q ),
    .X(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N1BEG0 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0662_ (.S0(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit4.Q ),
    .A0(Tile_X0Y1_E1END[0]),
    .A1(Tile_X0Y1_E6END[8]),
    .A2(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.J_NS4_BEG12 ),
    .A3(_0010_),
    .S1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit5.Q ),
    .X(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.S1BEG0 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0663_ (.S0(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit6.Q ),
    .A0(Tile_X0Y1_E1END[1]),
    .A1(Tile_X0Y1_E6END[9]),
    .A2(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.J_NS4_BEG13 ),
    .A3(_0314_),
    .S1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit7.Q ),
    .X(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.S1BEG1 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0664_ (.S0(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit8.Q ),
    .A0(Tile_X0Y1_E1END[2]),
    .A1(Tile_X0Y1_E6END[10]),
    .A2(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.J_NS4_BEG14 ),
    .A3(_0321_),
    .S1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit9.Q ),
    .X(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.S1BEG2 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0665_ (.S0(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit10.Q ),
    .A0(Tile_X0Y1_E1END[3]),
    .A1(Tile_X0Y1_E6END[11]),
    .A2(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.J_NS4_BEG15 ),
    .A3(_0328_),
    .S1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit11.Q ),
    .X(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.S1BEG3 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0666_ (.S0(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit12.Q ),
    .A0(Tile_X0Y1_E2MID[7]),
    .A1(Tile_X0Y1_E2END[7]),
    .A2(Tile_X0Y1_E6END[8]),
    .A3(_0335_),
    .S1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit13.Q ),
    .X(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.S2BEG0 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0667_ (.S0(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit14.Q ),
    .A0(Tile_X0Y1_E2MID[6]),
    .A1(Tile_X0Y1_E2END[6]),
    .A2(Tile_X0Y1_E6END[9]),
    .A3(_0342_),
    .S1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit15.Q ),
    .X(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.S2BEG1 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0668_ (.S0(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit16.Q ),
    .A0(Tile_X0Y1_E2MID[5]),
    .A1(Tile_X0Y1_E2END[5]),
    .A2(Tile_X0Y1_E6END[10]),
    .A3(_0349_),
    .S1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit17.Q ),
    .X(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.S2BEG2 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0669_ (.S0(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit18.Q ),
    .A0(Tile_X0Y1_E2MID[4]),
    .A1(Tile_X0Y1_E2END[4]),
    .A2(Tile_X0Y1_E6END[11]),
    .A3(_0356_),
    .S1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit19.Q ),
    .X(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.S2BEG3 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0670_ (.S0(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit21.Q ),
    .A0(Tile_X0Y1_E1END[0]),
    .A1(Tile_X0Y1_E2END[3]),
    .A2(Tile_X0Y1_E2MID[3]),
    .A3(_0000_),
    .S1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit20.Q ),
    .X(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.S2BEG4 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0671_ (.S0(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit23.Q ),
    .A0(Tile_X0Y1_E1END[1]),
    .A1(Tile_X0Y1_E2END[2]),
    .A2(Tile_X0Y1_E2MID[2]),
    .A3(_0001_),
    .S1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit22.Q ),
    .X(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.S2BEG5 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0672_ (.S0(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit25.Q ),
    .A0(Tile_X0Y1_E1END[2]),
    .A1(Tile_X0Y1_E2END[1]),
    .A2(Tile_X0Y1_E2MID[1]),
    .A3(_0002_),
    .S1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit24.Q ),
    .X(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.S2BEG6 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0673_ (.S0(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit27.Q ),
    .A0(Tile_X0Y1_E1END[3]),
    .A1(Tile_X0Y1_E2END[0]),
    .A2(Tile_X0Y1_E2MID[0]),
    .A3(_0003_),
    .S1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit26.Q ),
    .X(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.S2BEG7 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0674_ (.S0(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit9.Q ),
    .A0(Tile_X0Y1_N1END[0]),
    .A1(UO_OUT_TT_PROJECT2),
    .A2(_0007_),
    .A3(UO_OUT_TT_PROJECT7),
    .S1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit8.Q ),
    .X(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W1BEG0 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0675_ (.S0(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit11.Q ),
    .A0(Tile_X0Y1_N1END[1]),
    .A1(UO_OUT_TT_PROJECT3),
    .A2(_0311_),
    .A3(UO_OUT_TT_PROJECT6),
    .S1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit10.Q ),
    .X(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W1BEG1 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0676_ (.S0(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit13.Q ),
    .A0(Tile_X0Y1_N1END[2]),
    .A1(UO_OUT_TT_PROJECT0),
    .A2(_0318_),
    .A3(UO_OUT_TT_PROJECT5),
    .S1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit12.Q ),
    .X(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W1BEG2 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0677_ (.S0(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit15.Q ),
    .A0(Tile_X0Y1_N1END[3]),
    .A1(UO_OUT_TT_PROJECT1),
    .A2(_0325_),
    .A3(UO_OUT_TT_PROJECT4),
    .S1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit14.Q ),
    .X(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W1BEG3 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _0678_ (.Y(_0115_),
    .B(_0003_),
    .A_N(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit16.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _0679_ (.A(UO_OUT_TT_PROJECT0),
    .B(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit16.Q ),
    .C(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit17.Q ),
    .Y(_0116_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _0680_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit17.Q ),
    .C1(_0116_),
    .B1(_0115_),
    .A1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit16.Q ),
    .Y(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W2BEG0 ),
    .A2(_0334_));
 sg13g2_nand2b_1 _0681_ (.Y(_0117_),
    .B(_0002_),
    .A_N(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit18.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _0682_ (.A(UO_OUT_TT_PROJECT1),
    .B(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit18.Q ),
    .C(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit19.Q ),
    .Y(_0118_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _0683_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit19.Q ),
    .C1(_0118_),
    .B1(_0117_),
    .A1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit18.Q ),
    .Y(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W2BEG1 ),
    .A2(_0341_));
 sg13g2_nand2b_1 _0684_ (.Y(_0119_),
    .B(_0001_),
    .A_N(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit20.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _0685_ (.A(UO_OUT_TT_PROJECT2),
    .B(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit20.Q ),
    .C(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit21.Q ),
    .Y(_0120_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _0686_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit21.Q ),
    .C1(_0120_),
    .B1(_0119_),
    .A1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit20.Q ),
    .Y(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W2BEG2 ),
    .A2(_0348_));
 sg13g2_nand2b_1 _0687_ (.Y(_0121_),
    .B(_0000_),
    .A_N(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit22.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _0688_ (.A(UO_OUT_TT_PROJECT3),
    .B(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit22.Q ),
    .C(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit23.Q ),
    .Y(_0122_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _0689_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit23.Q ),
    .C1(_0122_),
    .B1(_0121_),
    .A1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit22.Q ),
    .Y(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W2BEG3 ),
    .A2(_0355_));
 sg13g2_nand2b_1 _0690_ (.Y(_0123_),
    .B(_0000_),
    .A_N(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit24.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _0691_ (.A(UO_OUT_TT_PROJECT4),
    .B(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit24.Q ),
    .C(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit25.Q ),
    .Y(_0124_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _0692_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit25.Q ),
    .C1(_0124_),
    .B1(_0123_),
    .A1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit24.Q ),
    .Y(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W2BEG4 ),
    .A2(_0355_));
 sg13g2_nand2b_1 _0693_ (.Y(_0125_),
    .B(_0001_),
    .A_N(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit26.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _0694_ (.A(UO_OUT_TT_PROJECT5),
    .B(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit26.Q ),
    .C(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit27.Q ),
    .Y(_0126_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _0695_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit27.Q ),
    .C1(_0126_),
    .B1(_0125_),
    .A1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit26.Q ),
    .Y(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W2BEG5 ),
    .A2(_0348_));
 sg13g2_nand2b_1 _0696_ (.Y(_0127_),
    .B(_0002_),
    .A_N(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit28.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _0697_ (.A(UO_OUT_TT_PROJECT6),
    .B(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit28.Q ),
    .C(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit29.Q ),
    .Y(_0128_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _0698_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit29.Q ),
    .C1(_0128_),
    .B1(_0127_),
    .A1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit28.Q ),
    .Y(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W2BEG6 ),
    .A2(_0341_));
 sg13g2_nand2b_1 _0699_ (.Y(_0129_),
    .B(_0003_),
    .A_N(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit30.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _0700_ (.A(UO_OUT_TT_PROJECT7),
    .B(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit30.Q ),
    .C(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit31.Q ),
    .Y(_0130_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _0701_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit31.Q ),
    .C1(_0130_),
    .B1(_0129_),
    .A1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit30.Q ),
    .Y(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W2BEG7 ),
    .A2(_0334_));
 sg13g2_nand2b_1 _0702_ (.Y(_0131_),
    .B(_0003_),
    .A_N(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit0.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _0703_ (.A(UO_OUT_TT_PROJECT0),
    .B(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit0.Q ),
    .C(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit1.Q ),
    .Y(_0132_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _0704_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit1.Q ),
    .C1(_0132_),
    .B1(_0131_),
    .A1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit0.Q ),
    .Y(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W2BEGb0 ),
    .A2(_0334_));
 sg13g2_nand2b_1 _0705_ (.Y(_0133_),
    .B(_0002_),
    .A_N(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit2.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _0706_ (.A(UO_OUT_TT_PROJECT1),
    .B(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit2.Q ),
    .C(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit3.Q ),
    .Y(_0134_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _0707_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit3.Q ),
    .C1(_0134_),
    .B1(_0133_),
    .A1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit2.Q ),
    .Y(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W2BEGb1 ),
    .A2(_0341_));
 sg13g2_nand2b_1 _0708_ (.Y(_0135_),
    .B(_0001_),
    .A_N(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit4.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _0709_ (.A(UO_OUT_TT_PROJECT2),
    .B(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit4.Q ),
    .C(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit5.Q ),
    .Y(_0136_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _0710_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit5.Q ),
    .C1(_0136_),
    .B1(_0135_),
    .A1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit4.Q ),
    .Y(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W2BEGb2 ),
    .A2(_0348_));
 sg13g2_nand2b_1 _0711_ (.Y(_0137_),
    .B(_0000_),
    .A_N(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit6.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _0712_ (.A(UO_OUT_TT_PROJECT3),
    .B(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit6.Q ),
    .C(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit7.Q ),
    .Y(_0138_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _0713_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit7.Q ),
    .C1(_0138_),
    .B1(_0137_),
    .A1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit6.Q ),
    .Y(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W2BEGb3 ),
    .A2(_0355_));
 sg13g2_nand2b_1 _0714_ (.Y(_0139_),
    .B(_0000_),
    .A_N(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit8.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _0715_ (.A(UO_OUT_TT_PROJECT4),
    .B(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit8.Q ),
    .C(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit9.Q ),
    .Y(_0140_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _0716_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit9.Q ),
    .C1(_0140_),
    .B1(_0139_),
    .A1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit8.Q ),
    .Y(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W2BEGb4 ),
    .A2(_0355_));
 sg13g2_nand2b_1 _0717_ (.Y(_0141_),
    .B(_0001_),
    .A_N(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit10.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _0718_ (.A(UO_OUT_TT_PROJECT5),
    .B(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit10.Q ),
    .C(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit11.Q ),
    .Y(_0142_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _0719_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit11.Q ),
    .C1(_0142_),
    .B1(_0141_),
    .A1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit10.Q ),
    .Y(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W2BEGb5 ),
    .A2(_0348_));
 sg13g2_nand2b_1 _0720_ (.Y(_0143_),
    .B(_0002_),
    .A_N(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit12.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _0721_ (.A(UO_OUT_TT_PROJECT6),
    .B(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit12.Q ),
    .C(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit13.Q ),
    .Y(_0144_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _0722_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit13.Q ),
    .C1(_0144_),
    .B1(_0143_),
    .A1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit12.Q ),
    .Y(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W2BEGb6 ),
    .A2(_0341_));
 sg13g2_nand2b_1 _0723_ (.Y(_0145_),
    .B(_0003_),
    .A_N(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit14.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _0724_ (.A(UO_OUT_TT_PROJECT7),
    .B(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit14.Q ),
    .C(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit15.Q ),
    .Y(_0146_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _0725_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit15.Q ),
    .C1(_0146_),
    .B1(_0145_),
    .A1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit14.Q ),
    .Y(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W2BEGb7 ),
    .A2(_0334_));
 sg13g2_mux4_1 _0726_ (.S0(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit16.Q ),
    .A0(UO_OUT_TT_PROJECT0),
    .A1(UO_OUT_TT_PROJECT4),
    .A2(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.J_NS4_BEG15 ),
    .A3(_0003_),
    .S1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit17.Q ),
    .X(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.WW4BEG0 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0727_ (.S0(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit19.Q ),
    .A0(UO_OUT_TT_PROJECT1),
    .A1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.J_NS4_BEG14 ),
    .A2(UO_OUT_TT_PROJECT5),
    .A3(_0002_),
    .S1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit18.Q ),
    .X(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.WW4BEG1 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0728_ (.S0(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit20.Q ),
    .A0(UO_OUT_TT_PROJECT2),
    .A1(UO_OUT_TT_PROJECT6),
    .A2(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.J_NS4_BEG13 ),
    .A3(_0001_),
    .S1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit21.Q ),
    .X(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.WW4BEG2 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0729_ (.S0(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit23.Q ),
    .A0(UO_OUT_TT_PROJECT3),
    .A1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.J_NS4_BEG12 ),
    .A2(UO_OUT_TT_PROJECT7),
    .A3(_0000_),
    .S1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit22.Q ),
    .X(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.WW4BEG3 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0730_ (.S0(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit30.Q ),
    .A0(Tile_X0Y1_N1END[3]),
    .A1(Tile_X0Y1_N4END[3]),
    .A2(_0325_),
    .A3(Tile_X0Y0_S4END[7]),
    .S1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit31.Q ),
    .X(_0147_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0731_ (.S0(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit24.Q ),
    .A0(UO_OUT_TT_PROJECT0),
    .A1(UO_OUT_TT_PROJECT4),
    .A2(_0147_),
    .A3(_0356_),
    .S1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit25.Q ),
    .X(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.WW4BEG4 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0732_ (.S0(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit28.Q ),
    .A0(Tile_X0Y1_N1END[2]),
    .A1(Tile_X0Y1_N4END[2]),
    .A2(_0318_),
    .A3(Tile_X0Y0_S4END[6]),
    .S1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit29.Q ),
    .X(_0148_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0733_ (.S0(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit27.Q ),
    .A0(UO_OUT_TT_PROJECT1),
    .A1(_0148_),
    .A2(UO_OUT_TT_PROJECT5),
    .A3(_0349_),
    .S1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit26.Q ),
    .X(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.WW4BEG5 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0734_ (.S0(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit26.Q ),
    .A0(Tile_X0Y1_N1END[1]),
    .A1(Tile_X0Y1_N4END[1]),
    .A2(_0311_),
    .A3(Tile_X0Y0_S4END[5]),
    .S1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit27.Q ),
    .X(_0149_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0735_ (.S0(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit28.Q ),
    .A0(UO_OUT_TT_PROJECT2),
    .A1(UO_OUT_TT_PROJECT6),
    .A2(_0149_),
    .A3(_0342_),
    .S1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit29.Q ),
    .X(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.WW4BEG6 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0736_ (.S0(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit24.Q ),
    .A0(Tile_X0Y1_N1END[0]),
    .A1(Tile_X0Y1_N4END[0]),
    .A2(_0007_),
    .A3(Tile_X0Y0_S4END[4]),
    .S1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit25.Q ),
    .X(_0150_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0737_ (.S0(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit31.Q ),
    .A0(UO_OUT_TT_PROJECT3),
    .A1(_0150_),
    .A2(UO_OUT_TT_PROJECT7),
    .A3(_0335_),
    .S1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit30.Q ),
    .X(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.WW4BEG7 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0738_ (.S0(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit22.Q ),
    .A0(Tile_X0Y1_N1END[3]),
    .A1(Tile_X0Y1_N4END[3]),
    .A2(_0325_),
    .A3(Tile_X0Y0_S4END[7]),
    .S1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit23.Q ),
    .X(_0151_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0739_ (.S0(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit0.Q ),
    .A0(UO_OUT_TT_PROJECT0),
    .A1(UO_OUT_TT_PROJECT4),
    .A2(_0151_),
    .A3(_0003_),
    .S1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit1.Q ),
    .X(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.WW4BEG8 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0740_ (.S0(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit20.Q ),
    .A0(Tile_X0Y1_N1END[2]),
    .A1(Tile_X0Y1_N4END[2]),
    .A2(_0318_),
    .A3(Tile_X0Y0_S4END[6]),
    .S1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit21.Q ),
    .X(_0152_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0741_ (.S0(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit3.Q ),
    .A0(UO_OUT_TT_PROJECT1),
    .A1(_0152_),
    .A2(UO_OUT_TT_PROJECT5),
    .A3(_0002_),
    .S1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit2.Q ),
    .X(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.WW4BEG9 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0742_ (.S0(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit18.Q ),
    .A0(Tile_X0Y1_N1END[1]),
    .A1(Tile_X0Y1_N4END[1]),
    .A2(_0311_),
    .A3(Tile_X0Y0_S4END[5]),
    .S1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit19.Q ),
    .X(_0153_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0743_ (.S0(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit4.Q ),
    .A0(UO_OUT_TT_PROJECT2),
    .A1(UO_OUT_TT_PROJECT6),
    .A2(_0153_),
    .A3(_0001_),
    .S1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit5.Q ),
    .X(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.WW4BEG10 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0744_ (.S0(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit16.Q ),
    .A0(Tile_X0Y1_N1END[0]),
    .A1(Tile_X0Y1_N4END[0]),
    .A2(_0007_),
    .A3(Tile_X0Y0_S4END[4]),
    .S1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit17.Q ),
    .X(_0154_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0745_ (.S0(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit7.Q ),
    .A0(UO_OUT_TT_PROJECT3),
    .A1(_0154_),
    .A2(UO_OUT_TT_PROJECT7),
    .A3(_0000_),
    .S1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit6.Q ),
    .X(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.WW4BEG11 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0746_ (.S0(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit14.Q ),
    .A0(Tile_X0Y1_N1END[3]),
    .A1(Tile_X0Y1_N4END[3]),
    .A2(_0325_),
    .A3(Tile_X0Y0_S4END[7]),
    .S1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit15.Q ),
    .X(_0155_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0747_ (.S0(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit8.Q ),
    .A0(UO_OUT_TT_PROJECT0),
    .A1(UO_OUT_TT_PROJECT4),
    .A2(_0155_),
    .A3(_0356_),
    .S1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit9.Q ),
    .X(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.WW4BEG12 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0748_ (.S0(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit12.Q ),
    .A0(Tile_X0Y1_N1END[2]),
    .A1(Tile_X0Y1_N4END[2]),
    .A2(_0318_),
    .A3(Tile_X0Y0_S4END[6]),
    .S1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit13.Q ),
    .X(_0156_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0749_ (.S0(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit11.Q ),
    .A0(UO_OUT_TT_PROJECT1),
    .A1(_0156_),
    .A2(UO_OUT_TT_PROJECT5),
    .A3(_0349_),
    .S1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit10.Q ),
    .X(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.WW4BEG13 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0750_ (.S0(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit10.Q ),
    .A0(Tile_X0Y1_N1END[1]),
    .A1(Tile_X0Y1_N4END[1]),
    .A2(_0311_),
    .A3(Tile_X0Y0_S4END[5]),
    .S1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit11.Q ),
    .X(_0157_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0751_ (.S0(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit12.Q ),
    .A0(UO_OUT_TT_PROJECT2),
    .A1(UO_OUT_TT_PROJECT6),
    .A2(_0157_),
    .A3(_0342_),
    .S1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit13.Q ),
    .X(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.WW4BEG14 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0752_ (.S0(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit8.Q ),
    .A0(Tile_X0Y1_N1END[0]),
    .A1(Tile_X0Y1_N4END[0]),
    .A2(_0007_),
    .A3(Tile_X0Y0_S4END[4]),
    .S1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit9.Q ),
    .X(_0158_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0753_ (.S0(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit15.Q ),
    .A0(UO_OUT_TT_PROJECT3),
    .A1(_0158_),
    .A2(UO_OUT_TT_PROJECT7),
    .A3(_0335_),
    .S1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit14.Q ),
    .X(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.WW4BEG15 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0754_ (.S0(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit16.Q ),
    .A0(Tile_X0Y1_N4END[0]),
    .A1(Tile_X0Y0_S4END[4]),
    .A2(_0147_),
    .A3(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.J_NS4_BEG15 ),
    .S1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit17.Q ),
    .X(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W6BEG0 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0755_ (.S0(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit18.Q ),
    .A0(Tile_X0Y1_N4END[1]),
    .A1(Tile_X0Y0_S4END[5]),
    .A2(_0148_),
    .A3(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.J_NS4_BEG14 ),
    .S1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit19.Q ),
    .X(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W6BEG1 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0756_ (.S0(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit20.Q ),
    .A0(Tile_X0Y1_N4END[2]),
    .A1(Tile_X0Y0_S4END[6]),
    .A2(_0149_),
    .A3(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.J_NS4_BEG13 ),
    .S1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit21.Q ),
    .X(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W6BEG2 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0757_ (.S0(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit22.Q ),
    .A0(Tile_X0Y1_N4END[3]),
    .A1(Tile_X0Y0_S4END[7]),
    .A2(_0150_),
    .A3(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.J_NS4_BEG12 ),
    .S1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit23.Q ),
    .X(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W6BEG3 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0758_ (.S0(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit25.Q ),
    .A0(UO_OUT_TT_PROJECT4),
    .A1(_0147_),
    .A2(_0151_),
    .A3(_0335_),
    .S1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit24.Q ),
    .X(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W6BEG4 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0759_ (.S0(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit27.Q ),
    .A0(UO_OUT_TT_PROJECT5),
    .A1(_0148_),
    .A2(_0152_),
    .A3(_0342_),
    .S1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit26.Q ),
    .X(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W6BEG5 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0760_ (.S0(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit29.Q ),
    .A0(UO_OUT_TT_PROJECT6),
    .A1(_0149_),
    .A2(_0153_),
    .A3(_0349_),
    .S1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit28.Q ),
    .X(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W6BEG6 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0761_ (.S0(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit31.Q ),
    .A0(UO_OUT_TT_PROJECT7),
    .A1(_0150_),
    .A2(_0154_),
    .A3(_0356_),
    .S1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit30.Q ),
    .X(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W6BEG7 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0762_ (.S0(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit1.Q ),
    .A0(UO_OUT_TT_PROJECT0),
    .A1(_0151_),
    .A2(_0155_),
    .A3(_0000_),
    .S1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit0.Q ),
    .X(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W6BEG8 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0763_ (.S0(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit3.Q ),
    .A0(UO_OUT_TT_PROJECT1),
    .A1(_0152_),
    .A2(_0156_),
    .A3(_0001_),
    .S1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit2.Q ),
    .X(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W6BEG9 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0764_ (.S0(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit5.Q ),
    .A0(UO_OUT_TT_PROJECT2),
    .A1(_0153_),
    .A2(_0157_),
    .A3(_0002_),
    .S1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit4.Q ),
    .X(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W6BEG10 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0765_ (.S0(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit7.Q ),
    .A0(UO_OUT_TT_PROJECT3),
    .A1(_0154_),
    .A2(_0158_),
    .A3(_0003_),
    .S1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit6.Q ),
    .X(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W6BEG11 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _0766_ (.A0(_0154_),
    .A1(_0150_),
    .S(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit24.Q ),
    .X(_0159_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _0767_ (.Y(_0160_),
    .B(_0159_),
    .A_N(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit25.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _0768_ (.B1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit25.Q ),
    .VDD(VPWR),
    .Y(_0161_),
    .VSS(VGND),
    .A1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit24.Q ),
    .A2(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.J_NS4_BEG12 ));
 sg13g2_a21oi_1 _0769_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit24.Q ),
    .A2(_0334_),
    .Y(_0162_),
    .B1(_0161_));
 sg13g2_nor2b_1 _0770_ (.A(_0162_),
    .B_N(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit26.Q ),
    .Y(_0163_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0771_ (.S0(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit25.Q ),
    .A0(Tile_X0Y1_E1END[0]),
    .A1(Tile_X0Y1_E6END[8]),
    .A2(Tile_X0Y1_EE4END[0]),
    .A3(_0158_),
    .S1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit24.Q ),
    .X(_0164_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _0772_ (.A(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit26.Q ),
    .B(_0164_),
    .Y(_0165_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _0773_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0160_),
    .A2(_0163_),
    .Y(\Tile_X0Y0_E_TT_IF2_top.N4BEG_outbuf_8.A ),
    .B1(_0165_));
 sg13g2_mux2_1 _0774_ (.A0(_0153_),
    .A1(_0149_),
    .S(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit27.Q ),
    .X(_0166_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _0775_ (.Y(_0167_),
    .B(_0166_),
    .A_N(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit28.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _0776_ (.B1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit28.Q ),
    .VDD(VPWR),
    .Y(_0168_),
    .VSS(VGND),
    .A1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit27.Q ),
    .A2(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.J_NS4_BEG13 ));
 sg13g2_a21oi_1 _0777_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit27.Q ),
    .A2(_0341_),
    .Y(_0169_),
    .B1(_0168_));
 sg13g2_nor2b_1 _0778_ (.A(_0169_),
    .B_N(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit29.Q ),
    .Y(_0170_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0779_ (.S0(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit28.Q ),
    .A0(Tile_X0Y1_E1END[1]),
    .A1(Tile_X0Y1_E6END[9]),
    .A2(Tile_X0Y1_EE4END[1]),
    .A3(_0157_),
    .S1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit27.Q ),
    .X(_0171_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _0780_ (.A(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit29.Q ),
    .B(_0171_),
    .Y(_0172_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _0781_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0167_),
    .A2(_0170_),
    .Y(\Tile_X0Y0_E_TT_IF2_top.N4BEG_outbuf_9.A ),
    .B1(_0172_));
 sg13g2_mux2_1 _0782_ (.A0(_0152_),
    .A1(_0148_),
    .S(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit30.Q ),
    .X(_0173_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _0783_ (.Y(_0174_),
    .B(_0173_),
    .A_N(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit31.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _0784_ (.B1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit31.Q ),
    .VDD(VPWR),
    .Y(_0175_),
    .VSS(VGND),
    .A1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit30.Q ),
    .A2(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.J_NS4_BEG14 ));
 sg13g2_a21oi_1 _0785_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit30.Q ),
    .A2(_0348_),
    .Y(_0176_),
    .B1(_0175_));
 sg13g2_nor2b_1 _0786_ (.A(_0176_),
    .B_N(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit0.Q ),
    .Y(_0177_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0787_ (.S0(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit31.Q ),
    .A0(Tile_X0Y1_E1END[2]),
    .A1(Tile_X0Y1_E6END[10]),
    .A2(Tile_X0Y1_EE4END[2]),
    .A3(_0156_),
    .S1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit30.Q ),
    .X(_0178_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _0788_ (.A(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit0.Q ),
    .B(_0178_),
    .Y(_0179_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _0789_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0174_),
    .A2(_0177_),
    .Y(\Tile_X0Y0_E_TT_IF2_top.N4BEG_outbuf_10.A ),
    .B1(_0179_));
 sg13g2_mux2_1 _0790_ (.A0(_0151_),
    .A1(_0147_),
    .S(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit1.Q ),
    .X(_0180_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _0791_ (.Y(_0181_),
    .B(_0180_),
    .A_N(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit2.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _0792_ (.B1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit2.Q ),
    .VDD(VPWR),
    .Y(_0182_),
    .VSS(VGND),
    .A1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit1.Q ),
    .A2(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.J_NS4_BEG15 ));
 sg13g2_a21oi_1 _0793_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit1.Q ),
    .A2(_0355_),
    .Y(_0183_),
    .B1(_0182_));
 sg13g2_nor2b_1 _0794_ (.A(_0183_),
    .B_N(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit3.Q ),
    .Y(_0184_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0795_ (.S0(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit2.Q ),
    .A0(Tile_X0Y1_E1END[3]),
    .A1(Tile_X0Y1_E6END[11]),
    .A2(Tile_X0Y1_EE4END[3]),
    .A3(_0155_),
    .S1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit1.Q ),
    .X(_0185_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _0796_ (.A(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit3.Q ),
    .B(_0185_),
    .Y(_0186_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _0797_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0181_),
    .A2(_0184_),
    .Y(\Tile_X0Y0_E_TT_IF2_top.N4BEG_outbuf_11.A ),
    .B1(_0186_));
 sg13g2_mux2_1 _0798_ (.A0(_0154_),
    .A1(_0150_),
    .S(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit28.Q ),
    .X(_0187_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _0799_ (.Y(_0188_),
    .B(_0187_),
    .A_N(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit29.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _0800_ (.A0(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.J_NS4_BEG12 ),
    .A1(_0000_),
    .S(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit28.Q ),
    .X(_0189_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _0801_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit29.Q ),
    .A2(_0189_),
    .Y(_0190_),
    .B1(_0301_));
 sg13g2_mux4_1 _0802_ (.S0(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit28.Q ),
    .A0(Tile_X0Y1_E1END[0]),
    .A1(Tile_X0Y1_EE4END[12]),
    .A2(Tile_X0Y1_E6END[4]),
    .A3(_0158_),
    .S1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit29.Q ),
    .X(_0191_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _0803_ (.A(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit30.Q ),
    .B(_0191_),
    .Y(_0192_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _0804_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0188_),
    .A2(_0190_),
    .Y(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.S4BEG0 ),
    .B1(_0192_));
 sg13g2_mux2_1 _0805_ (.A0(_0153_),
    .A1(_0149_),
    .S(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit31.Q ),
    .X(_0193_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _0806_ (.Y(_0194_),
    .B(_0193_),
    .A_N(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit0.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _0807_ (.A0(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.J_NS4_BEG13 ),
    .A1(_0001_),
    .S(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit31.Q ),
    .X(_0195_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _0808_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit0.Q ),
    .A2(_0195_),
    .Y(_0196_),
    .B1(_0302_));
 sg13g2_mux4_1 _0809_ (.S0(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit31.Q ),
    .A0(Tile_X0Y1_E1END[1]),
    .A1(Tile_X0Y1_EE4END[13]),
    .A2(Tile_X0Y1_E6END[5]),
    .A3(_0157_),
    .S1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit0.Q ),
    .X(_0197_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _0810_ (.A(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit1.Q ),
    .B(_0197_),
    .Y(_0198_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _0811_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0194_),
    .A2(_0196_),
    .Y(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.S4BEG1 ),
    .B1(_0198_));
 sg13g2_mux2_1 _0812_ (.A0(_0152_),
    .A1(_0148_),
    .S(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit2.Q ),
    .X(_0199_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _0813_ (.Y(_0200_),
    .B(_0199_),
    .A_N(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit3.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _0814_ (.A0(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.J_NS4_BEG14 ),
    .A1(_0002_),
    .S(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit2.Q ),
    .X(_0201_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _0815_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit3.Q ),
    .A2(_0201_),
    .Y(_0202_),
    .B1(_0303_));
 sg13g2_mux4_1 _0816_ (.S0(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit2.Q ),
    .A0(Tile_X0Y1_E1END[2]),
    .A1(Tile_X0Y1_EE4END[14]),
    .A2(Tile_X0Y1_E6END[6]),
    .A3(_0156_),
    .S1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit3.Q ),
    .X(_0203_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _0817_ (.A(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit4.Q ),
    .B(_0203_),
    .Y(_0204_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _0818_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0200_),
    .A2(_0202_),
    .Y(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.S4BEG2 ),
    .B1(_0204_));
 sg13g2_mux2_1 _0819_ (.A0(_0151_),
    .A1(_0147_),
    .S(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit5.Q ),
    .X(_0205_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _0820_ (.Y(_0206_),
    .B(_0205_),
    .A_N(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit6.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _0821_ (.A0(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.J_NS4_BEG15 ),
    .A1(_0003_),
    .S(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit5.Q ),
    .X(_0207_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _0822_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit6.Q ),
    .A2(_0207_),
    .Y(_0208_),
    .B1(_0304_));
 sg13g2_mux4_1 _0823_ (.S0(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit5.Q ),
    .A0(Tile_X0Y1_E1END[3]),
    .A1(Tile_X0Y1_EE4END[15]),
    .A2(Tile_X0Y1_E6END[7]),
    .A3(_0155_),
    .S1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit6.Q ),
    .X(_0209_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _0824_ (.A(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit7.Q ),
    .B(_0209_),
    .Y(_0210_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _0825_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0206_),
    .A2(_0208_),
    .Y(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.S4BEG3 ),
    .B1(_0210_));
 sg13g2_nor2_1 _0826_ (.A(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit8.Q ),
    .B(_0158_),
    .Y(_0211_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _0827_ (.A(_0150_),
    .B_N(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit8.Q ),
    .Y(_0212_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0828_ (.S0(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit8.Q ),
    .A0(Tile_X0Y1_EE4END[0]),
    .A1(Tile_X0Y1_EE4END[8]),
    .A2(Tile_X0Y1_E6END[0]),
    .A3(Tile_X0Y1_E6END[8]),
    .S1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit9.Q ),
    .X(_0213_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _0829_ (.A(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit9.Q ),
    .B(_0211_),
    .C(_0212_),
    .Y(_0214_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _0830_ (.A0(_0213_),
    .A1(_0214_),
    .S(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit10.Q ),
    .X(UI_IN_TT_PROJECT0),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _0831_ (.A0(_0157_),
    .A1(_0149_),
    .S(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit11.Q ),
    .X(_0215_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3b_1 _0832_ (.B(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit13.Q ),
    .C(_0215_),
    .Y(_0216_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit12.Q ));
 sg13g2_mux4_1 _0833_ (.S0(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit11.Q ),
    .A0(Tile_X0Y1_EE4END[1]),
    .A1(Tile_X0Y1_EE4END[9]),
    .A2(Tile_X0Y1_E6END[1]),
    .A3(Tile_X0Y1_E6END[9]),
    .S1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit12.Q ),
    .X(_0217_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _0834_ (.VDD(VPWR),
    .Y(_0218_),
    .A(_0217_),
    .VSS(VGND));
 sg13g2_o21ai_1 _0835_ (.B1(_0216_),
    .VDD(VPWR),
    .Y(UI_IN_TT_PROJECT1),
    .VSS(VGND),
    .A1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit13.Q ),
    .A2(_0218_));
 sg13g2_nor2b_1 _0836_ (.A(_0148_),
    .B_N(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit14.Q ),
    .Y(_0219_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _0837_ (.A(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit14.Q ),
    .B(_0156_),
    .Y(_0220_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0838_ (.S0(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit14.Q ),
    .A0(Tile_X0Y1_EE4END[2]),
    .A1(Tile_X0Y1_EE4END[10]),
    .A2(Tile_X0Y1_E6END[2]),
    .A3(Tile_X0Y1_E6END[10]),
    .S1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit15.Q ),
    .X(_0221_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _0839_ (.A(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit15.Q ),
    .B(_0219_),
    .C(_0220_),
    .Y(_0222_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _0840_ (.A0(_0221_),
    .A1(_0222_),
    .S(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit16.Q ),
    .X(UI_IN_TT_PROJECT2),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _0841_ (.A(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit17.Q ),
    .B(_0155_),
    .Y(_0223_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _0842_ (.A(_0147_),
    .B_N(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit17.Q ),
    .Y(_0224_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0843_ (.S0(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit17.Q ),
    .A0(Tile_X0Y1_EE4END[3]),
    .A1(Tile_X0Y1_EE4END[11]),
    .A2(Tile_X0Y1_E6END[3]),
    .A3(Tile_X0Y1_E6END[11]),
    .S1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit18.Q ),
    .X(_0225_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _0844_ (.A(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit18.Q ),
    .B(_0223_),
    .C(_0224_),
    .Y(_0226_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _0845_ (.A0(_0225_),
    .A1(_0226_),
    .S(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit19.Q ),
    .X(UI_IN_TT_PROJECT3),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0846_ (.S0(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit21.Q ),
    .A0(Tile_X0Y1_E1END[0]),
    .A1(Tile_X0Y1_EE4END[12]),
    .A2(Tile_X0Y1_EE4END[4]),
    .A3(Tile_X0Y1_E6END[4]),
    .S1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit20.Q ),
    .X(_0227_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _0847_ (.Y(_0228_),
    .B(_0227_),
    .A_N(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit22.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _0848_ (.Y(_0229_),
    .B(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit22.Q ),
    .A_N(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit21.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _0849_ (.Y(_0230_),
    .B(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit20.Q ),
    .A_N(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.J_NS4_BEG12 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _0850_ (.B1(_0230_),
    .VDD(VPWR),
    .Y(_0231_),
    .VSS(VGND),
    .A1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit20.Q ),
    .A2(_0154_));
 sg13g2_o21ai_1 _0851_ (.B1(_0228_),
    .VDD(VPWR),
    .Y(UI_IN_TT_PROJECT4),
    .VSS(VGND),
    .A1(_0229_),
    .A2(_0231_));
 sg13g2_mux4_1 _0852_ (.S0(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit24.Q ),
    .A0(Tile_X0Y1_E1END[1]),
    .A1(Tile_X0Y1_EE4END[13]),
    .A2(Tile_X0Y1_EE4END[5]),
    .A3(Tile_X0Y1_E6END[5]),
    .S1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit23.Q ),
    .X(_0232_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _0853_ (.Y(_0233_),
    .B(_0232_),
    .A_N(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit25.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _0854_ (.Y(_0234_),
    .B(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit25.Q ),
    .A_N(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit24.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _0855_ (.Y(_0235_),
    .B(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit23.Q ),
    .A_N(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.J_NS4_BEG13 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _0856_ (.B1(_0235_),
    .VDD(VPWR),
    .Y(_0236_),
    .VSS(VGND),
    .A1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit23.Q ),
    .A2(_0153_));
 sg13g2_o21ai_1 _0857_ (.B1(_0233_),
    .VDD(VPWR),
    .Y(UI_IN_TT_PROJECT5),
    .VSS(VGND),
    .A1(_0234_),
    .A2(_0236_));
 sg13g2_nand2b_1 _0858_ (.Y(_0237_),
    .B(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit28.Q ),
    .A_N(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit27.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _0859_ (.Y(_0238_),
    .B(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit26.Q ),
    .A_N(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.J_NS4_BEG14 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _0860_ (.B1(_0238_),
    .VDD(VPWR),
    .Y(_0239_),
    .VSS(VGND),
    .A1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit26.Q ),
    .A2(_0152_));
 sg13g2_mux4_1 _0861_ (.S0(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit27.Q ),
    .A0(Tile_X0Y1_E1END[2]),
    .A1(Tile_X0Y1_EE4END[14]),
    .A2(Tile_X0Y1_EE4END[6]),
    .A3(Tile_X0Y1_E6END[6]),
    .S1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit26.Q ),
    .X(_0240_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _0862_ (.Y(_0241_),
    .B(_0240_),
    .A_N(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit28.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _0863_ (.B1(_0241_),
    .VDD(VPWR),
    .Y(UI_IN_TT_PROJECT6),
    .VSS(VGND),
    .A1(_0237_),
    .A2(_0239_));
 sg13g2_mux4_1 _0864_ (.S0(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit30.Q ),
    .A0(Tile_X0Y1_E1END[3]),
    .A1(Tile_X0Y1_EE4END[15]),
    .A2(Tile_X0Y1_EE4END[7]),
    .A3(Tile_X0Y1_E6END[7]),
    .S1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit29.Q ),
    .X(_0242_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _0865_ (.Y(_0243_),
    .B(_0242_),
    .A_N(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit31.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _0866_ (.Y(_0244_),
    .B(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit31.Q ),
    .A_N(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit30.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _0867_ (.Y(_0245_),
    .B(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit29.Q ),
    .A_N(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.J_NS4_BEG15 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _0868_ (.B1(_0245_),
    .VDD(VPWR),
    .Y(_0246_),
    .VSS(VGND),
    .A1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit29.Q ),
    .A2(_0151_));
 sg13g2_o21ai_1 _0869_ (.B1(_0243_),
    .VDD(VPWR),
    .Y(UI_IN_TT_PROJECT7),
    .VSS(VGND),
    .A1(_0244_),
    .A2(_0246_));
 sg13g2_nor2b_1 _0870_ (.A(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit0.Q ),
    .B_N(Tile_X0Y1_E2MID[3]),
    .Y(_0247_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _0871_ (.A(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit1.Q ),
    .B(_0306_),
    .Y(_0248_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _0872_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(Tile_X0Y1_E2MID[6]),
    .A2(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit0.Q ),
    .Y(_0249_),
    .B1(_0247_));
 sg13g2_mux2_1 _0873_ (.A0(Tile_X0Y1_N2MID[6]),
    .A1(Tile_X0Y1_N2END[2]),
    .S(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit0.Q ),
    .X(_0250_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _0874_ (.A(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit1.Q ),
    .B(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit2.Q ),
    .C(_0250_),
    .Y(_0251_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _0875_ (.S0(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit2.Q ),
    .A0(Tile_X0Y1_N2END[3]),
    .A1(Tile_X0Y1_E2END[1]),
    .A2(Tile_X0Y1_E2MID[0]),
    .A3(Tile_X0Y1_E2END[2]),
    .S1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit0.Q ),
    .X(_0252_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _0876_ (.VDD(VPWR),
    .Y(_0253_),
    .A(_0252_),
    .VSS(VGND));
 sg13g2_a221oi_1 _0877_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit1.Q ),
    .C1(_0251_),
    .B1(_0253_),
    .A1(_0248_),
    .Y(_0254_),
    .A2(_0249_));
 sg13g2_nor3_1 _0878_ (.A(_0305_),
    .B(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit2.Q ),
    .C(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.S2BEG0 ),
    .Y(_0255_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _0879_ (.A0(Tile_X0Y1_E2END[4]),
    .A1(Tile_X0Y0_S2MID[3]),
    .S(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit2.Q ),
    .X(_0256_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _0880_ (.B1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit0.Q ),
    .VDD(VPWR),
    .Y(_0257_),
    .VSS(VGND),
    .A1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit1.Q ),
    .A2(_0256_));
 sg13g2_nand2b_1 _0881_ (.Y(_0258_),
    .B(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit2.Q ),
    .A_N(Tile_X0Y0_S2MID[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _0882_ (.Y(_0259_),
    .B1(_0258_),
    .B2(_0305_),
    .A2(_0306_),
    .A1(Tile_X0Y1_E2END[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _0883_ (.A(Tile_X0Y1_E2END[3]),
    .B(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit1.Q ),
    .C(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit2.Q ),
    .Y(_0260_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _0884_ (.A(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit0.Q ),
    .B(_0259_),
    .C(_0260_),
    .Y(_0261_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _0885_ (.A(_0261_),
    .B_N(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit3.Q ),
    .Y(_0262_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _0886_ (.B1(_0262_),
    .VDD(VPWR),
    .Y(_0263_),
    .VSS(VGND),
    .A1(_0255_),
    .A2(_0257_));
 sg13g2_o21ai_1 _0887_ (.B1(_0263_),
    .VDD(VPWR),
    .Y(_0264_),
    .VSS(VGND),
    .A1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit3.Q ),
    .A2(_0254_));
 sg13g2_inv_1 _0888_ (.VDD(VPWR),
    .Y(ENA_TT_PROJECT),
    .A(_0264_),
    .VSS(VGND));
 sg13g2_nor2b_1 _0889_ (.A(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit6.Q ),
    .B_N(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit5.Q ),
    .Y(_0265_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _0890_ (.A(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit5.Q ),
    .B_N(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit6.Q ),
    .Y(_0266_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _0891_ (.A(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit4.Q ),
    .B_N(Tile_X0Y1_E2END[1]),
    .Y(_0267_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _0892_ (.Y(_0268_),
    .A(Tile_X0Y1_E2END[2]),
    .B(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit4.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _0893_ (.B(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit6.Q ),
    .C(_0268_),
    .A(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit5.Q ),
    .Y(_0269_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _0894_ (.A0(Tile_X0Y1_N2MID[6]),
    .A1(Tile_X0Y1_N2END[2]),
    .S(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit4.Q ),
    .X(_0270_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _0895_ (.A(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit5.Q ),
    .B(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit6.Q ),
    .C(_0270_),
    .Y(_0271_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _0896_ (.A(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit4.Q ),
    .B_N(Tile_X0Y1_E2MID[3]),
    .Y(_0272_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _0897_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(Tile_X0Y1_E2MID[6]),
    .A2(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit4.Q ),
    .Y(_0273_),
    .B1(_0272_));
 sg13g2_nor2b_1 _0898_ (.A(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit4.Q ),
    .B_N(Tile_X0Y1_N2END[3]),
    .Y(_0274_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _0899_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(Tile_X0Y1_E2MID[0]),
    .A2(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit4.Q ),
    .Y(_0275_),
    .B1(_0274_));
 sg13g2_a221oi_1 _0900_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_0265_),
    .C1(_0271_),
    .B1(_0275_),
    .A1(_0266_),
    .Y(_0276_),
    .A2(_0273_));
 sg13g2_o21ai_1 _0901_ (.B1(_0276_),
    .VDD(VPWR),
    .Y(_0277_),
    .VSS(VGND),
    .A1(_0267_),
    .A2(_0269_));
 sg13g2_nand2b_1 _0902_ (.Y(_0278_),
    .B(_0265_),
    .A_N(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.S2BEG0 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _0903_ (.A(Tile_X0Y1_E2END[4]),
    .B(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit5.Q ),
    .C(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit6.Q ),
    .Y(_0279_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _0904_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0296_),
    .A2(_0266_),
    .Y(_0280_),
    .B1(_0279_));
 sg13g2_nand3_1 _0905_ (.B(_0278_),
    .C(_0280_),
    .A(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit4.Q ),
    .Y(_0281_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _0906_ (.A(Tile_X0Y1_E2END[3]),
    .B(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit5.Q ),
    .C(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit6.Q ),
    .Y(_0282_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _0907_ (.B1(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit5.Q ),
    .VDD(VPWR),
    .Y(_0283_),
    .VSS(VGND),
    .A1(_0295_),
    .A2(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit6.Q ));
 sg13g2_nor2b_1 _0908_ (.A(Tile_X0Y0_S2MID[2]),
    .B_N(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit6.Q ),
    .Y(_0284_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _0909_ (.A(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit4.Q ),
    .B(_0282_),
    .C(_0284_),
    .Y(_0285_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _0910_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0283_),
    .A2(_0285_),
    .Y(_0286_),
    .B1(_0307_));
 sg13g2_a22oi_1 _0911_ (.Y(RST_N_TT_PROJECT),
    .B1(_0281_),
    .B2(_0286_),
    .A2(_0277_),
    .A1(_0307_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _0912_ (.D(Tile_X0Y0_FrameData[31]),
    .GATE(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit31.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _0913_ (.D(Tile_X0Y0_FrameData[30]),
    .GATE(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit30.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _0914_ (.D(Tile_X0Y0_FrameData[29]),
    .GATE(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit29.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _0915_ (.D(Tile_X0Y0_FrameData[28]),
    .GATE(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit28.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _0916_ (.D(Tile_X0Y0_FrameData[27]),
    .GATE(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit27.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _0917_ (.D(Tile_X0Y0_FrameData[26]),
    .GATE(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit26.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _0918_ (.D(Tile_X0Y0_FrameData[25]),
    .GATE(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit25.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _0919_ (.D(Tile_X0Y0_FrameData[24]),
    .GATE(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit24.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _0920_ (.D(Tile_X0Y0_FrameData[23]),
    .GATE(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit23.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _0921_ (.D(Tile_X0Y0_FrameData[22]),
    .GATE(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit22.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _0922_ (.D(Tile_X0Y0_FrameData[21]),
    .GATE(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit21.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _0923_ (.D(Tile_X0Y0_FrameData[20]),
    .GATE(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit20.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _0924_ (.D(Tile_X0Y0_FrameData[19]),
    .GATE(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit19.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _0925_ (.D(Tile_X0Y0_FrameData[18]),
    .GATE(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit18.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _0926_ (.D(Tile_X0Y0_FrameData[17]),
    .GATE(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit17.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _0927_ (.D(Tile_X0Y0_FrameData[16]),
    .GATE(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit16.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _0928_ (.D(Tile_X0Y0_FrameData[15]),
    .GATE(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit15.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _0929_ (.D(Tile_X0Y0_FrameData[14]),
    .GATE(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit14.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _0930_ (.D(Tile_X0Y0_FrameData[13]),
    .GATE(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit13.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _0931_ (.D(Tile_X0Y0_FrameData[12]),
    .GATE(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit12.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _0932_ (.D(Tile_X0Y0_FrameData[11]),
    .GATE(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit11.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _0933_ (.D(Tile_X0Y0_FrameData[10]),
    .GATE(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit10.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _0934_ (.D(Tile_X0Y0_FrameData[9]),
    .GATE(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit9.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _0935_ (.D(Tile_X0Y0_FrameData[8]),
    .GATE(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit8.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _0936_ (.D(Tile_X0Y0_FrameData[7]),
    .GATE(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit7.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _0937_ (.D(Tile_X0Y0_FrameData[6]),
    .GATE(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit6.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _0938_ (.D(Tile_X0Y0_FrameData[5]),
    .GATE(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit5.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _0939_ (.D(Tile_X0Y0_FrameData[4]),
    .GATE(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit4.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _0940_ (.D(Tile_X0Y0_FrameData[3]),
    .GATE(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit3.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _0941_ (.D(Tile_X0Y0_FrameData[2]),
    .GATE(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit2.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _0942_ (.D(Tile_X0Y0_FrameData[1]),
    .GATE(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit1.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _0943_ (.D(Tile_X0Y0_FrameData[0]),
    .GATE(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit0.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _0944_ (.D(Tile_X0Y0_FrameData[31]),
    .GATE(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit31.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _0945_ (.D(Tile_X0Y0_FrameData[30]),
    .GATE(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit30.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _0946_ (.D(Tile_X0Y0_FrameData[29]),
    .GATE(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit29.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _0947_ (.D(Tile_X0Y0_FrameData[28]),
    .GATE(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit28.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _0948_ (.D(Tile_X0Y0_FrameData[27]),
    .GATE(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit27.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _0949_ (.D(Tile_X0Y0_FrameData[26]),
    .GATE(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit26.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _0950_ (.D(Tile_X0Y0_FrameData[25]),
    .GATE(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit25.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _0951_ (.D(Tile_X0Y0_FrameData[24]),
    .GATE(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit24.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _0952_ (.D(Tile_X0Y0_FrameData[23]),
    .GATE(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit23.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _0953_ (.D(Tile_X0Y0_FrameData[22]),
    .GATE(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit22.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _0954_ (.D(Tile_X0Y0_FrameData[21]),
    .GATE(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit21.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _0955_ (.D(Tile_X0Y0_FrameData[20]),
    .GATE(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit20.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _0956_ (.D(Tile_X0Y0_FrameData[19]),
    .GATE(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit19.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _0957_ (.D(Tile_X0Y0_FrameData[18]),
    .GATE(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit18.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _0958_ (.D(Tile_X0Y0_FrameData[17]),
    .GATE(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit17.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _0959_ (.D(Tile_X0Y0_FrameData[16]),
    .GATE(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit16.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _0960_ (.D(Tile_X0Y0_FrameData[15]),
    .GATE(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit15.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _0961_ (.D(Tile_X0Y0_FrameData[14]),
    .GATE(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit14.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _0962_ (.D(Tile_X0Y0_FrameData[13]),
    .GATE(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit13.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _0963_ (.D(Tile_X0Y0_FrameData[12]),
    .GATE(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit12.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _0964_ (.D(Tile_X0Y0_FrameData[11]),
    .GATE(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit11.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _0965_ (.D(Tile_X0Y0_FrameData[10]),
    .GATE(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit10.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _0966_ (.D(Tile_X0Y0_FrameData[9]),
    .GATE(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit9.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _0967_ (.D(Tile_X0Y0_FrameData[8]),
    .GATE(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit8.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _0968_ (.D(Tile_X0Y0_FrameData[7]),
    .GATE(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit7.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _0969_ (.D(Tile_X0Y0_FrameData[6]),
    .GATE(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit6.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _0970_ (.D(Tile_X0Y0_FrameData[5]),
    .GATE(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit5.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _0971_ (.D(Tile_X0Y0_FrameData[4]),
    .GATE(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit4.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _0972_ (.D(Tile_X0Y0_FrameData[3]),
    .GATE(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit3.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _0973_ (.D(Tile_X0Y0_FrameData[2]),
    .GATE(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit2.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _0974_ (.D(Tile_X0Y0_FrameData[1]),
    .GATE(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit1.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _0975_ (.D(Tile_X0Y0_FrameData[0]),
    .GATE(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit0.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _0976_ (.D(Tile_X0Y0_FrameData[31]),
    .GATE(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit31.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _0977_ (.D(Tile_X0Y0_FrameData[30]),
    .GATE(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit30.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _0978_ (.D(Tile_X0Y0_FrameData[29]),
    .GATE(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit29.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _0979_ (.D(Tile_X0Y0_FrameData[28]),
    .GATE(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit28.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _0980_ (.D(Tile_X0Y0_FrameData[27]),
    .GATE(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit27.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _0981_ (.D(Tile_X0Y0_FrameData[26]),
    .GATE(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit26.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _0982_ (.D(Tile_X0Y0_FrameData[25]),
    .GATE(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit25.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _0983_ (.D(Tile_X0Y0_FrameData[24]),
    .GATE(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit24.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _0984_ (.D(Tile_X0Y0_FrameData[23]),
    .GATE(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit23.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _0985_ (.D(Tile_X0Y0_FrameData[22]),
    .GATE(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit22.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _0986_ (.D(Tile_X0Y0_FrameData[21]),
    .GATE(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit21.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _0987_ (.D(Tile_X0Y0_FrameData[20]),
    .GATE(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit20.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _0988_ (.D(Tile_X0Y0_FrameData[19]),
    .GATE(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit19.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _0989_ (.D(Tile_X0Y0_FrameData[18]),
    .GATE(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit18.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _0990_ (.D(Tile_X0Y0_FrameData[17]),
    .GATE(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit17.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _0991_ (.D(Tile_X0Y0_FrameData[16]),
    .GATE(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit16.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _0992_ (.D(Tile_X0Y0_FrameData[15]),
    .GATE(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit15.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _0993_ (.D(Tile_X0Y0_FrameData[14]),
    .GATE(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit14.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _0994_ (.D(Tile_X0Y0_FrameData[13]),
    .GATE(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit13.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _0995_ (.D(Tile_X0Y0_FrameData[12]),
    .GATE(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit12.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _0996_ (.D(Tile_X0Y0_FrameData[11]),
    .GATE(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit11.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _0997_ (.D(Tile_X0Y0_FrameData[10]),
    .GATE(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit10.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _0998_ (.D(Tile_X0Y0_FrameData[9]),
    .GATE(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit9.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _0999_ (.D(Tile_X0Y0_FrameData[8]),
    .GATE(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit8.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1000_ (.D(Tile_X0Y0_FrameData[7]),
    .GATE(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit7.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1001_ (.D(Tile_X0Y0_FrameData[6]),
    .GATE(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit6.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1002_ (.D(Tile_X0Y0_FrameData[5]),
    .GATE(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit5.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1003_ (.D(Tile_X0Y0_FrameData[4]),
    .GATE(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit4.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1004_ (.D(Tile_X0Y0_FrameData[3]),
    .GATE(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit3.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1005_ (.D(Tile_X0Y0_FrameData[2]),
    .GATE(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit2.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1006_ (.D(Tile_X0Y0_FrameData[1]),
    .GATE(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit1.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1007_ (.D(Tile_X0Y0_FrameData[0]),
    .GATE(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit0.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1008_ (.D(Tile_X0Y0_FrameData[31]),
    .GATE(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit31.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1009_ (.D(Tile_X0Y0_FrameData[30]),
    .GATE(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit30.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1010_ (.D(Tile_X0Y0_FrameData[29]),
    .GATE(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit29.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1011_ (.D(Tile_X0Y0_FrameData[28]),
    .GATE(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit28.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1012_ (.D(Tile_X0Y0_FrameData[27]),
    .GATE(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit27.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1013_ (.D(Tile_X0Y0_FrameData[26]),
    .GATE(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit26.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1014_ (.D(Tile_X0Y0_FrameData[25]),
    .GATE(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit25.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1015_ (.D(Tile_X0Y0_FrameData[24]),
    .GATE(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit24.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1016_ (.D(Tile_X0Y0_FrameData[23]),
    .GATE(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit23.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1017_ (.D(Tile_X0Y0_FrameData[22]),
    .GATE(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit22.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1018_ (.D(Tile_X0Y0_FrameData[21]),
    .GATE(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit21.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1019_ (.D(Tile_X0Y0_FrameData[20]),
    .GATE(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit20.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1020_ (.D(Tile_X0Y0_FrameData[19]),
    .GATE(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit19.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1021_ (.D(Tile_X0Y0_FrameData[18]),
    .GATE(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit18.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1022_ (.D(Tile_X0Y0_FrameData[17]),
    .GATE(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit17.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1023_ (.D(Tile_X0Y0_FrameData[16]),
    .GATE(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit16.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1024_ (.D(Tile_X0Y0_FrameData[15]),
    .GATE(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit15.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1025_ (.D(Tile_X0Y0_FrameData[14]),
    .GATE(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit14.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1026_ (.D(Tile_X0Y0_FrameData[13]),
    .GATE(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit13.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1027_ (.D(Tile_X0Y0_FrameData[12]),
    .GATE(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit12.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1028_ (.D(Tile_X0Y0_FrameData[11]),
    .GATE(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit11.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1029_ (.D(Tile_X0Y0_FrameData[10]),
    .GATE(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit10.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1030_ (.D(Tile_X0Y0_FrameData[9]),
    .GATE(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit9.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1031_ (.D(Tile_X0Y0_FrameData[8]),
    .GATE(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit8.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1032_ (.D(Tile_X0Y0_FrameData[7]),
    .GATE(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit7.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1033_ (.D(Tile_X0Y0_FrameData[6]),
    .GATE(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit6.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1034_ (.D(Tile_X0Y0_FrameData[5]),
    .GATE(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit5.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1035_ (.D(Tile_X0Y0_FrameData[4]),
    .GATE(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit4.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1036_ (.D(Tile_X0Y0_FrameData[3]),
    .GATE(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit3.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1037_ (.D(Tile_X0Y0_FrameData[2]),
    .GATE(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit2.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1038_ (.D(Tile_X0Y0_FrameData[1]),
    .GATE(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit1.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1039_ (.D(Tile_X0Y0_FrameData[0]),
    .GATE(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit0.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1040_ (.D(Tile_X0Y0_FrameData[31]),
    .GATE(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit31.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1041_ (.D(Tile_X0Y0_FrameData[30]),
    .GATE(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit30.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1042_ (.D(Tile_X0Y0_FrameData[29]),
    .GATE(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit29.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1043_ (.D(Tile_X0Y0_FrameData[28]),
    .GATE(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit28.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1044_ (.D(Tile_X0Y0_FrameData[27]),
    .GATE(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit27.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1045_ (.D(Tile_X0Y0_FrameData[26]),
    .GATE(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit26.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1046_ (.D(Tile_X0Y0_FrameData[25]),
    .GATE(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit25.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1047_ (.D(Tile_X0Y0_FrameData[24]),
    .GATE(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit24.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1048_ (.D(Tile_X0Y0_FrameData[23]),
    .GATE(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit23.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1049_ (.D(Tile_X0Y0_FrameData[22]),
    .GATE(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit22.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1050_ (.D(Tile_X0Y0_FrameData[21]),
    .GATE(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit21.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1051_ (.D(Tile_X0Y0_FrameData[20]),
    .GATE(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit20.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1052_ (.D(Tile_X0Y0_FrameData[19]),
    .GATE(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit19.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1053_ (.D(Tile_X0Y0_FrameData[18]),
    .GATE(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit18.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1054_ (.D(Tile_X0Y0_FrameData[17]),
    .GATE(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit17.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1055_ (.D(Tile_X0Y0_FrameData[16]),
    .GATE(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit16.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1056_ (.D(Tile_X0Y0_FrameData[15]),
    .GATE(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit15.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1057_ (.D(Tile_X0Y0_FrameData[14]),
    .GATE(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit14.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1058_ (.D(Tile_X0Y0_FrameData[13]),
    .GATE(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit13.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1059_ (.D(Tile_X0Y0_FrameData[12]),
    .GATE(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit12.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1060_ (.D(Tile_X0Y0_FrameData[11]),
    .GATE(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit11.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1061_ (.D(Tile_X0Y0_FrameData[10]),
    .GATE(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit10.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1062_ (.D(Tile_X0Y0_FrameData[9]),
    .GATE(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit9.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1063_ (.D(Tile_X0Y0_FrameData[8]),
    .GATE(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit8.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1064_ (.D(Tile_X0Y0_FrameData[7]),
    .GATE(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit7.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1065_ (.D(Tile_X0Y0_FrameData[6]),
    .GATE(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit6.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1066_ (.D(Tile_X0Y0_FrameData[5]),
    .GATE(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit5.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1067_ (.D(Tile_X0Y0_FrameData[4]),
    .GATE(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit4.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1068_ (.D(Tile_X0Y0_FrameData[3]),
    .GATE(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit3.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1069_ (.D(Tile_X0Y0_FrameData[2]),
    .GATE(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit2.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1070_ (.D(Tile_X0Y0_FrameData[1]),
    .GATE(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit1.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1071_ (.D(Tile_X0Y0_FrameData[0]),
    .GATE(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit0.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1072_ (.D(Tile_X0Y0_FrameData[31]),
    .GATE(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit31.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1073_ (.D(Tile_X0Y0_FrameData[30]),
    .GATE(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit30.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1074_ (.D(Tile_X0Y0_FrameData[29]),
    .GATE(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit29.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1075_ (.D(Tile_X0Y0_FrameData[28]),
    .GATE(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit28.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1076_ (.D(Tile_X0Y0_FrameData[27]),
    .GATE(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit27.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1077_ (.D(Tile_X0Y0_FrameData[26]),
    .GATE(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit26.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1078_ (.D(Tile_X0Y0_FrameData[25]),
    .GATE(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit25.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1079_ (.D(Tile_X0Y0_FrameData[24]),
    .GATE(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit24.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1080_ (.D(Tile_X0Y0_FrameData[23]),
    .GATE(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit23.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1081_ (.D(Tile_X0Y0_FrameData[22]),
    .GATE(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit22.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1082_ (.D(Tile_X0Y0_FrameData[21]),
    .GATE(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit21.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1083_ (.D(Tile_X0Y0_FrameData[20]),
    .GATE(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit20.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1084_ (.D(Tile_X0Y0_FrameData[19]),
    .GATE(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit19.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1085_ (.D(Tile_X0Y0_FrameData[18]),
    .GATE(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit18.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1086_ (.D(Tile_X0Y0_FrameData[17]),
    .GATE(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit17.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1087_ (.D(Tile_X0Y0_FrameData[16]),
    .GATE(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit16.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1088_ (.D(Tile_X0Y0_FrameData[15]),
    .GATE(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit15.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1089_ (.D(Tile_X0Y0_FrameData[14]),
    .GATE(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit14.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1090_ (.D(Tile_X0Y0_FrameData[13]),
    .GATE(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit13.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1091_ (.D(Tile_X0Y0_FrameData[12]),
    .GATE(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit12.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1092_ (.D(Tile_X0Y0_FrameData[11]),
    .GATE(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit11.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1093_ (.D(Tile_X0Y0_FrameData[10]),
    .GATE(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit10.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1094_ (.D(Tile_X0Y0_FrameData[9]),
    .GATE(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit9.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1095_ (.D(Tile_X0Y0_FrameData[8]),
    .GATE(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit8.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1096_ (.D(Tile_X0Y0_FrameData[7]),
    .GATE(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit7.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1097_ (.D(Tile_X0Y0_FrameData[6]),
    .GATE(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit6.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1098_ (.D(Tile_X0Y0_FrameData[5]),
    .GATE(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit5.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1099_ (.D(Tile_X0Y0_FrameData[4]),
    .GATE(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit4.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1100_ (.D(Tile_X0Y0_FrameData[3]),
    .GATE(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit3.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1101_ (.D(Tile_X0Y0_FrameData[2]),
    .GATE(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit2.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1102_ (.D(Tile_X0Y0_FrameData[1]),
    .GATE(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit1.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1103_ (.D(Tile_X0Y0_FrameData[0]),
    .GATE(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit0.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1104_ (.D(Tile_X0Y0_FrameData[31]),
    .GATE(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit31.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1105_ (.D(Tile_X0Y0_FrameData[30]),
    .GATE(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit30.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1106_ (.D(Tile_X0Y0_FrameData[29]),
    .GATE(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit29.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1107_ (.D(Tile_X0Y0_FrameData[28]),
    .GATE(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit28.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1108_ (.D(Tile_X0Y0_FrameData[27]),
    .GATE(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit27.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1109_ (.D(Tile_X0Y0_FrameData[26]),
    .GATE(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit26.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1110_ (.D(Tile_X0Y0_FrameData[25]),
    .GATE(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit25.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1111_ (.D(Tile_X0Y0_FrameData[24]),
    .GATE(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit24.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1112_ (.D(Tile_X0Y0_FrameData[23]),
    .GATE(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit23.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1113_ (.D(Tile_X0Y0_FrameData[22]),
    .GATE(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit22.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1114_ (.D(Tile_X0Y0_FrameData[21]),
    .GATE(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit21.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1115_ (.D(Tile_X0Y0_FrameData[20]),
    .GATE(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit20.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1116_ (.D(Tile_X0Y0_FrameData[19]),
    .GATE(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit19.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1117_ (.D(Tile_X0Y0_FrameData[18]),
    .GATE(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit18.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1118_ (.D(Tile_X0Y0_FrameData[17]),
    .GATE(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit17.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1119_ (.D(Tile_X0Y0_FrameData[16]),
    .GATE(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit16.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1120_ (.D(Tile_X0Y0_FrameData[15]),
    .GATE(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit15.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1121_ (.D(Tile_X0Y0_FrameData[14]),
    .GATE(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit14.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1122_ (.D(Tile_X0Y0_FrameData[13]),
    .GATE(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit13.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1123_ (.D(Tile_X0Y0_FrameData[12]),
    .GATE(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit12.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1124_ (.D(Tile_X0Y0_FrameData[11]),
    .GATE(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit11.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1125_ (.D(Tile_X0Y0_FrameData[10]),
    .GATE(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit10.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1126_ (.D(Tile_X0Y0_FrameData[9]),
    .GATE(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit9.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1127_ (.D(Tile_X0Y0_FrameData[8]),
    .GATE(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit8.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1128_ (.D(Tile_X0Y0_FrameData[7]),
    .GATE(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit7.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1129_ (.D(Tile_X0Y0_FrameData[6]),
    .GATE(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit6.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1130_ (.D(Tile_X0Y0_FrameData[5]),
    .GATE(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit5.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1131_ (.D(Tile_X0Y0_FrameData[4]),
    .GATE(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit4.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1132_ (.D(Tile_X0Y0_FrameData[3]),
    .GATE(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit3.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1133_ (.D(Tile_X0Y0_FrameData[2]),
    .GATE(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit2.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1134_ (.D(Tile_X0Y0_FrameData[1]),
    .GATE(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit1.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1135_ (.D(Tile_X0Y0_FrameData[0]),
    .GATE(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit0.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1136_ (.D(Tile_X0Y0_FrameData[31]),
    .GATE(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit31.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1137_ (.D(Tile_X0Y0_FrameData[30]),
    .GATE(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit30.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1138_ (.D(Tile_X0Y0_FrameData[29]),
    .GATE(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit29.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1139_ (.D(Tile_X0Y0_FrameData[28]),
    .GATE(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit28.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1140_ (.D(Tile_X0Y0_FrameData[27]),
    .GATE(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit27.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1141_ (.D(Tile_X0Y0_FrameData[26]),
    .GATE(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit26.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1142_ (.D(Tile_X0Y0_FrameData[25]),
    .GATE(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit25.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1143_ (.D(Tile_X0Y0_FrameData[24]),
    .GATE(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit24.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1144_ (.D(Tile_X0Y0_FrameData[23]),
    .GATE(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit23.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1145_ (.D(Tile_X0Y0_FrameData[22]),
    .GATE(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit22.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1146_ (.D(Tile_X0Y0_FrameData[21]),
    .GATE(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit21.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1147_ (.D(Tile_X0Y0_FrameData[20]),
    .GATE(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit20.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1148_ (.D(Tile_X0Y0_FrameData[19]),
    .GATE(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit19.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1149_ (.D(Tile_X0Y0_FrameData[18]),
    .GATE(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit18.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1150_ (.D(Tile_X0Y0_FrameData[17]),
    .GATE(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit17.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1151_ (.D(Tile_X0Y0_FrameData[16]),
    .GATE(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit16.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1152_ (.D(Tile_X0Y0_FrameData[15]),
    .GATE(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit15.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1153_ (.D(Tile_X0Y0_FrameData[14]),
    .GATE(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit14.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1154_ (.D(Tile_X0Y0_FrameData[13]),
    .GATE(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit13.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1155_ (.D(Tile_X0Y0_FrameData[12]),
    .GATE(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit12.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1156_ (.D(Tile_X0Y0_FrameData[11]),
    .GATE(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit11.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1157_ (.D(Tile_X0Y0_FrameData[10]),
    .GATE(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit10.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1158_ (.D(Tile_X0Y0_FrameData[9]),
    .GATE(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit9.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1159_ (.D(Tile_X0Y0_FrameData[8]),
    .GATE(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit8.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1160_ (.D(Tile_X0Y1_FrameData[31]),
    .GATE(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit31.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1161_ (.D(Tile_X0Y1_FrameData[30]),
    .GATE(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit30.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1162_ (.D(Tile_X0Y1_FrameData[29]),
    .GATE(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit29.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1163_ (.D(Tile_X0Y1_FrameData[28]),
    .GATE(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit28.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1164_ (.D(Tile_X0Y1_FrameData[27]),
    .GATE(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit27.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1165_ (.D(Tile_X0Y1_FrameData[26]),
    .GATE(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit26.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1166_ (.D(Tile_X0Y1_FrameData[25]),
    .GATE(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit25.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1167_ (.D(Tile_X0Y1_FrameData[24]),
    .GATE(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit24.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1168_ (.D(Tile_X0Y1_FrameData[23]),
    .GATE(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit23.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1169_ (.D(Tile_X0Y1_FrameData[22]),
    .GATE(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit22.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1170_ (.D(Tile_X0Y1_FrameData[21]),
    .GATE(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit21.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1171_ (.D(Tile_X0Y1_FrameData[20]),
    .GATE(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit20.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1172_ (.D(Tile_X0Y1_FrameData[19]),
    .GATE(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit19.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1173_ (.D(Tile_X0Y1_FrameData[18]),
    .GATE(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit18.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1174_ (.D(Tile_X0Y1_FrameData[17]),
    .GATE(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit17.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1175_ (.D(Tile_X0Y1_FrameData[16]),
    .GATE(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit16.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1176_ (.D(Tile_X0Y1_FrameData[15]),
    .GATE(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit15.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1177_ (.D(Tile_X0Y1_FrameData[14]),
    .GATE(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit14.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1178_ (.D(Tile_X0Y1_FrameData[13]),
    .GATE(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit13.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1179_ (.D(Tile_X0Y1_FrameData[12]),
    .GATE(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit12.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1180_ (.D(Tile_X0Y1_FrameData[11]),
    .GATE(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit11.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1181_ (.D(Tile_X0Y1_FrameData[10]),
    .GATE(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit10.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1182_ (.D(Tile_X0Y1_FrameData[9]),
    .GATE(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit9.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1183_ (.D(Tile_X0Y1_FrameData[8]),
    .GATE(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit8.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1184_ (.D(Tile_X0Y1_FrameData[7]),
    .GATE(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit7.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1185_ (.D(Tile_X0Y1_FrameData[6]),
    .GATE(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit6.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1186_ (.D(Tile_X0Y1_FrameData[5]),
    .GATE(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit5.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1187_ (.D(Tile_X0Y1_FrameData[4]),
    .GATE(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit4.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1188_ (.D(Tile_X0Y1_FrameData[3]),
    .GATE(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit3.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1189_ (.D(Tile_X0Y1_FrameData[2]),
    .GATE(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit2.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1190_ (.D(Tile_X0Y1_FrameData[1]),
    .GATE(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit1.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1191_ (.D(Tile_X0Y1_FrameData[0]),
    .GATE(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit0.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1192_ (.D(Tile_X0Y1_FrameData[31]),
    .GATE(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit31.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1193_ (.D(Tile_X0Y1_FrameData[30]),
    .GATE(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit30.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1194_ (.D(Tile_X0Y1_FrameData[29]),
    .GATE(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit29.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1195_ (.D(Tile_X0Y1_FrameData[28]),
    .GATE(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit28.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1196_ (.D(Tile_X0Y1_FrameData[27]),
    .GATE(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit27.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1197_ (.D(Tile_X0Y1_FrameData[26]),
    .GATE(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit26.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1198_ (.D(Tile_X0Y1_FrameData[25]),
    .GATE(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit25.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1199_ (.D(Tile_X0Y1_FrameData[24]),
    .GATE(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit24.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1200_ (.D(Tile_X0Y1_FrameData[23]),
    .GATE(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit23.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1201_ (.D(Tile_X0Y1_FrameData[22]),
    .GATE(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit22.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1202_ (.D(Tile_X0Y1_FrameData[21]),
    .GATE(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit21.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1203_ (.D(Tile_X0Y1_FrameData[20]),
    .GATE(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit20.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1204_ (.D(Tile_X0Y1_FrameData[19]),
    .GATE(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit19.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1205_ (.D(Tile_X0Y1_FrameData[18]),
    .GATE(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit18.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1206_ (.D(Tile_X0Y1_FrameData[17]),
    .GATE(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit17.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1207_ (.D(Tile_X0Y1_FrameData[16]),
    .GATE(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit16.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1208_ (.D(Tile_X0Y1_FrameData[15]),
    .GATE(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit15.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1209_ (.D(Tile_X0Y1_FrameData[14]),
    .GATE(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit14.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1210_ (.D(Tile_X0Y1_FrameData[13]),
    .GATE(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit13.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1211_ (.D(Tile_X0Y1_FrameData[12]),
    .GATE(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit12.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1212_ (.D(Tile_X0Y1_FrameData[11]),
    .GATE(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit11.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1213_ (.D(Tile_X0Y1_FrameData[10]),
    .GATE(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit10.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1214_ (.D(Tile_X0Y1_FrameData[9]),
    .GATE(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit9.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1215_ (.D(Tile_X0Y1_FrameData[8]),
    .GATE(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit8.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1216_ (.D(Tile_X0Y1_FrameData[7]),
    .GATE(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit7.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1217_ (.D(Tile_X0Y1_FrameData[6]),
    .GATE(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit6.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1218_ (.D(Tile_X0Y1_FrameData[5]),
    .GATE(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit5.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1219_ (.D(Tile_X0Y1_FrameData[4]),
    .GATE(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit4.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1220_ (.D(Tile_X0Y1_FrameData[3]),
    .GATE(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit3.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1221_ (.D(Tile_X0Y1_FrameData[2]),
    .GATE(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit2.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1222_ (.D(Tile_X0Y1_FrameData[1]),
    .GATE(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit1.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1223_ (.D(Tile_X0Y1_FrameData[0]),
    .GATE(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit0.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1224_ (.D(Tile_X0Y1_FrameData[31]),
    .GATE(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit31.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1225_ (.D(Tile_X0Y1_FrameData[30]),
    .GATE(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit30.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1226_ (.D(Tile_X0Y1_FrameData[29]),
    .GATE(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit29.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1227_ (.D(Tile_X0Y1_FrameData[28]),
    .GATE(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit28.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1228_ (.D(Tile_X0Y1_FrameData[27]),
    .GATE(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit27.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1229_ (.D(Tile_X0Y1_FrameData[26]),
    .GATE(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit26.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1230_ (.D(Tile_X0Y1_FrameData[25]),
    .GATE(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit25.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1231_ (.D(Tile_X0Y1_FrameData[24]),
    .GATE(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit24.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1232_ (.D(Tile_X0Y1_FrameData[23]),
    .GATE(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit23.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1233_ (.D(Tile_X0Y1_FrameData[22]),
    .GATE(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit22.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1234_ (.D(Tile_X0Y1_FrameData[21]),
    .GATE(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit21.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1235_ (.D(Tile_X0Y1_FrameData[20]),
    .GATE(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit20.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1236_ (.D(Tile_X0Y1_FrameData[19]),
    .GATE(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit19.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1237_ (.D(Tile_X0Y1_FrameData[18]),
    .GATE(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit18.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1238_ (.D(Tile_X0Y1_FrameData[17]),
    .GATE(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit17.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1239_ (.D(Tile_X0Y1_FrameData[16]),
    .GATE(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit16.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1240_ (.D(Tile_X0Y1_FrameData[15]),
    .GATE(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit15.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1241_ (.D(Tile_X0Y1_FrameData[14]),
    .GATE(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit14.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1242_ (.D(Tile_X0Y1_FrameData[13]),
    .GATE(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit13.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1243_ (.D(Tile_X0Y1_FrameData[12]),
    .GATE(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit12.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1244_ (.D(Tile_X0Y1_FrameData[11]),
    .GATE(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit11.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1245_ (.D(Tile_X0Y1_FrameData[10]),
    .GATE(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit10.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1246_ (.D(Tile_X0Y1_FrameData[9]),
    .GATE(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit9.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1247_ (.D(Tile_X0Y1_FrameData[8]),
    .GATE(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit8.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1248_ (.D(Tile_X0Y1_FrameData[7]),
    .GATE(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit7.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1249_ (.D(Tile_X0Y1_FrameData[6]),
    .GATE(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit6.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1250_ (.D(Tile_X0Y1_FrameData[5]),
    .GATE(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit5.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1251_ (.D(Tile_X0Y1_FrameData[4]),
    .GATE(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit4.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1252_ (.D(Tile_X0Y1_FrameData[3]),
    .GATE(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit3.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1253_ (.D(Tile_X0Y1_FrameData[2]),
    .GATE(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit2.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1254_ (.D(Tile_X0Y1_FrameData[1]),
    .GATE(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit1.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1255_ (.D(Tile_X0Y1_FrameData[0]),
    .GATE(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit0.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1256_ (.D(Tile_X0Y1_FrameData[31]),
    .GATE(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit31.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1257_ (.D(Tile_X0Y1_FrameData[30]),
    .GATE(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit30.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1258_ (.D(Tile_X0Y1_FrameData[29]),
    .GATE(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit29.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1259_ (.D(Tile_X0Y1_FrameData[28]),
    .GATE(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit28.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1260_ (.D(Tile_X0Y1_FrameData[27]),
    .GATE(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit27.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1261_ (.D(Tile_X0Y1_FrameData[26]),
    .GATE(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit26.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1262_ (.D(Tile_X0Y1_FrameData[25]),
    .GATE(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit25.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1263_ (.D(Tile_X0Y1_FrameData[24]),
    .GATE(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit24.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1264_ (.D(Tile_X0Y1_FrameData[23]),
    .GATE(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit23.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1265_ (.D(Tile_X0Y1_FrameData[22]),
    .GATE(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit22.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1266_ (.D(Tile_X0Y1_FrameData[21]),
    .GATE(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit21.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1267_ (.D(Tile_X0Y1_FrameData[20]),
    .GATE(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit20.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1268_ (.D(Tile_X0Y1_FrameData[19]),
    .GATE(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit19.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1269_ (.D(Tile_X0Y1_FrameData[18]),
    .GATE(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit18.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1270_ (.D(Tile_X0Y1_FrameData[17]),
    .GATE(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit17.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1271_ (.D(Tile_X0Y1_FrameData[16]),
    .GATE(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit16.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1272_ (.D(Tile_X0Y1_FrameData[15]),
    .GATE(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit15.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1273_ (.D(Tile_X0Y1_FrameData[14]),
    .GATE(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit14.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1274_ (.D(Tile_X0Y1_FrameData[13]),
    .GATE(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit13.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1275_ (.D(Tile_X0Y1_FrameData[12]),
    .GATE(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit12.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1276_ (.D(Tile_X0Y1_FrameData[11]),
    .GATE(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit11.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1277_ (.D(Tile_X0Y1_FrameData[10]),
    .GATE(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit10.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1278_ (.D(Tile_X0Y1_FrameData[9]),
    .GATE(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit9.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1279_ (.D(Tile_X0Y1_FrameData[8]),
    .GATE(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit8.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1280_ (.D(Tile_X0Y1_FrameData[7]),
    .GATE(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit7.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1281_ (.D(Tile_X0Y1_FrameData[6]),
    .GATE(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit6.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1282_ (.D(Tile_X0Y1_FrameData[5]),
    .GATE(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit5.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1283_ (.D(Tile_X0Y1_FrameData[4]),
    .GATE(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit4.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1284_ (.D(Tile_X0Y1_FrameData[3]),
    .GATE(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit3.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1285_ (.D(Tile_X0Y1_FrameData[2]),
    .GATE(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit2.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1286_ (.D(Tile_X0Y1_FrameData[1]),
    .GATE(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit1.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1287_ (.D(Tile_X0Y1_FrameData[0]),
    .GATE(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit0.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1288_ (.D(Tile_X0Y1_FrameData[31]),
    .GATE(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit31.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1289_ (.D(Tile_X0Y1_FrameData[30]),
    .GATE(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit30.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1290_ (.D(Tile_X0Y1_FrameData[29]),
    .GATE(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit29.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1291_ (.D(Tile_X0Y1_FrameData[28]),
    .GATE(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit28.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1292_ (.D(Tile_X0Y1_FrameData[27]),
    .GATE(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit27.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1293_ (.D(Tile_X0Y1_FrameData[26]),
    .GATE(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit26.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1294_ (.D(Tile_X0Y1_FrameData[25]),
    .GATE(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit25.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1295_ (.D(Tile_X0Y1_FrameData[24]),
    .GATE(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit24.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1296_ (.D(Tile_X0Y1_FrameData[23]),
    .GATE(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit23.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1297_ (.D(Tile_X0Y1_FrameData[22]),
    .GATE(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit22.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1298_ (.D(Tile_X0Y1_FrameData[21]),
    .GATE(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit21.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1299_ (.D(Tile_X0Y1_FrameData[20]),
    .GATE(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit20.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1300_ (.D(Tile_X0Y1_FrameData[19]),
    .GATE(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit19.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1301_ (.D(Tile_X0Y1_FrameData[18]),
    .GATE(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit18.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1302_ (.D(Tile_X0Y1_FrameData[17]),
    .GATE(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit17.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1303_ (.D(Tile_X0Y1_FrameData[16]),
    .GATE(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit16.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1304_ (.D(Tile_X0Y1_FrameData[15]),
    .GATE(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit15.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1305_ (.D(Tile_X0Y1_FrameData[14]),
    .GATE(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit14.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1306_ (.D(Tile_X0Y1_FrameData[13]),
    .GATE(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit13.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1307_ (.D(Tile_X0Y1_FrameData[12]),
    .GATE(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit12.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1308_ (.D(Tile_X0Y1_FrameData[11]),
    .GATE(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit11.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1309_ (.D(Tile_X0Y1_FrameData[10]),
    .GATE(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit10.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1310_ (.D(Tile_X0Y1_FrameData[9]),
    .GATE(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit9.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1311_ (.D(Tile_X0Y1_FrameData[8]),
    .GATE(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit8.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1312_ (.D(Tile_X0Y1_FrameData[7]),
    .GATE(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit7.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1313_ (.D(Tile_X0Y1_FrameData[6]),
    .GATE(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit6.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1314_ (.D(Tile_X0Y1_FrameData[5]),
    .GATE(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit5.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1315_ (.D(Tile_X0Y1_FrameData[4]),
    .GATE(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit4.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1316_ (.D(Tile_X0Y1_FrameData[3]),
    .GATE(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit3.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1317_ (.D(Tile_X0Y1_FrameData[2]),
    .GATE(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit2.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1318_ (.D(Tile_X0Y1_FrameData[1]),
    .GATE(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit1.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1319_ (.D(Tile_X0Y1_FrameData[0]),
    .GATE(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit0.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1320_ (.D(Tile_X0Y1_FrameData[31]),
    .GATE(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit31.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1321_ (.D(Tile_X0Y1_FrameData[30]),
    .GATE(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit30.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1322_ (.D(Tile_X0Y1_FrameData[29]),
    .GATE(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit29.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1323_ (.D(Tile_X0Y1_FrameData[28]),
    .GATE(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit28.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1324_ (.D(Tile_X0Y1_FrameData[27]),
    .GATE(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit27.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1325_ (.D(Tile_X0Y1_FrameData[26]),
    .GATE(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit26.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1326_ (.D(Tile_X0Y1_FrameData[25]),
    .GATE(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit25.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1327_ (.D(Tile_X0Y1_FrameData[24]),
    .GATE(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit24.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1328_ (.D(Tile_X0Y1_FrameData[23]),
    .GATE(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit23.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1329_ (.D(Tile_X0Y1_FrameData[22]),
    .GATE(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit22.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1330_ (.D(Tile_X0Y1_FrameData[21]),
    .GATE(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit21.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1331_ (.D(Tile_X0Y1_FrameData[20]),
    .GATE(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit20.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1332_ (.D(Tile_X0Y1_FrameData[19]),
    .GATE(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit19.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1333_ (.D(Tile_X0Y1_FrameData[18]),
    .GATE(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit18.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1334_ (.D(Tile_X0Y1_FrameData[17]),
    .GATE(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit17.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1335_ (.D(Tile_X0Y1_FrameData[16]),
    .GATE(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit16.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1336_ (.D(Tile_X0Y1_FrameData[15]),
    .GATE(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit15.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1337_ (.D(Tile_X0Y1_FrameData[14]),
    .GATE(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit14.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1338_ (.D(Tile_X0Y1_FrameData[13]),
    .GATE(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit13.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1339_ (.D(Tile_X0Y1_FrameData[12]),
    .GATE(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit12.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1340_ (.D(Tile_X0Y1_FrameData[11]),
    .GATE(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit11.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1341_ (.D(Tile_X0Y1_FrameData[10]),
    .GATE(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit10.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1342_ (.D(Tile_X0Y1_FrameData[9]),
    .GATE(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit9.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1343_ (.D(Tile_X0Y1_FrameData[8]),
    .GATE(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit8.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1344_ (.D(Tile_X0Y1_FrameData[7]),
    .GATE(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit7.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1345_ (.D(Tile_X0Y1_FrameData[6]),
    .GATE(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit6.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1346_ (.D(Tile_X0Y1_FrameData[5]),
    .GATE(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit5.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1347_ (.D(Tile_X0Y1_FrameData[4]),
    .GATE(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit4.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1348_ (.D(Tile_X0Y1_FrameData[3]),
    .GATE(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit3.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1349_ (.D(Tile_X0Y1_FrameData[2]),
    .GATE(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit2.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1350_ (.D(Tile_X0Y1_FrameData[1]),
    .GATE(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit1.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1351_ (.D(Tile_X0Y1_FrameData[0]),
    .GATE(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit0.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1352_ (.D(Tile_X0Y1_FrameData[31]),
    .GATE(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit31.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1353_ (.D(Tile_X0Y1_FrameData[30]),
    .GATE(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit30.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1354_ (.D(Tile_X0Y1_FrameData[29]),
    .GATE(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit29.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1355_ (.D(Tile_X0Y1_FrameData[28]),
    .GATE(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit28.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1356_ (.D(Tile_X0Y1_FrameData[27]),
    .GATE(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit27.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1357_ (.D(Tile_X0Y1_FrameData[26]),
    .GATE(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit26.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1358_ (.D(Tile_X0Y1_FrameData[25]),
    .GATE(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit25.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1359_ (.D(Tile_X0Y1_FrameData[24]),
    .GATE(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit24.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1360_ (.D(Tile_X0Y1_FrameData[23]),
    .GATE(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit23.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1361_ (.D(Tile_X0Y1_FrameData[22]),
    .GATE(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit22.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1362_ (.D(Tile_X0Y1_FrameData[21]),
    .GATE(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit21.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1363_ (.D(Tile_X0Y1_FrameData[20]),
    .GATE(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit20.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1364_ (.D(Tile_X0Y1_FrameData[19]),
    .GATE(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit19.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1365_ (.D(Tile_X0Y1_FrameData[18]),
    .GATE(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit18.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1366_ (.D(Tile_X0Y1_FrameData[17]),
    .GATE(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit17.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1367_ (.D(Tile_X0Y1_FrameData[16]),
    .GATE(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit16.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1368_ (.D(Tile_X0Y1_FrameData[15]),
    .GATE(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit15.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1369_ (.D(Tile_X0Y1_FrameData[14]),
    .GATE(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit14.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1370_ (.D(Tile_X0Y1_FrameData[13]),
    .GATE(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit13.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1371_ (.D(Tile_X0Y1_FrameData[12]),
    .GATE(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit12.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1372_ (.D(Tile_X0Y1_FrameData[11]),
    .GATE(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit11.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1373_ (.D(Tile_X0Y1_FrameData[10]),
    .GATE(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit10.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1374_ (.D(Tile_X0Y1_FrameData[9]),
    .GATE(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit9.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1375_ (.D(Tile_X0Y1_FrameData[8]),
    .GATE(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit8.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1376_ (.D(Tile_X0Y1_FrameData[7]),
    .GATE(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit7.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1377_ (.D(Tile_X0Y1_FrameData[6]),
    .GATE(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit6.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1378_ (.D(Tile_X0Y1_FrameData[5]),
    .GATE(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit5.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1379_ (.D(Tile_X0Y1_FrameData[4]),
    .GATE(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit4.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1380_ (.D(Tile_X0Y1_FrameData[3]),
    .GATE(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit3.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1381_ (.D(Tile_X0Y1_FrameData[2]),
    .GATE(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit2.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1382_ (.D(Tile_X0Y1_FrameData[1]),
    .GATE(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit1.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1383_ (.D(Tile_X0Y1_FrameData[0]),
    .GATE(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit0.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1384_ (.D(Tile_X0Y1_FrameData[31]),
    .GATE(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit31.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1385_ (.D(Tile_X0Y1_FrameData[30]),
    .GATE(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit30.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1386_ (.D(Tile_X0Y1_FrameData[29]),
    .GATE(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit29.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1387_ (.D(Tile_X0Y1_FrameData[28]),
    .GATE(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit28.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1388_ (.D(Tile_X0Y1_FrameData[27]),
    .GATE(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit27.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1389_ (.D(Tile_X0Y1_FrameData[26]),
    .GATE(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit26.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1390_ (.D(Tile_X0Y1_FrameData[25]),
    .GATE(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit25.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1391_ (.D(Tile_X0Y1_FrameData[24]),
    .GATE(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit24.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1392_ (.D(Tile_X0Y1_FrameData[23]),
    .GATE(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit23.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1393_ (.D(Tile_X0Y1_FrameData[22]),
    .GATE(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit22.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1394_ (.D(Tile_X0Y1_FrameData[21]),
    .GATE(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit21.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1395_ (.D(Tile_X0Y1_FrameData[20]),
    .GATE(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit20.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1396_ (.D(Tile_X0Y1_FrameData[19]),
    .GATE(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit19.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1397_ (.D(Tile_X0Y1_FrameData[18]),
    .GATE(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit18.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1398_ (.D(Tile_X0Y1_FrameData[17]),
    .GATE(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit17.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1399_ (.D(Tile_X0Y1_FrameData[16]),
    .GATE(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit16.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1400_ (.D(Tile_X0Y1_FrameData[15]),
    .GATE(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit15.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1401_ (.D(Tile_X0Y1_FrameData[14]),
    .GATE(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit14.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1402_ (.D(Tile_X0Y1_FrameData[13]),
    .GATE(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit13.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1403_ (.D(Tile_X0Y1_FrameData[12]),
    .GATE(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit12.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1404_ (.D(Tile_X0Y1_FrameData[11]),
    .GATE(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit11.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1405_ (.D(Tile_X0Y1_FrameData[10]),
    .GATE(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit10.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1406_ (.D(Tile_X0Y1_FrameData[9]),
    .GATE(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit9.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1407_ (.D(Tile_X0Y1_FrameData[8]),
    .GATE(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit8.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1408_ (.D(Tile_X0Y1_FrameData[7]),
    .GATE(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit7.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1409_ (.D(Tile_X0Y1_FrameData[6]),
    .GATE(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit6.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1410_ (.D(Tile_X0Y1_FrameData[5]),
    .GATE(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit5.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1411_ (.D(Tile_X0Y1_FrameData[4]),
    .GATE(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit4.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1412_ (.D(Tile_X0Y1_FrameData[3]),
    .GATE(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit3.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1413_ (.D(Tile_X0Y1_FrameData[2]),
    .GATE(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit2.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1414_ (.D(Tile_X0Y1_FrameData[1]),
    .GATE(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit1.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _1415_ (.D(Tile_X0Y1_FrameData[0]),
    .GATE(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit0.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1416_ (.A(clknet_1_0__leaf_Tile_X0Y1_UserCLK),
    .X(CLK_TT_PROJECT),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1417_ (.A(Tile_X0Y0_FrameData[0]),
    .X(Tile_X0Y0_FrameData_O[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1418_ (.A(Tile_X0Y0_FrameData[1]),
    .X(Tile_X0Y0_FrameData_O[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1419_ (.A(Tile_X0Y0_FrameData[2]),
    .X(Tile_X0Y0_FrameData_O[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1420_ (.A(Tile_X0Y0_FrameData[3]),
    .X(Tile_X0Y0_FrameData_O[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1421_ (.A(Tile_X0Y0_FrameData[4]),
    .X(Tile_X0Y0_FrameData_O[4]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1422_ (.A(Tile_X0Y0_FrameData[5]),
    .X(Tile_X0Y0_FrameData_O[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1423_ (.A(Tile_X0Y0_FrameData[6]),
    .X(Tile_X0Y0_FrameData_O[6]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1424_ (.A(Tile_X0Y0_FrameData[7]),
    .X(Tile_X0Y0_FrameData_O[7]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1425_ (.A(Tile_X0Y0_FrameData[8]),
    .X(Tile_X0Y0_FrameData_O[8]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1426_ (.A(Tile_X0Y0_FrameData[9]),
    .X(Tile_X0Y0_FrameData_O[9]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1427_ (.A(Tile_X0Y0_FrameData[10]),
    .X(Tile_X0Y0_FrameData_O[10]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1428_ (.A(Tile_X0Y0_FrameData[11]),
    .X(Tile_X0Y0_FrameData_O[11]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1429_ (.A(Tile_X0Y0_FrameData[12]),
    .X(Tile_X0Y0_FrameData_O[12]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1430_ (.A(Tile_X0Y0_FrameData[13]),
    .X(Tile_X0Y0_FrameData_O[13]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1431_ (.A(Tile_X0Y0_FrameData[14]),
    .X(Tile_X0Y0_FrameData_O[14]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1432_ (.A(Tile_X0Y0_FrameData[15]),
    .X(Tile_X0Y0_FrameData_O[15]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1433_ (.A(Tile_X0Y0_FrameData[16]),
    .X(Tile_X0Y0_FrameData_O[16]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1434_ (.A(Tile_X0Y0_FrameData[17]),
    .X(Tile_X0Y0_FrameData_O[17]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1435_ (.A(Tile_X0Y0_FrameData[18]),
    .X(Tile_X0Y0_FrameData_O[18]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1436_ (.A(Tile_X0Y0_FrameData[19]),
    .X(Tile_X0Y0_FrameData_O[19]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1437_ (.A(Tile_X0Y0_FrameData[20]),
    .X(Tile_X0Y0_FrameData_O[20]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1438_ (.A(Tile_X0Y0_FrameData[21]),
    .X(Tile_X0Y0_FrameData_O[21]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1439_ (.A(Tile_X0Y0_FrameData[22]),
    .X(Tile_X0Y0_FrameData_O[22]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1440_ (.A(Tile_X0Y0_FrameData[23]),
    .X(Tile_X0Y0_FrameData_O[23]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1441_ (.A(Tile_X0Y0_FrameData[24]),
    .X(Tile_X0Y0_FrameData_O[24]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1442_ (.A(Tile_X0Y0_FrameData[25]),
    .X(Tile_X0Y0_FrameData_O[25]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1443_ (.A(Tile_X0Y0_FrameData[26]),
    .X(Tile_X0Y0_FrameData_O[26]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1444_ (.A(Tile_X0Y0_FrameData[27]),
    .X(Tile_X0Y0_FrameData_O[27]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1445_ (.A(Tile_X0Y0_FrameData[28]),
    .X(Tile_X0Y0_FrameData_O[28]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1446_ (.A(Tile_X0Y0_FrameData[29]),
    .X(Tile_X0Y0_FrameData_O[29]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1447_ (.A(Tile_X0Y0_FrameData[30]),
    .X(Tile_X0Y0_FrameData_O[30]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1448_ (.A(Tile_X0Y0_FrameData[31]),
    .X(Tile_X0Y0_FrameData_O[31]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1449_ (.A(Tile_X0Y1_FrameStrobe[0]),
    .X(Tile_X0Y0_FrameStrobe_O[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1450_ (.A(Tile_X0Y1_FrameStrobe[1]),
    .X(Tile_X0Y0_FrameStrobe_O[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1451_ (.A(Tile_X0Y1_FrameStrobe[2]),
    .X(Tile_X0Y0_FrameStrobe_O[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1452_ (.A(Tile_X0Y1_FrameStrobe[3]),
    .X(Tile_X0Y0_FrameStrobe_O[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1453_ (.A(Tile_X0Y1_FrameStrobe[4]),
    .X(Tile_X0Y0_FrameStrobe_O[4]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1454_ (.A(Tile_X0Y1_FrameStrobe[5]),
    .X(Tile_X0Y0_FrameStrobe_O[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1455_ (.A(Tile_X0Y1_FrameStrobe[6]),
    .X(Tile_X0Y0_FrameStrobe_O[6]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1456_ (.A(Tile_X0Y1_FrameStrobe[7]),
    .X(Tile_X0Y0_FrameStrobe_O[7]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1457_ (.A(Tile_X0Y1_FrameStrobe[8]),
    .X(Tile_X0Y0_FrameStrobe_O[8]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1458_ (.A(Tile_X0Y1_FrameStrobe[9]),
    .X(Tile_X0Y0_FrameStrobe_O[9]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1459_ (.A(Tile_X0Y1_FrameStrobe[10]),
    .X(Tile_X0Y0_FrameStrobe_O[10]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1460_ (.A(Tile_X0Y1_FrameStrobe[11]),
    .X(Tile_X0Y0_FrameStrobe_O[11]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1461_ (.A(Tile_X0Y1_FrameStrobe[12]),
    .X(Tile_X0Y0_FrameStrobe_O[12]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1462_ (.A(Tile_X0Y1_FrameStrobe[13]),
    .X(Tile_X0Y0_FrameStrobe_O[13]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1463_ (.A(Tile_X0Y1_FrameStrobe[14]),
    .X(Tile_X0Y0_FrameStrobe_O[14]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1464_ (.A(Tile_X0Y1_FrameStrobe[15]),
    .X(Tile_X0Y0_FrameStrobe_O[15]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1465_ (.A(Tile_X0Y1_FrameStrobe[16]),
    .X(Tile_X0Y0_FrameStrobe_O[16]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1466_ (.A(Tile_X0Y1_FrameStrobe[17]),
    .X(Tile_X0Y0_FrameStrobe_O[17]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1467_ (.A(Tile_X0Y1_FrameStrobe[18]),
    .X(Tile_X0Y0_FrameStrobe_O[18]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1468_ (.A(Tile_X0Y1_FrameStrobe[19]),
    .X(Tile_X0Y0_FrameStrobe_O[19]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1469_ (.A(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N1BEG0 ),
    .X(Tile_X0Y0_N1BEG[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1470_ (.A(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N1BEG1 ),
    .X(Tile_X0Y0_N1BEG[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1471_ (.A(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N1BEG2 ),
    .X(Tile_X0Y0_N1BEG[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1472_ (.A(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N1BEG3 ),
    .X(Tile_X0Y0_N1BEG[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1473_ (.A(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N2BEG0 ),
    .X(Tile_X0Y0_N2BEG[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1474_ (.A(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N2BEG1 ),
    .X(Tile_X0Y0_N2BEG[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1475_ (.A(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N2BEG2 ),
    .X(Tile_X0Y0_N2BEG[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1476_ (.A(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N2BEG3 ),
    .X(Tile_X0Y0_N2BEG[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1477_ (.A(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N2BEG4 ),
    .X(Tile_X0Y0_N2BEG[4]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1478_ (.A(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N2BEG5 ),
    .X(Tile_X0Y0_N2BEG[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1479_ (.A(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N2BEG6 ),
    .X(Tile_X0Y0_N2BEG[6]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1480_ (.A(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N2BEG7 ),
    .X(Tile_X0Y0_N2BEG[7]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1481_ (.A(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N2BEGb0 ),
    .X(Tile_X0Y0_N2BEGb[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1482_ (.A(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N2BEGb1 ),
    .X(Tile_X0Y0_N2BEGb[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1483_ (.A(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N2BEGb2 ),
    .X(Tile_X0Y0_N2BEGb[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1484_ (.A(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N2BEGb3 ),
    .X(Tile_X0Y0_N2BEGb[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1485_ (.A(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N2BEGb4 ),
    .X(Tile_X0Y0_N2BEGb[4]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1486_ (.A(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N2BEGb5 ),
    .X(Tile_X0Y0_N2BEGb[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1487_ (.A(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N2BEGb6 ),
    .X(Tile_X0Y0_N2BEGb[6]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1488_ (.A(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N2BEGb7 ),
    .X(Tile_X0Y0_N2BEGb[7]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1489_ (.A(Tile_X0Y1_N4END[8]),
    .X(Tile_X0Y0_N4BEG[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1490_ (.A(Tile_X0Y1_N4END[9]),
    .X(Tile_X0Y0_N4BEG[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1491_ (.A(Tile_X0Y1_N4END[10]),
    .X(Tile_X0Y0_N4BEG[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1492_ (.A(Tile_X0Y1_N4END[11]),
    .X(Tile_X0Y0_N4BEG[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1493_ (.A(Tile_X0Y1_N4END[12]),
    .X(Tile_X0Y0_N4BEG[4]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1494_ (.A(Tile_X0Y1_N4END[13]),
    .X(Tile_X0Y0_N4BEG[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1495_ (.A(Tile_X0Y1_N4END[14]),
    .X(Tile_X0Y0_N4BEG[6]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1496_ (.A(Tile_X0Y1_N4END[15]),
    .X(Tile_X0Y0_N4BEG[7]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1497_ (.A(\Tile_X0Y0_E_TT_IF2_top.N4BEG_outbuf_8.A ),
    .X(Tile_X0Y0_N4BEG[8]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1498_ (.A(\Tile_X0Y0_E_TT_IF2_top.N4BEG_outbuf_9.A ),
    .X(Tile_X0Y0_N4BEG[9]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1499_ (.A(\Tile_X0Y0_E_TT_IF2_top.N4BEG_outbuf_10.A ),
    .X(Tile_X0Y0_N4BEG[10]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1500_ (.A(\Tile_X0Y0_E_TT_IF2_top.N4BEG_outbuf_11.A ),
    .X(Tile_X0Y0_N4BEG[11]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1501_ (.A(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N4BEG0 ),
    .X(Tile_X0Y0_N4BEG[12]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1502_ (.A(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N4BEG1 ),
    .X(Tile_X0Y0_N4BEG[13]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1503_ (.A(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N4BEG2 ),
    .X(Tile_X0Y0_N4BEG[14]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1504_ (.A(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N4BEG3 ),
    .X(Tile_X0Y0_N4BEG[15]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1505_ (.A(clknet_1_1__leaf_Tile_X0Y1_UserCLK),
    .X(Tile_X0Y0_UserCLKo),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1506_ (.A(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W1BEG0 ),
    .X(Tile_X0Y0_W1BEG[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1507_ (.A(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W1BEG1 ),
    .X(Tile_X0Y0_W1BEG[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1508_ (.A(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W1BEG2 ),
    .X(Tile_X0Y0_W1BEG[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1509_ (.A(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W1BEG3 ),
    .X(Tile_X0Y0_W1BEG[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1510_ (.A(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W2BEG0 ),
    .X(Tile_X0Y0_W2BEG[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1511_ (.A(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W2BEG1 ),
    .X(Tile_X0Y0_W2BEG[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1512_ (.A(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W2BEG2 ),
    .X(Tile_X0Y0_W2BEG[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1513_ (.A(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W2BEG3 ),
    .X(Tile_X0Y0_W2BEG[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1514_ (.A(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W2BEG4 ),
    .X(Tile_X0Y0_W2BEG[4]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1515_ (.A(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W2BEG5 ),
    .X(Tile_X0Y0_W2BEG[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1516_ (.A(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W2BEG6 ),
    .X(Tile_X0Y0_W2BEG[6]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1517_ (.A(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W2BEG7 ),
    .X(Tile_X0Y0_W2BEG[7]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1518_ (.A(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W2BEGb0 ),
    .X(Tile_X0Y0_W2BEGb[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1519_ (.A(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W2BEGb1 ),
    .X(Tile_X0Y0_W2BEGb[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1520_ (.A(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W2BEGb2 ),
    .X(Tile_X0Y0_W2BEGb[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1521_ (.A(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W2BEGb3 ),
    .X(Tile_X0Y0_W2BEGb[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1522_ (.A(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W2BEGb4 ),
    .X(Tile_X0Y0_W2BEGb[4]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1523_ (.A(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W2BEGb5 ),
    .X(Tile_X0Y0_W2BEGb[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1524_ (.A(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W2BEGb6 ),
    .X(Tile_X0Y0_W2BEGb[6]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1525_ (.A(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W2BEGb7 ),
    .X(Tile_X0Y0_W2BEGb[7]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1526_ (.A(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W6BEG0 ),
    .X(Tile_X0Y0_W6BEG[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1527_ (.A(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W6BEG1 ),
    .X(Tile_X0Y0_W6BEG[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1528_ (.A(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W6BEG2 ),
    .X(Tile_X0Y0_W6BEG[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1529_ (.A(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W6BEG3 ),
    .X(Tile_X0Y0_W6BEG[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1530_ (.A(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W6BEG4 ),
    .X(Tile_X0Y0_W6BEG[4]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1531_ (.A(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W6BEG5 ),
    .X(Tile_X0Y0_W6BEG[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1532_ (.A(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W6BEG6 ),
    .X(Tile_X0Y0_W6BEG[6]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1533_ (.A(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W6BEG7 ),
    .X(Tile_X0Y0_W6BEG[7]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1534_ (.A(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W6BEG8 ),
    .X(Tile_X0Y0_W6BEG[8]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1535_ (.A(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W6BEG9 ),
    .X(Tile_X0Y0_W6BEG[9]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1536_ (.A(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W6BEG10 ),
    .X(Tile_X0Y0_W6BEG[10]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1537_ (.A(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W6BEG11 ),
    .X(Tile_X0Y0_W6BEG[11]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1538_ (.A(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.WW4BEG0 ),
    .X(Tile_X0Y0_WW4BEG[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1539_ (.A(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.WW4BEG1 ),
    .X(Tile_X0Y0_WW4BEG[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1540_ (.A(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.WW4BEG2 ),
    .X(Tile_X0Y0_WW4BEG[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1541_ (.A(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.WW4BEG3 ),
    .X(Tile_X0Y0_WW4BEG[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1542_ (.A(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.WW4BEG4 ),
    .X(Tile_X0Y0_WW4BEG[4]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1543_ (.A(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.WW4BEG5 ),
    .X(Tile_X0Y0_WW4BEG[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1544_ (.A(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.WW4BEG6 ),
    .X(Tile_X0Y0_WW4BEG[6]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1545_ (.A(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.WW4BEG7 ),
    .X(Tile_X0Y0_WW4BEG[7]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1546_ (.A(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.WW4BEG8 ),
    .X(Tile_X0Y0_WW4BEG[8]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1547_ (.A(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.WW4BEG9 ),
    .X(Tile_X0Y0_WW4BEG[9]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1548_ (.A(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.WW4BEG10 ),
    .X(Tile_X0Y0_WW4BEG[10]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1549_ (.A(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.WW4BEG11 ),
    .X(Tile_X0Y0_WW4BEG[11]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1550_ (.A(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.WW4BEG12 ),
    .X(Tile_X0Y0_WW4BEG[12]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1551_ (.A(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.WW4BEG13 ),
    .X(Tile_X0Y0_WW4BEG[13]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1552_ (.A(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.WW4BEG14 ),
    .X(Tile_X0Y0_WW4BEG[14]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1553_ (.A(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.WW4BEG15 ),
    .X(Tile_X0Y0_WW4BEG[15]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1554_ (.A(Tile_X0Y1_FrameData[0]),
    .X(Tile_X0Y1_FrameData_O[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1555_ (.A(Tile_X0Y1_FrameData[1]),
    .X(Tile_X0Y1_FrameData_O[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1556_ (.A(Tile_X0Y1_FrameData[2]),
    .X(Tile_X0Y1_FrameData_O[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1557_ (.A(Tile_X0Y1_FrameData[3]),
    .X(Tile_X0Y1_FrameData_O[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1558_ (.A(Tile_X0Y1_FrameData[4]),
    .X(Tile_X0Y1_FrameData_O[4]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1559_ (.A(Tile_X0Y1_FrameData[5]),
    .X(Tile_X0Y1_FrameData_O[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1560_ (.A(Tile_X0Y1_FrameData[6]),
    .X(Tile_X0Y1_FrameData_O[6]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1561_ (.A(Tile_X0Y1_FrameData[7]),
    .X(Tile_X0Y1_FrameData_O[7]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1562_ (.A(Tile_X0Y1_FrameData[8]),
    .X(Tile_X0Y1_FrameData_O[8]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1563_ (.A(Tile_X0Y1_FrameData[9]),
    .X(Tile_X0Y1_FrameData_O[9]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1564_ (.A(Tile_X0Y1_FrameData[10]),
    .X(Tile_X0Y1_FrameData_O[10]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1565_ (.A(Tile_X0Y1_FrameData[11]),
    .X(Tile_X0Y1_FrameData_O[11]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1566_ (.A(Tile_X0Y1_FrameData[12]),
    .X(Tile_X0Y1_FrameData_O[12]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1567_ (.A(Tile_X0Y1_FrameData[13]),
    .X(Tile_X0Y1_FrameData_O[13]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1568_ (.A(Tile_X0Y1_FrameData[14]),
    .X(Tile_X0Y1_FrameData_O[14]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1569_ (.A(Tile_X0Y1_FrameData[15]),
    .X(Tile_X0Y1_FrameData_O[15]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1570_ (.A(Tile_X0Y1_FrameData[16]),
    .X(Tile_X0Y1_FrameData_O[16]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1571_ (.A(Tile_X0Y1_FrameData[17]),
    .X(Tile_X0Y1_FrameData_O[17]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1572_ (.A(Tile_X0Y1_FrameData[18]),
    .X(Tile_X0Y1_FrameData_O[18]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1573_ (.A(Tile_X0Y1_FrameData[19]),
    .X(Tile_X0Y1_FrameData_O[19]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1574_ (.A(Tile_X0Y1_FrameData[20]),
    .X(Tile_X0Y1_FrameData_O[20]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1575_ (.A(Tile_X0Y1_FrameData[21]),
    .X(Tile_X0Y1_FrameData_O[21]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1576_ (.A(Tile_X0Y1_FrameData[22]),
    .X(Tile_X0Y1_FrameData_O[22]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1577_ (.A(Tile_X0Y1_FrameData[23]),
    .X(Tile_X0Y1_FrameData_O[23]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1578_ (.A(Tile_X0Y1_FrameData[24]),
    .X(Tile_X0Y1_FrameData_O[24]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1579_ (.A(Tile_X0Y1_FrameData[25]),
    .X(Tile_X0Y1_FrameData_O[25]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1580_ (.A(Tile_X0Y1_FrameData[26]),
    .X(Tile_X0Y1_FrameData_O[26]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1581_ (.A(Tile_X0Y1_FrameData[27]),
    .X(Tile_X0Y1_FrameData_O[27]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1582_ (.A(Tile_X0Y1_FrameData[28]),
    .X(Tile_X0Y1_FrameData_O[28]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1583_ (.A(Tile_X0Y1_FrameData[29]),
    .X(Tile_X0Y1_FrameData_O[29]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1584_ (.A(Tile_X0Y1_FrameData[30]),
    .X(Tile_X0Y1_FrameData_O[30]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1585_ (.A(Tile_X0Y1_FrameData[31]),
    .X(Tile_X0Y1_FrameData_O[31]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1586_ (.A(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.S1BEG0 ),
    .X(Tile_X0Y1_S1BEG[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1587_ (.A(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.S1BEG1 ),
    .X(Tile_X0Y1_S1BEG[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1588_ (.A(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.S1BEG2 ),
    .X(Tile_X0Y1_S1BEG[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1589_ (.A(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.S1BEG3 ),
    .X(Tile_X0Y1_S1BEG[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1590_ (.A(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.S2BEG0 ),
    .X(Tile_X0Y1_S2BEG[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1591_ (.A(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.S2BEG1 ),
    .X(Tile_X0Y1_S2BEG[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1592_ (.A(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.S2BEG2 ),
    .X(Tile_X0Y1_S2BEG[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1593_ (.A(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.S2BEG3 ),
    .X(Tile_X0Y1_S2BEG[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1594_ (.A(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.S2BEG4 ),
    .X(Tile_X0Y1_S2BEG[4]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1595_ (.A(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.S2BEG5 ),
    .X(Tile_X0Y1_S2BEG[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1596_ (.A(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.S2BEG6 ),
    .X(Tile_X0Y1_S2BEG[6]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1597_ (.A(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.S2BEG7 ),
    .X(Tile_X0Y1_S2BEG[7]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1598_ (.A(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.S2BEG0 ),
    .X(Tile_X0Y1_S2BEGb[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1599_ (.A(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.S2BEG1 ),
    .X(Tile_X0Y1_S2BEGb[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1600_ (.A(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.S2BEG2 ),
    .X(Tile_X0Y1_S2BEGb[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1601_ (.A(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.S2BEG3 ),
    .X(Tile_X0Y1_S2BEGb[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1602_ (.A(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.S2BEG4 ),
    .X(Tile_X0Y1_S2BEGb[4]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1603_ (.A(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.S2BEG5 ),
    .X(Tile_X0Y1_S2BEGb[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1604_ (.A(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.S2BEG6 ),
    .X(Tile_X0Y1_S2BEGb[6]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1605_ (.A(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.S2BEG7 ),
    .X(Tile_X0Y1_S2BEGb[7]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1606_ (.A(Tile_X0Y0_S4END[8]),
    .X(Tile_X0Y1_S4BEG[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1607_ (.A(Tile_X0Y0_S4END[9]),
    .X(Tile_X0Y1_S4BEG[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1608_ (.A(Tile_X0Y0_S4END[10]),
    .X(Tile_X0Y1_S4BEG[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1609_ (.A(Tile_X0Y0_S4END[11]),
    .X(Tile_X0Y1_S4BEG[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1610_ (.A(Tile_X0Y0_S4END[12]),
    .X(Tile_X0Y1_S4BEG[4]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1611_ (.A(Tile_X0Y0_S4END[13]),
    .X(Tile_X0Y1_S4BEG[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1612_ (.A(Tile_X0Y0_S4END[14]),
    .X(Tile_X0Y1_S4BEG[6]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1613_ (.A(Tile_X0Y0_S4END[15]),
    .X(Tile_X0Y1_S4BEG[7]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1614_ (.A(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.S4BEG0 ),
    .X(Tile_X0Y1_S4BEG[8]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1615_ (.A(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.S4BEG1 ),
    .X(Tile_X0Y1_S4BEG[9]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1616_ (.A(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.S4BEG2 ),
    .X(Tile_X0Y1_S4BEG[10]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1617_ (.A(\Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.S4BEG3 ),
    .X(Tile_X0Y1_S4BEG[11]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1618_ (.A(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.S4BEG0 ),
    .X(Tile_X0Y1_S4BEG[12]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1619_ (.A(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.S4BEG1 ),
    .X(Tile_X0Y1_S4BEG[13]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1620_ (.A(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.S4BEG2 ),
    .X(Tile_X0Y1_S4BEG[14]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1621_ (.A(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.S4BEG3 ),
    .X(Tile_X0Y1_S4BEG[15]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1622_ (.A(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W1BEG0 ),
    .X(Tile_X0Y1_W1BEG[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1623_ (.A(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W1BEG1 ),
    .X(Tile_X0Y1_W1BEG[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1624_ (.A(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W1BEG2 ),
    .X(Tile_X0Y1_W1BEG[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1625_ (.A(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W1BEG3 ),
    .X(Tile_X0Y1_W1BEG[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1626_ (.A(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W2BEG0 ),
    .X(Tile_X0Y1_W2BEG[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1627_ (.A(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W2BEG1 ),
    .X(Tile_X0Y1_W2BEG[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1628_ (.A(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W2BEG2 ),
    .X(Tile_X0Y1_W2BEG[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1629_ (.A(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W2BEG3 ),
    .X(Tile_X0Y1_W2BEG[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1630_ (.A(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W2BEG4 ),
    .X(Tile_X0Y1_W2BEG[4]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1631_ (.A(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W2BEG5 ),
    .X(Tile_X0Y1_W2BEG[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1632_ (.A(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W2BEG6 ),
    .X(Tile_X0Y1_W2BEG[6]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1633_ (.A(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W2BEG7 ),
    .X(Tile_X0Y1_W2BEG[7]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1634_ (.A(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W2BEGb0 ),
    .X(Tile_X0Y1_W2BEGb[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1635_ (.A(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W2BEGb1 ),
    .X(Tile_X0Y1_W2BEGb[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1636_ (.A(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W2BEGb2 ),
    .X(Tile_X0Y1_W2BEGb[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1637_ (.A(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W2BEGb3 ),
    .X(Tile_X0Y1_W2BEGb[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1638_ (.A(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W2BEGb4 ),
    .X(Tile_X0Y1_W2BEGb[4]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1639_ (.A(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W2BEGb5 ),
    .X(Tile_X0Y1_W2BEGb[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1640_ (.A(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W2BEGb6 ),
    .X(Tile_X0Y1_W2BEGb[6]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1641_ (.A(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W2BEGb7 ),
    .X(Tile_X0Y1_W2BEGb[7]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1642_ (.A(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W6BEG0 ),
    .X(Tile_X0Y1_W6BEG[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1643_ (.A(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W6BEG1 ),
    .X(Tile_X0Y1_W6BEG[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1644_ (.A(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W6BEG2 ),
    .X(Tile_X0Y1_W6BEG[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1645_ (.A(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W6BEG3 ),
    .X(Tile_X0Y1_W6BEG[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1646_ (.A(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W6BEG4 ),
    .X(Tile_X0Y1_W6BEG[4]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1647_ (.A(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W6BEG5 ),
    .X(Tile_X0Y1_W6BEG[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1648_ (.A(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W6BEG6 ),
    .X(Tile_X0Y1_W6BEG[6]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1649_ (.A(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W6BEG7 ),
    .X(Tile_X0Y1_W6BEG[7]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1650_ (.A(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W6BEG8 ),
    .X(Tile_X0Y1_W6BEG[8]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1651_ (.A(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W6BEG9 ),
    .X(Tile_X0Y1_W6BEG[9]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1652_ (.A(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W6BEG10 ),
    .X(Tile_X0Y1_W6BEG[10]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1653_ (.A(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W6BEG11 ),
    .X(Tile_X0Y1_W6BEG[11]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1654_ (.A(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.WW4BEG0 ),
    .X(Tile_X0Y1_WW4BEG[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1655_ (.A(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.WW4BEG1 ),
    .X(Tile_X0Y1_WW4BEG[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1656_ (.A(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.WW4BEG2 ),
    .X(Tile_X0Y1_WW4BEG[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1657_ (.A(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.WW4BEG3 ),
    .X(Tile_X0Y1_WW4BEG[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1658_ (.A(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.WW4BEG4 ),
    .X(Tile_X0Y1_WW4BEG[4]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1659_ (.A(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.WW4BEG5 ),
    .X(Tile_X0Y1_WW4BEG[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1660_ (.A(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.WW4BEG6 ),
    .X(Tile_X0Y1_WW4BEG[6]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1661_ (.A(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.WW4BEG7 ),
    .X(Tile_X0Y1_WW4BEG[7]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1662_ (.A(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.WW4BEG8 ),
    .X(Tile_X0Y1_WW4BEG[8]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1663_ (.A(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.WW4BEG9 ),
    .X(Tile_X0Y1_WW4BEG[9]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1664_ (.A(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.WW4BEG10 ),
    .X(Tile_X0Y1_WW4BEG[10]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1665_ (.A(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.WW4BEG11 ),
    .X(Tile_X0Y1_WW4BEG[11]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1666_ (.A(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.WW4BEG12 ),
    .X(Tile_X0Y1_WW4BEG[12]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1667_ (.A(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.WW4BEG13 ),
    .X(Tile_X0Y1_WW4BEG[13]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1668_ (.A(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.WW4BEG14 ),
    .X(Tile_X0Y1_WW4BEG[14]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _1669_ (.A(\Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.WW4BEG15 ),
    .X(Tile_X0Y1_WW4BEG[15]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_0_Tile_X0Y1_UserCLK (.A(Tile_X0Y1_UserCLK),
    .X(clknet_0_Tile_X0Y1_UserCLK),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_1_0__f_Tile_X0Y1_UserCLK (.A(clknet_0_Tile_X0Y1_UserCLK),
    .X(clknet_1_0__leaf_Tile_X0Y1_UserCLK),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_1_1__f_Tile_X0Y1_UserCLK (.A(clknet_0_Tile_X0Y1_UserCLK),
    .X(clknet_1_1__leaf_Tile_X0Y1_UserCLK),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_antennanp ANTENNA_1 (.VDD(VPWR),
    .VSS(VGND),
    .A(Tile_X0Y0_S2END[4]));
 sg13g2_antennanp ANTENNA_2 (.VDD(VPWR),
    .VSS(VGND),
    .A(Tile_X0Y1_FrameStrobe[10]));
 sg13g2_antennanp ANTENNA_3 (.VDD(VPWR),
    .VSS(VGND),
    .A(Tile_X0Y1_FrameStrobe[11]));
 sg13g2_antennanp ANTENNA_4 (.VDD(VPWR),
    .VSS(VGND),
    .A(Tile_X0Y1_FrameStrobe[12]));
 sg13g2_antennanp ANTENNA_5 (.VDD(VPWR),
    .VSS(VGND),
    .A(Tile_X0Y1_FrameStrobe[13]));
 sg13g2_antennanp ANTENNA_6 (.VDD(VPWR),
    .VSS(VGND),
    .A(Tile_X0Y1_FrameStrobe[14]));
 sg13g2_antennanp ANTENNA_7 (.VDD(VPWR),
    .VSS(VGND),
    .A(Tile_X0Y1_FrameStrobe[15]));
 sg13g2_antennanp ANTENNA_8 (.VDD(VPWR),
    .VSS(VGND),
    .A(Tile_X0Y1_FrameStrobe[16]));
 sg13g2_antennanp ANTENNA_9 (.VDD(VPWR),
    .VSS(VGND),
    .A(Tile_X0Y1_FrameStrobe[17]));
 sg13g2_antennanp ANTENNA_10 (.VDD(VPWR),
    .VSS(VGND),
    .A(Tile_X0Y1_FrameStrobe[18]));
 sg13g2_antennanp ANTENNA_11 (.VDD(VPWR),
    .VSS(VGND),
    .A(Tile_X0Y1_FrameStrobe[8]));
 sg13g2_antennanp ANTENNA_12 (.VDD(VPWR),
    .VSS(VGND),
    .A(Tile_X0Y1_FrameStrobe[9]));
 sg13g2_antennanp ANTENNA_13 (.VDD(VPWR),
    .VSS(VGND),
    .A(Tile_X0Y1_N2MID[5]));
 sg13g2_antennanp ANTENNA_14 (.VDD(VPWR),
    .VSS(VGND),
    .A(Tile_X0Y1_N2MID[5]));
 sg13g2_antennanp ANTENNA_15 (.VDD(VPWR),
    .VSS(VGND),
    .A(Tile_X0Y1_N2MID[5]));
 sg13g2_antennanp ANTENNA_16 (.VDD(VPWR),
    .VSS(VGND),
    .A(Tile_X0Y1_N2MID[5]));
 sg13g2_antennanp ANTENNA_17 (.VDD(VPWR),
    .VSS(VGND),
    .A(Tile_X0Y1_FrameStrobe[19]));
 sg13g2_fill_2 FILLER_0_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_2 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_15 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_22 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_29 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_0_36 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_40 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_48 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_61 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_72 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_79 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_142 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_0_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_156 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_163 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_170 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_177 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_184 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_191 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_198 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_2 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_19 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_51 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_117 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_124 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_129 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_131 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_160 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_167 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_174 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_181 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_188 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_1_195 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_2 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_16 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_23 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_2_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_107 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_114 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_121 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_139 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_141 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_159 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_166 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_173 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_180 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_187 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_2_194 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_198 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_2 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_23 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_3_50 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_76 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_141 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_2 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_15 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_22 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_24 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_44 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_50 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_57 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_72 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_79 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_86 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_92 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_4_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_120 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_160 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_167 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_174 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_181 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_188 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_4_195 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_45 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_72 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_97 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_5_125 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_129 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_148 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_166 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_173 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_180 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_187 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_5_194 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_198 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_19 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_75 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_6_101 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_6_139 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_143 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_22 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_24 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_138 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_145 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_183 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_190 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_197 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_2 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_80 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_82 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_100 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_141 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_185 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_192 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_2 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_10_68 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_72 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_120 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_127 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_134 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_152 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_159 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_166 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_10_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_2 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_15 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_11_26 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_43 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_50 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_52 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_92 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_94 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_11_146 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_150 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_169 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_171 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_11_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_12_78 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_12_120 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_145 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_184 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_191 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_198 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_13_26 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_30 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_13_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_100 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_107 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_13_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_14_69 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_94 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_96 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_101 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_103 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_121 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_190 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_197 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_15_30 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_34 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_15_124 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_128 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_55 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_57 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_79 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_86 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_106 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_113 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_16_120 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_124 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_146 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_170 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_177 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_184 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_191 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_198 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_48 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_55 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_62 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_83 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_17_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_17_128 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_170 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_17_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_50 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_57 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_64 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_66 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_18_106 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_148 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_155 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_162 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_185 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_192 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_80 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_87 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_19_94 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_153 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_177 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_184 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_191 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_198 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_20_26 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_68 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_75 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_82 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_104 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_20_111 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_115 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_20_134 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_181 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_188 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_20_195 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_43 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_122 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_184 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_191 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_198 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_44 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_97 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_104 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_106 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_22_124 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_22_167 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_188 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_22_195 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_22 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_29 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_31 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_122 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_129 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_156 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_184 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_191 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_198 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_24_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_29 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_69 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_97 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_24_121 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_125 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_148 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_155 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_162 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_25_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_30 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_149 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_177 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_184 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_191 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_198 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_26_83 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_104 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_26_111 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_26_132 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_136 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_184 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_191 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_198 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_27_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_22 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_45 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_104 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_27_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_148 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_187 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_27_194 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_198 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_28_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_76 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_83 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_90 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_97 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_28_104 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_128 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_163 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_167 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_174 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_181 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_188 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_28_195 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_45 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_83 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_90 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_132 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_160 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_184 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_197 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_17 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_30_103 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_148 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_173 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_198 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_37 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_55 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_121 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_31_141 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_145 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_31_169 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_173 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_192 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_9 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_32_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_106 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_113 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_32_120 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_141 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_159 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_170 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_177 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_184 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_191 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_198 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_2 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_33_20 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_33_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_50 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_33_106 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_110 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_33_129 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_89 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_107 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_34_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_134 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_157 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_164 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_166 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_198 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_48 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_66 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_73 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_75 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_35_97 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_35_118 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_122 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_149 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_35_170 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_174 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_198 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_17 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_19 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_68 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_33 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_40 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_79 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_108 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_131 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_155 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_174 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_17 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_52 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_59 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_78 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_80 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_118 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_124 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_157 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_164 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_39_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_50 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_39_57 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_111 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_127 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_39_155 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_176 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_198 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_30 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_54 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_40_76 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_80 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_198 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_41_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_68 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_80 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_41_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_41_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_164 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_171 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_178 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_185 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_192 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_78 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_85 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_92 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_99 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_106 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_113 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_42_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_42_150 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_173 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_180 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_187 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_42_194 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_198 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_43_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_22 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_29 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_48 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_43_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_113 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_115 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_157 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_164 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_171 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_178 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_185 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_192 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_44_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_156 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_163 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_170 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_177 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_44_184 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_188 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_44_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_33 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_51 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_93 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_120 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_132 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_162 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_169 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_176 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_183 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_104 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_184 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_197 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_47_43 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_47 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_82 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_47_89 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_93 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_139 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_146 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_153 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_160 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_167 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_174 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_47_181 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_48_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_48_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_48_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_128 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_146 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_153 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_160 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_167 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_174 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_48_181 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_48_197 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_49_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_49_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_64 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_49_73 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_96 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_49_103 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_49_141 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_49_145 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_49_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_49_185 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_50_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_97 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_50_104 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_50_106 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_129 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_50_136 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_142 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_149 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_156 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_163 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_170 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_177 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_50_184 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_50_188 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_51_62 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_51_66 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_87 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_51_94 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_51_113 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_51_117 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_124 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_131 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_138 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_145 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_152 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_159 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_166 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_173 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_51_180 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_51_184 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_51_197 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_51_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_17 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_52_24 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_52_45 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_52_83 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_52_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_127 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_134 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_141 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_148 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_155 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_162 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_169 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_176 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_52_183 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_53_24 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_53_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_87 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_53_94 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_53_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_124 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_131 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_138 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_145 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_152 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_159 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_166 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_173 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_53_180 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_53_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_54_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_54_36 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_54_41 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_59 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_117 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_124 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_131 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_138 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_145 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_152 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_54_159 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_54_163 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_54_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_54_177 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_54_198 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_55_17 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_59 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_55_66 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_55_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_89 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_96 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_103 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_55_110 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_55_114 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_55_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_55_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_55_197 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_55_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_56_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_56_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_34 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_41 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_56_48 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_56_90 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_56_129 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_56_131 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_56_136 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_56_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_56_146 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_56_150 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_177 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_56_184 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_57_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_57_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_65 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_72 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_57_79 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_57_85 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_57_87 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_57_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_57_132 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_57_171 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_57_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_57_197 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_57_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_58_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_58_2 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_58_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_33 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_58_40 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_58_44 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_58_66 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_104 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_58_111 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_134 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_58_141 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_58_145 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_58_167 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_58_171 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_58_198 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_59_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_59_2 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_59_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_59_47 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_59_51 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_59_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_110 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_59_117 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_59_121 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_59_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_59_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_59_195 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_59_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_17 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_24 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_60_31 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_60_33 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_60_68 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_60_110 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_60_115 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_138 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_60_145 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_163 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_60_170 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_60_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_60_198 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_61_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_61_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_31 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_59 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_61_66 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_61_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_61_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_61_97 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_61_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_61_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_61_141 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_61_198 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_62_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_62_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_62_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_62_89 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_62_93 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_111 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_118 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_62_125 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_146 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_62_153 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_62_155 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_62_198 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_63_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_63_57 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_63_75 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_63_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_99 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_63_106 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_63_145 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_63_149 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_167 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_63_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_64_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_64_2 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_64_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_82 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_64_89 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_64_145 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_64_184 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_64_197 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_64_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_65_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_57 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_65_64 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_100 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_65_107 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_65_129 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_65_150 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_65_198 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_66_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_66_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_66_41 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_66_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_86 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_66_93 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_66_120 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_145 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_66_152 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_66_173 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_66_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_67_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_67_2 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_67_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_33 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_40 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_67_47 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_66 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_67_73 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_67_145 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_67_149 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_67_171 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_67_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_67_198 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_68_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_44 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_51 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_79 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_86 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_68_93 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_68_115 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_68_117 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_156 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_68_163 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_68_167 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_68_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_68_188 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_68_197 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_68_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_69_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_69_2 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_41 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_169 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_69_176 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_69_197 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_69_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_70_17 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_70_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_70_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_70_148 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_70_170 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_70_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_70_198 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_71_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_71_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_31 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_71_38 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_71_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_61 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_71_68 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_71_104 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_71_164 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_71_166 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_72_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_61 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_72_68 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_72_94 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_72_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_72_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_72_141 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_72_143 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_178 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_72_185 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_73_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_40 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_85 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_73_92 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_73_94 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_73_120 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_73_124 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_73_167 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_74_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_74_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_74_82 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_74_128 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_74_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_74_156 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_74_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_45 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_75_52 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_75_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_75_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_75_104 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_143 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_75_150 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_75_152 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_173 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_180 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_187 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_75_194 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_75_198 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_17 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_76_24 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_76_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_76_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_76_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_76_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_76_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_76_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_77_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_34 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_77_83 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_77_85 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_77_103 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_190 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_77_197 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_77_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_78_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_36 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_103 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_78_110 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_190 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_78_197 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_78_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_79_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_79_37 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_79_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_79_125 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_79_129 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_79_157 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_79_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_79_194 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_79_198 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_80_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_30 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_37 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_80_44 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_80_83 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_80_87 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_80_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_80_131 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_80_135 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_80_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_81_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_81_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_22 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_81_29 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_81_92 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_132 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_81_139 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_81_156 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_81_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_176 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_183 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_190 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_81_197 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_81_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_82_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_36 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_82_43 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_82_47 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_82_87 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_106 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_82_113 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_82_117 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_82_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_181 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_188 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_82_195 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_82_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_83_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_83_9 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_31 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_83_38 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_83_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_83_64 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_83_68 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_83_96 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_83_127 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_83_129 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_83_166 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_180 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_187 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_83_194 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_83_198 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_17 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_84_79 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_84_85 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_176 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_183 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_190 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_84_197 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_84_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_85_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_85_2 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_24 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_85_31 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_85_59 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_85_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_176 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_183 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_190 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_85_197 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_85_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_86_17 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_86_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_86_64 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_86_66 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_86_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_86_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_166 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_86_173 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_86_177 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_86_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_87_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_87_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_87_22 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_87_75 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_87_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_87_93 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_87_111 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_87_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_87_174 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_87_197 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_87_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_88_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_88_66 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_88_68 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_88_107 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_88_111 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_88_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_88_138 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_88_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_88_167 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_89_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_89_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_89_29 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_97 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_89_104 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_89_106 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_89_124 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_89_128 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_191 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_89_198 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_90_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_90_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_66 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_90_111 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_90_129 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_90_157 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_90_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_90_197 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_90_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_91_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_62 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_91_69 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_128 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_91_135 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_91_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_92_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_92_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_92_33 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_92_37 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_92_69 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_92_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_92_93 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_92_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_92_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_92_170 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_92_198 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_34 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_93_41 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_93_43 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_93_66 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_93_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_93_113 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_93_148 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_93_187 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_192 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_93_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_97 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_94_104 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_94_108 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_94_131 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_171 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_178 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_185 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_192 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_94_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_95_51 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_118 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_125 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_132 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_139 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_146 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_95_153 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_96_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_96_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_26 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_96_33 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_96_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_96_57 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_96_66 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_96_90 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_117 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_124 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_131 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_138 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_145 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_152 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_159 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_166 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_173 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_180 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_187 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_96_194 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_96_198 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_34 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_97_41 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_97_43 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_69 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_97_76 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_97_97 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_97_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_97_104 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_122 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_129 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_136 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_143 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_150 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_157 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_164 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_171 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_178 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_185 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_192 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_97_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_17 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_24 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_69 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_98_76 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_98_80 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_120 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_127 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_134 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_141 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_148 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_155 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_162 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_169 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_176 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_183 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_190 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_98_197 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_98_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_99_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_23 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_30 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_99_37 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_99_69 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_99_92 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_99_94 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_99_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_100_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_26 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_100_55 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_100_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_100_163 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_100_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_101_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_101_37 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_101_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_102_17 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_102_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_102_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_24 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_103_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_103_78 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_97 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_104 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_111 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_118 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_125 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_132 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_139 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_146 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_153 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_103_160 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_166 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_173 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_180 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_187 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_103_194 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_103_198 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_17 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_104_66 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_87 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_94 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_101 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_108 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_115 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_122 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_129 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_136 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_143 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_104_150 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_156 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_163 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_170 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_177 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_184 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_191 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_104_198 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_105_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_105_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_105_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_64 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_71 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_78 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_85 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_92 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_99 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_106 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_113 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_120 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_127 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_134 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_141 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_148 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_155 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_162 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_169 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_176 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_183 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_190 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_105_197 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_105_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_68 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_75 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_82 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_89 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_96 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_103 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_110 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_117 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_124 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_131 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_138 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_106_145 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_106_149 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_106_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_107_17 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_107_24 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_107_43 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_107_50 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_107_57 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_107_64 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_107_71 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_107_78 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_107_85 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_107_92 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_107_99 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_107_106 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_107_113 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_107_120 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_107_127 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_107_134 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_107_141 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_107_148 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_107_155 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_107_162 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_107_169 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_107_173 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_107_178 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_107_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_107_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_107_190 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_107_197 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_107_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_108_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_108_24 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_108_29 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_108_47 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_108_54 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_108_61 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_108_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_108_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_108_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_108_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_108_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_108_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_108_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_108_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_108_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_108_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_108_134 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_108_143 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_108_150 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_108_157 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_108_164 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_108_171 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_108_191 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_108_195 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_108_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_109_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_109_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_109_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_109_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_109_83 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_109_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_109_100 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_109_104 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_109_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_109_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_109_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_109_148 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_109_150 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_109_155 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_109_159 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_110_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_110_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_110_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_110_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_110_27 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_110_34 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_110_41 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_110_48 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_110_55 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_110_62 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_110_69 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_110_76 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_110_83 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_110_90 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_110_97 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_110_104 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_110_111 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_110_118 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_110_125 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_110_132 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_110_139 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_110_146 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_110_153 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_110_160 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_110_167 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_110_174 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_110_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_110_183 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_110_187 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_110_191 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_110_198 (.VDD(VPWR),
    .VSS(VGND));
endmodule
