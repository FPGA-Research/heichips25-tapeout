module LUT4AB (Ci,
    Co,
    UserCLK,
    UserCLKo,
    VPWR,
    VGND,
    E1BEG,
    E1END,
    E2BEG,
    E2BEGb,
    E2END,
    E2MID,
    E6BEG,
    E6END,
    EE4BEG,
    EE4END,
    FrameData,
    FrameData_O,
    FrameStrobe,
    FrameStrobe_O,
    N1BEG,
    N1END,
    N2BEG,
    N2BEGb,
    N2END,
    N2MID,
    N4BEG,
    N4END,
    NN4BEG,
    NN4END,
    S1BEG,
    S1END,
    S2BEG,
    S2BEGb,
    S2END,
    S2MID,
    S4BEG,
    S4END,
    SS4BEG,
    SS4END,
    W1BEG,
    W1END,
    W2BEG,
    W2BEGb,
    W2END,
    W2MID,
    W6BEG,
    W6END,
    WW4BEG,
    WW4END);
 input Ci;
 output Co;
 input UserCLK;
 output UserCLKo;
 inout VPWR;
 inout VGND;
 output [3:0] E1BEG;
 input [3:0] E1END;
 output [7:0] E2BEG;
 output [7:0] E2BEGb;
 input [7:0] E2END;
 input [7:0] E2MID;
 output [11:0] E6BEG;
 input [11:0] E6END;
 output [15:0] EE4BEG;
 input [15:0] EE4END;
 input [31:0] FrameData;
 output [31:0] FrameData_O;
 input [19:0] FrameStrobe;
 output [19:0] FrameStrobe_O;
 output [3:0] N1BEG;
 input [3:0] N1END;
 output [7:0] N2BEG;
 output [7:0] N2BEGb;
 input [7:0] N2END;
 input [7:0] N2MID;
 output [15:0] N4BEG;
 input [15:0] N4END;
 output [15:0] NN4BEG;
 input [15:0] NN4END;
 output [3:0] S1BEG;
 input [3:0] S1END;
 output [7:0] S2BEG;
 output [7:0] S2BEGb;
 input [7:0] S2END;
 input [7:0] S2MID;
 output [15:0] S4BEG;
 input [15:0] S4END;
 output [15:0] SS4BEG;
 input [15:0] SS4END;
 output [3:0] W1BEG;
 input [3:0] W1END;
 output [7:0] W2BEG;
 output [7:0] W2BEGb;
 input [7:0] W2END;
 input [7:0] W2MID;
 output [11:0] W6BEG;
 input [11:0] W6END;
 output [15:0] WW4BEG;
 input [15:0] WW4END;

 wire A;
 wire B;
 wire C;
 wire D;
 wire E;
 wire F;
 wire G;
 wire H;
 wire \Inst_LA_LUT4c_frame_config_dffesr.LUT_flop ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.c_I0mux ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.c_out_mux ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.c_reset_value ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.LUT_flop ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.c_I0mux ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.c_out_mux ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.c_reset_value ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.LUT_flop ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.c_I0mux ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.c_out_mux ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.c_reset_value ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.LUT_flop ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.c_I0mux ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.c_out_mux ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.c_reset_value ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.LUT_flop ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.c_I0mux ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.c_out_mux ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.c_reset_value ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.LUT_flop ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.c_I0mux ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.c_out_mux ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.c_reset_value ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.LUT_flop ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.c_I0mux ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.c_out_mux ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.c_reset_value ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.LUT_flop ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.c_I0mux ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.c_out_mux ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.c_reset_value ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit0.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit1.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit10.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit11.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit12.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit13.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit14.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit15.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit16.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit17.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit18.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit19.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit2.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit20.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit21.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit22.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit23.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit24.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit25.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit26.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit27.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit28.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit29.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit3.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit30.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit31.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit4.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit5.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit6.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit7.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit8.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit9.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit0.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit1.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit10.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit11.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit12.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit13.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit14.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit15.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit16.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit17.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit18.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit19.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit2.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit20.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit21.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit22.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit23.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit24.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit25.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit26.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit27.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit28.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit29.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit3.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit30.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit31.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit4.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit5.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit6.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit7.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit8.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit9.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit0.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit1.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit10.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit11.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit12.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit13.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit14.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit15.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit16.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit17.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit18.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit19.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit2.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit20.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit21.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit22.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit23.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit24.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit25.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit26.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit27.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit28.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit29.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit3.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit30.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit31.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit4.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit5.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit6.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit7.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit8.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit9.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit0.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit1.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit10.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit11.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit12.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit13.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit14.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit15.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit16.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit17.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit18.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit19.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit2.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit20.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit21.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit22.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit23.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit24.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit25.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit26.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit27.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit28.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit29.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit3.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit30.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit31.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit4.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit5.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit6.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit7.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit8.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit9.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit0.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit1.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit10.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit11.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit12.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit13.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit14.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit15.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit16.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit17.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit18.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit19.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit2.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit20.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit21.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit22.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit23.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit24.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit25.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit26.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit27.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit28.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit29.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit3.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit30.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit31.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit4.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit5.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit6.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit7.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit8.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit9.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame14_bit16.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame14_bit17.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame14_bit18.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame14_bit19.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame14_bit20.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame14_bit21.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame14_bit22.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame14_bit23.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame14_bit24.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame14_bit25.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame14_bit26.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame14_bit27.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame14_bit28.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame14_bit29.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame14_bit30.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame14_bit31.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit0.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit1.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit10.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit11.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit12.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit13.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit14.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit15.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit16.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit17.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit18.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit19.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit2.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit20.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit21.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit22.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit23.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit24.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit25.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit26.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit27.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit28.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit29.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit3.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit30.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit31.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit4.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit5.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit6.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit7.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit8.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit9.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit0.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit1.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit10.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit11.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit12.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit13.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit14.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit15.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit16.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit17.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit18.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit19.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit2.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit20.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit21.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit22.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit23.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit24.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit25.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit26.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit27.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit28.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit29.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit3.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit30.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit31.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit4.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit5.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit6.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit7.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit8.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit9.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit0.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit1.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit10.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit11.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit12.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit13.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit14.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit15.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit16.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit17.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit18.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit19.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit2.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit20.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit21.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit22.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit23.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit24.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit25.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit26.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit27.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit28.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit29.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit3.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit30.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit31.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit4.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit5.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit6.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit7.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit8.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit9.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit0.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit1.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit10.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit11.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit12.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit13.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit14.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit15.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit16.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit17.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit18.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit19.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit2.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit20.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit21.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit22.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit23.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit24.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit25.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit26.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit27.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit28.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit29.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit3.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit30.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit31.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit4.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit5.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit6.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit7.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit8.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit9.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit0.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit1.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit10.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit11.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit12.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit13.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit14.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit15.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit16.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit17.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit18.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit19.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit2.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit20.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit21.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit22.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit23.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit24.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit25.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit26.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit27.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit28.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit29.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit3.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit30.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit31.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit4.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit5.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit6.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit7.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit8.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit9.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit0.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit1.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit10.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit11.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit12.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit13.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit14.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit15.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit16.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit17.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit18.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit19.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit2.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit20.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit21.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit22.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit23.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit24.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit25.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit26.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit27.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit28.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit29.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit3.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit30.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit31.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit4.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit5.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit6.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit7.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit8.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit9.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit0.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit1.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit10.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit11.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit12.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit13.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit14.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit15.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit16.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit17.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit18.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit19.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit2.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit20.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit21.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit22.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit23.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit24.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit25.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit26.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit27.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit28.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit29.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit3.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit30.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit31.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit4.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit5.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit6.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit7.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit8.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit9.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit0.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit1.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit10.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit11.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit12.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit13.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit14.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit15.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit16.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit17.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit18.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit19.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit2.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit20.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit21.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit22.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit23.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit24.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit25.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit26.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit27.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit28.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit29.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit3.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit30.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit31.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit4.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit5.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit6.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit7.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit8.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit9.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit0.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit1.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit10.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit11.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit12.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit13.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit14.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit15.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit16.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit17.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit18.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit19.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit2.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit20.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit21.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit22.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit23.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit24.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit25.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit26.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit27.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit28.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit29.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit3.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit30.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit31.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit4.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit5.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit6.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit7.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit8.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit9.Q ;
 wire \Inst_LUT4AB_switch_matrix.E1BEG0 ;
 wire \Inst_LUT4AB_switch_matrix.E1BEG1 ;
 wire \Inst_LUT4AB_switch_matrix.E1BEG2 ;
 wire \Inst_LUT4AB_switch_matrix.E1BEG3 ;
 wire \Inst_LUT4AB_switch_matrix.E2BEG0 ;
 wire \Inst_LUT4AB_switch_matrix.E2BEG1 ;
 wire \Inst_LUT4AB_switch_matrix.E2BEG2 ;
 wire \Inst_LUT4AB_switch_matrix.E2BEG3 ;
 wire \Inst_LUT4AB_switch_matrix.E2BEG4 ;
 wire \Inst_LUT4AB_switch_matrix.E2BEG5 ;
 wire \Inst_LUT4AB_switch_matrix.E2BEG6 ;
 wire \Inst_LUT4AB_switch_matrix.E2BEG7 ;
 wire \Inst_LUT4AB_switch_matrix.E6BEG0 ;
 wire \Inst_LUT4AB_switch_matrix.E6BEG1 ;
 wire \Inst_LUT4AB_switch_matrix.EE4BEG0 ;
 wire \Inst_LUT4AB_switch_matrix.EE4BEG1 ;
 wire \Inst_LUT4AB_switch_matrix.EE4BEG2 ;
 wire \Inst_LUT4AB_switch_matrix.EE4BEG3 ;
 wire \Inst_LUT4AB_switch_matrix.JN2BEG0 ;
 wire \Inst_LUT4AB_switch_matrix.JN2BEG1 ;
 wire \Inst_LUT4AB_switch_matrix.JN2BEG2 ;
 wire \Inst_LUT4AB_switch_matrix.JN2BEG3 ;
 wire \Inst_LUT4AB_switch_matrix.JN2BEG4 ;
 wire \Inst_LUT4AB_switch_matrix.JN2BEG5 ;
 wire \Inst_LUT4AB_switch_matrix.JN2BEG6 ;
 wire \Inst_LUT4AB_switch_matrix.JN2BEG7 ;
 wire \Inst_LUT4AB_switch_matrix.JS2BEG0 ;
 wire \Inst_LUT4AB_switch_matrix.JS2BEG1 ;
 wire \Inst_LUT4AB_switch_matrix.JS2BEG2 ;
 wire \Inst_LUT4AB_switch_matrix.JS2BEG3 ;
 wire \Inst_LUT4AB_switch_matrix.JS2BEG4 ;
 wire \Inst_LUT4AB_switch_matrix.JS2BEG5 ;
 wire \Inst_LUT4AB_switch_matrix.JS2BEG6 ;
 wire \Inst_LUT4AB_switch_matrix.JS2BEG7 ;
 wire \Inst_LUT4AB_switch_matrix.JW2BEG0 ;
 wire \Inst_LUT4AB_switch_matrix.JW2BEG1 ;
 wire \Inst_LUT4AB_switch_matrix.JW2BEG2 ;
 wire \Inst_LUT4AB_switch_matrix.JW2BEG3 ;
 wire \Inst_LUT4AB_switch_matrix.JW2BEG4 ;
 wire \Inst_LUT4AB_switch_matrix.JW2BEG5 ;
 wire \Inst_LUT4AB_switch_matrix.JW2BEG6 ;
 wire \Inst_LUT4AB_switch_matrix.JW2BEG7 ;
 wire \Inst_LUT4AB_switch_matrix.M_AB ;
 wire \Inst_LUT4AB_switch_matrix.M_AD ;
 wire \Inst_LUT4AB_switch_matrix.M_AH ;
 wire \Inst_LUT4AB_switch_matrix.M_EF ;
 wire \Inst_LUT4AB_switch_matrix.N1BEG0 ;
 wire \Inst_LUT4AB_switch_matrix.N1BEG1 ;
 wire \Inst_LUT4AB_switch_matrix.N1BEG2 ;
 wire \Inst_LUT4AB_switch_matrix.N1BEG3 ;
 wire \Inst_LUT4AB_switch_matrix.N4BEG0 ;
 wire \Inst_LUT4AB_switch_matrix.N4BEG1 ;
 wire \Inst_LUT4AB_switch_matrix.N4BEG2 ;
 wire \Inst_LUT4AB_switch_matrix.N4BEG3 ;
 wire \Inst_LUT4AB_switch_matrix.NN4BEG0 ;
 wire \Inst_LUT4AB_switch_matrix.NN4BEG1 ;
 wire \Inst_LUT4AB_switch_matrix.NN4BEG2 ;
 wire \Inst_LUT4AB_switch_matrix.NN4BEG3 ;
 wire \Inst_LUT4AB_switch_matrix.S1BEG0 ;
 wire \Inst_LUT4AB_switch_matrix.S1BEG1 ;
 wire \Inst_LUT4AB_switch_matrix.S1BEG2 ;
 wire \Inst_LUT4AB_switch_matrix.S1BEG3 ;
 wire \Inst_LUT4AB_switch_matrix.S4BEG0 ;
 wire \Inst_LUT4AB_switch_matrix.S4BEG1 ;
 wire \Inst_LUT4AB_switch_matrix.S4BEG2 ;
 wire \Inst_LUT4AB_switch_matrix.S4BEG3 ;
 wire \Inst_LUT4AB_switch_matrix.SS4BEG0 ;
 wire \Inst_LUT4AB_switch_matrix.SS4BEG1 ;
 wire \Inst_LUT4AB_switch_matrix.SS4BEG2 ;
 wire \Inst_LUT4AB_switch_matrix.SS4BEG3 ;
 wire \Inst_LUT4AB_switch_matrix.W1BEG0 ;
 wire \Inst_LUT4AB_switch_matrix.W1BEG1 ;
 wire \Inst_LUT4AB_switch_matrix.W1BEG2 ;
 wire \Inst_LUT4AB_switch_matrix.W1BEG3 ;
 wire \Inst_LUT4AB_switch_matrix.W6BEG0 ;
 wire \Inst_LUT4AB_switch_matrix.W6BEG1 ;
 wire \Inst_LUT4AB_switch_matrix.WW4BEG0 ;
 wire \Inst_LUT4AB_switch_matrix.WW4BEG1 ;
 wire \Inst_LUT4AB_switch_matrix.WW4BEG2 ;
 wire \Inst_LUT4AB_switch_matrix.WW4BEG3 ;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire UserCLK_regs;
 wire clknet_0_UserCLK;
 wire clknet_1_0__leaf_UserCLK;
 wire clknet_0_UserCLK_regs;
 wire clknet_1_0__leaf_UserCLK_regs;
 wire clknet_1_1__leaf_UserCLK_regs;

 sg13g2_inv_1 _1171_ (.VDD(VPWR),
    .Y(_1012_),
    .A(N4END[0]),
    .VSS(VGND));
 sg13g2_inv_1 _1172_ (.VDD(VPWR),
    .Y(_1013_),
    .A(E1END[2]),
    .VSS(VGND));
 sg13g2_inv_1 _1173_ (.VDD(VPWR),
    .Y(_1014_),
    .A(E6END[0]),
    .VSS(VGND));
 sg13g2_inv_1 _1174_ (.VDD(VPWR),
    .Y(_1015_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit8.Q ),
    .VSS(VGND));
 sg13g2_inv_1 _1175_ (.VDD(VPWR),
    .Y(_1016_),
    .A(E1END[0]),
    .VSS(VGND));
 sg13g2_inv_1 _1176_ (.VDD(VPWR),
    .Y(_1017_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit7.Q ),
    .VSS(VGND));
 sg13g2_inv_1 _1177_ (.VDD(VPWR),
    .Y(_1018_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit8.Q ),
    .VSS(VGND));
 sg13g2_inv_1 _1178_ (.VDD(VPWR),
    .Y(_1019_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit9.Q ),
    .VSS(VGND));
 sg13g2_inv_1 _1179_ (.VDD(VPWR),
    .Y(_1020_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit0.Q ),
    .VSS(VGND));
 sg13g2_inv_1 _1180_ (.VDD(VPWR),
    .Y(_1021_),
    .A(N2MID[4]),
    .VSS(VGND));
 sg13g2_inv_1 _1181_ (.VDD(VPWR),
    .Y(_1022_),
    .A(S4END[0]),
    .VSS(VGND));
 sg13g2_inv_1 _1182_ (.VDD(VPWR),
    .Y(_1023_),
    .A(WW4END[2]),
    .VSS(VGND));
 sg13g2_inv_1 _1183_ (.VDD(VPWR),
    .Y(_1024_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit8.Q ),
    .VSS(VGND));
 sg13g2_inv_1 _1184_ (.VDD(VPWR),
    .Y(_1025_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit9.Q ),
    .VSS(VGND));
 sg13g2_inv_1 _1185_ (.VDD(VPWR),
    .Y(_1026_),
    .A(W2MID[4]),
    .VSS(VGND));
 sg13g2_inv_1 _1186_ (.VDD(VPWR),
    .Y(_1027_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit0.Q ),
    .VSS(VGND));
 sg13g2_inv_1 _1187_ (.VDD(VPWR),
    .Y(_1028_),
    .A(W6END[1]),
    .VSS(VGND));
 sg13g2_inv_1 _1188_ (.VDD(VPWR),
    .Y(_1029_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit8.Q ),
    .VSS(VGND));
 sg13g2_inv_1 _1189_ (.VDD(VPWR),
    .Y(_1030_),
    .A(WW4END[1]),
    .VSS(VGND));
 sg13g2_inv_1 _1190_ (.VDD(VPWR),
    .Y(_1031_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit4.Q ),
    .VSS(VGND));
 sg13g2_inv_1 _1191_ (.VDD(VPWR),
    .Y(_1032_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit4.Q ),
    .VSS(VGND));
 sg13g2_inv_1 _1192_ (.VDD(VPWR),
    .Y(_1033_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit5.Q ),
    .VSS(VGND));
 sg13g2_inv_1 _1193_ (.VDD(VPWR),
    .Y(_1034_),
    .A(S2MID[4]),
    .VSS(VGND));
 sg13g2_inv_1 _1194_ (.VDD(VPWR),
    .Y(_1035_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit13.Q ),
    .VSS(VGND));
 sg13g2_inv_1 _1195_ (.VDD(VPWR),
    .Y(_1036_),
    .A(S4END[1]),
    .VSS(VGND));
 sg13g2_inv_1 _1196_ (.VDD(VPWR),
    .Y(_1037_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit4.Q ),
    .VSS(VGND));
 sg13g2_inv_1 _1197_ (.VDD(VPWR),
    .Y(_1038_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit5.Q ),
    .VSS(VGND));
 sg13g2_inv_1 _1198_ (.VDD(VPWR),
    .Y(_1039_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit12.Q ),
    .VSS(VGND));
 sg13g2_inv_1 _1199_ (.VDD(VPWR),
    .Y(_1040_),
    .A(EE4END[3]),
    .VSS(VGND));
 sg13g2_inv_1 _1200_ (.VDD(VPWR),
    .Y(_1041_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit13.Q ),
    .VSS(VGND));
 sg13g2_inv_1 _1201_ (.VDD(VPWR),
    .Y(_1042_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit16.Q ),
    .VSS(VGND));
 sg13g2_inv_1 _1202_ (.VDD(VPWR),
    .Y(_1043_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit17.Q ),
    .VSS(VGND));
 sg13g2_inv_1 _1203_ (.VDD(VPWR),
    .Y(_1044_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit20.Q ),
    .VSS(VGND));
 sg13g2_inv_1 _1204_ (.VDD(VPWR),
    .Y(_1045_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit24.Q ),
    .VSS(VGND));
 sg13g2_inv_1 _1205_ (.VDD(VPWR),
    .Y(_1046_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit25.Q ),
    .VSS(VGND));
 sg13g2_inv_1 _1206_ (.VDD(VPWR),
    .Y(_1047_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit21.Q ),
    .VSS(VGND));
 sg13g2_inv_1 _1207_ (.VDD(VPWR),
    .Y(_1048_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit19.Q ),
    .VSS(VGND));
 sg13g2_inv_1 _1208_ (.VDD(VPWR),
    .Y(_1049_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit8.Q ),
    .VSS(VGND));
 sg13g2_inv_1 _1209_ (.VDD(VPWR),
    .Y(_1050_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit7.Q ),
    .VSS(VGND));
 sg13g2_inv_1 _1210_ (.VDD(VPWR),
    .Y(_1051_),
    .A(G),
    .VSS(VGND));
 sg13g2_inv_1 _1211_ (.VDD(VPWR),
    .Y(_1052_),
    .A(H),
    .VSS(VGND));
 sg13g2_mux4_1 _1212_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit30.Q ),
    .A0(F),
    .A1(G),
    .A2(H),
    .A3(\Inst_LUT4AB_switch_matrix.M_AB ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit31.Q ),
    .X(_1053_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _1213_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit31.Q ),
    .A0(A),
    .A1(D),
    .A2(C),
    .A3(E),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit30.Q ),
    .X(_1054_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _1214_ (.A0(_1053_),
    .A1(_1054_),
    .S(_1020_),
    .X(_1055_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1215_ (.Y(_1056_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit1.Q ),
    .B(_1055_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _1216_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit30.Q ),
    .A0(N1END[0]),
    .A1(N2END[2]),
    .A2(N4END[2]),
    .A3(E2END[2]),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit31.Q ),
    .X(_1057_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _1217_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit0.Q ),
    .B(_1057_),
    .Y(_1058_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _1218_ (.A0(E6END[0]),
    .A1(S2END[2]),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit30.Q ),
    .X(_1059_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _1219_ (.Y(_1060_),
    .B(_1059_),
    .A_N(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit31.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _1220_ (.A0(W2END[2]),
    .A1(WW4END[3]),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit30.Q ),
    .X(_1061_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1221_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit31.Q ),
    .A2(_1061_),
    .Y(_1062_),
    .B1(_1020_));
 sg13g2_a21o_1 _1222_ (.A2(_1062_),
    .A1(_1060_),
    .B1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit1.Q ),
    .X(_1063_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1223_ (.B1(_1056_),
    .VDD(VPWR),
    .Y(\Inst_LUT4AB_switch_matrix.E2BEG1 ),
    .VSS(VGND),
    .A1(_1058_),
    .A2(_1063_));
 sg13g2_inv_1 _1224_ (.VDD(VPWR),
    .Y(_1064_),
    .A(\Inst_LUT4AB_switch_matrix.E2BEG1 ),
    .VSS(VGND));
 sg13g2_mux4_1 _1225_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit28.Q ),
    .A0(EE4END[2]),
    .A1(S4END[2]),
    .A2(W2END[7]),
    .A3(\Inst_LUT4AB_switch_matrix.E2BEG1 ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit29.Q ),
    .X(_1065_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _1226_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit29.Q ),
    .A0(NN4END[0]),
    .A1(S2END[2]),
    .A2(E2END[2]),
    .A3(W2END[2]),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit28.Q ),
    .X(_1066_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _1227_ (.A0(H),
    .A1(\Inst_LUT4AB_switch_matrix.M_AH ),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit6.Q ),
    .X(_1067_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1228_ (.Y(_1068_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit7.Q ),
    .B(_1067_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _1229_ (.A0(F),
    .A1(G),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit6.Q ),
    .X(_1069_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1230_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1017_),
    .A2(_1069_),
    .Y(_1070_),
    .B1(_1018_));
 sg13g2_mux2_1 _1231_ (.A0(C),
    .A1(E),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit6.Q ),
    .X(_1071_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1232_ (.Y(_1072_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit7.Q ),
    .B(_1071_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _1233_ (.A0(A),
    .A1(B),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit6.Q ),
    .X(_1073_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1234_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1017_),
    .A2(_1073_),
    .Y(_1074_),
    .B1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit8.Q ));
 sg13g2_a221oi_1 _1235_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_1074_),
    .C1(_1019_),
    .B1(_1072_),
    .A1(_1068_),
    .Y(_1075_),
    .A2(_1070_));
 sg13g2_mux4_1 _1236_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit6.Q ),
    .A0(N1END[2]),
    .A1(N2END[4]),
    .A2(N4END[0]),
    .A3(E2END[4]),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit7.Q ),
    .X(_1076_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _1237_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit8.Q ),
    .B(_1076_),
    .Y(_1077_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _1238_ (.A0(W2END[4]),
    .A1(W6END[0]),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit6.Q ),
    .X(_1078_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _1239_ (.A0(E6END[0]),
    .A1(S2END[4]),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit6.Q ),
    .X(_1079_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1240_ (.Y(_1080_),
    .A(_1017_),
    .B(_1079_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1241_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit7.Q ),
    .A2(_1078_),
    .Y(_1081_),
    .B1(_1018_));
 sg13g2_a21oi_1 _1242_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1080_),
    .A2(_1081_),
    .Y(_1082_),
    .B1(_1077_));
 sg13g2_a21o_1 _1243_ (.A2(_1082_),
    .A1(_1019_),
    .B1(_1075_),
    .X(\Inst_LUT4AB_switch_matrix.E2BEG3 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _1244_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit28.Q ),
    .A0(E2MID[2]),
    .A1(S2MID[2]),
    .A2(W2MID[2]),
    .A3(\Inst_LUT4AB_switch_matrix.E2BEG3 ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit29.Q ),
    .X(_1083_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _1245_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit28.Q ),
    .A0(N2MID[3]),
    .A1(E2MID[3]),
    .A2(S2MID[3]),
    .A3(W2MID[3]),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit29.Q ),
    .X(_1084_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _1246_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit4.Q ),
    .A0(_1083_),
    .A1(_1084_),
    .A2(_1066_),
    .A3(_1065_),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit5.Q ),
    .X(_1085_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _1247_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit6.Q ),
    .A0(A),
    .A1(B),
    .A2(C),
    .A3(E),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit7.Q ),
    .X(_1086_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _1248_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit6.Q ),
    .B(F),
    .Y(_1087_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1249_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit6.Q ),
    .A2(_1051_),
    .Y(_1088_),
    .B1(_1087_));
 sg13g2_nand2b_1 _1250_ (.Y(_1089_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit6.Q ),
    .A_N(\Inst_LUT4AB_switch_matrix.M_EF ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1251_ (.B1(_1089_),
    .VDD(VPWR),
    .Y(_1090_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit6.Q ),
    .A2(H));
 sg13g2_o21ai_1 _1252_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit8.Q ),
    .VDD(VPWR),
    .Y(_1091_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit7.Q ),
    .A2(_1088_));
 sg13g2_a21oi_1 _1253_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit7.Q ),
    .A2(_1090_),
    .Y(_1092_),
    .B1(_1091_));
 sg13g2_nand2b_1 _1254_ (.Y(_1093_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit9.Q ),
    .A_N(_1092_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1255_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1015_),
    .A2(_1086_),
    .Y(_1094_),
    .B1(_1093_));
 sg13g2_mux2_1 _1256_ (.A0(E6END[0]),
    .A1(S2END[4]),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit6.Q ),
    .X(_1095_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _1257_ (.A0(W2END[4]),
    .A1(W6END[0]),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit6.Q ),
    .X(_1096_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _1258_ (.A0(E1END[2]),
    .A1(E2END[4]),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit6.Q ),
    .X(_1097_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _1259_ (.A(N2END[4]),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit6.Q ),
    .Y(_1098_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1260_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1012_),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit6.Q ),
    .Y(_1099_),
    .B1(_1098_));
 sg13g2_mux4_1 _1261_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit7.Q ),
    .A0(_1095_),
    .A1(_1096_),
    .A2(_1099_),
    .A3(_1097_),
    .S1(_1015_),
    .X(_1100_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _1262_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit9.Q ),
    .B(_1100_),
    .Y(_1101_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _1263_ (.A(_1094_),
    .B(_1101_),
    .Y(\Inst_LUT4AB_switch_matrix.JN2BEG3 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _1264_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit26.Q ),
    .A0(N2MID[6]),
    .A1(S2MID[6]),
    .A2(W2MID[6]),
    .A3(\Inst_LUT4AB_switch_matrix.JN2BEG3 ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit27.Q ),
    .X(_1102_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _1265_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit26.Q ),
    .A0(N2MID[7]),
    .A1(E2MID[7]),
    .A2(S2MID[7]),
    .A3(W2MID[7]),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit27.Q ),
    .X(_1103_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _1266_ (.VDD(VPWR),
    .Y(_1104_),
    .A(_1103_),
    .VSS(VGND));
 sg13g2_mux4_1 _1267_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit30.Q ),
    .A0(F),
    .A1(G),
    .A2(H),
    .A3(\Inst_LUT4AB_switch_matrix.M_AD ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit31.Q ),
    .X(_1105_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _1268_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit31.Q ),
    .A0(A),
    .A1(D),
    .A2(C),
    .A3(E),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit30.Q ),
    .X(_1106_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _1269_ (.Y(_1107_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit0.Q ),
    .A_N(_1105_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1270_ (.B1(_1107_),
    .VDD(VPWR),
    .Y(_1108_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit0.Q ),
    .A2(_1106_));
 sg13g2_mux4_1 _1271_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit31.Q ),
    .A0(N2END[2]),
    .A1(E1END[0]),
    .A2(N4END[2]),
    .A3(E2END[2]),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit30.Q ),
    .X(_1109_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _1272_ (.Y(_1110_),
    .B(_1109_),
    .A_N(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit0.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1273_ (.Y(_1111_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit30.Q ),
    .B(S2END[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1274_ (.B1(_1111_),
    .VDD(VPWR),
    .Y(_1112_),
    .VSS(VGND),
    .A1(_1014_),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit30.Q ));
 sg13g2_nand2b_1 _1275_ (.Y(_1113_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit30.Q ),
    .A_N(W6END[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1276_ (.B1(_1113_),
    .VDD(VPWR),
    .Y(_1114_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit30.Q ),
    .A2(W2END[2]));
 sg13g2_o21ai_1 _1277_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit0.Q ),
    .VDD(VPWR),
    .Y(_1115_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit31.Q ),
    .A2(_1112_));
 sg13g2_a21oi_1 _1278_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit31.Q ),
    .A2(_1114_),
    .Y(_1116_),
    .B1(_1115_));
 sg13g2_nor2_1 _1279_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit1.Q ),
    .B(_1116_),
    .Y(_1117_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _1280_ (.Y(\Inst_LUT4AB_switch_matrix.JN2BEG1 ),
    .B1(_1110_),
    .B2(_1117_),
    .A2(_1108_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit1.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _1281_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit27.Q ),
    .A0(NN4END[3]),
    .A1(WW4END[0]),
    .A2(S4END[3]),
    .A3(\Inst_LUT4AB_switch_matrix.JN2BEG1 ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit26.Q ),
    .X(_1118_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _1282_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit27.Q ),
    .A0(N2END[6]),
    .A1(SS4END[3]),
    .A2(E2END[6]),
    .A3(W2END[6]),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit26.Q ),
    .X(_1119_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _1283_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit2.Q ),
    .A0(_1102_),
    .A1(_1103_),
    .A2(_1119_),
    .A3(_1118_),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit3.Q ),
    .X(_1120_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _1284_ (.A0(_1120_),
    .A1(Ci),
    .S(\Inst_LA_LUT4c_frame_config_dffesr.c_I0mux ),
    .X(_1121_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _1285_ (.Y(_1122_),
    .B(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ),
    .A_N(_1121_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1286_ (.Y(_1123_),
    .A(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ),
    .B(_1121_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _1287_ (.B(_1122_),
    .C(_1123_),
    .A(_1085_),
    .Y(_1124_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _1288_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit30.Q ),
    .B_N(F),
    .Y(_1125_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1289_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit30.Q ),
    .A2(G),
    .Y(_1126_),
    .B1(_1125_));
 sg13g2_mux2_1 _1290_ (.A0(H),
    .A1(\Inst_LUT4AB_switch_matrix.M_EF ),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit30.Q ),
    .X(_1127_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1291_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit31.Q ),
    .A2(_1127_),
    .Y(_1128_),
    .B1(_1027_));
 sg13g2_o21ai_1 _1292_ (.B1(_1128_),
    .VDD(VPWR),
    .Y(_1129_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit31.Q ),
    .A2(_1126_));
 sg13g2_mux4_1 _1293_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit31.Q ),
    .A0(A),
    .A1(D),
    .A2(C),
    .A3(E),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit30.Q ),
    .X(_1130_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _1294_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit0.Q ),
    .B(_1130_),
    .Y(_1131_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _1295_ (.A(_1131_),
    .B_N(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit1.Q ),
    .Y(_1132_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _1296_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit31.Q ),
    .A0(NN4END[2]),
    .A1(EE4END[2]),
    .A2(E1END[0]),
    .A3(E6END[0]),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit30.Q ),
    .X(_1133_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _1297_ (.VDD(VPWR),
    .Y(_1134_),
    .A(_1133_),
    .VSS(VGND));
 sg13g2_mux2_1 _1298_ (.A0(S4END[2]),
    .A1(SS4END[2]),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit30.Q ),
    .X(_1135_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _1299_ (.Y(_1136_),
    .B(_1135_),
    .A_N(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit31.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _1300_ (.A0(W2END[2]),
    .A1(W6END[0]),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit30.Q ),
    .X(_1137_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1301_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit31.Q ),
    .A2(_1137_),
    .Y(_1138_),
    .B1(_1027_));
 sg13g2_a221oi_1 _1302_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_1138_),
    .C1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit1.Q ),
    .B1(_1136_),
    .A1(_1027_),
    .Y(_1139_),
    .A2(_1134_));
 sg13g2_a21o_1 _1303_ (.A2(_1132_),
    .A1(_1129_),
    .B1(_1139_),
    .X(\Inst_LUT4AB_switch_matrix.JS2BEG1 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _1304_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit30.Q ),
    .A0(N4END[1]),
    .A1(E6END[1]),
    .A2(W6END[1]),
    .A3(\Inst_LUT4AB_switch_matrix.JS2BEG1 ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit31.Q ),
    .X(_1140_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _1305_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit31.Q ),
    .A0(N2END[4]),
    .A1(S2END[4]),
    .A2(EE4END[0]),
    .A3(W2END[4]),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit30.Q ),
    .X(_1141_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _1306_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit6.Q ),
    .A0(A),
    .A1(B),
    .A2(C),
    .A3(E),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit7.Q ),
    .X(_1142_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _1307_ (.VDD(VPWR),
    .Y(_1143_),
    .A(_1142_),
    .VSS(VGND));
 sg13g2_mux2_1 _1308_ (.A0(F),
    .A1(G),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit6.Q ),
    .X(_1144_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _1309_ (.Y(_1145_),
    .B(_1144_),
    .A_N(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit7.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _1310_ (.A0(H),
    .A1(\Inst_LUT4AB_switch_matrix.M_AD ),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit6.Q ),
    .X(_1146_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1311_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit7.Q ),
    .A2(_1146_),
    .Y(_1147_),
    .B1(_1024_));
 sg13g2_a221oi_1 _1312_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_1147_),
    .C1(_1025_),
    .B1(_1145_),
    .A1(_1024_),
    .Y(_1148_),
    .A2(_1143_));
 sg13g2_nor2b_1 _1313_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit6.Q ),
    .B_N(S2END[4]),
    .Y(_1149_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1314_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit6.Q ),
    .A2(S4END[0]),
    .Y(_1150_),
    .B1(_1149_));
 sg13g2_mux2_1 _1315_ (.A0(W2END[4]),
    .A1(WW4END[2]),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit6.Q ),
    .X(_1151_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1316_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit7.Q ),
    .A2(_1151_),
    .Y(_1152_),
    .B1(_1024_));
 sg13g2_o21ai_1 _1317_ (.B1(_1152_),
    .VDD(VPWR),
    .Y(_1153_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit7.Q ),
    .A2(_1150_));
 sg13g2_mux4_1 _1318_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit6.Q ),
    .A0(N2END[4]),
    .A1(E1END[2]),
    .A2(E2END[4]),
    .A3(E6END[0]),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit7.Q ),
    .X(_1154_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _1319_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit8.Q ),
    .B(_1154_),
    .Y(_1155_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _1320_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit9.Q ),
    .B(_1155_),
    .Y(_1156_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _1321_ (.A2(_1156_),
    .A1(_1153_),
    .B1(_1148_),
    .X(\Inst_LUT4AB_switch_matrix.JS2BEG3 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _1322_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit30.Q ),
    .A0(N2MID[4]),
    .A1(E2MID[4]),
    .A2(W2MID[4]),
    .A3(\Inst_LUT4AB_switch_matrix.JS2BEG3 ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit31.Q ),
    .X(_1157_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _1323_ (.VDD(VPWR),
    .Y(_1158_),
    .A(_1157_),
    .VSS(VGND));
 sg13g2_mux4_1 _1324_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit30.Q ),
    .A0(N2MID[5]),
    .A1(E2MID[5]),
    .A2(S2MID[5]),
    .A3(W2MID[5]),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit31.Q ),
    .X(_1159_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _1325_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit6.Q ),
    .A0(_1157_),
    .A1(_1159_),
    .A2(_1141_),
    .A3(_1140_),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit7.Q ),
    .X(_1160_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _1326_ (.A0(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ),
    .A1(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ),
    .S(_1121_),
    .X(_1161_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _1327_ (.A(_1085_),
    .B(_1161_),
    .Y(_1162_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _1328_ (.A(_1160_),
    .B(_1162_),
    .Y(_0008_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _1329_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit30.Q ),
    .A0(F),
    .A1(G),
    .A2(H),
    .A3(\Inst_LUT4AB_switch_matrix.M_AH ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit31.Q ),
    .X(_0009_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _1330_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit31.Q ),
    .A0(A),
    .A1(D),
    .A2(C),
    .A3(E),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit30.Q ),
    .X(_0010_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _1331_ (.Y(_0011_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit0.Q ),
    .A_N(_0009_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1332_ (.B1(_0011_),
    .VDD(VPWR),
    .Y(_0012_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit0.Q ),
    .A2(_0010_));
 sg13g2_mux4_1 _1333_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit31.Q ),
    .A0(N1END[0]),
    .A1(E2END[2]),
    .A2(N2END[2]),
    .A3(E6END[0]),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit30.Q ),
    .X(_0013_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _1334_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit0.Q ),
    .B_N(_0013_),
    .Y(_0014_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _1335_ (.A0(S2END[2]),
    .A1(S4END[2]),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit30.Q ),
    .X(_0015_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _1336_ (.Y(_0016_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit30.Q ),
    .A_N(W6END[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1337_ (.B1(_0016_),
    .VDD(VPWR),
    .Y(_0017_),
    .VSS(VGND),
    .A1(W2END[2]),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit30.Q ));
 sg13g2_o21ai_1 _1338_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit0.Q ),
    .VDD(VPWR),
    .Y(_0018_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit31.Q ),
    .A2(_0015_));
 sg13g2_a21oi_1 _1339_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit31.Q ),
    .A2(_0017_),
    .Y(_0019_),
    .B1(_0018_));
 sg13g2_nor3_1 _1340_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit1.Q ),
    .B(_0014_),
    .C(_0019_),
    .Y(_0020_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _1341_ (.A2(_0012_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit1.Q ),
    .B1(_0020_),
    .X(_0021_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _1342_ (.VDD(VPWR),
    .Y(\Inst_LUT4AB_switch_matrix.JW2BEG1 ),
    .A(_0021_),
    .VSS(VGND));
 sg13g2_mux4_1 _1343_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit0.Q ),
    .A0(_1012_),
    .A1(_1014_),
    .A2(_1022_),
    .A3(_0021_),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit1.Q ),
    .X(_0022_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _1344_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit1.Q ),
    .A0(N2END[0]),
    .A1(S2END[0]),
    .A2(E2END[0]),
    .A3(WW4END[3]),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit0.Q ),
    .X(_0023_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _1345_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit6.Q ),
    .A0(A),
    .A1(B),
    .A2(C),
    .A3(E),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit7.Q ),
    .X(_0024_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _1346_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit6.Q ),
    .A0(F),
    .A1(G),
    .A2(H),
    .A3(\Inst_LUT4AB_switch_matrix.M_AB ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit7.Q ),
    .X(_0025_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _1347_ (.Y(_0026_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit8.Q ),
    .A_N(_0025_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1348_ (.B1(_0026_),
    .VDD(VPWR),
    .Y(_0027_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit8.Q ),
    .A2(_0024_));
 sg13g2_mux4_1 _1349_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit7.Q ),
    .A0(N1END[2]),
    .A1(E2END[4]),
    .A2(N2END[4]),
    .A3(E6END[0]),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit6.Q ),
    .X(_0028_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _1350_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit8.Q ),
    .B_N(_0028_),
    .Y(_0029_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _1351_ (.A(S2END[4]),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit6.Q ),
    .Y(_0030_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1352_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1022_),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit6.Q ),
    .Y(_0031_),
    .B1(_0030_));
 sg13g2_nand2_1 _1353_ (.Y(_0032_),
    .A(_1023_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit6.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1354_ (.B1(_0032_),
    .VDD(VPWR),
    .Y(_0033_),
    .VSS(VGND),
    .A1(W2END[4]),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit6.Q ));
 sg13g2_o21ai_1 _1355_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit8.Q ),
    .VDD(VPWR),
    .Y(_0034_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit7.Q ),
    .A2(_0031_));
 sg13g2_a21oi_1 _1356_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit7.Q ),
    .A2(_0033_),
    .Y(_0035_),
    .B1(_0034_));
 sg13g2_nor3_1 _1357_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit9.Q ),
    .B(_0029_),
    .C(_0035_),
    .Y(_0036_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _1358_ (.A2(_0027_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit9.Q ),
    .B1(_0036_),
    .X(_0037_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _1359_ (.VDD(VPWR),
    .Y(\Inst_LUT4AB_switch_matrix.JW2BEG3 ),
    .A(_0037_),
    .VSS(VGND));
 sg13g2_o21ai_1 _1360_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit1.Q ),
    .VDD(VPWR),
    .Y(_0038_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit0.Q ),
    .A2(S2MID[0]));
 sg13g2_a21oi_1 _1361_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit0.Q ),
    .A2(_0037_),
    .Y(_0039_),
    .B1(_0038_));
 sg13g2_nor2b_1 _1362_ (.A(E2MID[0]),
    .B_N(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit0.Q ),
    .Y(_0040_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _1363_ (.A(N2MID[0]),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit0.Q ),
    .Y(_0041_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _1364_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit1.Q ),
    .B(_0040_),
    .C(_0041_),
    .Y(_0042_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _1365_ (.A(_0039_),
    .B(_0042_),
    .Y(_0043_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _1366_ (.A0(N2MID[1]),
    .A1(E2MID[1]),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit0.Q ),
    .X(_0044_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _1367_ (.Y(_0045_),
    .B(S2MID[1]),
    .A_N(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit0.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1368_ (.Y(_0046_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit0.Q ),
    .B(W2MID[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _1369_ (.B(_0045_),
    .C(_0046_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit1.Q ),
    .Y(_0047_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1370_ (.B1(_0047_),
    .VDD(VPWR),
    .Y(_0048_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit1.Q ),
    .A2(_0044_));
 sg13g2_nand2_1 _1371_ (.Y(_0049_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit8.Q ),
    .B(_0048_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1372_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1029_),
    .A2(_0043_),
    .Y(_0050_),
    .B1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit9.Q ));
 sg13g2_o21ai_1 _1373_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit9.Q ),
    .VDD(VPWR),
    .Y(_0051_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit8.Q ),
    .A2(_0023_));
 sg13g2_a21oi_1 _1374_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit8.Q ),
    .A2(_0022_),
    .Y(_0052_),
    .B1(_0051_));
 sg13g2_a21oi_1 _1375_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0049_),
    .A2(_0050_),
    .Y(_0053_),
    .B1(_0052_));
 sg13g2_mux2_1 _1376_ (.A0(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ),
    .A1(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ),
    .S(_1121_),
    .X(_0054_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _1377_ (.A0(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ),
    .A1(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ),
    .S(_1121_),
    .X(_0055_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _1378_ (.A0(_0055_),
    .A1(_0054_),
    .S(_1085_),
    .X(_0056_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _1379_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_1160_),
    .C1(_0053_),
    .B1(_0056_),
    .A1(_1124_),
    .Y(_0057_),
    .A2(_0008_));
 sg13g2_mux2_1 _1380_ (.A0(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ),
    .A1(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ),
    .S(_1121_),
    .X(_0058_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _1381_ (.A0(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ),
    .A1(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ),
    .S(_1121_),
    .X(_0059_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _1382_ (.A0(_0059_),
    .A1(_0058_),
    .S(_1085_),
    .X(_0060_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _1383_ (.Y(_0061_),
    .B(_0060_),
    .A_N(_1160_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _1384_ (.Y(_0062_),
    .B(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ),
    .A_N(_1121_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1385_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ),
    .A2(_1121_),
    .Y(_0063_),
    .B1(_1085_));
 sg13g2_nand2_1 _1386_ (.Y(_0064_),
    .A(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ),
    .B(_1121_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _1387_ (.Y(_0065_),
    .B(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ),
    .A_N(_1121_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _1388_ (.A(_1085_),
    .B(_0065_),
    .X(_0066_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _1389_ (.Y(_0067_),
    .B1(_0064_),
    .B2(_0066_),
    .A2(_0063_),
    .A1(_0062_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _1390_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_1160_),
    .C1(_0052_),
    .B1(_0067_),
    .A1(_0049_),
    .Y(_0068_),
    .A2(_0050_));
 sg13g2_a21oi_1 _1391_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0061_),
    .A2(_0068_),
    .Y(_0069_),
    .B1(_0057_));
 sg13g2_mux2_1 _1392_ (.A0(_0069_),
    .A1(\Inst_LA_LUT4c_frame_config_dffesr.LUT_flop ),
    .S(\Inst_LA_LUT4c_frame_config_dffesr.c_out_mux ),
    .X(A),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1393_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit19.Q ),
    .VDD(VPWR),
    .Y(_0070_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit18.Q ),
    .A2(_0023_));
 sg13g2_a21o_1 _1394_ (.A2(_0022_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit18.Q ),
    .B1(_0070_),
    .X(_0071_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _1395_ (.A0(_0043_),
    .A1(_0048_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit18.Q ),
    .X(_0072_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1396_ (.B1(_0071_),
    .VDD(VPWR),
    .Y(_0073_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit19.Q ),
    .A2(_0072_));
 sg13g2_mux4_1 _1397_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit14.Q ),
    .A0(_1083_),
    .A1(_1084_),
    .A2(_1066_),
    .A3(_1065_),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit15.Q ),
    .X(_0074_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _1398_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit16.Q ),
    .A0(_1157_),
    .A1(_1159_),
    .A2(_1141_),
    .A3(_1140_),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit17.Q ),
    .X(_0075_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _1399_ (.Y(_0076_),
    .B(_0075_),
    .A_N(_0074_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1400_ (.B1(_0073_),
    .VDD(VPWR),
    .Y(_0077_),
    .VSS(VGND),
    .A1(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ),
    .A2(_0076_));
 sg13g2_nor2b_1 _1401_ (.A(_0075_),
    .B_N(_0074_),
    .Y(_0078_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _1402_ (.A(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ),
    .B_N(_0078_),
    .Y(_0079_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _1403_ (.A(_0074_),
    .B(_0075_),
    .X(_0080_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1404_ (.Y(_0081_),
    .A(_0074_),
    .B(_0075_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _1405_ (.A(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ),
    .B(_0081_),
    .Y(_0082_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _1406_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0083_),
    .B(_0075_),
    .A(_0074_));
 sg13g2_nor2_1 _1407_ (.A(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ),
    .B(_0083_),
    .Y(_0084_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or4_1 _1408_ (.A(_0077_),
    .B(_0079_),
    .C(_0082_),
    .D(_0084_),
    .X(_0085_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _1409_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit12.Q ),
    .A0(_1102_),
    .A1(_1103_),
    .A2(_1119_),
    .A3(_1118_),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit13.Q ),
    .X(_0086_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1410_ (.Y(_0087_),
    .A(Ci),
    .B(_1160_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1411_ (.B1(_1085_),
    .VDD(VPWR),
    .Y(_0088_),
    .VSS(VGND),
    .A1(Ci),
    .A2(_1160_));
 sg13g2_nand2_1 _1412_ (.Y(_0089_),
    .A(_0087_),
    .B(_0088_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _1413_ (.A(\Inst_LB_LUT4c_frame_config_dffesr.c_I0mux ),
    .B_N(_0086_),
    .Y(_0090_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1414_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_LB_LUT4c_frame_config_dffesr.c_I0mux ),
    .A2(_0089_),
    .Y(_0091_),
    .B1(_0090_));
 sg13g2_nor2b_1 _1415_ (.A(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ),
    .B_N(_0078_),
    .Y(_0092_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _1416_ (.A(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ),
    .B(_0081_),
    .Y(_0093_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _1417_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0094_),
    .B(_0076_),
    .A(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ));
 sg13g2_o21ai_1 _1418_ (.B1(_0094_),
    .VDD(VPWR),
    .Y(_0095_),
    .VSS(VGND),
    .A1(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ),
    .A2(_0083_));
 sg13g2_or4_1 _1419_ (.A(_0073_),
    .B(_0092_),
    .C(_0093_),
    .D(_0095_),
    .X(_0096_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _1420_ (.A(_0091_),
    .B(_0096_),
    .X(_0097_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1421_ (.B1(_0073_),
    .VDD(VPWR),
    .Y(_0098_),
    .VSS(VGND),
    .A1(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ),
    .A2(_0081_));
 sg13g2_nor2_1 _1422_ (.A(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ),
    .B(_0083_),
    .Y(_0099_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _1423_ (.Y(_0100_),
    .B(_0078_),
    .A_N(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1424_ (.B1(_0100_),
    .VDD(VPWR),
    .Y(_0101_),
    .VSS(VGND),
    .A1(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ),
    .A2(_0076_));
 sg13g2_nor3_1 _1425_ (.A(_0098_),
    .B(_0099_),
    .C(_0101_),
    .Y(_0102_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _1426_ (.A(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ),
    .B(_0076_),
    .Y(_0103_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _1427_ (.A(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ),
    .B(_0081_),
    .Y(_0104_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _1428_ (.Y(_0105_),
    .B(_0078_),
    .A_N(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1429_ (.B1(_0105_),
    .VDD(VPWR),
    .Y(_0106_),
    .VSS(VGND),
    .A1(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ),
    .A2(_0083_));
 sg13g2_nor4_1 _1430_ (.A(_0073_),
    .B(_0103_),
    .C(_0104_),
    .D(_0106_),
    .Y(_0107_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _1431_ (.A(_0091_),
    .B(_0102_),
    .C(_0107_),
    .Y(_0108_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1432_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0085_),
    .A2(_0097_),
    .Y(_0109_),
    .B1(_0108_));
 sg13g2_mux2_1 _1433_ (.A0(_0109_),
    .A1(\Inst_LB_LUT4c_frame_config_dffesr.LUT_flop ),
    .S(\Inst_LB_LUT4c_frame_config_dffesr.c_out_mux ),
    .X(B),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _1434_ (.Y(_0110_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit2.Q ),
    .A_N(\Inst_LUT4AB_switch_matrix.M_AD ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1435_ (.B1(_0110_),
    .VDD(VPWR),
    .Y(_0111_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit2.Q ),
    .A2(H));
 sg13g2_mux2_1 _1436_ (.A0(F),
    .A1(G),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit2.Q ),
    .X(_0112_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1437_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit4.Q ),
    .VDD(VPWR),
    .Y(_0113_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit3.Q ),
    .A2(_0112_));
 sg13g2_a21oi_1 _1438_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit3.Q ),
    .A2(_0111_),
    .Y(_0114_),
    .B1(_0113_));
 sg13g2_nand2b_1 _1439_ (.Y(_0115_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit2.Q ),
    .A_N(E),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1440_ (.B1(_0115_),
    .VDD(VPWR),
    .Y(_0116_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit2.Q ),
    .A2(D));
 sg13g2_mux2_1 _1441_ (.A0(A),
    .A1(B),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit2.Q ),
    .X(_0117_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1442_ (.B1(_1032_),
    .VDD(VPWR),
    .Y(_0118_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit3.Q ),
    .A2(_0117_));
 sg13g2_a21oi_1 _1443_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit3.Q ),
    .A2(_0116_),
    .Y(_0119_),
    .B1(_0118_));
 sg13g2_nor3_1 _1444_ (.A(_1033_),
    .B(_0114_),
    .C(_0119_),
    .Y(_0120_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _1445_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit3.Q ),
    .A0(N1END[1]),
    .A1(N4END[3]),
    .A2(N2END[3]),
    .A3(E2END[3]),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit2.Q ),
    .X(_0121_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1446_ (.Y(_0122_),
    .A(_1032_),
    .B(_0121_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _1447_ (.Y(_0123_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit2.Q ),
    .A_N(W6END[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1448_ (.B1(_0123_),
    .VDD(VPWR),
    .Y(_0124_),
    .VSS(VGND),
    .A1(W2END[3]),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit2.Q ));
 sg13g2_mux2_1 _1449_ (.A0(E6END[1]),
    .A1(S2END[3]),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit2.Q ),
    .X(_0125_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1450_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit4.Q ),
    .VDD(VPWR),
    .Y(_0126_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit3.Q ),
    .A2(_0125_));
 sg13g2_a21oi_1 _1451_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit3.Q ),
    .A2(_0124_),
    .Y(_0127_),
    .B1(_0126_));
 sg13g2_nor2_1 _1452_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit5.Q ),
    .B(_0127_),
    .Y(_0128_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1453_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0122_),
    .A2(_0128_),
    .Y(\Inst_LUT4AB_switch_matrix.E2BEG2 ),
    .B1(_0120_));
 sg13g2_mux4_1 _1454_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit4.Q ),
    .A0(N4END[2]),
    .A1(E2END[2]),
    .A2(W2END[7]),
    .A3(\Inst_LUT4AB_switch_matrix.E2BEG2 ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit5.Q ),
    .X(_0129_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _1455_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit4.Q ),
    .A0(N2END[2]),
    .A1(E2END[2]),
    .A2(S2END[2]),
    .A3(WW4END[2]),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit5.Q ),
    .X(_0130_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _1456_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit10.Q ),
    .A0(A),
    .A1(B),
    .A2(C),
    .A3(D),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit11.Q ),
    .X(_0131_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _1457_ (.Y(_0132_),
    .B(_0131_),
    .A_N(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit12.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _1458_ (.A0(F),
    .A1(G),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit10.Q ),
    .X(_0133_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _1459_ (.Y(_0134_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit10.Q ),
    .A_N(\Inst_LUT4AB_switch_matrix.M_EF ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1460_ (.B1(_0134_),
    .VDD(VPWR),
    .Y(_0135_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit10.Q ),
    .A2(H));
 sg13g2_o21ai_1 _1461_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit12.Q ),
    .VDD(VPWR),
    .Y(_0136_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit11.Q ),
    .A2(_0133_));
 sg13g2_a21oi_1 _1462_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit11.Q ),
    .A2(_0135_),
    .Y(_0137_),
    .B1(_0136_));
 sg13g2_nor2b_1 _1463_ (.A(_0137_),
    .B_N(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit13.Q ),
    .Y(_0138_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _1464_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit10.Q ),
    .A0(N1END[1]),
    .A1(N2END[5]),
    .A2(E1END[1]),
    .A3(E2END[5]),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit11.Q ),
    .X(_0139_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _1465_ (.Y(_0140_),
    .B(_0139_),
    .A_N(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit12.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _1466_ (.Y(_0141_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit10.Q ),
    .A_N(W1END[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1467_ (.B1(_0141_),
    .VDD(VPWR),
    .Y(_0142_),
    .VSS(VGND),
    .A1(S2END[5]),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit10.Q ));
 sg13g2_mux2_1 _1468_ (.A0(S1END[1]),
    .A1(S1END[3]),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit10.Q ),
    .X(_0143_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1469_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit12.Q ),
    .VDD(VPWR),
    .Y(_0144_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit11.Q ),
    .A2(_0143_));
 sg13g2_a21oi_1 _1470_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit11.Q ),
    .A2(_0142_),
    .Y(_0145_),
    .B1(_0144_));
 sg13g2_nor2_1 _1471_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit13.Q ),
    .B(_0145_),
    .Y(_0146_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _1472_ (.Y(\Inst_LUT4AB_switch_matrix.E2BEG4 ),
    .B1(_0140_),
    .B2(_0146_),
    .A2(_0138_),
    .A1(_0132_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _1473_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit5.Q ),
    .A0(N2MID[2]),
    .A1(W2MID[2]),
    .A2(E2MID[2]),
    .A3(\Inst_LUT4AB_switch_matrix.E2BEG4 ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit4.Q ),
    .X(_0147_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _1474_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit4.Q ),
    .A0(N2MID[3]),
    .A1(E2MID[3]),
    .A2(S2MID[3]),
    .A3(W2MID[3]),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit5.Q ),
    .X(_0148_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _1475_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit2.Q ),
    .A0(_0147_),
    .A1(_0148_),
    .A2(_0130_),
    .A3(_0129_),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit3.Q ),
    .X(_0149_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _1476_ (.Y(_0150_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit2.Q ),
    .A_N(E),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1477_ (.B1(_0150_),
    .VDD(VPWR),
    .Y(_0151_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit2.Q ),
    .A2(D));
 sg13g2_mux2_1 _1478_ (.A0(A),
    .A1(B),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit2.Q ),
    .X(_0152_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1479_ (.B1(_1037_),
    .VDD(VPWR),
    .Y(_0153_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit3.Q ),
    .A2(_0152_));
 sg13g2_a21oi_1 _1480_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit3.Q ),
    .A2(_0151_),
    .Y(_0154_),
    .B1(_0153_));
 sg13g2_nor2_1 _1481_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit2.Q ),
    .B(F),
    .Y(_0155_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1482_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit2.Q ),
    .A2(_1051_),
    .Y(_0156_),
    .B1(_0155_));
 sg13g2_nand2b_1 _1483_ (.Y(_0157_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit2.Q ),
    .A_N(\Inst_LUT4AB_switch_matrix.M_AB ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1484_ (.B1(_0157_),
    .VDD(VPWR),
    .Y(_0158_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit2.Q ),
    .A2(H));
 sg13g2_a21oi_1 _1485_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit3.Q ),
    .A2(_0158_),
    .Y(_0159_),
    .B1(_1037_));
 sg13g2_o21ai_1 _1486_ (.B1(_0159_),
    .VDD(VPWR),
    .Y(_0160_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit3.Q ),
    .A2(_0156_));
 sg13g2_nor2_1 _1487_ (.A(_1038_),
    .B(_0154_),
    .Y(_0161_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _1488_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit2.Q ),
    .A0(NN4END[3]),
    .A1(E1END[1]),
    .A2(E2END[3]),
    .A3(E6END[1]),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit3.Q ),
    .X(_0162_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _1489_ (.Y(_0163_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit2.Q ),
    .A_N(W6END[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1490_ (.B1(_0163_),
    .VDD(VPWR),
    .Y(_0164_),
    .VSS(VGND),
    .A1(W2END[3]),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit2.Q ));
 sg13g2_mux2_1 _1491_ (.A0(S2END[3]),
    .A1(S4END[3]),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit2.Q ),
    .X(_0165_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1492_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit4.Q ),
    .VDD(VPWR),
    .Y(_0166_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit3.Q ),
    .A2(_0165_));
 sg13g2_a21oi_1 _1493_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit3.Q ),
    .A2(_0164_),
    .Y(_0167_),
    .B1(_0166_));
 sg13g2_a21oi_1 _1494_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1037_),
    .A2(_0162_),
    .Y(_0168_),
    .B1(_0167_));
 sg13g2_a22oi_1 _1495_ (.Y(\Inst_LUT4AB_switch_matrix.JS2BEG2 ),
    .B1(_0168_),
    .B2(_1038_),
    .A2(_0161_),
    .A1(_0160_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _1496_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit6.Q ),
    .A0(NN4END[1]),
    .A1(EE4END[1]),
    .A2(S4END[1]),
    .A3(\Inst_LUT4AB_switch_matrix.JS2BEG2 ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit7.Q ),
    .X(_0169_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _1497_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit6.Q ),
    .A0(N2END[4]),
    .A1(E2END[4]),
    .A2(SS4END[2]),
    .A3(W2END[4]),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit7.Q ),
    .X(_0170_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _1498_ (.VDD(VPWR),
    .Y(_0171_),
    .A(_0170_),
    .VSS(VGND));
 sg13g2_nand2b_1 _1499_ (.Y(_0172_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit10.Q ),
    .A_N(D),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1500_ (.B1(_0172_),
    .VDD(VPWR),
    .Y(_0173_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit10.Q ),
    .A2(C));
 sg13g2_mux2_1 _1501_ (.A0(A),
    .A1(B),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit10.Q ),
    .X(_0174_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1502_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit11.Q ),
    .A2(_0173_),
    .Y(_0175_),
    .B1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit12.Q ));
 sg13g2_o21ai_1 _1503_ (.B1(_0175_),
    .VDD(VPWR),
    .Y(_0176_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit11.Q ),
    .A2(_0174_));
 sg13g2_mux2_1 _1504_ (.A0(F),
    .A1(G),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit10.Q ),
    .X(_0177_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _1505_ (.Y(_0178_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit10.Q ),
    .A_N(\Inst_LUT4AB_switch_matrix.M_AH ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1506_ (.B1(_0178_),
    .VDD(VPWR),
    .Y(_0179_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit10.Q ),
    .A2(H));
 sg13g2_o21ai_1 _1507_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit12.Q ),
    .VDD(VPWR),
    .Y(_0180_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit11.Q ),
    .A2(_0177_));
 sg13g2_a21oi_1 _1508_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit11.Q ),
    .A2(_0179_),
    .Y(_0181_),
    .B1(_0180_));
 sg13g2_nor2_1 _1509_ (.A(_1035_),
    .B(_0181_),
    .Y(_0182_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _1510_ (.Y(_0183_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit10.Q ),
    .A_N(S2END[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1511_ (.B1(_0183_),
    .VDD(VPWR),
    .Y(_0184_),
    .VSS(VGND),
    .A1(S1END[1]),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit10.Q ));
 sg13g2_nand2b_1 _1512_ (.Y(_0185_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit10.Q ),
    .A_N(W1END[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1513_ (.B1(_0185_),
    .VDD(VPWR),
    .Y(_0186_),
    .VSS(VGND),
    .A1(W1END[1]),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit10.Q ));
 sg13g2_nand2b_1 _1514_ (.Y(_0187_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit10.Q ),
    .A_N(E2END[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1515_ (.B1(_0187_),
    .VDD(VPWR),
    .Y(_0188_),
    .VSS(VGND),
    .A1(E1END[1]),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit10.Q ));
 sg13g2_nand2b_1 _1516_ (.Y(_0189_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit10.Q ),
    .A_N(N2END[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1517_ (.B1(_0189_),
    .VDD(VPWR),
    .Y(_0190_),
    .VSS(VGND),
    .A1(N1END[1]),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit10.Q ));
 sg13g2_mux4_1 _1518_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit11.Q ),
    .A0(_0190_),
    .A1(_0188_),
    .A2(_0184_),
    .A3(_0186_),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit12.Q ),
    .X(_0191_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _1519_ (.Y(\Inst_LUT4AB_switch_matrix.JS2BEG4 ),
    .B1(_0191_),
    .B2(_1035_),
    .A2(_0182_),
    .A1(_0176_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1520_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit7.Q ),
    .VDD(VPWR),
    .Y(_0192_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit6.Q ),
    .A2(_1034_));
 sg13g2_a21o_1 _1521_ (.A2(\Inst_LUT4AB_switch_matrix.JS2BEG4 ),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit6.Q ),
    .B1(_0192_),
    .X(_0193_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1522_ (.Y(_0194_),
    .A(E2MID[4]),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit6.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1523_ (.B1(_0194_),
    .VDD(VPWR),
    .Y(_0195_),
    .VSS(VGND),
    .A1(_1021_),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit6.Q ));
 sg13g2_o21ai_1 _1524_ (.B1(_0193_),
    .VDD(VPWR),
    .Y(_0196_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit7.Q ),
    .A2(_0195_));
 sg13g2_mux4_1 _1525_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit6.Q ),
    .A0(N2MID[4]),
    .A1(E2MID[4]),
    .A2(S2MID[4]),
    .A3(\Inst_LUT4AB_switch_matrix.JS2BEG4 ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit7.Q ),
    .X(_0197_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _1526_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit6.Q ),
    .A0(N2MID[5]),
    .A1(E2MID[5]),
    .A2(S2MID[5]),
    .A3(W2MID[5]),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit7.Q ),
    .X(_0198_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _1527_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit4.Q ),
    .A0(_0197_),
    .A1(_0198_),
    .A2(_0170_),
    .A3(_0169_),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit5.Q ),
    .X(_0199_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _1528_ (.A(_0149_),
    .B(_0199_),
    .Y(_0200_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1529_ (.Y(_0201_),
    .A(_0149_),
    .B(_0199_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _1530_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit24.Q ),
    .A0(_0147_),
    .A1(_0148_),
    .A2(_0130_),
    .A3(_0129_),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit25.Q ),
    .X(_0202_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _1531_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit26.Q ),
    .A0(_0197_),
    .A1(_0198_),
    .A2(_0170_),
    .A3(_0169_),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit27.Q ),
    .X(_0203_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _1532_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0204_),
    .B(_0203_),
    .A(_0202_));
 sg13g2_nand2_1 _1533_ (.Y(_0205_),
    .A(_0202_),
    .B(_0203_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _1534_ (.VDD(VPWR),
    .Y(_0206_),
    .A(_0205_),
    .VSS(VGND));
 sg13g2_a21o_1 _1535_ (.A2(_0089_),
    .A1(_0083_),
    .B1(_0080_),
    .X(_0207_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1536_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0204_),
    .A2(_0207_),
    .Y(_0208_),
    .B1(_0206_));
 sg13g2_o21ai_1 _1537_ (.B1(_0201_),
    .VDD(VPWR),
    .Y(_0209_),
    .VSS(VGND),
    .A1(_0200_),
    .A2(_0208_));
 sg13g2_o21ai_1 _1538_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit15.Q ),
    .VDD(VPWR),
    .Y(_0210_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit14.Q ),
    .A2(_1052_));
 sg13g2_a21oi_1 _1539_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit14.Q ),
    .A2(\Inst_LUT4AB_switch_matrix.M_AD ),
    .Y(_0211_),
    .B1(_0210_));
 sg13g2_nor2_1 _1540_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit14.Q ),
    .B(E),
    .Y(_0212_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1541_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit14.Q ),
    .A2(_1051_),
    .Y(_0213_),
    .B1(_0212_));
 sg13g2_o21ai_1 _1542_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit16.Q ),
    .VDD(VPWR),
    .Y(_0214_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit15.Q ),
    .A2(_0213_));
 sg13g2_nor2_1 _1543_ (.A(_0211_),
    .B(_0214_),
    .Y(_0215_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _1544_ (.Y(_0216_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit14.Q ),
    .A_N(D),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1545_ (.B1(_0216_),
    .VDD(VPWR),
    .Y(_0217_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit14.Q ),
    .A2(C));
 sg13g2_mux2_1 _1546_ (.A0(A),
    .A1(B),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit14.Q ),
    .X(_0218_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1547_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit15.Q ),
    .A2(_0217_),
    .Y(_0219_),
    .B1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit16.Q ));
 sg13g2_o21ai_1 _1548_ (.B1(_0219_),
    .VDD(VPWR),
    .Y(_0220_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit15.Q ),
    .A2(_0218_));
 sg13g2_nand2_1 _1549_ (.Y(_0221_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit17.Q ),
    .B(_0220_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _1550_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit14.Q ),
    .A0(N1END[2]),
    .A1(N2END[6]),
    .A2(E1END[2]),
    .A3(E2END[6]),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit15.Q ),
    .X(_0222_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _1551_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit16.Q ),
    .B_N(_0222_),
    .Y(_0223_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _1552_ (.Y(_0224_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit14.Q ),
    .A_N(W1END[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1553_ (.B1(_0224_),
    .VDD(VPWR),
    .Y(_0225_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit14.Q ),
    .A2(W1END[0]));
 sg13g2_mux2_1 _1554_ (.A0(S1END[2]),
    .A1(S2END[6]),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit14.Q ),
    .X(_0226_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1555_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit16.Q ),
    .VDD(VPWR),
    .Y(_0227_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit15.Q ),
    .A2(_0226_));
 sg13g2_a21oi_1 _1556_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit15.Q ),
    .A2(_0225_),
    .Y(_0228_),
    .B1(_0227_));
 sg13g2_or3_1 _1557_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit17.Q ),
    .B(_0223_),
    .C(_0228_),
    .X(_0229_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1558_ (.B1(_0229_),
    .VDD(VPWR),
    .Y(_0230_),
    .VSS(VGND),
    .A1(_0215_),
    .A2(_0221_));
 sg13g2_inv_1 _1559_ (.VDD(VPWR),
    .Y(\Inst_LUT4AB_switch_matrix.JN2BEG5 ),
    .A(_0230_),
    .VSS(VGND));
 sg13g2_o21ai_1 _1560_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit11.Q ),
    .VDD(VPWR),
    .Y(_0231_),
    .VSS(VGND),
    .A1(W2MID[6]),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit10.Q ));
 sg13g2_a21oi_1 _1561_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit10.Q ),
    .A2(_0230_),
    .Y(_0232_),
    .B1(_0231_));
 sg13g2_nor2b_1 _1562_ (.A(E2MID[6]),
    .B_N(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit10.Q ),
    .Y(_0233_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _1563_ (.A(N2MID[6]),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit10.Q ),
    .Y(_0234_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _1564_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit11.Q ),
    .B(_0233_),
    .C(_0234_),
    .Y(_0235_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _1565_ (.A(_0232_),
    .B(_0235_),
    .Y(_0236_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _1566_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit10.Q ),
    .A0(N2MID[7]),
    .A1(E2MID[7]),
    .A2(S2MID[7]),
    .A3(W2MID[7]),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit11.Q ),
    .X(_0237_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _1567_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit11.Q ),
    .A0(N4END[3]),
    .A1(W2END[3]),
    .A2(E2END[3]),
    .A3(\Inst_LUT4AB_switch_matrix.JN2BEG3 ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit10.Q ),
    .X(_0238_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _1568_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit11.Q ),
    .A0(N2END[7]),
    .A1(S2END[7]),
    .A2(EE4END[2]),
    .A3(W2END[7]),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit10.Q ),
    .X(_0239_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1569_ (.Y(_0240_),
    .A(\Inst_LE_LUT4c_frame_config_dffesr.c_I0mux ),
    .B(_0209_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1570_ (.Y(_0241_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit10.Q ),
    .B(_0237_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1571_ (.B1(_0241_),
    .VDD(VPWR),
    .Y(_0242_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit10.Q ),
    .A2(_0236_));
 sg13g2_nor2b_1 _1572_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit10.Q ),
    .B_N(_0239_),
    .Y(_0243_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1573_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit10.Q ),
    .A2(_0238_),
    .Y(_0244_),
    .B1(_0243_));
 sg13g2_a21oi_1 _1574_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit11.Q ),
    .A2(_0244_),
    .Y(_0245_),
    .B1(\Inst_LE_LUT4c_frame_config_dffesr.c_I0mux ));
 sg13g2_o21ai_1 _1575_ (.B1(_0245_),
    .VDD(VPWR),
    .Y(_0246_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit11.Q ),
    .A2(_0242_));
 sg13g2_nand2_1 _1576_ (.Y(_0247_),
    .A(_0240_),
    .B(_0246_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _1577_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit14.Q ),
    .A0(N4END[1]),
    .A1(SS4END[1]),
    .A2(W2END[4]),
    .A3(\Inst_LUT4AB_switch_matrix.JS2BEG3 ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit15.Q ),
    .X(_0248_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _1578_ (.A0(N2END[5]),
    .A1(E2END[5]),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit14.Q ),
    .X(_0249_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _1579_ (.Y(_0250_),
    .B(SS4END[1]),
    .A_N(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit14.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1580_ (.Y(_0251_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit14.Q ),
    .B(W2END[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _1581_ (.B(_0250_),
    .C(_0251_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit15.Q ),
    .Y(_0252_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1582_ (.B1(_0252_),
    .VDD(VPWR),
    .Y(_0253_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit15.Q ),
    .A2(_0249_));
 sg13g2_o21ai_1 _1583_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit15.Q ),
    .VDD(VPWR),
    .Y(_0254_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit14.Q ),
    .A2(_0253_));
 sg13g2_a21oi_1 _1584_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit14.Q ),
    .A2(_0248_),
    .Y(_0255_),
    .B1(_0254_));
 sg13g2_mux4_1 _1585_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit14.Q ),
    .A0(A),
    .A1(B),
    .A2(C),
    .A3(D),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit15.Q ),
    .X(_0256_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _1586_ (.A(_1042_),
    .B(_0256_),
    .X(_0257_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _1587_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit14.Q ),
    .B(E),
    .Y(_0258_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1588_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit14.Q ),
    .A2(_1051_),
    .Y(_0259_),
    .B1(_0258_));
 sg13g2_mux2_1 _1589_ (.A0(H),
    .A1(\Inst_LUT4AB_switch_matrix.M_EF ),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit14.Q ),
    .X(_0260_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _1590_ (.A(_0260_),
    .B_N(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit15.Q ),
    .Y(_0261_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1591_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit16.Q ),
    .VDD(VPWR),
    .Y(_0262_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit15.Q ),
    .A2(_0259_));
 sg13g2_o21ai_1 _1592_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit17.Q ),
    .VDD(VPWR),
    .Y(_0263_),
    .VSS(VGND),
    .A1(_0261_),
    .A2(_0262_));
 sg13g2_o21ai_1 _1593_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit15.Q ),
    .VDD(VPWR),
    .Y(_0264_),
    .VSS(VGND),
    .A1(_1013_),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit14.Q ));
 sg13g2_a21oi_1 _1594_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(E2END[6]),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit14.Q ),
    .Y(_0265_),
    .B1(_0264_));
 sg13g2_mux2_1 _1595_ (.A0(N1END[2]),
    .A1(N2END[6]),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit14.Q ),
    .X(_0266_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1596_ (.B1(_1042_),
    .VDD(VPWR),
    .Y(_0267_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit15.Q ),
    .A2(_0266_));
 sg13g2_nor2_1 _1597_ (.A(_0265_),
    .B(_0267_),
    .Y(_0268_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _1598_ (.Y(_0269_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit14.Q ),
    .A_N(W1END[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1599_ (.B1(_0269_),
    .VDD(VPWR),
    .Y(_0270_),
    .VSS(VGND),
    .A1(W1END[0]),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit14.Q ));
 sg13g2_mux2_1 _1600_ (.A0(S1END[2]),
    .A1(S2END[6]),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit14.Q ),
    .X(_0271_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1601_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit16.Q ),
    .VDD(VPWR),
    .Y(_0272_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit15.Q ),
    .A2(_0271_));
 sg13g2_a21oi_1 _1602_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit15.Q ),
    .A2(_0270_),
    .Y(_0273_),
    .B1(_0272_));
 sg13g2_or3_1 _1603_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit17.Q ),
    .B(_0268_),
    .C(_0273_),
    .X(_0274_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1604_ (.B1(_0274_),
    .VDD(VPWR),
    .Y(_0275_),
    .VSS(VGND),
    .A1(_0257_),
    .A2(_0263_));
 sg13g2_inv_1 _1605_ (.VDD(VPWR),
    .Y(\Inst_LUT4AB_switch_matrix.JS2BEG5 ),
    .A(_0275_),
    .VSS(VGND));
 sg13g2_mux4_1 _1606_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit15.Q ),
    .A0(_1021_),
    .A1(_1026_),
    .A2(_1034_),
    .A3(_0275_),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit14.Q ),
    .X(_0276_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _1607_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit14.Q ),
    .A0(N2MID[5]),
    .A1(E2MID[5]),
    .A2(S2MID[5]),
    .A3(W2MID[5]),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit15.Q ),
    .X(_0277_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1608_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit14.Q ),
    .A2(_0277_),
    .Y(_0278_),
    .B1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit15.Q ));
 sg13g2_o21ai_1 _1609_ (.B1(_0278_),
    .VDD(VPWR),
    .Y(_0279_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit14.Q ),
    .A2(_0276_));
 sg13g2_nor2b_1 _1610_ (.A(_0255_),
    .B_N(_0279_),
    .Y(_0280_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _1611_ (.VDD(VPWR),
    .Y(_0281_),
    .A(_0280_),
    .VSS(VGND));
 sg13g2_mux2_1 _1612_ (.A0(NN4END[2]),
    .A1(E2END[2]),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit12.Q ),
    .X(_0282_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _1613_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit12.Q ),
    .B_N(S4END[2]),
    .Y(_0283_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1614_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit12.Q ),
    .A2(\Inst_LUT4AB_switch_matrix.E2BEG3 ),
    .Y(_0284_),
    .B1(_0283_));
 sg13g2_nand2_1 _1615_ (.Y(_0285_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit13.Q ),
    .B(_0284_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1616_ (.B1(_0285_),
    .VDD(VPWR),
    .Y(_0286_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit13.Q ),
    .A2(_0282_));
 sg13g2_o21ai_1 _1617_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit13.Q ),
    .VDD(VPWR),
    .Y(_0287_),
    .VSS(VGND),
    .A1(S2END[3]),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit12.Q ));
 sg13g2_a21oi_1 _1618_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1030_),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit12.Q ),
    .Y(_0288_),
    .B1(_0287_));
 sg13g2_mux2_1 _1619_ (.A0(N2END[3]),
    .A1(E2END[3]),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit12.Q ),
    .X(_0289_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1620_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1041_),
    .A2(_0289_),
    .Y(_0290_),
    .B1(_0288_));
 sg13g2_mux4_1 _1621_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit14.Q ),
    .A0(A),
    .A1(B),
    .A2(C),
    .A3(D),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit15.Q ),
    .X(_0291_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _1622_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit14.Q ),
    .A0(E),
    .A1(G),
    .A2(H),
    .A3(\Inst_LUT4AB_switch_matrix.M_AB ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit15.Q ),
    .X(_0292_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _1623_ (.Y(_0293_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit16.Q ),
    .A_N(_0292_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1624_ (.B1(_0293_),
    .VDD(VPWR),
    .Y(_0294_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit16.Q ),
    .A2(_0291_));
 sg13g2_mux4_1 _1625_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit14.Q ),
    .A0(N1END[2]),
    .A1(N2END[6]),
    .A2(E1END[2]),
    .A3(E2END[6]),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit15.Q ),
    .X(_0295_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _1626_ (.Y(_0296_),
    .B(_0295_),
    .A_N(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit16.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _1627_ (.A0(S1END[0]),
    .A1(S1END[2]),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit14.Q ),
    .X(_0297_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _1628_ (.Y(_0298_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit14.Q ),
    .A_N(W1END[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1629_ (.B1(_0298_),
    .VDD(VPWR),
    .Y(_0299_),
    .VSS(VGND),
    .A1(S2END[6]),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit14.Q ));
 sg13g2_o21ai_1 _1630_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit16.Q ),
    .VDD(VPWR),
    .Y(_0300_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit15.Q ),
    .A2(_0297_));
 sg13g2_a21oi_1 _1631_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit15.Q ),
    .A2(_0299_),
    .Y(_0301_),
    .B1(_0300_));
 sg13g2_nor2_1 _1632_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit17.Q ),
    .B(_0301_),
    .Y(_0302_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _1633_ (.Y(\Inst_LUT4AB_switch_matrix.E2BEG5 ),
    .B1(_0296_),
    .B2(_0302_),
    .A2(_0294_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit17.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _1634_ (.A0(N2MID[2]),
    .A1(E2MID[2]),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit12.Q ),
    .X(_0303_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1635_ (.Y(_0304_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit12.Q ),
    .B(\Inst_LUT4AB_switch_matrix.E2BEG5 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _1636_ (.Y(_0305_),
    .B(S2MID[2]),
    .A_N(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit12.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _1637_ (.B(_0304_),
    .C(_0305_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit13.Q ),
    .Y(_0306_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1638_ (.B1(_0306_),
    .VDD(VPWR),
    .Y(_0307_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit13.Q ),
    .A2(_0303_));
 sg13g2_mux4_1 _1639_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit12.Q ),
    .A0(N2MID[3]),
    .A1(E2MID[3]),
    .A2(S2MID[3]),
    .A3(W2MID[3]),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit13.Q ),
    .X(_0308_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _1640_ (.VDD(VPWR),
    .Y(_0309_),
    .A(_0308_),
    .VSS(VGND));
 sg13g2_mux4_1 _1641_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit12.Q ),
    .A0(_0307_),
    .A1(_0309_),
    .A2(_0290_),
    .A3(_0286_),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit13.Q ),
    .X(_0310_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1642_ (.Y(_0311_),
    .A(_0281_),
    .B(_0310_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _1643_ (.A(_0281_),
    .B(_0310_),
    .Y(_0312_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _1644_ (.S0(_0280_),
    .A0(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ),
    .A1(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ),
    .A2(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ),
    .A3(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ),
    .S1(_0310_),
    .X(_0313_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _1645_ (.A(_0313_),
    .B_N(_0247_),
    .Y(_0314_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _1646_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit17.Q ),
    .A0(_1040_),
    .A1(_1030_),
    .A2(_1022_),
    .A3(_0037_),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit16.Q ),
    .X(_0315_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _1647_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit16.Q ),
    .A0(NN4END[2]),
    .A1(E2END[1]),
    .A2(S2END[1]),
    .A3(W2END[1]),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit17.Q ),
    .X(_0316_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _1648_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit14.Q ),
    .A0(A),
    .A1(B),
    .A2(C),
    .A3(D),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit15.Q ),
    .X(_0317_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _1649_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit14.Q ),
    .A0(E),
    .A1(G),
    .A2(H),
    .A3(\Inst_LUT4AB_switch_matrix.M_AH ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit15.Q ),
    .X(_0318_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _1650_ (.Y(_0319_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit16.Q ),
    .A_N(_0318_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1651_ (.B1(_0319_),
    .VDD(VPWR),
    .Y(_0320_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit16.Q ),
    .A2(_0317_));
 sg13g2_mux4_1 _1652_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit14.Q ),
    .A0(N1END[2]),
    .A1(N2END[6]),
    .A2(E1END[2]),
    .A3(E2END[6]),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit15.Q ),
    .X(_0321_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _1653_ (.Y(_0322_),
    .B(_0321_),
    .A_N(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit16.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _1654_ (.Y(_0323_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit14.Q ),
    .A_N(W1END[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1655_ (.B1(_0323_),
    .VDD(VPWR),
    .Y(_0324_),
    .VSS(VGND),
    .A1(S2END[6]),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit14.Q ));
 sg13g2_mux2_1 _1656_ (.A0(S1END[0]),
    .A1(S1END[2]),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit14.Q ),
    .X(_0325_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1657_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit16.Q ),
    .VDD(VPWR),
    .Y(_0326_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit15.Q ),
    .A2(_0325_));
 sg13g2_a21oi_1 _1658_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit15.Q ),
    .A2(_0324_),
    .Y(_0327_),
    .B1(_0326_));
 sg13g2_nor2_1 _1659_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit17.Q ),
    .B(_0327_),
    .Y(_0328_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _1660_ (.Y(\Inst_LUT4AB_switch_matrix.JW2BEG5 ),
    .B1(_0322_),
    .B2(_0328_),
    .A2(_0320_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit17.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _1661_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit16.Q ),
    .A0(E2MID[0]),
    .A1(S2MID[0]),
    .A2(W2MID[0]),
    .A3(\Inst_LUT4AB_switch_matrix.JW2BEG5 ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit17.Q ),
    .X(_0329_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _1662_ (.A0(N2MID[1]),
    .A1(E2MID[1]),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit16.Q ),
    .X(_0330_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _1663_ (.Y(_0331_),
    .B(S2MID[1]),
    .A_N(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit16.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1664_ (.Y(_0332_),
    .A(W2MID[1]),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit16.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _1665_ (.B(_0331_),
    .C(_0332_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit17.Q ),
    .Y(_0333_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1666_ (.B1(_0333_),
    .VDD(VPWR),
    .Y(_0334_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit17.Q ),
    .A2(_0330_));
 sg13g2_a21oi_1 _1667_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit16.Q ),
    .A2(_0315_),
    .Y(_0335_),
    .B1(_1043_));
 sg13g2_o21ai_1 _1668_ (.B1(_0335_),
    .VDD(VPWR),
    .Y(_0336_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit16.Q ),
    .A2(_0316_));
 sg13g2_nand2_1 _1669_ (.Y(_0337_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit16.Q ),
    .B(_0334_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1670_ (.B1(_0337_),
    .VDD(VPWR),
    .Y(_0338_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit16.Q ),
    .A2(_0329_));
 sg13g2_o21ai_1 _1671_ (.B1(_0336_),
    .VDD(VPWR),
    .Y(_0339_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit17.Q ),
    .A2(_0338_));
 sg13g2_mux4_1 _1672_ (.S0(_0280_),
    .A0(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ),
    .A1(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ),
    .A2(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ),
    .A3(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ),
    .S1(_0310_),
    .X(_0340_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _1673_ (.A(_0247_),
    .B(_0340_),
    .Y(_0341_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _1674_ (.A(_0314_),
    .B(_0339_),
    .C(_0341_),
    .Y(_0342_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _1675_ (.S0(_0280_),
    .A0(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ),
    .A1(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ),
    .A2(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ),
    .A3(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ),
    .S1(_0310_),
    .X(_0343_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _1676_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0344_),
    .B(_0343_),
    .A(_0247_));
 sg13g2_mux4_1 _1677_ (.S0(_0280_),
    .A0(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ),
    .A1(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ),
    .A2(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ),
    .A3(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ),
    .S1(_0310_),
    .X(_0345_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _1678_ (.Y(_0346_),
    .B(_0247_),
    .A_N(_0345_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _1679_ (.B(_0344_),
    .C(_0346_),
    .A(_0339_),
    .Y(_0347_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _1680_ (.Y(_0348_),
    .B(_0347_),
    .A_N(_0342_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _1681_ (.A0(_0348_),
    .A1(\Inst_LE_LUT4c_frame_config_dffesr.LUT_flop ),
    .S(\Inst_LE_LUT4c_frame_config_dffesr.c_out_mux ),
    .X(E),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _1682_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit2.Q ),
    .A0(A),
    .A1(B),
    .A2(D),
    .A3(E),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit3.Q ),
    .X(_0349_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _1683_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit2.Q ),
    .A0(F),
    .A1(G),
    .A2(H),
    .A3(\Inst_LUT4AB_switch_matrix.M_AH ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit3.Q ),
    .X(_0350_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _1684_ (.Y(_0351_),
    .B(_1031_),
    .A_N(_0349_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1685_ (.B1(_0351_),
    .VDD(VPWR),
    .Y(_0352_),
    .VSS(VGND),
    .A1(_1031_),
    .A2(_0350_));
 sg13g2_mux4_1 _1686_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit2.Q ),
    .A0(N2END[3]),
    .A1(N4END[3]),
    .A2(E1END[1]),
    .A3(E2END[3]),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit3.Q ),
    .X(_0353_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1687_ (.Y(_0354_),
    .A(_1031_),
    .B(_0353_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _1688_ (.A0(E6END[1]),
    .A1(S2END[3]),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit2.Q ),
    .X(_0355_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _1689_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0356_),
    .B(_0355_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit3.Q ));
 sg13g2_nand2_1 _1690_ (.Y(_0357_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit2.Q ),
    .B(_1030_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1691_ (.B1(_0357_),
    .VDD(VPWR),
    .Y(_0358_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit2.Q ),
    .A2(W2END[3]));
 sg13g2_a21oi_1 _1692_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit3.Q ),
    .A2(_0358_),
    .Y(_0359_),
    .B1(_1031_));
 sg13g2_a21oi_1 _1693_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0356_),
    .A2(_0359_),
    .Y(_0360_),
    .B1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit5.Q ));
 sg13g2_a22oi_1 _1694_ (.Y(\Inst_LUT4AB_switch_matrix.JN2BEG2 ),
    .B1(_0354_),
    .B2(_0360_),
    .A2(_0352_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit5.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _1695_ (.A0(E2END[3]),
    .A1(SS4END[3]),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit2.Q ),
    .X(_0361_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _1696_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit3.Q ),
    .B(_0361_),
    .Y(_0362_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1697_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit3.Q ),
    .VDD(VPWR),
    .Y(_0363_),
    .VSS(VGND),
    .A1(_1023_),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit2.Q ));
 sg13g2_a21oi_1 _1698_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit2.Q ),
    .A2(\Inst_LUT4AB_switch_matrix.JN2BEG2 ),
    .Y(_0364_),
    .B1(_0363_));
 sg13g2_or2_1 _1699_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0365_),
    .B(_0364_),
    .A(_0362_));
 sg13g2_mux4_1 _1700_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit3.Q ),
    .A0(NN4END[3]),
    .A1(S2END[6]),
    .A2(E2END[6]),
    .A3(W2END[6]),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit2.Q ),
    .X(_0366_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1701_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit23.Q ),
    .VDD(VPWR),
    .Y(_0367_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit22.Q ),
    .A2(_0366_));
 sg13g2_a21oi_1 _1702_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit22.Q ),
    .A2(_0365_),
    .Y(_0368_),
    .B1(_0367_));
 sg13g2_mux4_1 _1703_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit10.Q ),
    .A0(A),
    .A1(B),
    .A2(C),
    .A3(D),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit11.Q ),
    .X(_0369_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _1704_ (.Y(_0370_),
    .B(_0369_),
    .A_N(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit12.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _1705_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit10.Q ),
    .B(F),
    .Y(_0371_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1706_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit10.Q ),
    .A2(_1051_),
    .Y(_0372_),
    .B1(_0371_));
 sg13g2_nand2b_1 _1707_ (.Y(_0373_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit10.Q ),
    .A_N(\Inst_LUT4AB_switch_matrix.M_AB ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1708_ (.B1(_0373_),
    .VDD(VPWR),
    .Y(_0374_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit10.Q ),
    .A2(H));
 sg13g2_o21ai_1 _1709_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit12.Q ),
    .VDD(VPWR),
    .Y(_0375_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit11.Q ),
    .A2(_0372_));
 sg13g2_a21oi_1 _1710_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit11.Q ),
    .A2(_0374_),
    .Y(_0376_),
    .B1(_0375_));
 sg13g2_nor2b_1 _1711_ (.A(_0376_),
    .B_N(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit13.Q ),
    .Y(_0377_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _1712_ (.Y(_0378_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit10.Q ),
    .A_N(E2END[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1713_ (.B1(_0378_),
    .VDD(VPWR),
    .Y(_0379_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit10.Q ),
    .A2(E1END[1]));
 sg13g2_mux2_1 _1714_ (.A0(N1END[1]),
    .A1(N2END[5]),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit10.Q ),
    .X(_0380_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1715_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit11.Q ),
    .A2(_0379_),
    .Y(_0381_),
    .B1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit12.Q ));
 sg13g2_o21ai_1 _1716_ (.B1(_0381_),
    .VDD(VPWR),
    .Y(_0382_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit11.Q ),
    .A2(_0380_));
 sg13g2_nand2b_1 _1717_ (.Y(_0383_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit10.Q ),
    .A_N(W1END[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1718_ (.B1(_0383_),
    .VDD(VPWR),
    .Y(_0384_),
    .VSS(VGND),
    .A1(W1END[1]),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit10.Q ));
 sg13g2_mux2_1 _1719_ (.A0(S1END[1]),
    .A1(S2END[5]),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit10.Q ),
    .X(_0385_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1720_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit12.Q ),
    .VDD(VPWR),
    .Y(_0386_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit11.Q ),
    .A2(_0385_));
 sg13g2_a21oi_1 _1721_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit11.Q ),
    .A2(_0384_),
    .Y(_0387_),
    .B1(_0386_));
 sg13g2_nor2_1 _1722_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit13.Q ),
    .B(_0387_),
    .Y(_0388_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _1723_ (.Y(\Inst_LUT4AB_switch_matrix.JN2BEG4 ),
    .B1(_0382_),
    .B2(_0388_),
    .A2(_0377_),
    .A1(_0370_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _1724_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit3.Q ),
    .A0(E2MID[6]),
    .A1(W2MID[6]),
    .A2(S2MID[6]),
    .A3(\Inst_LUT4AB_switch_matrix.JN2BEG4 ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit2.Q ),
    .X(_0389_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _1725_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit2.Q ),
    .A0(N2MID[7]),
    .A1(E2MID[7]),
    .A2(S2MID[7]),
    .A3(W2MID[7]),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit3.Q ),
    .X(_0390_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _1726_ (.VDD(VPWR),
    .Y(_0391_),
    .A(_0390_),
    .VSS(VGND));
 sg13g2_a21oi_1 _1727_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit22.Q ),
    .A2(_0391_),
    .Y(_0392_),
    .B1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit23.Q ));
 sg13g2_o21ai_1 _1728_ (.B1(_0392_),
    .VDD(VPWR),
    .Y(_0393_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit22.Q ),
    .A2(_0389_));
 sg13g2_nand2b_1 _1729_ (.Y(_0394_),
    .B(_0393_),
    .A_N(_0368_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _1730_ (.A0(_0394_),
    .A1(_0207_),
    .S(\Inst_LC_LUT4c_frame_config_dffesr.c_I0mux ),
    .X(_0395_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1731_ (.Y(_0396_),
    .A(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ),
    .B(_0395_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _1732_ (.Y(_0397_),
    .B(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ),
    .A_N(_0395_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _1733_ (.B(_0396_),
    .C(_0397_),
    .A(_0206_),
    .Y(_0398_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _1734_ (.Y(_0399_),
    .B(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ),
    .A_N(_0395_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3b_1 _1735_ (.B(_0203_),
    .C(_0399_),
    .Y(_0400_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(_0202_));
 sg13g2_a21oi_1 _1736_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ),
    .A2(_0395_),
    .Y(_0401_),
    .B1(_0400_));
 sg13g2_mux4_1 _1737_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit2.Q ),
    .A0(A),
    .A1(B),
    .A2(D),
    .A3(E),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit3.Q ),
    .X(_0402_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _1738_ (.Y(_0403_),
    .B(_0402_),
    .A_N(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit4.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _1739_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit2.Q ),
    .B(F),
    .Y(_0404_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1740_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit2.Q ),
    .A2(_1051_),
    .Y(_0405_),
    .B1(_0404_));
 sg13g2_nand2b_1 _1741_ (.Y(_0406_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit2.Q ),
    .A_N(\Inst_LUT4AB_switch_matrix.M_EF ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1742_ (.B1(_0406_),
    .VDD(VPWR),
    .Y(_0407_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit2.Q ),
    .A2(H));
 sg13g2_o21ai_1 _1743_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit4.Q ),
    .VDD(VPWR),
    .Y(_0408_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit3.Q ),
    .A2(_0405_));
 sg13g2_a21oi_1 _1744_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit3.Q ),
    .A2(_0407_),
    .Y(_0409_),
    .B1(_0408_));
 sg13g2_nor2b_1 _1745_ (.A(_0409_),
    .B_N(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit5.Q ),
    .Y(_0410_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _1746_ (.A0(S4END[3]),
    .A1(SS4END[3]),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit2.Q ),
    .X(_0411_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1747_ (.Y(_0412_),
    .A(_1028_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit2.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1748_ (.B1(_0412_),
    .VDD(VPWR),
    .Y(_0413_),
    .VSS(VGND),
    .A1(W2END[3]),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit2.Q ));
 sg13g2_o21ai_1 _1749_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit4.Q ),
    .VDD(VPWR),
    .Y(_0414_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit3.Q ),
    .A2(_0411_));
 sg13g2_a21oi_1 _1750_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit3.Q ),
    .A2(_0413_),
    .Y(_0415_),
    .B1(_0414_));
 sg13g2_mux4_1 _1751_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit2.Q ),
    .A0(N1END[1]),
    .A1(N2END[3]),
    .A2(EE4END[3]),
    .A3(E6END[1]),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit3.Q ),
    .X(_0416_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _1752_ (.Y(_0417_),
    .B(_0416_),
    .A_N(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit4.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _1753_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit5.Q ),
    .B(_0415_),
    .Y(_0418_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _1754_ (.Y(\Inst_LUT4AB_switch_matrix.JW2BEG2 ),
    .B1(_0417_),
    .B2(_0418_),
    .A2(_0410_),
    .A1(_0403_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1755_ (.Y(_0419_),
    .A(SS4END[0]),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit8.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1756_ (.B1(_0419_),
    .VDD(VPWR),
    .Y(_0420_),
    .VSS(VGND),
    .A1(_1012_),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit8.Q ));
 sg13g2_nand2_1 _1757_ (.Y(_0421_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit8.Q ),
    .B(\Inst_LUT4AB_switch_matrix.JW2BEG2 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _1758_ (.Y(_0422_),
    .B(W6END[0]),
    .A_N(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit8.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _1759_ (.B(_0421_),
    .C(_0422_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit9.Q ),
    .Y(_0423_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1760_ (.B1(_0423_),
    .VDD(VPWR),
    .Y(_0424_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit9.Q ),
    .A2(_0420_));
 sg13g2_inv_1 _1761_ (.VDD(VPWR),
    .Y(_0425_),
    .A(_0424_),
    .VSS(VGND));
 sg13g2_mux2_1 _1762_ (.A0(N2END[0]),
    .A1(EE4END[1]),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit8.Q ),
    .X(_0426_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _1763_ (.Y(_0427_),
    .B(S2END[0]),
    .A_N(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit8.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1764_ (.Y(_0428_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit8.Q ),
    .B(W2END[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _1765_ (.B(_0427_),
    .C(_0428_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit9.Q ),
    .Y(_0429_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1766_ (.B1(_0429_),
    .VDD(VPWR),
    .Y(_0430_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit9.Q ),
    .A2(_0426_));
 sg13g2_o21ai_1 _1767_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit29.Q ),
    .VDD(VPWR),
    .Y(_0431_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit28.Q ),
    .A2(_0430_));
 sg13g2_a21oi_1 _1768_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit28.Q ),
    .A2(_0425_),
    .Y(_0432_),
    .B1(_0431_));
 sg13g2_mux4_1 _1769_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit10.Q ),
    .A0(A),
    .A1(B),
    .A2(C),
    .A3(D),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit11.Q ),
    .X(_0433_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _1770_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit10.Q ),
    .B(F),
    .Y(_0434_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1771_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit10.Q ),
    .A2(_1051_),
    .Y(_0435_),
    .B1(_0434_));
 sg13g2_o21ai_1 _1772_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit11.Q ),
    .VDD(VPWR),
    .Y(_0436_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit10.Q ),
    .A2(_1052_));
 sg13g2_a21oi_1 _1773_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit10.Q ),
    .A2(\Inst_LUT4AB_switch_matrix.M_AD ),
    .Y(_0437_),
    .B1(_0436_));
 sg13g2_o21ai_1 _1774_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit12.Q ),
    .VDD(VPWR),
    .Y(_0438_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit11.Q ),
    .A2(_0435_));
 sg13g2_o21ai_1 _1775_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit13.Q ),
    .VDD(VPWR),
    .Y(_0439_),
    .VSS(VGND),
    .A1(_0437_),
    .A2(_0438_));
 sg13g2_a21oi_1 _1776_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1039_),
    .A2(_0433_),
    .Y(_0440_),
    .B1(_0439_));
 sg13g2_mux4_1 _1777_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit10.Q ),
    .A0(N1END[1]),
    .A1(N2END[5]),
    .A2(E1END[1]),
    .A3(E2END[5]),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit11.Q ),
    .X(_0441_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _1778_ (.Y(_0442_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit10.Q ),
    .A_N(W1END[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1779_ (.B1(_0442_),
    .VDD(VPWR),
    .Y(_0443_),
    .VSS(VGND),
    .A1(S2END[5]),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit10.Q ));
 sg13g2_mux2_1 _1780_ (.A0(S1END[1]),
    .A1(S1END[3]),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit10.Q ),
    .X(_0444_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _1781_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0445_),
    .B(_0444_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit11.Q ));
 sg13g2_a21oi_1 _1782_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit11.Q ),
    .A2(_0443_),
    .Y(_0446_),
    .B1(_1039_));
 sg13g2_a221oi_1 _1783_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_0446_),
    .C1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit13.Q ),
    .B1(_0445_),
    .A1(_1039_),
    .Y(_0447_),
    .A2(_0441_));
 sg13g2_nor2_1 _1784_ (.A(_0440_),
    .B(_0447_),
    .Y(\Inst_LUT4AB_switch_matrix.JW2BEG4 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _1785_ (.A(\Inst_LUT4AB_switch_matrix.JW2BEG4 ),
    .B_N(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit8.Q ),
    .Y(_0448_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _1786_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit8.Q ),
    .B(W2MID[0]),
    .Y(_0449_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1787_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit9.Q ),
    .VDD(VPWR),
    .Y(_0450_),
    .VSS(VGND),
    .A1(_0448_),
    .A2(_0449_));
 sg13g2_mux2_1 _1788_ (.A0(N2MID[0]),
    .A1(S2MID[0]),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit8.Q ),
    .X(_0451_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1789_ (.B1(_0450_),
    .VDD(VPWR),
    .Y(_0452_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit9.Q ),
    .A2(_0451_));
 sg13g2_mux4_1 _1790_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit8.Q ),
    .A0(N2MID[1]),
    .A1(E2MID[1]),
    .A2(S2MID[1]),
    .A3(W2MID[1]),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit9.Q ),
    .X(_0453_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _1791_ (.VDD(VPWR),
    .Y(_0454_),
    .A(_0453_),
    .VSS(VGND));
 sg13g2_a21oi_1 _1792_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit28.Q ),
    .A2(_0453_),
    .Y(_0455_),
    .B1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit29.Q ));
 sg13g2_o21ai_1 _1793_ (.B1(_0455_),
    .VDD(VPWR),
    .Y(_0456_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit28.Q ),
    .A2(_0452_));
 sg13g2_nor2b_1 _1794_ (.A(_0432_),
    .B_N(_0456_),
    .Y(_0457_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _1795_ (.Y(_0458_),
    .B(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ),
    .A_N(_0395_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3b_1 _1796_ (.B(_0458_),
    .C(_0202_),
    .Y(_0459_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(_0203_));
 sg13g2_a21oi_1 _1797_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ),
    .A2(_0395_),
    .Y(_0460_),
    .B1(_0459_));
 sg13g2_mux2_1 _1798_ (.A0(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ),
    .A1(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ),
    .S(_0395_),
    .X(_0461_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1799_ (.B1(_0398_),
    .VDD(VPWR),
    .Y(_0462_),
    .VSS(VGND),
    .A1(_0204_),
    .A2(_0461_));
 sg13g2_nor4_1 _1800_ (.A(_0401_),
    .B(_0457_),
    .C(_0460_),
    .D(_0462_),
    .Y(_0463_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _1801_ (.S0(_0202_),
    .A0(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ),
    .A1(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ),
    .A2(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ),
    .A3(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ),
    .S1(_0395_),
    .X(_0464_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _1802_ (.S0(_0202_),
    .A0(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ),
    .A1(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ),
    .A2(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ),
    .A3(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ),
    .S1(_0395_),
    .X(_0465_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _1803_ (.A0(_0464_),
    .A1(_0465_),
    .S(_0203_),
    .X(_0466_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _1804_ (.A2(_0466_),
    .A1(_0457_),
    .B1(_0463_),
    .X(_0467_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _1805_ (.A0(_0467_),
    .A1(\Inst_LC_LUT4c_frame_config_dffesr.LUT_flop ),
    .S(\Inst_LC_LUT4c_frame_config_dffesr.c_out_mux ),
    .X(C),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _1806_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit26.Q ),
    .B(_0316_),
    .Y(_0468_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1807_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit26.Q ),
    .A2(_0315_),
    .Y(_0469_),
    .B1(_0468_));
 sg13g2_nand2_1 _1808_ (.Y(_0470_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit26.Q ),
    .B(_0334_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _1809_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit26.Q ),
    .B(_0329_),
    .Y(_0471_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _1810_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit27.Q ),
    .B(_0471_),
    .Y(_0472_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _1811_ (.Y(_0473_),
    .B1(_0470_),
    .B2(_0472_),
    .A2(_0469_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit27.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1812_ (.Y(_0474_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit20.Q ),
    .B(_0237_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1813_ (.B1(_0474_),
    .VDD(VPWR),
    .Y(_0475_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit20.Q ),
    .A2(_0236_));
 sg13g2_or2_1 _1814_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0476_),
    .B(_0475_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit21.Q ));
 sg13g2_nor2b_1 _1815_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit20.Q ),
    .B_N(_0239_),
    .Y(_0477_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1816_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit20.Q ),
    .A2(_0238_),
    .Y(_0478_),
    .B1(_0477_));
 sg13g2_a21o_1 _1817_ (.A2(_0311_),
    .A1(_0209_),
    .B1(_0312_),
    .X(_0479_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1818_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit21.Q ),
    .A2(_0478_),
    .Y(_0480_),
    .B1(\Inst_LF_LUT4c_frame_config_dffesr.c_I0mux ));
 sg13g2_a22oi_1 _1819_ (.Y(_0481_),
    .B1(_0480_),
    .B2(_0476_),
    .A2(_0479_),
    .A1(\Inst_LF_LUT4c_frame_config_dffesr.c_I0mux ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1820_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit25.Q ),
    .VDD(VPWR),
    .Y(_0482_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit24.Q ),
    .A2(_0253_));
 sg13g2_a21oi_1 _1821_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit24.Q ),
    .A2(_0248_),
    .Y(_0483_),
    .B1(_0482_));
 sg13g2_a21oi_1 _1822_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit24.Q ),
    .A2(_0277_),
    .Y(_0484_),
    .B1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit25.Q ));
 sg13g2_o21ai_1 _1823_ (.B1(_0484_),
    .VDD(VPWR),
    .Y(_0485_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit24.Q ),
    .A2(_0276_));
 sg13g2_nand2b_1 _1824_ (.Y(_0486_),
    .B(_0485_),
    .A_N(_0483_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _1825_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit22.Q ),
    .A0(_0307_),
    .A1(_0309_),
    .A2(_0290_),
    .A3(_0286_),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit23.Q ),
    .X(_0487_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _1826_ (.A(_0486_),
    .B(_0487_),
    .Y(_0488_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _1827_ (.S0(_0481_),
    .A0(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ),
    .A1(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ),
    .A2(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ),
    .A3(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ),
    .S1(_0487_),
    .X(_0489_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1828_ (.Y(_0490_),
    .A(_0486_),
    .B(_0487_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _1829_ (.S0(_0481_),
    .A0(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ),
    .A1(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ),
    .A2(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ),
    .A3(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ),
    .S1(_0487_),
    .X(_0491_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _1830_ (.A0(_0489_),
    .A1(_0491_),
    .S(_0486_),
    .X(_0492_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _1831_ (.S0(_0481_),
    .A0(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ),
    .A1(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ),
    .A2(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ),
    .A3(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ),
    .S1(_0487_),
    .X(_0493_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _1832_ (.S0(_0481_),
    .A0(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ),
    .A1(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ),
    .A2(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ),
    .A3(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ),
    .S1(_0487_),
    .X(_0494_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _1833_ (.A0(_0493_),
    .A1(_0494_),
    .S(_0486_),
    .X(_0495_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _1834_ (.A0(_0492_),
    .A1(_0495_),
    .S(_0473_),
    .X(_0496_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _1835_ (.A0(_0496_),
    .A1(\Inst_LF_LUT4c_frame_config_dffesr.LUT_flop ),
    .S(\Inst_LF_LUT4c_frame_config_dffesr.c_out_mux ),
    .X(F),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1836_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit19.Q ),
    .VDD(VPWR),
    .Y(_0497_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit18.Q ),
    .A2(_1052_));
 sg13g2_a21oi_1 _1837_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit18.Q ),
    .A2(\Inst_LUT4AB_switch_matrix.M_AH ),
    .Y(_0498_),
    .B1(_0497_));
 sg13g2_mux2_1 _1838_ (.A0(E),
    .A1(F),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit18.Q ),
    .X(_0499_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1839_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit20.Q ),
    .VDD(VPWR),
    .Y(_0500_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit19.Q ),
    .A2(_0499_));
 sg13g2_or2_1 _1840_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0501_),
    .B(_0500_),
    .A(_0498_));
 sg13g2_nand2b_1 _1841_ (.Y(_0502_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit18.Q ),
    .A_N(D),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1842_ (.B1(_0502_),
    .VDD(VPWR),
    .Y(_0503_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit18.Q ),
    .A2(C));
 sg13g2_mux2_1 _1843_ (.A0(A),
    .A1(B),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit18.Q ),
    .X(_0504_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1844_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit19.Q ),
    .A2(_0503_),
    .Y(_0505_),
    .B1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit20.Q ));
 sg13g2_o21ai_1 _1845_ (.B1(_0505_),
    .VDD(VPWR),
    .Y(_0506_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit19.Q ),
    .A2(_0504_));
 sg13g2_and2_1 _1846_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit21.Q ),
    .B(_0506_),
    .X(_0507_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _1847_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit18.Q ),
    .A0(N1END[3]),
    .A1(N2END[7]),
    .A2(E1END[3]),
    .A3(E2END[7]),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit19.Q ),
    .X(_0508_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _1848_ (.Y(_0509_),
    .B(_0508_),
    .A_N(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit20.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _1849_ (.Y(_0510_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit18.Q ),
    .A_N(W1END[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1850_ (.B1(_0510_),
    .VDD(VPWR),
    .Y(_0511_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit18.Q ),
    .A2(W1END[1]));
 sg13g2_mux2_1 _1851_ (.A0(S1END[3]),
    .A1(S2END[7]),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit18.Q ),
    .X(_0512_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1852_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit20.Q ),
    .VDD(VPWR),
    .Y(_0513_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit19.Q ),
    .A2(_0512_));
 sg13g2_a21oi_1 _1853_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit19.Q ),
    .A2(_0511_),
    .Y(_0514_),
    .B1(_0513_));
 sg13g2_nor2_1 _1854_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit21.Q ),
    .B(_0514_),
    .Y(_0515_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _1855_ (.Y(\Inst_LUT4AB_switch_matrix.JN2BEG6 ),
    .B1(_0509_),
    .B2(_0515_),
    .A2(_0507_),
    .A1(_0501_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _1856_ (.A(\Inst_LUT4AB_switch_matrix.JN2BEG6 ),
    .B_N(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit18.Q ),
    .Y(_0516_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _1857_ (.A(S2MID[6]),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit18.Q ),
    .Y(_0517_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1858_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit19.Q ),
    .VDD(VPWR),
    .Y(_0518_),
    .VSS(VGND),
    .A1(_0516_),
    .A2(_0517_));
 sg13g2_mux2_1 _1859_ (.A0(N2MID[6]),
    .A1(E2MID[6]),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit18.Q ),
    .X(_0519_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1860_ (.B1(_0518_),
    .VDD(VPWR),
    .Y(_0520_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit19.Q ),
    .A2(_0519_));
 sg13g2_mux2_1 _1861_ (.A0(N2MID[7]),
    .A1(E2MID[7]),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit18.Q ),
    .X(_0521_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _1862_ (.Y(_0522_),
    .B(S2MID[7]),
    .A_N(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit18.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1863_ (.Y(_0523_),
    .A(W2MID[7]),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit18.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _1864_ (.B(_0522_),
    .C(_0523_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit19.Q ),
    .Y(_0524_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1865_ (.B1(_0524_),
    .VDD(VPWR),
    .Y(_0525_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit19.Q ),
    .A2(_0521_));
 sg13g2_mux4_1 _1866_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit18.Q ),
    .A0(N4END[3]),
    .A1(EE4END[0]),
    .A2(S4END[3]),
    .A3(\Inst_LUT4AB_switch_matrix.JN2BEG4 ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit19.Q ),
    .X(_0526_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _1867_ (.VDD(VPWR),
    .Y(_0527_),
    .A(_0526_),
    .VSS(VGND));
 sg13g2_mux4_1 _1868_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit18.Q ),
    .A0(N2END[7]),
    .A1(E2END[7]),
    .A2(S2END[7]),
    .A3(WW4END[0]),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit19.Q ),
    .X(_0528_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _1869_ (.VDD(VPWR),
    .Y(_0529_),
    .A(_0528_),
    .VSS(VGND));
 sg13g2_mux4_1 _1870_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit30.Q ),
    .A0(_0520_),
    .A1(_0525_),
    .A2(_0529_),
    .A3(_0527_),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit31.Q ),
    .X(_0530_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1871_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0479_),
    .A2(_0490_),
    .Y(_0531_),
    .B1(_0488_));
 sg13g2_mux2_1 _1872_ (.A0(_0530_),
    .A1(_0531_),
    .S(\Inst_LG_LUT4c_frame_config_dffesr.c_I0mux ),
    .X(_0532_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _1873_ (.A0(E6END[1]),
    .A1(S4END[1]),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit22.Q ),
    .X(_0533_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1874_ (.Y(_0534_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit22.Q ),
    .B(\Inst_LUT4AB_switch_matrix.JS2BEG4 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _1875_ (.Y(_0535_),
    .B(WW4END[3]),
    .A_N(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit22.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _1876_ (.B(_0534_),
    .C(_0535_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit23.Q ),
    .Y(_0536_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1877_ (.B1(_0536_),
    .VDD(VPWR),
    .Y(_0537_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit23.Q ),
    .A2(_0533_));
 sg13g2_mux4_1 _1878_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit23.Q ),
    .A0(NN4END[1]),
    .A1(S2END[5]),
    .A2(E2END[5]),
    .A3(W2END[5]),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit22.Q ),
    .X(_0538_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _1879_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit18.Q ),
    .A0(A),
    .A1(B),
    .A2(C),
    .A3(D),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit19.Q ),
    .X(_0539_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _1880_ (.A0(E),
    .A1(F),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit18.Q ),
    .X(_0540_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1881_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit19.Q ),
    .VDD(VPWR),
    .Y(_0541_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit18.Q ),
    .A2(_1052_));
 sg13g2_a21oi_1 _1882_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit18.Q ),
    .A2(\Inst_LUT4AB_switch_matrix.M_AB ),
    .Y(_0542_),
    .B1(_0541_));
 sg13g2_o21ai_1 _1883_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit20.Q ),
    .VDD(VPWR),
    .Y(_0543_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit19.Q ),
    .A2(_0540_));
 sg13g2_o21ai_1 _1884_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit21.Q ),
    .VDD(VPWR),
    .Y(_0544_),
    .VSS(VGND),
    .A1(_0542_),
    .A2(_0543_));
 sg13g2_a21oi_1 _1885_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1044_),
    .A2(_0539_),
    .Y(_0545_),
    .B1(_0544_));
 sg13g2_mux4_1 _1886_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit18.Q ),
    .A0(N1END[3]),
    .A1(N2END[7]),
    .A2(E1END[3]),
    .A3(E2END[7]),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit19.Q ),
    .X(_0546_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _1887_ (.Y(_0547_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit18.Q ),
    .A_N(W1END[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1888_ (.B1(_0547_),
    .VDD(VPWR),
    .Y(_0548_),
    .VSS(VGND),
    .A1(W1END[1]),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit18.Q ));
 sg13g2_mux2_1 _1889_ (.A0(S1END[3]),
    .A1(S2END[7]),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit18.Q ),
    .X(_0549_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _1890_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0550_),
    .B(_0549_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit19.Q ));
 sg13g2_a21oi_1 _1891_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit19.Q ),
    .A2(_0548_),
    .Y(_0551_),
    .B1(_1044_));
 sg13g2_a221oi_1 _1892_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_0551_),
    .C1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit21.Q ),
    .B1(_0550_),
    .A1(_1044_),
    .Y(_0552_),
    .A2(_0546_));
 sg13g2_nor2_1 _1893_ (.A(_0545_),
    .B(_0552_),
    .Y(\Inst_LUT4AB_switch_matrix.JS2BEG6 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1894_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit23.Q ),
    .VDD(VPWR),
    .Y(_0553_),
    .VSS(VGND),
    .A1(_1026_),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit22.Q ));
 sg13g2_a21o_1 _1895_ (.A2(\Inst_LUT4AB_switch_matrix.JS2BEG6 ),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit22.Q ),
    .B1(_0553_),
    .X(_0554_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _1896_ (.A0(E2MID[4]),
    .A1(S2MID[4]),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit22.Q ),
    .X(_0555_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1897_ (.B1(_0554_),
    .VDD(VPWR),
    .Y(_0556_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit23.Q ),
    .A2(_0555_));
 sg13g2_mux2_1 _1898_ (.A0(N2MID[5]),
    .A1(E2MID[5]),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit22.Q ),
    .X(_0557_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _1899_ (.Y(_0558_),
    .B(S2MID[5]),
    .A_N(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit22.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1900_ (.Y(_0559_),
    .A(W2MID[5]),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit22.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _1901_ (.B(_0558_),
    .C(_0559_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit23.Q ),
    .Y(_0560_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1902_ (.B1(_0560_),
    .VDD(VPWR),
    .Y(_0561_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit23.Q ),
    .A2(_0557_));
 sg13g2_mux2_1 _1903_ (.A0(_0556_),
    .A1(_0561_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit2.Q ),
    .X(_0562_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1904_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit3.Q ),
    .VDD(VPWR),
    .Y(_0563_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit2.Q ),
    .A2(_0538_));
 sg13g2_a21o_1 _1905_ (.A2(_0537_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit2.Q ),
    .B1(_0563_),
    .X(_0564_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1906_ (.B1(_0564_),
    .VDD(VPWR),
    .Y(_0565_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit3.Q ),
    .A2(_0562_));
 sg13g2_mux4_1 _1907_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit18.Q ),
    .A0(A),
    .A1(B),
    .A2(C),
    .A3(D),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit19.Q ),
    .X(_0566_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _1908_ (.Y(_0567_),
    .B(_0566_),
    .A_N(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit20.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _1909_ (.A0(E),
    .A1(F),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit18.Q ),
    .X(_0568_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _1910_ (.Y(_0569_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit18.Q ),
    .A_N(\Inst_LUT4AB_switch_matrix.M_AD ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1911_ (.B1(_0569_),
    .VDD(VPWR),
    .Y(_0570_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit18.Q ),
    .A2(H));
 sg13g2_o21ai_1 _1912_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit20.Q ),
    .VDD(VPWR),
    .Y(_0571_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit19.Q ),
    .A2(_0568_));
 sg13g2_a21oi_1 _1913_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit19.Q ),
    .A2(_0570_),
    .Y(_0572_),
    .B1(_0571_));
 sg13g2_nor2b_1 _1914_ (.A(_0572_),
    .B_N(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit21.Q ),
    .Y(_0573_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _1915_ (.Y(_0574_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit18.Q ),
    .A_N(E2END[7]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1916_ (.B1(_0574_),
    .VDD(VPWR),
    .Y(_0575_),
    .VSS(VGND),
    .A1(E1END[3]),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit18.Q ));
 sg13g2_mux2_1 _1917_ (.A0(N1END[3]),
    .A1(N2END[7]),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit18.Q ),
    .X(_0576_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1918_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit19.Q ),
    .A2(_0575_),
    .Y(_0577_),
    .B1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit20.Q ));
 sg13g2_o21ai_1 _1919_ (.B1(_0577_),
    .VDD(VPWR),
    .Y(_0578_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit19.Q ),
    .A2(_0576_));
 sg13g2_nand2b_1 _1920_ (.Y(_0579_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit18.Q ),
    .A_N(W1END[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1921_ (.B1(_0579_),
    .VDD(VPWR),
    .Y(_0580_),
    .VSS(VGND),
    .A1(S2END[7]),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit18.Q ));
 sg13g2_mux2_1 _1922_ (.A0(S1END[1]),
    .A1(S1END[3]),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit18.Q ),
    .X(_0581_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1923_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit20.Q ),
    .VDD(VPWR),
    .Y(_0582_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit19.Q ),
    .A2(_0581_));
 sg13g2_a21oi_1 _1924_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit19.Q ),
    .A2(_0580_),
    .Y(_0583_),
    .B1(_0582_));
 sg13g2_nor2_1 _1925_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit21.Q ),
    .B(_0583_),
    .Y(_0584_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _1926_ (.Y(\Inst_LUT4AB_switch_matrix.E2BEG6 ),
    .B1(_0578_),
    .B2(_0584_),
    .A2(_0573_),
    .A1(_0567_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _1927_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit21.Q ),
    .A0(N2MID[2]),
    .A1(W2MID[2]),
    .A2(S2MID[2]),
    .A3(\Inst_LUT4AB_switch_matrix.E2BEG6 ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit20.Q ),
    .X(_0585_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _1928_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit20.Q ),
    .A0(N2MID[3]),
    .A1(E2MID[3]),
    .A2(S2MID[3]),
    .A3(W2MID[3]),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit21.Q ),
    .X(_0586_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _1929_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit21.Q ),
    .A0(N4END[2]),
    .A1(W2END[2]),
    .A2(SS4END[2]),
    .A3(\Inst_LUT4AB_switch_matrix.E2BEG4 ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit20.Q ),
    .X(_0587_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _1930_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit21.Q ),
    .A0(N2END[3]),
    .A1(SS4END[0]),
    .A2(E2END[3]),
    .A3(W2END[3]),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit20.Q ),
    .X(_0588_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _1931_ (.VDD(VPWR),
    .Y(_0589_),
    .A(_0588_),
    .VSS(VGND));
 sg13g2_mux4_1 _1932_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit0.Q ),
    .A0(_0585_),
    .A1(_0586_),
    .A2(_0588_),
    .A3(_0587_),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit1.Q ),
    .X(_0590_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _1933_ (.A(_0565_),
    .B(_0590_),
    .Y(_0591_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _1934_ (.S0(_0590_),
    .A0(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ),
    .A1(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ),
    .A2(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ),
    .A3(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ),
    .S1(_0565_),
    .X(_0592_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _1935_ (.VDD(VPWR),
    .Y(_0593_),
    .A(_0592_),
    .VSS(VGND));
 sg13g2_o21ai_1 _1936_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit19.Q ),
    .VDD(VPWR),
    .Y(_0594_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit18.Q ),
    .A2(_1052_));
 sg13g2_a21oi_1 _1937_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit18.Q ),
    .A2(\Inst_LUT4AB_switch_matrix.M_EF ),
    .Y(_0595_),
    .B1(_0594_));
 sg13g2_mux2_1 _1938_ (.A0(E),
    .A1(F),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit18.Q ),
    .X(_0596_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1939_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit20.Q ),
    .VDD(VPWR),
    .Y(_0597_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit19.Q ),
    .A2(_0596_));
 sg13g2_or2_1 _1940_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0598_),
    .B(_0597_),
    .A(_0595_));
 sg13g2_nand2b_1 _1941_ (.Y(_0599_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit18.Q ),
    .A_N(D),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1942_ (.B1(_0599_),
    .VDD(VPWR),
    .Y(_0600_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit18.Q ),
    .A2(C));
 sg13g2_mux2_1 _1943_ (.A0(A),
    .A1(B),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit18.Q ),
    .X(_0601_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1944_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit19.Q ),
    .A2(_0600_),
    .Y(_0602_),
    .B1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit20.Q ));
 sg13g2_o21ai_1 _1945_ (.B1(_0602_),
    .VDD(VPWR),
    .Y(_0603_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit19.Q ),
    .A2(_0601_));
 sg13g2_and2_1 _1946_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit21.Q ),
    .B(_0603_),
    .X(_0604_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _1947_ (.A0(S1END[1]),
    .A1(S1END[3]),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit18.Q ),
    .X(_0605_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _1948_ (.Y(_0606_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit18.Q ),
    .A_N(W1END[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1949_ (.B1(_0606_),
    .VDD(VPWR),
    .Y(_0607_),
    .VSS(VGND),
    .A1(S2END[7]),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit18.Q ));
 sg13g2_o21ai_1 _1950_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit20.Q ),
    .VDD(VPWR),
    .Y(_0608_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit19.Q ),
    .A2(_0605_));
 sg13g2_a21oi_1 _1951_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit19.Q ),
    .A2(_0607_),
    .Y(_0609_),
    .B1(_0608_));
 sg13g2_mux4_1 _1952_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit18.Q ),
    .A0(N1END[3]),
    .A1(N2END[7]),
    .A2(E1END[3]),
    .A3(E2END[7]),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit19.Q ),
    .X(_0610_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _1953_ (.Y(_0611_),
    .B(_0610_),
    .A_N(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit20.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _1954_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit21.Q ),
    .B(_0609_),
    .Y(_0612_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _1955_ (.Y(\Inst_LUT4AB_switch_matrix.JW2BEG6 ),
    .B1(_0611_),
    .B2(_0612_),
    .A2(_0604_),
    .A1(_0598_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _1956_ (.A(\Inst_LUT4AB_switch_matrix.JW2BEG6 ),
    .B_N(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit24.Q ),
    .Y(_0613_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _1957_ (.A(W2MID[0]),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit24.Q ),
    .Y(_0614_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1958_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit25.Q ),
    .VDD(VPWR),
    .Y(_0615_),
    .VSS(VGND),
    .A1(_0613_),
    .A2(_0614_));
 sg13g2_mux2_1 _1959_ (.A0(N2MID[0]),
    .A1(E2MID[0]),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit24.Q ),
    .X(_0616_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1960_ (.B1(_0615_),
    .VDD(VPWR),
    .Y(_0617_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit25.Q ),
    .A2(_0616_));
 sg13g2_mux2_1 _1961_ (.A0(N2MID[1]),
    .A1(E2MID[1]),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit24.Q ),
    .X(_0618_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _1962_ (.Y(_0619_),
    .B(S2MID[1]),
    .A_N(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit24.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1963_ (.Y(_0620_),
    .A(W2MID[1]),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit24.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _1964_ (.B(_0619_),
    .C(_0620_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit25.Q ),
    .Y(_0621_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1965_ (.B1(_0621_),
    .VDD(VPWR),
    .Y(_0622_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit25.Q ),
    .A2(_0618_));
 sg13g2_mux4_1 _1966_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit25.Q ),
    .A0(NN4END[0]),
    .A1(W2END[0]),
    .A2(E6END[0]),
    .A3(\Inst_LUT4AB_switch_matrix.JW2BEG4 ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit24.Q ),
    .X(_0623_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _1967_ (.VDD(VPWR),
    .Y(_0624_),
    .A(_0623_),
    .VSS(VGND));
 sg13g2_mux4_1 _1968_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit25.Q ),
    .A0(N2END[1]),
    .A1(S2END[1]),
    .A2(EE4END[3]),
    .A3(W2END[1]),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit24.Q ),
    .X(_0625_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _1969_ (.VDD(VPWR),
    .Y(_0626_),
    .A(_0625_),
    .VSS(VGND));
 sg13g2_mux4_1 _1970_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit4.Q ),
    .A0(_0617_),
    .A1(_0622_),
    .A2(_0626_),
    .A3(_0624_),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit5.Q ),
    .X(_0627_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _1971_ (.S0(_0590_),
    .A0(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ),
    .A1(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ),
    .A2(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ),
    .A3(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ),
    .S1(_0565_),
    .X(_0628_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1972_ (.B1(_0627_),
    .VDD(VPWR),
    .Y(_0629_),
    .VSS(VGND),
    .A1(_0532_),
    .A2(_0628_));
 sg13g2_a21oi_1 _1973_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0532_),
    .A2(_0593_),
    .Y(_0630_),
    .B1(_0629_));
 sg13g2_mux4_1 _1974_ (.S0(_0590_),
    .A0(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ),
    .A1(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ),
    .A2(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ),
    .A3(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ),
    .S1(_0565_),
    .X(_0631_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _1975_ (.Y(_0632_),
    .B(_0532_),
    .A_N(_0631_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _1976_ (.S0(_0590_),
    .A0(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ),
    .A1(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ),
    .A2(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ),
    .A3(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ),
    .S1(_0565_),
    .X(_0633_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _1977_ (.A(_0532_),
    .B(_0633_),
    .Y(_0634_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _1978_ (.A(_0627_),
    .B(_0634_),
    .Y(_0635_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1979_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0632_),
    .A2(_0635_),
    .Y(_0636_),
    .B1(_0630_));
 sg13g2_nand2_1 _1980_ (.Y(_0637_),
    .A(\Inst_LG_LUT4c_frame_config_dffesr.LUT_flop ),
    .B(\Inst_LG_LUT4c_frame_config_dffesr.c_out_mux ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1981_ (.B1(_0637_),
    .VDD(VPWR),
    .Y(G),
    .VSS(VGND),
    .A1(\Inst_LG_LUT4c_frame_config_dffesr.c_out_mux ),
    .A2(_0636_));
 sg13g2_a221oi_1 _1982_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_0590_),
    .C1(_0488_),
    .B1(_0565_),
    .A1(_0479_),
    .Y(_0638_),
    .A2(_0490_));
 sg13g2_or2_1 _1983_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0639_),
    .B(_0638_),
    .A(_0591_));
 sg13g2_o21ai_1 _1984_ (.B1(\Inst_LH_LUT4c_frame_config_dffesr.c_I0mux ),
    .VDD(VPWR),
    .Y(_0640_),
    .VSS(VGND),
    .A1(_0591_),
    .A2(_0638_));
 sg13g2_o21ai_1 _1985_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit9.Q ),
    .VDD(VPWR),
    .Y(_0641_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit8.Q ),
    .A2(_0528_));
 sg13g2_a21oi_1 _1986_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit8.Q ),
    .A2(_0527_),
    .Y(_0642_),
    .B1(_0641_));
 sg13g2_mux2_1 _1987_ (.A0(_0520_),
    .A1(_0525_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit8.Q ),
    .X(_0643_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _1988_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit9.Q ),
    .B(_0643_),
    .Y(_0644_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or3_1 _1989_ (.A(\Inst_LH_LUT4c_frame_config_dffesr.c_I0mux ),
    .B(_0642_),
    .C(_0644_),
    .X(_0645_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _1990_ (.A0(_0556_),
    .A1(_0561_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit12.Q ),
    .X(_0646_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1991_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit13.Q ),
    .VDD(VPWR),
    .Y(_0647_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit12.Q ),
    .A2(_0538_));
 sg13g2_a21o_1 _1992_ (.A2(_0537_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit12.Q ),
    .B1(_0647_),
    .X(_0648_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1993_ (.B1(_0648_),
    .VDD(VPWR),
    .Y(_0649_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit13.Q ),
    .A2(_0646_));
 sg13g2_mux4_1 _1994_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit10.Q ),
    .A0(_0585_),
    .A1(_0586_),
    .A2(_0588_),
    .A3(_0587_),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit11.Q ),
    .X(_0650_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1995_ (.Y(_0651_),
    .A(_0649_),
    .B(_0650_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _1996_ (.A(_0649_),
    .B(_0650_),
    .Y(_0652_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _1997_ (.S0(_0650_),
    .A0(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ),
    .A1(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ),
    .A2(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ),
    .A3(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ),
    .S1(_0649_),
    .X(_0653_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _1998_ (.A2(_0645_),
    .A1(_0640_),
    .B1(_0653_),
    .X(_0654_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _1999_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit14.Q ),
    .A0(_0617_),
    .A1(_0622_),
    .A2(_0626_),
    .A3(_0624_),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit15.Q ),
    .X(_0655_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _2000_ (.S0(_0650_),
    .A0(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ),
    .A1(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ),
    .A2(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ),
    .A3(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ),
    .S1(_0649_),
    .X(_0656_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _2001_ (.VDD(VPWR),
    .Y(_0657_),
    .A(_0656_),
    .VSS(VGND));
 sg13g2_nand3_1 _2002_ (.B(_0645_),
    .C(_0657_),
    .A(_0640_),
    .Y(_0658_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_1 _2003_ (.X(_0659_),
    .A(_0654_),
    .B(_0655_),
    .C(_0658_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _2004_ (.S0(_0650_),
    .A0(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ),
    .A1(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ),
    .A2(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ),
    .A3(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ),
    .S1(_0649_),
    .X(_0660_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _2005_ (.A2(_0645_),
    .A1(_0640_),
    .B1(_0660_),
    .X(_0661_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _2006_ (.S0(_0650_),
    .A0(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ),
    .A1(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ),
    .A2(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ),
    .A3(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ),
    .S1(_0649_),
    .X(_0662_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _2007_ (.VDD(VPWR),
    .Y(_0663_),
    .A(_0662_),
    .VSS(VGND));
 sg13g2_nand3_1 _2008_ (.B(_0645_),
    .C(_0663_),
    .A(_0640_),
    .Y(_0664_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _2009_ (.A(_0655_),
    .B_N(_0664_),
    .Y(_0665_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2010_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0661_),
    .A2(_0665_),
    .Y(_0666_),
    .B1(_0659_));
 sg13g2_nand2_1 _2011_ (.Y(_0667_),
    .A(\Inst_LH_LUT4c_frame_config_dffesr.LUT_flop ),
    .B(\Inst_LH_LUT4c_frame_config_dffesr.c_out_mux ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2012_ (.B1(_0667_),
    .VDD(VPWR),
    .Y(H),
    .VSS(VGND),
    .A1(\Inst_LH_LUT4c_frame_config_dffesr.c_out_mux ),
    .A2(_0666_));
 sg13g2_mux4_1 _2013_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit23.Q ),
    .A0(\Inst_LUT4AB_switch_matrix.JN2BEG6 ),
    .A1(\Inst_LUT4AB_switch_matrix.JS2BEG6 ),
    .A2(\Inst_LUT4AB_switch_matrix.E2BEG6 ),
    .A3(\Inst_LUT4AB_switch_matrix.JW2BEG6 ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit22.Q ),
    .X(_0668_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _2014_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit19.Q ),
    .A0(\Inst_LUT4AB_switch_matrix.JN2BEG4 ),
    .A1(\Inst_LUT4AB_switch_matrix.JS2BEG4 ),
    .A2(\Inst_LUT4AB_switch_matrix.E2BEG4 ),
    .A3(\Inst_LUT4AB_switch_matrix.JW2BEG4 ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit18.Q ),
    .X(_0669_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _2015_ (.A0(_0668_),
    .A1(_0669_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit17.Q ),
    .X(_0670_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _2016_ (.A0(E),
    .A1(F),
    .S(_0670_),
    .X(\Inst_LUT4AB_switch_matrix.M_EF ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2017_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit1.Q ),
    .VDD(VPWR),
    .Y(_0671_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit0.Q ),
    .A2(_0366_));
 sg13g2_a21o_1 _2018_ (.A2(_0365_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit0.Q ),
    .B1(_0671_),
    .X(_0672_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2019_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit0.Q ),
    .A2(_0391_),
    .Y(_0673_),
    .B1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit1.Q ));
 sg13g2_o21ai_1 _2020_ (.B1(_0673_),
    .VDD(VPWR),
    .Y(_0674_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit0.Q ),
    .A2(_0389_));
 sg13g2_nor2b_1 _2021_ (.A(\Inst_LD_LUT4c_frame_config_dffesr.c_I0mux ),
    .B_N(_0674_),
    .Y(_0675_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2022_ (.Y(_0676_),
    .B1(_0672_),
    .B2(_0675_),
    .A2(_0208_),
    .A1(\Inst_LD_LUT4c_frame_config_dffesr.c_I0mux ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _2023_ (.S0(_0149_),
    .A0(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ),
    .A1(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ),
    .A2(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ),
    .A3(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ),
    .S1(_0199_),
    .X(_0677_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2024_ (.A(_0676_),
    .B(_0677_),
    .Y(_0678_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _2025_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit6.Q ),
    .A0(_0452_),
    .A1(_0454_),
    .A2(_0430_),
    .A3(_0424_),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit7.Q ),
    .X(_0679_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _2026_ (.S0(_0149_),
    .A0(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ),
    .A1(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ),
    .A2(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ),
    .A3(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ),
    .S1(_0199_),
    .X(_0680_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _2027_ (.A(_0680_),
    .B_N(_0676_),
    .Y(_0681_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _2028_ (.A(_0678_),
    .B(_0679_),
    .C(_0681_),
    .Y(_0682_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _2029_ (.S0(_0149_),
    .A0(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ),
    .A1(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ),
    .A2(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ),
    .A3(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ),
    .S1(_0199_),
    .X(_0683_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _2030_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0684_),
    .B(_0683_),
    .A(_0676_));
 sg13g2_mux4_1 _2031_ (.S0(_0149_),
    .A0(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ),
    .A1(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ),
    .A2(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ),
    .A3(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ),
    .S1(_0199_),
    .X(_0685_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _2032_ (.Y(_0686_),
    .B(_0676_),
    .A_N(_0685_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _2033_ (.A(_0679_),
    .B(_0686_),
    .X(_0687_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _2034_ (.A2(_0687_),
    .A1(_0684_),
    .B1(_0682_),
    .X(_0688_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _2035_ (.A0(_0688_),
    .A1(\Inst_LD_LUT4c_frame_config_dffesr.LUT_flop ),
    .S(\Inst_LD_LUT4c_frame_config_dffesr.c_out_mux ),
    .X(D),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2036_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit20.Q ),
    .A2(\Inst_LUT4AB_switch_matrix.E2BEG5 ),
    .Y(_0689_),
    .B1(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit21.Q ));
 sg13g2_o21ai_1 _2037_ (.B1(_0689_),
    .VDD(VPWR),
    .Y(_0690_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit20.Q ),
    .A2(_0230_));
 sg13g2_a21oi_1 _2038_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit20.Q ),
    .A2(\Inst_LUT4AB_switch_matrix.JW2BEG5 ),
    .Y(_0691_),
    .B1(_1047_));
 sg13g2_o21ai_1 _2039_ (.B1(_0691_),
    .VDD(VPWR),
    .Y(_0692_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit20.Q ),
    .A2(_0275_));
 sg13g2_nand2_1 _2040_ (.Y(_0693_),
    .A(_0690_),
    .B(_0692_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2041_ (.Y(_0694_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit16.Q ),
    .B(_0669_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2042_ (.B1(_0694_),
    .VDD(VPWR),
    .Y(_0695_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit16.Q ),
    .A2(_0693_));
 sg13g2_mux2_1 _2043_ (.A0(C),
    .A1(D),
    .S(_0695_),
    .X(_0696_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _2044_ (.A0(_0696_),
    .A1(\Inst_LUT4AB_switch_matrix.M_AB ),
    .S(_0693_),
    .X(_0697_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _2045_ (.A0(_0696_),
    .A1(_0697_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit16.Q ),
    .X(\Inst_LUT4AB_switch_matrix.M_AD ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2046_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit23.Q ),
    .VDD(VPWR),
    .Y(_0698_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit22.Q ),
    .A2(_1051_));
 sg13g2_a21oi_1 _2047_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit22.Q ),
    .A2(\Inst_LUT4AB_switch_matrix.M_AD ),
    .Y(_0699_),
    .B1(_0698_));
 sg13g2_mux2_1 _2048_ (.A0(E),
    .A1(F),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit22.Q ),
    .X(_0700_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2049_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit24.Q ),
    .VDD(VPWR),
    .Y(_0701_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit23.Q ),
    .A2(_0700_));
 sg13g2_mux4_1 _2050_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit22.Q ),
    .A0(A),
    .A1(B),
    .A2(C),
    .A3(D),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit23.Q ),
    .X(_0702_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2051_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit25.Q ),
    .VDD(VPWR),
    .Y(_0703_),
    .VSS(VGND),
    .A1(_0699_),
    .A2(_0701_));
 sg13g2_a21oi_1 _2052_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1045_),
    .A2(_0702_),
    .Y(_0704_),
    .B1(_0703_));
 sg13g2_mux4_1 _2053_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit22.Q ),
    .A0(N1END[0]),
    .A1(N2END[0]),
    .A2(E1END[0]),
    .A3(E2END[0]),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit23.Q ),
    .X(_0705_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _2054_ (.Y(_0706_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit22.Q ),
    .A_N(W1END[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2055_ (.B1(_0706_),
    .VDD(VPWR),
    .Y(_0707_),
    .VSS(VGND),
    .A1(W1END[0]),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit22.Q ));
 sg13g2_mux2_1 _2056_ (.A0(S1END[0]),
    .A1(S2END[0]),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit22.Q ),
    .X(_0708_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2057_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit24.Q ),
    .VDD(VPWR),
    .Y(_0709_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit23.Q ),
    .A2(_0708_));
 sg13g2_a21oi_1 _2058_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit23.Q ),
    .A2(_0707_),
    .Y(_0710_),
    .B1(_0709_));
 sg13g2_a21oi_1 _2059_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1045_),
    .A2(_0705_),
    .Y(_0711_),
    .B1(_0710_));
 sg13g2_a21oi_1 _2060_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1046_),
    .A2(_0711_),
    .Y(\Inst_LUT4AB_switch_matrix.JS2BEG7 ),
    .B1(_0704_));
 sg13g2_mux4_1 _2061_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit23.Q ),
    .A0(E),
    .A1(G),
    .A2(F),
    .A3(\Inst_LUT4AB_switch_matrix.M_AB ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit22.Q ),
    .X(_0712_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _2062_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit22.Q ),
    .A0(A),
    .A1(B),
    .A2(C),
    .A3(D),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit23.Q ),
    .X(_0713_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _2063_ (.Y(_0714_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit24.Q ),
    .A_N(_0712_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2064_ (.B1(_0714_),
    .VDD(VPWR),
    .Y(_0715_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit24.Q ),
    .A2(_0713_));
 sg13g2_mux4_1 _2065_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit22.Q ),
    .A0(N1END[0]),
    .A1(NN4END[0]),
    .A2(E1END[0]),
    .A3(E2END[0]),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit23.Q ),
    .X(_0716_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _2066_ (.Y(_0717_),
    .B(_0716_),
    .A_N(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit24.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _2067_ (.A0(S1END[0]),
    .A1(S1END[2]),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit22.Q ),
    .X(_0718_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _2068_ (.Y(_0719_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit22.Q ),
    .A_N(W1END[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2069_ (.B1(_0719_),
    .VDD(VPWR),
    .Y(_0720_),
    .VSS(VGND),
    .A1(S2END[0]),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit22.Q ));
 sg13g2_o21ai_1 _2070_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit24.Q ),
    .VDD(VPWR),
    .Y(_0721_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit23.Q ),
    .A2(_0718_));
 sg13g2_a21oi_1 _2071_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit23.Q ),
    .A2(_0720_),
    .Y(_0722_),
    .B1(_0721_));
 sg13g2_nor2_1 _2072_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit25.Q ),
    .B(_0722_),
    .Y(_0723_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2073_ (.Y(\Inst_LUT4AB_switch_matrix.JW2BEG7 ),
    .B1(_0717_),
    .B2(_0723_),
    .A2(_0715_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit25.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _2074_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit22.Q ),
    .A0(A),
    .A1(B),
    .A2(C),
    .A3(D),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit23.Q ),
    .X(_0724_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _2075_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit23.Q ),
    .A0(E),
    .A1(G),
    .A2(F),
    .A3(\Inst_LUT4AB_switch_matrix.M_EF ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit22.Q ),
    .X(_0725_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _2076_ (.Y(_0726_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit24.Q ),
    .A_N(_0725_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2077_ (.B1(_0726_),
    .VDD(VPWR),
    .Y(_0727_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit24.Q ),
    .A2(_0724_));
 sg13g2_nand2b_1 _2078_ (.Y(_0728_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit22.Q ),
    .A_N(W1END[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2079_ (.B1(_0728_),
    .VDD(VPWR),
    .Y(_0729_),
    .VSS(VGND),
    .A1(W1END[0]),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit22.Q ));
 sg13g2_mux2_1 _2080_ (.A0(S1END[0]),
    .A1(S2END[0]),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit22.Q ),
    .X(_0730_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2081_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit24.Q ),
    .VDD(VPWR),
    .Y(_0731_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit23.Q ),
    .A2(_0730_));
 sg13g2_a21oi_1 _2082_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit23.Q ),
    .A2(_0729_),
    .Y(_0732_),
    .B1(_0731_));
 sg13g2_mux4_1 _2083_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit22.Q ),
    .A0(N1END[0]),
    .A1(N2END[0]),
    .A2(E1END[0]),
    .A3(EE4END[0]),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit23.Q ),
    .X(_0733_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _2084_ (.Y(_0734_),
    .B(_0733_),
    .A_N(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit24.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2085_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit25.Q ),
    .B(_0732_),
    .Y(_0735_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2086_ (.Y(\Inst_LUT4AB_switch_matrix.JN2BEG7 ),
    .B1(_0734_),
    .B2(_0735_),
    .A2(_0727_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit25.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _2087_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit22.Q ),
    .A0(A),
    .A1(B),
    .A2(C),
    .A3(D),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit23.Q ),
    .X(_0736_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _2088_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit23.Q ),
    .A0(E),
    .A1(G),
    .A2(F),
    .A3(\Inst_LUT4AB_switch_matrix.M_AH ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit22.Q ),
    .X(_0737_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _2089_ (.Y(_0738_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit24.Q ),
    .A_N(_0737_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2090_ (.B1(_0738_),
    .VDD(VPWR),
    .Y(_0739_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit24.Q ),
    .A2(_0736_));
 sg13g2_mux4_1 _2091_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit22.Q ),
    .A0(N1END[0]),
    .A1(N2END[0]),
    .A2(E1END[0]),
    .A3(E2END[0]),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit23.Q ),
    .X(_0740_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _2092_ (.Y(_0741_),
    .B(_0740_),
    .A_N(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit24.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _2093_ (.Y(_0742_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit22.Q ),
    .A_N(WW4END[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2094_ (.B1(_0742_),
    .VDD(VPWR),
    .Y(_0743_),
    .VSS(VGND),
    .A1(SS4END[0]),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit22.Q ));
 sg13g2_mux2_1 _2095_ (.A0(S1END[0]),
    .A1(S1END[2]),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit22.Q ),
    .X(_0744_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2096_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit24.Q ),
    .VDD(VPWR),
    .Y(_0745_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit23.Q ),
    .A2(_0744_));
 sg13g2_a21oi_1 _2097_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit23.Q ),
    .A2(_0743_),
    .Y(_0746_),
    .B1(_0745_));
 sg13g2_nor2_1 _2098_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit25.Q ),
    .B(_0746_),
    .Y(_0747_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2099_ (.Y(\Inst_LUT4AB_switch_matrix.E2BEG7 ),
    .B1(_0741_),
    .B2(_0747_),
    .A2(_0739_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit25.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _2100_ (.A0(\Inst_LUT4AB_switch_matrix.JN2BEG7 ),
    .A1(\Inst_LUT4AB_switch_matrix.E2BEG7 ),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit24.Q ),
    .X(_0748_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2101_ (.Y(_0749_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit24.Q ),
    .B(\Inst_LUT4AB_switch_matrix.JW2BEG7 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _2102_ (.Y(_0750_),
    .B(\Inst_LUT4AB_switch_matrix.JS2BEG7 ),
    .A_N(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit24.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2103_ (.B(_0749_),
    .C(_0750_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit25.Q ),
    .Y(_0751_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2104_ (.B1(_0751_),
    .VDD(VPWR),
    .Y(_0752_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit25.Q ),
    .A2(_0748_));
 sg13g2_mux2_1 _2105_ (.A0(_0752_),
    .A1(_0693_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit17.Q ),
    .X(_0753_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2106_ (.Y(_0754_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit16.Q ),
    .B(_0670_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2107_ (.B1(_0754_),
    .VDD(VPWR),
    .Y(_0755_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit16.Q ),
    .A2(_0753_));
 sg13g2_nor2_1 _2108_ (.A(G),
    .B(_0755_),
    .Y(_0756_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2109_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1052_),
    .A2(_0755_),
    .Y(_0757_),
    .B1(_0756_));
 sg13g2_mux2_1 _2110_ (.A0(_0757_),
    .A1(\Inst_LUT4AB_switch_matrix.M_EF ),
    .S(_0753_),
    .X(_0758_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _2111_ (.A(_0758_),
    .B_N(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit16.Q ),
    .Y(_0759_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2112_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit16.Q ),
    .B(_0757_),
    .Y(_0760_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _2113_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit17.Q ),
    .B(_0759_),
    .C(_0760_),
    .Y(_0761_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _2114_ (.A0(_0758_),
    .A1(_0697_),
    .S(_0752_),
    .X(_0762_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _2115_ (.A2(_0762_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit17.Q ),
    .B1(_0761_),
    .X(\Inst_LUT4AB_switch_matrix.M_AH ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _2116_ (.A0(A),
    .A1(B),
    .S(_0669_),
    .X(\Inst_LUT4AB_switch_matrix.M_AB ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _2117_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit27.Q ),
    .A0(B),
    .A1(D),
    .A2(C),
    .A3(E),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit26.Q ),
    .X(_0763_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _2118_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit26.Q ),
    .B_N(F),
    .Y(_0764_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2119_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit26.Q ),
    .A2(G),
    .Y(_0765_),
    .B1(_0764_));
 sg13g2_nand2_1 _2120_ (.Y(_0766_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit26.Q ),
    .B(\Inst_LUT4AB_switch_matrix.M_AD ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2121_ (.B1(_0766_),
    .VDD(VPWR),
    .Y(_0767_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit26.Q ),
    .A2(_1052_));
 sg13g2_o21ai_1 _2122_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit28.Q ),
    .VDD(VPWR),
    .Y(_0768_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit27.Q ),
    .A2(_0765_));
 sg13g2_a21oi_1 _2123_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit27.Q ),
    .A2(_0767_),
    .Y(_0769_),
    .B1(_0768_));
 sg13g2_nor2b_1 _2124_ (.A(_0769_),
    .B_N(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit29.Q ),
    .Y(_0770_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2125_ (.B1(_0770_),
    .VDD(VPWR),
    .Y(_0771_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit28.Q ),
    .A2(_0763_));
 sg13g2_mux4_1 _2126_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit27.Q ),
    .A0(N1END[3]),
    .A1(E2END[1]),
    .A2(N2END[1]),
    .A3(E6END[1]),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit26.Q ),
    .X(_0772_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _2127_ (.A0(W2END[1]),
    .A1(W6END[1]),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit26.Q ),
    .X(_0773_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _2128_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit26.Q ),
    .B_N(S2END[1]),
    .Y(_0774_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2129_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(S4END[1]),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit26.Q ),
    .Y(_0775_),
    .B1(_0774_));
 sg13g2_o21ai_1 _2130_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit28.Q ),
    .VDD(VPWR),
    .Y(_0776_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit27.Q ),
    .A2(_0775_));
 sg13g2_a21o_1 _2131_ (.A2(_0773_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit27.Q ),
    .B1(_0776_),
    .X(_0777_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2132_ (.B1(_0777_),
    .VDD(VPWR),
    .Y(_0778_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit28.Q ),
    .A2(_0772_));
 sg13g2_o21ai_1 _2133_ (.B1(_0771_),
    .VDD(VPWR),
    .Y(\Inst_LUT4AB_switch_matrix.JW2BEG0 ),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit29.Q ),
    .A2(_0778_));
 sg13g2_mux4_1 _2134_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit27.Q ),
    .A0(B),
    .A1(D),
    .A2(C),
    .A3(E),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit26.Q ),
    .X(_0779_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2135_ (.Y(_0780_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit26.Q ),
    .B(\Inst_LUT4AB_switch_matrix.M_AH ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2136_ (.B1(_0780_),
    .VDD(VPWR),
    .Y(_0781_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit26.Q ),
    .A2(_1052_));
 sg13g2_nor2b_1 _2137_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit26.Q ),
    .B_N(F),
    .Y(_0782_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2138_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit26.Q ),
    .A2(G),
    .Y(_0783_),
    .B1(_0782_));
 sg13g2_o21ai_1 _2139_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit28.Q ),
    .VDD(VPWR),
    .Y(_0784_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit27.Q ),
    .A2(_0783_));
 sg13g2_a21oi_1 _2140_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit27.Q ),
    .A2(_0781_),
    .Y(_0785_),
    .B1(_0784_));
 sg13g2_o21ai_1 _2141_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit29.Q ),
    .VDD(VPWR),
    .Y(_0786_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit28.Q ),
    .A2(_0779_));
 sg13g2_mux4_1 _2142_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit27.Q ),
    .A0(NN4END[1]),
    .A1(E2END[1]),
    .A2(E1END[3]),
    .A3(E6END[1]),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit26.Q ),
    .X(_0787_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2143_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1036_),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit26.Q ),
    .Y(_0788_),
    .B1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit27.Q ));
 sg13g2_o21ai_1 _2144_ (.B1(_0788_),
    .VDD(VPWR),
    .Y(_0789_),
    .VSS(VGND),
    .A1(S2END[1]),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit26.Q ));
 sg13g2_o21ai_1 _2145_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit27.Q ),
    .VDD(VPWR),
    .Y(_0790_),
    .VSS(VGND),
    .A1(W2END[1]),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit26.Q ));
 sg13g2_a21oi_1 _2146_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1028_),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit26.Q ),
    .Y(_0791_),
    .B1(_0790_));
 sg13g2_nor2b_1 _2147_ (.A(_0791_),
    .B_N(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit28.Q ),
    .Y(_0792_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2148_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0789_),
    .A2(_0792_),
    .Y(_0793_),
    .B1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit29.Q ));
 sg13g2_o21ai_1 _2149_ (.B1(_0793_),
    .VDD(VPWR),
    .Y(_0794_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit28.Q ),
    .A2(_0787_));
 sg13g2_o21ai_1 _2150_ (.B1(_0794_),
    .VDD(VPWR),
    .Y(\Inst_LUT4AB_switch_matrix.JS2BEG0 ),
    .VSS(VGND),
    .A1(_0785_),
    .A2(_0786_));
 sg13g2_nor2b_1 _2151_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit26.Q ),
    .B_N(F),
    .Y(_0795_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2152_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit26.Q ),
    .A2(G),
    .Y(_0796_),
    .B1(_0795_));
 sg13g2_nand2_1 _2153_ (.Y(_0797_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit26.Q ),
    .B(\Inst_LUT4AB_switch_matrix.M_EF ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2154_ (.B1(_0797_),
    .VDD(VPWR),
    .Y(_0798_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit26.Q ),
    .A2(_1052_));
 sg13g2_o21ai_1 _2155_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit28.Q ),
    .VDD(VPWR),
    .Y(_0799_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit27.Q ),
    .A2(_0796_));
 sg13g2_a21o_1 _2156_ (.A2(_0798_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit27.Q ),
    .B1(_0799_),
    .X(_0800_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _2157_ (.A0(D),
    .A1(E),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit26.Q ),
    .X(_0801_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _2158_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit26.Q ),
    .B_N(B),
    .Y(_0802_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2159_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit26.Q ),
    .A2(C),
    .Y(_0803_),
    .B1(_0802_));
 sg13g2_a21oi_1 _2160_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit27.Q ),
    .A2(_0801_),
    .Y(_0804_),
    .B1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit28.Q ));
 sg13g2_o21ai_1 _2161_ (.B1(_0804_),
    .VDD(VPWR),
    .Y(_0805_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit27.Q ),
    .A2(_0803_));
 sg13g2_nand3_1 _2162_ (.B(_0800_),
    .C(_0805_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit29.Q ),
    .Y(_0806_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _2163_ (.A0(N4END[1]),
    .A1(EE4END[1]),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit26.Q ),
    .X(_0807_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _2164_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit26.Q ),
    .B_N(N1END[3]),
    .Y(_0808_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2165_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(N2END[1]),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit26.Q ),
    .Y(_0809_),
    .B1(_0808_));
 sg13g2_a21oi_1 _2166_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit27.Q ),
    .A2(_0807_),
    .Y(_0810_),
    .B1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit28.Q ));
 sg13g2_o21ai_1 _2167_ (.B1(_0810_),
    .VDD(VPWR),
    .Y(_0811_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit27.Q ),
    .A2(_0809_));
 sg13g2_nor2b_1 _2168_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit26.Q ),
    .B_N(E6END[1]),
    .Y(_0812_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2169_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(S2END[1]),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit26.Q ),
    .Y(_0813_),
    .B1(_0812_));
 sg13g2_mux2_1 _2170_ (.A0(W2END[1]),
    .A1(W6END[1]),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit26.Q ),
    .X(_0814_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2171_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit28.Q ),
    .VDD(VPWR),
    .Y(_0815_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit27.Q ),
    .A2(_0813_));
 sg13g2_a21oi_1 _2172_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit27.Q ),
    .A2(_0814_),
    .Y(_0816_),
    .B1(_0815_));
 sg13g2_nand2b_1 _2173_ (.Y(_0817_),
    .B(_0811_),
    .A_N(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit29.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2174_ (.B1(_0806_),
    .VDD(VPWR),
    .Y(\Inst_LUT4AB_switch_matrix.E2BEG0 ),
    .VSS(VGND),
    .A1(_0816_),
    .A2(_0817_));
 sg13g2_mux4_1 _2175_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit27.Q ),
    .A0(B),
    .A1(D),
    .A2(C),
    .A3(E),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit26.Q ),
    .X(_0818_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _2176_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit26.Q ),
    .B_N(F),
    .Y(_0819_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2177_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit26.Q ),
    .A2(G),
    .Y(_0820_),
    .B1(_0819_));
 sg13g2_nand2_1 _2178_ (.Y(_0821_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit26.Q ),
    .B(\Inst_LUT4AB_switch_matrix.M_AB ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2179_ (.B1(_0821_),
    .VDD(VPWR),
    .Y(_0822_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit26.Q ),
    .A2(_1052_));
 sg13g2_o21ai_1 _2180_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit28.Q ),
    .VDD(VPWR),
    .Y(_0823_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit27.Q ),
    .A2(_0820_));
 sg13g2_a21oi_1 _2181_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit27.Q ),
    .A2(_0822_),
    .Y(_0824_),
    .B1(_0823_));
 sg13g2_nor2b_1 _2182_ (.A(_0824_),
    .B_N(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit29.Q ),
    .Y(_0825_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2183_ (.B1(_0825_),
    .VDD(VPWR),
    .Y(_0826_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit28.Q ),
    .A2(_0818_));
 sg13g2_mux2_1 _2184_ (.A0(E1END[3]),
    .A1(E2END[1]),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit26.Q ),
    .X(_0827_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _2185_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit26.Q ),
    .B_N(N2END[1]),
    .Y(_0828_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2186_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(N4END[1]),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit26.Q ),
    .Y(_0829_),
    .B1(_0828_));
 sg13g2_a21oi_1 _2187_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit27.Q ),
    .A2(_0827_),
    .Y(_0830_),
    .B1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit28.Q ));
 sg13g2_o21ai_1 _2188_ (.B1(_0830_),
    .VDD(VPWR),
    .Y(_0831_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit27.Q ),
    .A2(_0829_));
 sg13g2_o21ai_1 _2189_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit27.Q ),
    .VDD(VPWR),
    .Y(_0832_),
    .VSS(VGND),
    .A1(W2END[1]),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit26.Q ));
 sg13g2_a21oi_1 _2190_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1028_),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit26.Q ),
    .Y(_0833_),
    .B1(_0832_));
 sg13g2_nor2b_1 _2191_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit26.Q ),
    .B_N(E6END[1]),
    .Y(_0834_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2192_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(SS4END[1]),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit26.Q ),
    .Y(_0835_),
    .B1(_0834_));
 sg13g2_o21ai_1 _2193_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit28.Q ),
    .VDD(VPWR),
    .Y(_0836_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit27.Q ),
    .A2(_0835_));
 sg13g2_o21ai_1 _2194_ (.B1(_0831_),
    .VDD(VPWR),
    .Y(_0837_),
    .VSS(VGND),
    .A1(_0833_),
    .A2(_0836_));
 sg13g2_o21ai_1 _2195_ (.B1(_0826_),
    .VDD(VPWR),
    .Y(\Inst_LUT4AB_switch_matrix.JN2BEG0 ),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit29.Q ),
    .A2(_0837_));
 sg13g2_mux4_1 _2196_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit30.Q ),
    .A0(_1158_),
    .A1(_0196_),
    .A2(_0276_),
    .A3(_0556_),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit31.Q ),
    .X(_0838_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _2197_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit30.Q ),
    .A0(G),
    .A1(H),
    .A2(\Inst_LUT4AB_switch_matrix.M_AD ),
    .A3(\Inst_LUT4AB_switch_matrix.M_EF ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit31.Q ),
    .X(_0839_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2198_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit1.Q ),
    .VDD(VPWR),
    .Y(_0840_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit0.Q ),
    .A2(_0839_));
 sg13g2_a21oi_1 _2199_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit0.Q ),
    .A2(_0838_),
    .Y(_0841_),
    .B1(_0840_));
 sg13g2_mux4_1 _2200_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit30.Q ),
    .A0(E1END[2]),
    .A1(W1END[2]),
    .A2(A),
    .A3(B),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit31.Q ),
    .X(_0842_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _2201_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit30.Q ),
    .A0(C),
    .A1(D),
    .A2(E),
    .A3(F),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit31.Q ),
    .X(_0843_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _2202_ (.VDD(VPWR),
    .Y(_0844_),
    .A(_0843_),
    .VSS(VGND));
 sg13g2_a21oi_1 _2203_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit0.Q ),
    .A2(_0844_),
    .Y(_0845_),
    .B1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit1.Q ));
 sg13g2_o21ai_1 _2204_ (.B1(_0845_),
    .VDD(VPWR),
    .Y(_0846_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit0.Q ),
    .A2(_0842_));
 sg13g2_nand2b_1 _2205_ (.Y(\Inst_LUT4AB_switch_matrix.W6BEG1 ),
    .B(_0846_),
    .A_N(_0841_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _2206_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit26.Q ),
    .A0(E1END[3]),
    .A1(W1END[3]),
    .A2(A),
    .A3(B),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit27.Q ),
    .X(_0847_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _2207_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit26.Q ),
    .A0(C),
    .A1(D),
    .A2(E),
    .A3(F),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit27.Q ),
    .X(_0848_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _2208_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit26.Q ),
    .A0(G),
    .A1(H),
    .A2(\Inst_LUT4AB_switch_matrix.M_AB ),
    .A3(\Inst_LUT4AB_switch_matrix.M_AH ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit27.Q ),
    .X(_0849_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _2209_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit26.Q ),
    .A0(_1084_),
    .A1(_0148_),
    .A2(_0308_),
    .A3(_0586_),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit27.Q ),
    .X(_0850_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _2210_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit28.Q ),
    .A0(_0847_),
    .A1(_0848_),
    .A2(_0849_),
    .A3(_0850_),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit29.Q ),
    .X(\Inst_LUT4AB_switch_matrix.W6BEG0 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _2211_ (.A0(N1END[1]),
    .A1(S1END[1]),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit23.Q ),
    .X(_0851_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _2212_ (.A0(W1END[1]),
    .A1(D),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit23.Q ),
    .X(_0852_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2213_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit23.Q ),
    .B(E),
    .Y(_0853_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2214_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit23.Q ),
    .A2(_0276_),
    .Y(_0854_),
    .B1(_0853_));
 sg13g2_nand2_1 _2215_ (.Y(_0855_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit23.Q ),
    .B(_1141_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2216_ (.B1(_0855_),
    .VDD(VPWR),
    .Y(_0856_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit23.Q ),
    .A2(_0556_));
 sg13g2_mux4_1 _2217_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit24.Q ),
    .A0(_0851_),
    .A1(_0852_),
    .A2(_0854_),
    .A3(_0856_),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit25.Q ),
    .X(\Inst_LUT4AB_switch_matrix.WW4BEG3 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2218_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit21.Q ),
    .VDD(VPWR),
    .Y(_0857_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit20.Q ),
    .A2(_0586_));
 sg13g2_a21oi_1 _2219_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit20.Q ),
    .A2(_0171_),
    .Y(_0858_),
    .B1(_0857_));
 sg13g2_nor2b_1 _2220_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit20.Q ),
    .B_N(C),
    .Y(_0859_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2221_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit20.Q ),
    .A2(_0308_),
    .Y(_0860_),
    .B1(_0859_));
 sg13g2_o21ai_1 _2222_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit22.Q ),
    .VDD(VPWR),
    .Y(_0861_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit21.Q ),
    .A2(_0860_));
 sg13g2_nor2_1 _2223_ (.A(_0858_),
    .B(_0861_),
    .Y(_0862_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _2224_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit21.Q ),
    .A0(N1END[0]),
    .A1(W1END[0]),
    .A2(S1END[0]),
    .A3(B),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit20.Q ),
    .X(_0863_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2225_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit22.Q ),
    .B(_0863_),
    .Y(_0864_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2226_ (.A(_0862_),
    .B(_0864_),
    .Y(\Inst_LUT4AB_switch_matrix.WW4BEG2 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _2227_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit17.Q ),
    .A0(_1052_),
    .A1(_1158_),
    .A2(_0196_),
    .A3(_0253_),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit18.Q ),
    .X(_0865_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _2228_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit17.Q ),
    .A0(N1END[3]),
    .A1(S1END[3]),
    .A2(W1END[3]),
    .A3(A),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit18.Q ),
    .X(_0866_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2229_ (.Y(_0867_),
    .A(_1048_),
    .B(_0866_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2230_ (.B1(_0867_),
    .VDD(VPWR),
    .Y(\Inst_LUT4AB_switch_matrix.WW4BEG1 ),
    .VSS(VGND),
    .A1(_1048_),
    .A2(_0865_));
 sg13g2_mux4_1 _2231_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit14.Q ),
    .A0(N1END[2]),
    .A1(S1END[2]),
    .A2(W1END[2]),
    .A3(F),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit15.Q ),
    .X(_0868_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _2232_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit14.Q ),
    .A0(G),
    .A1(_1084_),
    .A2(_0148_),
    .A3(_0538_),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit15.Q ),
    .X(_0869_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _2233_ (.A0(_0868_),
    .A1(_0869_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit16.Q ),
    .X(\Inst_LUT4AB_switch_matrix.WW4BEG0 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _2234_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit3.Q ),
    .A0(N1END[1]),
    .A1(E1END[1]),
    .A2(W1END[1]),
    .A3(D),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit4.Q ),
    .X(_0870_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2235_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit5.Q ),
    .B(_0870_),
    .Y(_0871_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2236_ (.Y(_0872_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit3.Q ),
    .B(_0276_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2237_ (.B1(_0872_),
    .VDD(VPWR),
    .Y(_0873_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit3.Q ),
    .A2(E));
 sg13g2_nand2_1 _2238_ (.Y(_0874_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit3.Q ),
    .B(_0023_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2239_ (.B1(_0874_),
    .VDD(VPWR),
    .Y(_0875_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit3.Q ),
    .A2(_0556_));
 sg13g2_o21ai_1 _2240_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit5.Q ),
    .VDD(VPWR),
    .Y(_0876_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit4.Q ),
    .A2(_0873_));
 sg13g2_a21oi_1 _2241_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit4.Q ),
    .A2(_0875_),
    .Y(_0877_),
    .B1(_0876_));
 sg13g2_nor2_1 _2242_ (.A(_0871_),
    .B(_0877_),
    .Y(\Inst_LUT4AB_switch_matrix.SS4BEG3 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2243_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit1.Q ),
    .VDD(VPWR),
    .Y(_0878_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit0.Q ),
    .A2(_0586_));
 sg13g2_a21oi_1 _2244_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit0.Q ),
    .A2(_0430_),
    .Y(_0879_),
    .B1(_0878_));
 sg13g2_nor2b_1 _2245_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit0.Q ),
    .B_N(C),
    .Y(_0880_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2246_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit0.Q ),
    .A2(_0308_),
    .Y(_0881_),
    .B1(_0880_));
 sg13g2_o21ai_1 _2247_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit2.Q ),
    .VDD(VPWR),
    .Y(_0882_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit1.Q ),
    .A2(_0881_));
 sg13g2_nor2_1 _2248_ (.A(_0879_),
    .B(_0882_),
    .Y(_0883_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _2249_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit1.Q ),
    .A0(N1END[0]),
    .A1(W1END[0]),
    .A2(E1END[0]),
    .A3(B),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit0.Q ),
    .X(_0884_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2250_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit2.Q ),
    .B(_0884_),
    .Y(_0885_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2251_ (.A(_0883_),
    .B(_0885_),
    .Y(\Inst_LUT4AB_switch_matrix.SS4BEG2 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _2252_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit29.Q ),
    .A0(N1END[3]),
    .A1(E1END[3]),
    .A2(W1END[3]),
    .A3(A),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit30.Q ),
    .X(_0886_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2253_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit31.Q ),
    .B(_0886_),
    .Y(_0887_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _2254_ (.A0(_0197_),
    .A1(_0316_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit29.Q ),
    .X(_0888_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2255_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit29.Q ),
    .B(_1052_),
    .Y(_0889_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2256_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit29.Q ),
    .A2(_1157_),
    .Y(_0890_),
    .B1(_0889_));
 sg13g2_o21ai_1 _2257_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit31.Q ),
    .VDD(VPWR),
    .Y(_0891_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit30.Q ),
    .A2(_0890_));
 sg13g2_a21oi_1 _2258_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit30.Q ),
    .A2(_0888_),
    .Y(_0892_),
    .B1(_0891_));
 sg13g2_nor2_1 _2259_ (.A(_0887_),
    .B(_0892_),
    .Y(\Inst_LUT4AB_switch_matrix.SS4BEG1 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2260_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit27.Q ),
    .VDD(VPWR),
    .Y(_0893_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit26.Q ),
    .A2(_0148_));
 sg13g2_a21oi_1 _2261_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit26.Q ),
    .A2(_0626_),
    .Y(_0894_),
    .B1(_0893_));
 sg13g2_nor2b_1 _2262_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit26.Q ),
    .B_N(G),
    .Y(_0895_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2263_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit26.Q ),
    .A2(_1084_),
    .Y(_0896_),
    .B1(_0895_));
 sg13g2_o21ai_1 _2264_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit28.Q ),
    .VDD(VPWR),
    .Y(_0897_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit27.Q ),
    .A2(_0896_));
 sg13g2_nor2_1 _2265_ (.A(_0894_),
    .B(_0897_),
    .Y(_0898_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _2266_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit27.Q ),
    .A0(N1END[2]),
    .A1(W1END[2]),
    .A2(E1END[2]),
    .A3(F),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit26.Q ),
    .X(_0899_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2267_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit28.Q ),
    .B(_0899_),
    .Y(_0900_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2268_ (.A(_0898_),
    .B(_0900_),
    .Y(\Inst_LUT4AB_switch_matrix.SS4BEG0 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2269_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(W1END[2]),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit6.Q ),
    .Y(_0901_),
    .B1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit7.Q ));
 sg13g2_o21ai_1 _2270_ (.B1(_0901_),
    .VDD(VPWR),
    .Y(_0902_),
    .VSS(VGND),
    .A1(_1013_),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit6.Q ));
 sg13g2_nor2b_1 _2271_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit6.Q ),
    .B_N(A),
    .Y(_0903_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2272_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit6.Q ),
    .A2(B),
    .Y(_0904_),
    .B1(_0903_));
 sg13g2_a21oi_1 _2273_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit7.Q ),
    .A2(_0904_),
    .Y(_0905_),
    .B1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit8.Q ));
 sg13g2_mux4_1 _2274_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit6.Q ),
    .A0(C),
    .A1(D),
    .A2(E),
    .A3(F),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit7.Q ),
    .X(_0906_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _2275_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit8.Q ),
    .C1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit9.Q ),
    .B1(_0906_),
    .A1(_0902_),
    .Y(_0907_),
    .A2(_0905_));
 sg13g2_mux4_1 _2276_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit6.Q ),
    .A0(_1158_),
    .A1(_0196_),
    .A2(_0276_),
    .A3(_0556_),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit7.Q ),
    .X(_0908_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _2277_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit6.Q ),
    .A0(G),
    .A1(H),
    .A2(\Inst_LUT4AB_switch_matrix.M_AD ),
    .A3(\Inst_LUT4AB_switch_matrix.M_EF ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit7.Q ),
    .X(_0909_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2278_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit9.Q ),
    .VDD(VPWR),
    .Y(_0910_),
    .VSS(VGND),
    .A1(_1049_),
    .A2(_0908_));
 sg13g2_a21oi_1 _2279_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1049_),
    .A2(_0909_),
    .Y(_0911_),
    .B1(_0910_));
 sg13g2_nor2_1 _2280_ (.A(_0907_),
    .B(_0911_),
    .Y(\Inst_LUT4AB_switch_matrix.E6BEG1 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _2281_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit2.Q ),
    .A0(E1END[3]),
    .A1(W1END[3]),
    .A2(A),
    .A3(B),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit3.Q ),
    .X(_0912_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _2282_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit2.Q ),
    .A0(C),
    .A1(D),
    .A2(E),
    .A3(F),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit3.Q ),
    .X(_0913_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _2283_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit2.Q ),
    .A0(G),
    .A1(H),
    .A2(\Inst_LUT4AB_switch_matrix.M_AB ),
    .A3(\Inst_LUT4AB_switch_matrix.M_AH ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit3.Q ),
    .X(_0914_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _2284_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit2.Q ),
    .A0(_1084_),
    .A1(_0148_),
    .A2(_0308_),
    .A3(_0586_),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit3.Q ),
    .X(_0915_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _2285_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit4.Q ),
    .A0(_0912_),
    .A1(_0913_),
    .A2(_0914_),
    .A3(_0915_),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit5.Q ),
    .X(\Inst_LUT4AB_switch_matrix.E6BEG0 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _2286_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit31.Q ),
    .A0(N1END[1]),
    .A1(E1END[1]),
    .A2(S1END[1]),
    .A3(D),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit0.Q ),
    .X(_0916_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2287_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit1.Q ),
    .B(_0916_),
    .Y(_0917_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2288_ (.Y(_0918_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit31.Q ),
    .B(_1119_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2289_ (.B1(_0918_),
    .VDD(VPWR),
    .Y(_0919_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit31.Q ),
    .A2(_0556_));
 sg13g2_nand2_1 _2290_ (.Y(_0920_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit31.Q ),
    .B(_0276_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2291_ (.B1(_0920_),
    .VDD(VPWR),
    .Y(_0921_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit31.Q ),
    .A2(E));
 sg13g2_o21ai_1 _2292_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit1.Q ),
    .VDD(VPWR),
    .Y(_0922_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit0.Q ),
    .A2(_0921_));
 sg13g2_a21oi_1 _2293_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit0.Q ),
    .A2(_0919_),
    .Y(_0923_),
    .B1(_0922_));
 sg13g2_nor2_1 _2294_ (.A(_0917_),
    .B(_0923_),
    .Y(\Inst_LUT4AB_switch_matrix.EE4BEG3 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _2295_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit28.Q ),
    .A0(C),
    .A1(_0308_),
    .A2(_0586_),
    .A3(_0366_),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit29.Q ),
    .X(_0924_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _2296_ (.VDD(VPWR),
    .Y(_0925_),
    .A(_0924_),
    .VSS(VGND));
 sg13g2_a21oi_1 _2297_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1016_),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit28.Q ),
    .Y(_0926_),
    .B1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit29.Q ));
 sg13g2_o21ai_1 _2298_ (.B1(_0926_),
    .VDD(VPWR),
    .Y(_0927_),
    .VSS(VGND),
    .A1(N1END[0]),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit28.Q ));
 sg13g2_mux2_1 _2299_ (.A0(S1END[0]),
    .A1(B),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit28.Q ),
    .X(_0928_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2300_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit29.Q ),
    .A2(_0928_),
    .Y(_0929_),
    .B1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit30.Q ));
 sg13g2_a22oi_1 _2301_ (.Y(\Inst_LUT4AB_switch_matrix.EE4BEG2 ),
    .B1(_0927_),
    .B2(_0929_),
    .A2(_0925_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit30.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _2302_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit25.Q ),
    .A0(H),
    .A1(_1157_),
    .A2(_0197_),
    .A3(_0239_),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit26.Q ),
    .X(_0930_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _2303_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit25.Q ),
    .A0(N1END[3]),
    .A1(E1END[3]),
    .A2(S1END[3]),
    .A3(A),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit26.Q ),
    .X(_0931_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _2304_ (.A0(_0931_),
    .A1(_0930_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit27.Q ),
    .X(\Inst_LUT4AB_switch_matrix.EE4BEG1 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2305_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit23.Q ),
    .VDD(VPWR),
    .Y(_0932_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit22.Q ),
    .A2(_0148_));
 sg13g2_a21oi_1 _2306_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit22.Q ),
    .A2(_0529_),
    .Y(_0933_),
    .B1(_0932_));
 sg13g2_nor2b_1 _2307_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit22.Q ),
    .B_N(G),
    .Y(_0934_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2308_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit22.Q ),
    .A2(_1084_),
    .Y(_0935_),
    .B1(_0934_));
 sg13g2_o21ai_1 _2309_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit24.Q ),
    .VDD(VPWR),
    .Y(_0936_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit23.Q ),
    .A2(_0935_));
 sg13g2_nor2_1 _2310_ (.A(_0933_),
    .B(_0936_),
    .Y(_0937_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _2311_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit23.Q ),
    .A0(N1END[2]),
    .A1(S1END[2]),
    .A2(E1END[2]),
    .A3(F),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit22.Q ),
    .X(_0938_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2312_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit24.Q ),
    .B(_0938_),
    .Y(_0939_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2313_ (.A(_0937_),
    .B(_0939_),
    .Y(\Inst_LUT4AB_switch_matrix.EE4BEG0 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _2314_ (.A0(N1END[1]),
    .A1(E1END[1]),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit11.Q ),
    .X(_0940_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _2315_ (.A0(W1END[1]),
    .A1(D),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit11.Q ),
    .X(_0941_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2316_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit11.Q ),
    .B(E),
    .Y(_0942_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2317_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit11.Q ),
    .A2(_0276_),
    .Y(_0943_),
    .B1(_0942_));
 sg13g2_nand2_1 _2318_ (.Y(_0944_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit11.Q ),
    .B(_1066_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2319_ (.B1(_0944_),
    .VDD(VPWR),
    .Y(_0945_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit11.Q ),
    .A2(_0556_));
 sg13g2_mux4_1 _2320_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit12.Q ),
    .A0(_0940_),
    .A1(_0941_),
    .A2(_0943_),
    .A3(_0945_),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit13.Q ),
    .X(\Inst_LUT4AB_switch_matrix.NN4BEG3 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _2321_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0946_),
    .B(_0586_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit8.Q ));
 sg13g2_nand2b_1 _2322_ (.Y(_0947_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit8.Q ),
    .A_N(_0130_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2323_ (.B(_0946_),
    .C(_0947_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit9.Q ),
    .Y(_0948_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _2324_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit8.Q ),
    .B_N(C),
    .Y(_0949_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2325_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit8.Q ),
    .A2(_0308_),
    .Y(_0950_),
    .B1(_0949_));
 sg13g2_o21ai_1 _2326_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit10.Q ),
    .VDD(VPWR),
    .Y(_0951_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit9.Q ),
    .A2(_0950_));
 sg13g2_inv_1 _2327_ (.VDD(VPWR),
    .Y(_0952_),
    .A(_0951_),
    .VSS(VGND));
 sg13g2_mux4_1 _2328_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit9.Q ),
    .A0(N1END[0]),
    .A1(W1END[0]),
    .A2(E1END[0]),
    .A3(B),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit8.Q ),
    .X(_0953_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2329_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit10.Q ),
    .B(_0953_),
    .Y(_0954_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2330_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0948_),
    .A2(_0952_),
    .Y(\Inst_LUT4AB_switch_matrix.NN4BEG2 ),
    .B1(_0954_));
 sg13g2_mux4_1 _2331_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit5.Q ),
    .A0(_1052_),
    .A1(_1158_),
    .A2(_0196_),
    .A3(_0290_),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit6.Q ),
    .X(_0955_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _2332_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit5.Q ),
    .A0(N1END[3]),
    .A1(E1END[3]),
    .A2(W1END[3]),
    .A3(A),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit6.Q ),
    .X(_0956_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2333_ (.Y(_0957_),
    .A(_1050_),
    .B(_0956_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2334_ (.B1(_0957_),
    .VDD(VPWR),
    .Y(\Inst_LUT4AB_switch_matrix.NN4BEG1 ),
    .VSS(VGND),
    .A1(_1050_),
    .A2(_0955_));
 sg13g2_o21ai_1 _2335_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit3.Q ),
    .VDD(VPWR),
    .Y(_0958_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit2.Q ),
    .A2(_0148_));
 sg13g2_a21oi_1 _2336_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit2.Q ),
    .A2(_0589_),
    .Y(_0959_),
    .B1(_0958_));
 sg13g2_nor2b_1 _2337_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit2.Q ),
    .B_N(G),
    .Y(_0960_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2338_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit2.Q ),
    .A2(_1084_),
    .Y(_0961_),
    .B1(_0960_));
 sg13g2_o21ai_1 _2339_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit4.Q ),
    .VDD(VPWR),
    .Y(_0962_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit3.Q ),
    .A2(_0961_));
 sg13g2_nor2_1 _2340_ (.A(_0959_),
    .B(_0962_),
    .Y(_0963_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _2341_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit3.Q ),
    .A0(N1END[2]),
    .A1(W1END[2]),
    .A2(E1END[2]),
    .A3(F),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit2.Q ),
    .X(_0964_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2342_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit4.Q ),
    .B(_0964_),
    .Y(_0965_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2343_ (.A(_0963_),
    .B(_0965_),
    .Y(\Inst_LUT4AB_switch_matrix.NN4BEG0 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _2344_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit12.Q ),
    .A0(A),
    .A1(_1159_),
    .A2(\Inst_LUT4AB_switch_matrix.JS2BEG2 ),
    .A3(_1118_),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit13.Q ),
    .X(\Inst_LUT4AB_switch_matrix.W1BEG3 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _2345_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit11.Q ),
    .A0(H),
    .A1(\Inst_LUT4AB_switch_matrix.JS2BEG1 ),
    .A2(_0586_),
    .A3(_0623_),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit10.Q ),
    .X(\Inst_LUT4AB_switch_matrix.W1BEG2 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _2346_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit8.Q ),
    .A0(G),
    .A1(_0237_),
    .A2(\Inst_LUT4AB_switch_matrix.JS2BEG0 ),
    .A3(_0248_),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit9.Q ),
    .X(\Inst_LUT4AB_switch_matrix.W1BEG1 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _2347_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit7.Q ),
    .A0(F),
    .A1(\Inst_LUT4AB_switch_matrix.JS2BEG3 ),
    .A2(_0453_),
    .A3(_0129_),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit6.Q ),
    .X(\Inst_LUT4AB_switch_matrix.W1BEG0 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _2348_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit24.Q ),
    .A0(S2END[1]),
    .A1(S4END[0]),
    .A2(W6END[0]),
    .A3(D),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit25.Q ),
    .X(\Inst_LUT4AB_switch_matrix.S4BEG3 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _2349_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit23.Q ),
    .A0(S2END[0]),
    .A1(W6END[1]),
    .A2(S4END[3]),
    .A3(C),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit22.Q ),
    .X(\Inst_LUT4AB_switch_matrix.S4BEG2 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _2350_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit21.Q ),
    .A0(E6END[0]),
    .A1(S4END[2]),
    .A2(S2END[3]),
    .A3(B),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit20.Q ),
    .X(\Inst_LUT4AB_switch_matrix.S4BEG1 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _2351_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit19.Q ),
    .A0(E6END[1]),
    .A1(S4END[1]),
    .A2(S2END[2]),
    .A3(A),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit18.Q ),
    .X(\Inst_LUT4AB_switch_matrix.S4BEG0 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _2352_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit16.Q ),
    .A0(H),
    .A1(_1159_),
    .A2(\Inst_LUT4AB_switch_matrix.E2BEG2 ),
    .A3(_1118_),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit17.Q ),
    .X(\Inst_LUT4AB_switch_matrix.S1BEG3 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _2353_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit15.Q ),
    .A0(G),
    .A1(\Inst_LUT4AB_switch_matrix.E2BEG1 ),
    .A2(_0586_),
    .A3(_0623_),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit14.Q ),
    .X(\Inst_LUT4AB_switch_matrix.S1BEG2 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _2354_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit12.Q ),
    .A0(F),
    .A1(_0237_),
    .A2(\Inst_LUT4AB_switch_matrix.E2BEG0 ),
    .A3(_0248_),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit13.Q ),
    .X(\Inst_LUT4AB_switch_matrix.S1BEG1 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _2355_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit11.Q ),
    .A0(E),
    .A1(\Inst_LUT4AB_switch_matrix.E2BEG3 ),
    .A2(_0453_),
    .A3(_0129_),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit10.Q ),
    .X(\Inst_LUT4AB_switch_matrix.S1BEG0 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _2356_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit20.Q ),
    .A0(G),
    .A1(_1159_),
    .A2(\Inst_LUT4AB_switch_matrix.JN2BEG2 ),
    .A3(_1118_),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit21.Q ),
    .X(\Inst_LUT4AB_switch_matrix.E1BEG3 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _2357_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit19.Q ),
    .A0(F),
    .A1(\Inst_LUT4AB_switch_matrix.JN2BEG1 ),
    .A2(_0586_),
    .A3(_0623_),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit18.Q ),
    .X(\Inst_LUT4AB_switch_matrix.E1BEG2 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _2358_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit16.Q ),
    .A0(E),
    .A1(_0237_),
    .A2(\Inst_LUT4AB_switch_matrix.JN2BEG0 ),
    .A3(_0248_),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit17.Q ),
    .X(\Inst_LUT4AB_switch_matrix.E1BEG1 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _2359_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit15.Q ),
    .A0(D),
    .A1(\Inst_LUT4AB_switch_matrix.JN2BEG3 ),
    .A2(_0453_),
    .A3(_0129_),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit14.Q ),
    .X(\Inst_LUT4AB_switch_matrix.E1BEG0 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _2360_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit1.Q ),
    .A0(N2END[1]),
    .A1(W6END[0]),
    .A2(N4END[0]),
    .A3(H),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit0.Q ),
    .X(\Inst_LUT4AB_switch_matrix.N4BEG3 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _2361_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit30.Q ),
    .A0(N2END[0]),
    .A1(N4END[3]),
    .A2(W6END[1]),
    .A3(G),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit31.Q ),
    .X(\Inst_LUT4AB_switch_matrix.N4BEG2 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _2362_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit28.Q ),
    .A0(N2END[3]),
    .A1(N4END[2]),
    .A2(E6END[0]),
    .A3(F),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit29.Q ),
    .X(\Inst_LUT4AB_switch_matrix.N4BEG1 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _2363_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit26.Q ),
    .A0(N2END[2]),
    .A1(N4END[1]),
    .A2(E6END[1]),
    .A3(E),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit27.Q ),
    .X(\Inst_LUT4AB_switch_matrix.N4BEG0 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _2364_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit24.Q ),
    .A0(F),
    .A1(_1159_),
    .A2(\Inst_LUT4AB_switch_matrix.JW2BEG2 ),
    .A3(_1118_),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit25.Q ),
    .X(\Inst_LUT4AB_switch_matrix.N1BEG3 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _2365_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit23.Q ),
    .A0(E),
    .A1(\Inst_LUT4AB_switch_matrix.JW2BEG1 ),
    .A2(_0586_),
    .A3(_0623_),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit22.Q ),
    .X(\Inst_LUT4AB_switch_matrix.N1BEG2 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _2366_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit20.Q ),
    .A0(D),
    .A1(_0237_),
    .A2(\Inst_LUT4AB_switch_matrix.JW2BEG0 ),
    .A3(_0248_),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit21.Q ),
    .X(\Inst_LUT4AB_switch_matrix.N1BEG1 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _2367_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit19.Q ),
    .A0(C),
    .A1(\Inst_LUT4AB_switch_matrix.JW2BEG3 ),
    .A2(_0453_),
    .A3(_0129_),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit18.Q ),
    .X(\Inst_LUT4AB_switch_matrix.N1BEG0 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2368_ (.B1(_0651_),
    .VDD(VPWR),
    .Y(Co),
    .VSS(VGND),
    .A1(_0639_),
    .A2(_0652_));
 sg13g2_nand2b_1 _2369_ (.Y(_0966_),
    .B(_0617_),
    .A_N(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit29.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2370_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit29.Q ),
    .A2(_0048_),
    .Y(_0967_),
    .B1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit30.Q ));
 sg13g2_nor2_1 _2371_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit29.Q ),
    .B(_0453_),
    .Y(_0968_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2372_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit29.Q ),
    .A2(_0334_),
    .Y(_0969_),
    .B1(_0968_));
 sg13g2_mux4_1 _2373_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit30.Q ),
    .A0(\Inst_LUT4AB_switch_matrix.JN2BEG2 ),
    .A1(\Inst_LUT4AB_switch_matrix.JS2BEG2 ),
    .A2(\Inst_LUT4AB_switch_matrix.E2BEG2 ),
    .A3(\Inst_LUT4AB_switch_matrix.JW2BEG2 ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit29.Q ),
    .X(_0970_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2374_ (.Y(_0971_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit31.Q ),
    .B(_0970_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2375_ (.Y(_0972_),
    .B1(_0969_),
    .B2(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit30.Q ),
    .A2(_0967_),
    .A1(_0966_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2376_ (.B1(_0971_),
    .VDD(VPWR),
    .Y(_0973_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit31.Q ),
    .A2(_0972_));
 sg13g2_nand2b_1 _2377_ (.Y(_0974_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit17.Q ),
    .A_N(_0973_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3b_1 _2378_ (.B(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit17.Q ),
    .C(\Inst_LH_LUT4c_frame_config_dffesr.LUT_flop ),
    .Y(_0975_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(_0973_));
 sg13g2_nand2b_1 _2379_ (.Y(_0976_),
    .B(_0520_),
    .A_N(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit26.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2380_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit26.Q ),
    .A2(_1104_),
    .Y(_0977_),
    .B1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit27.Q ));
 sg13g2_mux2_1 _2381_ (.A0(_0390_),
    .A1(_0237_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit26.Q ),
    .X(_0978_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _2382_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit27.Q ),
    .C1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit28.Q ),
    .B1(_0978_),
    .A1(_0976_),
    .Y(_0979_),
    .A2(_0977_));
 sg13g2_o21ai_1 _2383_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit27.Q ),
    .VDD(VPWR),
    .Y(_0980_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit26.Q ),
    .A2(\Inst_LUT4AB_switch_matrix.JS2BEG1 ));
 sg13g2_a21oi_1 _2384_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit26.Q ),
    .A2(_0021_),
    .Y(_0981_),
    .B1(_0980_));
 sg13g2_a21oi_1 _2385_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit26.Q ),
    .A2(_1064_),
    .Y(_0982_),
    .B1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit27.Q ));
 sg13g2_o21ai_1 _2386_ (.B1(_0982_),
    .VDD(VPWR),
    .Y(_0983_),
    .VSS(VGND),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit26.Q ),
    .A2(\Inst_LUT4AB_switch_matrix.JN2BEG1 ));
 sg13g2_nor2b_1 _2387_ (.A(_0981_),
    .B_N(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit28.Q ),
    .Y(_0984_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2388_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0983_),
    .A2(_0984_),
    .Y(_0985_),
    .B1(_0979_));
 sg13g2_nand2_1 _2389_ (.Y(_0986_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit16.Q ),
    .B(_0985_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _2390_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit16.Q ),
    .C1(_0659_),
    .B1(_0985_),
    .A1(_0661_),
    .Y(_0987_),
    .A2(_0665_));
 sg13g2_o21ai_1 _2391_ (.B1(_0974_),
    .VDD(VPWR),
    .Y(_0988_),
    .VSS(VGND),
    .A1(\Inst_LH_LUT4c_frame_config_dffesr.c_reset_value ),
    .A2(_0986_));
 sg13g2_o21ai_1 _2392_ (.B1(_0975_),
    .VDD(VPWR),
    .Y(_0000_),
    .VSS(VGND),
    .A1(_0987_),
    .A2(_0988_));
 sg13g2_nand2_1 _2393_ (.Y(_0989_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit10.Q ),
    .B(_0985_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _2394_ (.Y(_0990_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit11.Q ),
    .A_N(_0973_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _2395_ (.A0(\Inst_LA_LUT4c_frame_config_dffesr.c_reset_value ),
    .A1(_0069_),
    .S(_0989_),
    .X(_0991_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _2396_ (.A0(\Inst_LA_LUT4c_frame_config_dffesr.LUT_flop ),
    .A1(_0991_),
    .S(_0990_),
    .X(_0001_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _2397_ (.Y(_0992_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit21.Q ),
    .A_N(_0973_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2398_ (.Y(_0993_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit20.Q ),
    .B(_0985_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _2399_ (.A0(\Inst_LB_LUT4c_frame_config_dffesr.c_reset_value ),
    .A1(_0109_),
    .S(_0993_),
    .X(_0994_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _2400_ (.A0(\Inst_LB_LUT4c_frame_config_dffesr.LUT_flop ),
    .A1(_0994_),
    .S(_0992_),
    .X(_0002_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _2401_ (.Y(_0995_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit31.Q ),
    .A_N(_0973_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2402_ (.Y(_0996_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit30.Q ),
    .B(_0985_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _2403_ (.A0(\Inst_LC_LUT4c_frame_config_dffesr.c_reset_value ),
    .A1(_0467_),
    .S(_0996_),
    .X(_0997_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _2404_ (.A0(\Inst_LC_LUT4c_frame_config_dffesr.LUT_flop ),
    .A1(_0997_),
    .S(_0995_),
    .X(_0003_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _2405_ (.Y(_0998_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit9.Q ),
    .A_N(_0973_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2406_ (.Y(_0999_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit8.Q ),
    .B(_0985_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _2407_ (.A0(\Inst_LD_LUT4c_frame_config_dffesr.c_reset_value ),
    .A1(_0688_),
    .S(_0999_),
    .X(_1000_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _2408_ (.A0(\Inst_LD_LUT4c_frame_config_dffesr.LUT_flop ),
    .A1(_1000_),
    .S(_0998_),
    .X(_0004_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _2409_ (.Y(_1001_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit19.Q ),
    .A_N(_0973_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2410_ (.Y(_1002_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit18.Q ),
    .B(_0985_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _2411_ (.A0(\Inst_LE_LUT4c_frame_config_dffesr.c_reset_value ),
    .A1(_0348_),
    .S(_1002_),
    .X(_1003_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _2412_ (.A0(\Inst_LE_LUT4c_frame_config_dffesr.LUT_flop ),
    .A1(_1003_),
    .S(_1001_),
    .X(_0005_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _2413_ (.Y(_1004_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit29.Q ),
    .A_N(_0973_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2414_ (.Y(_1005_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit28.Q ),
    .B(_0985_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _2415_ (.A0(\Inst_LF_LUT4c_frame_config_dffesr.c_reset_value ),
    .A1(_0496_),
    .S(_1005_),
    .X(_1006_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _2416_ (.A0(\Inst_LF_LUT4c_frame_config_dffesr.LUT_flop ),
    .A1(_1006_),
    .S(_1004_),
    .X(_0006_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _2417_ (.Y(_1007_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit7.Q ),
    .A_N(_0973_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3b_1 _2418_ (.B(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit7.Q ),
    .C(\Inst_LG_LUT4c_frame_config_dffesr.LUT_flop ),
    .Y(_1008_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(_0973_));
 sg13g2_nand2_1 _2419_ (.Y(_1009_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit6.Q ),
    .B(_0985_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _2420_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit6.Q ),
    .C1(_0630_),
    .B1(_0985_),
    .A1(_0632_),
    .Y(_1010_),
    .A2(_0635_));
 sg13g2_o21ai_1 _2421_ (.B1(_1007_),
    .VDD(VPWR),
    .Y(_1011_),
    .VSS(VGND),
    .A1(\Inst_LG_LUT4c_frame_config_dffesr.c_reset_value ),
    .A2(_1009_));
 sg13g2_o21ai_1 _2422_ (.B1(_1008_),
    .VDD(VPWR),
    .Y(_0007_),
    .VSS(VGND),
    .A1(_1010_),
    .A2(_1011_));
 sg13g2_dlhq_1 _2423_ (.D(FrameData[24]),
    .GATE(FrameStrobe[19]),
    .Q(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2424_ (.D(FrameData[25]),
    .GATE(FrameStrobe[19]),
    .Q(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2425_ (.D(FrameData[26]),
    .GATE(FrameStrobe[19]),
    .Q(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2426_ (.D(FrameData[27]),
    .GATE(FrameStrobe[19]),
    .Q(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2427_ (.D(FrameData[28]),
    .GATE(FrameStrobe[19]),
    .Q(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2428_ (.D(FrameData[29]),
    .GATE(FrameStrobe[19]),
    .Q(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2429_ (.D(FrameData[30]),
    .GATE(FrameStrobe[19]),
    .Q(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2430_ (.D(FrameData[31]),
    .GATE(FrameStrobe[19]),
    .Q(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2431_ (.D(FrameData[0]),
    .GATE(FrameStrobe[18]),
    .Q(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2432_ (.D(FrameData[1]),
    .GATE(FrameStrobe[18]),
    .Q(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2433_ (.D(FrameData[2]),
    .GATE(FrameStrobe[18]),
    .Q(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2434_ (.D(FrameData[3]),
    .GATE(FrameStrobe[18]),
    .Q(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2435_ (.D(FrameData[4]),
    .GATE(FrameStrobe[18]),
    .Q(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2436_ (.D(FrameData[5]),
    .GATE(FrameStrobe[18]),
    .Q(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2437_ (.D(FrameData[6]),
    .GATE(FrameStrobe[18]),
    .Q(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2438_ (.D(FrameData[7]),
    .GATE(FrameStrobe[18]),
    .Q(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2439_ (.D(FrameData[8]),
    .GATE(FrameStrobe[18]),
    .Q(\Inst_LA_LUT4c_frame_config_dffesr.c_out_mux ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2440_ (.D(FrameData[9]),
    .GATE(FrameStrobe[18]),
    .Q(\Inst_LA_LUT4c_frame_config_dffesr.c_I0mux ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2441_ (.D(FrameData[10]),
    .GATE(FrameStrobe[18]),
    .Q(\Inst_LA_LUT4c_frame_config_dffesr.c_reset_value ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2442_ (.D(FrameData[11]),
    .GATE(FrameStrobe[18]),
    .Q(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2443_ (.D(FrameData[12]),
    .GATE(FrameStrobe[18]),
    .Q(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2444_ (.D(FrameData[13]),
    .GATE(FrameStrobe[18]),
    .Q(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2445_ (.D(FrameData[14]),
    .GATE(FrameStrobe[18]),
    .Q(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2446_ (.D(FrameData[15]),
    .GATE(FrameStrobe[18]),
    .Q(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2447_ (.D(FrameData[16]),
    .GATE(FrameStrobe[18]),
    .Q(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2448_ (.D(FrameData[17]),
    .GATE(FrameStrobe[18]),
    .Q(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2449_ (.D(FrameData[18]),
    .GATE(FrameStrobe[18]),
    .Q(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2450_ (.D(FrameData[19]),
    .GATE(FrameStrobe[18]),
    .Q(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2451_ (.D(FrameData[20]),
    .GATE(FrameStrobe[18]),
    .Q(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2452_ (.D(FrameData[21]),
    .GATE(FrameStrobe[18]),
    .Q(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2453_ (.D(FrameData[22]),
    .GATE(FrameStrobe[18]),
    .Q(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2454_ (.D(FrameData[23]),
    .GATE(FrameStrobe[18]),
    .Q(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2455_ (.D(FrameData[24]),
    .GATE(FrameStrobe[18]),
    .Q(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2456_ (.D(FrameData[25]),
    .GATE(FrameStrobe[18]),
    .Q(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2457_ (.D(FrameData[26]),
    .GATE(FrameStrobe[18]),
    .Q(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2458_ (.D(FrameData[27]),
    .GATE(FrameStrobe[18]),
    .Q(\Inst_LB_LUT4c_frame_config_dffesr.c_out_mux ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2459_ (.D(FrameData[28]),
    .GATE(FrameStrobe[18]),
    .Q(\Inst_LB_LUT4c_frame_config_dffesr.c_I0mux ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2460_ (.D(FrameData[29]),
    .GATE(FrameStrobe[18]),
    .Q(\Inst_LB_LUT4c_frame_config_dffesr.c_reset_value ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2461_ (.D(FrameData[30]),
    .GATE(FrameStrobe[18]),
    .Q(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2462_ (.D(FrameData[31]),
    .GATE(FrameStrobe[18]),
    .Q(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2463_ (.D(FrameData[0]),
    .GATE(FrameStrobe[17]),
    .Q(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2464_ (.D(FrameData[1]),
    .GATE(FrameStrobe[17]),
    .Q(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2465_ (.D(FrameData[2]),
    .GATE(FrameStrobe[17]),
    .Q(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2466_ (.D(FrameData[3]),
    .GATE(FrameStrobe[17]),
    .Q(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2467_ (.D(FrameData[4]),
    .GATE(FrameStrobe[17]),
    .Q(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2468_ (.D(FrameData[5]),
    .GATE(FrameStrobe[17]),
    .Q(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2469_ (.D(FrameData[6]),
    .GATE(FrameStrobe[17]),
    .Q(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2470_ (.D(FrameData[7]),
    .GATE(FrameStrobe[17]),
    .Q(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2471_ (.D(FrameData[8]),
    .GATE(FrameStrobe[17]),
    .Q(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2472_ (.D(FrameData[9]),
    .GATE(FrameStrobe[17]),
    .Q(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2473_ (.D(FrameData[10]),
    .GATE(FrameStrobe[17]),
    .Q(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2474_ (.D(FrameData[11]),
    .GATE(FrameStrobe[17]),
    .Q(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2475_ (.D(FrameData[12]),
    .GATE(FrameStrobe[17]),
    .Q(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2476_ (.D(FrameData[13]),
    .GATE(FrameStrobe[17]),
    .Q(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2477_ (.D(FrameData[14]),
    .GATE(FrameStrobe[17]),
    .Q(\Inst_LC_LUT4c_frame_config_dffesr.c_out_mux ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2478_ (.D(FrameData[15]),
    .GATE(FrameStrobe[17]),
    .Q(\Inst_LC_LUT4c_frame_config_dffesr.c_I0mux ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2479_ (.D(FrameData[16]),
    .GATE(FrameStrobe[17]),
    .Q(\Inst_LC_LUT4c_frame_config_dffesr.c_reset_value ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2480_ (.D(FrameData[17]),
    .GATE(FrameStrobe[17]),
    .Q(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2481_ (.D(FrameData[18]),
    .GATE(FrameStrobe[17]),
    .Q(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2482_ (.D(FrameData[19]),
    .GATE(FrameStrobe[17]),
    .Q(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2483_ (.D(FrameData[20]),
    .GATE(FrameStrobe[17]),
    .Q(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2484_ (.D(FrameData[21]),
    .GATE(FrameStrobe[17]),
    .Q(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2485_ (.D(FrameData[22]),
    .GATE(FrameStrobe[17]),
    .Q(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2486_ (.D(FrameData[23]),
    .GATE(FrameStrobe[17]),
    .Q(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2487_ (.D(FrameData[24]),
    .GATE(FrameStrobe[17]),
    .Q(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2488_ (.D(FrameData[25]),
    .GATE(FrameStrobe[17]),
    .Q(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2489_ (.D(FrameData[26]),
    .GATE(FrameStrobe[17]),
    .Q(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2490_ (.D(FrameData[27]),
    .GATE(FrameStrobe[17]),
    .Q(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2491_ (.D(FrameData[28]),
    .GATE(FrameStrobe[17]),
    .Q(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2492_ (.D(FrameData[29]),
    .GATE(FrameStrobe[17]),
    .Q(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2493_ (.D(FrameData[30]),
    .GATE(FrameStrobe[17]),
    .Q(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2494_ (.D(FrameData[31]),
    .GATE(FrameStrobe[17]),
    .Q(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2495_ (.D(FrameData[0]),
    .GATE(FrameStrobe[16]),
    .Q(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2496_ (.D(FrameData[1]),
    .GATE(FrameStrobe[16]),
    .Q(\Inst_LD_LUT4c_frame_config_dffesr.c_out_mux ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2497_ (.D(FrameData[2]),
    .GATE(FrameStrobe[16]),
    .Q(\Inst_LD_LUT4c_frame_config_dffesr.c_I0mux ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2498_ (.D(FrameData[3]),
    .GATE(FrameStrobe[16]),
    .Q(\Inst_LD_LUT4c_frame_config_dffesr.c_reset_value ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2499_ (.D(FrameData[4]),
    .GATE(FrameStrobe[16]),
    .Q(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2500_ (.D(FrameData[5]),
    .GATE(FrameStrobe[16]),
    .Q(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2501_ (.D(FrameData[6]),
    .GATE(FrameStrobe[16]),
    .Q(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2502_ (.D(FrameData[7]),
    .GATE(FrameStrobe[16]),
    .Q(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2503_ (.D(FrameData[8]),
    .GATE(FrameStrobe[16]),
    .Q(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2504_ (.D(FrameData[9]),
    .GATE(FrameStrobe[16]),
    .Q(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2505_ (.D(FrameData[10]),
    .GATE(FrameStrobe[16]),
    .Q(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2506_ (.D(FrameData[11]),
    .GATE(FrameStrobe[16]),
    .Q(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2507_ (.D(FrameData[12]),
    .GATE(FrameStrobe[16]),
    .Q(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2508_ (.D(FrameData[13]),
    .GATE(FrameStrobe[16]),
    .Q(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2509_ (.D(FrameData[14]),
    .GATE(FrameStrobe[16]),
    .Q(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2510_ (.D(FrameData[15]),
    .GATE(FrameStrobe[16]),
    .Q(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2511_ (.D(FrameData[16]),
    .GATE(FrameStrobe[16]),
    .Q(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2512_ (.D(FrameData[17]),
    .GATE(FrameStrobe[16]),
    .Q(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2513_ (.D(FrameData[18]),
    .GATE(FrameStrobe[16]),
    .Q(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2514_ (.D(FrameData[19]),
    .GATE(FrameStrobe[16]),
    .Q(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2515_ (.D(FrameData[20]),
    .GATE(FrameStrobe[16]),
    .Q(\Inst_LE_LUT4c_frame_config_dffesr.c_out_mux ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2516_ (.D(FrameData[21]),
    .GATE(FrameStrobe[16]),
    .Q(\Inst_LE_LUT4c_frame_config_dffesr.c_I0mux ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2517_ (.D(FrameData[22]),
    .GATE(FrameStrobe[16]),
    .Q(\Inst_LE_LUT4c_frame_config_dffesr.c_reset_value ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2518_ (.D(FrameData[23]),
    .GATE(FrameStrobe[16]),
    .Q(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2519_ (.D(FrameData[24]),
    .GATE(FrameStrobe[16]),
    .Q(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2520_ (.D(FrameData[25]),
    .GATE(FrameStrobe[16]),
    .Q(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2521_ (.D(FrameData[26]),
    .GATE(FrameStrobe[16]),
    .Q(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2522_ (.D(FrameData[27]),
    .GATE(FrameStrobe[16]),
    .Q(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2523_ (.D(FrameData[28]),
    .GATE(FrameStrobe[16]),
    .Q(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2524_ (.D(FrameData[29]),
    .GATE(FrameStrobe[16]),
    .Q(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2525_ (.D(FrameData[30]),
    .GATE(FrameStrobe[16]),
    .Q(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2526_ (.D(FrameData[31]),
    .GATE(FrameStrobe[16]),
    .Q(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2527_ (.D(FrameData[0]),
    .GATE(FrameStrobe[15]),
    .Q(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2528_ (.D(FrameData[1]),
    .GATE(FrameStrobe[15]),
    .Q(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2529_ (.D(FrameData[2]),
    .GATE(FrameStrobe[15]),
    .Q(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2530_ (.D(FrameData[3]),
    .GATE(FrameStrobe[15]),
    .Q(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2531_ (.D(FrameData[4]),
    .GATE(FrameStrobe[15]),
    .Q(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2532_ (.D(FrameData[5]),
    .GATE(FrameStrobe[15]),
    .Q(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2533_ (.D(FrameData[6]),
    .GATE(FrameStrobe[15]),
    .Q(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2534_ (.D(FrameData[7]),
    .GATE(FrameStrobe[15]),
    .Q(\Inst_LF_LUT4c_frame_config_dffesr.c_out_mux ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2535_ (.D(FrameData[8]),
    .GATE(FrameStrobe[15]),
    .Q(\Inst_LF_LUT4c_frame_config_dffesr.c_I0mux ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2536_ (.D(FrameData[9]),
    .GATE(FrameStrobe[15]),
    .Q(\Inst_LF_LUT4c_frame_config_dffesr.c_reset_value ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2537_ (.D(FrameData[10]),
    .GATE(FrameStrobe[15]),
    .Q(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2538_ (.D(FrameData[11]),
    .GATE(FrameStrobe[15]),
    .Q(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2539_ (.D(FrameData[12]),
    .GATE(FrameStrobe[15]),
    .Q(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2540_ (.D(FrameData[13]),
    .GATE(FrameStrobe[15]),
    .Q(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2541_ (.D(FrameData[14]),
    .GATE(FrameStrobe[15]),
    .Q(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2542_ (.D(FrameData[15]),
    .GATE(FrameStrobe[15]),
    .Q(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2543_ (.D(FrameData[16]),
    .GATE(FrameStrobe[15]),
    .Q(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2544_ (.D(FrameData[17]),
    .GATE(FrameStrobe[15]),
    .Q(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2545_ (.D(FrameData[18]),
    .GATE(FrameStrobe[15]),
    .Q(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2546_ (.D(FrameData[19]),
    .GATE(FrameStrobe[15]),
    .Q(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2547_ (.D(FrameData[20]),
    .GATE(FrameStrobe[15]),
    .Q(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2548_ (.D(FrameData[21]),
    .GATE(FrameStrobe[15]),
    .Q(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2549_ (.D(FrameData[22]),
    .GATE(FrameStrobe[15]),
    .Q(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2550_ (.D(FrameData[23]),
    .GATE(FrameStrobe[15]),
    .Q(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2551_ (.D(FrameData[24]),
    .GATE(FrameStrobe[15]),
    .Q(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2552_ (.D(FrameData[25]),
    .GATE(FrameStrobe[15]),
    .Q(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2553_ (.D(FrameData[26]),
    .GATE(FrameStrobe[15]),
    .Q(\Inst_LG_LUT4c_frame_config_dffesr.c_out_mux ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2554_ (.D(FrameData[27]),
    .GATE(FrameStrobe[15]),
    .Q(\Inst_LG_LUT4c_frame_config_dffesr.c_I0mux ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2555_ (.D(FrameData[28]),
    .GATE(FrameStrobe[15]),
    .Q(\Inst_LG_LUT4c_frame_config_dffesr.c_reset_value ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2556_ (.D(FrameData[29]),
    .GATE(FrameStrobe[15]),
    .Q(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2557_ (.D(FrameData[30]),
    .GATE(FrameStrobe[15]),
    .Q(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2558_ (.D(FrameData[31]),
    .GATE(FrameStrobe[15]),
    .Q(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2559_ (.D(FrameData[0]),
    .GATE(FrameStrobe[14]),
    .Q(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2560_ (.D(FrameData[1]),
    .GATE(FrameStrobe[14]),
    .Q(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2561_ (.D(FrameData[2]),
    .GATE(FrameStrobe[14]),
    .Q(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2562_ (.D(FrameData[3]),
    .GATE(FrameStrobe[14]),
    .Q(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2563_ (.D(FrameData[4]),
    .GATE(FrameStrobe[14]),
    .Q(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2564_ (.D(FrameData[5]),
    .GATE(FrameStrobe[14]),
    .Q(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2565_ (.D(FrameData[6]),
    .GATE(FrameStrobe[14]),
    .Q(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2566_ (.D(FrameData[7]),
    .GATE(FrameStrobe[14]),
    .Q(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2567_ (.D(FrameData[8]),
    .GATE(FrameStrobe[14]),
    .Q(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2568_ (.D(FrameData[9]),
    .GATE(FrameStrobe[14]),
    .Q(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2569_ (.D(FrameData[10]),
    .GATE(FrameStrobe[14]),
    .Q(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2570_ (.D(FrameData[11]),
    .GATE(FrameStrobe[14]),
    .Q(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2571_ (.D(FrameData[12]),
    .GATE(FrameStrobe[14]),
    .Q(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2572_ (.D(FrameData[13]),
    .GATE(FrameStrobe[14]),
    .Q(\Inst_LH_LUT4c_frame_config_dffesr.c_out_mux ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2573_ (.D(FrameData[14]),
    .GATE(FrameStrobe[14]),
    .Q(\Inst_LH_LUT4c_frame_config_dffesr.c_I0mux ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2574_ (.D(FrameData[15]),
    .GATE(FrameStrobe[14]),
    .Q(\Inst_LH_LUT4c_frame_config_dffesr.c_reset_value ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2575_ (.D(FrameData[16]),
    .GATE(FrameStrobe[14]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit16.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2576_ (.D(FrameData[17]),
    .GATE(FrameStrobe[14]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit17.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2577_ (.D(FrameData[18]),
    .GATE(FrameStrobe[14]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit18.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2578_ (.D(FrameData[19]),
    .GATE(FrameStrobe[14]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit19.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2579_ (.D(FrameData[20]),
    .GATE(FrameStrobe[14]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit20.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2580_ (.D(FrameData[21]),
    .GATE(FrameStrobe[14]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit21.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2581_ (.D(FrameData[22]),
    .GATE(FrameStrobe[14]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit22.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2582_ (.D(FrameData[23]),
    .GATE(FrameStrobe[14]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit23.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2583_ (.D(FrameData[24]),
    .GATE(FrameStrobe[14]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit24.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2584_ (.D(FrameData[25]),
    .GATE(FrameStrobe[14]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit25.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2585_ (.D(FrameData[26]),
    .GATE(FrameStrobe[14]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit26.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2586_ (.D(FrameData[27]),
    .GATE(FrameStrobe[14]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit27.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2587_ (.D(FrameData[28]),
    .GATE(FrameStrobe[14]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit28.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2588_ (.D(FrameData[29]),
    .GATE(FrameStrobe[14]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit29.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2589_ (.D(FrameData[30]),
    .GATE(FrameStrobe[14]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit30.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2590_ (.D(FrameData[31]),
    .GATE(FrameStrobe[14]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit31.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2591_ (.D(FrameData[0]),
    .GATE(FrameStrobe[13]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit0.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2592_ (.D(FrameData[1]),
    .GATE(FrameStrobe[13]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit1.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2593_ (.D(FrameData[2]),
    .GATE(FrameStrobe[13]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit2.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2594_ (.D(FrameData[3]),
    .GATE(FrameStrobe[13]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit3.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2595_ (.D(FrameData[4]),
    .GATE(FrameStrobe[13]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit4.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2596_ (.D(FrameData[5]),
    .GATE(FrameStrobe[13]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit5.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2597_ (.D(FrameData[6]),
    .GATE(FrameStrobe[13]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit6.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2598_ (.D(FrameData[7]),
    .GATE(FrameStrobe[13]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit7.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2599_ (.D(FrameData[8]),
    .GATE(FrameStrobe[13]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit8.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2600_ (.D(FrameData[9]),
    .GATE(FrameStrobe[13]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit9.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2601_ (.D(FrameData[10]),
    .GATE(FrameStrobe[13]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit10.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2602_ (.D(FrameData[11]),
    .GATE(FrameStrobe[13]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit11.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2603_ (.D(FrameData[12]),
    .GATE(FrameStrobe[13]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit12.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2604_ (.D(FrameData[13]),
    .GATE(FrameStrobe[13]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit13.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2605_ (.D(FrameData[14]),
    .GATE(FrameStrobe[13]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit14.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2606_ (.D(FrameData[15]),
    .GATE(FrameStrobe[13]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit15.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2607_ (.D(FrameData[16]),
    .GATE(FrameStrobe[13]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit16.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2608_ (.D(FrameData[17]),
    .GATE(FrameStrobe[13]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit17.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2609_ (.D(FrameData[18]),
    .GATE(FrameStrobe[13]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit18.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2610_ (.D(FrameData[19]),
    .GATE(FrameStrobe[13]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit19.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2611_ (.D(FrameData[20]),
    .GATE(FrameStrobe[13]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit20.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2612_ (.D(FrameData[21]),
    .GATE(FrameStrobe[13]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit21.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2613_ (.D(FrameData[22]),
    .GATE(FrameStrobe[13]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit22.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2614_ (.D(FrameData[23]),
    .GATE(FrameStrobe[13]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit23.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2615_ (.D(FrameData[24]),
    .GATE(FrameStrobe[13]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit24.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2616_ (.D(FrameData[25]),
    .GATE(FrameStrobe[13]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit25.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2617_ (.D(FrameData[26]),
    .GATE(FrameStrobe[13]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit26.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2618_ (.D(FrameData[27]),
    .GATE(FrameStrobe[13]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit27.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2619_ (.D(FrameData[28]),
    .GATE(FrameStrobe[13]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit28.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2620_ (.D(FrameData[29]),
    .GATE(FrameStrobe[13]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit29.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2621_ (.D(FrameData[30]),
    .GATE(FrameStrobe[13]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit30.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2622_ (.D(FrameData[31]),
    .GATE(FrameStrobe[13]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit31.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2623_ (.D(FrameData[0]),
    .GATE(FrameStrobe[12]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit0.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2624_ (.D(FrameData[1]),
    .GATE(FrameStrobe[12]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit1.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2625_ (.D(FrameData[2]),
    .GATE(FrameStrobe[12]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit2.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2626_ (.D(FrameData[3]),
    .GATE(FrameStrobe[12]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit3.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2627_ (.D(FrameData[4]),
    .GATE(FrameStrobe[12]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit4.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2628_ (.D(FrameData[5]),
    .GATE(FrameStrobe[12]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit5.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2629_ (.D(FrameData[6]),
    .GATE(FrameStrobe[12]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit6.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2630_ (.D(FrameData[7]),
    .GATE(FrameStrobe[12]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit7.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2631_ (.D(FrameData[8]),
    .GATE(FrameStrobe[12]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit8.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2632_ (.D(FrameData[9]),
    .GATE(FrameStrobe[12]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit9.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2633_ (.D(FrameData[10]),
    .GATE(FrameStrobe[12]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit10.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2634_ (.D(FrameData[11]),
    .GATE(FrameStrobe[12]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit11.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2635_ (.D(FrameData[12]),
    .GATE(FrameStrobe[12]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit12.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2636_ (.D(FrameData[13]),
    .GATE(FrameStrobe[12]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit13.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2637_ (.D(FrameData[14]),
    .GATE(FrameStrobe[12]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit14.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2638_ (.D(FrameData[15]),
    .GATE(FrameStrobe[12]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit15.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2639_ (.D(FrameData[16]),
    .GATE(FrameStrobe[12]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit16.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2640_ (.D(FrameData[17]),
    .GATE(FrameStrobe[12]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit17.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2641_ (.D(FrameData[18]),
    .GATE(FrameStrobe[12]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit18.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2642_ (.D(FrameData[19]),
    .GATE(FrameStrobe[12]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit19.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2643_ (.D(FrameData[20]),
    .GATE(FrameStrobe[12]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit20.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2644_ (.D(FrameData[21]),
    .GATE(FrameStrobe[12]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit21.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2645_ (.D(FrameData[22]),
    .GATE(FrameStrobe[12]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit22.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2646_ (.D(FrameData[23]),
    .GATE(FrameStrobe[12]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit23.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2647_ (.D(FrameData[24]),
    .GATE(FrameStrobe[12]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit24.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2648_ (.D(FrameData[25]),
    .GATE(FrameStrobe[12]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit25.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2649_ (.D(FrameData[26]),
    .GATE(FrameStrobe[12]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit26.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2650_ (.D(FrameData[27]),
    .GATE(FrameStrobe[12]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit27.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2651_ (.D(FrameData[28]),
    .GATE(FrameStrobe[12]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit28.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2652_ (.D(FrameData[29]),
    .GATE(FrameStrobe[12]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit29.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2653_ (.D(FrameData[30]),
    .GATE(FrameStrobe[12]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit30.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2654_ (.D(FrameData[31]),
    .GATE(FrameStrobe[12]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit31.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2655_ (.D(FrameData[0]),
    .GATE(FrameStrobe[11]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit0.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2656_ (.D(FrameData[1]),
    .GATE(FrameStrobe[11]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit1.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2657_ (.D(FrameData[2]),
    .GATE(FrameStrobe[11]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit2.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2658_ (.D(FrameData[3]),
    .GATE(FrameStrobe[11]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit3.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2659_ (.D(FrameData[4]),
    .GATE(FrameStrobe[11]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit4.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2660_ (.D(FrameData[5]),
    .GATE(FrameStrobe[11]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit5.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2661_ (.D(FrameData[6]),
    .GATE(FrameStrobe[11]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit6.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2662_ (.D(FrameData[7]),
    .GATE(FrameStrobe[11]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit7.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2663_ (.D(FrameData[8]),
    .GATE(FrameStrobe[11]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit8.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2664_ (.D(FrameData[9]),
    .GATE(FrameStrobe[11]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit9.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2665_ (.D(FrameData[10]),
    .GATE(FrameStrobe[11]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit10.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2666_ (.D(FrameData[11]),
    .GATE(FrameStrobe[11]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit11.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2667_ (.D(FrameData[12]),
    .GATE(FrameStrobe[11]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit12.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2668_ (.D(FrameData[13]),
    .GATE(FrameStrobe[11]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit13.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2669_ (.D(FrameData[14]),
    .GATE(FrameStrobe[11]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit14.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2670_ (.D(FrameData[15]),
    .GATE(FrameStrobe[11]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit15.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2671_ (.D(FrameData[16]),
    .GATE(FrameStrobe[11]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit16.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2672_ (.D(FrameData[17]),
    .GATE(FrameStrobe[11]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit17.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2673_ (.D(FrameData[18]),
    .GATE(FrameStrobe[11]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit18.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2674_ (.D(FrameData[19]),
    .GATE(FrameStrobe[11]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit19.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2675_ (.D(FrameData[20]),
    .GATE(FrameStrobe[11]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit20.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2676_ (.D(FrameData[21]),
    .GATE(FrameStrobe[11]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit21.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2677_ (.D(FrameData[22]),
    .GATE(FrameStrobe[11]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit22.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2678_ (.D(FrameData[23]),
    .GATE(FrameStrobe[11]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit23.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2679_ (.D(FrameData[24]),
    .GATE(FrameStrobe[11]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit24.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2680_ (.D(FrameData[25]),
    .GATE(FrameStrobe[11]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit25.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2681_ (.D(FrameData[26]),
    .GATE(FrameStrobe[11]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit26.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2682_ (.D(FrameData[27]),
    .GATE(FrameStrobe[11]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit27.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2683_ (.D(FrameData[28]),
    .GATE(FrameStrobe[11]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit28.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2684_ (.D(FrameData[29]),
    .GATE(FrameStrobe[11]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit29.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2685_ (.D(FrameData[30]),
    .GATE(FrameStrobe[11]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit30.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2686_ (.D(FrameData[31]),
    .GATE(FrameStrobe[11]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit31.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2687_ (.D(FrameData[0]),
    .GATE(FrameStrobe[10]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit0.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2688_ (.D(FrameData[1]),
    .GATE(FrameStrobe[10]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit1.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2689_ (.D(FrameData[2]),
    .GATE(FrameStrobe[10]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit2.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2690_ (.D(FrameData[3]),
    .GATE(FrameStrobe[10]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit3.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2691_ (.D(FrameData[4]),
    .GATE(FrameStrobe[10]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit4.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2692_ (.D(FrameData[5]),
    .GATE(FrameStrobe[10]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit5.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2693_ (.D(FrameData[6]),
    .GATE(FrameStrobe[10]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit6.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2694_ (.D(FrameData[7]),
    .GATE(FrameStrobe[10]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit7.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2695_ (.D(FrameData[8]),
    .GATE(FrameStrobe[10]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit8.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2696_ (.D(FrameData[9]),
    .GATE(FrameStrobe[10]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit9.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2697_ (.D(FrameData[10]),
    .GATE(FrameStrobe[10]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit10.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2698_ (.D(FrameData[11]),
    .GATE(FrameStrobe[10]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit11.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2699_ (.D(FrameData[12]),
    .GATE(FrameStrobe[10]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit12.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2700_ (.D(FrameData[13]),
    .GATE(FrameStrobe[10]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit13.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2701_ (.D(FrameData[14]),
    .GATE(FrameStrobe[10]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit14.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2702_ (.D(FrameData[15]),
    .GATE(FrameStrobe[10]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit15.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2703_ (.D(FrameData[16]),
    .GATE(FrameStrobe[10]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit16.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2704_ (.D(FrameData[17]),
    .GATE(FrameStrobe[10]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit17.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2705_ (.D(FrameData[18]),
    .GATE(FrameStrobe[10]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit18.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2706_ (.D(FrameData[19]),
    .GATE(FrameStrobe[10]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit19.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2707_ (.D(FrameData[20]),
    .GATE(FrameStrobe[10]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit20.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2708_ (.D(FrameData[21]),
    .GATE(FrameStrobe[10]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit21.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2709_ (.D(FrameData[22]),
    .GATE(FrameStrobe[10]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit22.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2710_ (.D(FrameData[23]),
    .GATE(FrameStrobe[10]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit23.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2711_ (.D(FrameData[24]),
    .GATE(FrameStrobe[10]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit24.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2712_ (.D(FrameData[25]),
    .GATE(FrameStrobe[10]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit25.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2713_ (.D(FrameData[26]),
    .GATE(FrameStrobe[10]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit26.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2714_ (.D(FrameData[27]),
    .GATE(FrameStrobe[10]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit27.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2715_ (.D(FrameData[28]),
    .GATE(FrameStrobe[10]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit28.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2716_ (.D(FrameData[29]),
    .GATE(FrameStrobe[10]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit29.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2717_ (.D(FrameData[30]),
    .GATE(FrameStrobe[10]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit30.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2718_ (.D(FrameData[31]),
    .GATE(FrameStrobe[10]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit31.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2719_ (.D(FrameData[0]),
    .GATE(FrameStrobe[9]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit0.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2720_ (.D(FrameData[1]),
    .GATE(FrameStrobe[9]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit1.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2721_ (.D(FrameData[2]),
    .GATE(FrameStrobe[9]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit2.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2722_ (.D(FrameData[3]),
    .GATE(FrameStrobe[9]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit3.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2723_ (.D(FrameData[4]),
    .GATE(FrameStrobe[9]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit4.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2724_ (.D(FrameData[5]),
    .GATE(FrameStrobe[9]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit5.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2725_ (.D(FrameData[6]),
    .GATE(FrameStrobe[9]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit6.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2726_ (.D(FrameData[7]),
    .GATE(FrameStrobe[9]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit7.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2727_ (.D(FrameData[8]),
    .GATE(FrameStrobe[9]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit8.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2728_ (.D(FrameData[9]),
    .GATE(FrameStrobe[9]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit9.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2729_ (.D(FrameData[10]),
    .GATE(FrameStrobe[9]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit10.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2730_ (.D(FrameData[11]),
    .GATE(FrameStrobe[9]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit11.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2731_ (.D(FrameData[12]),
    .GATE(FrameStrobe[9]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit12.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2732_ (.D(FrameData[13]),
    .GATE(FrameStrobe[9]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit13.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2733_ (.D(FrameData[14]),
    .GATE(FrameStrobe[9]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit14.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2734_ (.D(FrameData[15]),
    .GATE(FrameStrobe[9]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit15.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2735_ (.D(FrameData[16]),
    .GATE(FrameStrobe[9]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit16.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2736_ (.D(FrameData[17]),
    .GATE(FrameStrobe[9]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit17.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2737_ (.D(FrameData[18]),
    .GATE(FrameStrobe[9]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit18.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2738_ (.D(FrameData[19]),
    .GATE(FrameStrobe[9]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit19.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2739_ (.D(FrameData[20]),
    .GATE(FrameStrobe[9]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit20.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2740_ (.D(FrameData[21]),
    .GATE(FrameStrobe[9]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit21.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2741_ (.D(FrameData[22]),
    .GATE(FrameStrobe[9]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit22.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2742_ (.D(FrameData[23]),
    .GATE(FrameStrobe[9]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit23.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2743_ (.D(FrameData[24]),
    .GATE(FrameStrobe[9]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit24.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2744_ (.D(FrameData[25]),
    .GATE(FrameStrobe[9]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit25.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2745_ (.D(FrameData[26]),
    .GATE(FrameStrobe[9]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit26.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2746_ (.D(FrameData[27]),
    .GATE(FrameStrobe[9]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit27.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2747_ (.D(FrameData[28]),
    .GATE(FrameStrobe[9]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit28.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2748_ (.D(FrameData[29]),
    .GATE(FrameStrobe[9]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit29.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2749_ (.D(FrameData[30]),
    .GATE(FrameStrobe[9]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit30.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2750_ (.D(FrameData[31]),
    .GATE(FrameStrobe[9]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit31.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2751_ (.D(FrameData[0]),
    .GATE(FrameStrobe[8]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit0.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2752_ (.D(FrameData[1]),
    .GATE(FrameStrobe[8]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit1.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2753_ (.D(FrameData[2]),
    .GATE(FrameStrobe[8]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit2.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2754_ (.D(FrameData[3]),
    .GATE(FrameStrobe[8]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit3.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2755_ (.D(FrameData[4]),
    .GATE(FrameStrobe[8]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit4.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2756_ (.D(FrameData[5]),
    .GATE(FrameStrobe[8]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit5.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2757_ (.D(FrameData[6]),
    .GATE(FrameStrobe[8]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit6.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2758_ (.D(FrameData[7]),
    .GATE(FrameStrobe[8]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit7.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2759_ (.D(FrameData[8]),
    .GATE(FrameStrobe[8]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit8.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2760_ (.D(FrameData[9]),
    .GATE(FrameStrobe[8]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit9.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2761_ (.D(FrameData[10]),
    .GATE(FrameStrobe[8]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit10.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2762_ (.D(FrameData[11]),
    .GATE(FrameStrobe[8]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit11.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2763_ (.D(FrameData[12]),
    .GATE(FrameStrobe[8]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit12.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2764_ (.D(FrameData[13]),
    .GATE(FrameStrobe[8]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit13.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2765_ (.D(FrameData[14]),
    .GATE(FrameStrobe[8]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit14.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2766_ (.D(FrameData[15]),
    .GATE(FrameStrobe[8]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit15.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2767_ (.D(FrameData[16]),
    .GATE(FrameStrobe[8]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit16.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2768_ (.D(FrameData[17]),
    .GATE(FrameStrobe[8]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit17.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2769_ (.D(FrameData[18]),
    .GATE(FrameStrobe[8]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit18.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2770_ (.D(FrameData[19]),
    .GATE(FrameStrobe[8]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit19.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2771_ (.D(FrameData[20]),
    .GATE(FrameStrobe[8]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit20.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2772_ (.D(FrameData[21]),
    .GATE(FrameStrobe[8]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit21.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2773_ (.D(FrameData[22]),
    .GATE(FrameStrobe[8]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit22.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2774_ (.D(FrameData[23]),
    .GATE(FrameStrobe[8]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit23.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2775_ (.D(FrameData[24]),
    .GATE(FrameStrobe[8]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit24.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2776_ (.D(FrameData[25]),
    .GATE(FrameStrobe[8]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit25.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2777_ (.D(FrameData[26]),
    .GATE(FrameStrobe[8]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit26.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2778_ (.D(FrameData[27]),
    .GATE(FrameStrobe[8]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit27.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2779_ (.D(FrameData[28]),
    .GATE(FrameStrobe[8]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit28.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2780_ (.D(FrameData[29]),
    .GATE(FrameStrobe[8]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit29.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2781_ (.D(FrameData[30]),
    .GATE(FrameStrobe[8]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit30.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2782_ (.D(FrameData[31]),
    .GATE(FrameStrobe[8]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit31.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2783_ (.D(FrameData[0]),
    .GATE(FrameStrobe[7]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit0.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2784_ (.D(FrameData[1]),
    .GATE(FrameStrobe[7]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit1.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2785_ (.D(FrameData[2]),
    .GATE(FrameStrobe[7]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit2.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2786_ (.D(FrameData[3]),
    .GATE(FrameStrobe[7]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit3.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2787_ (.D(FrameData[4]),
    .GATE(FrameStrobe[7]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit4.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2788_ (.D(FrameData[5]),
    .GATE(FrameStrobe[7]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit5.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2789_ (.D(FrameData[6]),
    .GATE(FrameStrobe[7]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit6.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2790_ (.D(FrameData[7]),
    .GATE(FrameStrobe[7]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit7.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2791_ (.D(FrameData[8]),
    .GATE(FrameStrobe[7]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit8.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2792_ (.D(FrameData[9]),
    .GATE(FrameStrobe[7]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit9.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2793_ (.D(FrameData[10]),
    .GATE(FrameStrobe[7]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit10.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2794_ (.D(FrameData[11]),
    .GATE(FrameStrobe[7]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit11.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2795_ (.D(FrameData[12]),
    .GATE(FrameStrobe[7]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit12.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2796_ (.D(FrameData[13]),
    .GATE(FrameStrobe[7]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit13.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2797_ (.D(FrameData[14]),
    .GATE(FrameStrobe[7]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit14.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2798_ (.D(FrameData[15]),
    .GATE(FrameStrobe[7]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit15.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2799_ (.D(FrameData[16]),
    .GATE(FrameStrobe[7]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit16.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2800_ (.D(FrameData[17]),
    .GATE(FrameStrobe[7]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit17.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2801_ (.D(FrameData[18]),
    .GATE(FrameStrobe[7]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit18.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2802_ (.D(FrameData[19]),
    .GATE(FrameStrobe[7]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit19.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2803_ (.D(FrameData[20]),
    .GATE(FrameStrobe[7]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit20.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2804_ (.D(FrameData[21]),
    .GATE(FrameStrobe[7]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit21.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2805_ (.D(FrameData[22]),
    .GATE(FrameStrobe[7]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit22.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2806_ (.D(FrameData[23]),
    .GATE(FrameStrobe[7]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit23.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2807_ (.D(FrameData[24]),
    .GATE(FrameStrobe[7]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit24.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2808_ (.D(FrameData[25]),
    .GATE(FrameStrobe[7]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit25.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2809_ (.D(FrameData[26]),
    .GATE(FrameStrobe[7]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit26.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2810_ (.D(FrameData[27]),
    .GATE(FrameStrobe[7]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit27.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2811_ (.D(FrameData[28]),
    .GATE(FrameStrobe[7]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit28.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2812_ (.D(FrameData[29]),
    .GATE(FrameStrobe[7]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit29.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2813_ (.D(FrameData[30]),
    .GATE(FrameStrobe[7]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit30.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2814_ (.D(FrameData[31]),
    .GATE(FrameStrobe[7]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit31.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2815_ (.D(FrameData[0]),
    .GATE(FrameStrobe[6]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit0.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2816_ (.D(FrameData[1]),
    .GATE(FrameStrobe[6]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit1.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2817_ (.D(FrameData[2]),
    .GATE(FrameStrobe[6]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit2.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2818_ (.D(FrameData[3]),
    .GATE(FrameStrobe[6]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit3.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2819_ (.D(FrameData[4]),
    .GATE(FrameStrobe[6]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit4.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2820_ (.D(FrameData[5]),
    .GATE(FrameStrobe[6]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit5.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2821_ (.D(FrameData[6]),
    .GATE(FrameStrobe[6]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit6.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2822_ (.D(FrameData[7]),
    .GATE(FrameStrobe[6]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit7.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2823_ (.D(FrameData[8]),
    .GATE(FrameStrobe[6]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit8.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2824_ (.D(FrameData[9]),
    .GATE(FrameStrobe[6]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit9.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2825_ (.D(FrameData[10]),
    .GATE(FrameStrobe[6]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit10.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2826_ (.D(FrameData[11]),
    .GATE(FrameStrobe[6]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit11.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2827_ (.D(FrameData[12]),
    .GATE(FrameStrobe[6]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit12.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2828_ (.D(FrameData[13]),
    .GATE(FrameStrobe[6]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit13.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2829_ (.D(FrameData[14]),
    .GATE(FrameStrobe[6]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit14.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2830_ (.D(FrameData[15]),
    .GATE(FrameStrobe[6]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit15.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2831_ (.D(FrameData[16]),
    .GATE(FrameStrobe[6]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit16.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2832_ (.D(FrameData[17]),
    .GATE(FrameStrobe[6]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit17.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2833_ (.D(FrameData[18]),
    .GATE(FrameStrobe[6]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit18.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2834_ (.D(FrameData[19]),
    .GATE(FrameStrobe[6]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit19.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2835_ (.D(FrameData[20]),
    .GATE(FrameStrobe[6]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit20.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2836_ (.D(FrameData[21]),
    .GATE(FrameStrobe[6]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit21.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2837_ (.D(FrameData[22]),
    .GATE(FrameStrobe[6]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit22.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2838_ (.D(FrameData[23]),
    .GATE(FrameStrobe[6]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit23.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2839_ (.D(FrameData[24]),
    .GATE(FrameStrobe[6]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit24.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2840_ (.D(FrameData[25]),
    .GATE(FrameStrobe[6]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit25.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2841_ (.D(FrameData[26]),
    .GATE(FrameStrobe[6]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit26.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2842_ (.D(FrameData[27]),
    .GATE(FrameStrobe[6]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit27.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2843_ (.D(FrameData[28]),
    .GATE(FrameStrobe[6]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit28.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2844_ (.D(FrameData[29]),
    .GATE(FrameStrobe[6]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit29.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2845_ (.D(FrameData[30]),
    .GATE(FrameStrobe[6]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit30.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2846_ (.D(FrameData[31]),
    .GATE(FrameStrobe[6]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit31.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2847_ (.D(FrameData[0]),
    .GATE(FrameStrobe[5]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit0.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2848_ (.D(FrameData[1]),
    .GATE(FrameStrobe[5]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit1.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2849_ (.D(FrameData[2]),
    .GATE(FrameStrobe[5]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit2.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2850_ (.D(FrameData[3]),
    .GATE(FrameStrobe[5]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit3.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2851_ (.D(FrameData[4]),
    .GATE(FrameStrobe[5]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit4.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2852_ (.D(FrameData[5]),
    .GATE(FrameStrobe[5]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit5.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2853_ (.D(FrameData[6]),
    .GATE(FrameStrobe[5]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit6.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2854_ (.D(FrameData[7]),
    .GATE(FrameStrobe[5]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit7.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2855_ (.D(FrameData[8]),
    .GATE(FrameStrobe[5]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit8.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2856_ (.D(FrameData[9]),
    .GATE(FrameStrobe[5]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit9.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2857_ (.D(FrameData[10]),
    .GATE(FrameStrobe[5]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit10.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2858_ (.D(FrameData[11]),
    .GATE(FrameStrobe[5]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit11.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2859_ (.D(FrameData[12]),
    .GATE(FrameStrobe[5]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit12.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2860_ (.D(FrameData[13]),
    .GATE(FrameStrobe[5]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit13.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2861_ (.D(FrameData[14]),
    .GATE(FrameStrobe[5]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit14.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2862_ (.D(FrameData[15]),
    .GATE(FrameStrobe[5]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit15.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2863_ (.D(FrameData[16]),
    .GATE(FrameStrobe[5]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit16.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2864_ (.D(FrameData[17]),
    .GATE(FrameStrobe[5]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit17.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2865_ (.D(FrameData[18]),
    .GATE(FrameStrobe[5]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit18.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2866_ (.D(FrameData[19]),
    .GATE(FrameStrobe[5]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit19.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2867_ (.D(FrameData[20]),
    .GATE(FrameStrobe[5]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit20.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2868_ (.D(FrameData[21]),
    .GATE(FrameStrobe[5]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit21.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2869_ (.D(FrameData[22]),
    .GATE(FrameStrobe[5]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit22.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2870_ (.D(FrameData[23]),
    .GATE(FrameStrobe[5]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit23.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2871_ (.D(FrameData[24]),
    .GATE(FrameStrobe[5]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit24.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2872_ (.D(FrameData[25]),
    .GATE(FrameStrobe[5]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit25.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2873_ (.D(FrameData[26]),
    .GATE(FrameStrobe[5]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit26.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2874_ (.D(FrameData[27]),
    .GATE(FrameStrobe[5]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit27.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2875_ (.D(FrameData[28]),
    .GATE(FrameStrobe[5]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit28.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2876_ (.D(FrameData[29]),
    .GATE(FrameStrobe[5]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit29.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2877_ (.D(FrameData[30]),
    .GATE(FrameStrobe[5]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit30.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2878_ (.D(FrameData[31]),
    .GATE(FrameStrobe[5]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit31.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2879_ (.D(FrameData[0]),
    .GATE(FrameStrobe[4]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit0.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2880_ (.D(FrameData[1]),
    .GATE(FrameStrobe[4]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit1.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2881_ (.D(FrameData[2]),
    .GATE(FrameStrobe[4]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit2.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2882_ (.D(FrameData[3]),
    .GATE(FrameStrobe[4]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit3.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2883_ (.D(FrameData[4]),
    .GATE(FrameStrobe[4]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit4.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2884_ (.D(FrameData[5]),
    .GATE(FrameStrobe[4]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit5.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2885_ (.D(FrameData[6]),
    .GATE(FrameStrobe[4]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit6.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2886_ (.D(FrameData[7]),
    .GATE(FrameStrobe[4]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit7.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2887_ (.D(FrameData[8]),
    .GATE(FrameStrobe[4]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit8.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2888_ (.D(FrameData[9]),
    .GATE(FrameStrobe[4]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit9.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2889_ (.D(FrameData[10]),
    .GATE(FrameStrobe[4]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit10.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2890_ (.D(FrameData[11]),
    .GATE(FrameStrobe[4]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit11.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2891_ (.D(FrameData[12]),
    .GATE(FrameStrobe[4]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit12.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2892_ (.D(FrameData[13]),
    .GATE(FrameStrobe[4]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit13.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2893_ (.D(FrameData[14]),
    .GATE(FrameStrobe[4]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit14.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2894_ (.D(FrameData[15]),
    .GATE(FrameStrobe[4]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit15.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2895_ (.D(FrameData[16]),
    .GATE(FrameStrobe[4]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit16.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2896_ (.D(FrameData[17]),
    .GATE(FrameStrobe[4]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit17.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2897_ (.D(FrameData[18]),
    .GATE(FrameStrobe[4]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit18.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2898_ (.D(FrameData[19]),
    .GATE(FrameStrobe[4]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit19.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2899_ (.D(FrameData[20]),
    .GATE(FrameStrobe[4]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit20.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2900_ (.D(FrameData[21]),
    .GATE(FrameStrobe[4]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit21.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2901_ (.D(FrameData[22]),
    .GATE(FrameStrobe[4]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit22.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2902_ (.D(FrameData[23]),
    .GATE(FrameStrobe[4]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit23.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2903_ (.D(FrameData[24]),
    .GATE(FrameStrobe[4]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit24.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2904_ (.D(FrameData[25]),
    .GATE(FrameStrobe[4]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit25.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2905_ (.D(FrameData[26]),
    .GATE(FrameStrobe[4]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit26.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2906_ (.D(FrameData[27]),
    .GATE(FrameStrobe[4]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit27.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2907_ (.D(FrameData[28]),
    .GATE(FrameStrobe[4]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit28.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2908_ (.D(FrameData[29]),
    .GATE(FrameStrobe[4]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit29.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2909_ (.D(FrameData[30]),
    .GATE(FrameStrobe[4]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit30.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2910_ (.D(FrameData[31]),
    .GATE(FrameStrobe[4]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit31.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2911_ (.D(FrameData[0]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit0.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2912_ (.D(FrameData[1]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit1.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2913_ (.D(FrameData[2]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit2.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2914_ (.D(FrameData[3]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit3.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2915_ (.D(FrameData[4]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit4.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2916_ (.D(FrameData[5]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit5.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2917_ (.D(FrameData[6]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit6.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2918_ (.D(FrameData[7]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit7.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2919_ (.D(FrameData[8]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit8.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2920_ (.D(FrameData[9]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit9.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2921_ (.D(FrameData[10]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit10.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2922_ (.D(FrameData[11]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit11.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2923_ (.D(FrameData[12]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit12.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2924_ (.D(FrameData[13]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit13.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2925_ (.D(FrameData[14]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit14.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2926_ (.D(FrameData[15]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit15.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2927_ (.D(FrameData[16]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit16.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2928_ (.D(FrameData[17]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit17.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2929_ (.D(FrameData[18]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit18.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2930_ (.D(FrameData[19]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit19.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2931_ (.D(FrameData[20]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit20.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2932_ (.D(FrameData[21]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit21.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2933_ (.D(FrameData[22]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit22.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2934_ (.D(FrameData[23]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit23.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2935_ (.D(FrameData[24]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit24.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2936_ (.D(FrameData[25]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit25.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2937_ (.D(FrameData[26]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit26.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2938_ (.D(FrameData[27]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit27.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2939_ (.D(FrameData[28]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit28.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2940_ (.D(FrameData[29]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit29.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2941_ (.D(FrameData[30]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit30.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2942_ (.D(FrameData[31]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit31.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2943_ (.D(FrameData[0]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit0.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2944_ (.D(FrameData[1]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit1.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2945_ (.D(FrameData[2]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit2.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2946_ (.D(FrameData[3]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit3.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2947_ (.D(FrameData[4]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit4.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2948_ (.D(FrameData[5]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit5.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2949_ (.D(FrameData[6]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit6.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2950_ (.D(FrameData[7]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit7.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2951_ (.D(FrameData[8]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit8.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2952_ (.D(FrameData[9]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit9.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2953_ (.D(FrameData[10]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit10.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2954_ (.D(FrameData[11]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit11.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2955_ (.D(FrameData[12]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit12.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2956_ (.D(FrameData[13]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit13.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2957_ (.D(FrameData[14]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit14.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2958_ (.D(FrameData[15]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit15.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2959_ (.D(FrameData[16]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit16.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2960_ (.D(FrameData[17]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit17.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2961_ (.D(FrameData[18]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit18.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2962_ (.D(FrameData[19]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit19.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2963_ (.D(FrameData[20]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit20.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2964_ (.D(FrameData[21]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit21.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2965_ (.D(FrameData[22]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit22.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2966_ (.D(FrameData[23]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit23.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2967_ (.D(FrameData[24]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit24.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2968_ (.D(FrameData[25]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit25.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2969_ (.D(FrameData[26]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit26.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2970_ (.D(FrameData[27]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit27.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2971_ (.D(FrameData[28]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit28.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2972_ (.D(FrameData[29]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit29.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2973_ (.D(FrameData[30]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit30.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2974_ (.D(FrameData[31]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit31.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2975_ (.D(FrameData[0]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit0.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2976_ (.D(FrameData[1]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit1.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2977_ (.D(FrameData[2]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit2.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2978_ (.D(FrameData[3]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit3.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2979_ (.D(FrameData[4]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit4.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2980_ (.D(FrameData[5]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit5.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2981_ (.D(FrameData[6]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit6.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2982_ (.D(FrameData[7]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit7.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2983_ (.D(FrameData[8]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit8.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2984_ (.D(FrameData[9]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit9.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2985_ (.D(FrameData[10]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit10.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2986_ (.D(FrameData[11]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit11.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2987_ (.D(FrameData[12]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit12.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2988_ (.D(FrameData[13]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit13.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2989_ (.D(FrameData[14]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit14.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2990_ (.D(FrameData[15]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit15.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2991_ (.D(FrameData[16]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit16.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2992_ (.D(FrameData[17]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit17.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2993_ (.D(FrameData[18]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit18.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2994_ (.D(FrameData[19]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit19.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2995_ (.D(FrameData[20]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit20.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2996_ (.D(FrameData[21]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit21.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2997_ (.D(FrameData[22]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit22.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2998_ (.D(FrameData[23]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit23.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _2999_ (.D(FrameData[24]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit24.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _3000_ (.D(FrameData[25]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit25.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _3001_ (.D(FrameData[26]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit26.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _3002_ (.D(FrameData[27]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit27.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _3003_ (.D(FrameData[28]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit28.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _3004_ (.D(FrameData[29]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit29.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _3005_ (.D(FrameData[30]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit30.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _3006_ (.D(FrameData[31]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit31.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _3007_ (.D(FrameData[0]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit0.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _3008_ (.D(FrameData[1]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit1.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _3009_ (.D(FrameData[2]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit2.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _3010_ (.D(FrameData[3]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit3.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _3011_ (.D(FrameData[4]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit4.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _3012_ (.D(FrameData[5]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit5.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _3013_ (.D(FrameData[6]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit6.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _3014_ (.D(FrameData[7]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit7.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _3015_ (.D(FrameData[8]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit8.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _3016_ (.D(FrameData[9]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit9.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _3017_ (.D(FrameData[10]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit10.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _3018_ (.D(FrameData[11]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit11.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _3019_ (.D(FrameData[12]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit12.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _3020_ (.D(FrameData[13]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit13.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _3021_ (.D(FrameData[14]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit14.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _3022_ (.D(FrameData[15]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit15.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _3023_ (.D(FrameData[16]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit16.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _3024_ (.D(FrameData[17]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit17.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _3025_ (.D(FrameData[18]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit18.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _3026_ (.D(FrameData[19]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit19.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _3027_ (.D(FrameData[20]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit20.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _3028_ (.D(FrameData[21]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit21.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _3029_ (.D(FrameData[22]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit22.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _3030_ (.D(FrameData[23]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit23.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _3031_ (.D(FrameData[24]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit24.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _3032_ (.D(FrameData[25]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit25.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _3033_ (.D(FrameData[26]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit26.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _3034_ (.D(FrameData[27]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit27.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _3035_ (.D(FrameData[28]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit28.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _3036_ (.D(FrameData[29]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit29.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _3037_ (.D(FrameData[30]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit30.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _3038_ (.D(FrameData[31]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit31.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dfrbpq_1 _3039_ (.RESET_B(_1168_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0000_),
    .Q(\Inst_LH_LUT4c_frame_config_dffesr.LUT_flop ),
    .CLK(clknet_1_1__leaf_UserCLK_regs));
 sg13g2_dfrbpq_1 _3040_ (.RESET_B(_1167_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0001_),
    .Q(\Inst_LA_LUT4c_frame_config_dffesr.LUT_flop ),
    .CLK(clknet_1_0__leaf_UserCLK_regs));
 sg13g2_dfrbpq_1 _3041_ (.RESET_B(_1166_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0002_),
    .Q(\Inst_LB_LUT4c_frame_config_dffesr.LUT_flop ),
    .CLK(clknet_1_0__leaf_UserCLK_regs));
 sg13g2_dfrbpq_1 _3042_ (.RESET_B(_1165_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0003_),
    .Q(\Inst_LC_LUT4c_frame_config_dffesr.LUT_flop ),
    .CLK(clknet_1_0__leaf_UserCLK_regs));
 sg13g2_dfrbpq_1 _3043_ (.RESET_B(_1164_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0004_),
    .Q(\Inst_LD_LUT4c_frame_config_dffesr.LUT_flop ),
    .CLK(clknet_1_0__leaf_UserCLK_regs));
 sg13g2_dfrbpq_1 _3044_ (.RESET_B(_1163_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0005_),
    .Q(\Inst_LE_LUT4c_frame_config_dffesr.LUT_flop ),
    .CLK(clknet_1_1__leaf_UserCLK_regs));
 sg13g2_dfrbpq_1 _3045_ (.RESET_B(_1170_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0006_),
    .Q(\Inst_LF_LUT4c_frame_config_dffesr.LUT_flop ),
    .CLK(clknet_1_1__leaf_UserCLK_regs));
 sg13g2_dfrbpq_1 _3046_ (.RESET_B(_1169_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0007_),
    .Q(\Inst_LG_LUT4c_frame_config_dffesr.LUT_flop ),
    .CLK(clknet_1_1__leaf_UserCLK_regs));
 sg13g2_tiehi _3047_ (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(_1163_));
 sg13g2_tiehi _3048_ (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(_1164_));
 sg13g2_tiehi _3049_ (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(_1165_));
 sg13g2_tiehi _3050_ (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(_1166_));
 sg13g2_tiehi _3051_ (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(_1167_));
 sg13g2_tiehi _3052_ (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(_1168_));
 sg13g2_tiehi _3053_ (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(_1169_));
 sg13g2_tiehi _3054_ (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(_1170_));
 sg13g2_buf_1 _3055_ (.A(\Inst_LUT4AB_switch_matrix.E1BEG0 ),
    .X(E1BEG[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3056_ (.A(\Inst_LUT4AB_switch_matrix.E1BEG1 ),
    .X(E1BEG[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3057_ (.A(\Inst_LUT4AB_switch_matrix.E1BEG2 ),
    .X(E1BEG[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3058_ (.A(\Inst_LUT4AB_switch_matrix.E1BEG3 ),
    .X(E1BEG[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3059_ (.A(\Inst_LUT4AB_switch_matrix.E2BEG0 ),
    .X(E2BEG[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3060_ (.A(\Inst_LUT4AB_switch_matrix.E2BEG1 ),
    .X(E2BEG[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3061_ (.A(\Inst_LUT4AB_switch_matrix.E2BEG2 ),
    .X(E2BEG[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3062_ (.A(\Inst_LUT4AB_switch_matrix.E2BEG3 ),
    .X(E2BEG[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3063_ (.A(\Inst_LUT4AB_switch_matrix.E2BEG4 ),
    .X(E2BEG[4]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3064_ (.A(\Inst_LUT4AB_switch_matrix.E2BEG5 ),
    .X(E2BEG[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3065_ (.A(\Inst_LUT4AB_switch_matrix.E2BEG6 ),
    .X(E2BEG[6]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3066_ (.A(\Inst_LUT4AB_switch_matrix.E2BEG7 ),
    .X(E2BEG[7]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3067_ (.A(E2MID[0]),
    .X(E2BEGb[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3068_ (.A(E2MID[1]),
    .X(E2BEGb[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3069_ (.A(E2MID[2]),
    .X(E2BEGb[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3070_ (.A(E2MID[3]),
    .X(E2BEGb[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3071_ (.A(E2MID[4]),
    .X(E2BEGb[4]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3072_ (.A(E2MID[5]),
    .X(E2BEGb[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3073_ (.A(E2MID[6]),
    .X(E2BEGb[6]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3074_ (.A(E2MID[7]),
    .X(E2BEGb[7]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3075_ (.A(E6END[2]),
    .X(E6BEG[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3076_ (.A(E6END[3]),
    .X(E6BEG[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3077_ (.A(E6END[4]),
    .X(E6BEG[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3078_ (.A(E6END[5]),
    .X(E6BEG[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3079_ (.A(E6END[6]),
    .X(E6BEG[4]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3080_ (.A(E6END[7]),
    .X(E6BEG[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3081_ (.A(E6END[8]),
    .X(E6BEG[6]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3082_ (.A(E6END[9]),
    .X(E6BEG[7]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3083_ (.A(E6END[10]),
    .X(E6BEG[8]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3084_ (.A(E6END[11]),
    .X(E6BEG[9]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3085_ (.A(\Inst_LUT4AB_switch_matrix.E6BEG0 ),
    .X(E6BEG[10]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3086_ (.A(\Inst_LUT4AB_switch_matrix.E6BEG1 ),
    .X(E6BEG[11]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3087_ (.A(EE4END[4]),
    .X(EE4BEG[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3088_ (.A(EE4END[5]),
    .X(EE4BEG[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3089_ (.A(EE4END[6]),
    .X(EE4BEG[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3090_ (.A(EE4END[7]),
    .X(EE4BEG[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3091_ (.A(EE4END[8]),
    .X(EE4BEG[4]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3092_ (.A(EE4END[9]),
    .X(EE4BEG[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3093_ (.A(EE4END[10]),
    .X(EE4BEG[6]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3094_ (.A(EE4END[11]),
    .X(EE4BEG[7]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3095_ (.A(EE4END[12]),
    .X(EE4BEG[8]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3096_ (.A(EE4END[13]),
    .X(EE4BEG[9]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3097_ (.A(EE4END[14]),
    .X(EE4BEG[10]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3098_ (.A(EE4END[15]),
    .X(EE4BEG[11]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3099_ (.A(\Inst_LUT4AB_switch_matrix.EE4BEG0 ),
    .X(EE4BEG[12]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3100_ (.A(\Inst_LUT4AB_switch_matrix.EE4BEG1 ),
    .X(EE4BEG[13]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3101_ (.A(\Inst_LUT4AB_switch_matrix.EE4BEG2 ),
    .X(EE4BEG[14]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3102_ (.A(\Inst_LUT4AB_switch_matrix.EE4BEG3 ),
    .X(EE4BEG[15]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3103_ (.A(FrameData[0]),
    .X(FrameData_O[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3104_ (.A(FrameData[1]),
    .X(FrameData_O[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3105_ (.A(FrameData[2]),
    .X(FrameData_O[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3106_ (.A(FrameData[3]),
    .X(FrameData_O[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3107_ (.A(FrameData[4]),
    .X(FrameData_O[4]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3108_ (.A(FrameData[5]),
    .X(FrameData_O[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3109_ (.A(FrameData[6]),
    .X(FrameData_O[6]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3110_ (.A(FrameData[7]),
    .X(FrameData_O[7]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3111_ (.A(FrameData[8]),
    .X(FrameData_O[8]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3112_ (.A(FrameData[9]),
    .X(FrameData_O[9]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3113_ (.A(FrameData[10]),
    .X(FrameData_O[10]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3114_ (.A(FrameData[11]),
    .X(FrameData_O[11]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3115_ (.A(FrameData[12]),
    .X(FrameData_O[12]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3116_ (.A(FrameData[13]),
    .X(FrameData_O[13]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3117_ (.A(FrameData[14]),
    .X(FrameData_O[14]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3118_ (.A(FrameData[15]),
    .X(FrameData_O[15]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3119_ (.A(FrameData[16]),
    .X(FrameData_O[16]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3120_ (.A(FrameData[17]),
    .X(FrameData_O[17]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3121_ (.A(FrameData[18]),
    .X(FrameData_O[18]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3122_ (.A(FrameData[19]),
    .X(FrameData_O[19]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3123_ (.A(FrameData[20]),
    .X(FrameData_O[20]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3124_ (.A(FrameData[21]),
    .X(FrameData_O[21]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3125_ (.A(FrameData[22]),
    .X(FrameData_O[22]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3126_ (.A(FrameData[23]),
    .X(FrameData_O[23]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3127_ (.A(FrameData[24]),
    .X(FrameData_O[24]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3128_ (.A(FrameData[25]),
    .X(FrameData_O[25]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3129_ (.A(FrameData[26]),
    .X(FrameData_O[26]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3130_ (.A(FrameData[27]),
    .X(FrameData_O[27]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3131_ (.A(FrameData[28]),
    .X(FrameData_O[28]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3132_ (.A(FrameData[29]),
    .X(FrameData_O[29]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3133_ (.A(FrameData[30]),
    .X(FrameData_O[30]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3134_ (.A(FrameData[31]),
    .X(FrameData_O[31]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3135_ (.A(FrameStrobe[0]),
    .X(FrameStrobe_O[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3136_ (.A(FrameStrobe[1]),
    .X(FrameStrobe_O[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3137_ (.A(FrameStrobe[2]),
    .X(FrameStrobe_O[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3138_ (.A(FrameStrobe[3]),
    .X(FrameStrobe_O[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3139_ (.A(FrameStrobe[4]),
    .X(FrameStrobe_O[4]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3140_ (.A(FrameStrobe[5]),
    .X(FrameStrobe_O[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3141_ (.A(FrameStrobe[6]),
    .X(FrameStrobe_O[6]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3142_ (.A(FrameStrobe[7]),
    .X(FrameStrobe_O[7]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3143_ (.A(FrameStrobe[8]),
    .X(FrameStrobe_O[8]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3144_ (.A(FrameStrobe[9]),
    .X(FrameStrobe_O[9]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3145_ (.A(FrameStrobe[10]),
    .X(FrameStrobe_O[10]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3146_ (.A(FrameStrobe[11]),
    .X(FrameStrobe_O[11]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3147_ (.A(FrameStrobe[12]),
    .X(FrameStrobe_O[12]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3148_ (.A(FrameStrobe[13]),
    .X(FrameStrobe_O[13]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3149_ (.A(FrameStrobe[14]),
    .X(FrameStrobe_O[14]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3150_ (.A(FrameStrobe[15]),
    .X(FrameStrobe_O[15]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3151_ (.A(FrameStrobe[16]),
    .X(FrameStrobe_O[16]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3152_ (.A(FrameStrobe[17]),
    .X(FrameStrobe_O[17]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3153_ (.A(FrameStrobe[18]),
    .X(FrameStrobe_O[18]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3154_ (.A(FrameStrobe[19]),
    .X(FrameStrobe_O[19]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3155_ (.A(\Inst_LUT4AB_switch_matrix.N1BEG0 ),
    .X(N1BEG[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3156_ (.A(\Inst_LUT4AB_switch_matrix.N1BEG1 ),
    .X(N1BEG[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3157_ (.A(\Inst_LUT4AB_switch_matrix.N1BEG2 ),
    .X(N1BEG[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3158_ (.A(\Inst_LUT4AB_switch_matrix.N1BEG3 ),
    .X(N1BEG[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3159_ (.A(\Inst_LUT4AB_switch_matrix.JN2BEG0 ),
    .X(N2BEG[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3160_ (.A(\Inst_LUT4AB_switch_matrix.JN2BEG1 ),
    .X(N2BEG[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3161_ (.A(\Inst_LUT4AB_switch_matrix.JN2BEG2 ),
    .X(N2BEG[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3162_ (.A(\Inst_LUT4AB_switch_matrix.JN2BEG3 ),
    .X(N2BEG[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3163_ (.A(\Inst_LUT4AB_switch_matrix.JN2BEG4 ),
    .X(N2BEG[4]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3164_ (.A(\Inst_LUT4AB_switch_matrix.JN2BEG5 ),
    .X(N2BEG[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3165_ (.A(\Inst_LUT4AB_switch_matrix.JN2BEG6 ),
    .X(N2BEG[6]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3166_ (.A(\Inst_LUT4AB_switch_matrix.JN2BEG7 ),
    .X(N2BEG[7]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3167_ (.A(N2MID[0]),
    .X(N2BEGb[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3168_ (.A(N2MID[1]),
    .X(N2BEGb[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3169_ (.A(N2MID[2]),
    .X(N2BEGb[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3170_ (.A(N2MID[3]),
    .X(N2BEGb[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3171_ (.A(N2MID[4]),
    .X(N2BEGb[4]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3172_ (.A(N2MID[5]),
    .X(N2BEGb[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3173_ (.A(N2MID[6]),
    .X(N2BEGb[6]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3174_ (.A(N2MID[7]),
    .X(N2BEGb[7]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3175_ (.A(N4END[4]),
    .X(N4BEG[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3176_ (.A(N4END[5]),
    .X(N4BEG[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3177_ (.A(N4END[6]),
    .X(N4BEG[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3178_ (.A(N4END[7]),
    .X(N4BEG[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3179_ (.A(N4END[8]),
    .X(N4BEG[4]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3180_ (.A(N4END[9]),
    .X(N4BEG[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3181_ (.A(N4END[10]),
    .X(N4BEG[6]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3182_ (.A(N4END[11]),
    .X(N4BEG[7]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3183_ (.A(N4END[12]),
    .X(N4BEG[8]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3184_ (.A(N4END[13]),
    .X(N4BEG[9]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3185_ (.A(N4END[14]),
    .X(N4BEG[10]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3186_ (.A(N4END[15]),
    .X(N4BEG[11]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3187_ (.A(\Inst_LUT4AB_switch_matrix.N4BEG0 ),
    .X(N4BEG[12]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3188_ (.A(\Inst_LUT4AB_switch_matrix.N4BEG1 ),
    .X(N4BEG[13]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3189_ (.A(\Inst_LUT4AB_switch_matrix.N4BEG2 ),
    .X(N4BEG[14]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3190_ (.A(\Inst_LUT4AB_switch_matrix.N4BEG3 ),
    .X(N4BEG[15]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3191_ (.A(NN4END[4]),
    .X(NN4BEG[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3192_ (.A(NN4END[5]),
    .X(NN4BEG[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3193_ (.A(NN4END[6]),
    .X(NN4BEG[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3194_ (.A(NN4END[7]),
    .X(NN4BEG[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3195_ (.A(NN4END[8]),
    .X(NN4BEG[4]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3196_ (.A(NN4END[9]),
    .X(NN4BEG[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3197_ (.A(NN4END[10]),
    .X(NN4BEG[6]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3198_ (.A(NN4END[11]),
    .X(NN4BEG[7]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3199_ (.A(NN4END[12]),
    .X(NN4BEG[8]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3200_ (.A(NN4END[13]),
    .X(NN4BEG[9]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3201_ (.A(NN4END[14]),
    .X(NN4BEG[10]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3202_ (.A(NN4END[15]),
    .X(NN4BEG[11]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3203_ (.A(\Inst_LUT4AB_switch_matrix.NN4BEG0 ),
    .X(NN4BEG[12]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3204_ (.A(\Inst_LUT4AB_switch_matrix.NN4BEG1 ),
    .X(NN4BEG[13]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3205_ (.A(\Inst_LUT4AB_switch_matrix.NN4BEG2 ),
    .X(NN4BEG[14]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3206_ (.A(\Inst_LUT4AB_switch_matrix.NN4BEG3 ),
    .X(NN4BEG[15]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3207_ (.A(\Inst_LUT4AB_switch_matrix.S1BEG0 ),
    .X(S1BEG[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3208_ (.A(\Inst_LUT4AB_switch_matrix.S1BEG1 ),
    .X(S1BEG[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3209_ (.A(\Inst_LUT4AB_switch_matrix.S1BEG2 ),
    .X(S1BEG[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3210_ (.A(\Inst_LUT4AB_switch_matrix.S1BEG3 ),
    .X(S1BEG[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3211_ (.A(\Inst_LUT4AB_switch_matrix.JS2BEG0 ),
    .X(S2BEG[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3212_ (.A(\Inst_LUT4AB_switch_matrix.JS2BEG1 ),
    .X(S2BEG[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3213_ (.A(\Inst_LUT4AB_switch_matrix.JS2BEG2 ),
    .X(S2BEG[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3214_ (.A(\Inst_LUT4AB_switch_matrix.JS2BEG3 ),
    .X(S2BEG[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3215_ (.A(\Inst_LUT4AB_switch_matrix.JS2BEG4 ),
    .X(S2BEG[4]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3216_ (.A(\Inst_LUT4AB_switch_matrix.JS2BEG5 ),
    .X(S2BEG[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3217_ (.A(\Inst_LUT4AB_switch_matrix.JS2BEG6 ),
    .X(S2BEG[6]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3218_ (.A(\Inst_LUT4AB_switch_matrix.JS2BEG7 ),
    .X(S2BEG[7]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3219_ (.A(S2MID[0]),
    .X(S2BEGb[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3220_ (.A(S2MID[1]),
    .X(S2BEGb[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3221_ (.A(S2MID[2]),
    .X(S2BEGb[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3222_ (.A(S2MID[3]),
    .X(S2BEGb[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3223_ (.A(S2MID[4]),
    .X(S2BEGb[4]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3224_ (.A(S2MID[5]),
    .X(S2BEGb[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3225_ (.A(S2MID[6]),
    .X(S2BEGb[6]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3226_ (.A(S2MID[7]),
    .X(S2BEGb[7]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3227_ (.A(S4END[4]),
    .X(S4BEG[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3228_ (.A(S4END[5]),
    .X(S4BEG[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3229_ (.A(S4END[6]),
    .X(S4BEG[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3230_ (.A(S4END[7]),
    .X(S4BEG[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3231_ (.A(S4END[8]),
    .X(S4BEG[4]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3232_ (.A(S4END[9]),
    .X(S4BEG[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3233_ (.A(S4END[10]),
    .X(S4BEG[6]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3234_ (.A(S4END[11]),
    .X(S4BEG[7]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3235_ (.A(S4END[12]),
    .X(S4BEG[8]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3236_ (.A(S4END[13]),
    .X(S4BEG[9]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3237_ (.A(S4END[14]),
    .X(S4BEG[10]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3238_ (.A(S4END[15]),
    .X(S4BEG[11]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3239_ (.A(\Inst_LUT4AB_switch_matrix.S4BEG0 ),
    .X(S4BEG[12]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3240_ (.A(\Inst_LUT4AB_switch_matrix.S4BEG1 ),
    .X(S4BEG[13]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3241_ (.A(\Inst_LUT4AB_switch_matrix.S4BEG2 ),
    .X(S4BEG[14]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3242_ (.A(\Inst_LUT4AB_switch_matrix.S4BEG3 ),
    .X(S4BEG[15]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3243_ (.A(SS4END[4]),
    .X(SS4BEG[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3244_ (.A(SS4END[5]),
    .X(SS4BEG[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3245_ (.A(SS4END[6]),
    .X(SS4BEG[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3246_ (.A(SS4END[7]),
    .X(SS4BEG[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3247_ (.A(SS4END[8]),
    .X(SS4BEG[4]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3248_ (.A(SS4END[9]),
    .X(SS4BEG[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3249_ (.A(SS4END[10]),
    .X(SS4BEG[6]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3250_ (.A(SS4END[11]),
    .X(SS4BEG[7]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3251_ (.A(SS4END[12]),
    .X(SS4BEG[8]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3252_ (.A(SS4END[13]),
    .X(SS4BEG[9]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3253_ (.A(SS4END[14]),
    .X(SS4BEG[10]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3254_ (.A(SS4END[15]),
    .X(SS4BEG[11]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3255_ (.A(\Inst_LUT4AB_switch_matrix.SS4BEG0 ),
    .X(SS4BEG[12]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3256_ (.A(\Inst_LUT4AB_switch_matrix.SS4BEG1 ),
    .X(SS4BEG[13]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3257_ (.A(\Inst_LUT4AB_switch_matrix.SS4BEG2 ),
    .X(SS4BEG[14]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3258_ (.A(\Inst_LUT4AB_switch_matrix.SS4BEG3 ),
    .X(SS4BEG[15]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3259_ (.A(clknet_1_0__leaf_UserCLK),
    .X(UserCLKo),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3260_ (.A(\Inst_LUT4AB_switch_matrix.W1BEG0 ),
    .X(W1BEG[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3261_ (.A(\Inst_LUT4AB_switch_matrix.W1BEG1 ),
    .X(W1BEG[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3262_ (.A(\Inst_LUT4AB_switch_matrix.W1BEG2 ),
    .X(W1BEG[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3263_ (.A(\Inst_LUT4AB_switch_matrix.W1BEG3 ),
    .X(W1BEG[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3264_ (.A(\Inst_LUT4AB_switch_matrix.JW2BEG0 ),
    .X(W2BEG[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3265_ (.A(\Inst_LUT4AB_switch_matrix.JW2BEG1 ),
    .X(W2BEG[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3266_ (.A(\Inst_LUT4AB_switch_matrix.JW2BEG2 ),
    .X(W2BEG[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3267_ (.A(\Inst_LUT4AB_switch_matrix.JW2BEG3 ),
    .X(W2BEG[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3268_ (.A(\Inst_LUT4AB_switch_matrix.JW2BEG4 ),
    .X(W2BEG[4]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3269_ (.A(\Inst_LUT4AB_switch_matrix.JW2BEG5 ),
    .X(W2BEG[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3270_ (.A(\Inst_LUT4AB_switch_matrix.JW2BEG6 ),
    .X(W2BEG[6]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3271_ (.A(\Inst_LUT4AB_switch_matrix.JW2BEG7 ),
    .X(W2BEG[7]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3272_ (.A(W2MID[0]),
    .X(W2BEGb[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3273_ (.A(W2MID[1]),
    .X(W2BEGb[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3274_ (.A(W2MID[2]),
    .X(W2BEGb[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3275_ (.A(W2MID[3]),
    .X(W2BEGb[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3276_ (.A(W2MID[4]),
    .X(W2BEGb[4]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3277_ (.A(W2MID[5]),
    .X(W2BEGb[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3278_ (.A(W2MID[6]),
    .X(W2BEGb[6]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3279_ (.A(W2MID[7]),
    .X(W2BEGb[7]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3280_ (.A(W6END[2]),
    .X(W6BEG[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3281_ (.A(W6END[3]),
    .X(W6BEG[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3282_ (.A(W6END[4]),
    .X(W6BEG[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3283_ (.A(W6END[5]),
    .X(W6BEG[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3284_ (.A(W6END[6]),
    .X(W6BEG[4]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3285_ (.A(W6END[7]),
    .X(W6BEG[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3286_ (.A(W6END[8]),
    .X(W6BEG[6]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3287_ (.A(W6END[9]),
    .X(W6BEG[7]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3288_ (.A(W6END[10]),
    .X(W6BEG[8]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3289_ (.A(W6END[11]),
    .X(W6BEG[9]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3290_ (.A(\Inst_LUT4AB_switch_matrix.W6BEG0 ),
    .X(W6BEG[10]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3291_ (.A(\Inst_LUT4AB_switch_matrix.W6BEG1 ),
    .X(W6BEG[11]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3292_ (.A(WW4END[4]),
    .X(WW4BEG[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3293_ (.A(WW4END[5]),
    .X(WW4BEG[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3294_ (.A(WW4END[6]),
    .X(WW4BEG[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3295_ (.A(WW4END[7]),
    .X(WW4BEG[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3296_ (.A(WW4END[8]),
    .X(WW4BEG[4]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3297_ (.A(WW4END[9]),
    .X(WW4BEG[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3298_ (.A(WW4END[10]),
    .X(WW4BEG[6]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3299_ (.A(WW4END[11]),
    .X(WW4BEG[7]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3300_ (.A(WW4END[12]),
    .X(WW4BEG[8]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3301_ (.A(WW4END[13]),
    .X(WW4BEG[9]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3302_ (.A(WW4END[14]),
    .X(WW4BEG[10]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3303_ (.A(WW4END[15]),
    .X(WW4BEG[11]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3304_ (.A(\Inst_LUT4AB_switch_matrix.WW4BEG0 ),
    .X(WW4BEG[12]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3305_ (.A(\Inst_LUT4AB_switch_matrix.WW4BEG1 ),
    .X(WW4BEG[13]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3306_ (.A(\Inst_LUT4AB_switch_matrix.WW4BEG2 ),
    .X(WW4BEG[14]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3307_ (.A(\Inst_LUT4AB_switch_matrix.WW4BEG3 ),
    .X(WW4BEG[15]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_regs_0_UserCLK (.A(UserCLK),
    .X(UserCLK_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_0_UserCLK (.A(UserCLK),
    .X(clknet_0_UserCLK),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_1_0__f_UserCLK (.A(clknet_0_UserCLK),
    .X(clknet_1_0__leaf_UserCLK),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_0_UserCLK_regs (.A(UserCLK_regs),
    .X(clknet_0_UserCLK_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_1_0__f_UserCLK_regs (.A(clknet_0_UserCLK_regs),
    .X(clknet_1_0__leaf_UserCLK_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_1_1__f_UserCLK_regs (.A(clknet_0_UserCLK_regs),
    .X(clknet_1_1__leaf_UserCLK_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_antennanp ANTENNA_1 (.VDD(VPWR),
    .VSS(VGND),
    .A(EE4END[10]));
 sg13g2_antennanp ANTENNA_2 (.VDD(VPWR),
    .VSS(VGND),
    .A(EE4END[11]));
 sg13g2_antennanp ANTENNA_3 (.VDD(VPWR),
    .VSS(VGND),
    .A(EE4END[12]));
 sg13g2_antennanp ANTENNA_4 (.VDD(VPWR),
    .VSS(VGND),
    .A(EE4END[13]));
 sg13g2_antennanp ANTENNA_5 (.VDD(VPWR),
    .VSS(VGND),
    .A(EE4END[14]));
 sg13g2_antennanp ANTENNA_6 (.VDD(VPWR),
    .VSS(VGND),
    .A(EE4END[15]));
 sg13g2_antennanp ANTENNA_7 (.VDD(VPWR),
    .VSS(VGND),
    .A(EE4END[5]));
 sg13g2_antennanp ANTENNA_8 (.VDD(VPWR),
    .VSS(VGND),
    .A(EE4END[6]));
 sg13g2_antennanp ANTENNA_9 (.VDD(VPWR),
    .VSS(VGND),
    .A(EE4END[7]));
 sg13g2_antennanp ANTENNA_10 (.VDD(VPWR),
    .VSS(VGND),
    .A(N4END[12]));
 sg13g2_antennanp ANTENNA_11 (.VDD(VPWR),
    .VSS(VGND),
    .A(N4END[14]));
 sg13g2_antennanp ANTENNA_12 (.VDD(VPWR),
    .VSS(VGND),
    .A(N4END[5]));
 sg13g2_antennanp ANTENNA_13 (.VDD(VPWR),
    .VSS(VGND),
    .A(N4END[9]));
 sg13g2_antennanp ANTENNA_14 (.VDD(VPWR),
    .VSS(VGND),
    .A(NN4END[10]));
 sg13g2_antennanp ANTENNA_15 (.VDD(VPWR),
    .VSS(VGND),
    .A(NN4END[14]));
 sg13g2_antennanp ANTENNA_16 (.VDD(VPWR),
    .VSS(VGND),
    .A(NN4END[4]));
 sg13g2_antennanp ANTENNA_17 (.VDD(VPWR),
    .VSS(VGND),
    .A(NN4END[6]));
 sg13g2_antennanp ANTENNA_18 (.VDD(VPWR),
    .VSS(VGND),
    .A(NN4END[7]));
 sg13g2_antennanp ANTENNA_19 (.VDD(VPWR),
    .VSS(VGND),
    .A(S2END[1]));
 sg13g2_antennanp ANTENNA_20 (.VDD(VPWR),
    .VSS(VGND),
    .A(S2END[1]));
 sg13g2_antennanp ANTENNA_21 (.VDD(VPWR),
    .VSS(VGND),
    .A(S2END[1]));
 sg13g2_antennanp ANTENNA_22 (.VDD(VPWR),
    .VSS(VGND),
    .A(S2END[1]));
 sg13g2_antennanp ANTENNA_23 (.VDD(VPWR),
    .VSS(VGND),
    .A(S2END[1]));
 sg13g2_antennanp ANTENNA_24 (.VDD(VPWR),
    .VSS(VGND),
    .A(S2END[1]));
 sg13g2_antennanp ANTENNA_25 (.VDD(VPWR),
    .VSS(VGND),
    .A(S4END[0]));
 sg13g2_antennanp ANTENNA_26 (.VDD(VPWR),
    .VSS(VGND),
    .A(S4END[0]));
 sg13g2_antennanp ANTENNA_27 (.VDD(VPWR),
    .VSS(VGND),
    .A(S4END[0]));
 sg13g2_antennanp ANTENNA_28 (.VDD(VPWR),
    .VSS(VGND),
    .A(EE4END[8]));
 sg13g2_antennanp ANTENNA_29 (.VDD(VPWR),
    .VSS(VGND),
    .A(EE4END[9]));
 sg13g2_antennanp ANTENNA_30 (.VDD(VPWR),
    .VSS(VGND),
    .A(N2MID[6]));
 sg13g2_antennanp ANTENNA_31 (.VDD(VPWR),
    .VSS(VGND),
    .A(N2MID[6]));
 sg13g2_antennanp ANTENNA_32 (.VDD(VPWR),
    .VSS(VGND),
    .A(N2MID[6]));
 sg13g2_antennanp ANTENNA_33 (.VDD(VPWR),
    .VSS(VGND),
    .A(N2MID[6]));
 sg13g2_antennanp ANTENNA_34 (.VDD(VPWR),
    .VSS(VGND),
    .A(N4END[10]));
 sg13g2_antennanp ANTENNA_35 (.VDD(VPWR),
    .VSS(VGND),
    .A(N4END[11]));
 sg13g2_antennanp ANTENNA_36 (.VDD(VPWR),
    .VSS(VGND),
    .A(N4END[11]));
 sg13g2_antennanp ANTENNA_37 (.VDD(VPWR),
    .VSS(VGND),
    .A(N4END[15]));
 sg13g2_antennanp ANTENNA_38 (.VDD(VPWR),
    .VSS(VGND),
    .A(NN4END[11]));
 sg13g2_antennanp ANTENNA_39 (.VDD(VPWR),
    .VSS(VGND),
    .A(NN4END[13]));
 sg13g2_antennanp ANTENNA_40 (.VDD(VPWR),
    .VSS(VGND),
    .A(NN4END[15]));
 sg13g2_antennanp ANTENNA_41 (.VDD(VPWR),
    .VSS(VGND),
    .A(NN4END[15]));
 sg13g2_antennanp ANTENNA_42 (.VDD(VPWR),
    .VSS(VGND),
    .A(W2MID[6]));
 sg13g2_antennanp ANTENNA_43 (.VDD(VPWR),
    .VSS(VGND),
    .A(W2MID[6]));
 sg13g2_antennanp ANTENNA_44 (.VDD(VPWR),
    .VSS(VGND),
    .A(W2MID[6]));
 sg13g2_antennanp ANTENNA_45 (.VDD(VPWR),
    .VSS(VGND),
    .A(W2MID[6]));
 sg13g2_antennanp ANTENNA_46 (.VDD(VPWR),
    .VSS(VGND),
    .A(W2MID[6]));
 sg13g2_antennanp ANTENNA_47 (.VDD(VPWR),
    .VSS(VGND),
    .A(W2MID[6]));
 sg13g2_antennanp ANTENNA_48 (.VDD(VPWR),
    .VSS(VGND),
    .A(W2MID[6]));
 sg13g2_antennanp ANTENNA_49 (.VDD(VPWR),
    .VSS(VGND),
    .A(W2MID[6]));
 sg13g2_antennanp ANTENNA_50 (.VDD(VPWR),
    .VSS(VGND),
    .A(W2MID[6]));
 sg13g2_antennanp ANTENNA_51 (.VDD(VPWR),
    .VSS(VGND),
    .A(W2MID[6]));
 sg13g2_antennanp ANTENNA_52 (.VDD(VPWR),
    .VSS(VGND),
    .A(W2MID[6]));
 sg13g2_antennanp ANTENNA_53 (.VDD(VPWR),
    .VSS(VGND),
    .A(W2MID[6]));
 sg13g2_antennanp ANTENNA_54 (.VDD(VPWR),
    .VSS(VGND),
    .A(W2MID[6]));
 sg13g2_antennanp ANTENNA_55 (.VDD(VPWR),
    .VSS(VGND),
    .A(W2MID[6]));
 sg13g2_antennanp ANTENNA_56 (.VDD(VPWR),
    .VSS(VGND),
    .A(W2MID[6]));
 sg13g2_antennanp ANTENNA_57 (.VDD(VPWR),
    .VSS(VGND),
    .A(W2MID[6]));
 sg13g2_antennanp ANTENNA_58 (.VDD(VPWR),
    .VSS(VGND),
    .A(NN4END[5]));
 sg13g2_antennanp ANTENNA_59 (.VDD(VPWR),
    .VSS(VGND),
    .A(NN4END[8]));
 sg13g2_antennanp ANTENNA_60 (.VDD(VPWR),
    .VSS(VGND),
    .A(NN4END[9]));
 sg13g2_fill_1 FILLER_0_65 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_145 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_275 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_307 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_409 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_87 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_143 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_285 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_304 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_423 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_57 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_92 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_136 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_173 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_401 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_65 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_234 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_306 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_366 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_97 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_129 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_275 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_303 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_321 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_345 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_129 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_204 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_222 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_297 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_401 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_41 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_106 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_121 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_195 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_264 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_269 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_289 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_344 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_369 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_226 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_317 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_345 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_391 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_393 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_258 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_318 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_163 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_205 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_244 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_68 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_110 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_358 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_369 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_398 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_167 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_211 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_267 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_374 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_397 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_163 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_185 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_243 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_267 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_398 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_419 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_89 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_142 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_162 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_164 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_220 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_222 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_401 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_47 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_139 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_188 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_215 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_227 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_250 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_337 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_339 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_5 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_64 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_138 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_156 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_240 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_251 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_289 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_323 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_349 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_351 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_374 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_423 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_68 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_90 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_114 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_120 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_159 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_279 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_318 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_423 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_23 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_114 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_131 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_149 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_254 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_360 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_422 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_19 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_89 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_107 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_208 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_253 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_386 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_388 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_423 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_69 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_141 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_233 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_268 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_400 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_423 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_38 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_107 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_423 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_58 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_170 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_218 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_220 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_21_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_302 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_321 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_29 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_89 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_141 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_197 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_276 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_311 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_390 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_422 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_89 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_173 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_219 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_241 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_285 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_423 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_89 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_160 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_191 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_216 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_222 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_244 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_423 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_86 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_155 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_25_192 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_236 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_254 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_422 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_48 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_108 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_141 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_174 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_296 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_321 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_360 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_20 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_117 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_234 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_253 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_297 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_320 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_345 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_386 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_22 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_128 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_155 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_197 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_215 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_379 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_397 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_423 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_38 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_40 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_131 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_313 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_321 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_2 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_13 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_82 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_152 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_171 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_197 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_216 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_360 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_400 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_422 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_22 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_68 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_94 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_180 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_187 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_278 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_296 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_320 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_339 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_344 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_367 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_422 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_22 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_48 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_50 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_72 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_108 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_110 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_160 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_257 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_339 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_422 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_38 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_114 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_153 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_278 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_289 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_359 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_400 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_422 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_55 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_57 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_92 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_208 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_233 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_274 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_278 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_344 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_404 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_423 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_20 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_92 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_127 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_141 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_202 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_248 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_269 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_2 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_13 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_307 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_309 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_327 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_356 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_401 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_2 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_387 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_2 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_37 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_43 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_68 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_183 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_202 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_225 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_251 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_352 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_62 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_90 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_206 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_27 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_43 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_45 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_250 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_349 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_57 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_75 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_129 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_141 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_219 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_337 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_356 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_372 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_170 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_236 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_290 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_314 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_337 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_418 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_48 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_271 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_341 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_72 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_236 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_346 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_381 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_400 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_423 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_20 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_206 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_422 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_93 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_115 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_219 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_33 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_124 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_198 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_230 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_289 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_302 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_304 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_339 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_358 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_422 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_72 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_83 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_48_180 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_187 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_48_234 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_236 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_262 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_48_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_48_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_419 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_49_33 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_49_40 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_49_206 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_49_303 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_49_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_324 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_49_330 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_332 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_49_391 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_49_422 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_50_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_50_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_50_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_50_92 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_50_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_50_160 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_50_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_50_229 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_50_247 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_50_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_50_260 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_50_352 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_50_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_50_377 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_50_379 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_50_414 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_50_423 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_51_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_51_72 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_51_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_51_106 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_51_236 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_51_254 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_51_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_51_275 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_51_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_51_283 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_51_289 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_51_337 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_51_339 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_51_412 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_51_422 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_52_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_52_94 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_52_121 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_52_185 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_52_212 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_52_278 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_52_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_52_285 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_52_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_52_401 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_52_423 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_53_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_53_36 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_53_79 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_53_155 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_53_178 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_53_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_53_317 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_53_335 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_53_337 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_53_376 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_53_394 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_53_396 (.VDD(VPWR),
    .VSS(VGND));
endmodule
