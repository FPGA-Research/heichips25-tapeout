magic
tech ihp-sg13g2
magscale 1 2
timestamp 1752761838
<< metal1 >>
rect 1152 9848 41856 9872
rect 1152 9808 4928 9848
rect 4968 9808 5010 9848
rect 5050 9808 5092 9848
rect 5132 9808 5174 9848
rect 5214 9808 5256 9848
rect 5296 9808 20048 9848
rect 20088 9808 20130 9848
rect 20170 9808 20212 9848
rect 20252 9808 20294 9848
rect 20334 9808 20376 9848
rect 20416 9808 35168 9848
rect 35208 9808 35250 9848
rect 35290 9808 35332 9848
rect 35372 9808 35414 9848
rect 35454 9808 35496 9848
rect 35536 9808 41856 9848
rect 1152 9784 41856 9808
rect 4003 9680 4061 9681
rect 4003 9640 4012 9680
rect 4052 9640 4061 9680
rect 4003 9639 4061 9640
rect 5731 9680 5789 9681
rect 5731 9640 5740 9680
rect 5780 9640 5789 9680
rect 5731 9639 5789 9640
rect 9003 9680 9045 9689
rect 9003 9640 9004 9680
rect 9044 9640 9045 9680
rect 9003 9631 9045 9640
rect 10155 9680 10197 9689
rect 10155 9640 10156 9680
rect 10196 9640 10197 9680
rect 10155 9631 10197 9640
rect 10731 9680 10773 9689
rect 10731 9640 10732 9680
rect 10772 9640 10773 9680
rect 10731 9631 10773 9640
rect 14187 9680 14229 9689
rect 14187 9640 14188 9680
rect 14228 9640 14229 9680
rect 14187 9631 14229 9640
rect 17067 9680 17109 9689
rect 17067 9640 17068 9680
rect 17108 9640 17109 9680
rect 17067 9631 17109 9640
rect 18987 9680 19029 9689
rect 18987 9640 18988 9680
rect 19028 9640 19029 9680
rect 18987 9631 19029 9640
rect 22251 9680 22293 9689
rect 22251 9640 22252 9680
rect 22292 9640 22293 9680
rect 22251 9631 22293 9640
rect 29835 9680 29877 9689
rect 29835 9640 29836 9680
rect 29876 9640 29877 9680
rect 29835 9631 29877 9640
rect 30027 9680 30069 9689
rect 30027 9640 30028 9680
rect 30068 9640 30069 9680
rect 30027 9631 30069 9640
rect 30411 9680 30453 9689
rect 30411 9640 30412 9680
rect 30452 9640 30453 9680
rect 30411 9631 30453 9640
rect 30795 9680 30837 9689
rect 30795 9640 30796 9680
rect 30836 9640 30837 9680
rect 30795 9631 30837 9640
rect 41451 9680 41493 9689
rect 41451 9640 41452 9680
rect 41492 9640 41493 9680
rect 41451 9631 41493 9640
rect 3531 9596 3573 9605
rect 3531 9556 3532 9596
rect 3572 9556 3573 9596
rect 3531 9547 3573 9556
rect 1891 9512 1949 9513
rect 1891 9472 1900 9512
rect 1940 9472 1949 9512
rect 1891 9471 1949 9472
rect 3139 9512 3197 9513
rect 3139 9472 3148 9512
rect 3188 9472 3197 9512
rect 3139 9471 3197 9472
rect 3627 9512 3669 9521
rect 3627 9472 3628 9512
rect 3668 9472 3669 9512
rect 3627 9463 3669 9472
rect 3723 9512 3765 9521
rect 3723 9472 3724 9512
rect 3764 9472 3765 9512
rect 3723 9463 3765 9472
rect 3819 9512 3861 9521
rect 3819 9472 3820 9512
rect 3860 9472 3861 9512
rect 3819 9463 3861 9472
rect 4203 9512 4245 9521
rect 4203 9472 4204 9512
rect 4244 9472 4245 9512
rect 4203 9463 4245 9472
rect 4299 9512 4341 9521
rect 4299 9472 4300 9512
rect 4340 9472 4341 9512
rect 4299 9463 4341 9472
rect 4483 9512 4541 9513
rect 4483 9472 4492 9512
rect 4532 9472 4541 9512
rect 4483 9471 4541 9472
rect 4579 9512 4637 9513
rect 4579 9472 4588 9512
rect 4628 9472 4637 9512
rect 4579 9471 4637 9472
rect 4779 9512 4821 9521
rect 4779 9472 4780 9512
rect 4820 9472 4821 9512
rect 4779 9463 4821 9472
rect 4875 9512 4917 9521
rect 4875 9472 4876 9512
rect 4916 9472 4917 9512
rect 5259 9512 5301 9521
rect 4875 9463 4917 9472
rect 5032 9497 5074 9506
rect 5032 9457 5033 9497
rect 5073 9457 5074 9497
rect 5259 9472 5260 9512
rect 5300 9472 5301 9512
rect 5259 9463 5301 9472
rect 5355 9512 5397 9521
rect 5355 9472 5356 9512
rect 5396 9472 5397 9512
rect 5355 9463 5397 9472
rect 5451 9512 5493 9521
rect 5451 9472 5452 9512
rect 5492 9472 5493 9512
rect 5451 9463 5493 9472
rect 5547 9512 5589 9521
rect 5547 9472 5548 9512
rect 5588 9472 5589 9512
rect 5547 9463 5589 9472
rect 5835 9512 5877 9521
rect 5835 9472 5836 9512
rect 5876 9472 5877 9512
rect 5835 9463 5877 9472
rect 5931 9512 5973 9521
rect 5931 9472 5932 9512
rect 5972 9472 5973 9512
rect 5931 9463 5973 9472
rect 6027 9512 6069 9521
rect 6027 9472 6028 9512
rect 6068 9472 6069 9512
rect 6027 9463 6069 9472
rect 6211 9512 6269 9513
rect 6211 9472 6220 9512
rect 6260 9472 6269 9512
rect 6211 9471 6269 9472
rect 6411 9512 6453 9521
rect 6411 9472 6412 9512
rect 6452 9472 6453 9512
rect 6411 9463 6453 9472
rect 6891 9512 6933 9521
rect 6891 9472 6892 9512
rect 6932 9472 6933 9512
rect 6891 9463 6933 9472
rect 6987 9512 7029 9521
rect 6987 9472 6988 9512
rect 7028 9472 7029 9512
rect 6987 9463 7029 9472
rect 7267 9512 7325 9513
rect 7267 9472 7276 9512
rect 7316 9472 7325 9512
rect 7267 9471 7325 9472
rect 7555 9512 7613 9513
rect 7555 9472 7564 9512
rect 7604 9472 7613 9512
rect 7555 9471 7613 9472
rect 8803 9512 8861 9513
rect 8803 9472 8812 9512
rect 8852 9472 8861 9512
rect 8803 9471 8861 9472
rect 9483 9512 9525 9521
rect 9483 9472 9484 9512
rect 9524 9472 9525 9512
rect 9483 9463 9525 9472
rect 9579 9512 9621 9521
rect 9579 9472 9580 9512
rect 9620 9472 9621 9512
rect 9579 9463 9621 9472
rect 9859 9512 9917 9513
rect 9859 9472 9868 9512
rect 9908 9472 9917 9512
rect 9859 9471 9917 9472
rect 10915 9512 10973 9513
rect 10915 9472 10924 9512
rect 10964 9472 10973 9512
rect 10915 9471 10973 9472
rect 12163 9512 12221 9513
rect 12163 9472 12172 9512
rect 12212 9472 12221 9512
rect 12163 9471 12221 9472
rect 14947 9512 15005 9513
rect 14947 9472 14956 9512
rect 14996 9472 15005 9512
rect 14947 9471 15005 9472
rect 16195 9512 16253 9513
rect 16195 9472 16204 9512
rect 16244 9472 16253 9512
rect 16195 9471 16253 9472
rect 19171 9512 19229 9513
rect 19171 9472 19180 9512
rect 19220 9472 19229 9512
rect 19171 9471 19229 9472
rect 20419 9512 20477 9513
rect 20419 9472 20428 9512
rect 20468 9472 20477 9512
rect 20419 9471 20477 9472
rect 22723 9512 22781 9513
rect 22723 9472 22732 9512
rect 22772 9472 22781 9512
rect 22723 9471 22781 9472
rect 23971 9512 24029 9513
rect 23971 9472 23980 9512
rect 24020 9472 24029 9512
rect 23971 9471 24029 9472
rect 24355 9512 24413 9513
rect 24355 9472 24364 9512
rect 24404 9472 24413 9512
rect 24355 9471 24413 9472
rect 25603 9512 25661 9513
rect 25603 9472 25612 9512
rect 25652 9472 25661 9512
rect 25603 9471 25661 9472
rect 27139 9512 27197 9513
rect 27139 9472 27148 9512
rect 27188 9472 27197 9512
rect 27139 9471 27197 9472
rect 28387 9512 28445 9513
rect 28387 9472 28396 9512
rect 28436 9472 28445 9512
rect 28387 9471 28445 9472
rect 31171 9512 31229 9513
rect 31171 9472 31180 9512
rect 31220 9472 31229 9512
rect 31171 9471 31229 9472
rect 32419 9512 32477 9513
rect 32419 9472 32428 9512
rect 32468 9472 32477 9512
rect 32419 9471 32477 9472
rect 32899 9512 32957 9513
rect 32899 9472 32908 9512
rect 32948 9472 32957 9512
rect 32899 9471 32957 9472
rect 34147 9512 34205 9513
rect 34147 9472 34156 9512
rect 34196 9472 34205 9512
rect 34147 9471 34205 9472
rect 35011 9512 35069 9513
rect 35011 9472 35020 9512
rect 35060 9472 35069 9512
rect 35011 9471 35069 9472
rect 36259 9512 36317 9513
rect 36259 9472 36268 9512
rect 36308 9472 36317 9512
rect 36259 9471 36317 9472
rect 38467 9512 38525 9513
rect 38467 9472 38476 9512
rect 38516 9472 38525 9512
rect 38467 9471 38525 9472
rect 39715 9512 39773 9513
rect 39715 9472 39724 9512
rect 39764 9472 39773 9512
rect 39715 9471 39773 9472
rect 5032 9448 5074 9457
rect 10339 9428 10397 9429
rect 10339 9388 10348 9428
rect 10388 9388 10397 9428
rect 10339 9387 10397 9388
rect 10531 9428 10589 9429
rect 10531 9388 10540 9428
rect 10580 9388 10589 9428
rect 10531 9387 10589 9388
rect 14371 9428 14429 9429
rect 14371 9388 14380 9428
rect 14420 9388 14429 9428
rect 14371 9387 14429 9388
rect 16867 9428 16925 9429
rect 16867 9388 16876 9428
rect 16916 9388 16925 9428
rect 16867 9387 16925 9388
rect 18787 9428 18845 9429
rect 18787 9388 18796 9428
rect 18836 9388 18845 9428
rect 18787 9387 18845 9388
rect 22435 9428 22493 9429
rect 22435 9388 22444 9428
rect 22484 9388 22493 9428
rect 22435 9387 22493 9388
rect 29635 9428 29693 9429
rect 29635 9388 29644 9428
rect 29684 9388 29693 9428
rect 29635 9387 29693 9388
rect 30211 9428 30269 9429
rect 30211 9388 30220 9428
rect 30260 9388 30269 9428
rect 30211 9387 30269 9388
rect 30595 9428 30653 9429
rect 30595 9388 30604 9428
rect 30644 9388 30653 9428
rect 30595 9387 30653 9388
rect 30979 9428 31037 9429
rect 30979 9388 30988 9428
rect 31028 9388 31037 9428
rect 30979 9387 31037 9388
rect 37219 9428 37277 9429
rect 37219 9388 37228 9428
rect 37268 9388 37277 9428
rect 37219 9387 37277 9388
rect 37795 9428 37853 9429
rect 37795 9388 37804 9428
rect 37844 9388 37853 9428
rect 37795 9387 37853 9388
rect 40867 9428 40925 9429
rect 40867 9388 40876 9428
rect 40916 9388 40925 9428
rect 40867 9387 40925 9388
rect 41251 9428 41309 9429
rect 41251 9388 41260 9428
rect 41300 9388 41309 9428
rect 41251 9387 41309 9388
rect 3339 9344 3381 9353
rect 3339 9304 3340 9344
rect 3380 9304 3381 9344
rect 3339 9295 3381 9304
rect 41067 9344 41109 9353
rect 41067 9304 41068 9344
rect 41108 9304 41109 9344
rect 41067 9295 41109 9304
rect 4491 9260 4533 9269
rect 4491 9220 4492 9260
rect 4532 9220 4533 9260
rect 4491 9211 4533 9220
rect 6315 9260 6357 9269
rect 6315 9220 6316 9260
rect 6356 9220 6357 9260
rect 6315 9211 6357 9220
rect 6595 9260 6653 9261
rect 6595 9220 6604 9260
rect 6644 9220 6653 9260
rect 6595 9219 6653 9220
rect 9187 9260 9245 9261
rect 9187 9220 9196 9260
rect 9236 9220 9245 9260
rect 9187 9219 9245 9220
rect 12363 9260 12405 9269
rect 12363 9220 12364 9260
rect 12404 9220 12405 9260
rect 12363 9211 12405 9220
rect 16395 9260 16437 9269
rect 16395 9220 16396 9260
rect 16436 9220 16437 9260
rect 16395 9211 16437 9220
rect 20619 9260 20661 9269
rect 20619 9220 20620 9260
rect 20660 9220 20661 9260
rect 20619 9211 20661 9220
rect 24171 9260 24213 9269
rect 24171 9220 24172 9260
rect 24212 9220 24213 9260
rect 24171 9211 24213 9220
rect 25803 9260 25845 9269
rect 25803 9220 25804 9260
rect 25844 9220 25845 9260
rect 25803 9211 25845 9220
rect 26955 9260 26997 9269
rect 26955 9220 26956 9260
rect 26996 9220 26997 9260
rect 26955 9211 26997 9220
rect 32619 9260 32661 9269
rect 32619 9220 32620 9260
rect 32660 9220 32661 9260
rect 32619 9211 32661 9220
rect 34347 9260 34389 9269
rect 34347 9220 34348 9260
rect 34388 9220 34389 9260
rect 34347 9211 34389 9220
rect 36459 9260 36501 9269
rect 36459 9220 36460 9260
rect 36500 9220 36501 9260
rect 36459 9211 36501 9220
rect 37035 9260 37077 9269
rect 37035 9220 37036 9260
rect 37076 9220 37077 9260
rect 37035 9211 37077 9220
rect 37611 9260 37653 9269
rect 37611 9220 37612 9260
rect 37652 9220 37653 9260
rect 37611 9211 37653 9220
rect 38283 9260 38325 9269
rect 38283 9220 38284 9260
rect 38324 9220 38325 9260
rect 38283 9211 38325 9220
rect 1152 9092 41856 9116
rect 1152 9052 3688 9092
rect 3728 9052 3770 9092
rect 3810 9052 3852 9092
rect 3892 9052 3934 9092
rect 3974 9052 4016 9092
rect 4056 9052 18808 9092
rect 18848 9052 18890 9092
rect 18930 9052 18972 9092
rect 19012 9052 19054 9092
rect 19094 9052 19136 9092
rect 19176 9052 33928 9092
rect 33968 9052 34010 9092
rect 34050 9052 34092 9092
rect 34132 9052 34174 9092
rect 34214 9052 34256 9092
rect 34296 9052 41856 9092
rect 1152 9028 41856 9052
rect 3531 8924 3573 8933
rect 3531 8884 3532 8924
rect 3572 8884 3573 8924
rect 3531 8875 3573 8884
rect 5163 8924 5205 8933
rect 5163 8884 5164 8924
rect 5204 8884 5205 8924
rect 5163 8875 5205 8884
rect 1707 8840 1749 8849
rect 1707 8800 1708 8840
rect 1748 8800 1749 8840
rect 1707 8791 1749 8800
rect 1899 8840 1941 8849
rect 1899 8800 1900 8840
rect 1940 8800 1941 8840
rect 1899 8791 1941 8800
rect 8619 8840 8661 8849
rect 8619 8800 8620 8840
rect 8660 8800 8661 8840
rect 8619 8791 8661 8800
rect 18411 8840 18453 8849
rect 18411 8800 18412 8840
rect 18452 8800 18453 8840
rect 18411 8791 18453 8800
rect 24555 8840 24597 8849
rect 24555 8800 24556 8840
rect 24596 8800 24597 8840
rect 24555 8791 24597 8800
rect 25035 8840 25077 8849
rect 25035 8800 25036 8840
rect 25076 8800 25077 8840
rect 25035 8791 25077 8800
rect 25515 8840 25557 8849
rect 25515 8800 25516 8840
rect 25556 8800 25557 8840
rect 25515 8791 25557 8800
rect 34339 8840 34397 8841
rect 34339 8800 34348 8840
rect 34388 8800 34397 8840
rect 34339 8799 34397 8800
rect 40299 8840 40341 8849
rect 40299 8800 40300 8840
rect 40340 8800 40341 8840
rect 40299 8791 40341 8800
rect 40683 8840 40725 8849
rect 40683 8800 40684 8840
rect 40724 8800 40725 8840
rect 40683 8791 40725 8800
rect 41451 8840 41493 8849
rect 41451 8800 41452 8840
rect 41492 8800 41493 8840
rect 41451 8791 41493 8800
rect 8419 8756 8477 8757
rect 8419 8716 8428 8756
rect 8468 8716 8477 8756
rect 22923 8756 22965 8765
rect 8419 8715 8477 8716
rect 3331 8714 3389 8715
rect 1707 8672 1749 8681
rect 3331 8674 3340 8714
rect 3380 8674 3389 8714
rect 11403 8714 11445 8723
rect 7659 8686 7701 8695
rect 3331 8673 3389 8674
rect 1707 8632 1708 8672
rect 1748 8632 1749 8672
rect 1707 8623 1749 8632
rect 2083 8672 2141 8673
rect 2083 8632 2092 8672
rect 2132 8632 2141 8672
rect 2083 8631 2141 8632
rect 3715 8672 3773 8673
rect 3715 8632 3724 8672
rect 3764 8632 3773 8672
rect 3715 8631 3773 8632
rect 4963 8672 5021 8673
rect 4963 8632 4972 8672
rect 5012 8632 5021 8672
rect 4963 8631 5021 8632
rect 5451 8672 5493 8681
rect 5451 8632 5452 8672
rect 5492 8632 5493 8672
rect 5451 8623 5493 8632
rect 5547 8672 5589 8681
rect 5547 8632 5548 8672
rect 5588 8632 5589 8672
rect 5547 8623 5589 8632
rect 6123 8672 6165 8681
rect 6123 8632 6124 8672
rect 6164 8632 6165 8672
rect 6123 8623 6165 8632
rect 6219 8672 6261 8681
rect 6219 8632 6220 8672
rect 6260 8632 6261 8672
rect 6219 8623 6261 8632
rect 6603 8672 6645 8681
rect 6603 8632 6604 8672
rect 6644 8632 6645 8672
rect 6603 8623 6645 8632
rect 6699 8672 6741 8681
rect 6699 8632 6700 8672
rect 6740 8632 6741 8672
rect 6699 8623 6741 8632
rect 7171 8672 7229 8673
rect 7171 8632 7180 8672
rect 7220 8632 7229 8672
rect 7659 8646 7660 8686
rect 7700 8646 7701 8686
rect 7659 8637 7701 8646
rect 8803 8672 8861 8673
rect 7171 8631 7229 8632
rect 8803 8632 8812 8672
rect 8852 8632 8861 8672
rect 8803 8631 8861 8632
rect 10051 8672 10109 8673
rect 10051 8632 10060 8672
rect 10100 8632 10109 8672
rect 10051 8631 10109 8632
rect 10827 8672 10869 8681
rect 10827 8632 10828 8672
rect 10868 8632 10869 8672
rect 10827 8623 10869 8632
rect 10923 8672 10965 8681
rect 10923 8632 10924 8672
rect 10964 8632 10965 8672
rect 10923 8623 10965 8632
rect 11307 8672 11349 8681
rect 11307 8632 11308 8672
rect 11348 8632 11349 8672
rect 11403 8674 11404 8714
rect 11444 8674 11445 8714
rect 20283 8714 20325 8723
rect 11403 8665 11445 8674
rect 12363 8686 12405 8695
rect 11875 8672 11933 8673
rect 11307 8623 11349 8632
rect 11875 8632 11884 8672
rect 11924 8632 11933 8672
rect 12363 8646 12364 8686
rect 12404 8646 12405 8686
rect 16299 8686 16341 8695
rect 12363 8637 12405 8646
rect 13027 8672 13085 8673
rect 11875 8631 11933 8632
rect 13027 8632 13036 8672
rect 13076 8632 13085 8672
rect 13027 8631 13085 8632
rect 14275 8672 14333 8673
rect 14275 8632 14284 8672
rect 14324 8632 14333 8672
rect 14275 8631 14333 8632
rect 14763 8672 14805 8681
rect 14763 8632 14764 8672
rect 14804 8632 14805 8672
rect 14763 8623 14805 8632
rect 14859 8672 14901 8681
rect 14859 8632 14860 8672
rect 14900 8632 14901 8672
rect 14859 8623 14901 8632
rect 15243 8672 15285 8681
rect 15243 8632 15244 8672
rect 15284 8632 15285 8672
rect 15243 8623 15285 8632
rect 15339 8672 15381 8681
rect 15339 8632 15340 8672
rect 15380 8632 15381 8672
rect 15339 8623 15381 8632
rect 15811 8672 15869 8673
rect 15811 8632 15820 8672
rect 15860 8632 15869 8672
rect 16299 8646 16300 8686
rect 16340 8646 16341 8686
rect 16299 8637 16341 8646
rect 16963 8672 17021 8673
rect 15811 8631 15869 8632
rect 16963 8632 16972 8672
rect 17012 8632 17021 8672
rect 16963 8631 17021 8632
rect 18211 8672 18269 8673
rect 18211 8632 18220 8672
rect 18260 8632 18269 8672
rect 18211 8631 18269 8632
rect 18699 8672 18741 8681
rect 18699 8632 18700 8672
rect 18740 8632 18741 8672
rect 18699 8623 18741 8632
rect 18795 8672 18837 8681
rect 18795 8632 18796 8672
rect 18836 8632 18837 8672
rect 18795 8623 18837 8632
rect 19179 8672 19221 8681
rect 19179 8632 19180 8672
rect 19220 8632 19221 8672
rect 19179 8623 19221 8632
rect 19275 8672 19317 8681
rect 20283 8674 20284 8714
rect 20324 8674 20325 8714
rect 22923 8716 22924 8756
rect 22964 8716 22965 8756
rect 22923 8707 22965 8716
rect 23019 8756 23061 8765
rect 23019 8716 23020 8756
rect 23060 8716 23061 8756
rect 24739 8756 24797 8757
rect 23019 8707 23061 8716
rect 24027 8714 24069 8723
rect 24739 8716 24748 8756
rect 24788 8716 24797 8756
rect 24739 8715 24797 8716
rect 25219 8756 25277 8757
rect 25219 8716 25228 8756
rect 25268 8716 25277 8756
rect 25219 8715 25277 8716
rect 25699 8756 25757 8757
rect 25699 8716 25708 8756
rect 25748 8716 25757 8756
rect 25699 8715 25757 8716
rect 26475 8756 26517 8765
rect 26475 8716 26476 8756
rect 26516 8716 26517 8756
rect 19275 8632 19276 8672
rect 19316 8632 19317 8672
rect 19275 8623 19317 8632
rect 19747 8672 19805 8673
rect 19747 8632 19756 8672
rect 19796 8632 19805 8672
rect 20283 8665 20325 8674
rect 20707 8672 20765 8673
rect 19747 8631 19805 8632
rect 20707 8632 20716 8672
rect 20756 8632 20765 8672
rect 20707 8631 20765 8632
rect 21955 8672 22013 8673
rect 21955 8632 21964 8672
rect 22004 8632 22013 8672
rect 21955 8631 22013 8632
rect 22443 8672 22485 8681
rect 22443 8632 22444 8672
rect 22484 8632 22485 8672
rect 22443 8623 22485 8632
rect 22539 8672 22581 8681
rect 24027 8674 24028 8714
rect 24068 8674 24069 8714
rect 26475 8707 26517 8716
rect 26571 8756 26613 8765
rect 26571 8716 26572 8756
rect 26612 8716 26613 8756
rect 26571 8707 26613 8716
rect 28099 8756 28157 8757
rect 28099 8716 28108 8756
rect 28148 8716 28157 8756
rect 28099 8715 28157 8716
rect 29547 8756 29589 8765
rect 29547 8716 29548 8756
rect 29588 8716 29589 8756
rect 29547 8707 29589 8716
rect 29643 8756 29685 8765
rect 29643 8716 29644 8756
rect 29684 8716 29685 8756
rect 29643 8707 29685 8716
rect 31171 8756 31229 8757
rect 31171 8716 31180 8756
rect 31220 8716 31229 8756
rect 31171 8715 31229 8716
rect 31555 8756 31613 8757
rect 31555 8716 31564 8756
rect 31604 8716 31613 8756
rect 31555 8715 31613 8716
rect 31939 8756 31997 8757
rect 31939 8716 31948 8756
rect 31988 8716 31997 8756
rect 31939 8715 31997 8716
rect 32811 8756 32853 8765
rect 32811 8716 32812 8756
rect 32852 8716 32853 8756
rect 32811 8707 32853 8716
rect 36267 8756 36309 8765
rect 36267 8716 36268 8756
rect 36308 8716 36309 8756
rect 36267 8707 36309 8716
rect 39907 8756 39965 8757
rect 39907 8716 39916 8756
rect 39956 8716 39965 8756
rect 39907 8715 39965 8716
rect 40099 8756 40157 8757
rect 40099 8716 40108 8756
rect 40148 8716 40157 8756
rect 40099 8715 40157 8716
rect 40483 8756 40541 8757
rect 40483 8716 40492 8756
rect 40532 8716 40541 8756
rect 40483 8715 40541 8716
rect 40867 8756 40925 8757
rect 40867 8716 40876 8756
rect 40916 8716 40925 8756
rect 40867 8715 40925 8716
rect 41251 8756 41309 8757
rect 41251 8716 41260 8756
rect 41300 8716 41309 8756
rect 41251 8715 41309 8716
rect 27531 8686 27573 8695
rect 22539 8632 22540 8672
rect 22580 8632 22581 8672
rect 22539 8623 22581 8632
rect 23491 8672 23549 8673
rect 23491 8632 23500 8672
rect 23540 8632 23549 8672
rect 24027 8665 24069 8674
rect 25995 8672 26037 8681
rect 23491 8631 23549 8632
rect 25995 8632 25996 8672
rect 26036 8632 26037 8672
rect 25995 8623 26037 8632
rect 26091 8672 26133 8681
rect 26091 8632 26092 8672
rect 26132 8632 26133 8672
rect 26091 8623 26133 8632
rect 27043 8672 27101 8673
rect 27043 8632 27052 8672
rect 27092 8632 27101 8672
rect 27531 8646 27532 8686
rect 27572 8646 27573 8686
rect 30603 8686 30645 8695
rect 27531 8637 27573 8646
rect 29067 8672 29109 8681
rect 27043 8631 27101 8632
rect 29067 8632 29068 8672
rect 29108 8632 29109 8672
rect 29067 8623 29109 8632
rect 29163 8672 29205 8681
rect 29163 8632 29164 8672
rect 29204 8632 29205 8672
rect 29163 8623 29205 8632
rect 30115 8672 30173 8673
rect 30115 8632 30124 8672
rect 30164 8632 30173 8672
rect 30603 8646 30604 8686
rect 30644 8646 30645 8686
rect 33867 8686 33909 8695
rect 30603 8637 30645 8646
rect 32331 8672 32373 8681
rect 30115 8631 30173 8632
rect 32331 8632 32332 8672
rect 32372 8632 32373 8672
rect 32331 8623 32373 8632
rect 32427 8672 32469 8681
rect 32427 8632 32428 8672
rect 32468 8632 32469 8672
rect 32427 8623 32469 8632
rect 32907 8672 32949 8681
rect 32907 8632 32908 8672
rect 32948 8632 32949 8672
rect 32907 8623 32949 8632
rect 33379 8672 33437 8673
rect 33379 8632 33388 8672
rect 33428 8632 33437 8672
rect 33867 8646 33868 8686
rect 33908 8646 33909 8686
rect 33867 8637 33909 8646
rect 34635 8672 34677 8681
rect 33379 8631 33437 8632
rect 34635 8632 34636 8672
rect 34676 8632 34677 8672
rect 34635 8623 34677 8632
rect 34731 8672 34773 8681
rect 34731 8632 34732 8672
rect 34772 8632 34773 8672
rect 34731 8623 34773 8632
rect 35011 8672 35069 8673
rect 35011 8632 35020 8672
rect 35060 8632 35069 8672
rect 35011 8631 35069 8632
rect 35691 8672 35733 8681
rect 35691 8632 35692 8672
rect 35732 8632 35733 8672
rect 35691 8623 35733 8632
rect 35787 8672 35829 8681
rect 35787 8632 35788 8672
rect 35828 8632 35829 8672
rect 35787 8623 35829 8632
rect 36171 8672 36213 8681
rect 37227 8677 37269 8686
rect 36171 8632 36172 8672
rect 36212 8632 36213 8672
rect 36171 8623 36213 8632
rect 36739 8672 36797 8673
rect 36739 8632 36748 8672
rect 36788 8632 36797 8672
rect 36739 8631 36797 8632
rect 37227 8637 37228 8677
rect 37268 8637 37269 8677
rect 37227 8628 37269 8637
rect 37795 8672 37853 8673
rect 37795 8632 37804 8672
rect 37844 8632 37853 8672
rect 37795 8631 37853 8632
rect 39043 8672 39101 8673
rect 39043 8632 39052 8672
rect 39092 8632 39101 8672
rect 39043 8631 39101 8632
rect 7851 8588 7893 8597
rect 7851 8548 7852 8588
rect 7892 8548 7893 8588
rect 7851 8539 7893 8548
rect 10251 8588 10293 8597
rect 10251 8548 10252 8588
rect 10292 8548 10293 8588
rect 10251 8539 10293 8548
rect 14475 8588 14517 8597
rect 14475 8548 14476 8588
rect 14516 8548 14517 8588
rect 14475 8539 14517 8548
rect 16491 8588 16533 8597
rect 16491 8548 16492 8588
rect 16532 8548 16533 8588
rect 16491 8539 16533 8548
rect 22155 8588 22197 8597
rect 22155 8548 22156 8588
rect 22196 8548 22197 8588
rect 22155 8539 22197 8548
rect 24171 8588 24213 8597
rect 24171 8548 24172 8588
rect 24212 8548 24213 8588
rect 24171 8539 24213 8548
rect 37419 8588 37461 8597
rect 37419 8548 37420 8588
rect 37460 8548 37461 8588
rect 37419 8539 37461 8548
rect 3531 8504 3573 8513
rect 3531 8464 3532 8504
rect 3572 8464 3573 8504
rect 3531 8455 3573 8464
rect 5731 8504 5789 8505
rect 5731 8464 5740 8504
rect 5780 8464 5789 8504
rect 5731 8463 5789 8464
rect 12555 8504 12597 8513
rect 12555 8464 12556 8504
rect 12596 8464 12597 8504
rect 12555 8455 12597 8464
rect 20427 8504 20469 8513
rect 20427 8464 20428 8504
rect 20468 8464 20469 8504
rect 20427 8455 20469 8464
rect 27723 8504 27765 8513
rect 27723 8464 27724 8504
rect 27764 8464 27765 8504
rect 27723 8455 27765 8464
rect 27915 8504 27957 8513
rect 27915 8464 27916 8504
rect 27956 8464 27957 8504
rect 30987 8504 31029 8513
rect 27915 8455 27957 8464
rect 30795 8462 30837 8471
rect 30795 8422 30796 8462
rect 30836 8422 30837 8462
rect 30987 8464 30988 8504
rect 31028 8464 31029 8504
rect 30987 8455 31029 8464
rect 31371 8504 31413 8513
rect 31371 8464 31372 8504
rect 31412 8464 31413 8504
rect 31371 8455 31413 8464
rect 31755 8504 31797 8513
rect 31755 8464 31756 8504
rect 31796 8464 31797 8504
rect 31755 8455 31797 8464
rect 34059 8504 34101 8513
rect 34059 8464 34060 8504
rect 34100 8464 34101 8504
rect 34059 8455 34101 8464
rect 37611 8504 37653 8513
rect 37611 8464 37612 8504
rect 37652 8464 37653 8504
rect 37611 8455 37653 8464
rect 39723 8504 39765 8513
rect 39723 8464 39724 8504
rect 39764 8464 39765 8504
rect 39723 8455 39765 8464
rect 41067 8504 41109 8513
rect 41067 8464 41068 8504
rect 41108 8464 41109 8504
rect 41067 8455 41109 8464
rect 30795 8413 30837 8422
rect 1152 8336 41856 8360
rect 1152 8296 4928 8336
rect 4968 8296 5010 8336
rect 5050 8296 5092 8336
rect 5132 8296 5174 8336
rect 5214 8296 5256 8336
rect 5296 8296 20048 8336
rect 20088 8296 20130 8336
rect 20170 8296 20212 8336
rect 20252 8296 20294 8336
rect 20334 8296 20376 8336
rect 20416 8296 35168 8336
rect 35208 8296 35250 8336
rect 35290 8296 35332 8336
rect 35372 8296 35414 8336
rect 35454 8296 35496 8336
rect 35536 8296 41856 8336
rect 1152 8272 41856 8296
rect 19275 8210 19317 8219
rect 3339 8168 3381 8177
rect 3339 8128 3340 8168
rect 3380 8128 3381 8168
rect 3339 8119 3381 8128
rect 3811 8168 3869 8169
rect 3811 8128 3820 8168
rect 3860 8128 3869 8168
rect 3811 8127 3869 8128
rect 7659 8168 7701 8177
rect 7659 8128 7660 8168
rect 7700 8128 7701 8168
rect 7659 8119 7701 8128
rect 9579 8168 9621 8177
rect 9579 8128 9580 8168
rect 9620 8128 9621 8168
rect 9579 8119 9621 8128
rect 11499 8168 11541 8177
rect 11499 8128 11500 8168
rect 11540 8128 11541 8168
rect 11499 8119 11541 8128
rect 11883 8168 11925 8177
rect 11883 8128 11884 8168
rect 11924 8128 11925 8168
rect 11883 8119 11925 8128
rect 17067 8168 17109 8177
rect 17067 8128 17068 8168
rect 17108 8128 17109 8168
rect 19275 8170 19276 8210
rect 19316 8170 19317 8210
rect 19275 8161 19317 8170
rect 19459 8168 19517 8169
rect 17067 8119 17109 8128
rect 19459 8128 19468 8168
rect 19508 8128 19517 8168
rect 19459 8127 19517 8128
rect 20043 8168 20085 8177
rect 20043 8128 20044 8168
rect 20084 8128 20085 8168
rect 20043 8119 20085 8128
rect 22731 8168 22773 8177
rect 22731 8128 22732 8168
rect 22772 8128 22773 8168
rect 22731 8119 22773 8128
rect 22923 8168 22965 8177
rect 22923 8128 22924 8168
rect 22964 8128 22965 8168
rect 22923 8119 22965 8128
rect 27531 8168 27573 8177
rect 27531 8128 27532 8168
rect 27572 8128 27573 8168
rect 27531 8119 27573 8128
rect 29451 8168 29493 8177
rect 29451 8128 29452 8168
rect 29492 8128 29493 8168
rect 29451 8119 29493 8128
rect 31179 8168 31221 8177
rect 31179 8128 31180 8168
rect 31220 8128 31221 8168
rect 31179 8119 31221 8128
rect 32235 8168 32277 8177
rect 32235 8128 32236 8168
rect 32276 8128 32277 8168
rect 32235 8119 32277 8128
rect 34731 8168 34773 8177
rect 34731 8128 34732 8168
rect 34772 8128 34773 8168
rect 34731 8119 34773 8128
rect 37995 8168 38037 8177
rect 37995 8128 37996 8168
rect 38036 8128 38037 8168
rect 37995 8119 38037 8128
rect 40011 8168 40053 8177
rect 40011 8128 40012 8168
rect 40052 8128 40053 8168
rect 40011 8119 40053 8128
rect 40683 8168 40725 8177
rect 40683 8128 40684 8168
rect 40724 8128 40725 8168
rect 40683 8119 40725 8128
rect 41451 8168 41493 8177
rect 41451 8128 41452 8168
rect 41492 8128 41493 8168
rect 41451 8119 41493 8128
rect 14187 8084 14229 8093
rect 14187 8044 14188 8084
rect 14228 8044 14229 8084
rect 14187 8035 14229 8044
rect 16299 8084 16341 8093
rect 16299 8044 16300 8084
rect 16340 8044 16341 8084
rect 16299 8035 16341 8044
rect 1891 8000 1949 8001
rect 1891 7960 1900 8000
rect 1940 7960 1949 8000
rect 1891 7959 1949 7960
rect 3139 8000 3197 8001
rect 3139 7960 3148 8000
rect 3188 7960 3197 8000
rect 3139 7959 3197 7960
rect 3723 8000 3765 8009
rect 3723 7960 3724 8000
rect 3764 7960 3765 8000
rect 3723 7951 3765 7960
rect 3915 8000 3957 8009
rect 4291 8007 4349 8008
rect 3915 7960 3916 8000
rect 3956 7960 3957 8000
rect 3915 7951 3957 7960
rect 4003 8000 4061 8001
rect 4003 7960 4012 8000
rect 4052 7960 4061 8000
rect 4291 7967 4300 8007
rect 4340 7967 4349 8007
rect 4291 7966 4349 7967
rect 4587 8000 4629 8009
rect 4003 7959 4061 7960
rect 4587 7960 4588 8000
rect 4628 7960 4629 8000
rect 4587 7951 4629 7960
rect 4683 8000 4725 8009
rect 4683 7960 4684 8000
rect 4724 7960 4725 8000
rect 4683 7951 4725 7960
rect 5355 8000 5397 8009
rect 5355 7960 5356 8000
rect 5396 7960 5397 8000
rect 5355 7951 5397 7960
rect 5451 8000 5493 8009
rect 5451 7960 5452 8000
rect 5492 7960 5493 8000
rect 5451 7951 5493 7960
rect 5547 8000 5589 8009
rect 5547 7960 5548 8000
rect 5588 7960 5589 8000
rect 5547 7951 5589 7960
rect 5643 8000 5685 8009
rect 5643 7960 5644 8000
rect 5684 7960 5685 8000
rect 5643 7951 5685 7960
rect 5931 8000 5973 8009
rect 5931 7960 5932 8000
rect 5972 7960 5973 8000
rect 5931 7951 5973 7960
rect 6027 8000 6069 8009
rect 6027 7960 6028 8000
rect 6068 7960 6069 8000
rect 6027 7951 6069 7960
rect 6411 8000 6453 8009
rect 6411 7960 6412 8000
rect 6452 7960 6453 8000
rect 6411 7951 6453 7960
rect 6979 8000 7037 8001
rect 6979 7960 6988 8000
rect 7028 7960 7037 8000
rect 6979 7959 7037 7960
rect 7467 7995 7509 8004
rect 7467 7955 7468 7995
rect 7508 7955 7509 7995
rect 9763 8000 9821 8001
rect 9763 7960 9772 8000
rect 9812 7960 9821 8000
rect 9763 7959 9821 7960
rect 11011 8000 11069 8001
rect 11011 7960 11020 8000
rect 11060 7960 11069 8000
rect 11011 7959 11069 7960
rect 12739 8000 12797 8001
rect 12739 7960 12748 8000
rect 12788 7960 12797 8000
rect 12739 7959 12797 7960
rect 13987 8000 14045 8001
rect 13987 7960 13996 8000
rect 14036 7960 14045 8000
rect 13987 7959 14045 7960
rect 14571 8000 14613 8009
rect 14571 7960 14572 8000
rect 14612 7960 14613 8000
rect 7467 7946 7509 7955
rect 14571 7951 14613 7960
rect 14667 8000 14709 8009
rect 14667 7960 14668 8000
rect 14708 7960 14709 8000
rect 14667 7951 14709 7960
rect 15147 8000 15189 8009
rect 15147 7960 15148 8000
rect 15188 7960 15189 8000
rect 17547 8000 17589 8009
rect 15147 7951 15189 7960
rect 16107 7986 16149 7995
rect 15619 7958 15677 7959
rect 6507 7916 6549 7925
rect 6507 7876 6508 7916
rect 6548 7876 6549 7916
rect 6507 7867 6549 7876
rect 9379 7916 9437 7917
rect 9379 7876 9388 7916
rect 9428 7876 9437 7916
rect 9379 7875 9437 7876
rect 11683 7916 11741 7917
rect 11683 7876 11692 7916
rect 11732 7876 11741 7916
rect 11683 7875 11741 7876
rect 12067 7916 12125 7917
rect 12067 7876 12076 7916
rect 12116 7876 12125 7916
rect 12067 7875 12125 7876
rect 15051 7916 15093 7925
rect 15619 7918 15628 7958
rect 15668 7918 15677 7958
rect 16107 7946 16108 7986
rect 16148 7946 16149 7986
rect 17547 7960 17548 8000
rect 17588 7960 17589 8000
rect 17547 7951 17589 7960
rect 17643 8000 17685 8009
rect 17643 7960 17644 8000
rect 17684 7960 17685 8000
rect 17643 7951 17685 7960
rect 18123 8000 18165 8009
rect 18123 7960 18124 8000
rect 18164 7960 18165 8000
rect 18123 7951 18165 7960
rect 18595 8000 18653 8001
rect 18595 7960 18604 8000
rect 18644 7960 18653 8000
rect 21003 8000 21045 8009
rect 18595 7959 18653 7960
rect 19131 7958 19173 7967
rect 16107 7937 16149 7946
rect 15619 7917 15677 7918
rect 15051 7876 15052 7916
rect 15092 7876 15093 7916
rect 15051 7867 15093 7876
rect 16867 7916 16925 7917
rect 16867 7876 16876 7916
rect 16916 7876 16925 7916
rect 16867 7875 16925 7876
rect 18027 7916 18069 7925
rect 18027 7876 18028 7916
rect 18068 7876 18069 7916
rect 19131 7918 19132 7958
rect 19172 7918 19173 7958
rect 21003 7960 21004 8000
rect 21044 7960 21045 8000
rect 21003 7951 21045 7960
rect 21099 8000 21141 8009
rect 21099 7960 21100 8000
rect 21140 7960 21141 8000
rect 21099 7951 21141 7960
rect 21579 8000 21621 8009
rect 21579 7960 21580 8000
rect 21620 7960 21621 8000
rect 21579 7951 21621 7960
rect 22051 8000 22109 8001
rect 22051 7960 22060 8000
rect 22100 7960 22109 8000
rect 24067 8000 24125 8001
rect 22051 7959 22109 7960
rect 22587 7958 22629 7967
rect 24067 7960 24076 8000
rect 24116 7960 24125 8000
rect 24067 7959 24125 7960
rect 25315 8000 25373 8001
rect 25315 7960 25324 8000
rect 25364 7960 25373 8000
rect 25315 7959 25373 7960
rect 25803 8000 25845 8009
rect 25803 7960 25804 8000
rect 25844 7960 25845 8000
rect 19131 7909 19173 7918
rect 20227 7916 20285 7917
rect 18027 7867 18069 7876
rect 20227 7876 20236 7916
rect 20276 7876 20285 7916
rect 20227 7875 20285 7876
rect 21483 7916 21525 7925
rect 21483 7876 21484 7916
rect 21524 7876 21525 7916
rect 22587 7918 22588 7958
rect 22628 7918 22629 7958
rect 25803 7951 25845 7960
rect 25899 8000 25941 8009
rect 25899 7960 25900 8000
rect 25940 7960 25941 8000
rect 25899 7951 25941 7960
rect 26283 8000 26325 8009
rect 26283 7960 26284 8000
rect 26324 7960 26325 8000
rect 26283 7951 26325 7960
rect 26379 8000 26421 8009
rect 26379 7960 26380 8000
rect 26420 7960 26421 8000
rect 26379 7951 26421 7960
rect 26851 8000 26909 8001
rect 26851 7960 26860 8000
rect 26900 7960 26909 8000
rect 28003 8000 28061 8001
rect 26851 7959 26909 7960
rect 27387 7958 27429 7967
rect 28003 7960 28012 8000
rect 28052 7960 28061 8000
rect 28003 7959 28061 7960
rect 29251 8000 29309 8001
rect 29251 7960 29260 8000
rect 29300 7960 29309 8000
rect 29251 7959 29309 7960
rect 29731 8000 29789 8001
rect 29731 7960 29740 8000
rect 29780 7960 29789 8000
rect 29731 7959 29789 7960
rect 30979 8000 31037 8001
rect 30979 7960 30988 8000
rect 31028 7960 31037 8000
rect 30979 7959 31037 7960
rect 33283 8000 33341 8001
rect 33283 7960 33292 8000
rect 33332 7960 33341 8000
rect 33283 7959 33341 7960
rect 34531 8000 34589 8001
rect 34531 7960 34540 8000
rect 34580 7960 34589 8000
rect 34531 7959 34589 7960
rect 36267 8000 36309 8009
rect 36267 7960 36268 8000
rect 36308 7960 36309 8000
rect 22587 7909 22629 7918
rect 27387 7918 27388 7958
rect 27428 7918 27429 7958
rect 36267 7951 36309 7960
rect 36363 8000 36405 8009
rect 36363 7960 36364 8000
rect 36404 7960 36405 8000
rect 36363 7951 36405 7960
rect 37315 8000 37373 8001
rect 37315 7960 37324 8000
rect 37364 7960 37373 8000
rect 38283 8000 38325 8009
rect 37315 7959 37373 7960
rect 37851 7990 37893 7999
rect 37851 7950 37852 7990
rect 37892 7950 37893 7990
rect 38283 7960 38284 8000
rect 38324 7960 38325 8000
rect 38283 7951 38325 7960
rect 38379 8000 38421 8009
rect 38379 7960 38380 8000
rect 38420 7960 38421 8000
rect 38379 7951 38421 7960
rect 39331 8000 39389 8001
rect 39331 7960 39340 8000
rect 39380 7960 39389 8000
rect 39331 7959 39389 7960
rect 39819 7986 39861 7995
rect 37851 7941 37893 7950
rect 39819 7946 39820 7986
rect 39860 7946 39861 7986
rect 39819 7937 39861 7946
rect 23107 7916 23165 7917
rect 21483 7867 21525 7876
rect 23107 7876 23116 7916
rect 23156 7876 23165 7916
rect 27387 7909 27429 7918
rect 31555 7916 31613 7917
rect 23107 7875 23165 7876
rect 31555 7876 31564 7916
rect 31604 7876 31613 7916
rect 31555 7875 31613 7876
rect 32419 7916 32477 7917
rect 32419 7876 32428 7916
rect 32468 7876 32477 7916
rect 32419 7875 32477 7876
rect 32803 7916 32861 7917
rect 32803 7876 32812 7916
rect 32852 7876 32861 7916
rect 32803 7875 32861 7876
rect 36747 7916 36789 7925
rect 36747 7876 36748 7916
rect 36788 7876 36789 7916
rect 36747 7867 36789 7876
rect 36843 7916 36885 7925
rect 36843 7876 36844 7916
rect 36884 7876 36885 7916
rect 36843 7867 36885 7876
rect 38763 7916 38805 7925
rect 38763 7876 38764 7916
rect 38804 7876 38805 7916
rect 38763 7867 38805 7876
rect 38859 7916 38901 7925
rect 38859 7876 38860 7916
rect 38900 7876 38901 7916
rect 38859 7867 38901 7876
rect 40483 7916 40541 7917
rect 40483 7876 40492 7916
rect 40532 7876 40541 7916
rect 40483 7875 40541 7876
rect 40867 7916 40925 7917
rect 40867 7876 40876 7916
rect 40916 7876 40925 7916
rect 40867 7875 40925 7876
rect 41251 7916 41309 7917
rect 41251 7876 41260 7916
rect 41300 7876 41309 7916
rect 41251 7875 41309 7876
rect 4963 7832 5021 7833
rect 4963 7792 4972 7832
rect 5012 7792 5021 7832
rect 4963 7791 5021 7792
rect 41067 7832 41109 7841
rect 41067 7792 41068 7832
rect 41108 7792 41109 7832
rect 41067 7783 41109 7792
rect 11211 7748 11253 7757
rect 11211 7708 11212 7748
rect 11252 7708 11253 7748
rect 11211 7699 11253 7708
rect 25515 7748 25557 7757
rect 25515 7708 25516 7748
rect 25556 7708 25557 7748
rect 25515 7699 25557 7708
rect 31371 7748 31413 7757
rect 31371 7708 31372 7748
rect 31412 7708 31413 7748
rect 31371 7699 31413 7708
rect 32619 7748 32661 7757
rect 32619 7708 32620 7748
rect 32660 7708 32661 7748
rect 32619 7699 32661 7708
rect 1152 7580 41856 7604
rect 1152 7540 3688 7580
rect 3728 7540 3770 7580
rect 3810 7540 3852 7580
rect 3892 7540 3934 7580
rect 3974 7540 4016 7580
rect 4056 7540 18808 7580
rect 18848 7540 18890 7580
rect 18930 7540 18972 7580
rect 19012 7540 19054 7580
rect 19094 7540 19136 7580
rect 19176 7540 33928 7580
rect 33968 7540 34010 7580
rect 34050 7540 34092 7580
rect 34132 7540 34174 7580
rect 34214 7540 34256 7580
rect 34296 7540 41856 7580
rect 1152 7516 41856 7540
rect 3627 7412 3669 7421
rect 3627 7372 3628 7412
rect 3668 7372 3669 7412
rect 3627 7363 3669 7372
rect 4395 7412 4437 7421
rect 4395 7372 4396 7412
rect 4436 7372 4437 7412
rect 4395 7363 4437 7372
rect 11691 7412 11733 7421
rect 11691 7372 11692 7412
rect 11732 7372 11733 7412
rect 11691 7363 11733 7372
rect 12939 7412 12981 7421
rect 12939 7372 12940 7412
rect 12980 7372 12981 7412
rect 12939 7363 12981 7372
rect 13707 7412 13749 7421
rect 13707 7372 13708 7412
rect 13748 7372 13749 7412
rect 13707 7363 13749 7372
rect 15819 7412 15861 7421
rect 15819 7372 15820 7412
rect 15860 7372 15861 7412
rect 15819 7363 15861 7372
rect 17451 7412 17493 7421
rect 17451 7372 17452 7412
rect 17492 7372 17493 7412
rect 17451 7363 17493 7372
rect 19083 7412 19125 7421
rect 19083 7372 19084 7412
rect 19124 7372 19125 7412
rect 19083 7363 19125 7372
rect 21099 7412 21141 7421
rect 21099 7372 21100 7412
rect 21140 7372 21141 7412
rect 21099 7363 21141 7372
rect 22827 7412 22869 7421
rect 22827 7372 22828 7412
rect 22868 7372 22869 7412
rect 22827 7363 22869 7372
rect 27531 7412 27573 7421
rect 27531 7372 27532 7412
rect 27572 7372 27573 7412
rect 27531 7363 27573 7372
rect 35979 7412 36021 7421
rect 35979 7372 35980 7412
rect 36020 7372 36021 7412
rect 35979 7363 36021 7372
rect 37707 7412 37749 7421
rect 37707 7372 37708 7412
rect 37748 7372 37749 7412
rect 37707 7363 37749 7372
rect 40395 7412 40437 7421
rect 40395 7372 40396 7412
rect 40436 7372 40437 7412
rect 40395 7363 40437 7372
rect 41451 7412 41493 7421
rect 41451 7372 41452 7412
rect 41492 7372 41493 7412
rect 41451 7363 41493 7372
rect 10251 7244 10293 7253
rect 10251 7204 10252 7244
rect 10292 7204 10293 7244
rect 11875 7244 11933 7245
rect 10251 7195 10293 7204
rect 11355 7202 11397 7211
rect 11875 7204 11884 7244
rect 11924 7204 11933 7244
rect 11875 7203 11933 7204
rect 12739 7244 12797 7245
rect 12739 7204 12748 7244
rect 12788 7204 12797 7244
rect 12739 7203 12797 7204
rect 13891 7244 13949 7245
rect 13891 7204 13900 7244
rect 13940 7204 13949 7244
rect 13891 7203 13949 7204
rect 33859 7244 33917 7245
rect 33859 7204 33868 7244
rect 33908 7204 33917 7244
rect 33859 7203 33917 7204
rect 40867 7244 40925 7245
rect 40867 7204 40876 7244
rect 40916 7204 40925 7244
rect 40867 7203 40925 7204
rect 41251 7244 41309 7245
rect 41251 7204 41260 7244
rect 41300 7204 41309 7244
rect 41251 7203 41309 7204
rect 1699 7160 1757 7161
rect 1699 7120 1708 7160
rect 1748 7120 1757 7160
rect 1699 7119 1757 7120
rect 2947 7160 3005 7161
rect 2947 7120 2956 7160
rect 2996 7120 3005 7160
rect 2947 7119 3005 7120
rect 3627 7160 3669 7169
rect 3627 7120 3628 7160
rect 3668 7120 3669 7160
rect 3627 7111 3669 7120
rect 3819 7160 3861 7169
rect 3819 7120 3820 7160
rect 3860 7120 3861 7160
rect 3819 7111 3861 7120
rect 3907 7160 3965 7161
rect 3907 7120 3916 7160
rect 3956 7120 3965 7160
rect 3907 7119 3965 7120
rect 4107 7160 4149 7169
rect 4107 7120 4108 7160
rect 4148 7120 4149 7160
rect 4107 7111 4149 7120
rect 4395 7160 4437 7169
rect 4395 7120 4396 7160
rect 4436 7120 4437 7160
rect 4395 7111 4437 7120
rect 4579 7160 4637 7161
rect 4579 7120 4588 7160
rect 4628 7120 4637 7160
rect 4579 7119 4637 7120
rect 5827 7160 5885 7161
rect 5827 7120 5836 7160
rect 5876 7120 5885 7160
rect 5827 7119 5885 7120
rect 6411 7160 6453 7169
rect 6411 7120 6412 7160
rect 6452 7120 6453 7160
rect 6411 7111 6453 7120
rect 6507 7160 6549 7169
rect 6507 7120 6508 7160
rect 6548 7120 6549 7160
rect 6507 7111 6549 7120
rect 8035 7160 8093 7161
rect 8035 7120 8044 7160
rect 8084 7120 8093 7160
rect 8035 7119 8093 7120
rect 9283 7160 9341 7161
rect 9283 7120 9292 7160
rect 9332 7120 9341 7160
rect 9283 7119 9341 7120
rect 9771 7160 9813 7169
rect 9771 7120 9772 7160
rect 9812 7120 9813 7160
rect 9771 7111 9813 7120
rect 9867 7160 9909 7169
rect 9867 7120 9868 7160
rect 9908 7120 9909 7160
rect 9867 7111 9909 7120
rect 10347 7160 10389 7169
rect 11355 7162 11356 7202
rect 11396 7162 11397 7202
rect 10347 7120 10348 7160
rect 10388 7120 10389 7160
rect 10347 7111 10389 7120
rect 10819 7160 10877 7161
rect 10819 7120 10828 7160
rect 10868 7120 10877 7160
rect 11355 7153 11397 7162
rect 14371 7160 14429 7161
rect 10819 7119 10877 7120
rect 14371 7120 14380 7160
rect 14420 7120 14429 7160
rect 14371 7119 14429 7120
rect 15619 7160 15677 7161
rect 15619 7120 15628 7160
rect 15668 7120 15677 7160
rect 15619 7119 15677 7120
rect 16003 7160 16061 7161
rect 16003 7120 16012 7160
rect 16052 7120 16061 7160
rect 16003 7119 16061 7120
rect 17251 7160 17309 7161
rect 17251 7120 17260 7160
rect 17300 7120 17309 7160
rect 17251 7119 17309 7120
rect 17635 7160 17693 7161
rect 17635 7120 17644 7160
rect 17684 7120 17693 7160
rect 17635 7119 17693 7120
rect 18883 7160 18941 7161
rect 18883 7120 18892 7160
rect 18932 7120 18941 7160
rect 18883 7119 18941 7120
rect 19651 7160 19709 7161
rect 19651 7120 19660 7160
rect 19700 7120 19709 7160
rect 19651 7119 19709 7120
rect 20899 7160 20957 7161
rect 20899 7120 20908 7160
rect 20948 7120 20957 7160
rect 20899 7119 20957 7120
rect 21379 7160 21437 7161
rect 21379 7120 21388 7160
rect 21428 7120 21437 7160
rect 21379 7119 21437 7120
rect 22627 7160 22685 7161
rect 22627 7120 22636 7160
rect 22676 7120 22685 7160
rect 22627 7119 22685 7120
rect 24355 7160 24413 7161
rect 24355 7120 24364 7160
rect 24404 7120 24413 7160
rect 24355 7119 24413 7120
rect 25603 7160 25661 7161
rect 25603 7120 25612 7160
rect 25652 7120 25661 7160
rect 25603 7119 25661 7120
rect 26083 7160 26141 7161
rect 26083 7120 26092 7160
rect 26132 7120 26141 7160
rect 26083 7119 26141 7120
rect 27331 7160 27389 7161
rect 27331 7120 27340 7160
rect 27380 7120 27389 7160
rect 27331 7119 27389 7120
rect 27715 7160 27773 7161
rect 27715 7120 27724 7160
rect 27764 7120 27773 7160
rect 27715 7119 27773 7120
rect 28963 7160 29021 7161
rect 28963 7120 28972 7160
rect 29012 7120 29021 7160
rect 28963 7119 29021 7120
rect 30211 7160 30269 7161
rect 30211 7120 30220 7160
rect 30260 7120 30269 7160
rect 30211 7119 30269 7120
rect 31459 7160 31517 7161
rect 31459 7120 31468 7160
rect 31508 7120 31517 7160
rect 31459 7119 31517 7120
rect 31939 7160 31997 7161
rect 31939 7120 31948 7160
rect 31988 7120 31997 7160
rect 31939 7119 31997 7120
rect 33187 7160 33245 7161
rect 33187 7120 33196 7160
rect 33236 7120 33245 7160
rect 33187 7119 33245 7120
rect 34531 7160 34589 7161
rect 34531 7120 34540 7160
rect 34580 7120 34589 7160
rect 34531 7119 34589 7120
rect 35779 7160 35837 7161
rect 35779 7120 35788 7160
rect 35828 7120 35837 7160
rect 35779 7119 35837 7120
rect 36259 7160 36317 7161
rect 36259 7120 36268 7160
rect 36308 7120 36317 7160
rect 36259 7119 36317 7120
rect 37507 7160 37565 7161
rect 37507 7120 37516 7160
rect 37556 7120 37565 7160
rect 37507 7119 37565 7120
rect 38947 7160 39005 7161
rect 38947 7120 38956 7160
rect 38996 7120 39005 7160
rect 38947 7119 39005 7120
rect 40195 7160 40253 7161
rect 40195 7120 40204 7160
rect 40244 7120 40253 7160
rect 40195 7119 40253 7120
rect 9483 7076 9525 7085
rect 9483 7036 9484 7076
rect 9524 7036 9525 7076
rect 9483 7027 9525 7036
rect 11499 7076 11541 7085
rect 11499 7036 11500 7076
rect 11540 7036 11541 7076
rect 11499 7027 11541 7036
rect 3147 6992 3189 7001
rect 3147 6952 3148 6992
rect 3188 6952 3189 6992
rect 3147 6943 3189 6952
rect 6027 6992 6069 7001
rect 6027 6952 6028 6992
rect 6068 6952 6069 6992
rect 6027 6943 6069 6952
rect 6211 6992 6269 6993
rect 6211 6952 6220 6992
rect 6260 6952 6269 6992
rect 6211 6951 6269 6952
rect 25803 6992 25845 7001
rect 25803 6952 25804 6992
rect 25844 6952 25845 6992
rect 25803 6943 25845 6952
rect 29163 6992 29205 7001
rect 29163 6952 29164 6992
rect 29204 6952 29205 6992
rect 29163 6943 29205 6952
rect 31659 6992 31701 7001
rect 31659 6952 31660 6992
rect 31700 6952 31701 6992
rect 31659 6943 31701 6952
rect 33387 6992 33429 7001
rect 33387 6952 33388 6992
rect 33428 6952 33429 6992
rect 33387 6943 33429 6952
rect 33675 6992 33717 7001
rect 33675 6952 33676 6992
rect 33716 6952 33717 6992
rect 33675 6943 33717 6952
rect 41067 6992 41109 7001
rect 41067 6952 41068 6992
rect 41108 6952 41109 6992
rect 41067 6943 41109 6952
rect 1152 6824 41856 6848
rect 1152 6784 4928 6824
rect 4968 6784 5010 6824
rect 5050 6784 5092 6824
rect 5132 6784 5174 6824
rect 5214 6784 5256 6824
rect 5296 6784 20048 6824
rect 20088 6784 20130 6824
rect 20170 6784 20212 6824
rect 20252 6784 20294 6824
rect 20334 6784 20376 6824
rect 20416 6784 35168 6824
rect 35208 6784 35250 6824
rect 35290 6784 35332 6824
rect 35372 6784 35414 6824
rect 35454 6784 35496 6824
rect 35536 6784 41856 6824
rect 1152 6760 41856 6784
rect 7267 6656 7325 6657
rect 7267 6616 7276 6656
rect 7316 6616 7325 6656
rect 7267 6615 7325 6616
rect 10347 6656 10389 6665
rect 10347 6616 10348 6656
rect 10388 6616 10389 6656
rect 10347 6607 10389 6616
rect 14187 6656 14229 6665
rect 14187 6616 14188 6656
rect 14228 6616 14229 6656
rect 14187 6607 14229 6616
rect 14667 6656 14709 6665
rect 14667 6616 14668 6656
rect 14708 6616 14709 6656
rect 14667 6607 14709 6616
rect 19467 6656 19509 6665
rect 19467 6616 19468 6656
rect 19508 6616 19509 6656
rect 19467 6607 19509 6616
rect 21291 6656 21333 6665
rect 21291 6616 21292 6656
rect 21332 6616 21333 6656
rect 21291 6607 21333 6616
rect 23307 6656 23349 6665
rect 23307 6616 23308 6656
rect 23348 6616 23349 6656
rect 23307 6607 23349 6616
rect 25707 6656 25749 6665
rect 25707 6616 25708 6656
rect 25748 6616 25749 6656
rect 25707 6607 25749 6616
rect 30891 6656 30933 6665
rect 30891 6616 30892 6656
rect 30932 6616 30933 6656
rect 30891 6607 30933 6616
rect 33195 6656 33237 6665
rect 33195 6616 33196 6656
rect 33236 6616 33237 6656
rect 33195 6607 33237 6616
rect 37611 6656 37653 6665
rect 37611 6616 37612 6656
rect 37652 6616 37653 6656
rect 37611 6607 37653 6616
rect 41451 6656 41493 6665
rect 41451 6616 41452 6656
rect 41492 6616 41493 6656
rect 41451 6607 41493 6616
rect 4491 6572 4533 6581
rect 4491 6532 4492 6572
rect 4532 6532 4533 6572
rect 4491 6523 4533 6532
rect 8907 6572 8949 6581
rect 8907 6532 8908 6572
rect 8948 6532 8949 6572
rect 8907 6523 8949 6532
rect 12171 6572 12213 6581
rect 12171 6532 12172 6572
rect 12212 6532 12213 6572
rect 12171 6523 12213 6532
rect 28875 6572 28917 6581
rect 28875 6532 28876 6572
rect 28916 6532 28917 6572
rect 28875 6523 28917 6532
rect 40011 6572 40053 6581
rect 40011 6532 40012 6572
rect 40052 6532 40053 6572
rect 40011 6523 40053 6532
rect 2755 6488 2813 6489
rect 2755 6448 2764 6488
rect 2804 6448 2813 6488
rect 2755 6447 2813 6448
rect 4003 6488 4061 6489
rect 4003 6448 4012 6488
rect 4052 6448 4061 6488
rect 5155 6488 5213 6489
rect 4003 6447 4061 6448
rect 4683 6474 4725 6483
rect 4683 6434 4684 6474
rect 4724 6434 4725 6474
rect 5155 6448 5164 6488
rect 5204 6448 5213 6488
rect 5155 6447 5213 6448
rect 6123 6488 6165 6497
rect 6123 6448 6124 6488
rect 6164 6448 6165 6488
rect 6123 6439 6165 6448
rect 6219 6488 6261 6497
rect 6219 6448 6220 6488
rect 6260 6448 6261 6488
rect 6219 6439 6261 6448
rect 6507 6488 6549 6497
rect 6507 6448 6508 6488
rect 6548 6448 6549 6488
rect 6507 6439 6549 6448
rect 6603 6488 6645 6497
rect 6603 6448 6604 6488
rect 6644 6448 6645 6488
rect 6603 6439 6645 6448
rect 6699 6488 6741 6497
rect 6699 6448 6700 6488
rect 6740 6448 6741 6488
rect 6699 6439 6741 6448
rect 6795 6488 6837 6497
rect 6795 6448 6796 6488
rect 6836 6448 6837 6488
rect 6795 6439 6837 6448
rect 6987 6488 7029 6497
rect 6987 6448 6988 6488
rect 7028 6448 7029 6488
rect 6987 6439 7029 6448
rect 7083 6488 7125 6497
rect 7083 6448 7084 6488
rect 7124 6448 7125 6488
rect 7083 6439 7125 6448
rect 7179 6488 7221 6497
rect 7179 6448 7180 6488
rect 7220 6448 7221 6488
rect 7179 6439 7221 6448
rect 7459 6488 7517 6489
rect 7459 6448 7468 6488
rect 7508 6448 7517 6488
rect 7459 6447 7517 6448
rect 8707 6488 8765 6489
rect 8707 6448 8716 6488
rect 8756 6448 8765 6488
rect 8707 6447 8765 6448
rect 9187 6488 9245 6489
rect 9187 6448 9196 6488
rect 9236 6448 9245 6488
rect 9187 6447 9245 6448
rect 9483 6488 9525 6497
rect 9483 6448 9484 6488
rect 9524 6448 9525 6488
rect 9483 6439 9525 6448
rect 9579 6488 9621 6497
rect 9579 6448 9580 6488
rect 9620 6448 9621 6488
rect 9579 6439 9621 6448
rect 10723 6488 10781 6489
rect 10723 6448 10732 6488
rect 10772 6448 10781 6488
rect 10723 6447 10781 6448
rect 11971 6488 12029 6489
rect 11971 6448 11980 6488
rect 12020 6448 12029 6488
rect 11971 6447 12029 6448
rect 12459 6488 12501 6497
rect 12459 6448 12460 6488
rect 12500 6448 12501 6488
rect 12459 6439 12501 6448
rect 12555 6488 12597 6497
rect 12555 6448 12556 6488
rect 12596 6448 12597 6488
rect 12555 6439 12597 6448
rect 12939 6488 12981 6497
rect 12939 6448 12940 6488
rect 12980 6448 12981 6488
rect 12939 6439 12981 6448
rect 13507 6488 13565 6489
rect 13507 6448 13516 6488
rect 13556 6448 13565 6488
rect 15331 6488 15389 6489
rect 13507 6447 13565 6448
rect 13995 6474 14037 6483
rect 4683 6425 4725 6434
rect 13995 6434 13996 6474
rect 14036 6434 14037 6474
rect 13995 6425 14037 6434
rect 14811 6446 14853 6455
rect 15331 6448 15340 6488
rect 15380 6448 15389 6488
rect 15331 6447 15389 6448
rect 15915 6488 15957 6497
rect 15915 6448 15916 6488
rect 15956 6448 15957 6488
rect 5643 6404 5685 6413
rect 5643 6364 5644 6404
rect 5684 6364 5685 6404
rect 5643 6355 5685 6364
rect 5739 6404 5781 6413
rect 5739 6364 5740 6404
rect 5780 6364 5781 6404
rect 5739 6355 5781 6364
rect 10531 6404 10589 6405
rect 10531 6364 10540 6404
rect 10580 6364 10589 6404
rect 10531 6363 10589 6364
rect 13035 6404 13077 6413
rect 13035 6364 13036 6404
rect 13076 6364 13077 6404
rect 14811 6406 14812 6446
rect 14852 6406 14853 6446
rect 15915 6439 15957 6448
rect 16299 6488 16341 6497
rect 16299 6448 16300 6488
rect 16340 6448 16341 6488
rect 16299 6439 16341 6448
rect 16395 6488 16437 6497
rect 16395 6448 16396 6488
rect 16436 6448 16437 6488
rect 16395 6439 16437 6448
rect 17635 6488 17693 6489
rect 17635 6448 17644 6488
rect 17684 6448 17693 6488
rect 17635 6447 17693 6448
rect 18883 6488 18941 6489
rect 18883 6448 18892 6488
rect 18932 6448 18941 6488
rect 18883 6447 18941 6448
rect 19843 6488 19901 6489
rect 19843 6448 19852 6488
rect 19892 6448 19901 6488
rect 19843 6447 19901 6448
rect 21091 6488 21149 6489
rect 21091 6448 21100 6488
rect 21140 6448 21149 6488
rect 21091 6447 21149 6448
rect 21579 6488 21621 6497
rect 21579 6448 21580 6488
rect 21620 6448 21621 6488
rect 21579 6439 21621 6448
rect 21675 6488 21717 6497
rect 21675 6448 21676 6488
rect 21716 6448 21717 6488
rect 21675 6439 21717 6448
rect 22059 6488 22101 6497
rect 22059 6448 22060 6488
rect 22100 6448 22101 6488
rect 22059 6439 22101 6448
rect 22155 6488 22197 6497
rect 22155 6448 22156 6488
rect 22196 6448 22197 6488
rect 22155 6439 22197 6448
rect 22627 6488 22685 6489
rect 22627 6448 22636 6488
rect 22676 6448 22685 6488
rect 23979 6488 24021 6497
rect 22627 6447 22685 6448
rect 23115 6474 23157 6483
rect 23115 6434 23116 6474
rect 23156 6434 23157 6474
rect 23979 6448 23980 6488
rect 24020 6448 24021 6488
rect 23979 6439 24021 6448
rect 24075 6488 24117 6497
rect 24075 6448 24076 6488
rect 24116 6448 24117 6488
rect 24075 6439 24117 6448
rect 24459 6488 24501 6497
rect 24459 6448 24460 6488
rect 24500 6448 24501 6488
rect 24459 6439 24501 6448
rect 24555 6488 24597 6497
rect 24555 6448 24556 6488
rect 24596 6448 24597 6488
rect 24555 6439 24597 6448
rect 25027 6488 25085 6489
rect 25027 6448 25036 6488
rect 25076 6448 25085 6488
rect 25027 6447 25085 6448
rect 25515 6483 25557 6492
rect 25515 6443 25516 6483
rect 25556 6443 25557 6483
rect 25515 6434 25557 6443
rect 27147 6488 27189 6497
rect 27147 6448 27148 6488
rect 27188 6448 27189 6488
rect 27147 6439 27189 6448
rect 27243 6488 27285 6497
rect 27243 6448 27244 6488
rect 27284 6448 27285 6488
rect 27243 6439 27285 6448
rect 27627 6488 27669 6497
rect 27627 6448 27628 6488
rect 27668 6448 27669 6488
rect 27627 6439 27669 6448
rect 27723 6488 27765 6497
rect 27723 6448 27724 6488
rect 27764 6448 27765 6488
rect 27723 6439 27765 6448
rect 28195 6488 28253 6489
rect 28195 6448 28204 6488
rect 28244 6448 28253 6488
rect 28195 6447 28253 6448
rect 28683 6483 28725 6492
rect 28683 6443 28684 6483
rect 28724 6443 28725 6483
rect 28683 6434 28725 6443
rect 29163 6488 29205 6497
rect 29163 6448 29164 6488
rect 29204 6448 29205 6488
rect 29163 6439 29205 6448
rect 29259 6488 29301 6497
rect 29259 6448 29260 6488
rect 29300 6448 29301 6488
rect 29259 6439 29301 6448
rect 29643 6488 29685 6497
rect 29643 6448 29644 6488
rect 29684 6448 29685 6488
rect 29643 6439 29685 6448
rect 29739 6488 29781 6497
rect 29739 6448 29740 6488
rect 29780 6448 29781 6488
rect 29739 6439 29781 6448
rect 30211 6488 30269 6489
rect 30211 6448 30220 6488
rect 30260 6448 30269 6488
rect 31467 6488 31509 6497
rect 30211 6447 30269 6448
rect 30699 6474 30741 6483
rect 30699 6434 30700 6474
rect 30740 6434 30741 6474
rect 31467 6448 31468 6488
rect 31508 6448 31509 6488
rect 31467 6439 31509 6448
rect 31563 6488 31605 6497
rect 31563 6448 31564 6488
rect 31604 6448 31605 6488
rect 31563 6439 31605 6448
rect 31947 6488 31989 6497
rect 31947 6448 31948 6488
rect 31988 6448 31989 6488
rect 31947 6439 31989 6448
rect 32515 6488 32573 6489
rect 32515 6448 32524 6488
rect 32564 6448 32573 6488
rect 33379 6488 33437 6489
rect 32515 6447 32573 6448
rect 33051 6446 33093 6455
rect 33379 6448 33388 6488
rect 33428 6448 33437 6488
rect 33379 6447 33437 6448
rect 34627 6488 34685 6489
rect 34627 6448 34636 6488
rect 34676 6448 34685 6488
rect 34627 6447 34685 6448
rect 38283 6488 38325 6497
rect 38283 6448 38284 6488
rect 38324 6448 38325 6488
rect 23115 6425 23157 6434
rect 30699 6425 30741 6434
rect 14811 6397 14853 6406
rect 15819 6404 15861 6413
rect 13035 6355 13077 6364
rect 15819 6364 15820 6404
rect 15860 6364 15861 6404
rect 15819 6355 15861 6364
rect 19651 6404 19709 6405
rect 19651 6364 19660 6404
rect 19700 6364 19709 6404
rect 19651 6363 19709 6364
rect 32043 6404 32085 6413
rect 32043 6364 32044 6404
rect 32084 6364 32085 6404
rect 33051 6406 33052 6446
rect 33092 6406 33093 6446
rect 38283 6439 38325 6448
rect 38379 6488 38421 6497
rect 38379 6448 38380 6488
rect 38420 6448 38421 6488
rect 38379 6439 38421 6448
rect 38763 6488 38805 6497
rect 38763 6448 38764 6488
rect 38804 6448 38805 6488
rect 38763 6439 38805 6448
rect 38859 6488 38901 6497
rect 38859 6448 38860 6488
rect 38900 6448 38901 6488
rect 38859 6439 38901 6448
rect 39331 6488 39389 6489
rect 39331 6448 39340 6488
rect 39380 6448 39389 6488
rect 39331 6447 39389 6448
rect 39819 6474 39861 6483
rect 39819 6434 39820 6474
rect 39860 6434 39861 6474
rect 39819 6425 39861 6434
rect 33051 6397 33093 6406
rect 35875 6404 35933 6405
rect 32043 6355 32085 6364
rect 35875 6364 35884 6404
rect 35924 6364 35933 6404
rect 35875 6363 35933 6364
rect 37795 6404 37853 6405
rect 37795 6364 37804 6404
rect 37844 6364 37853 6404
rect 37795 6363 37853 6364
rect 40387 6404 40445 6405
rect 40387 6364 40396 6404
rect 40436 6364 40445 6404
rect 40387 6363 40445 6364
rect 40867 6404 40925 6405
rect 40867 6364 40876 6404
rect 40916 6364 40925 6404
rect 40867 6363 40925 6364
rect 41251 6404 41309 6405
rect 41251 6364 41260 6404
rect 41300 6364 41309 6404
rect 41251 6363 41309 6364
rect 4203 6320 4245 6329
rect 4203 6280 4204 6320
rect 4244 6280 4245 6320
rect 4203 6271 4245 6280
rect 9859 6320 9917 6321
rect 9859 6280 9868 6320
rect 9908 6280 9917 6320
rect 9859 6279 9917 6280
rect 19083 6320 19125 6329
rect 19083 6280 19084 6320
rect 19124 6280 19125 6320
rect 19083 6271 19125 6280
rect 35691 6320 35733 6329
rect 35691 6280 35692 6320
rect 35732 6280 35733 6320
rect 35691 6271 35733 6280
rect 40203 6320 40245 6329
rect 40203 6280 40204 6320
rect 40244 6280 40245 6320
rect 40203 6271 40245 6280
rect 41067 6320 41109 6329
rect 41067 6280 41068 6320
rect 41108 6280 41109 6320
rect 41067 6271 41109 6280
rect 34827 6236 34869 6245
rect 34827 6196 34828 6236
rect 34868 6196 34869 6236
rect 34827 6187 34869 6196
rect 1152 6068 41856 6092
rect 1152 6028 3688 6068
rect 3728 6028 3770 6068
rect 3810 6028 3852 6068
rect 3892 6028 3934 6068
rect 3974 6028 4016 6068
rect 4056 6028 18808 6068
rect 18848 6028 18890 6068
rect 18930 6028 18972 6068
rect 19012 6028 19054 6068
rect 19094 6028 19136 6068
rect 19176 6028 33928 6068
rect 33968 6028 34010 6068
rect 34050 6028 34092 6068
rect 34132 6028 34174 6068
rect 34214 6028 34256 6068
rect 34296 6028 41856 6068
rect 1152 6004 41856 6028
rect 4683 5900 4725 5909
rect 4683 5860 4684 5900
rect 4724 5860 4725 5900
rect 4683 5851 4725 5860
rect 10923 5900 10965 5909
rect 10923 5860 10924 5900
rect 10964 5860 10965 5900
rect 10923 5851 10965 5860
rect 12843 5900 12885 5909
rect 12843 5860 12844 5900
rect 12884 5860 12885 5900
rect 12843 5851 12885 5860
rect 14475 5900 14517 5909
rect 14475 5860 14476 5900
rect 14516 5860 14517 5900
rect 14475 5851 14517 5860
rect 14667 5900 14709 5909
rect 14667 5860 14668 5900
rect 14708 5860 14709 5900
rect 14667 5851 14709 5860
rect 22731 5900 22773 5909
rect 22731 5860 22732 5900
rect 22772 5860 22773 5900
rect 22731 5851 22773 5860
rect 27243 5900 27285 5909
rect 27243 5860 27244 5900
rect 27284 5860 27285 5900
rect 27243 5851 27285 5860
rect 40395 5900 40437 5909
rect 40395 5860 40396 5900
rect 40436 5860 40437 5900
rect 40395 5851 40437 5860
rect 41067 5900 41109 5909
rect 41067 5860 41068 5900
rect 41108 5860 41109 5900
rect 41067 5851 41109 5860
rect 4299 5816 4341 5825
rect 4299 5776 4300 5816
rect 4340 5776 4341 5816
rect 4299 5767 4341 5776
rect 19939 5816 19997 5817
rect 19939 5776 19948 5816
rect 19988 5776 19997 5816
rect 19939 5775 19997 5776
rect 24363 5816 24405 5825
rect 24363 5776 24364 5816
rect 24404 5776 24405 5816
rect 24363 5767 24405 5776
rect 41451 5816 41493 5825
rect 41451 5776 41452 5816
rect 41492 5776 41493 5816
rect 41451 5767 41493 5776
rect 11107 5732 11165 5733
rect 11107 5692 11116 5732
rect 11156 5692 11165 5732
rect 11107 5691 11165 5692
rect 12643 5732 12701 5733
rect 12643 5692 12652 5732
rect 12692 5692 12701 5732
rect 12643 5691 12701 5692
rect 28483 5732 28541 5733
rect 28483 5692 28492 5732
rect 28532 5692 28541 5732
rect 28483 5691 28541 5692
rect 29355 5732 29397 5741
rect 29355 5692 29356 5732
rect 29396 5692 29397 5732
rect 29355 5683 29397 5692
rect 29451 5732 29493 5741
rect 29451 5692 29452 5732
rect 29492 5692 29493 5732
rect 29451 5683 29493 5692
rect 32043 5732 32085 5741
rect 32043 5692 32044 5732
rect 32084 5692 32085 5732
rect 32043 5683 32085 5692
rect 32139 5732 32181 5741
rect 32139 5692 32140 5732
rect 32180 5692 32181 5732
rect 32139 5683 32181 5692
rect 34827 5732 34869 5741
rect 34827 5692 34828 5732
rect 34868 5692 34869 5732
rect 34827 5683 34869 5692
rect 36843 5732 36885 5741
rect 36843 5692 36844 5732
rect 36884 5692 36885 5732
rect 36843 5683 36885 5692
rect 40867 5732 40925 5733
rect 40867 5692 40876 5732
rect 40916 5692 40925 5732
rect 40867 5691 40925 5692
rect 41251 5732 41309 5733
rect 41251 5692 41260 5732
rect 41300 5692 41309 5732
rect 41251 5691 41309 5692
rect 7323 5657 7365 5666
rect 1603 5648 1661 5649
rect 1603 5608 1612 5648
rect 1652 5608 1661 5648
rect 1603 5607 1661 5608
rect 2851 5648 2909 5649
rect 2851 5608 2860 5648
rect 2900 5608 2909 5648
rect 2851 5607 2909 5608
rect 4299 5648 4341 5657
rect 4299 5608 4300 5648
rect 4340 5608 4341 5648
rect 4299 5599 4341 5608
rect 4771 5648 4829 5649
rect 4771 5608 4780 5648
rect 4820 5608 4829 5648
rect 4771 5607 4829 5608
rect 5163 5648 5205 5657
rect 5163 5608 5164 5648
rect 5204 5608 5205 5648
rect 5163 5599 5205 5608
rect 5259 5648 5301 5657
rect 5259 5608 5260 5648
rect 5300 5608 5301 5648
rect 5259 5599 5301 5608
rect 5739 5648 5781 5657
rect 5739 5608 5740 5648
rect 5780 5608 5781 5648
rect 5739 5599 5781 5608
rect 5835 5648 5877 5657
rect 5835 5608 5836 5648
rect 5876 5608 5877 5648
rect 5835 5599 5877 5608
rect 6219 5648 6261 5657
rect 6219 5608 6220 5648
rect 6260 5608 6261 5648
rect 6219 5599 6261 5608
rect 6315 5648 6357 5657
rect 6315 5608 6316 5648
rect 6356 5608 6357 5648
rect 6315 5599 6357 5608
rect 6787 5648 6845 5649
rect 6787 5608 6796 5648
rect 6836 5608 6845 5648
rect 7323 5617 7324 5657
rect 7364 5617 7365 5657
rect 7323 5608 7365 5617
rect 7651 5648 7709 5649
rect 7651 5608 7660 5648
rect 7700 5608 7709 5648
rect 6787 5607 6845 5608
rect 7651 5607 7709 5608
rect 8899 5648 8957 5649
rect 8899 5608 8908 5648
rect 8948 5608 8957 5648
rect 8899 5607 8957 5608
rect 9283 5648 9341 5649
rect 9283 5608 9292 5648
rect 9332 5608 9341 5648
rect 9283 5607 9341 5608
rect 10531 5648 10589 5649
rect 10531 5608 10540 5648
rect 10580 5608 10589 5648
rect 10531 5607 10589 5608
rect 13027 5648 13085 5649
rect 13027 5608 13036 5648
rect 13076 5608 13085 5648
rect 13027 5607 13085 5608
rect 14275 5648 14333 5649
rect 14275 5608 14284 5648
rect 14324 5608 14333 5648
rect 14275 5607 14333 5608
rect 14851 5648 14909 5649
rect 14851 5608 14860 5648
rect 14900 5608 14909 5648
rect 14851 5607 14909 5608
rect 16099 5648 16157 5649
rect 16099 5608 16108 5648
rect 16148 5608 16157 5648
rect 16099 5607 16157 5608
rect 16291 5648 16349 5649
rect 16291 5608 16300 5648
rect 16340 5608 16349 5648
rect 16291 5607 16349 5608
rect 17539 5648 17597 5649
rect 17539 5608 17548 5648
rect 17588 5608 17597 5648
rect 17539 5607 17597 5608
rect 18027 5648 18069 5657
rect 18027 5608 18028 5648
rect 18068 5608 18069 5648
rect 18027 5599 18069 5608
rect 18123 5648 18165 5657
rect 18123 5608 18124 5648
rect 18164 5608 18165 5648
rect 18123 5599 18165 5608
rect 18507 5648 18549 5657
rect 18507 5608 18508 5648
rect 18548 5608 18549 5648
rect 18507 5599 18549 5608
rect 18603 5648 18645 5657
rect 19563 5653 19605 5662
rect 30459 5657 30501 5666
rect 33147 5657 33189 5666
rect 18603 5608 18604 5648
rect 18644 5608 18645 5648
rect 18603 5599 18645 5608
rect 19075 5648 19133 5649
rect 19075 5608 19084 5648
rect 19124 5608 19133 5648
rect 19075 5607 19133 5608
rect 19563 5613 19564 5653
rect 19604 5613 19605 5653
rect 19563 5604 19605 5613
rect 20331 5648 20373 5657
rect 20331 5608 20332 5648
rect 20372 5608 20373 5648
rect 20331 5599 20373 5608
rect 20611 5648 20669 5649
rect 20611 5608 20620 5648
rect 20660 5608 20669 5648
rect 20611 5607 20669 5608
rect 21283 5648 21341 5649
rect 21283 5608 21292 5648
rect 21332 5608 21341 5648
rect 21283 5607 21341 5608
rect 22531 5648 22589 5649
rect 22531 5608 22540 5648
rect 22580 5608 22589 5648
rect 22531 5607 22589 5608
rect 22915 5648 22973 5649
rect 22915 5608 22924 5648
rect 22964 5608 22973 5648
rect 22915 5607 22973 5608
rect 24163 5648 24221 5649
rect 24163 5608 24172 5648
rect 24212 5608 24221 5648
rect 24163 5607 24221 5608
rect 25795 5648 25853 5649
rect 25795 5608 25804 5648
rect 25844 5608 25853 5648
rect 25795 5607 25853 5608
rect 27043 5648 27101 5649
rect 27043 5608 27052 5648
rect 27092 5608 27101 5648
rect 27043 5607 27101 5608
rect 28875 5648 28917 5657
rect 28875 5608 28876 5648
rect 28916 5608 28917 5648
rect 28875 5599 28917 5608
rect 28971 5648 29013 5657
rect 28971 5608 28972 5648
rect 29012 5608 29013 5648
rect 28971 5599 29013 5608
rect 29923 5639 29981 5640
rect 29923 5599 29932 5639
rect 29972 5599 29981 5639
rect 30459 5617 30460 5657
rect 30500 5617 30501 5657
rect 30459 5608 30501 5617
rect 31563 5648 31605 5657
rect 31563 5608 31564 5648
rect 31604 5608 31605 5648
rect 31563 5599 31605 5608
rect 31659 5648 31701 5657
rect 31659 5608 31660 5648
rect 31700 5608 31701 5648
rect 31659 5599 31701 5608
rect 32611 5648 32669 5649
rect 32611 5608 32620 5648
rect 32660 5608 32669 5648
rect 33147 5617 33148 5657
rect 33188 5617 33189 5657
rect 33147 5608 33189 5617
rect 34347 5648 34389 5657
rect 34347 5608 34348 5648
rect 34388 5608 34389 5648
rect 32611 5607 32669 5608
rect 34347 5599 34389 5608
rect 34443 5648 34485 5657
rect 34443 5608 34444 5648
rect 34484 5608 34485 5648
rect 34443 5599 34485 5608
rect 34923 5648 34965 5657
rect 35883 5653 35925 5662
rect 34923 5608 34924 5648
rect 34964 5608 34965 5648
rect 34923 5599 34965 5608
rect 35395 5648 35453 5649
rect 35395 5608 35404 5648
rect 35444 5608 35453 5648
rect 35395 5607 35453 5608
rect 35883 5613 35884 5653
rect 35924 5613 35925 5653
rect 35883 5604 35925 5613
rect 36363 5648 36405 5657
rect 36363 5608 36364 5648
rect 36404 5608 36405 5648
rect 36363 5599 36405 5608
rect 36459 5648 36501 5657
rect 36459 5608 36460 5648
rect 36500 5608 36501 5648
rect 36459 5599 36501 5608
rect 36939 5648 36981 5657
rect 37899 5653 37941 5662
rect 36939 5608 36940 5648
rect 36980 5608 36981 5648
rect 36939 5599 36981 5608
rect 37411 5648 37469 5649
rect 37411 5608 37420 5648
rect 37460 5608 37469 5648
rect 37411 5607 37469 5608
rect 37899 5613 37900 5653
rect 37940 5613 37941 5653
rect 37899 5604 37941 5613
rect 38947 5648 39005 5649
rect 38947 5608 38956 5648
rect 38996 5608 39005 5648
rect 38947 5607 39005 5608
rect 40195 5648 40253 5649
rect 40195 5608 40204 5648
rect 40244 5608 40253 5648
rect 40195 5607 40253 5608
rect 29923 5598 29981 5599
rect 17739 5564 17781 5573
rect 17739 5524 17740 5564
rect 17780 5524 17781 5564
rect 17739 5515 17781 5524
rect 19755 5564 19797 5573
rect 19755 5524 19756 5564
rect 19796 5524 19797 5564
rect 19755 5515 19797 5524
rect 20235 5564 20277 5573
rect 20235 5524 20236 5564
rect 20276 5524 20277 5564
rect 20235 5515 20277 5524
rect 30603 5564 30645 5573
rect 30603 5524 30604 5564
rect 30644 5524 30645 5564
rect 30603 5515 30645 5524
rect 36075 5564 36117 5573
rect 36075 5524 36076 5564
rect 36116 5524 36117 5564
rect 36075 5515 36117 5524
rect 38091 5564 38133 5573
rect 38091 5524 38092 5564
rect 38132 5524 38133 5564
rect 38091 5515 38133 5524
rect 3051 5480 3093 5489
rect 3051 5440 3052 5480
rect 3092 5440 3093 5480
rect 3051 5431 3093 5440
rect 4491 5480 4533 5489
rect 4491 5440 4492 5480
rect 4532 5440 4533 5480
rect 4491 5431 4533 5440
rect 5443 5480 5501 5481
rect 5443 5440 5452 5480
rect 5492 5440 5501 5480
rect 5443 5439 5501 5440
rect 7467 5480 7509 5489
rect 7467 5440 7468 5480
rect 7508 5440 7509 5480
rect 7467 5431 7509 5440
rect 9099 5480 9141 5489
rect 9099 5440 9100 5480
rect 9140 5440 9141 5480
rect 9099 5431 9141 5440
rect 10731 5480 10773 5489
rect 10731 5440 10732 5480
rect 10772 5440 10773 5480
rect 10731 5431 10773 5440
rect 28299 5480 28341 5489
rect 28299 5440 28300 5480
rect 28340 5440 28341 5480
rect 28299 5431 28341 5440
rect 33291 5480 33333 5489
rect 33291 5440 33292 5480
rect 33332 5440 33333 5480
rect 33291 5431 33333 5440
rect 1152 5312 41856 5336
rect 1152 5272 4928 5312
rect 4968 5272 5010 5312
rect 5050 5272 5092 5312
rect 5132 5272 5174 5312
rect 5214 5272 5256 5312
rect 5296 5272 20048 5312
rect 20088 5272 20130 5312
rect 20170 5272 20212 5312
rect 20252 5272 20294 5312
rect 20334 5272 20376 5312
rect 20416 5272 35168 5312
rect 35208 5272 35250 5312
rect 35290 5272 35332 5312
rect 35372 5272 35414 5312
rect 35454 5272 35496 5312
rect 35536 5272 41856 5312
rect 1152 5248 41856 5272
rect 3907 5144 3965 5145
rect 3907 5104 3916 5144
rect 3956 5104 3965 5144
rect 3907 5103 3965 5104
rect 11211 5144 11253 5153
rect 11211 5104 11212 5144
rect 11252 5104 11253 5144
rect 11211 5095 11253 5104
rect 19755 5144 19797 5153
rect 19755 5104 19756 5144
rect 19796 5104 19797 5144
rect 19755 5095 19797 5104
rect 28875 5144 28917 5153
rect 28875 5104 28876 5144
rect 28916 5104 28917 5144
rect 28875 5095 28917 5104
rect 33483 5144 33525 5153
rect 33483 5104 33484 5144
rect 33524 5104 33525 5144
rect 33483 5095 33525 5104
rect 35787 5144 35829 5153
rect 35787 5104 35788 5144
rect 35828 5104 35829 5144
rect 35787 5095 35829 5104
rect 5163 5060 5205 5069
rect 5163 5020 5164 5060
rect 5204 5020 5205 5060
rect 5163 5011 5205 5020
rect 5739 5060 5781 5069
rect 5739 5020 5740 5060
rect 5780 5020 5781 5060
rect 5739 5011 5781 5020
rect 7755 5060 7797 5069
rect 7755 5020 7756 5060
rect 7796 5020 7797 5060
rect 7755 5011 7797 5020
rect 13899 5060 13941 5069
rect 13899 5020 13900 5060
rect 13940 5020 13941 5060
rect 13899 5011 13941 5020
rect 23115 5060 23157 5069
rect 23115 5020 23116 5060
rect 23156 5020 23157 5060
rect 23115 5011 23157 5020
rect 30891 5060 30933 5069
rect 30891 5020 30892 5060
rect 30932 5020 30933 5060
rect 30891 5011 30933 5020
rect 38667 5060 38709 5069
rect 38667 5020 38668 5060
rect 38708 5020 38709 5060
rect 38667 5011 38709 5020
rect 1699 4976 1757 4977
rect 1699 4936 1708 4976
rect 1748 4936 1757 4976
rect 1699 4935 1757 4936
rect 2947 4976 3005 4977
rect 2947 4936 2956 4976
rect 2996 4936 3005 4976
rect 2947 4935 3005 4936
rect 3627 4976 3669 4985
rect 3627 4936 3628 4976
rect 3668 4936 3669 4976
rect 3627 4927 3669 4936
rect 3723 4976 3765 4985
rect 3723 4936 3724 4976
rect 3764 4936 3765 4976
rect 3723 4927 3765 4936
rect 4107 4976 4149 4985
rect 4107 4936 4108 4976
rect 4148 4936 4149 4976
rect 4107 4927 4149 4936
rect 4299 4976 4341 4985
rect 4299 4936 4300 4976
rect 4340 4936 4341 4976
rect 4299 4927 4341 4936
rect 4387 4976 4445 4977
rect 4387 4936 4396 4976
rect 4436 4936 4445 4976
rect 4387 4935 4445 4936
rect 4587 4976 4629 4985
rect 4587 4936 4588 4976
rect 4628 4936 4629 4976
rect 4587 4927 4629 4936
rect 4875 4976 4917 4985
rect 4875 4936 4876 4976
rect 4916 4936 4917 4976
rect 4875 4927 4917 4936
rect 5067 4976 5109 4985
rect 5067 4936 5068 4976
rect 5108 4936 5109 4976
rect 5067 4927 5109 4936
rect 5251 4976 5309 4977
rect 5251 4936 5260 4976
rect 5300 4936 5309 4976
rect 5251 4935 5309 4936
rect 5451 4976 5493 4985
rect 5451 4936 5452 4976
rect 5492 4936 5493 4976
rect 5451 4927 5493 4936
rect 5547 4976 5589 4985
rect 5547 4936 5548 4976
rect 5588 4936 5589 4976
rect 5547 4927 5589 4936
rect 5643 4976 5685 4985
rect 5643 4936 5644 4976
rect 5684 4936 5685 4976
rect 5643 4927 5685 4936
rect 6027 4976 6069 4985
rect 6027 4936 6028 4976
rect 6068 4936 6069 4976
rect 6027 4927 6069 4936
rect 6123 4976 6165 4985
rect 6123 4936 6124 4976
rect 6164 4936 6165 4976
rect 6123 4927 6165 4936
rect 6507 4976 6549 4985
rect 6507 4936 6508 4976
rect 6548 4936 6549 4976
rect 6507 4927 6549 4936
rect 6603 4976 6645 4985
rect 6603 4936 6604 4976
rect 6644 4936 6645 4976
rect 6603 4927 6645 4936
rect 7075 4976 7133 4977
rect 7075 4936 7084 4976
rect 7124 4936 7133 4976
rect 9483 4976 9525 4985
rect 7075 4935 7133 4936
rect 7563 4962 7605 4971
rect 7563 4922 7564 4962
rect 7604 4922 7605 4962
rect 9483 4936 9484 4976
rect 9524 4936 9525 4976
rect 9483 4927 9525 4936
rect 9579 4976 9621 4985
rect 9579 4936 9580 4976
rect 9620 4936 9621 4976
rect 9579 4927 9621 4936
rect 9963 4976 10005 4985
rect 9963 4936 9964 4976
rect 10004 4936 10005 4976
rect 9963 4927 10005 4936
rect 10059 4976 10101 4985
rect 10059 4936 10060 4976
rect 10100 4936 10101 4976
rect 10059 4927 10101 4936
rect 10531 4976 10589 4977
rect 10531 4936 10540 4976
rect 10580 4936 10589 4976
rect 10531 4935 10589 4936
rect 11019 4971 11061 4980
rect 11019 4931 11020 4971
rect 11060 4931 11061 4971
rect 12451 4976 12509 4977
rect 12451 4936 12460 4976
rect 12500 4936 12509 4976
rect 12451 4935 12509 4936
rect 13699 4976 13757 4977
rect 13699 4936 13708 4976
rect 13748 4936 13757 4976
rect 13699 4935 13757 4936
rect 18307 4976 18365 4977
rect 18307 4936 18316 4976
rect 18356 4936 18365 4976
rect 18307 4935 18365 4936
rect 19555 4976 19613 4977
rect 19555 4936 19564 4976
rect 19604 4936 19613 4976
rect 19555 4935 19613 4936
rect 21387 4976 21429 4985
rect 21387 4936 21388 4976
rect 21428 4936 21429 4976
rect 11019 4922 11061 4931
rect 21387 4927 21429 4936
rect 21483 4976 21525 4985
rect 21483 4936 21484 4976
rect 21524 4936 21525 4976
rect 21483 4927 21525 4936
rect 21963 4976 22005 4985
rect 21963 4936 21964 4976
rect 22004 4936 22005 4976
rect 21963 4927 22005 4936
rect 22435 4976 22493 4977
rect 22435 4936 22444 4976
rect 22484 4936 22493 4976
rect 23875 4976 23933 4977
rect 22435 4935 22493 4936
rect 22971 4966 23013 4975
rect 22971 4926 22972 4966
rect 23012 4926 23013 4966
rect 23875 4936 23884 4976
rect 23924 4936 23933 4976
rect 23875 4935 23933 4936
rect 25123 4976 25181 4977
rect 25123 4936 25132 4976
rect 25172 4936 25181 4976
rect 25123 4935 25181 4936
rect 27147 4976 27189 4985
rect 27147 4936 27148 4976
rect 27188 4936 27189 4976
rect 27147 4927 27189 4936
rect 27243 4976 27285 4985
rect 27243 4936 27244 4976
rect 27284 4936 27285 4976
rect 27243 4927 27285 4936
rect 27627 4976 27669 4985
rect 27627 4936 27628 4976
rect 27668 4936 27669 4976
rect 27627 4927 27669 4936
rect 27723 4976 27765 4985
rect 27723 4936 27724 4976
rect 27764 4936 27765 4976
rect 27723 4927 27765 4936
rect 28195 4976 28253 4977
rect 28195 4936 28204 4976
rect 28244 4936 28253 4976
rect 29259 4976 29301 4985
rect 28195 4935 28253 4936
rect 28731 4966 28773 4975
rect 7563 4913 7605 4922
rect 22971 4917 23013 4926
rect 28731 4926 28732 4966
rect 28772 4926 28773 4966
rect 28731 4917 28773 4926
rect 29163 4957 29205 4966
rect 29163 4917 29164 4957
rect 29204 4917 29205 4957
rect 29259 4936 29260 4976
rect 29300 4936 29301 4976
rect 29259 4927 29301 4936
rect 29643 4976 29685 4985
rect 29643 4936 29644 4976
rect 29684 4936 29685 4976
rect 29643 4927 29685 4936
rect 30211 4976 30269 4977
rect 30211 4936 30220 4976
rect 30260 4936 30269 4976
rect 32035 4976 32093 4977
rect 30211 4935 30269 4936
rect 30699 4962 30741 4971
rect 29163 4908 29205 4917
rect 30699 4922 30700 4962
rect 30740 4922 30741 4962
rect 32035 4936 32044 4976
rect 32084 4936 32093 4976
rect 32035 4935 32093 4936
rect 33283 4976 33341 4977
rect 33283 4936 33292 4976
rect 33332 4936 33341 4976
rect 33283 4935 33341 4936
rect 34339 4976 34397 4977
rect 34339 4936 34348 4976
rect 34388 4936 34397 4976
rect 34339 4935 34397 4936
rect 35587 4976 35645 4977
rect 35587 4936 35596 4976
rect 35636 4936 35645 4976
rect 35587 4935 35645 4936
rect 37219 4976 37277 4977
rect 37219 4936 37228 4976
rect 37268 4936 37277 4976
rect 37219 4935 37277 4936
rect 38467 4976 38525 4977
rect 38467 4936 38476 4976
rect 38516 4936 38525 4976
rect 38467 4935 38525 4936
rect 39043 4976 39101 4977
rect 39043 4936 39052 4976
rect 39092 4936 39101 4976
rect 39043 4935 39101 4936
rect 40291 4976 40349 4977
rect 40291 4936 40300 4976
rect 40340 4936 40349 4976
rect 40291 4935 40349 4936
rect 30699 4913 30741 4922
rect 11683 4892 11741 4893
rect 11683 4852 11692 4892
rect 11732 4852 11741 4892
rect 11683 4851 11741 4852
rect 12259 4892 12317 4893
rect 12259 4852 12268 4892
rect 12308 4852 12317 4892
rect 12259 4851 12317 4852
rect 14851 4892 14909 4893
rect 14851 4852 14860 4892
rect 14900 4852 14909 4892
rect 14851 4851 14909 4852
rect 16963 4892 17021 4893
rect 16963 4852 16972 4892
rect 17012 4852 17021 4892
rect 16963 4851 17021 4852
rect 17155 4892 17213 4893
rect 17155 4852 17164 4892
rect 17204 4852 17213 4892
rect 17155 4851 17213 4852
rect 21091 4892 21149 4893
rect 21091 4852 21100 4892
rect 21140 4852 21149 4892
rect 21091 4851 21149 4852
rect 21867 4892 21909 4901
rect 21867 4852 21868 4892
rect 21908 4852 21909 4892
rect 21867 4843 21909 4852
rect 29739 4892 29781 4901
rect 29739 4852 29740 4892
rect 29780 4852 29781 4892
rect 29739 4843 29781 4852
rect 36835 4892 36893 4893
rect 36835 4852 36844 4892
rect 36884 4852 36893 4892
rect 36835 4851 36893 4852
rect 40675 4892 40733 4893
rect 40675 4852 40684 4892
rect 40724 4852 40733 4892
rect 40675 4851 40733 4852
rect 40867 4892 40925 4893
rect 40867 4852 40876 4892
rect 40916 4852 40925 4892
rect 40867 4851 40925 4852
rect 41251 4892 41309 4893
rect 41251 4852 41260 4892
rect 41300 4852 41309 4892
rect 41251 4851 41309 4852
rect 3147 4808 3189 4817
rect 3147 4768 3148 4808
rect 3188 4768 3189 4808
rect 3147 4759 3189 4768
rect 11883 4808 11925 4817
rect 11883 4768 11884 4808
rect 11924 4768 11925 4808
rect 11883 4759 11925 4768
rect 14667 4808 14709 4817
rect 14667 4768 14668 4808
rect 14708 4768 14709 4808
rect 14667 4759 14709 4768
rect 16779 4808 16821 4817
rect 16779 4768 16780 4808
rect 16820 4768 16821 4808
rect 16779 4759 16821 4768
rect 17355 4808 17397 4817
rect 17355 4768 17356 4808
rect 17396 4768 17397 4808
rect 17355 4759 17397 4768
rect 20907 4808 20949 4817
rect 20907 4768 20908 4808
rect 20948 4768 20949 4808
rect 20907 4759 20949 4768
rect 36651 4808 36693 4817
rect 36651 4768 36652 4808
rect 36692 4768 36693 4808
rect 36651 4759 36693 4768
rect 41067 4808 41109 4817
rect 41067 4768 41068 4808
rect 41108 4768 41109 4808
rect 41067 4759 41109 4768
rect 41451 4808 41493 4817
rect 41451 4768 41452 4808
rect 41492 4768 41493 4808
rect 41451 4759 41493 4768
rect 4107 4724 4149 4733
rect 4107 4684 4108 4724
rect 4148 4684 4149 4724
rect 4107 4675 4149 4684
rect 4875 4724 4917 4733
rect 4875 4684 4876 4724
rect 4916 4684 4917 4724
rect 4875 4675 4917 4684
rect 12075 4724 12117 4733
rect 12075 4684 12076 4724
rect 12116 4684 12117 4724
rect 12075 4675 12117 4684
rect 25323 4724 25365 4733
rect 25323 4684 25324 4724
rect 25364 4684 25365 4724
rect 25323 4675 25365 4684
rect 38859 4724 38901 4733
rect 38859 4684 38860 4724
rect 38900 4684 38901 4724
rect 38859 4675 38901 4684
rect 40491 4724 40533 4733
rect 40491 4684 40492 4724
rect 40532 4684 40533 4724
rect 40491 4675 40533 4684
rect 1152 4556 41856 4580
rect 1152 4516 3688 4556
rect 3728 4516 3770 4556
rect 3810 4516 3852 4556
rect 3892 4516 3934 4556
rect 3974 4516 4016 4556
rect 4056 4516 18808 4556
rect 18848 4516 18890 4556
rect 18930 4516 18972 4556
rect 19012 4516 19054 4556
rect 19094 4516 19136 4556
rect 19176 4516 33928 4556
rect 33968 4516 34010 4556
rect 34050 4516 34092 4556
rect 34132 4516 34174 4556
rect 34214 4516 34256 4556
rect 34296 4516 41856 4556
rect 1152 4492 41856 4516
rect 28971 4388 29013 4397
rect 28971 4348 28972 4388
rect 29012 4348 29013 4388
rect 28971 4339 29013 4348
rect 32043 4388 32085 4397
rect 32043 4348 32044 4388
rect 32084 4348 32085 4388
rect 32043 4339 32085 4348
rect 40683 4388 40725 4397
rect 40683 4348 40684 4388
rect 40724 4348 40725 4388
rect 40683 4339 40725 4348
rect 41067 4388 41109 4397
rect 41067 4348 41068 4388
rect 41108 4348 41109 4388
rect 41067 4339 41109 4348
rect 4771 4304 4829 4305
rect 4771 4264 4780 4304
rect 4820 4264 4829 4304
rect 4771 4263 4829 4264
rect 29451 4304 29493 4313
rect 29451 4264 29452 4304
rect 29492 4264 29493 4304
rect 29451 4255 29493 4264
rect 7371 4220 7413 4229
rect 7371 4180 7372 4220
rect 7412 4180 7413 4220
rect 7371 4171 7413 4180
rect 7467 4220 7509 4229
rect 7467 4180 7468 4220
rect 7508 4180 7509 4220
rect 7467 4171 7509 4180
rect 11403 4220 11445 4229
rect 11403 4180 11404 4220
rect 11444 4180 11445 4220
rect 11403 4171 11445 4180
rect 11499 4220 11541 4229
rect 11499 4180 11500 4220
rect 11540 4180 11541 4220
rect 11499 4171 11541 4180
rect 13707 4220 13749 4229
rect 13707 4180 13708 4220
rect 13748 4180 13749 4220
rect 13707 4171 13749 4180
rect 20331 4220 20373 4229
rect 20331 4180 20332 4220
rect 20372 4180 20373 4220
rect 20331 4171 20373 4180
rect 23883 4220 23925 4229
rect 23883 4180 23884 4220
rect 23924 4180 23925 4220
rect 23883 4171 23925 4180
rect 23979 4220 24021 4229
rect 23979 4180 23980 4220
rect 24020 4180 24021 4220
rect 25899 4220 25941 4229
rect 23979 4171 24021 4180
rect 24987 4178 25029 4187
rect 1603 4136 1661 4137
rect 1603 4096 1612 4136
rect 1652 4096 1661 4136
rect 1603 4095 1661 4096
rect 2851 4136 2909 4137
rect 2851 4096 2860 4136
rect 2900 4096 2909 4136
rect 2851 4095 2909 4096
rect 3531 4136 3573 4145
rect 3531 4096 3532 4136
rect 3572 4096 3573 4136
rect 3531 4087 3573 4096
rect 3723 4136 3765 4145
rect 3723 4096 3724 4136
rect 3764 4096 3765 4136
rect 3723 4087 3765 4096
rect 3811 4136 3869 4137
rect 3811 4096 3820 4136
rect 3860 4096 3869 4136
rect 3811 4095 3869 4096
rect 4099 4136 4157 4137
rect 4099 4096 4108 4136
rect 4148 4096 4157 4136
rect 4099 4095 4157 4096
rect 4395 4136 4437 4145
rect 4395 4096 4396 4136
rect 4436 4096 4437 4136
rect 4395 4087 4437 4096
rect 4491 4136 4533 4145
rect 4491 4096 4492 4136
rect 4532 4096 4533 4136
rect 4491 4087 4533 4096
rect 5067 4136 5109 4145
rect 5067 4096 5068 4136
rect 5108 4096 5109 4136
rect 5067 4087 5109 4096
rect 5163 4136 5205 4145
rect 5163 4096 5164 4136
rect 5204 4096 5205 4136
rect 5163 4087 5205 4096
rect 5259 4136 5301 4145
rect 5259 4096 5260 4136
rect 5300 4096 5301 4136
rect 5259 4087 5301 4096
rect 5451 4136 5493 4145
rect 5451 4096 5452 4136
rect 5492 4096 5493 4136
rect 5451 4087 5493 4096
rect 5547 4136 5589 4145
rect 5547 4096 5548 4136
rect 5588 4096 5589 4136
rect 5547 4087 5589 4096
rect 5643 4136 5685 4145
rect 5643 4096 5644 4136
rect 5684 4096 5685 4136
rect 5643 4087 5685 4096
rect 5931 4136 5973 4145
rect 5931 4096 5932 4136
rect 5972 4096 5973 4136
rect 5931 4087 5973 4096
rect 6027 4136 6069 4145
rect 6027 4096 6028 4136
rect 6068 4096 6069 4136
rect 6027 4087 6069 4096
rect 6123 4136 6165 4145
rect 6123 4096 6124 4136
rect 6164 4096 6165 4136
rect 6123 4087 6165 4096
rect 6891 4136 6933 4145
rect 6891 4096 6892 4136
rect 6932 4096 6933 4136
rect 6891 4087 6933 4096
rect 6987 4136 7029 4145
rect 8427 4141 8469 4150
rect 6987 4096 6988 4136
rect 7028 4096 7029 4136
rect 6987 4087 7029 4096
rect 7939 4136 7997 4137
rect 7939 4096 7948 4136
rect 7988 4096 7997 4136
rect 7939 4095 7997 4096
rect 8427 4101 8428 4141
rect 8468 4101 8469 4141
rect 8427 4092 8469 4101
rect 10923 4136 10965 4145
rect 10923 4096 10924 4136
rect 10964 4096 10965 4136
rect 10923 4087 10965 4096
rect 11019 4136 11061 4145
rect 12459 4141 12501 4150
rect 11019 4096 11020 4136
rect 11060 4096 11061 4136
rect 11019 4087 11061 4096
rect 11971 4136 12029 4137
rect 11971 4096 11980 4136
rect 12020 4096 12029 4136
rect 11971 4095 12029 4096
rect 12459 4101 12460 4141
rect 12500 4101 12501 4141
rect 12459 4092 12501 4101
rect 13131 4136 13173 4145
rect 13131 4096 13132 4136
rect 13172 4096 13173 4136
rect 13131 4087 13173 4096
rect 13227 4136 13269 4145
rect 13227 4096 13228 4136
rect 13268 4096 13269 4136
rect 13227 4087 13269 4096
rect 13611 4136 13653 4145
rect 14667 4141 14709 4150
rect 13611 4096 13612 4136
rect 13652 4096 13653 4136
rect 13611 4087 13653 4096
rect 14179 4136 14237 4137
rect 14179 4096 14188 4136
rect 14228 4096 14237 4136
rect 14179 4095 14237 4096
rect 14667 4101 14668 4141
rect 14708 4101 14709 4141
rect 14667 4092 14709 4101
rect 15435 4136 15477 4145
rect 15435 4096 15436 4136
rect 15476 4096 15477 4136
rect 15435 4087 15477 4096
rect 15531 4136 15573 4145
rect 15531 4096 15532 4136
rect 15572 4096 15573 4136
rect 15531 4087 15573 4096
rect 15915 4136 15957 4145
rect 15915 4096 15916 4136
rect 15956 4096 15957 4136
rect 15915 4087 15957 4096
rect 16011 4136 16053 4145
rect 16971 4141 17013 4150
rect 16011 4096 16012 4136
rect 16052 4096 16053 4136
rect 16011 4087 16053 4096
rect 16483 4136 16541 4137
rect 16483 4096 16492 4136
rect 16532 4096 16541 4136
rect 16483 4095 16541 4096
rect 16971 4101 16972 4141
rect 17012 4101 17013 4141
rect 16971 4092 17013 4101
rect 19851 4136 19893 4145
rect 19851 4096 19852 4136
rect 19892 4096 19893 4136
rect 19851 4087 19893 4096
rect 19947 4136 19989 4145
rect 19947 4096 19948 4136
rect 19988 4096 19989 4136
rect 19947 4087 19989 4096
rect 20427 4136 20469 4145
rect 21387 4141 21429 4150
rect 20427 4096 20428 4136
rect 20468 4096 20469 4136
rect 20427 4087 20469 4096
rect 20899 4136 20957 4137
rect 20899 4096 20908 4136
rect 20948 4096 20957 4136
rect 20899 4095 20957 4096
rect 21387 4101 21388 4141
rect 21428 4101 21429 4141
rect 21387 4092 21429 4101
rect 23403 4136 23445 4145
rect 23403 4096 23404 4136
rect 23444 4096 23445 4136
rect 23403 4087 23445 4096
rect 23499 4136 23541 4145
rect 24987 4138 24988 4178
rect 25028 4138 25029 4178
rect 25899 4180 25900 4220
rect 25940 4180 25941 4220
rect 25899 4171 25941 4180
rect 25995 4220 26037 4229
rect 25995 4180 25996 4220
rect 26036 4180 26037 4220
rect 25995 4171 26037 4180
rect 34339 4220 34397 4221
rect 34339 4180 34348 4220
rect 34388 4180 34397 4220
rect 34339 4179 34397 4180
rect 35403 4220 35445 4229
rect 35403 4180 35404 4220
rect 35444 4180 35445 4220
rect 35403 4171 35445 4180
rect 37027 4220 37085 4221
rect 37027 4180 37036 4220
rect 37076 4180 37085 4220
rect 37027 4179 37085 4180
rect 38379 4220 38421 4229
rect 38379 4180 38380 4220
rect 38420 4180 38421 4220
rect 38379 4171 38421 4180
rect 38475 4220 38517 4229
rect 38475 4180 38476 4220
rect 38516 4180 38517 4220
rect 38475 4171 38517 4180
rect 40483 4220 40541 4221
rect 40483 4180 40492 4220
rect 40532 4180 40541 4220
rect 40483 4179 40541 4180
rect 40867 4220 40925 4221
rect 40867 4180 40876 4220
rect 40916 4180 40925 4220
rect 40867 4179 40925 4180
rect 41251 4220 41309 4221
rect 41251 4180 41260 4220
rect 41300 4180 41309 4220
rect 41251 4179 41309 4180
rect 23499 4096 23500 4136
rect 23540 4096 23541 4136
rect 23499 4087 23541 4096
rect 24451 4136 24509 4137
rect 24451 4096 24460 4136
rect 24500 4096 24509 4136
rect 24987 4129 25029 4138
rect 25419 4136 25461 4145
rect 24451 4095 24509 4096
rect 25419 4096 25420 4136
rect 25460 4096 25461 4136
rect 25419 4087 25461 4096
rect 25515 4136 25557 4145
rect 26955 4141 26997 4150
rect 36507 4145 36549 4154
rect 39435 4150 39477 4159
rect 25515 4096 25516 4136
rect 25556 4096 25557 4136
rect 25515 4087 25557 4096
rect 26467 4136 26525 4137
rect 26467 4096 26476 4136
rect 26516 4096 26525 4136
rect 26467 4095 26525 4096
rect 26955 4101 26956 4141
rect 26996 4101 26997 4141
rect 26955 4092 26997 4101
rect 27523 4136 27581 4137
rect 27523 4096 27532 4136
rect 27572 4096 27581 4136
rect 27523 4095 27581 4096
rect 28771 4136 28829 4137
rect 28771 4096 28780 4136
rect 28820 4096 28829 4136
rect 28771 4095 28829 4096
rect 30115 4136 30173 4137
rect 30115 4096 30124 4136
rect 30164 4096 30173 4136
rect 30115 4095 30173 4096
rect 30595 4136 30653 4137
rect 30595 4096 30604 4136
rect 30644 4096 30653 4136
rect 30595 4095 30653 4096
rect 31843 4136 31901 4137
rect 31843 4096 31852 4136
rect 31892 4096 31901 4136
rect 31843 4095 31901 4096
rect 32515 4136 32573 4137
rect 32515 4096 32524 4136
rect 32564 4096 32573 4136
rect 32515 4095 32573 4096
rect 33763 4136 33821 4137
rect 33763 4096 33772 4136
rect 33812 4096 33821 4136
rect 33763 4095 33821 4096
rect 34923 4136 34965 4145
rect 34923 4096 34924 4136
rect 34964 4096 34965 4136
rect 34923 4087 34965 4096
rect 35019 4136 35061 4145
rect 35019 4096 35020 4136
rect 35060 4096 35061 4136
rect 35019 4087 35061 4096
rect 35499 4136 35541 4145
rect 35499 4096 35500 4136
rect 35540 4096 35541 4136
rect 35499 4087 35541 4096
rect 35971 4136 36029 4137
rect 35971 4096 35980 4136
rect 36020 4096 36029 4136
rect 36507 4105 36508 4145
rect 36548 4105 36549 4145
rect 36507 4096 36549 4105
rect 37899 4136 37941 4145
rect 37899 4096 37900 4136
rect 37940 4096 37941 4136
rect 35971 4095 36029 4096
rect 37899 4087 37941 4096
rect 37995 4136 38037 4145
rect 37995 4096 37996 4136
rect 38036 4096 38037 4136
rect 37995 4087 38037 4096
rect 38947 4136 39005 4137
rect 38947 4096 38956 4136
rect 38996 4096 39005 4136
rect 39435 4110 39436 4150
rect 39476 4110 39477 4150
rect 39435 4101 39477 4110
rect 38947 4095 39005 4096
rect 12651 4052 12693 4061
rect 12651 4012 12652 4052
rect 12692 4012 12693 4052
rect 12651 4003 12693 4012
rect 14859 4052 14901 4061
rect 14859 4012 14860 4052
rect 14900 4012 14901 4052
rect 14859 4003 14901 4012
rect 17163 4052 17205 4061
rect 17163 4012 17164 4052
rect 17204 4012 17205 4052
rect 17163 4003 17205 4012
rect 21579 4052 21621 4061
rect 21579 4012 21580 4052
rect 21620 4012 21621 4052
rect 21579 4003 21621 4012
rect 25131 4052 25173 4061
rect 25131 4012 25132 4052
rect 25172 4012 25173 4052
rect 25131 4003 25173 4012
rect 36651 4052 36693 4061
rect 36651 4012 36652 4052
rect 36692 4012 36693 4052
rect 36651 4003 36693 4012
rect 39627 4052 39669 4061
rect 39627 4012 39628 4052
rect 39668 4012 39669 4052
rect 39627 4003 39669 4012
rect 3051 3968 3093 3977
rect 3051 3928 3052 3968
rect 3092 3928 3093 3968
rect 3051 3919 3093 3928
rect 3619 3968 3677 3969
rect 3619 3928 3628 3968
rect 3668 3928 3677 3968
rect 3619 3927 3677 3928
rect 4963 3968 5021 3969
rect 4963 3928 4972 3968
rect 5012 3928 5021 3968
rect 4963 3927 5021 3928
rect 5731 3968 5789 3969
rect 5731 3928 5740 3968
rect 5780 3928 5789 3968
rect 5731 3927 5789 3928
rect 6211 3968 6269 3969
rect 6211 3928 6220 3968
rect 6260 3928 6269 3968
rect 6211 3927 6269 3928
rect 8619 3968 8661 3977
rect 8619 3928 8620 3968
rect 8660 3928 8661 3968
rect 8619 3919 8661 3928
rect 27147 3968 27189 3977
rect 27147 3928 27148 3968
rect 27188 3928 27189 3968
rect 27147 3919 27189 3928
rect 33963 3968 34005 3977
rect 33963 3928 33964 3968
rect 34004 3928 34005 3968
rect 33963 3919 34005 3928
rect 34155 3968 34197 3977
rect 34155 3928 34156 3968
rect 34196 3928 34197 3968
rect 34155 3919 34197 3928
rect 36843 3968 36885 3977
rect 36843 3928 36844 3968
rect 36884 3928 36885 3968
rect 36843 3919 36885 3928
rect 41451 3968 41493 3977
rect 41451 3928 41452 3968
rect 41492 3928 41493 3968
rect 41451 3919 41493 3928
rect 1152 3800 41856 3824
rect 1152 3760 4928 3800
rect 4968 3760 5010 3800
rect 5050 3760 5092 3800
rect 5132 3760 5174 3800
rect 5214 3760 5256 3800
rect 5296 3760 20048 3800
rect 20088 3760 20130 3800
rect 20170 3760 20212 3800
rect 20252 3760 20294 3800
rect 20334 3760 20376 3800
rect 20416 3760 35168 3800
rect 35208 3760 35250 3800
rect 35290 3760 35332 3800
rect 35372 3760 35414 3800
rect 35454 3760 35496 3800
rect 35536 3760 41856 3800
rect 1152 3736 41856 3760
rect 4579 3632 4637 3633
rect 4579 3592 4588 3632
rect 4628 3592 4637 3632
rect 4579 3591 4637 3592
rect 4867 3632 4925 3633
rect 4867 3592 4876 3632
rect 4916 3592 4925 3632
rect 4867 3591 4925 3592
rect 11499 3632 11541 3641
rect 11499 3592 11500 3632
rect 11540 3592 11541 3632
rect 11499 3583 11541 3592
rect 13707 3632 13749 3641
rect 13707 3592 13708 3632
rect 13748 3592 13749 3632
rect 13707 3583 13749 3592
rect 15339 3632 15381 3641
rect 15339 3592 15340 3632
rect 15380 3592 15381 3632
rect 15339 3583 15381 3592
rect 16971 3632 17013 3641
rect 16971 3592 16972 3632
rect 17012 3592 17013 3632
rect 16971 3583 17013 3592
rect 17739 3632 17781 3641
rect 17739 3592 17740 3632
rect 17780 3592 17781 3632
rect 17739 3583 17781 3592
rect 17931 3632 17973 3641
rect 17931 3592 17932 3632
rect 17972 3592 17973 3632
rect 17931 3583 17973 3592
rect 19755 3632 19797 3641
rect 19755 3592 19756 3632
rect 19796 3592 19797 3632
rect 19755 3583 19797 3592
rect 21483 3632 21525 3641
rect 21483 3592 21484 3632
rect 21524 3592 21525 3632
rect 21483 3583 21525 3592
rect 27339 3632 27381 3641
rect 27339 3592 27340 3632
rect 27380 3592 27381 3632
rect 27339 3583 27381 3592
rect 30795 3632 30837 3641
rect 30795 3592 30796 3632
rect 30836 3592 30837 3632
rect 30795 3583 30837 3592
rect 31563 3632 31605 3641
rect 31563 3592 31564 3632
rect 31604 3592 31605 3632
rect 31563 3583 31605 3592
rect 34347 3632 34389 3641
rect 34347 3592 34348 3632
rect 34388 3592 34389 3632
rect 34347 3583 34389 3592
rect 37035 3632 37077 3641
rect 37035 3592 37036 3632
rect 37076 3592 37077 3632
rect 37035 3583 37077 3592
rect 37323 3632 37365 3641
rect 37323 3592 37324 3632
rect 37364 3592 37365 3632
rect 37323 3583 37365 3592
rect 41067 3632 41109 3641
rect 41067 3592 41068 3632
rect 41108 3592 41109 3632
rect 41067 3583 41109 3592
rect 3051 3548 3093 3557
rect 3051 3508 3052 3548
rect 3092 3508 3093 3548
rect 3051 3499 3093 3508
rect 6987 3548 7029 3557
rect 6987 3508 6988 3548
rect 7028 3508 7029 3548
rect 6987 3499 7029 3508
rect 24459 3548 24501 3557
rect 24459 3508 24460 3548
rect 24500 3508 24501 3548
rect 24459 3499 24501 3508
rect 1603 3464 1661 3465
rect 1603 3424 1612 3464
rect 1652 3424 1661 3464
rect 1603 3423 1661 3424
rect 2851 3464 2909 3465
rect 2851 3424 2860 3464
rect 2900 3424 2909 3464
rect 2851 3423 2909 3424
rect 3627 3464 3669 3473
rect 3627 3424 3628 3464
rect 3668 3424 3669 3464
rect 3627 3415 3669 3424
rect 3723 3464 3765 3473
rect 3723 3424 3724 3464
rect 3764 3424 3765 3464
rect 3723 3415 3765 3424
rect 3819 3464 3861 3473
rect 3819 3424 3820 3464
rect 3860 3424 3861 3464
rect 3819 3415 3861 3424
rect 3915 3464 3957 3473
rect 3915 3424 3916 3464
rect 3956 3424 3957 3464
rect 3915 3415 3957 3424
rect 4099 3464 4157 3465
rect 4099 3424 4108 3464
rect 4148 3424 4157 3464
rect 4099 3423 4157 3424
rect 4195 3464 4253 3465
rect 4195 3424 4204 3464
rect 4244 3424 4253 3464
rect 4195 3423 4253 3424
rect 4395 3464 4437 3473
rect 4395 3424 4396 3464
rect 4436 3424 4437 3464
rect 4395 3415 4437 3424
rect 4491 3464 4533 3473
rect 4491 3424 4492 3464
rect 4532 3424 4533 3464
rect 4491 3415 4533 3424
rect 4638 3464 4696 3465
rect 4638 3424 4647 3464
rect 4687 3424 4696 3464
rect 4638 3423 4696 3424
rect 5067 3464 5109 3473
rect 5067 3424 5068 3464
rect 5108 3424 5109 3464
rect 5067 3415 5109 3424
rect 5163 3464 5205 3473
rect 5163 3424 5164 3464
rect 5204 3424 5205 3464
rect 5163 3415 5205 3424
rect 7083 3464 7125 3473
rect 7083 3424 7084 3464
rect 7124 3424 7125 3464
rect 7083 3415 7125 3424
rect 7363 3464 7421 3465
rect 7363 3424 7372 3464
rect 7412 3424 7421 3464
rect 7363 3423 7421 3424
rect 9771 3464 9813 3473
rect 9771 3424 9772 3464
rect 9812 3424 9813 3464
rect 9771 3415 9813 3424
rect 9867 3464 9909 3473
rect 9867 3424 9868 3464
rect 9908 3424 9909 3464
rect 9867 3415 9909 3424
rect 10251 3464 10293 3473
rect 10251 3424 10252 3464
rect 10292 3424 10293 3464
rect 10251 3415 10293 3424
rect 10347 3464 10389 3473
rect 10347 3424 10348 3464
rect 10388 3424 10389 3464
rect 10347 3415 10389 3424
rect 10819 3464 10877 3465
rect 10819 3424 10828 3464
rect 10868 3424 10877 3464
rect 12259 3464 12317 3465
rect 10819 3423 10877 3424
rect 11307 3450 11349 3459
rect 11307 3410 11308 3450
rect 11348 3410 11349 3450
rect 12259 3424 12268 3464
rect 12308 3424 12317 3464
rect 12259 3423 12317 3424
rect 13507 3464 13565 3465
rect 13507 3424 13516 3464
rect 13556 3424 13565 3464
rect 13507 3423 13565 3424
rect 13891 3464 13949 3465
rect 13891 3424 13900 3464
rect 13940 3424 13949 3464
rect 13891 3423 13949 3424
rect 15139 3464 15197 3465
rect 15139 3424 15148 3464
rect 15188 3424 15197 3464
rect 15139 3423 15197 3424
rect 15523 3464 15581 3465
rect 15523 3424 15532 3464
rect 15572 3424 15581 3464
rect 15523 3423 15581 3424
rect 16771 3464 16829 3465
rect 16771 3424 16780 3464
rect 16820 3424 16829 3464
rect 16771 3423 16829 3424
rect 18307 3464 18365 3465
rect 18307 3424 18316 3464
rect 18356 3424 18365 3464
rect 18307 3423 18365 3424
rect 19555 3464 19613 3465
rect 19555 3424 19564 3464
rect 19604 3424 19613 3464
rect 19555 3423 19613 3424
rect 20035 3464 20093 3465
rect 20035 3424 20044 3464
rect 20084 3424 20093 3464
rect 20035 3423 20093 3424
rect 21283 3464 21341 3465
rect 21283 3424 21292 3464
rect 21332 3424 21341 3464
rect 21283 3423 21341 3424
rect 22731 3464 22773 3473
rect 22731 3424 22732 3464
rect 22772 3424 22773 3464
rect 22731 3415 22773 3424
rect 22827 3464 22869 3473
rect 22827 3424 22828 3464
rect 22868 3424 22869 3464
rect 22827 3415 22869 3424
rect 23211 3464 23253 3473
rect 23211 3424 23212 3464
rect 23252 3424 23253 3464
rect 23211 3415 23253 3424
rect 23307 3464 23349 3473
rect 23307 3424 23308 3464
rect 23348 3424 23349 3464
rect 23307 3415 23349 3424
rect 23779 3464 23837 3465
rect 23779 3424 23788 3464
rect 23828 3424 23837 3464
rect 24843 3464 24885 3473
rect 23779 3423 23837 3424
rect 24315 3422 24357 3431
rect 11307 3401 11349 3410
rect 24315 3382 24316 3422
rect 24356 3382 24357 3422
rect 24843 3424 24844 3464
rect 24884 3424 24885 3464
rect 24843 3415 24885 3424
rect 25699 3464 25757 3465
rect 25699 3424 25708 3464
rect 25748 3424 25757 3464
rect 25699 3423 25757 3424
rect 25891 3464 25949 3465
rect 25891 3424 25900 3464
rect 25940 3424 25949 3464
rect 25891 3423 25949 3424
rect 27139 3464 27197 3465
rect 27139 3424 27148 3464
rect 27188 3424 27197 3464
rect 27139 3423 27197 3424
rect 27619 3464 27677 3465
rect 27619 3424 27628 3464
rect 27668 3424 27677 3464
rect 27619 3423 27677 3424
rect 28579 3464 28637 3465
rect 28579 3424 28588 3464
rect 28628 3424 28637 3464
rect 28579 3423 28637 3424
rect 29347 3464 29405 3465
rect 29347 3424 29356 3464
rect 29396 3424 29405 3464
rect 29347 3423 29405 3424
rect 30595 3464 30653 3465
rect 30595 3424 30604 3464
rect 30644 3424 30653 3464
rect 30595 3423 30653 3424
rect 32619 3464 32661 3473
rect 32619 3424 32620 3464
rect 32660 3424 32661 3464
rect 32619 3415 32661 3424
rect 32715 3464 32757 3473
rect 32715 3424 32716 3464
rect 32756 3424 32757 3464
rect 32715 3415 32757 3424
rect 33099 3464 33141 3473
rect 33099 3424 33100 3464
rect 33140 3424 33141 3464
rect 33099 3415 33141 3424
rect 33195 3464 33237 3473
rect 33195 3424 33196 3464
rect 33236 3424 33237 3464
rect 33195 3415 33237 3424
rect 33667 3464 33725 3465
rect 33667 3424 33676 3464
rect 33716 3424 33725 3464
rect 33667 3423 33725 3424
rect 34155 3459 34197 3468
rect 34155 3419 34156 3459
rect 34196 3419 34197 3459
rect 34155 3410 34197 3419
rect 35307 3464 35349 3473
rect 35307 3424 35308 3464
rect 35348 3424 35349 3464
rect 35307 3415 35349 3424
rect 35403 3464 35445 3473
rect 35403 3424 35404 3464
rect 35444 3424 35445 3464
rect 35403 3415 35445 3424
rect 35787 3464 35829 3473
rect 35787 3424 35788 3464
rect 35828 3424 35829 3464
rect 35787 3415 35829 3424
rect 35883 3464 35925 3473
rect 35883 3424 35884 3464
rect 35924 3424 35925 3464
rect 35883 3415 35925 3424
rect 36355 3464 36413 3465
rect 36355 3424 36364 3464
rect 36404 3424 36413 3464
rect 37507 3464 37565 3465
rect 36355 3423 36413 3424
rect 36891 3422 36933 3431
rect 37507 3424 37516 3464
rect 37556 3424 37565 3464
rect 37507 3423 37565 3424
rect 38755 3464 38813 3465
rect 38755 3424 38764 3464
rect 38804 3424 38813 3464
rect 38755 3423 38813 3424
rect 17539 3380 17597 3381
rect 17539 3340 17548 3380
rect 17588 3340 17597 3380
rect 17539 3339 17597 3340
rect 18115 3380 18173 3381
rect 18115 3340 18124 3380
rect 18164 3340 18173 3380
rect 24315 3373 24357 3382
rect 36891 3382 36892 3422
rect 36932 3382 36933 3422
rect 28963 3380 29021 3381
rect 18115 3339 18173 3340
rect 28963 3340 28972 3380
rect 29012 3340 29021 3380
rect 28963 3339 29021 3340
rect 31363 3380 31421 3381
rect 31363 3340 31372 3380
rect 31412 3340 31421 3380
rect 31363 3339 31421 3340
rect 31747 3380 31805 3381
rect 31747 3340 31756 3380
rect 31796 3340 31805 3380
rect 36891 3373 36933 3382
rect 40483 3380 40541 3381
rect 31747 3339 31805 3340
rect 40483 3340 40492 3380
rect 40532 3340 40541 3380
rect 40483 3339 40541 3340
rect 40867 3380 40925 3381
rect 40867 3340 40876 3380
rect 40916 3340 40925 3380
rect 40867 3339 40925 3340
rect 6691 3296 6749 3297
rect 6691 3256 6700 3296
rect 6740 3256 6749 3296
rect 6691 3255 6749 3256
rect 31179 3296 31221 3305
rect 31179 3256 31180 3296
rect 31220 3256 31221 3296
rect 31179 3247 31221 3256
rect 40683 3296 40725 3305
rect 40683 3256 40684 3296
rect 40724 3256 40725 3296
rect 40683 3247 40725 3256
rect 27915 3212 27957 3221
rect 27915 3172 27916 3212
rect 27956 3172 27957 3212
rect 27915 3163 27957 3172
rect 28779 3212 28821 3221
rect 28779 3172 28780 3212
rect 28820 3172 28821 3212
rect 28779 3163 28821 3172
rect 1152 3044 41856 3068
rect 1152 3004 3688 3044
rect 3728 3004 3770 3044
rect 3810 3004 3852 3044
rect 3892 3004 3934 3044
rect 3974 3004 4016 3044
rect 4056 3004 18808 3044
rect 18848 3004 18890 3044
rect 18930 3004 18972 3044
rect 19012 3004 19054 3044
rect 19094 3004 19136 3044
rect 19176 3004 33928 3044
rect 33968 3004 34010 3044
rect 34050 3004 34092 3044
rect 34132 3004 34174 3044
rect 34214 3004 34256 3044
rect 34296 3004 41856 3044
rect 1152 2980 41856 3004
rect 7947 2876 7989 2885
rect 7947 2836 7948 2876
rect 7988 2836 7989 2876
rect 7947 2827 7989 2836
rect 10539 2876 10581 2885
rect 10539 2836 10540 2876
rect 10580 2836 10581 2876
rect 10539 2827 10581 2836
rect 12459 2876 12501 2885
rect 12459 2836 12460 2876
rect 12500 2836 12501 2876
rect 12459 2827 12501 2836
rect 12843 2876 12885 2885
rect 12843 2836 12844 2876
rect 12884 2836 12885 2876
rect 12843 2827 12885 2836
rect 23499 2876 23541 2885
rect 23499 2836 23500 2876
rect 23540 2836 23541 2876
rect 23499 2827 23541 2836
rect 28971 2876 29013 2885
rect 28971 2836 28972 2876
rect 29012 2836 29013 2876
rect 28971 2827 29013 2836
rect 31083 2876 31125 2885
rect 31083 2836 31084 2876
rect 31124 2836 31125 2876
rect 31083 2827 31125 2836
rect 32907 2876 32949 2885
rect 32907 2836 32908 2876
rect 32948 2836 32949 2876
rect 32907 2827 32949 2836
rect 35115 2876 35157 2885
rect 35115 2836 35116 2876
rect 35156 2836 35157 2876
rect 35115 2827 35157 2836
rect 36939 2876 36981 2885
rect 36939 2836 36940 2876
rect 36980 2836 36981 2876
rect 36939 2827 36981 2836
rect 38571 2876 38613 2885
rect 38571 2836 38572 2876
rect 38612 2836 38613 2876
rect 38571 2827 38613 2836
rect 41067 2876 41109 2885
rect 41067 2836 41068 2876
rect 41108 2836 41109 2876
rect 41067 2827 41109 2836
rect 19467 2792 19509 2801
rect 19467 2752 19468 2792
rect 19508 2752 19509 2792
rect 19467 2743 19509 2752
rect 40683 2792 40725 2801
rect 40683 2752 40684 2792
rect 40724 2752 40725 2792
rect 40683 2743 40725 2752
rect 13027 2708 13085 2709
rect 13027 2668 13036 2708
rect 13076 2668 13085 2708
rect 13027 2667 13085 2668
rect 16587 2708 16629 2717
rect 16587 2668 16588 2708
rect 16628 2668 16629 2708
rect 16587 2659 16629 2668
rect 16683 2708 16725 2717
rect 16683 2668 16684 2708
rect 16724 2668 16725 2708
rect 16683 2659 16725 2668
rect 20811 2708 20853 2717
rect 20811 2668 20812 2708
rect 20852 2668 20853 2708
rect 20811 2659 20853 2668
rect 20907 2708 20949 2717
rect 20907 2668 20908 2708
rect 20948 2668 20949 2708
rect 20907 2659 20949 2668
rect 25995 2708 26037 2717
rect 25995 2668 25996 2708
rect 26036 2668 26037 2708
rect 25995 2659 26037 2668
rect 26091 2708 26133 2717
rect 26091 2668 26092 2708
rect 26132 2668 26133 2708
rect 26091 2659 26133 2668
rect 40483 2708 40541 2709
rect 40483 2668 40492 2708
rect 40532 2668 40541 2708
rect 40483 2667 40541 2668
rect 40867 2708 40925 2709
rect 40867 2668 40876 2708
rect 40916 2668 40925 2708
rect 40867 2667 40925 2668
rect 41251 2708 41309 2709
rect 41251 2668 41260 2708
rect 41300 2668 41309 2708
rect 41251 2667 41309 2668
rect 17691 2633 17733 2642
rect 1795 2624 1853 2625
rect 1795 2584 1804 2624
rect 1844 2584 1853 2624
rect 1795 2583 1853 2584
rect 3043 2624 3101 2625
rect 3043 2584 3052 2624
rect 3092 2584 3101 2624
rect 3043 2583 3101 2584
rect 3427 2624 3485 2625
rect 3427 2584 3436 2624
rect 3476 2584 3485 2624
rect 3427 2583 3485 2584
rect 3531 2624 3573 2633
rect 3531 2584 3532 2624
rect 3572 2584 3573 2624
rect 3531 2575 3573 2584
rect 3715 2624 3773 2625
rect 3715 2584 3724 2624
rect 3764 2584 3773 2624
rect 3715 2583 3773 2584
rect 3819 2624 3861 2633
rect 3819 2584 3820 2624
rect 3860 2584 3861 2624
rect 3819 2575 3861 2584
rect 4003 2624 4061 2625
rect 4003 2584 4012 2624
rect 4052 2584 4061 2624
rect 4003 2583 4061 2584
rect 4299 2624 4341 2633
rect 4299 2584 4300 2624
rect 4340 2584 4341 2624
rect 4299 2575 4341 2584
rect 4395 2624 4437 2633
rect 4395 2584 4396 2624
rect 4436 2584 4437 2624
rect 4395 2575 4437 2584
rect 4491 2624 4533 2633
rect 4491 2584 4492 2624
rect 4532 2584 4533 2624
rect 4491 2575 4533 2584
rect 4875 2624 4917 2633
rect 4875 2584 4876 2624
rect 4916 2584 4917 2624
rect 4875 2575 4917 2584
rect 4971 2624 5013 2633
rect 4971 2584 4972 2624
rect 5012 2584 5013 2624
rect 4971 2575 5013 2584
rect 5451 2624 5493 2633
rect 5451 2584 5452 2624
rect 5492 2584 5493 2624
rect 5451 2575 5493 2584
rect 5547 2624 5589 2633
rect 5547 2584 5548 2624
rect 5588 2584 5589 2624
rect 5547 2575 5589 2584
rect 5643 2624 5685 2633
rect 5643 2584 5644 2624
rect 5684 2584 5685 2624
rect 5643 2575 5685 2584
rect 6499 2624 6557 2625
rect 6499 2584 6508 2624
rect 6548 2584 6557 2624
rect 6499 2583 6557 2584
rect 7747 2624 7805 2625
rect 7747 2584 7756 2624
rect 7796 2584 7805 2624
rect 7747 2583 7805 2584
rect 9091 2624 9149 2625
rect 9091 2584 9100 2624
rect 9140 2584 9149 2624
rect 9091 2583 9149 2584
rect 10339 2624 10397 2625
rect 10339 2584 10348 2624
rect 10388 2584 10397 2624
rect 10339 2583 10397 2584
rect 11011 2624 11069 2625
rect 11011 2584 11020 2624
rect 11060 2584 11069 2624
rect 11011 2583 11069 2584
rect 12259 2624 12317 2625
rect 12259 2584 12268 2624
rect 12308 2584 12317 2624
rect 12259 2583 12317 2584
rect 14371 2624 14429 2625
rect 14371 2584 14380 2624
rect 14420 2584 14429 2624
rect 14371 2583 14429 2584
rect 15619 2624 15677 2625
rect 15619 2584 15628 2624
rect 15668 2584 15677 2624
rect 15619 2583 15677 2584
rect 16107 2624 16149 2633
rect 16107 2584 16108 2624
rect 16148 2584 16149 2624
rect 16107 2575 16149 2584
rect 16203 2624 16245 2633
rect 16203 2584 16204 2624
rect 16244 2584 16245 2624
rect 16203 2575 16245 2584
rect 17155 2624 17213 2625
rect 17155 2584 17164 2624
rect 17204 2584 17213 2624
rect 17691 2593 17692 2633
rect 17732 2593 17733 2633
rect 19851 2629 19893 2638
rect 27099 2633 27141 2642
rect 17691 2584 17733 2593
rect 18019 2624 18077 2625
rect 18019 2584 18028 2624
rect 18068 2584 18077 2624
rect 17155 2583 17213 2584
rect 18019 2583 18077 2584
rect 19267 2624 19325 2625
rect 19267 2584 19276 2624
rect 19316 2584 19325 2624
rect 19267 2583 19325 2584
rect 19851 2589 19852 2629
rect 19892 2589 19893 2629
rect 19851 2580 19893 2589
rect 20323 2624 20381 2625
rect 20323 2584 20332 2624
rect 20372 2584 20381 2624
rect 20323 2583 20381 2584
rect 21291 2624 21333 2633
rect 21291 2584 21292 2624
rect 21332 2584 21333 2624
rect 21291 2575 21333 2584
rect 21387 2624 21429 2633
rect 21387 2584 21388 2624
rect 21428 2584 21429 2624
rect 21387 2575 21429 2584
rect 22051 2624 22109 2625
rect 22051 2584 22060 2624
rect 22100 2584 22109 2624
rect 22051 2583 22109 2584
rect 23299 2624 23357 2625
rect 23299 2584 23308 2624
rect 23348 2584 23357 2624
rect 23299 2583 23357 2584
rect 23683 2624 23741 2625
rect 23683 2584 23692 2624
rect 23732 2584 23741 2624
rect 23683 2583 23741 2584
rect 24643 2624 24701 2625
rect 24643 2584 24652 2624
rect 24692 2584 24701 2624
rect 24643 2583 24701 2584
rect 25515 2624 25557 2633
rect 25515 2584 25516 2624
rect 25556 2584 25557 2624
rect 25515 2575 25557 2584
rect 25611 2624 25653 2633
rect 25611 2584 25612 2624
rect 25652 2584 25653 2624
rect 25611 2575 25653 2584
rect 26563 2624 26621 2625
rect 26563 2584 26572 2624
rect 26612 2584 26621 2624
rect 27099 2593 27100 2633
rect 27140 2593 27141 2633
rect 27099 2584 27141 2593
rect 27523 2624 27581 2625
rect 27523 2584 27532 2624
rect 27572 2584 27581 2624
rect 26563 2583 26621 2584
rect 27523 2583 27581 2584
rect 28771 2624 28829 2625
rect 28771 2584 28780 2624
rect 28820 2584 28829 2624
rect 28771 2583 28829 2584
rect 29635 2624 29693 2625
rect 29635 2584 29644 2624
rect 29684 2584 29693 2624
rect 29635 2583 29693 2584
rect 30883 2624 30941 2625
rect 30883 2584 30892 2624
rect 30932 2584 30941 2624
rect 30883 2583 30941 2584
rect 32707 2624 32765 2625
rect 32707 2584 32716 2624
rect 32756 2584 32765 2624
rect 32707 2583 32765 2584
rect 33667 2624 33725 2625
rect 33667 2584 33676 2624
rect 33716 2584 33725 2624
rect 33667 2583 33725 2584
rect 34915 2624 34973 2625
rect 34915 2584 34924 2624
rect 34964 2584 34973 2624
rect 34915 2583 34973 2584
rect 35491 2624 35549 2625
rect 35491 2584 35500 2624
rect 35540 2584 35549 2624
rect 35491 2583 35549 2584
rect 36739 2624 36797 2625
rect 36739 2584 36748 2624
rect 36788 2584 36797 2624
rect 36739 2583 36797 2584
rect 37123 2624 37181 2625
rect 37123 2584 37132 2624
rect 37172 2584 37181 2624
rect 37123 2583 37181 2584
rect 38371 2624 38429 2625
rect 38371 2584 38380 2624
rect 38420 2584 38429 2624
rect 38371 2583 38429 2584
rect 31459 2582 31517 2583
rect 3243 2540 3285 2549
rect 3243 2500 3244 2540
rect 3284 2500 3285 2540
rect 3243 2491 3285 2500
rect 15819 2540 15861 2549
rect 15819 2500 15820 2540
rect 15860 2500 15861 2540
rect 15819 2491 15861 2500
rect 17835 2540 17877 2549
rect 17835 2500 17836 2540
rect 17876 2500 17877 2540
rect 17835 2491 17877 2500
rect 19659 2540 19701 2549
rect 19659 2500 19660 2540
rect 19700 2500 19701 2540
rect 19659 2491 19701 2500
rect 27243 2540 27285 2549
rect 31459 2542 31468 2582
rect 31508 2542 31517 2582
rect 31459 2541 31517 2542
rect 27243 2500 27244 2540
rect 27284 2500 27285 2540
rect 27243 2491 27285 2500
rect 4011 2456 4053 2465
rect 4011 2416 4012 2456
rect 4052 2416 4053 2456
rect 4011 2407 4053 2416
rect 4683 2456 4725 2465
rect 4683 2416 4684 2456
rect 4724 2416 4725 2456
rect 4683 2407 4725 2416
rect 5155 2456 5213 2457
rect 5155 2416 5164 2456
rect 5204 2416 5213 2456
rect 5155 2415 5213 2416
rect 5347 2456 5405 2457
rect 5347 2416 5356 2456
rect 5396 2416 5405 2456
rect 5347 2415 5405 2416
rect 41451 2456 41493 2465
rect 41451 2416 41452 2456
rect 41492 2416 41493 2456
rect 41451 2407 41493 2416
rect 1152 2288 41856 2312
rect 1152 2248 4928 2288
rect 4968 2248 5010 2288
rect 5050 2248 5092 2288
rect 5132 2248 5174 2288
rect 5214 2248 5256 2288
rect 5296 2248 20048 2288
rect 20088 2248 20130 2288
rect 20170 2248 20212 2288
rect 20252 2248 20294 2288
rect 20334 2248 20376 2288
rect 20416 2248 35168 2288
rect 35208 2248 35250 2288
rect 35290 2248 35332 2288
rect 35372 2248 35414 2288
rect 35454 2248 35496 2288
rect 35536 2248 41856 2288
rect 1152 2224 41856 2248
rect 4387 2120 4445 2121
rect 4387 2080 4396 2120
rect 4436 2080 4445 2120
rect 4387 2079 4445 2080
rect 6699 2120 6741 2129
rect 6699 2080 6700 2120
rect 6740 2080 6741 2120
rect 6699 2071 6741 2080
rect 19555 2120 19613 2121
rect 19555 2080 19564 2120
rect 19604 2080 19613 2120
rect 19555 2079 19613 2080
rect 22731 2120 22773 2129
rect 22731 2080 22732 2120
rect 22772 2080 22773 2120
rect 22731 2071 22773 2080
rect 24363 2120 24405 2129
rect 24363 2080 24364 2120
rect 24404 2080 24405 2120
rect 24363 2071 24405 2080
rect 25995 2120 26037 2129
rect 25995 2080 25996 2120
rect 26036 2080 26037 2120
rect 25995 2071 26037 2080
rect 29355 2120 29397 2129
rect 29355 2080 29356 2120
rect 29396 2080 29397 2120
rect 29355 2071 29397 2080
rect 30987 2120 31029 2129
rect 30987 2080 30988 2120
rect 31028 2080 31029 2120
rect 30987 2071 31029 2080
rect 31179 2120 31221 2129
rect 31179 2080 31180 2120
rect 31220 2080 31221 2120
rect 31179 2071 31221 2080
rect 31563 2120 31605 2129
rect 31563 2080 31564 2120
rect 31604 2080 31605 2120
rect 31563 2071 31605 2080
rect 32227 2120 32285 2121
rect 32227 2080 32236 2120
rect 32276 2080 32285 2120
rect 32227 2079 32285 2080
rect 34827 2120 34869 2129
rect 34827 2080 34828 2120
rect 34868 2080 34869 2120
rect 34827 2071 34869 2080
rect 36459 2120 36501 2129
rect 36459 2080 36460 2120
rect 36500 2080 36501 2120
rect 36459 2071 36501 2080
rect 39243 2120 39285 2129
rect 39243 2080 39244 2120
rect 39284 2080 39285 2120
rect 39243 2071 39285 2080
rect 40395 2120 40437 2129
rect 40395 2080 40396 2120
rect 40436 2080 40437 2120
rect 40395 2071 40437 2080
rect 41067 2120 41109 2129
rect 41067 2080 41068 2120
rect 41108 2080 41109 2120
rect 41067 2071 41109 2080
rect 4483 2036 4541 2037
rect 4483 1996 4492 2036
rect 4532 1996 4541 2036
rect 4483 1995 4541 1996
rect 17163 2036 17205 2045
rect 17163 1996 17164 2036
rect 17204 1996 17205 2036
rect 17163 1987 17205 1996
rect 34635 2036 34677 2045
rect 34635 1996 34636 2036
rect 34676 1996 34677 2036
rect 34635 1987 34677 1996
rect 1891 1952 1949 1953
rect 1891 1912 1900 1952
rect 1940 1912 1949 1952
rect 1891 1911 1949 1912
rect 3139 1952 3197 1953
rect 3139 1912 3148 1952
rect 3188 1912 3197 1952
rect 3139 1911 3197 1912
rect 3819 1952 3861 1961
rect 3819 1912 3820 1952
rect 3860 1912 3861 1952
rect 3819 1903 3861 1912
rect 3915 1952 3957 1961
rect 3915 1912 3916 1952
rect 3956 1912 3957 1952
rect 3915 1903 3957 1912
rect 4011 1952 4053 1961
rect 4011 1912 4012 1952
rect 4052 1912 4053 1952
rect 4011 1903 4053 1912
rect 4107 1952 4149 1961
rect 4107 1912 4108 1952
rect 4148 1912 4149 1952
rect 4107 1903 4149 1912
rect 4587 1952 4629 1961
rect 4587 1912 4588 1952
rect 4628 1912 4629 1952
rect 4587 1903 4629 1912
rect 4683 1952 4725 1961
rect 4683 1912 4684 1952
rect 4724 1912 4725 1952
rect 4683 1903 4725 1912
rect 4867 1952 4925 1953
rect 4867 1912 4876 1952
rect 4916 1912 4925 1952
rect 4867 1911 4925 1912
rect 5067 1952 5109 1961
rect 5067 1912 5068 1952
rect 5108 1912 5109 1952
rect 5067 1903 5109 1912
rect 5251 1952 5309 1953
rect 5251 1912 5260 1952
rect 5300 1912 5309 1952
rect 5251 1911 5309 1912
rect 6499 1952 6557 1953
rect 6499 1912 6508 1952
rect 6548 1912 6557 1952
rect 6499 1911 6557 1912
rect 7267 1952 7325 1953
rect 7267 1912 7276 1952
rect 7316 1912 7325 1952
rect 7267 1911 7325 1912
rect 8515 1952 8573 1953
rect 8515 1912 8524 1952
rect 8564 1912 8573 1952
rect 8515 1911 8573 1912
rect 8899 1952 8957 1953
rect 8899 1912 8908 1952
rect 8948 1912 8957 1952
rect 8899 1911 8957 1912
rect 10147 1952 10205 1953
rect 10147 1912 10156 1952
rect 10196 1912 10205 1952
rect 10147 1911 10205 1912
rect 10531 1952 10589 1953
rect 10531 1912 10540 1952
rect 10580 1912 10589 1952
rect 10531 1911 10589 1912
rect 11779 1952 11837 1953
rect 11779 1912 11788 1952
rect 11828 1912 11837 1952
rect 11779 1911 11837 1912
rect 12163 1952 12221 1953
rect 12163 1912 12172 1952
rect 12212 1912 12221 1952
rect 12163 1911 12221 1912
rect 13411 1952 13469 1953
rect 13411 1912 13420 1952
rect 13460 1912 13469 1952
rect 13411 1911 13469 1912
rect 13795 1952 13853 1953
rect 13795 1912 13804 1952
rect 13844 1912 13853 1952
rect 13795 1911 13853 1912
rect 15043 1952 15101 1953
rect 15043 1912 15052 1952
rect 15092 1912 15101 1952
rect 15043 1911 15101 1912
rect 15427 1952 15485 1953
rect 15427 1912 15436 1952
rect 15476 1912 15485 1952
rect 15427 1911 15485 1912
rect 16675 1952 16733 1953
rect 16675 1912 16684 1952
rect 16724 1912 16733 1952
rect 16675 1911 16733 1912
rect 17539 1952 17597 1953
rect 17539 1912 17548 1952
rect 17588 1912 17597 1952
rect 17539 1911 17597 1912
rect 18403 1952 18461 1953
rect 18403 1912 18412 1952
rect 18452 1912 18461 1952
rect 18403 1911 18461 1912
rect 21283 1952 21341 1953
rect 21283 1912 21292 1952
rect 21332 1912 21341 1952
rect 21283 1911 21341 1912
rect 22531 1952 22589 1953
rect 22531 1912 22540 1952
rect 22580 1912 22589 1952
rect 22531 1911 22589 1912
rect 22915 1952 22973 1953
rect 22915 1912 22924 1952
rect 22964 1912 22973 1952
rect 22915 1911 22973 1912
rect 24163 1952 24221 1953
rect 24163 1912 24172 1952
rect 24212 1912 24221 1952
rect 24163 1911 24221 1912
rect 24547 1952 24605 1953
rect 24547 1912 24556 1952
rect 24596 1912 24605 1952
rect 24547 1911 24605 1912
rect 25795 1952 25853 1953
rect 25795 1912 25804 1952
rect 25844 1912 25853 1952
rect 25795 1911 25853 1912
rect 26179 1952 26237 1953
rect 26179 1912 26188 1952
rect 26228 1912 26237 1952
rect 26179 1911 26237 1912
rect 27427 1952 27485 1953
rect 27427 1912 27436 1952
rect 27476 1912 27485 1952
rect 27427 1911 27485 1912
rect 27907 1952 27965 1953
rect 27907 1912 27916 1952
rect 27956 1912 27965 1952
rect 27907 1911 27965 1912
rect 29155 1952 29213 1953
rect 29155 1912 29164 1952
rect 29204 1912 29213 1952
rect 29155 1911 29213 1912
rect 29539 1952 29597 1953
rect 29539 1912 29548 1952
rect 29588 1912 29597 1952
rect 29539 1911 29597 1912
rect 30787 1952 30845 1953
rect 30787 1912 30796 1952
rect 30836 1912 30845 1952
rect 30787 1911 30845 1912
rect 33379 1952 33437 1953
rect 33379 1912 33388 1952
rect 33428 1912 33437 1952
rect 33379 1911 33437 1912
rect 34243 1952 34301 1953
rect 34243 1912 34252 1952
rect 34292 1912 34301 1952
rect 34243 1911 34301 1912
rect 35011 1952 35069 1953
rect 35011 1912 35020 1952
rect 35060 1912 35069 1952
rect 35011 1911 35069 1912
rect 36259 1952 36317 1953
rect 36259 1912 36268 1952
rect 36308 1912 36317 1952
rect 36259 1911 36317 1912
rect 36643 1952 36701 1953
rect 36643 1912 36652 1952
rect 36692 1912 36701 1952
rect 36643 1911 36701 1912
rect 37891 1952 37949 1953
rect 37891 1912 37900 1952
rect 37940 1912 37949 1952
rect 37891 1911 37949 1912
rect 31363 1868 31421 1869
rect 31363 1828 31372 1868
rect 31412 1828 31421 1868
rect 31363 1827 31421 1828
rect 31747 1868 31805 1869
rect 31747 1828 31756 1868
rect 31796 1828 31805 1868
rect 31747 1827 31805 1828
rect 38371 1868 38429 1869
rect 38371 1828 38380 1868
rect 38420 1828 38429 1868
rect 38371 1827 38429 1828
rect 39427 1868 39485 1869
rect 39427 1828 39436 1868
rect 39476 1828 39485 1868
rect 39427 1827 39485 1828
rect 39619 1868 39677 1869
rect 39619 1828 39628 1868
rect 39668 1828 39677 1868
rect 39619 1827 39677 1828
rect 40003 1868 40061 1869
rect 40003 1828 40012 1868
rect 40052 1828 40061 1868
rect 40003 1827 40061 1828
rect 40579 1868 40637 1869
rect 40579 1828 40588 1868
rect 40628 1828 40637 1868
rect 40579 1827 40637 1828
rect 40867 1868 40925 1869
rect 40867 1828 40876 1868
rect 40916 1828 40925 1868
rect 40867 1827 40925 1828
rect 41251 1868 41309 1869
rect 41251 1828 41260 1868
rect 41300 1828 41309 1868
rect 41251 1827 41309 1828
rect 4971 1784 5013 1793
rect 4971 1744 4972 1784
rect 5012 1744 5013 1784
rect 4971 1735 5013 1744
rect 41451 1784 41493 1793
rect 41451 1744 41452 1784
rect 41492 1744 41493 1784
rect 41451 1735 41493 1744
rect 3339 1700 3381 1709
rect 3339 1660 3340 1700
rect 3380 1660 3381 1700
rect 3339 1651 3381 1660
rect 4587 1700 4629 1709
rect 4587 1660 4588 1700
rect 4628 1660 4629 1700
rect 4587 1651 4629 1660
rect 8715 1700 8757 1709
rect 8715 1660 8716 1700
rect 8756 1660 8757 1700
rect 8715 1651 8757 1660
rect 10347 1700 10389 1709
rect 10347 1660 10348 1700
rect 10388 1660 10389 1700
rect 10347 1651 10389 1660
rect 11979 1700 12021 1709
rect 11979 1660 11980 1700
rect 12020 1660 12021 1700
rect 11979 1651 12021 1660
rect 13611 1700 13653 1709
rect 13611 1660 13612 1700
rect 13652 1660 13653 1700
rect 13611 1651 13653 1660
rect 15243 1700 15285 1709
rect 15243 1660 15244 1700
rect 15284 1660 15285 1700
rect 15243 1651 15285 1660
rect 16875 1700 16917 1709
rect 16875 1660 16876 1700
rect 16916 1660 16917 1700
rect 16875 1651 16917 1660
rect 27627 1700 27669 1709
rect 27627 1660 27628 1700
rect 27668 1660 27669 1700
rect 27627 1651 27669 1660
rect 38187 1700 38229 1709
rect 38187 1660 38188 1700
rect 38228 1660 38229 1700
rect 38187 1651 38229 1660
rect 39819 1700 39861 1709
rect 39819 1660 39820 1700
rect 39860 1660 39861 1700
rect 39819 1651 39861 1660
rect 40203 1700 40245 1709
rect 40203 1660 40204 1700
rect 40244 1660 40245 1700
rect 40203 1651 40245 1660
rect 1152 1532 41856 1556
rect 1152 1492 3688 1532
rect 3728 1492 3770 1532
rect 3810 1492 3852 1532
rect 3892 1492 3934 1532
rect 3974 1492 4016 1532
rect 4056 1492 18808 1532
rect 18848 1492 18890 1532
rect 18930 1492 18972 1532
rect 19012 1492 19054 1532
rect 19094 1492 19136 1532
rect 19176 1492 33928 1532
rect 33968 1492 34010 1532
rect 34050 1492 34092 1532
rect 34132 1492 34174 1532
rect 34214 1492 34256 1532
rect 34296 1492 41856 1532
rect 1152 1468 41856 1492
rect 9579 1280 9621 1289
rect 9579 1240 9580 1280
rect 9620 1240 9621 1280
rect 9579 1231 9621 1240
rect 11211 1280 11253 1289
rect 11211 1240 11212 1280
rect 11252 1240 11253 1280
rect 11211 1231 11253 1240
rect 14475 1280 14517 1289
rect 14475 1240 14476 1280
rect 14516 1240 14517 1280
rect 14475 1231 14517 1240
rect 17739 1280 17781 1289
rect 17739 1240 17740 1280
rect 17780 1240 17781 1280
rect 17739 1231 17781 1240
rect 17931 1280 17973 1289
rect 17931 1240 17932 1280
rect 17972 1240 17973 1280
rect 17931 1231 17973 1240
rect 19851 1280 19893 1289
rect 19851 1240 19852 1280
rect 19892 1240 19893 1280
rect 19851 1231 19893 1240
rect 21483 1280 21525 1289
rect 21483 1240 21484 1280
rect 21524 1240 21525 1280
rect 21483 1231 21525 1240
rect 23115 1280 23157 1289
rect 23115 1240 23116 1280
rect 23156 1240 23157 1280
rect 23115 1231 23157 1240
rect 25131 1280 25173 1289
rect 25131 1240 25132 1280
rect 25172 1240 25173 1280
rect 25131 1231 25173 1240
rect 26859 1280 26901 1289
rect 26859 1240 26860 1280
rect 26900 1240 26901 1280
rect 26859 1231 26901 1240
rect 29067 1280 29109 1289
rect 29067 1240 29068 1280
rect 29108 1240 29109 1280
rect 29067 1231 29109 1240
rect 29643 1280 29685 1289
rect 29643 1240 29644 1280
rect 29684 1240 29685 1280
rect 29643 1231 29685 1240
rect 31659 1280 31701 1289
rect 31659 1240 31660 1280
rect 31700 1240 31701 1280
rect 31659 1231 31701 1240
rect 32715 1280 32757 1289
rect 32715 1240 32716 1280
rect 32756 1240 32757 1280
rect 32715 1231 32757 1240
rect 33099 1280 33141 1289
rect 33099 1240 33100 1280
rect 33140 1240 33141 1280
rect 33099 1231 33141 1240
rect 33483 1280 33525 1289
rect 33483 1240 33484 1280
rect 33524 1240 33525 1280
rect 33483 1231 33525 1240
rect 34059 1280 34101 1289
rect 34059 1240 34060 1280
rect 34100 1240 34101 1280
rect 34059 1231 34101 1240
rect 37035 1280 37077 1289
rect 37035 1240 37036 1280
rect 37076 1240 37077 1280
rect 37035 1231 37077 1240
rect 37227 1280 37269 1289
rect 37227 1240 37228 1280
rect 37268 1240 37269 1280
rect 37227 1231 37269 1240
rect 37611 1280 37653 1289
rect 37611 1240 37612 1280
rect 37652 1240 37653 1280
rect 37611 1231 37653 1240
rect 29443 1196 29501 1197
rect 29443 1156 29452 1196
rect 29492 1156 29501 1196
rect 29443 1155 29501 1156
rect 32515 1196 32573 1197
rect 32515 1156 32524 1196
rect 32564 1156 32573 1196
rect 32515 1155 32573 1156
rect 32899 1196 32957 1197
rect 32899 1156 32908 1196
rect 32948 1156 32957 1196
rect 32899 1155 32957 1156
rect 33283 1196 33341 1197
rect 33283 1156 33292 1196
rect 33332 1156 33341 1196
rect 33283 1155 33341 1156
rect 33667 1196 33725 1197
rect 33667 1156 33676 1196
rect 33716 1156 33725 1196
rect 33667 1155 33725 1156
rect 34435 1196 34493 1197
rect 34435 1156 34444 1196
rect 34484 1156 34493 1196
rect 34435 1155 34493 1156
rect 34819 1196 34877 1197
rect 34819 1156 34828 1196
rect 34868 1156 34877 1196
rect 34819 1155 34877 1156
rect 35203 1196 35261 1197
rect 35203 1156 35212 1196
rect 35252 1156 35261 1196
rect 35203 1155 35261 1156
rect 37411 1196 37469 1197
rect 37411 1156 37420 1196
rect 37460 1156 37469 1196
rect 37411 1155 37469 1156
rect 37795 1196 37853 1197
rect 37795 1156 37804 1196
rect 37844 1156 37853 1196
rect 37795 1155 37853 1156
rect 40483 1196 40541 1197
rect 40483 1156 40492 1196
rect 40532 1156 40541 1196
rect 40483 1155 40541 1156
rect 40867 1196 40925 1197
rect 40867 1156 40876 1196
rect 40916 1156 40925 1196
rect 40867 1155 40925 1156
rect 41251 1196 41309 1197
rect 41251 1156 41260 1196
rect 41300 1156 41309 1196
rect 41251 1155 41309 1156
rect 2467 1112 2525 1113
rect 2467 1072 2476 1112
rect 2516 1072 2525 1112
rect 2467 1071 2525 1072
rect 3715 1112 3773 1113
rect 3715 1072 3724 1112
rect 3764 1072 3773 1112
rect 3715 1071 3773 1072
rect 4203 1112 4245 1121
rect 4203 1072 4204 1112
rect 4244 1072 4245 1112
rect 4203 1063 4245 1072
rect 4299 1112 4341 1121
rect 4299 1072 4300 1112
rect 4340 1072 4341 1112
rect 4299 1063 4341 1072
rect 4395 1112 4437 1121
rect 4395 1072 4396 1112
rect 4436 1072 4437 1112
rect 4395 1063 4437 1072
rect 4491 1112 4533 1121
rect 4491 1072 4492 1112
rect 4532 1072 4533 1112
rect 4491 1063 4533 1072
rect 4683 1112 4725 1121
rect 4683 1072 4684 1112
rect 4724 1072 4725 1112
rect 4683 1063 4725 1072
rect 4779 1112 4821 1121
rect 4779 1072 4780 1112
rect 4820 1072 4821 1112
rect 4779 1063 4821 1072
rect 4875 1112 4917 1121
rect 4875 1072 4876 1112
rect 4916 1072 4917 1112
rect 4875 1063 4917 1072
rect 6499 1112 6557 1113
rect 6499 1072 6508 1112
rect 6548 1072 6557 1112
rect 6499 1071 6557 1072
rect 7747 1112 7805 1113
rect 7747 1072 7756 1112
rect 7796 1072 7805 1112
rect 7747 1071 7805 1072
rect 8131 1112 8189 1113
rect 8131 1072 8140 1112
rect 8180 1072 8189 1112
rect 8131 1071 8189 1072
rect 9379 1112 9437 1113
rect 9379 1072 9388 1112
rect 9428 1072 9437 1112
rect 9379 1071 9437 1072
rect 9763 1112 9821 1113
rect 9763 1072 9772 1112
rect 9812 1072 9821 1112
rect 9763 1071 9821 1072
rect 11011 1112 11069 1113
rect 11011 1072 11020 1112
rect 11060 1072 11069 1112
rect 11011 1071 11069 1072
rect 11395 1112 11453 1113
rect 11395 1072 11404 1112
rect 11444 1072 11453 1112
rect 11395 1071 11453 1072
rect 12643 1112 12701 1113
rect 12643 1072 12652 1112
rect 12692 1072 12701 1112
rect 12643 1071 12701 1072
rect 13027 1112 13085 1113
rect 13027 1072 13036 1112
rect 13076 1072 13085 1112
rect 13027 1071 13085 1072
rect 14275 1112 14333 1113
rect 14275 1072 14284 1112
rect 14324 1072 14333 1112
rect 14275 1071 14333 1072
rect 16291 1112 16349 1113
rect 16291 1072 16300 1112
rect 16340 1072 16349 1112
rect 16291 1071 16349 1072
rect 17539 1112 17597 1113
rect 17539 1072 17548 1112
rect 17588 1072 17597 1112
rect 17539 1071 17597 1072
rect 18403 1112 18461 1113
rect 18403 1072 18412 1112
rect 18452 1072 18461 1112
rect 18403 1071 18461 1072
rect 19651 1112 19709 1113
rect 19651 1072 19660 1112
rect 19700 1072 19709 1112
rect 19651 1071 19709 1072
rect 20035 1112 20093 1113
rect 20035 1072 20044 1112
rect 20084 1072 20093 1112
rect 20035 1071 20093 1072
rect 21283 1112 21341 1113
rect 21283 1072 21292 1112
rect 21332 1072 21341 1112
rect 21283 1071 21341 1072
rect 21667 1112 21725 1113
rect 21667 1072 21676 1112
rect 21716 1072 21725 1112
rect 21667 1071 21725 1072
rect 22915 1112 22973 1113
rect 22915 1072 22924 1112
rect 22964 1072 22973 1112
rect 22915 1071 22973 1072
rect 23683 1112 23741 1113
rect 23683 1072 23692 1112
rect 23732 1072 23741 1112
rect 23683 1071 23741 1072
rect 24931 1112 24989 1113
rect 24931 1072 24940 1112
rect 24980 1072 24989 1112
rect 24931 1071 24989 1072
rect 25411 1112 25469 1113
rect 25411 1072 25420 1112
rect 25460 1072 25469 1112
rect 25411 1071 25469 1072
rect 26659 1112 26717 1113
rect 26659 1072 26668 1112
rect 26708 1072 26717 1112
rect 26659 1071 26717 1072
rect 27619 1112 27677 1113
rect 27619 1072 27628 1112
rect 27668 1072 27677 1112
rect 27619 1071 27677 1072
rect 28867 1112 28925 1113
rect 28867 1072 28876 1112
rect 28916 1072 28925 1112
rect 28867 1071 28925 1072
rect 29923 1112 29981 1113
rect 29923 1072 29932 1112
rect 29972 1072 29981 1112
rect 29923 1071 29981 1072
rect 30883 1112 30941 1113
rect 30883 1072 30892 1112
rect 30932 1072 30941 1112
rect 30883 1071 30941 1072
rect 31171 1112 31229 1113
rect 31171 1072 31180 1112
rect 31220 1072 31229 1112
rect 31171 1071 31229 1072
rect 35587 1112 35645 1113
rect 35587 1072 35596 1112
rect 35636 1072 35645 1112
rect 35587 1071 35645 1072
rect 36835 1112 36893 1113
rect 36835 1072 36844 1112
rect 36884 1072 36893 1112
rect 36835 1071 36893 1072
rect 3915 1028 3957 1037
rect 3915 988 3916 1028
rect 3956 988 3957 1028
rect 3915 979 3957 988
rect 4963 944 5021 945
rect 4963 904 4972 944
rect 5012 904 5021 944
rect 4963 903 5021 904
rect 7947 944 7989 953
rect 7947 904 7948 944
rect 7988 904 7989 944
rect 7947 895 7989 904
rect 12843 944 12885 953
rect 12843 904 12844 944
rect 12884 904 12885 944
rect 12843 895 12885 904
rect 32331 944 32373 953
rect 32331 904 32332 944
rect 32372 904 32373 944
rect 32331 895 32373 904
rect 34251 944 34293 953
rect 34251 904 34252 944
rect 34292 904 34293 944
rect 34251 895 34293 904
rect 34635 944 34677 953
rect 34635 904 34636 944
rect 34676 904 34677 944
rect 34635 895 34677 904
rect 35019 944 35061 953
rect 35019 904 35020 944
rect 35060 904 35061 944
rect 35019 895 35061 904
rect 40683 944 40725 953
rect 40683 904 40684 944
rect 40724 904 40725 944
rect 40683 895 40725 904
rect 41067 944 41109 953
rect 41067 904 41068 944
rect 41108 904 41109 944
rect 41067 895 41109 904
rect 41451 944 41493 953
rect 41451 904 41452 944
rect 41492 904 41493 944
rect 41451 895 41493 904
rect 1152 776 41856 800
rect 1152 736 4928 776
rect 4968 736 5010 776
rect 5050 736 5092 776
rect 5132 736 5174 776
rect 5214 736 5256 776
rect 5296 736 20048 776
rect 20088 736 20130 776
rect 20170 736 20212 776
rect 20252 736 20294 776
rect 20334 736 20376 776
rect 20416 736 35168 776
rect 35208 736 35250 776
rect 35290 736 35332 776
rect 35372 736 35414 776
rect 35454 736 35496 776
rect 35536 736 41856 776
rect 1152 712 41856 736
<< via1 >>
rect 4928 9808 4968 9848
rect 5010 9808 5050 9848
rect 5092 9808 5132 9848
rect 5174 9808 5214 9848
rect 5256 9808 5296 9848
rect 20048 9808 20088 9848
rect 20130 9808 20170 9848
rect 20212 9808 20252 9848
rect 20294 9808 20334 9848
rect 20376 9808 20416 9848
rect 35168 9808 35208 9848
rect 35250 9808 35290 9848
rect 35332 9808 35372 9848
rect 35414 9808 35454 9848
rect 35496 9808 35536 9848
rect 4012 9640 4052 9680
rect 5740 9640 5780 9680
rect 9004 9640 9044 9680
rect 10156 9640 10196 9680
rect 10732 9640 10772 9680
rect 14188 9640 14228 9680
rect 17068 9640 17108 9680
rect 18988 9640 19028 9680
rect 22252 9640 22292 9680
rect 29836 9640 29876 9680
rect 30028 9640 30068 9680
rect 30412 9640 30452 9680
rect 30796 9640 30836 9680
rect 41452 9640 41492 9680
rect 3532 9556 3572 9596
rect 1900 9472 1940 9512
rect 3148 9472 3188 9512
rect 3628 9472 3668 9512
rect 3724 9472 3764 9512
rect 3820 9472 3860 9512
rect 4204 9472 4244 9512
rect 4300 9472 4340 9512
rect 4492 9472 4532 9512
rect 4588 9472 4628 9512
rect 4780 9472 4820 9512
rect 4876 9472 4916 9512
rect 5033 9457 5073 9497
rect 5260 9472 5300 9512
rect 5356 9472 5396 9512
rect 5452 9472 5492 9512
rect 5548 9472 5588 9512
rect 5836 9472 5876 9512
rect 5932 9472 5972 9512
rect 6028 9472 6068 9512
rect 6220 9472 6260 9512
rect 6412 9472 6452 9512
rect 6892 9472 6932 9512
rect 6988 9472 7028 9512
rect 7276 9472 7316 9512
rect 7564 9472 7604 9512
rect 8812 9472 8852 9512
rect 9484 9472 9524 9512
rect 9580 9472 9620 9512
rect 9868 9472 9908 9512
rect 10924 9472 10964 9512
rect 12172 9472 12212 9512
rect 14956 9472 14996 9512
rect 16204 9472 16244 9512
rect 19180 9472 19220 9512
rect 20428 9472 20468 9512
rect 22732 9472 22772 9512
rect 23980 9472 24020 9512
rect 24364 9472 24404 9512
rect 25612 9472 25652 9512
rect 27148 9472 27188 9512
rect 28396 9472 28436 9512
rect 31180 9472 31220 9512
rect 32428 9472 32468 9512
rect 32908 9472 32948 9512
rect 34156 9472 34196 9512
rect 35020 9472 35060 9512
rect 36268 9472 36308 9512
rect 38476 9472 38516 9512
rect 39724 9472 39764 9512
rect 10348 9388 10388 9428
rect 10540 9388 10580 9428
rect 14380 9388 14420 9428
rect 16876 9388 16916 9428
rect 18796 9388 18836 9428
rect 22444 9388 22484 9428
rect 29644 9388 29684 9428
rect 30220 9388 30260 9428
rect 30604 9388 30644 9428
rect 30988 9388 31028 9428
rect 37228 9388 37268 9428
rect 37804 9388 37844 9428
rect 40876 9388 40916 9428
rect 41260 9388 41300 9428
rect 3340 9304 3380 9344
rect 41068 9304 41108 9344
rect 4492 9220 4532 9260
rect 6316 9220 6356 9260
rect 6604 9220 6644 9260
rect 9196 9220 9236 9260
rect 12364 9220 12404 9260
rect 16396 9220 16436 9260
rect 20620 9220 20660 9260
rect 24172 9220 24212 9260
rect 25804 9220 25844 9260
rect 26956 9220 26996 9260
rect 32620 9220 32660 9260
rect 34348 9220 34388 9260
rect 36460 9220 36500 9260
rect 37036 9220 37076 9260
rect 37612 9220 37652 9260
rect 38284 9220 38324 9260
rect 3688 9052 3728 9092
rect 3770 9052 3810 9092
rect 3852 9052 3892 9092
rect 3934 9052 3974 9092
rect 4016 9052 4056 9092
rect 18808 9052 18848 9092
rect 18890 9052 18930 9092
rect 18972 9052 19012 9092
rect 19054 9052 19094 9092
rect 19136 9052 19176 9092
rect 33928 9052 33968 9092
rect 34010 9052 34050 9092
rect 34092 9052 34132 9092
rect 34174 9052 34214 9092
rect 34256 9052 34296 9092
rect 3532 8884 3572 8924
rect 5164 8884 5204 8924
rect 1708 8800 1748 8840
rect 1900 8800 1940 8840
rect 8620 8800 8660 8840
rect 18412 8800 18452 8840
rect 24556 8800 24596 8840
rect 25036 8800 25076 8840
rect 25516 8800 25556 8840
rect 34348 8800 34388 8840
rect 40300 8800 40340 8840
rect 40684 8800 40724 8840
rect 41452 8800 41492 8840
rect 8428 8716 8468 8756
rect 3340 8674 3380 8714
rect 1708 8632 1748 8672
rect 2092 8632 2132 8672
rect 3724 8632 3764 8672
rect 4972 8632 5012 8672
rect 5452 8632 5492 8672
rect 5548 8632 5588 8672
rect 6124 8632 6164 8672
rect 6220 8632 6260 8672
rect 6604 8632 6644 8672
rect 6700 8632 6740 8672
rect 7180 8632 7220 8672
rect 7660 8646 7700 8686
rect 8812 8632 8852 8672
rect 10060 8632 10100 8672
rect 10828 8632 10868 8672
rect 10924 8632 10964 8672
rect 11308 8632 11348 8672
rect 11404 8674 11444 8714
rect 11884 8632 11924 8672
rect 12364 8646 12404 8686
rect 13036 8632 13076 8672
rect 14284 8632 14324 8672
rect 14764 8632 14804 8672
rect 14860 8632 14900 8672
rect 15244 8632 15284 8672
rect 15340 8632 15380 8672
rect 15820 8632 15860 8672
rect 16300 8646 16340 8686
rect 16972 8632 17012 8672
rect 18220 8632 18260 8672
rect 18700 8632 18740 8672
rect 18796 8632 18836 8672
rect 19180 8632 19220 8672
rect 20284 8674 20324 8714
rect 22924 8716 22964 8756
rect 23020 8716 23060 8756
rect 24748 8716 24788 8756
rect 25228 8716 25268 8756
rect 25708 8716 25748 8756
rect 26476 8716 26516 8756
rect 19276 8632 19316 8672
rect 19756 8632 19796 8672
rect 20716 8632 20756 8672
rect 21964 8632 22004 8672
rect 22444 8632 22484 8672
rect 24028 8674 24068 8714
rect 26572 8716 26612 8756
rect 28108 8716 28148 8756
rect 29548 8716 29588 8756
rect 29644 8716 29684 8756
rect 31180 8716 31220 8756
rect 31564 8716 31604 8756
rect 31948 8716 31988 8756
rect 32812 8716 32852 8756
rect 36268 8716 36308 8756
rect 39916 8716 39956 8756
rect 40108 8716 40148 8756
rect 40492 8716 40532 8756
rect 40876 8716 40916 8756
rect 41260 8716 41300 8756
rect 22540 8632 22580 8672
rect 23500 8632 23540 8672
rect 25996 8632 26036 8672
rect 26092 8632 26132 8672
rect 27052 8632 27092 8672
rect 27532 8646 27572 8686
rect 29068 8632 29108 8672
rect 29164 8632 29204 8672
rect 30124 8632 30164 8672
rect 30604 8646 30644 8686
rect 32332 8632 32372 8672
rect 32428 8632 32468 8672
rect 32908 8632 32948 8672
rect 33388 8632 33428 8672
rect 33868 8646 33908 8686
rect 34636 8632 34676 8672
rect 34732 8632 34772 8672
rect 35020 8632 35060 8672
rect 35692 8632 35732 8672
rect 35788 8632 35828 8672
rect 36172 8632 36212 8672
rect 36748 8632 36788 8672
rect 37228 8637 37268 8677
rect 37804 8632 37844 8672
rect 39052 8632 39092 8672
rect 7852 8548 7892 8588
rect 10252 8548 10292 8588
rect 14476 8548 14516 8588
rect 16492 8548 16532 8588
rect 22156 8548 22196 8588
rect 24172 8548 24212 8588
rect 37420 8548 37460 8588
rect 3532 8464 3572 8504
rect 5740 8464 5780 8504
rect 12556 8464 12596 8504
rect 20428 8464 20468 8504
rect 27724 8464 27764 8504
rect 27916 8464 27956 8504
rect 30796 8422 30836 8462
rect 30988 8464 31028 8504
rect 31372 8464 31412 8504
rect 31756 8464 31796 8504
rect 34060 8464 34100 8504
rect 37612 8464 37652 8504
rect 39724 8464 39764 8504
rect 41068 8464 41108 8504
rect 4928 8296 4968 8336
rect 5010 8296 5050 8336
rect 5092 8296 5132 8336
rect 5174 8296 5214 8336
rect 5256 8296 5296 8336
rect 20048 8296 20088 8336
rect 20130 8296 20170 8336
rect 20212 8296 20252 8336
rect 20294 8296 20334 8336
rect 20376 8296 20416 8336
rect 35168 8296 35208 8336
rect 35250 8296 35290 8336
rect 35332 8296 35372 8336
rect 35414 8296 35454 8336
rect 35496 8296 35536 8336
rect 3340 8128 3380 8168
rect 3820 8128 3860 8168
rect 7660 8128 7700 8168
rect 9580 8128 9620 8168
rect 11500 8128 11540 8168
rect 11884 8128 11924 8168
rect 17068 8128 17108 8168
rect 19276 8170 19316 8210
rect 19468 8128 19508 8168
rect 20044 8128 20084 8168
rect 22732 8128 22772 8168
rect 22924 8128 22964 8168
rect 27532 8128 27572 8168
rect 29452 8128 29492 8168
rect 31180 8128 31220 8168
rect 32236 8128 32276 8168
rect 34732 8128 34772 8168
rect 37996 8128 38036 8168
rect 40012 8128 40052 8168
rect 40684 8128 40724 8168
rect 41452 8128 41492 8168
rect 14188 8044 14228 8084
rect 16300 8044 16340 8084
rect 1900 7960 1940 8000
rect 3148 7960 3188 8000
rect 3724 7960 3764 8000
rect 3916 7960 3956 8000
rect 4012 7960 4052 8000
rect 4300 7967 4340 8007
rect 4588 7960 4628 8000
rect 4684 7960 4724 8000
rect 5356 7960 5396 8000
rect 5452 7960 5492 8000
rect 5548 7960 5588 8000
rect 5644 7960 5684 8000
rect 5932 7960 5972 8000
rect 6028 7960 6068 8000
rect 6412 7960 6452 8000
rect 6988 7960 7028 8000
rect 7468 7955 7508 7995
rect 9772 7960 9812 8000
rect 11020 7960 11060 8000
rect 12748 7960 12788 8000
rect 13996 7960 14036 8000
rect 14572 7960 14612 8000
rect 14668 7960 14708 8000
rect 15148 7960 15188 8000
rect 6508 7876 6548 7916
rect 9388 7876 9428 7916
rect 11692 7876 11732 7916
rect 12076 7876 12116 7916
rect 15628 7918 15668 7958
rect 16108 7946 16148 7986
rect 17548 7960 17588 8000
rect 17644 7960 17684 8000
rect 18124 7960 18164 8000
rect 18604 7960 18644 8000
rect 15052 7876 15092 7916
rect 16876 7876 16916 7916
rect 18028 7876 18068 7916
rect 19132 7918 19172 7958
rect 21004 7960 21044 8000
rect 21100 7960 21140 8000
rect 21580 7960 21620 8000
rect 22060 7960 22100 8000
rect 24076 7960 24116 8000
rect 25324 7960 25364 8000
rect 25804 7960 25844 8000
rect 20236 7876 20276 7916
rect 21484 7876 21524 7916
rect 22588 7918 22628 7958
rect 25900 7960 25940 8000
rect 26284 7960 26324 8000
rect 26380 7960 26420 8000
rect 26860 7960 26900 8000
rect 28012 7960 28052 8000
rect 29260 7960 29300 8000
rect 29740 7960 29780 8000
rect 30988 7960 31028 8000
rect 33292 7960 33332 8000
rect 34540 7960 34580 8000
rect 36268 7960 36308 8000
rect 27388 7918 27428 7958
rect 36364 7960 36404 8000
rect 37324 7960 37364 8000
rect 37852 7950 37892 7990
rect 38284 7960 38324 8000
rect 38380 7960 38420 8000
rect 39340 7960 39380 8000
rect 39820 7946 39860 7986
rect 23116 7876 23156 7916
rect 31564 7876 31604 7916
rect 32428 7876 32468 7916
rect 32812 7876 32852 7916
rect 36748 7876 36788 7916
rect 36844 7876 36884 7916
rect 38764 7876 38804 7916
rect 38860 7876 38900 7916
rect 40492 7876 40532 7916
rect 40876 7876 40916 7916
rect 41260 7876 41300 7916
rect 4972 7792 5012 7832
rect 41068 7792 41108 7832
rect 11212 7708 11252 7748
rect 25516 7708 25556 7748
rect 31372 7708 31412 7748
rect 32620 7708 32660 7748
rect 3688 7540 3728 7580
rect 3770 7540 3810 7580
rect 3852 7540 3892 7580
rect 3934 7540 3974 7580
rect 4016 7540 4056 7580
rect 18808 7540 18848 7580
rect 18890 7540 18930 7580
rect 18972 7540 19012 7580
rect 19054 7540 19094 7580
rect 19136 7540 19176 7580
rect 33928 7540 33968 7580
rect 34010 7540 34050 7580
rect 34092 7540 34132 7580
rect 34174 7540 34214 7580
rect 34256 7540 34296 7580
rect 3628 7372 3668 7412
rect 4396 7372 4436 7412
rect 11692 7372 11732 7412
rect 12940 7372 12980 7412
rect 13708 7372 13748 7412
rect 15820 7372 15860 7412
rect 17452 7372 17492 7412
rect 19084 7372 19124 7412
rect 21100 7372 21140 7412
rect 22828 7372 22868 7412
rect 27532 7372 27572 7412
rect 35980 7372 36020 7412
rect 37708 7372 37748 7412
rect 40396 7372 40436 7412
rect 41452 7372 41492 7412
rect 10252 7204 10292 7244
rect 11884 7204 11924 7244
rect 12748 7204 12788 7244
rect 13900 7204 13940 7244
rect 33868 7204 33908 7244
rect 40876 7204 40916 7244
rect 41260 7204 41300 7244
rect 1708 7120 1748 7160
rect 2956 7120 2996 7160
rect 3628 7120 3668 7160
rect 3820 7120 3860 7160
rect 3916 7120 3956 7160
rect 4108 7120 4148 7160
rect 4396 7120 4436 7160
rect 4588 7120 4628 7160
rect 5836 7120 5876 7160
rect 6412 7120 6452 7160
rect 6508 7120 6548 7160
rect 8044 7120 8084 7160
rect 9292 7120 9332 7160
rect 9772 7120 9812 7160
rect 9868 7120 9908 7160
rect 11356 7162 11396 7202
rect 10348 7120 10388 7160
rect 10828 7120 10868 7160
rect 14380 7120 14420 7160
rect 15628 7120 15668 7160
rect 16012 7120 16052 7160
rect 17260 7120 17300 7160
rect 17644 7120 17684 7160
rect 18892 7120 18932 7160
rect 19660 7120 19700 7160
rect 20908 7120 20948 7160
rect 21388 7120 21428 7160
rect 22636 7120 22676 7160
rect 24364 7120 24404 7160
rect 25612 7120 25652 7160
rect 26092 7120 26132 7160
rect 27340 7120 27380 7160
rect 27724 7120 27764 7160
rect 28972 7120 29012 7160
rect 30220 7120 30260 7160
rect 31468 7120 31508 7160
rect 31948 7120 31988 7160
rect 33196 7120 33236 7160
rect 34540 7120 34580 7160
rect 35788 7120 35828 7160
rect 36268 7120 36308 7160
rect 37516 7120 37556 7160
rect 38956 7120 38996 7160
rect 40204 7120 40244 7160
rect 9484 7036 9524 7076
rect 11500 7036 11540 7076
rect 3148 6952 3188 6992
rect 6028 6952 6068 6992
rect 6220 6952 6260 6992
rect 25804 6952 25844 6992
rect 29164 6952 29204 6992
rect 31660 6952 31700 6992
rect 33388 6952 33428 6992
rect 33676 6952 33716 6992
rect 41068 6952 41108 6992
rect 4928 6784 4968 6824
rect 5010 6784 5050 6824
rect 5092 6784 5132 6824
rect 5174 6784 5214 6824
rect 5256 6784 5296 6824
rect 20048 6784 20088 6824
rect 20130 6784 20170 6824
rect 20212 6784 20252 6824
rect 20294 6784 20334 6824
rect 20376 6784 20416 6824
rect 35168 6784 35208 6824
rect 35250 6784 35290 6824
rect 35332 6784 35372 6824
rect 35414 6784 35454 6824
rect 35496 6784 35536 6824
rect 7276 6616 7316 6656
rect 10348 6616 10388 6656
rect 14188 6616 14228 6656
rect 14668 6616 14708 6656
rect 19468 6616 19508 6656
rect 21292 6616 21332 6656
rect 23308 6616 23348 6656
rect 25708 6616 25748 6656
rect 30892 6616 30932 6656
rect 33196 6616 33236 6656
rect 37612 6616 37652 6656
rect 41452 6616 41492 6656
rect 4492 6532 4532 6572
rect 8908 6532 8948 6572
rect 12172 6532 12212 6572
rect 28876 6532 28916 6572
rect 40012 6532 40052 6572
rect 2764 6448 2804 6488
rect 4012 6448 4052 6488
rect 4684 6434 4724 6474
rect 5164 6448 5204 6488
rect 6124 6448 6164 6488
rect 6220 6448 6260 6488
rect 6508 6448 6548 6488
rect 6604 6448 6644 6488
rect 6700 6448 6740 6488
rect 6796 6448 6836 6488
rect 6988 6448 7028 6488
rect 7084 6448 7124 6488
rect 7180 6448 7220 6488
rect 7468 6448 7508 6488
rect 8716 6448 8756 6488
rect 9196 6448 9236 6488
rect 9484 6448 9524 6488
rect 9580 6448 9620 6488
rect 10732 6448 10772 6488
rect 11980 6448 12020 6488
rect 12460 6448 12500 6488
rect 12556 6448 12596 6488
rect 12940 6448 12980 6488
rect 13516 6448 13556 6488
rect 13996 6434 14036 6474
rect 15340 6448 15380 6488
rect 15916 6448 15956 6488
rect 5644 6364 5684 6404
rect 5740 6364 5780 6404
rect 10540 6364 10580 6404
rect 13036 6364 13076 6404
rect 14812 6406 14852 6446
rect 16300 6448 16340 6488
rect 16396 6448 16436 6488
rect 17644 6448 17684 6488
rect 18892 6448 18932 6488
rect 19852 6448 19892 6488
rect 21100 6448 21140 6488
rect 21580 6448 21620 6488
rect 21676 6448 21716 6488
rect 22060 6448 22100 6488
rect 22156 6448 22196 6488
rect 22636 6448 22676 6488
rect 23116 6434 23156 6474
rect 23980 6448 24020 6488
rect 24076 6448 24116 6488
rect 24460 6448 24500 6488
rect 24556 6448 24596 6488
rect 25036 6448 25076 6488
rect 25516 6443 25556 6483
rect 27148 6448 27188 6488
rect 27244 6448 27284 6488
rect 27628 6448 27668 6488
rect 27724 6448 27764 6488
rect 28204 6448 28244 6488
rect 28684 6443 28724 6483
rect 29164 6448 29204 6488
rect 29260 6448 29300 6488
rect 29644 6448 29684 6488
rect 29740 6448 29780 6488
rect 30220 6448 30260 6488
rect 30700 6434 30740 6474
rect 31468 6448 31508 6488
rect 31564 6448 31604 6488
rect 31948 6448 31988 6488
rect 32524 6448 32564 6488
rect 33388 6448 33428 6488
rect 34636 6448 34676 6488
rect 38284 6448 38324 6488
rect 15820 6364 15860 6404
rect 19660 6364 19700 6404
rect 32044 6364 32084 6404
rect 33052 6406 33092 6446
rect 38380 6448 38420 6488
rect 38764 6448 38804 6488
rect 38860 6448 38900 6488
rect 39340 6448 39380 6488
rect 39820 6434 39860 6474
rect 35884 6364 35924 6404
rect 37804 6364 37844 6404
rect 40396 6364 40436 6404
rect 40876 6364 40916 6404
rect 41260 6364 41300 6404
rect 4204 6280 4244 6320
rect 9868 6280 9908 6320
rect 19084 6280 19124 6320
rect 35692 6280 35732 6320
rect 40204 6280 40244 6320
rect 41068 6280 41108 6320
rect 34828 6196 34868 6236
rect 3688 6028 3728 6068
rect 3770 6028 3810 6068
rect 3852 6028 3892 6068
rect 3934 6028 3974 6068
rect 4016 6028 4056 6068
rect 18808 6028 18848 6068
rect 18890 6028 18930 6068
rect 18972 6028 19012 6068
rect 19054 6028 19094 6068
rect 19136 6028 19176 6068
rect 33928 6028 33968 6068
rect 34010 6028 34050 6068
rect 34092 6028 34132 6068
rect 34174 6028 34214 6068
rect 34256 6028 34296 6068
rect 4684 5860 4724 5900
rect 10924 5860 10964 5900
rect 12844 5860 12884 5900
rect 14476 5860 14516 5900
rect 14668 5860 14708 5900
rect 22732 5860 22772 5900
rect 27244 5860 27284 5900
rect 40396 5860 40436 5900
rect 41068 5860 41108 5900
rect 4300 5776 4340 5816
rect 19948 5776 19988 5816
rect 24364 5776 24404 5816
rect 41452 5776 41492 5816
rect 11116 5692 11156 5732
rect 12652 5692 12692 5732
rect 28492 5692 28532 5732
rect 29356 5692 29396 5732
rect 29452 5692 29492 5732
rect 32044 5692 32084 5732
rect 32140 5692 32180 5732
rect 34828 5692 34868 5732
rect 36844 5692 36884 5732
rect 40876 5692 40916 5732
rect 41260 5692 41300 5732
rect 1612 5608 1652 5648
rect 2860 5608 2900 5648
rect 4300 5608 4340 5648
rect 4780 5608 4820 5648
rect 5164 5608 5204 5648
rect 5260 5608 5300 5648
rect 5740 5608 5780 5648
rect 5836 5608 5876 5648
rect 6220 5608 6260 5648
rect 6316 5608 6356 5648
rect 6796 5608 6836 5648
rect 7324 5617 7364 5657
rect 7660 5608 7700 5648
rect 8908 5608 8948 5648
rect 9292 5608 9332 5648
rect 10540 5608 10580 5648
rect 13036 5608 13076 5648
rect 14284 5608 14324 5648
rect 14860 5608 14900 5648
rect 16108 5608 16148 5648
rect 16300 5608 16340 5648
rect 17548 5608 17588 5648
rect 18028 5608 18068 5648
rect 18124 5608 18164 5648
rect 18508 5608 18548 5648
rect 18604 5608 18644 5648
rect 19084 5608 19124 5648
rect 19564 5613 19604 5653
rect 20332 5608 20372 5648
rect 20620 5608 20660 5648
rect 21292 5608 21332 5648
rect 22540 5608 22580 5648
rect 22924 5608 22964 5648
rect 24172 5608 24212 5648
rect 25804 5608 25844 5648
rect 27052 5608 27092 5648
rect 28876 5608 28916 5648
rect 28972 5608 29012 5648
rect 29932 5599 29972 5639
rect 30460 5617 30500 5657
rect 31564 5608 31604 5648
rect 31660 5608 31700 5648
rect 32620 5608 32660 5648
rect 33148 5617 33188 5657
rect 34348 5608 34388 5648
rect 34444 5608 34484 5648
rect 34924 5608 34964 5648
rect 35404 5608 35444 5648
rect 35884 5613 35924 5653
rect 36364 5608 36404 5648
rect 36460 5608 36500 5648
rect 36940 5608 36980 5648
rect 37420 5608 37460 5648
rect 37900 5613 37940 5653
rect 38956 5608 38996 5648
rect 40204 5608 40244 5648
rect 17740 5524 17780 5564
rect 19756 5524 19796 5564
rect 20236 5524 20276 5564
rect 30604 5524 30644 5564
rect 36076 5524 36116 5564
rect 38092 5524 38132 5564
rect 3052 5440 3092 5480
rect 4492 5440 4532 5480
rect 5452 5440 5492 5480
rect 7468 5440 7508 5480
rect 9100 5440 9140 5480
rect 10732 5440 10772 5480
rect 28300 5440 28340 5480
rect 33292 5440 33332 5480
rect 4928 5272 4968 5312
rect 5010 5272 5050 5312
rect 5092 5272 5132 5312
rect 5174 5272 5214 5312
rect 5256 5272 5296 5312
rect 20048 5272 20088 5312
rect 20130 5272 20170 5312
rect 20212 5272 20252 5312
rect 20294 5272 20334 5312
rect 20376 5272 20416 5312
rect 35168 5272 35208 5312
rect 35250 5272 35290 5312
rect 35332 5272 35372 5312
rect 35414 5272 35454 5312
rect 35496 5272 35536 5312
rect 3916 5104 3956 5144
rect 11212 5104 11252 5144
rect 19756 5104 19796 5144
rect 28876 5104 28916 5144
rect 33484 5104 33524 5144
rect 35788 5104 35828 5144
rect 5164 5020 5204 5060
rect 5740 5020 5780 5060
rect 7756 5020 7796 5060
rect 13900 5020 13940 5060
rect 23116 5020 23156 5060
rect 30892 5020 30932 5060
rect 38668 5020 38708 5060
rect 1708 4936 1748 4976
rect 2956 4936 2996 4976
rect 3628 4936 3668 4976
rect 3724 4936 3764 4976
rect 4108 4936 4148 4976
rect 4300 4936 4340 4976
rect 4396 4936 4436 4976
rect 4588 4936 4628 4976
rect 4876 4936 4916 4976
rect 5068 4936 5108 4976
rect 5260 4936 5300 4976
rect 5452 4936 5492 4976
rect 5548 4936 5588 4976
rect 5644 4936 5684 4976
rect 6028 4936 6068 4976
rect 6124 4936 6164 4976
rect 6508 4936 6548 4976
rect 6604 4936 6644 4976
rect 7084 4936 7124 4976
rect 7564 4922 7604 4962
rect 9484 4936 9524 4976
rect 9580 4936 9620 4976
rect 9964 4936 10004 4976
rect 10060 4936 10100 4976
rect 10540 4936 10580 4976
rect 11020 4931 11060 4971
rect 12460 4936 12500 4976
rect 13708 4936 13748 4976
rect 18316 4936 18356 4976
rect 19564 4936 19604 4976
rect 21388 4936 21428 4976
rect 21484 4936 21524 4976
rect 21964 4936 22004 4976
rect 22444 4936 22484 4976
rect 22972 4926 23012 4966
rect 23884 4936 23924 4976
rect 25132 4936 25172 4976
rect 27148 4936 27188 4976
rect 27244 4936 27284 4976
rect 27628 4936 27668 4976
rect 27724 4936 27764 4976
rect 28204 4936 28244 4976
rect 28732 4926 28772 4966
rect 29164 4917 29204 4957
rect 29260 4936 29300 4976
rect 29644 4936 29684 4976
rect 30220 4936 30260 4976
rect 30700 4922 30740 4962
rect 32044 4936 32084 4976
rect 33292 4936 33332 4976
rect 34348 4936 34388 4976
rect 35596 4936 35636 4976
rect 37228 4936 37268 4976
rect 38476 4936 38516 4976
rect 39052 4936 39092 4976
rect 40300 4936 40340 4976
rect 11692 4852 11732 4892
rect 12268 4852 12308 4892
rect 14860 4852 14900 4892
rect 16972 4852 17012 4892
rect 17164 4852 17204 4892
rect 21100 4852 21140 4892
rect 21868 4852 21908 4892
rect 29740 4852 29780 4892
rect 36844 4852 36884 4892
rect 40684 4852 40724 4892
rect 40876 4852 40916 4892
rect 41260 4852 41300 4892
rect 3148 4768 3188 4808
rect 11884 4768 11924 4808
rect 14668 4768 14708 4808
rect 16780 4768 16820 4808
rect 17356 4768 17396 4808
rect 20908 4768 20948 4808
rect 36652 4768 36692 4808
rect 41068 4768 41108 4808
rect 41452 4768 41492 4808
rect 4108 4684 4148 4724
rect 4876 4684 4916 4724
rect 12076 4684 12116 4724
rect 25324 4684 25364 4724
rect 38860 4684 38900 4724
rect 40492 4684 40532 4724
rect 3688 4516 3728 4556
rect 3770 4516 3810 4556
rect 3852 4516 3892 4556
rect 3934 4516 3974 4556
rect 4016 4516 4056 4556
rect 18808 4516 18848 4556
rect 18890 4516 18930 4556
rect 18972 4516 19012 4556
rect 19054 4516 19094 4556
rect 19136 4516 19176 4556
rect 33928 4516 33968 4556
rect 34010 4516 34050 4556
rect 34092 4516 34132 4556
rect 34174 4516 34214 4556
rect 34256 4516 34296 4556
rect 28972 4348 29012 4388
rect 32044 4348 32084 4388
rect 40684 4348 40724 4388
rect 41068 4348 41108 4388
rect 4780 4264 4820 4304
rect 29452 4264 29492 4304
rect 7372 4180 7412 4220
rect 7468 4180 7508 4220
rect 11404 4180 11444 4220
rect 11500 4180 11540 4220
rect 13708 4180 13748 4220
rect 20332 4180 20372 4220
rect 23884 4180 23924 4220
rect 23980 4180 24020 4220
rect 1612 4096 1652 4136
rect 2860 4096 2900 4136
rect 3532 4096 3572 4136
rect 3724 4096 3764 4136
rect 3820 4096 3860 4136
rect 4108 4096 4148 4136
rect 4396 4096 4436 4136
rect 4492 4096 4532 4136
rect 5068 4096 5108 4136
rect 5164 4096 5204 4136
rect 5260 4096 5300 4136
rect 5452 4096 5492 4136
rect 5548 4096 5588 4136
rect 5644 4096 5684 4136
rect 5932 4096 5972 4136
rect 6028 4096 6068 4136
rect 6124 4096 6164 4136
rect 6892 4096 6932 4136
rect 6988 4096 7028 4136
rect 7948 4096 7988 4136
rect 8428 4101 8468 4141
rect 10924 4096 10964 4136
rect 11020 4096 11060 4136
rect 11980 4096 12020 4136
rect 12460 4101 12500 4141
rect 13132 4096 13172 4136
rect 13228 4096 13268 4136
rect 13612 4096 13652 4136
rect 14188 4096 14228 4136
rect 14668 4101 14708 4141
rect 15436 4096 15476 4136
rect 15532 4096 15572 4136
rect 15916 4096 15956 4136
rect 16012 4096 16052 4136
rect 16492 4096 16532 4136
rect 16972 4101 17012 4141
rect 19852 4096 19892 4136
rect 19948 4096 19988 4136
rect 20428 4096 20468 4136
rect 20908 4096 20948 4136
rect 21388 4101 21428 4141
rect 23404 4096 23444 4136
rect 24988 4138 25028 4178
rect 25900 4180 25940 4220
rect 25996 4180 26036 4220
rect 34348 4180 34388 4220
rect 35404 4180 35444 4220
rect 37036 4180 37076 4220
rect 38380 4180 38420 4220
rect 38476 4180 38516 4220
rect 40492 4180 40532 4220
rect 40876 4180 40916 4220
rect 41260 4180 41300 4220
rect 23500 4096 23540 4136
rect 24460 4096 24500 4136
rect 25420 4096 25460 4136
rect 25516 4096 25556 4136
rect 26476 4096 26516 4136
rect 26956 4101 26996 4141
rect 27532 4096 27572 4136
rect 28780 4096 28820 4136
rect 30124 4096 30164 4136
rect 30604 4096 30644 4136
rect 31852 4096 31892 4136
rect 32524 4096 32564 4136
rect 33772 4096 33812 4136
rect 34924 4096 34964 4136
rect 35020 4096 35060 4136
rect 35500 4096 35540 4136
rect 35980 4096 36020 4136
rect 36508 4105 36548 4145
rect 37900 4096 37940 4136
rect 37996 4096 38036 4136
rect 38956 4096 38996 4136
rect 39436 4110 39476 4150
rect 12652 4012 12692 4052
rect 14860 4012 14900 4052
rect 17164 4012 17204 4052
rect 21580 4012 21620 4052
rect 25132 4012 25172 4052
rect 36652 4012 36692 4052
rect 39628 4012 39668 4052
rect 3052 3928 3092 3968
rect 3628 3928 3668 3968
rect 4972 3928 5012 3968
rect 5740 3928 5780 3968
rect 6220 3928 6260 3968
rect 8620 3928 8660 3968
rect 27148 3928 27188 3968
rect 33964 3928 34004 3968
rect 34156 3928 34196 3968
rect 36844 3928 36884 3968
rect 41452 3928 41492 3968
rect 4928 3760 4968 3800
rect 5010 3760 5050 3800
rect 5092 3760 5132 3800
rect 5174 3760 5214 3800
rect 5256 3760 5296 3800
rect 20048 3760 20088 3800
rect 20130 3760 20170 3800
rect 20212 3760 20252 3800
rect 20294 3760 20334 3800
rect 20376 3760 20416 3800
rect 35168 3760 35208 3800
rect 35250 3760 35290 3800
rect 35332 3760 35372 3800
rect 35414 3760 35454 3800
rect 35496 3760 35536 3800
rect 4588 3592 4628 3632
rect 4876 3592 4916 3632
rect 11500 3592 11540 3632
rect 13708 3592 13748 3632
rect 15340 3592 15380 3632
rect 16972 3592 17012 3632
rect 17740 3592 17780 3632
rect 17932 3592 17972 3632
rect 19756 3592 19796 3632
rect 21484 3592 21524 3632
rect 27340 3592 27380 3632
rect 30796 3592 30836 3632
rect 31564 3592 31604 3632
rect 34348 3592 34388 3632
rect 37036 3592 37076 3632
rect 37324 3592 37364 3632
rect 41068 3592 41108 3632
rect 3052 3508 3092 3548
rect 6988 3508 7028 3548
rect 24460 3508 24500 3548
rect 1612 3424 1652 3464
rect 2860 3424 2900 3464
rect 3628 3424 3668 3464
rect 3724 3424 3764 3464
rect 3820 3424 3860 3464
rect 3916 3424 3956 3464
rect 4108 3424 4148 3464
rect 4204 3424 4244 3464
rect 4396 3424 4436 3464
rect 4492 3424 4532 3464
rect 4647 3424 4687 3464
rect 5068 3424 5108 3464
rect 5164 3424 5204 3464
rect 7084 3424 7124 3464
rect 7372 3424 7412 3464
rect 9772 3424 9812 3464
rect 9868 3424 9908 3464
rect 10252 3424 10292 3464
rect 10348 3424 10388 3464
rect 10828 3424 10868 3464
rect 11308 3410 11348 3450
rect 12268 3424 12308 3464
rect 13516 3424 13556 3464
rect 13900 3424 13940 3464
rect 15148 3424 15188 3464
rect 15532 3424 15572 3464
rect 16780 3424 16820 3464
rect 18316 3424 18356 3464
rect 19564 3424 19604 3464
rect 20044 3424 20084 3464
rect 21292 3424 21332 3464
rect 22732 3424 22772 3464
rect 22828 3424 22868 3464
rect 23212 3424 23252 3464
rect 23308 3424 23348 3464
rect 23788 3424 23828 3464
rect 24316 3382 24356 3422
rect 24844 3424 24884 3464
rect 25708 3424 25748 3464
rect 25900 3424 25940 3464
rect 27148 3424 27188 3464
rect 27628 3424 27668 3464
rect 28588 3424 28628 3464
rect 29356 3424 29396 3464
rect 30604 3424 30644 3464
rect 32620 3424 32660 3464
rect 32716 3424 32756 3464
rect 33100 3424 33140 3464
rect 33196 3424 33236 3464
rect 33676 3424 33716 3464
rect 34156 3419 34196 3459
rect 35308 3424 35348 3464
rect 35404 3424 35444 3464
rect 35788 3424 35828 3464
rect 35884 3424 35924 3464
rect 36364 3424 36404 3464
rect 37516 3424 37556 3464
rect 38764 3424 38804 3464
rect 17548 3340 17588 3380
rect 18124 3340 18164 3380
rect 36892 3382 36932 3422
rect 28972 3340 29012 3380
rect 31372 3340 31412 3380
rect 31756 3340 31796 3380
rect 40492 3340 40532 3380
rect 40876 3340 40916 3380
rect 6700 3256 6740 3296
rect 31180 3256 31220 3296
rect 40684 3256 40724 3296
rect 27916 3172 27956 3212
rect 28780 3172 28820 3212
rect 3688 3004 3728 3044
rect 3770 3004 3810 3044
rect 3852 3004 3892 3044
rect 3934 3004 3974 3044
rect 4016 3004 4056 3044
rect 18808 3004 18848 3044
rect 18890 3004 18930 3044
rect 18972 3004 19012 3044
rect 19054 3004 19094 3044
rect 19136 3004 19176 3044
rect 33928 3004 33968 3044
rect 34010 3004 34050 3044
rect 34092 3004 34132 3044
rect 34174 3004 34214 3044
rect 34256 3004 34296 3044
rect 7948 2836 7988 2876
rect 10540 2836 10580 2876
rect 12460 2836 12500 2876
rect 12844 2836 12884 2876
rect 23500 2836 23540 2876
rect 28972 2836 29012 2876
rect 31084 2836 31124 2876
rect 32908 2836 32948 2876
rect 35116 2836 35156 2876
rect 36940 2836 36980 2876
rect 38572 2836 38612 2876
rect 41068 2836 41108 2876
rect 19468 2752 19508 2792
rect 40684 2752 40724 2792
rect 13036 2668 13076 2708
rect 16588 2668 16628 2708
rect 16684 2668 16724 2708
rect 20812 2668 20852 2708
rect 20908 2668 20948 2708
rect 25996 2668 26036 2708
rect 26092 2668 26132 2708
rect 40492 2668 40532 2708
rect 40876 2668 40916 2708
rect 41260 2668 41300 2708
rect 1804 2584 1844 2624
rect 3052 2584 3092 2624
rect 3436 2584 3476 2624
rect 3532 2584 3572 2624
rect 3724 2584 3764 2624
rect 3820 2584 3860 2624
rect 4012 2584 4052 2624
rect 4300 2584 4340 2624
rect 4396 2584 4436 2624
rect 4492 2584 4532 2624
rect 4876 2584 4916 2624
rect 4972 2584 5012 2624
rect 5452 2584 5492 2624
rect 5548 2584 5588 2624
rect 5644 2584 5684 2624
rect 6508 2584 6548 2624
rect 7756 2584 7796 2624
rect 9100 2584 9140 2624
rect 10348 2584 10388 2624
rect 11020 2584 11060 2624
rect 12268 2584 12308 2624
rect 14380 2584 14420 2624
rect 15628 2584 15668 2624
rect 16108 2584 16148 2624
rect 16204 2584 16244 2624
rect 17164 2584 17204 2624
rect 17692 2593 17732 2633
rect 18028 2584 18068 2624
rect 19276 2584 19316 2624
rect 19852 2589 19892 2629
rect 20332 2584 20372 2624
rect 21292 2584 21332 2624
rect 21388 2584 21428 2624
rect 22060 2584 22100 2624
rect 23308 2584 23348 2624
rect 23692 2584 23732 2624
rect 24652 2584 24692 2624
rect 25516 2584 25556 2624
rect 25612 2584 25652 2624
rect 26572 2584 26612 2624
rect 27100 2593 27140 2633
rect 27532 2584 27572 2624
rect 28780 2584 28820 2624
rect 29644 2584 29684 2624
rect 30892 2584 30932 2624
rect 32716 2584 32756 2624
rect 33676 2584 33716 2624
rect 34924 2584 34964 2624
rect 35500 2584 35540 2624
rect 36748 2584 36788 2624
rect 37132 2584 37172 2624
rect 38380 2584 38420 2624
rect 3244 2500 3284 2540
rect 15820 2500 15860 2540
rect 17836 2500 17876 2540
rect 19660 2500 19700 2540
rect 31468 2542 31508 2582
rect 27244 2500 27284 2540
rect 4012 2416 4052 2456
rect 4684 2416 4724 2456
rect 5164 2416 5204 2456
rect 5356 2416 5396 2456
rect 41452 2416 41492 2456
rect 4928 2248 4968 2288
rect 5010 2248 5050 2288
rect 5092 2248 5132 2288
rect 5174 2248 5214 2288
rect 5256 2248 5296 2288
rect 20048 2248 20088 2288
rect 20130 2248 20170 2288
rect 20212 2248 20252 2288
rect 20294 2248 20334 2288
rect 20376 2248 20416 2288
rect 35168 2248 35208 2288
rect 35250 2248 35290 2288
rect 35332 2248 35372 2288
rect 35414 2248 35454 2288
rect 35496 2248 35536 2288
rect 4396 2080 4436 2120
rect 6700 2080 6740 2120
rect 19564 2080 19604 2120
rect 22732 2080 22772 2120
rect 24364 2080 24404 2120
rect 25996 2080 26036 2120
rect 29356 2080 29396 2120
rect 30988 2080 31028 2120
rect 31180 2080 31220 2120
rect 31564 2080 31604 2120
rect 32236 2080 32276 2120
rect 34828 2080 34868 2120
rect 36460 2080 36500 2120
rect 39244 2080 39284 2120
rect 40396 2080 40436 2120
rect 41068 2080 41108 2120
rect 4492 1996 4532 2036
rect 17164 1996 17204 2036
rect 34636 1996 34676 2036
rect 1900 1912 1940 1952
rect 3148 1912 3188 1952
rect 3820 1912 3860 1952
rect 3916 1912 3956 1952
rect 4012 1912 4052 1952
rect 4108 1912 4148 1952
rect 4588 1912 4628 1952
rect 4684 1912 4724 1952
rect 4876 1912 4916 1952
rect 5068 1912 5108 1952
rect 5260 1912 5300 1952
rect 6508 1912 6548 1952
rect 7276 1912 7316 1952
rect 8524 1912 8564 1952
rect 8908 1912 8948 1952
rect 10156 1912 10196 1952
rect 10540 1912 10580 1952
rect 11788 1912 11828 1952
rect 12172 1912 12212 1952
rect 13420 1912 13460 1952
rect 13804 1912 13844 1952
rect 15052 1912 15092 1952
rect 15436 1912 15476 1952
rect 16684 1912 16724 1952
rect 17548 1912 17588 1952
rect 18412 1912 18452 1952
rect 21292 1912 21332 1952
rect 22540 1912 22580 1952
rect 22924 1912 22964 1952
rect 24172 1912 24212 1952
rect 24556 1912 24596 1952
rect 25804 1912 25844 1952
rect 26188 1912 26228 1952
rect 27436 1912 27476 1952
rect 27916 1912 27956 1952
rect 29164 1912 29204 1952
rect 29548 1912 29588 1952
rect 30796 1912 30836 1952
rect 33388 1912 33428 1952
rect 34252 1912 34292 1952
rect 35020 1912 35060 1952
rect 36268 1912 36308 1952
rect 36652 1912 36692 1952
rect 37900 1912 37940 1952
rect 31372 1828 31412 1868
rect 31756 1828 31796 1868
rect 38380 1828 38420 1868
rect 39436 1828 39476 1868
rect 39628 1828 39668 1868
rect 40012 1828 40052 1868
rect 40588 1828 40628 1868
rect 40876 1828 40916 1868
rect 41260 1828 41300 1868
rect 4972 1744 5012 1784
rect 41452 1744 41492 1784
rect 3340 1660 3380 1700
rect 4588 1660 4628 1700
rect 8716 1660 8756 1700
rect 10348 1660 10388 1700
rect 11980 1660 12020 1700
rect 13612 1660 13652 1700
rect 15244 1660 15284 1700
rect 16876 1660 16916 1700
rect 27628 1660 27668 1700
rect 38188 1660 38228 1700
rect 39820 1660 39860 1700
rect 40204 1660 40244 1700
rect 3688 1492 3728 1532
rect 3770 1492 3810 1532
rect 3852 1492 3892 1532
rect 3934 1492 3974 1532
rect 4016 1492 4056 1532
rect 18808 1492 18848 1532
rect 18890 1492 18930 1532
rect 18972 1492 19012 1532
rect 19054 1492 19094 1532
rect 19136 1492 19176 1532
rect 33928 1492 33968 1532
rect 34010 1492 34050 1532
rect 34092 1492 34132 1532
rect 34174 1492 34214 1532
rect 34256 1492 34296 1532
rect 9580 1240 9620 1280
rect 11212 1240 11252 1280
rect 14476 1240 14516 1280
rect 17740 1240 17780 1280
rect 17932 1240 17972 1280
rect 19852 1240 19892 1280
rect 21484 1240 21524 1280
rect 23116 1240 23156 1280
rect 25132 1240 25172 1280
rect 26860 1240 26900 1280
rect 29068 1240 29108 1280
rect 29644 1240 29684 1280
rect 31660 1240 31700 1280
rect 32716 1240 32756 1280
rect 33100 1240 33140 1280
rect 33484 1240 33524 1280
rect 34060 1240 34100 1280
rect 37036 1240 37076 1280
rect 37228 1240 37268 1280
rect 37612 1240 37652 1280
rect 29452 1156 29492 1196
rect 32524 1156 32564 1196
rect 32908 1156 32948 1196
rect 33292 1156 33332 1196
rect 33676 1156 33716 1196
rect 34444 1156 34484 1196
rect 34828 1156 34868 1196
rect 35212 1156 35252 1196
rect 37420 1156 37460 1196
rect 37804 1156 37844 1196
rect 40492 1156 40532 1196
rect 40876 1156 40916 1196
rect 41260 1156 41300 1196
rect 2476 1072 2516 1112
rect 3724 1072 3764 1112
rect 4204 1072 4244 1112
rect 4300 1072 4340 1112
rect 4396 1072 4436 1112
rect 4492 1072 4532 1112
rect 4684 1072 4724 1112
rect 4780 1072 4820 1112
rect 4876 1072 4916 1112
rect 6508 1072 6548 1112
rect 7756 1072 7796 1112
rect 8140 1072 8180 1112
rect 9388 1072 9428 1112
rect 9772 1072 9812 1112
rect 11020 1072 11060 1112
rect 11404 1072 11444 1112
rect 12652 1072 12692 1112
rect 13036 1072 13076 1112
rect 14284 1072 14324 1112
rect 16300 1072 16340 1112
rect 17548 1072 17588 1112
rect 18412 1072 18452 1112
rect 19660 1072 19700 1112
rect 20044 1072 20084 1112
rect 21292 1072 21332 1112
rect 21676 1072 21716 1112
rect 22924 1072 22964 1112
rect 23692 1072 23732 1112
rect 24940 1072 24980 1112
rect 25420 1072 25460 1112
rect 26668 1072 26708 1112
rect 27628 1072 27668 1112
rect 28876 1072 28916 1112
rect 29932 1072 29972 1112
rect 30892 1072 30932 1112
rect 31180 1072 31220 1112
rect 35596 1072 35636 1112
rect 36844 1072 36884 1112
rect 3916 988 3956 1028
rect 4972 904 5012 944
rect 7948 904 7988 944
rect 12844 904 12884 944
rect 32332 904 32372 944
rect 34252 904 34292 944
rect 34636 904 34676 944
rect 35020 904 35060 944
rect 40684 904 40724 944
rect 41068 904 41108 944
rect 41452 904 41492 944
rect 4928 736 4968 776
rect 5010 736 5050 776
rect 5092 736 5132 776
rect 5174 736 5214 776
rect 5256 736 5296 776
rect 20048 736 20088 776
rect 20130 736 20170 776
rect 20212 736 20252 776
rect 20294 736 20334 776
rect 20376 736 20416 776
rect 35168 736 35208 776
rect 35250 736 35290 776
rect 35332 736 35372 776
rect 35414 736 35454 776
rect 35496 736 35536 776
<< metal2 >>
rect 8907 10688 8949 10697
rect 8907 10648 8908 10688
rect 8948 10648 8949 10688
rect 9464 10688 9544 10752
rect 9464 10672 9484 10688
rect 8907 10639 8949 10648
rect 9483 10648 9484 10672
rect 9524 10672 9544 10688
rect 9656 10672 9736 10752
rect 9848 10672 9928 10752
rect 10040 10672 10120 10752
rect 10232 10672 10312 10752
rect 10424 10672 10504 10752
rect 10616 10672 10696 10752
rect 10808 10672 10888 10752
rect 11000 10672 11080 10752
rect 11192 10672 11272 10752
rect 11384 10672 11464 10752
rect 11576 10672 11656 10752
rect 11768 10672 11848 10752
rect 11960 10672 12040 10752
rect 12152 10672 12232 10752
rect 12344 10672 12424 10752
rect 12536 10672 12616 10752
rect 12728 10672 12808 10752
rect 12920 10672 13000 10752
rect 13112 10672 13192 10752
rect 13304 10672 13384 10752
rect 13496 10672 13576 10752
rect 13688 10672 13768 10752
rect 13880 10672 13960 10752
rect 14072 10672 14152 10752
rect 14264 10672 14344 10752
rect 14456 10672 14536 10752
rect 14648 10672 14728 10752
rect 14840 10672 14920 10752
rect 15032 10672 15112 10752
rect 15224 10672 15304 10752
rect 15416 10672 15496 10752
rect 15608 10672 15688 10752
rect 15800 10672 15880 10752
rect 15992 10672 16072 10752
rect 16184 10672 16264 10752
rect 16376 10672 16456 10752
rect 16568 10672 16648 10752
rect 16760 10672 16840 10752
rect 16952 10672 17032 10752
rect 17144 10672 17224 10752
rect 17336 10672 17416 10752
rect 17528 10672 17608 10752
rect 17720 10672 17800 10752
rect 17912 10672 17992 10752
rect 18104 10672 18184 10752
rect 18296 10672 18376 10752
rect 18488 10672 18568 10752
rect 18680 10672 18760 10752
rect 18872 10672 18952 10752
rect 19064 10672 19144 10752
rect 19256 10672 19336 10752
rect 19448 10672 19528 10752
rect 19640 10672 19720 10752
rect 19832 10672 19912 10752
rect 20024 10672 20104 10752
rect 20216 10672 20296 10752
rect 20408 10672 20488 10752
rect 20600 10688 20680 10752
rect 20600 10672 20620 10688
rect 9524 10648 9525 10672
rect 9483 10639 9525 10648
rect 2763 10184 2805 10193
rect 2763 10144 2764 10184
rect 2804 10144 2805 10184
rect 2763 10135 2805 10144
rect 1899 9932 1941 9941
rect 1899 9892 1900 9932
rect 1940 9892 1941 9932
rect 1899 9883 1941 9892
rect 1900 9512 1940 9883
rect 1900 9185 1940 9472
rect 1899 9176 1941 9185
rect 1899 9136 1900 9176
rect 1940 9136 1941 9176
rect 1899 9127 1941 9136
rect 1803 9008 1845 9017
rect 1803 8968 1804 9008
rect 1844 8968 1845 9008
rect 1803 8959 1845 8968
rect 1708 8840 1748 8849
rect 1612 8800 1708 8840
rect 1419 8168 1461 8177
rect 1419 8128 1420 8168
rect 1460 8128 1461 8168
rect 1419 8119 1461 8128
rect 1227 6488 1269 6497
rect 1227 6448 1228 6488
rect 1268 6448 1269 6488
rect 1227 6439 1269 6448
rect 1228 5489 1268 6439
rect 1227 5480 1269 5489
rect 1227 5440 1228 5480
rect 1268 5440 1269 5480
rect 1227 5431 1269 5440
rect 1420 5405 1460 8119
rect 1515 6824 1557 6833
rect 1515 6784 1516 6824
rect 1556 6784 1557 6824
rect 1515 6775 1557 6784
rect 1516 5909 1556 6775
rect 1612 6474 1652 8800
rect 1708 8791 1748 8800
rect 1708 8672 1748 8681
rect 1708 8177 1748 8632
rect 1707 8168 1749 8177
rect 1707 8128 1708 8168
rect 1748 8128 1749 8168
rect 1707 8119 1749 8128
rect 1708 7160 1748 7169
rect 1804 7160 1844 8959
rect 1899 8840 1941 8849
rect 1899 8800 1900 8840
rect 1940 8800 1941 8840
rect 1899 8791 1941 8800
rect 1900 8706 1940 8791
rect 2092 8765 2132 8796
rect 2091 8756 2133 8765
rect 2091 8716 2092 8756
rect 2132 8716 2133 8756
rect 2091 8707 2133 8716
rect 2092 8672 2132 8707
rect 1899 8504 1941 8513
rect 1899 8464 1900 8504
rect 1940 8464 1941 8504
rect 1899 8455 1941 8464
rect 1748 7120 1844 7160
rect 1900 8000 1940 8455
rect 2092 8429 2132 8632
rect 2091 8420 2133 8429
rect 2091 8380 2092 8420
rect 2132 8380 2133 8420
rect 2091 8371 2133 8380
rect 1708 6581 1748 7120
rect 1900 6917 1940 7960
rect 2475 7160 2517 7169
rect 2475 7120 2476 7160
rect 2516 7120 2517 7160
rect 2475 7111 2517 7120
rect 1899 6908 1941 6917
rect 1899 6868 1900 6908
rect 1940 6868 1941 6908
rect 1899 6859 1941 6868
rect 1707 6572 1749 6581
rect 1707 6532 1708 6572
rect 1748 6532 1749 6572
rect 1707 6523 1749 6532
rect 1612 6434 1748 6474
rect 1611 6320 1653 6329
rect 1611 6280 1612 6320
rect 1652 6280 1653 6320
rect 1611 6271 1653 6280
rect 1515 5900 1557 5909
rect 1515 5860 1516 5900
rect 1556 5860 1557 5900
rect 1515 5851 1557 5860
rect 1419 5396 1461 5405
rect 1419 5356 1420 5396
rect 1460 5356 1461 5396
rect 1419 5347 1461 5356
rect 1420 2624 1460 5347
rect 1516 4136 1556 5851
rect 1612 5648 1652 6271
rect 1708 5993 1748 6434
rect 1899 6320 1941 6329
rect 1899 6280 1900 6320
rect 1940 6280 1941 6320
rect 1899 6271 1941 6280
rect 1707 5984 1749 5993
rect 1707 5944 1708 5984
rect 1748 5944 1749 5984
rect 1707 5935 1749 5944
rect 1612 5599 1652 5608
rect 1803 5228 1845 5237
rect 1803 5188 1804 5228
rect 1844 5188 1845 5228
rect 1803 5179 1845 5188
rect 1707 4976 1749 4985
rect 1707 4936 1708 4976
rect 1748 4936 1749 4976
rect 1707 4927 1749 4936
rect 1708 4842 1748 4927
rect 1612 4136 1652 4145
rect 1516 4096 1612 4136
rect 1612 4087 1652 4096
rect 1612 3464 1652 3473
rect 1804 3464 1844 5179
rect 1652 3424 1844 3464
rect 1612 3415 1652 3424
rect 1804 2624 1844 2633
rect 1420 2584 1804 2624
rect 1804 2575 1844 2584
rect 1900 1952 1940 6271
rect 2476 5489 2516 7111
rect 2764 7001 2804 10135
rect 4928 9848 5296 9857
rect 4968 9808 5010 9848
rect 5050 9808 5092 9848
rect 5132 9808 5174 9848
rect 5214 9808 5256 9848
rect 4928 9799 5296 9808
rect 3723 9680 3765 9689
rect 3723 9640 3724 9680
rect 3764 9640 3765 9680
rect 3723 9631 3765 9640
rect 4012 9680 4052 9689
rect 5739 9680 5781 9689
rect 4052 9640 4148 9680
rect 4012 9631 4052 9640
rect 3531 9596 3573 9605
rect 3531 9556 3532 9596
rect 3572 9556 3573 9596
rect 3531 9547 3573 9556
rect 3148 9512 3188 9521
rect 3148 8714 3188 9472
rect 3435 9512 3477 9521
rect 3435 9472 3436 9512
rect 3476 9472 3477 9512
rect 3435 9463 3477 9472
rect 3339 9428 3381 9437
rect 3339 9388 3340 9428
rect 3380 9388 3381 9428
rect 3339 9379 3381 9388
rect 3340 9344 3380 9379
rect 3340 9293 3380 9304
rect 3340 8714 3380 8723
rect 3148 8674 3340 8714
rect 3148 8000 3188 8674
rect 3244 8597 3284 8674
rect 3340 8665 3380 8674
rect 3436 8672 3476 9463
rect 3532 9462 3572 9547
rect 3628 9512 3668 9523
rect 3628 9437 3668 9472
rect 3724 9512 3764 9631
rect 3724 9463 3764 9472
rect 3819 9512 3861 9521
rect 3819 9472 3820 9512
rect 3860 9472 3861 9512
rect 3819 9463 3861 9472
rect 3627 9428 3669 9437
rect 3627 9388 3628 9428
rect 3668 9388 3669 9428
rect 3627 9379 3669 9388
rect 3820 9378 3860 9463
rect 3531 9344 3573 9353
rect 3531 9304 3532 9344
rect 3572 9304 3573 9344
rect 3531 9295 3573 9304
rect 3532 8924 3572 9295
rect 3688 9092 4056 9101
rect 3728 9052 3770 9092
rect 3810 9052 3852 9092
rect 3892 9052 3934 9092
rect 3974 9052 4016 9092
rect 3688 9043 4056 9052
rect 3532 8875 3572 8884
rect 3724 8681 3764 8766
rect 3723 8672 3765 8681
rect 3436 8632 3724 8672
rect 3764 8632 3765 8672
rect 3723 8623 3765 8632
rect 3243 8588 3285 8597
rect 3243 8548 3244 8588
rect 3284 8548 3285 8588
rect 3243 8539 3285 8548
rect 3532 8504 3572 8513
rect 3819 8504 3861 8513
rect 3436 8464 3532 8504
rect 3572 8464 3764 8504
rect 3339 8168 3381 8177
rect 3339 8128 3340 8168
rect 3380 8128 3381 8168
rect 3339 8119 3381 8128
rect 3340 8034 3380 8119
rect 2956 7160 2996 7169
rect 3148 7160 3188 7960
rect 2860 7120 2956 7160
rect 2996 7120 3188 7160
rect 3436 7160 3476 8464
rect 3532 8455 3572 8464
rect 3531 8252 3573 8261
rect 3531 8212 3532 8252
rect 3572 8212 3573 8252
rect 3531 8203 3573 8212
rect 3532 7412 3572 8203
rect 3724 8000 3764 8464
rect 3819 8464 3820 8504
rect 3860 8464 3861 8504
rect 3819 8455 3861 8464
rect 3820 8168 3860 8455
rect 3820 8119 3860 8128
rect 3915 8168 3957 8177
rect 3915 8128 3916 8168
rect 3956 8128 3957 8168
rect 3915 8119 3957 8128
rect 3724 7951 3764 7960
rect 3916 8000 3956 8119
rect 3916 7951 3956 7960
rect 4012 8000 4052 8009
rect 4108 8000 4148 9640
rect 5739 9640 5740 9680
rect 5780 9640 5781 9680
rect 5739 9631 5781 9640
rect 5355 9596 5397 9605
rect 5355 9556 5356 9596
rect 5396 9556 5397 9596
rect 5355 9547 5397 9556
rect 4204 9512 4244 9521
rect 4204 8681 4244 9472
rect 4300 9512 4340 9521
rect 4203 8672 4245 8681
rect 4203 8632 4204 8672
rect 4244 8632 4245 8672
rect 4203 8623 4245 8632
rect 4300 8345 4340 9472
rect 4395 9512 4437 9521
rect 4395 9472 4396 9512
rect 4436 9472 4437 9512
rect 4395 9463 4437 9472
rect 4492 9512 4532 9523
rect 4299 8336 4341 8345
rect 4299 8296 4300 8336
rect 4340 8296 4341 8336
rect 4299 8287 4341 8296
rect 4300 8168 4340 8287
rect 4300 8128 4348 8168
rect 4308 8016 4348 8128
rect 4052 7960 4148 8000
rect 4300 8007 4348 8016
rect 4340 7967 4348 8007
rect 4300 7960 4348 7967
rect 4012 7951 4052 7960
rect 4300 7958 4340 7960
rect 3688 7580 4056 7589
rect 3728 7540 3770 7580
rect 3810 7540 3852 7580
rect 3892 7540 3934 7580
rect 3974 7540 4016 7580
rect 3688 7531 4056 7540
rect 3628 7412 3668 7421
rect 3532 7372 3628 7412
rect 3628 7363 3668 7372
rect 4396 7412 4436 9463
rect 4492 9437 4532 9472
rect 4588 9512 4628 9521
rect 4780 9512 4820 9521
rect 4491 9428 4533 9437
rect 4491 9388 4492 9428
rect 4532 9388 4533 9428
rect 4491 9379 4533 9388
rect 4492 9260 4532 9269
rect 4492 8009 4532 9220
rect 4588 8261 4628 9472
rect 4684 9472 4780 9512
rect 4684 8849 4724 9472
rect 4780 9463 4820 9472
rect 4876 9512 4916 9521
rect 5260 9512 5300 9521
rect 4876 9353 4916 9472
rect 5033 9497 5073 9506
rect 4875 9344 4917 9353
rect 4875 9304 4876 9344
rect 4916 9304 4917 9344
rect 4875 9295 4917 9304
rect 5033 9176 5073 9457
rect 5033 9136 5108 9176
rect 4683 8840 4725 8849
rect 5068 8840 5108 9136
rect 5163 9008 5205 9017
rect 5163 8968 5164 9008
rect 5204 8968 5205 9008
rect 5163 8959 5205 8968
rect 5164 8924 5204 8959
rect 5164 8873 5204 8884
rect 4683 8800 4684 8840
rect 4724 8800 4725 8840
rect 4683 8791 4725 8800
rect 4780 8800 5108 8840
rect 4587 8252 4629 8261
rect 4587 8212 4588 8252
rect 4628 8212 4629 8252
rect 4587 8203 4629 8212
rect 4491 8000 4533 8009
rect 4491 7960 4492 8000
rect 4532 7960 4533 8000
rect 4491 7951 4533 7960
rect 4588 8000 4628 8009
rect 4588 7412 4628 7960
rect 4684 8000 4724 8009
rect 4684 7673 4724 7960
rect 4780 7832 4820 8800
rect 4972 8672 5012 8683
rect 4972 8597 5012 8632
rect 4971 8588 5013 8597
rect 4971 8548 4972 8588
rect 5012 8548 5013 8588
rect 4971 8539 5013 8548
rect 5260 8513 5300 9472
rect 5356 9512 5396 9547
rect 5740 9546 5780 9631
rect 5931 9596 5973 9605
rect 5931 9556 5932 9596
rect 5972 9556 5973 9596
rect 5931 9547 5973 9556
rect 5356 9461 5396 9472
rect 5452 9512 5492 9521
rect 5452 9017 5492 9472
rect 5548 9512 5588 9521
rect 5836 9512 5876 9521
rect 5588 9472 5684 9512
rect 5548 9463 5588 9472
rect 5451 9008 5493 9017
rect 5451 8968 5452 9008
rect 5492 8968 5493 9008
rect 5451 8959 5493 8968
rect 5452 8672 5492 8959
rect 5547 8840 5589 8849
rect 5547 8800 5548 8840
rect 5588 8800 5589 8840
rect 5547 8791 5589 8800
rect 5452 8623 5492 8632
rect 5548 8672 5588 8791
rect 5548 8623 5588 8632
rect 5259 8504 5301 8513
rect 5644 8504 5684 9472
rect 5836 9353 5876 9472
rect 5932 9512 5972 9547
rect 5932 9461 5972 9472
rect 6028 9512 6068 9521
rect 6220 9512 6260 9521
rect 6068 9472 6220 9512
rect 5835 9344 5877 9353
rect 6028 9344 6068 9472
rect 6220 9463 6260 9472
rect 6412 9512 6452 9521
rect 5835 9304 5836 9344
rect 5876 9304 5877 9344
rect 5835 9295 5877 9304
rect 5932 9304 6068 9344
rect 5932 8681 5972 9304
rect 6316 9260 6356 9269
rect 6028 9220 6316 9260
rect 5931 8672 5973 8681
rect 5931 8632 5932 8672
rect 5972 8632 5973 8672
rect 5931 8623 5973 8632
rect 5259 8464 5260 8504
rect 5300 8464 5301 8504
rect 5259 8455 5301 8464
rect 5452 8464 5684 8504
rect 5740 8504 5780 8513
rect 4928 8336 5296 8345
rect 4968 8296 5010 8336
rect 5050 8296 5092 8336
rect 5132 8296 5174 8336
rect 5214 8296 5256 8336
rect 4928 8287 5296 8296
rect 5355 8000 5397 8009
rect 5355 7960 5356 8000
rect 5396 7960 5397 8000
rect 5355 7951 5397 7960
rect 5452 8000 5492 8464
rect 5740 8252 5780 8464
rect 5835 8336 5877 8345
rect 5835 8296 5836 8336
rect 5876 8296 5877 8336
rect 5835 8287 5877 8296
rect 5452 7951 5492 7960
rect 5548 8212 5780 8252
rect 5548 8000 5588 8212
rect 5548 7951 5588 7960
rect 5643 8000 5685 8009
rect 5643 7960 5644 8000
rect 5684 7960 5685 8000
rect 5643 7951 5685 7960
rect 5356 7866 5396 7951
rect 5644 7866 5684 7951
rect 4972 7832 5012 7841
rect 4780 7792 4972 7832
rect 4972 7783 5012 7792
rect 5451 7832 5493 7841
rect 5451 7792 5452 7832
rect 5492 7792 5493 7832
rect 5451 7783 5493 7792
rect 5355 7748 5397 7757
rect 5355 7708 5356 7748
rect 5396 7708 5397 7748
rect 5355 7699 5397 7708
rect 4683 7664 4725 7673
rect 4683 7624 4684 7664
rect 4724 7624 4725 7664
rect 4683 7615 4725 7624
rect 4396 7363 4436 7372
rect 4492 7372 4628 7412
rect 3628 7160 3668 7169
rect 3436 7120 3628 7160
rect 2763 6992 2805 7001
rect 2763 6952 2764 6992
rect 2804 6952 2805 6992
rect 2763 6943 2805 6952
rect 2764 6488 2804 6943
rect 2860 6497 2900 7120
rect 2956 7111 2996 7120
rect 3628 7111 3668 7120
rect 3819 7160 3861 7169
rect 3819 7120 3820 7160
rect 3860 7120 3861 7160
rect 3819 7111 3861 7120
rect 3916 7160 3956 7169
rect 3820 7026 3860 7111
rect 3148 6992 3188 7001
rect 2764 6439 2804 6448
rect 2859 6488 2901 6497
rect 2859 6448 2860 6488
rect 2900 6448 2901 6488
rect 2859 6439 2901 6448
rect 2860 5648 2900 6439
rect 2475 5480 2517 5489
rect 2475 5440 2476 5480
rect 2516 5440 2517 5480
rect 2475 5431 2517 5440
rect 2476 5237 2516 5431
rect 2475 5228 2517 5237
rect 2475 5188 2476 5228
rect 2516 5188 2517 5228
rect 2475 5179 2517 5188
rect 2860 4976 2900 5608
rect 3052 5480 3092 5489
rect 3052 5237 3092 5440
rect 3051 5228 3093 5237
rect 3051 5188 3052 5228
rect 3092 5188 3093 5228
rect 3051 5179 3093 5188
rect 3148 4985 3188 6952
rect 3916 6749 3956 7120
rect 4107 7160 4149 7169
rect 4107 7120 4108 7160
rect 4148 7120 4149 7160
rect 4107 7111 4149 7120
rect 4395 7160 4437 7169
rect 4395 7120 4396 7160
rect 4436 7120 4437 7160
rect 4395 7111 4437 7120
rect 4011 7076 4053 7085
rect 4011 7036 4012 7076
rect 4052 7036 4053 7076
rect 4011 7027 4053 7036
rect 3915 6740 3957 6749
rect 3915 6700 3916 6740
rect 3956 6700 3957 6740
rect 3915 6691 3957 6700
rect 4012 6497 4052 7027
rect 4108 7026 4148 7111
rect 4396 7026 4436 7111
rect 4492 6740 4532 7372
rect 4587 7244 4629 7253
rect 4587 7204 4588 7244
rect 4628 7204 4629 7244
rect 4587 7195 4629 7204
rect 4588 7160 4628 7195
rect 4588 7109 4628 7120
rect 4396 6700 4532 6740
rect 4587 6740 4629 6749
rect 4587 6700 4588 6740
rect 4628 6700 4629 6740
rect 4011 6488 4053 6497
rect 4011 6448 4012 6488
rect 4052 6448 4053 6488
rect 4011 6439 4053 6448
rect 4012 6354 4052 6439
rect 4203 6320 4245 6329
rect 4203 6280 4204 6320
rect 4244 6280 4245 6320
rect 4203 6271 4245 6280
rect 4204 6186 4244 6271
rect 3688 6068 4056 6077
rect 3728 6028 3770 6068
rect 3810 6028 3852 6068
rect 3892 6028 3934 6068
rect 3974 6028 4016 6068
rect 3688 6019 4056 6028
rect 4396 5993 4436 6700
rect 4587 6691 4629 6700
rect 4491 6572 4533 6581
rect 4491 6532 4492 6572
rect 4532 6532 4533 6572
rect 4491 6523 4533 6532
rect 4492 6438 4532 6523
rect 4203 5984 4245 5993
rect 4203 5944 4204 5984
rect 4244 5944 4245 5984
rect 4203 5935 4245 5944
rect 4395 5984 4437 5993
rect 4395 5944 4396 5984
rect 4436 5944 4437 5984
rect 4395 5935 4437 5944
rect 4204 5732 4244 5935
rect 4300 5825 4340 5910
rect 4588 5900 4628 6691
rect 4684 6572 4724 7615
rect 4779 7160 4821 7169
rect 4779 7120 4780 7160
rect 4820 7120 4821 7160
rect 4779 7111 4821 7120
rect 4780 6656 4820 7111
rect 4928 6824 5296 6833
rect 4968 6784 5010 6824
rect 5050 6784 5092 6824
rect 5132 6784 5174 6824
rect 5214 6784 5256 6824
rect 4928 6775 5296 6784
rect 5356 6656 5396 7699
rect 4780 6616 4916 6656
rect 4684 6532 4820 6572
rect 4684 6474 4724 6483
rect 4684 6329 4724 6434
rect 4683 6320 4725 6329
rect 4683 6280 4684 6320
rect 4724 6280 4725 6320
rect 4683 6271 4725 6280
rect 4780 6245 4820 6532
rect 4779 6236 4821 6245
rect 4779 6196 4780 6236
rect 4820 6196 4821 6236
rect 4779 6187 4821 6196
rect 4779 6068 4821 6077
rect 4779 6028 4780 6068
rect 4820 6028 4821 6068
rect 4779 6019 4821 6028
rect 4684 5900 4724 5909
rect 4588 5860 4684 5900
rect 4299 5816 4341 5825
rect 4299 5776 4300 5816
rect 4340 5776 4341 5816
rect 4299 5767 4341 5776
rect 4588 5732 4628 5860
rect 4684 5851 4724 5860
rect 4204 5692 4271 5732
rect 4231 5667 4271 5692
rect 4396 5692 4628 5732
rect 4231 5648 4340 5667
rect 4231 5627 4300 5648
rect 4300 5599 4340 5608
rect 4396 5480 4436 5692
rect 4780 5657 4820 6019
rect 4779 5648 4821 5657
rect 4779 5608 4780 5648
rect 4820 5608 4821 5648
rect 4779 5599 4821 5608
rect 4300 5440 4436 5480
rect 4492 5480 4532 5489
rect 4876 5480 4916 6616
rect 5260 6616 5396 6656
rect 5164 6497 5204 6582
rect 5163 6488 5205 6497
rect 5163 6448 5164 6488
rect 5204 6448 5205 6488
rect 5163 6439 5205 6448
rect 5163 6320 5205 6329
rect 5163 6280 5164 6320
rect 5204 6280 5205 6320
rect 5163 6271 5205 6280
rect 5164 5657 5204 6271
rect 5163 5648 5205 5657
rect 5163 5608 5164 5648
rect 5204 5608 5205 5648
rect 5163 5599 5205 5608
rect 5260 5648 5300 6616
rect 5452 5648 5492 7783
rect 5836 7328 5876 8287
rect 5932 8261 5972 8623
rect 5931 8252 5973 8261
rect 5931 8212 5932 8252
rect 5972 8212 5973 8252
rect 5931 8203 5973 8212
rect 5932 8000 5972 8203
rect 6028 8177 6068 9220
rect 6316 9211 6356 9220
rect 6412 8840 6452 9472
rect 6892 9512 6932 9521
rect 6604 9260 6644 9269
rect 6604 8849 6644 9220
rect 6892 8849 6932 9472
rect 6987 9512 7029 9521
rect 6987 9472 6988 9512
rect 7028 9472 7029 9512
rect 6987 9463 7029 9472
rect 7276 9512 7316 9521
rect 6988 9378 7028 9463
rect 7179 9428 7221 9437
rect 7276 9428 7316 9472
rect 7564 9512 7604 9523
rect 7564 9437 7604 9472
rect 7851 9512 7893 9521
rect 7851 9472 7852 9512
rect 7892 9472 7893 9512
rect 7851 9463 7893 9472
rect 8812 9512 8852 9521
rect 7179 9388 7180 9428
rect 7220 9388 7316 9428
rect 7563 9428 7605 9437
rect 7563 9388 7564 9428
rect 7604 9388 7605 9428
rect 7179 9379 7221 9388
rect 7563 9379 7605 9388
rect 7467 9344 7509 9353
rect 7467 9304 7468 9344
rect 7508 9304 7509 9344
rect 7467 9295 7509 9304
rect 7468 9008 7508 9295
rect 7468 8968 7700 9008
rect 6316 8800 6452 8840
rect 6603 8840 6645 8849
rect 6603 8800 6604 8840
rect 6644 8800 6645 8840
rect 6123 8672 6165 8681
rect 6123 8632 6124 8672
rect 6164 8632 6165 8672
rect 6123 8623 6165 8632
rect 6220 8672 6260 8681
rect 6124 8538 6164 8623
rect 6220 8345 6260 8632
rect 6219 8336 6261 8345
rect 6219 8296 6220 8336
rect 6260 8296 6261 8336
rect 6219 8287 6261 8296
rect 6027 8168 6069 8177
rect 6027 8128 6028 8168
rect 6068 8128 6069 8168
rect 6027 8119 6069 8128
rect 5932 7951 5972 7960
rect 6028 8000 6068 8009
rect 6028 7757 6068 7960
rect 6316 7841 6356 8800
rect 6603 8791 6645 8800
rect 6891 8840 6933 8849
rect 6891 8800 6892 8840
rect 6932 8800 6933 8840
rect 6891 8791 6933 8800
rect 6604 8672 6644 8681
rect 6604 8261 6644 8632
rect 6699 8672 6741 8681
rect 6699 8632 6700 8672
rect 6740 8632 6741 8672
rect 6699 8623 6741 8632
rect 7180 8672 7220 8681
rect 6700 8538 6740 8623
rect 6603 8252 6645 8261
rect 6603 8212 6604 8252
rect 6644 8212 6645 8252
rect 6603 8203 6645 8212
rect 6412 8044 6932 8084
rect 6412 8000 6452 8044
rect 6412 7951 6452 7960
rect 6508 7916 6548 7925
rect 6315 7832 6357 7841
rect 6315 7792 6316 7832
rect 6356 7792 6357 7832
rect 6315 7783 6357 7792
rect 6027 7748 6069 7757
rect 6027 7708 6028 7748
rect 6068 7708 6069 7748
rect 6027 7699 6069 7708
rect 6508 7328 6548 7876
rect 5740 7288 5876 7328
rect 6316 7288 6548 7328
rect 5643 6824 5685 6833
rect 5643 6784 5644 6824
rect 5684 6784 5685 6824
rect 5643 6775 5685 6784
rect 5644 6404 5684 6775
rect 5740 6572 5780 7288
rect 5836 7160 5876 7171
rect 5836 7085 5876 7120
rect 5835 7076 5877 7085
rect 5835 7036 5836 7076
rect 5876 7036 5877 7076
rect 5835 7027 5877 7036
rect 6028 6992 6068 7001
rect 5740 6532 5876 6572
rect 5644 6245 5684 6364
rect 5739 6404 5781 6413
rect 5739 6364 5740 6404
rect 5780 6364 5781 6404
rect 5739 6355 5781 6364
rect 5740 6270 5780 6355
rect 5643 6236 5685 6245
rect 5643 6196 5644 6236
rect 5684 6196 5685 6236
rect 5643 6187 5685 6196
rect 5836 5993 5876 6532
rect 6028 6497 6068 6952
rect 6219 6992 6261 7001
rect 6219 6952 6220 6992
rect 6260 6952 6261 6992
rect 6219 6943 6261 6952
rect 6220 6858 6260 6943
rect 6027 6488 6069 6497
rect 6027 6448 6028 6488
rect 6068 6448 6069 6488
rect 6027 6439 6069 6448
rect 6124 6488 6164 6497
rect 6124 6329 6164 6448
rect 6220 6488 6260 6497
rect 6220 6413 6260 6448
rect 6219 6404 6261 6413
rect 6219 6364 6220 6404
rect 6260 6364 6261 6404
rect 6219 6355 6261 6364
rect 6123 6320 6165 6329
rect 6123 6280 6124 6320
rect 6164 6280 6165 6320
rect 6123 6271 6165 6280
rect 6220 6152 6260 6355
rect 6316 6329 6356 7288
rect 6412 7160 6452 7169
rect 6315 6320 6357 6329
rect 6315 6280 6316 6320
rect 6356 6280 6357 6320
rect 6315 6271 6357 6280
rect 6028 6112 6260 6152
rect 5835 5984 5877 5993
rect 5835 5944 5836 5984
rect 5876 5944 5877 5984
rect 5835 5935 5877 5944
rect 5739 5816 5781 5825
rect 5739 5776 5740 5816
rect 5780 5776 5781 5816
rect 5739 5767 5781 5776
rect 5164 5514 5204 5599
rect 5260 5489 5300 5608
rect 5356 5608 5492 5648
rect 5547 5648 5589 5657
rect 5547 5608 5548 5648
rect 5588 5608 5589 5648
rect 3916 5144 3956 5153
rect 3531 5060 3573 5069
rect 3531 5020 3532 5060
rect 3572 5020 3573 5060
rect 3531 5011 3573 5020
rect 2956 4976 2996 4985
rect 2860 4936 2956 4976
rect 2763 4388 2805 4397
rect 2763 4348 2764 4388
rect 2804 4348 2805 4388
rect 2763 4339 2805 4348
rect 2667 3968 2709 3977
rect 2667 3928 2668 3968
rect 2708 3928 2709 3968
rect 2667 3919 2709 3928
rect 2668 2540 2708 3919
rect 2764 3809 2804 4339
rect 2860 4136 2900 4936
rect 2956 4927 2996 4936
rect 3147 4976 3189 4985
rect 3147 4936 3148 4976
rect 3188 4936 3189 4976
rect 3147 4927 3189 4936
rect 3339 4892 3381 4901
rect 3339 4852 3340 4892
rect 3380 4852 3381 4892
rect 3339 4843 3381 4852
rect 3147 4808 3189 4817
rect 3147 4768 3148 4808
rect 3188 4768 3189 4808
rect 3147 4759 3189 4768
rect 3148 4674 3188 4759
rect 3340 4229 3380 4843
rect 3435 4724 3477 4733
rect 3435 4684 3436 4724
rect 3476 4684 3477 4724
rect 3435 4675 3477 4684
rect 3339 4220 3381 4229
rect 3339 4180 3340 4220
rect 3380 4180 3381 4220
rect 3339 4171 3381 4180
rect 2763 3800 2805 3809
rect 2763 3760 2764 3800
rect 2804 3760 2805 3800
rect 2763 3751 2805 3760
rect 2860 3464 2900 4096
rect 3052 3968 3092 3977
rect 3052 3809 3092 3928
rect 3051 3800 3093 3809
rect 3051 3760 3052 3800
rect 3092 3760 3093 3800
rect 3051 3751 3093 3760
rect 3052 3548 3092 3559
rect 3052 3473 3092 3508
rect 3436 3473 3476 4675
rect 3532 4388 3572 5011
rect 3628 4976 3668 4985
rect 3628 4733 3668 4936
rect 3724 4976 3764 4987
rect 3724 4901 3764 4936
rect 3723 4892 3765 4901
rect 3723 4852 3724 4892
rect 3764 4852 3765 4892
rect 3723 4843 3765 4852
rect 3916 4733 3956 5104
rect 4108 4985 4148 5070
rect 4107 4976 4149 4985
rect 4107 4936 4108 4976
rect 4148 4936 4149 4976
rect 4107 4927 4149 4936
rect 4300 4976 4340 5440
rect 4300 4927 4340 4936
rect 4396 4976 4436 4985
rect 4396 4817 4436 4936
rect 4395 4808 4437 4817
rect 4395 4768 4396 4808
rect 4436 4768 4437 4808
rect 4395 4759 4437 4768
rect 3627 4724 3669 4733
rect 3627 4684 3628 4724
rect 3668 4684 3669 4724
rect 3627 4675 3669 4684
rect 3915 4724 3957 4733
rect 3915 4684 3916 4724
rect 3956 4684 3957 4724
rect 3915 4675 3957 4684
rect 4108 4724 4148 4733
rect 4148 4684 4244 4724
rect 4108 4675 4148 4684
rect 3688 4556 4056 4565
rect 3728 4516 3770 4556
rect 3810 4516 3852 4556
rect 3892 4516 3934 4556
rect 3974 4516 4016 4556
rect 3688 4507 4056 4516
rect 3532 4348 3764 4388
rect 3531 4220 3573 4229
rect 3531 4180 3532 4220
rect 3572 4180 3573 4220
rect 3531 4171 3573 4180
rect 3532 4136 3572 4171
rect 3532 4085 3572 4096
rect 3724 4136 3764 4348
rect 4011 4220 4053 4229
rect 4011 4180 4012 4220
rect 4052 4180 4053 4220
rect 4011 4171 4053 4180
rect 3724 4087 3764 4096
rect 3820 4136 3860 4145
rect 3628 3968 3668 3977
rect 2860 2624 2900 3424
rect 3051 3464 3093 3473
rect 3051 3424 3052 3464
rect 3092 3424 3093 3464
rect 3051 3415 3093 3424
rect 3435 3464 3477 3473
rect 3435 3424 3436 3464
rect 3476 3424 3477 3464
rect 3435 3415 3477 3424
rect 3628 3464 3668 3928
rect 3820 3641 3860 4096
rect 4012 3893 4052 4171
rect 4107 4136 4149 4145
rect 4107 4096 4108 4136
rect 4148 4096 4149 4136
rect 4107 4087 4149 4096
rect 4108 4002 4148 4087
rect 4011 3884 4053 3893
rect 4011 3844 4012 3884
rect 4052 3844 4053 3884
rect 4011 3835 4053 3844
rect 4107 3800 4149 3809
rect 4107 3760 4108 3800
rect 4148 3760 4149 3800
rect 4107 3751 4149 3760
rect 3819 3632 3861 3641
rect 3819 3592 3820 3632
rect 3860 3592 3861 3632
rect 3819 3583 3861 3592
rect 3723 3548 3765 3557
rect 3723 3508 3724 3548
rect 3764 3508 3765 3548
rect 3723 3499 3765 3508
rect 3628 3415 3668 3424
rect 3724 3464 3764 3499
rect 3724 3413 3764 3424
rect 3819 3464 3861 3473
rect 3819 3424 3820 3464
rect 3860 3424 3861 3464
rect 3819 3415 3861 3424
rect 3916 3464 3956 3475
rect 4108 3473 4148 3751
rect 3820 3330 3860 3415
rect 3916 3389 3956 3424
rect 4107 3464 4149 3473
rect 4107 3424 4108 3464
rect 4148 3424 4149 3464
rect 4107 3415 4149 3424
rect 4204 3464 4244 4684
rect 4395 4640 4437 4649
rect 4395 4600 4396 4640
rect 4436 4600 4437 4640
rect 4395 4591 4437 4600
rect 4299 4556 4341 4565
rect 4299 4516 4300 4556
rect 4340 4516 4341 4556
rect 4299 4507 4341 4516
rect 4300 3464 4340 4507
rect 4396 4136 4436 4591
rect 4492 4565 4532 5440
rect 4780 5440 4916 5480
rect 5259 5480 5301 5489
rect 5259 5440 5260 5480
rect 5300 5440 5301 5480
rect 4588 4976 4628 4985
rect 4780 4976 4820 5440
rect 5259 5431 5301 5440
rect 4928 5312 5296 5321
rect 4968 5272 5010 5312
rect 5050 5272 5092 5312
rect 5132 5272 5174 5312
rect 5214 5272 5256 5312
rect 4928 5263 5296 5272
rect 5163 5060 5205 5069
rect 5163 5020 5164 5060
rect 5204 5020 5205 5060
rect 5163 5011 5205 5020
rect 4876 4976 4916 4985
rect 4780 4936 4876 4976
rect 4588 4817 4628 4936
rect 4876 4927 4916 4936
rect 5068 4976 5108 4985
rect 5068 4817 5108 4936
rect 5164 4926 5204 5011
rect 5259 4976 5301 4985
rect 5259 4936 5260 4976
rect 5300 4936 5301 4976
rect 5259 4927 5301 4936
rect 5356 4976 5396 5608
rect 5547 5599 5589 5608
rect 5740 5648 5780 5767
rect 5740 5599 5780 5608
rect 5835 5648 5877 5657
rect 5835 5608 5836 5648
rect 5876 5608 5877 5648
rect 5835 5599 5877 5608
rect 5451 5480 5493 5489
rect 5451 5440 5452 5480
rect 5492 5440 5493 5480
rect 5451 5431 5493 5440
rect 5452 5346 5492 5431
rect 5548 5312 5588 5599
rect 5836 5514 5876 5599
rect 6028 5564 6068 6112
rect 6123 5984 6165 5993
rect 6123 5944 6124 5984
rect 6164 5944 6165 5984
rect 6123 5935 6165 5944
rect 5932 5524 6068 5564
rect 5545 5272 5588 5312
rect 5545 5228 5585 5272
rect 5932 5237 5972 5524
rect 5643 5228 5685 5237
rect 5545 5188 5588 5228
rect 5452 4976 5492 4985
rect 5356 4936 5452 4976
rect 5260 4842 5300 4927
rect 4587 4808 4629 4817
rect 4587 4768 4588 4808
rect 4628 4768 4629 4808
rect 4587 4759 4629 4768
rect 5067 4808 5109 4817
rect 5067 4768 5068 4808
rect 5108 4768 5204 4808
rect 5067 4759 5109 4768
rect 4491 4556 4533 4565
rect 4491 4516 4492 4556
rect 4532 4516 4533 4556
rect 4491 4507 4533 4516
rect 4491 4304 4533 4313
rect 4491 4264 4492 4304
rect 4532 4264 4533 4304
rect 4491 4255 4533 4264
rect 4396 4087 4436 4096
rect 4492 4136 4532 4255
rect 4588 4145 4628 4759
rect 4876 4724 4916 4733
rect 4780 4304 4820 4313
rect 4684 4264 4780 4304
rect 4492 4087 4532 4096
rect 4587 4136 4629 4145
rect 4587 4096 4588 4136
rect 4628 4096 4629 4136
rect 4587 4087 4629 4096
rect 4491 3800 4533 3809
rect 4491 3760 4492 3800
rect 4532 3760 4533 3800
rect 4491 3751 4533 3760
rect 4396 3464 4436 3473
rect 4300 3424 4396 3464
rect 4204 3415 4244 3424
rect 4396 3415 4436 3424
rect 4492 3464 4532 3751
rect 4587 3716 4629 3725
rect 4587 3676 4588 3716
rect 4628 3676 4629 3716
rect 4587 3667 4629 3676
rect 4588 3632 4628 3667
rect 4588 3581 4628 3592
rect 4684 3473 4724 4264
rect 4780 4255 4820 4264
rect 4876 4145 4916 4684
rect 5067 4220 5109 4229
rect 5067 4180 5068 4220
rect 5108 4180 5109 4220
rect 5067 4171 5109 4180
rect 4875 4136 4917 4145
rect 4875 4096 4876 4136
rect 4916 4096 4917 4136
rect 4875 4087 4917 4096
rect 5068 4136 5108 4171
rect 5068 4085 5108 4096
rect 5164 4136 5204 4768
rect 5356 4481 5396 4936
rect 5452 4927 5492 4936
rect 5548 4976 5588 5188
rect 5643 5188 5644 5228
rect 5684 5188 5685 5228
rect 5643 5179 5685 5188
rect 5931 5228 5973 5237
rect 5931 5188 5932 5228
rect 5972 5188 5973 5228
rect 5931 5179 5973 5188
rect 5548 4927 5588 4936
rect 5644 4976 5684 5179
rect 5739 5060 5781 5069
rect 5739 5020 5740 5060
rect 5780 5020 5781 5060
rect 5739 5011 5781 5020
rect 5644 4927 5684 4936
rect 5740 4926 5780 5011
rect 6028 4976 6068 4985
rect 6028 4817 6068 4936
rect 6124 4976 6164 5935
rect 6220 5648 6260 5657
rect 6220 5237 6260 5608
rect 6316 5648 6356 6271
rect 6316 5321 6356 5608
rect 6315 5312 6357 5321
rect 6315 5272 6316 5312
rect 6356 5272 6357 5312
rect 6315 5263 6357 5272
rect 6219 5228 6261 5237
rect 6219 5188 6220 5228
rect 6260 5188 6261 5228
rect 6219 5179 6261 5188
rect 6412 5069 6452 7120
rect 6507 7160 6549 7169
rect 6507 7120 6508 7160
rect 6548 7120 6549 7160
rect 6507 7111 6549 7120
rect 6508 7026 6548 7111
rect 6699 6992 6741 7001
rect 6699 6952 6700 6992
rect 6740 6952 6741 6992
rect 6699 6943 6741 6952
rect 6603 6572 6645 6581
rect 6603 6532 6604 6572
rect 6644 6532 6645 6572
rect 6603 6523 6645 6532
rect 6507 6488 6549 6497
rect 6507 6448 6508 6488
rect 6548 6448 6549 6488
rect 6507 6439 6549 6448
rect 6604 6488 6644 6523
rect 6508 6354 6548 6439
rect 6604 6437 6644 6448
rect 6700 6488 6740 6943
rect 6700 6439 6740 6448
rect 6796 6488 6836 6497
rect 6796 6329 6836 6448
rect 6795 6320 6837 6329
rect 6795 6280 6796 6320
rect 6836 6280 6837 6320
rect 6795 6271 6837 6280
rect 6603 6236 6645 6245
rect 6603 6196 6604 6236
rect 6644 6196 6645 6236
rect 6603 6187 6645 6196
rect 6507 6152 6549 6161
rect 6507 6112 6508 6152
rect 6548 6112 6549 6152
rect 6507 6103 6549 6112
rect 6411 5060 6453 5069
rect 6411 5020 6412 5060
rect 6452 5020 6453 5060
rect 6411 5011 6453 5020
rect 6124 4927 6164 4936
rect 6508 4976 6548 6103
rect 6027 4808 6069 4817
rect 6027 4768 6028 4808
rect 6068 4768 6069 4808
rect 6027 4759 6069 4768
rect 6123 4724 6165 4733
rect 6123 4684 6124 4724
rect 6164 4684 6165 4724
rect 6123 4675 6165 4684
rect 5355 4472 5397 4481
rect 5355 4432 5356 4472
rect 5396 4432 5397 4472
rect 5355 4423 5397 4432
rect 5164 4087 5204 4096
rect 5260 4136 5300 4145
rect 5356 4136 5396 4423
rect 5452 4145 5492 4230
rect 5300 4096 5396 4136
rect 5451 4136 5493 4145
rect 5451 4096 5452 4136
rect 5492 4096 5493 4136
rect 5260 4087 5300 4096
rect 5451 4087 5493 4096
rect 5548 4136 5588 4145
rect 4972 3968 5012 3977
rect 5548 3968 5588 4096
rect 5012 3928 5588 3968
rect 5644 4136 5684 4145
rect 4972 3919 5012 3928
rect 4928 3800 5296 3809
rect 4968 3760 5010 3800
rect 5050 3760 5092 3800
rect 5132 3760 5174 3800
rect 5214 3760 5256 3800
rect 4928 3751 5296 3760
rect 4875 3632 4917 3641
rect 4875 3592 4876 3632
rect 4916 3592 4917 3632
rect 4875 3583 4917 3592
rect 5067 3632 5109 3641
rect 5067 3592 5068 3632
rect 5108 3592 5109 3632
rect 5067 3583 5109 3592
rect 4876 3498 4916 3583
rect 4492 3415 4532 3424
rect 4647 3464 4724 3473
rect 4687 3424 4724 3464
rect 5068 3464 5108 3583
rect 5644 3473 5684 4096
rect 5932 4136 5972 4145
rect 5740 3968 5780 3977
rect 5740 3557 5780 3928
rect 5932 3725 5972 4096
rect 6028 4136 6068 4145
rect 5931 3716 5973 3725
rect 5931 3676 5932 3716
rect 5972 3676 5973 3716
rect 5931 3667 5973 3676
rect 5739 3548 5781 3557
rect 5739 3508 5740 3548
rect 5780 3508 5781 3548
rect 5739 3499 5781 3508
rect 4647 3415 4687 3424
rect 3915 3380 3957 3389
rect 3915 3340 3916 3380
rect 3956 3340 3957 3380
rect 3915 3331 3957 3340
rect 4108 3330 4148 3415
rect 3339 3296 3381 3305
rect 3339 3256 3340 3296
rect 3380 3256 3381 3296
rect 3339 3247 3381 3256
rect 3340 2801 3380 3247
rect 4107 3212 4149 3221
rect 4107 3172 4108 3212
rect 4148 3172 4149 3212
rect 4107 3163 4149 3172
rect 3688 3044 4056 3053
rect 3728 3004 3770 3044
rect 3810 3004 3852 3044
rect 3892 3004 3934 3044
rect 3974 3004 4016 3044
rect 3688 2995 4056 3004
rect 4108 2876 4148 3163
rect 4395 2960 4437 2969
rect 4395 2920 4396 2960
rect 4436 2920 4437 2960
rect 4395 2911 4437 2920
rect 4012 2836 4148 2876
rect 3339 2792 3381 2801
rect 3339 2752 3340 2792
rect 3380 2752 3381 2792
rect 3339 2743 3381 2752
rect 3436 2717 3476 2748
rect 3435 2708 3477 2717
rect 3435 2668 3436 2708
rect 3476 2668 3477 2708
rect 3435 2659 3477 2668
rect 3052 2624 3092 2633
rect 2860 2584 3052 2624
rect 2668 2500 2996 2540
rect 1900 1903 1940 1912
rect 1803 1868 1845 1877
rect 1803 1828 1804 1868
rect 1844 1828 1845 1868
rect 1803 1819 1845 1828
rect 1804 80 1844 1819
rect 2475 1112 2517 1121
rect 2475 1072 2476 1112
rect 2516 1072 2517 1112
rect 2475 1063 2517 1072
rect 2476 978 2516 1063
rect 2956 80 2996 2500
rect 3052 2204 3092 2584
rect 3436 2624 3476 2659
rect 3724 2633 3764 2718
rect 3244 2540 3284 2549
rect 3436 2540 3476 2584
rect 3532 2624 3572 2633
rect 3723 2624 3765 2633
rect 3572 2584 3724 2624
rect 3764 2584 3765 2624
rect 3532 2575 3572 2584
rect 3723 2575 3765 2584
rect 3820 2624 3860 2633
rect 3284 2500 3476 2540
rect 3244 2491 3284 2500
rect 3147 2204 3189 2213
rect 3052 2164 3148 2204
rect 3188 2164 3189 2204
rect 3147 2155 3189 2164
rect 3531 2204 3573 2213
rect 3531 2164 3532 2204
rect 3572 2164 3573 2204
rect 3531 2155 3573 2164
rect 3148 1952 3188 2155
rect 3148 1903 3188 1912
rect 3339 1700 3381 1709
rect 3339 1660 3340 1700
rect 3380 1660 3381 1700
rect 3339 1651 3381 1660
rect 3340 1566 3380 1651
rect 3532 1364 3572 2155
rect 3820 1952 3860 2584
rect 4012 2624 4052 2836
rect 4012 2575 4052 2584
rect 4300 2624 4340 2633
rect 4012 2456 4052 2465
rect 3820 1709 3860 1912
rect 3915 1952 3957 1961
rect 3915 1912 3916 1952
rect 3956 1912 3957 1952
rect 3915 1903 3957 1912
rect 4012 1952 4052 2416
rect 4203 2288 4245 2297
rect 4203 2248 4204 2288
rect 4244 2248 4245 2288
rect 4203 2239 4245 2248
rect 4012 1903 4052 1912
rect 4108 1952 4148 1961
rect 3916 1818 3956 1903
rect 3819 1700 3861 1709
rect 3819 1660 3820 1700
rect 3860 1660 3861 1700
rect 3819 1651 3861 1660
rect 3688 1532 4056 1541
rect 3728 1492 3770 1532
rect 3810 1492 3852 1532
rect 3892 1492 3934 1532
rect 3974 1492 4016 1532
rect 3688 1483 4056 1492
rect 3532 1324 3764 1364
rect 3724 1112 3764 1324
rect 4108 1121 4148 1912
rect 3724 1063 3764 1072
rect 4107 1112 4149 1121
rect 4107 1072 4108 1112
rect 4148 1072 4149 1112
rect 4107 1063 4149 1072
rect 4204 1112 4244 2239
rect 4300 1709 4340 2584
rect 4396 2624 4436 2911
rect 4492 2633 4532 2718
rect 4876 2633 4916 2718
rect 4971 2708 5013 2717
rect 4971 2668 4972 2708
rect 5012 2668 5013 2708
rect 4971 2659 5013 2668
rect 4396 2575 4436 2584
rect 4491 2624 4533 2633
rect 4491 2584 4492 2624
rect 4532 2584 4533 2624
rect 4491 2575 4533 2584
rect 4875 2624 4917 2633
rect 4875 2584 4876 2624
rect 4916 2584 4917 2624
rect 4875 2575 4917 2584
rect 4972 2624 5012 2659
rect 4972 2573 5012 2584
rect 4684 2456 4724 2465
rect 5068 2456 5108 3424
rect 5164 3464 5204 3473
rect 5164 3221 5204 3424
rect 5643 3464 5685 3473
rect 5643 3424 5644 3464
rect 5684 3424 5685 3464
rect 5643 3415 5685 3424
rect 6028 3389 6068 4096
rect 6124 4136 6164 4675
rect 6508 4145 6548 4936
rect 6604 4976 6644 6187
rect 6795 5648 6837 5657
rect 6795 5608 6796 5648
rect 6836 5608 6837 5648
rect 6795 5599 6837 5608
rect 6796 5514 6836 5599
rect 6892 5237 6932 8044
rect 6988 8000 7028 8011
rect 6988 7925 7028 7960
rect 6987 7916 7029 7925
rect 6987 7876 6988 7916
rect 7028 7876 7029 7916
rect 6987 7867 7029 7876
rect 7180 6749 7220 8632
rect 7371 8672 7413 8681
rect 7371 8632 7372 8672
rect 7412 8632 7413 8672
rect 7371 8623 7413 8632
rect 7275 7160 7317 7169
rect 7275 7120 7276 7160
rect 7316 7120 7317 7160
rect 7275 7111 7317 7120
rect 7179 6740 7221 6749
rect 7179 6700 7180 6740
rect 7220 6700 7221 6740
rect 7179 6691 7221 6700
rect 7276 6656 7316 7111
rect 7276 6607 7316 6616
rect 6988 6488 7028 6499
rect 6988 6413 7028 6448
rect 7084 6488 7124 6497
rect 6987 6404 7029 6413
rect 6987 6364 6988 6404
rect 7028 6364 7029 6404
rect 6987 6355 7029 6364
rect 6987 5984 7029 5993
rect 6987 5944 6988 5984
rect 7028 5944 7029 5984
rect 6987 5935 7029 5944
rect 6988 5825 7028 5935
rect 6987 5816 7029 5825
rect 6987 5776 6988 5816
rect 7028 5776 7029 5816
rect 6987 5767 7029 5776
rect 6891 5228 6933 5237
rect 6891 5188 6892 5228
rect 6932 5188 6933 5228
rect 6891 5179 6933 5188
rect 6988 4976 7028 5767
rect 7084 5489 7124 6448
rect 7179 6488 7221 6497
rect 7179 6448 7180 6488
rect 7220 6448 7221 6488
rect 7179 6439 7221 6448
rect 7180 6354 7220 6439
rect 7372 6245 7412 8623
rect 7468 7995 7508 8968
rect 7563 8840 7605 8849
rect 7563 8800 7564 8840
rect 7604 8800 7605 8840
rect 7563 8791 7605 8800
rect 7564 8168 7604 8791
rect 7660 8686 7700 8968
rect 7660 8637 7700 8646
rect 7852 8588 7892 9463
rect 8812 9101 8852 9472
rect 8811 9092 8853 9101
rect 8811 9052 8812 9092
rect 8852 9052 8853 9092
rect 8811 9043 8853 9052
rect 8620 8840 8660 8849
rect 8908 8840 8948 10639
rect 9676 9857 9716 10672
rect 9675 9848 9717 9857
rect 9675 9808 9676 9848
rect 9716 9808 9717 9848
rect 9675 9799 9717 9808
rect 9868 9764 9908 10672
rect 9868 9724 10004 9764
rect 9004 9680 9044 9689
rect 9044 9640 9908 9680
rect 9004 9631 9044 9640
rect 9484 9512 9524 9521
rect 9292 9472 9484 9512
rect 8660 8800 8948 8840
rect 9196 9260 9236 9269
rect 8620 8791 8660 8800
rect 9196 8765 9236 9220
rect 8427 8756 8469 8765
rect 8427 8716 8428 8756
rect 8468 8716 8469 8756
rect 8427 8707 8469 8716
rect 9195 8756 9237 8765
rect 9195 8716 9196 8756
rect 9236 8716 9237 8756
rect 9195 8707 9237 8716
rect 8428 8622 8468 8707
rect 8811 8672 8853 8681
rect 8811 8632 8812 8672
rect 8852 8632 8853 8672
rect 8811 8623 8853 8632
rect 7852 8539 7892 8548
rect 8812 8538 8852 8623
rect 7660 8168 7700 8177
rect 7564 8128 7660 8168
rect 7660 8119 7700 8128
rect 7468 7946 7508 7955
rect 9292 7748 9332 9472
rect 9484 9463 9524 9472
rect 9580 9512 9620 9521
rect 9580 9344 9620 9472
rect 9868 9512 9908 9640
rect 9868 9463 9908 9472
rect 9484 9304 9620 9344
rect 9196 7708 9332 7748
rect 9388 7916 9428 7925
rect 7467 7496 7509 7505
rect 7467 7456 7468 7496
rect 7508 7456 7509 7496
rect 7467 7447 7509 7456
rect 7468 6665 7508 7447
rect 8043 7160 8085 7169
rect 8043 7120 8044 7160
rect 8084 7120 8085 7160
rect 8043 7111 8085 7120
rect 8044 7026 8084 7111
rect 7467 6656 7509 6665
rect 7467 6616 7468 6656
rect 7508 6616 7509 6656
rect 9196 6656 9236 7708
rect 9291 7580 9333 7589
rect 9291 7540 9292 7580
rect 9332 7540 9333 7580
rect 9291 7531 9333 7540
rect 9292 7160 9332 7531
rect 9292 7111 9332 7120
rect 9196 6616 9332 6656
rect 7467 6607 7509 6616
rect 7468 6488 7508 6607
rect 8908 6572 8948 6581
rect 8948 6532 9236 6572
rect 8908 6523 8948 6532
rect 7468 6439 7508 6448
rect 8716 6488 8756 6497
rect 8716 6329 8756 6448
rect 8811 6488 8853 6497
rect 8811 6448 8812 6488
rect 8852 6448 8853 6488
rect 8811 6439 8853 6448
rect 9196 6488 9236 6532
rect 9196 6439 9236 6448
rect 7563 6320 7605 6329
rect 7563 6280 7564 6320
rect 7604 6280 7605 6320
rect 7563 6271 7605 6280
rect 8715 6320 8757 6329
rect 8715 6280 8716 6320
rect 8756 6280 8757 6320
rect 8715 6271 8757 6280
rect 7371 6236 7413 6245
rect 7371 6196 7372 6236
rect 7412 6196 7413 6236
rect 7371 6187 7413 6196
rect 7324 5657 7364 5666
rect 7364 5617 7412 5648
rect 7324 5608 7412 5617
rect 7083 5480 7125 5489
rect 7275 5480 7317 5489
rect 7083 5440 7084 5480
rect 7124 5440 7125 5480
rect 7083 5431 7125 5440
rect 7180 5440 7276 5480
rect 7316 5440 7317 5480
rect 7084 4976 7124 4985
rect 6988 4936 7084 4976
rect 6604 4927 6644 4936
rect 6699 4892 6741 4901
rect 6699 4852 6700 4892
rect 6740 4852 6741 4892
rect 6699 4843 6741 4852
rect 6124 4087 6164 4096
rect 6507 4136 6549 4145
rect 6507 4096 6508 4136
rect 6548 4096 6549 4136
rect 6507 4087 6549 4096
rect 6219 3968 6261 3977
rect 6219 3928 6220 3968
rect 6260 3928 6261 3968
rect 6219 3919 6261 3928
rect 6220 3834 6260 3919
rect 6027 3380 6069 3389
rect 6027 3340 6028 3380
rect 6068 3340 6069 3380
rect 6027 3331 6069 3340
rect 6603 3380 6645 3389
rect 6603 3340 6604 3380
rect 6644 3340 6645 3380
rect 6603 3331 6645 3340
rect 5163 3212 5205 3221
rect 5163 3172 5164 3212
rect 5204 3172 5205 3212
rect 5163 3163 5205 3172
rect 5548 2717 5588 2719
rect 5547 2708 5589 2717
rect 5547 2668 5548 2708
rect 5588 2668 5589 2708
rect 5547 2659 5589 2668
rect 5452 2624 5492 2633
rect 4492 2416 4684 2456
rect 4396 2120 4436 2129
rect 4396 1784 4436 2080
rect 4492 2036 4532 2416
rect 4684 2407 4724 2416
rect 4780 2416 5108 2456
rect 5164 2584 5452 2624
rect 5164 2456 5204 2584
rect 5452 2575 5492 2584
rect 5548 2624 5588 2659
rect 4587 2288 4629 2297
rect 4587 2248 4588 2288
rect 4628 2248 4629 2288
rect 4587 2239 4629 2248
rect 4492 1987 4532 1996
rect 4588 1952 4628 2239
rect 4588 1903 4628 1912
rect 4684 1952 4724 1961
rect 4780 1952 4820 2416
rect 5164 2407 5204 2416
rect 5356 2456 5396 2465
rect 4928 2288 5296 2297
rect 4968 2248 5010 2288
rect 5050 2248 5092 2288
rect 5132 2248 5174 2288
rect 5214 2248 5256 2288
rect 4928 2239 5296 2248
rect 5067 2036 5109 2045
rect 5067 1996 5068 2036
rect 5108 1996 5109 2036
rect 5067 1987 5109 1996
rect 4876 1952 4916 1961
rect 4780 1912 4876 1952
rect 4684 1784 4724 1912
rect 4876 1903 4916 1912
rect 5068 1952 5108 1987
rect 5356 1961 5396 2416
rect 5451 2204 5493 2213
rect 5451 2164 5452 2204
rect 5492 2164 5493 2204
rect 5451 2155 5493 2164
rect 4972 1784 5012 1793
rect 4396 1744 4532 1784
rect 4684 1744 4972 1784
rect 4299 1700 4341 1709
rect 4299 1660 4300 1700
rect 4340 1660 4341 1700
rect 4299 1651 4341 1660
rect 4204 1063 4244 1072
rect 4300 1112 4340 1651
rect 4395 1616 4437 1625
rect 4395 1576 4396 1616
rect 4436 1576 4437 1616
rect 4395 1567 4437 1576
rect 4396 1448 4436 1567
rect 4492 1532 4532 1744
rect 4972 1735 5012 1744
rect 4588 1700 4628 1709
rect 4628 1660 4916 1700
rect 4588 1651 4628 1660
rect 4492 1492 4724 1532
rect 4396 1408 4532 1448
rect 4395 1196 4437 1205
rect 4395 1156 4396 1196
rect 4436 1156 4437 1196
rect 4395 1147 4437 1156
rect 4300 1063 4340 1072
rect 4396 1112 4436 1147
rect 4396 1061 4436 1072
rect 4492 1112 4532 1408
rect 4492 1063 4532 1072
rect 4684 1112 4724 1492
rect 4684 1037 4724 1072
rect 4779 1112 4821 1121
rect 4779 1072 4780 1112
rect 4820 1072 4821 1112
rect 4779 1063 4821 1072
rect 4876 1112 4916 1660
rect 5068 1205 5108 1912
rect 5260 1952 5300 1961
rect 5067 1196 5109 1205
rect 5067 1156 5068 1196
rect 5108 1156 5109 1196
rect 5067 1147 5109 1156
rect 4876 1063 4916 1072
rect 3915 1028 3957 1037
rect 3915 988 3916 1028
rect 3956 988 3957 1028
rect 3915 979 3957 988
rect 4683 1028 4725 1037
rect 4683 988 4684 1028
rect 4724 988 4725 1028
rect 4683 979 4725 988
rect 3916 894 3956 979
rect 4780 978 4820 1063
rect 4972 953 5012 1038
rect 5260 1028 5300 1912
rect 5355 1952 5397 1961
rect 5355 1912 5356 1952
rect 5396 1912 5397 1952
rect 5355 1903 5397 1912
rect 5355 1028 5397 1037
rect 5260 988 5356 1028
rect 5396 988 5397 1028
rect 5355 979 5397 988
rect 4107 944 4149 953
rect 4107 904 4108 944
rect 4148 904 4149 944
rect 4107 895 4149 904
rect 4971 944 5013 953
rect 4971 904 4972 944
rect 5012 904 5013 944
rect 4971 895 5013 904
rect 4108 80 4148 895
rect 4928 776 5296 785
rect 4968 736 5010 776
rect 5050 736 5092 776
rect 5132 736 5174 776
rect 5214 736 5256 776
rect 4928 727 5296 736
rect 5356 449 5396 979
rect 5355 440 5397 449
rect 5355 400 5356 440
rect 5396 400 5397 440
rect 5355 391 5397 400
rect 5452 188 5492 2155
rect 5548 2045 5588 2584
rect 5643 2624 5685 2633
rect 5643 2584 5644 2624
rect 5684 2584 5685 2624
rect 5643 2575 5685 2584
rect 6508 2624 6548 2652
rect 6604 2624 6644 3331
rect 6700 3296 6740 4843
rect 7084 4313 7124 4936
rect 7083 4304 7125 4313
rect 7083 4264 7084 4304
rect 7124 4264 7125 4304
rect 7083 4255 7125 4264
rect 6988 4145 7028 4230
rect 6700 3247 6740 3256
rect 6892 4136 6932 4145
rect 6548 2584 6644 2624
rect 6508 2575 6548 2584
rect 5644 2490 5684 2575
rect 5739 2288 5781 2297
rect 5739 2248 5740 2288
rect 5780 2248 5781 2288
rect 5739 2239 5781 2248
rect 5740 2045 5780 2239
rect 6411 2120 6453 2129
rect 6411 2080 6412 2120
rect 6452 2080 6453 2120
rect 6411 2071 6453 2080
rect 5547 2036 5589 2045
rect 5547 1996 5548 2036
rect 5588 1996 5589 2036
rect 5547 1987 5589 1996
rect 5739 2036 5781 2045
rect 5739 1996 5740 2036
rect 5780 1996 5781 2036
rect 5739 1987 5781 1996
rect 6412 1112 6452 2071
rect 6507 1952 6549 1961
rect 6507 1912 6508 1952
rect 6548 1912 6549 1952
rect 6507 1903 6549 1912
rect 6508 1818 6548 1903
rect 6508 1112 6548 1121
rect 6412 1072 6508 1112
rect 6508 1063 6548 1072
rect 6411 944 6453 953
rect 6411 904 6412 944
rect 6452 904 6453 944
rect 6411 895 6453 904
rect 5259 148 5492 188
rect 5259 104 5299 148
rect 5259 80 5300 104
rect 6412 80 6452 895
rect 6604 113 6644 2584
rect 6700 2120 6740 2129
rect 6892 2120 6932 4096
rect 6987 4136 7029 4145
rect 6987 4096 6988 4136
rect 7028 4096 7029 4136
rect 6987 4087 7029 4096
rect 7180 3968 7220 5440
rect 7275 5431 7317 5440
rect 7275 5228 7317 5237
rect 7275 5188 7276 5228
rect 7316 5188 7317 5228
rect 7275 5179 7317 5188
rect 7276 4220 7316 5179
rect 7372 4976 7412 5608
rect 7467 5480 7509 5489
rect 7467 5440 7468 5480
rect 7508 5440 7509 5480
rect 7467 5431 7509 5440
rect 7468 5346 7508 5431
rect 7564 5060 7604 6271
rect 7659 5900 7701 5909
rect 7659 5860 7660 5900
rect 7700 5860 7701 5900
rect 7659 5851 7701 5860
rect 7660 5648 7700 5851
rect 7660 5599 7700 5608
rect 7947 5648 7989 5657
rect 7947 5608 7948 5648
rect 7988 5608 7989 5648
rect 7947 5599 7989 5608
rect 7659 5480 7701 5489
rect 7659 5440 7660 5480
rect 7700 5440 7701 5480
rect 7659 5431 7701 5440
rect 7660 5237 7700 5431
rect 7659 5228 7701 5237
rect 7659 5188 7660 5228
rect 7700 5188 7701 5228
rect 7659 5179 7701 5188
rect 7756 5060 7796 5069
rect 7564 5020 7700 5060
rect 7372 4962 7604 4976
rect 7372 4936 7564 4962
rect 7467 4304 7509 4313
rect 7467 4264 7468 4304
rect 7508 4264 7509 4304
rect 7467 4255 7509 4264
rect 7372 4220 7412 4229
rect 7276 4180 7372 4220
rect 7372 4171 7412 4180
rect 7468 4220 7508 4255
rect 7564 4229 7604 4922
rect 7468 4169 7508 4180
rect 7563 4220 7605 4229
rect 7563 4180 7564 4220
rect 7604 4180 7605 4220
rect 7563 4171 7605 4180
rect 6988 3928 7220 3968
rect 6988 3548 7028 3928
rect 7083 3800 7125 3809
rect 7083 3760 7084 3800
rect 7124 3760 7125 3800
rect 7083 3751 7125 3760
rect 6988 3499 7028 3508
rect 7084 3464 7124 3751
rect 7084 3415 7124 3424
rect 7371 3464 7413 3473
rect 7371 3424 7372 3464
rect 7412 3424 7413 3464
rect 7371 3415 7413 3424
rect 7372 3330 7412 3415
rect 7467 3212 7509 3221
rect 7467 3172 7468 3212
rect 7508 3172 7509 3212
rect 7467 3163 7509 3172
rect 7275 2456 7317 2465
rect 7275 2416 7276 2456
rect 7316 2416 7317 2456
rect 7275 2407 7317 2416
rect 6740 2080 6932 2120
rect 6700 2071 6740 2080
rect 7276 1952 7316 2407
rect 7468 2129 7508 3163
rect 7660 2540 7700 5020
rect 7756 3809 7796 5020
rect 7948 4313 7988 5599
rect 7947 4304 7989 4313
rect 7947 4264 7948 4304
rect 7988 4264 7989 4304
rect 7947 4255 7989 4264
rect 7948 4136 7988 4255
rect 7852 4096 7948 4136
rect 7755 3800 7797 3809
rect 7755 3760 7756 3800
rect 7796 3760 7797 3800
rect 7755 3751 7797 3760
rect 7755 3044 7797 3053
rect 7755 3004 7756 3044
rect 7796 3004 7797 3044
rect 7755 2995 7797 3004
rect 7564 2500 7700 2540
rect 7756 2624 7796 2995
rect 7852 2633 7892 4096
rect 7948 4087 7988 4096
rect 8428 4141 8468 4150
rect 8428 3380 8468 4101
rect 8619 3968 8661 3977
rect 8619 3928 8620 3968
rect 8660 3928 8661 3968
rect 8619 3919 8661 3928
rect 8620 3834 8660 3919
rect 7948 3340 8468 3380
rect 7948 2876 7988 3340
rect 7948 2827 7988 2836
rect 7467 2120 7509 2129
rect 7467 2080 7468 2120
rect 7508 2080 7509 2120
rect 7467 2071 7509 2080
rect 7276 1709 7316 1912
rect 7275 1700 7317 1709
rect 7275 1660 7276 1700
rect 7316 1660 7317 1700
rect 7275 1651 7317 1660
rect 6603 104 6645 113
rect 1784 0 1864 80
rect 2936 0 3016 80
rect 4088 0 4168 80
rect 5240 0 5320 80
rect 6392 0 6472 80
rect 6603 64 6604 104
rect 6644 64 6645 104
rect 7564 80 7604 2500
rect 7756 1961 7796 2584
rect 7851 2624 7893 2633
rect 7851 2584 7852 2624
rect 7892 2584 7893 2624
rect 7851 2575 7893 2584
rect 8812 2213 8852 6439
rect 8907 6320 8949 6329
rect 8907 6280 8908 6320
rect 8948 6280 8949 6320
rect 8907 6271 8949 6280
rect 8908 5648 8948 6271
rect 9292 6152 9332 6616
rect 9388 6320 9428 7876
rect 9484 7253 9524 9304
rect 9964 9260 10004 9724
rect 9580 9220 10004 9260
rect 9580 8168 9620 9220
rect 10060 9185 10100 10672
rect 10155 9848 10197 9857
rect 10155 9808 10156 9848
rect 10196 9808 10197 9848
rect 10155 9799 10197 9808
rect 10156 9680 10196 9799
rect 10156 9631 10196 9640
rect 10059 9176 10101 9185
rect 10059 9136 10060 9176
rect 10100 9136 10101 9176
rect 10059 9127 10101 9136
rect 9963 9092 10005 9101
rect 9963 9052 9964 9092
rect 10004 9052 10005 9092
rect 9963 9043 10005 9052
rect 9964 8756 10004 9043
rect 10252 8849 10292 10672
rect 10347 9428 10389 9437
rect 10347 9388 10348 9428
rect 10388 9388 10389 9428
rect 10347 9379 10389 9388
rect 10348 9294 10388 9379
rect 10347 9008 10389 9017
rect 10347 8968 10348 9008
rect 10388 8968 10389 9008
rect 10347 8959 10389 8968
rect 10251 8840 10293 8849
rect 10251 8800 10252 8840
rect 10292 8800 10293 8840
rect 10251 8791 10293 8800
rect 9964 8716 10100 8756
rect 9771 8672 9813 8681
rect 9771 8632 9772 8672
rect 9812 8632 9813 8672
rect 9771 8623 9813 8632
rect 10060 8672 10100 8716
rect 10251 8714 10293 8723
rect 10251 8674 10252 8714
rect 10292 8674 10293 8714
rect 10251 8665 10293 8674
rect 9580 8119 9620 8128
rect 9772 8000 9812 8623
rect 9772 7951 9812 7960
rect 10060 7328 10100 8632
rect 10252 8588 10292 8665
rect 10252 8539 10292 8548
rect 10348 7328 10388 8959
rect 10444 7421 10484 10672
rect 10539 10016 10581 10025
rect 10539 9976 10540 10016
rect 10580 9976 10581 10016
rect 10539 9967 10581 9976
rect 10540 9428 10580 9967
rect 10540 9379 10580 9388
rect 10539 9176 10581 9185
rect 10539 9136 10540 9176
rect 10580 9136 10581 9176
rect 10539 9127 10581 9136
rect 10443 7412 10485 7421
rect 10443 7372 10444 7412
rect 10484 7372 10485 7412
rect 10443 7363 10485 7372
rect 9964 7288 10100 7328
rect 10252 7288 10388 7328
rect 9483 7244 9525 7253
rect 9483 7204 9484 7244
rect 9524 7204 9525 7244
rect 9483 7195 9525 7204
rect 9867 7244 9909 7253
rect 9867 7204 9868 7244
rect 9908 7204 9909 7244
rect 9867 7195 9909 7204
rect 9772 7160 9812 7169
rect 9484 7076 9524 7085
rect 9772 7076 9812 7120
rect 9524 7036 9812 7076
rect 9868 7160 9908 7195
rect 9484 7027 9524 7036
rect 9868 6749 9908 7120
rect 9867 6740 9909 6749
rect 9867 6700 9868 6740
rect 9908 6700 9909 6740
rect 9867 6691 9909 6700
rect 9483 6656 9525 6665
rect 9483 6616 9484 6656
rect 9524 6616 9525 6656
rect 9483 6607 9525 6616
rect 9484 6488 9524 6607
rect 9580 6497 9620 6582
rect 9484 6439 9524 6448
rect 9579 6488 9621 6497
rect 9579 6448 9580 6488
rect 9620 6448 9621 6488
rect 9579 6439 9621 6448
rect 9964 6329 10004 7288
rect 10252 7244 10292 7288
rect 10060 7204 10252 7244
rect 9868 6320 9908 6329
rect 9388 6280 9868 6320
rect 9868 6271 9908 6280
rect 9963 6320 10005 6329
rect 9963 6280 9964 6320
rect 10004 6280 10005 6320
rect 9963 6271 10005 6280
rect 9292 6112 9428 6152
rect 9291 5984 9333 5993
rect 9291 5944 9292 5984
rect 9332 5944 9333 5984
rect 9291 5935 9333 5944
rect 9292 5657 9332 5935
rect 8908 5599 8948 5608
rect 9291 5648 9333 5657
rect 9291 5608 9292 5648
rect 9332 5608 9333 5648
rect 9291 5599 9333 5608
rect 9100 5480 9140 5489
rect 9100 4985 9140 5440
rect 9099 4976 9141 4985
rect 9099 4936 9100 4976
rect 9140 4936 9141 4976
rect 9099 4927 9141 4936
rect 9099 4052 9141 4061
rect 9099 4012 9100 4052
rect 9140 4012 9141 4052
rect 9099 4003 9141 4012
rect 8907 3296 8949 3305
rect 8907 3256 8908 3296
rect 8948 3256 8949 3296
rect 8907 3247 8949 3256
rect 8908 2633 8948 3247
rect 9100 2717 9140 4003
rect 9388 3641 9428 6112
rect 9771 5816 9813 5825
rect 9771 5776 9772 5816
rect 9812 5776 9813 5816
rect 9771 5767 9813 5776
rect 9579 5648 9621 5657
rect 9579 5608 9580 5648
rect 9620 5608 9621 5648
rect 9579 5599 9621 5608
rect 9580 5321 9620 5599
rect 9772 5321 9812 5767
rect 9579 5312 9621 5321
rect 9579 5272 9580 5312
rect 9620 5272 9621 5312
rect 9579 5263 9621 5272
rect 9771 5312 9813 5321
rect 9771 5272 9772 5312
rect 9812 5272 9813 5312
rect 9771 5263 9813 5272
rect 9483 4976 9525 4985
rect 9483 4936 9484 4976
rect 9524 4936 9525 4976
rect 9483 4927 9525 4936
rect 9580 4976 9620 5263
rect 10060 5144 10100 7204
rect 10252 7195 10292 7204
rect 10348 7160 10388 7169
rect 10388 7120 10484 7160
rect 10348 7111 10388 7120
rect 10347 6992 10389 7001
rect 10347 6952 10348 6992
rect 10388 6952 10389 6992
rect 10347 6943 10389 6952
rect 10348 6656 10388 6943
rect 10348 6607 10388 6616
rect 10060 5104 10388 5144
rect 9580 4927 9620 4936
rect 9963 4976 10005 4985
rect 9963 4936 9964 4976
rect 10004 4936 10005 4976
rect 9963 4927 10005 4936
rect 10060 4976 10100 5104
rect 10060 4927 10100 4936
rect 10251 4976 10293 4985
rect 10251 4936 10252 4976
rect 10292 4936 10293 4976
rect 10251 4927 10293 4936
rect 9484 4842 9524 4927
rect 9964 4842 10004 4927
rect 9867 4472 9909 4481
rect 9867 4432 9868 4472
rect 9908 4432 9909 4472
rect 9867 4423 9909 4432
rect 9387 3632 9429 3641
rect 9387 3592 9388 3632
rect 9428 3592 9429 3632
rect 9387 3583 9429 3592
rect 9099 2708 9141 2717
rect 9099 2668 9100 2708
rect 9140 2668 9141 2708
rect 9099 2659 9141 2668
rect 8907 2624 8949 2633
rect 8907 2584 8908 2624
rect 8948 2584 8949 2624
rect 8907 2575 8949 2584
rect 9100 2624 9140 2659
rect 8811 2204 8853 2213
rect 8811 2164 8812 2204
rect 8852 2164 8853 2204
rect 8811 2155 8853 2164
rect 7755 1952 7797 1961
rect 7755 1912 7756 1952
rect 7796 1912 7797 1952
rect 7755 1903 7797 1912
rect 8523 1952 8565 1961
rect 8523 1912 8524 1952
rect 8564 1912 8565 1952
rect 8523 1903 8565 1912
rect 8908 1952 8948 2575
rect 9100 2574 9140 2584
rect 9388 2540 9428 3583
rect 9772 3464 9812 3473
rect 9772 2540 9812 3424
rect 9868 3464 9908 4423
rect 10252 3809 10292 4927
rect 10251 3800 10293 3809
rect 10251 3760 10252 3800
rect 10292 3760 10293 3800
rect 10251 3751 10293 3760
rect 9868 3415 9908 3424
rect 10252 3464 10292 3751
rect 10252 3415 10292 3424
rect 10348 3464 10388 5104
rect 10444 4985 10484 7120
rect 10540 7001 10580 9127
rect 10636 8765 10676 10672
rect 10732 9680 10772 9689
rect 10828 9680 10868 10672
rect 10772 9640 10868 9680
rect 10732 9631 10772 9640
rect 10924 9512 10964 9521
rect 10732 9472 10924 9512
rect 10635 8756 10677 8765
rect 10635 8716 10636 8756
rect 10676 8716 10677 8756
rect 10635 8707 10677 8716
rect 10732 7337 10772 9472
rect 10924 9463 10964 9472
rect 11020 8849 11060 10672
rect 11115 10604 11157 10613
rect 11115 10564 11116 10604
rect 11156 10564 11157 10604
rect 11115 10555 11157 10564
rect 11116 9017 11156 10555
rect 11115 9008 11157 9017
rect 11115 8968 11116 9008
rect 11156 8968 11157 9008
rect 11115 8959 11157 8968
rect 11212 8849 11252 10672
rect 11404 9101 11444 10672
rect 11499 10436 11541 10445
rect 11499 10396 11500 10436
rect 11540 10396 11541 10436
rect 11499 10387 11541 10396
rect 11403 9092 11445 9101
rect 11403 9052 11404 9092
rect 11444 9052 11445 9092
rect 11403 9043 11445 9052
rect 11019 8840 11061 8849
rect 11019 8800 11020 8840
rect 11060 8800 11061 8840
rect 11019 8791 11061 8800
rect 11211 8840 11253 8849
rect 11500 8840 11540 10387
rect 11211 8800 11212 8840
rect 11252 8800 11253 8840
rect 11211 8791 11253 8800
rect 11404 8800 11540 8840
rect 11404 8714 11444 8800
rect 10827 8672 10869 8681
rect 10827 8632 10828 8672
rect 10868 8632 10869 8672
rect 10827 8623 10869 8632
rect 10924 8672 10964 8683
rect 10828 8538 10868 8623
rect 10924 8597 10964 8632
rect 11308 8672 11348 8681
rect 10923 8588 10965 8597
rect 10923 8548 10924 8588
rect 10964 8548 10965 8588
rect 10923 8539 10965 8548
rect 10924 8261 10964 8539
rect 10923 8252 10965 8261
rect 10923 8212 10924 8252
rect 10964 8212 10965 8252
rect 10923 8203 10965 8212
rect 11020 8000 11060 8009
rect 11020 7589 11060 7960
rect 11308 7916 11348 8632
rect 11116 7876 11348 7916
rect 11019 7580 11061 7589
rect 11019 7540 11020 7580
rect 11060 7540 11061 7580
rect 11019 7531 11061 7540
rect 10923 7412 10965 7421
rect 10923 7372 10924 7412
rect 10964 7372 10965 7412
rect 10923 7363 10965 7372
rect 10731 7328 10773 7337
rect 10731 7288 10732 7328
rect 10772 7288 10773 7328
rect 10731 7279 10773 7288
rect 10827 7160 10869 7169
rect 10827 7120 10828 7160
rect 10868 7120 10869 7160
rect 10827 7111 10869 7120
rect 10539 6992 10581 7001
rect 10539 6952 10540 6992
rect 10580 6952 10581 6992
rect 10539 6943 10581 6952
rect 10828 6497 10868 7111
rect 10732 6488 10772 6497
rect 10732 6413 10772 6448
rect 10827 6488 10869 6497
rect 10827 6448 10828 6488
rect 10868 6448 10869 6488
rect 10827 6439 10869 6448
rect 10540 6404 10580 6413
rect 10540 5825 10580 6364
rect 10731 6404 10773 6413
rect 10731 6364 10732 6404
rect 10772 6364 10773 6404
rect 10731 6355 10773 6364
rect 10635 6320 10677 6329
rect 10635 6280 10636 6320
rect 10676 6280 10677 6320
rect 10635 6271 10677 6280
rect 10539 5816 10581 5825
rect 10539 5776 10540 5816
rect 10580 5776 10581 5816
rect 10539 5767 10581 5776
rect 10540 5648 10580 5657
rect 10636 5648 10676 6271
rect 10732 5909 10772 6355
rect 10827 6320 10869 6329
rect 10827 6280 10828 6320
rect 10868 6280 10869 6320
rect 10827 6271 10869 6280
rect 10731 5900 10773 5909
rect 10731 5860 10732 5900
rect 10772 5860 10773 5900
rect 10731 5851 10773 5860
rect 10580 5608 10676 5648
rect 10540 5599 10580 5608
rect 10443 4976 10485 4985
rect 10443 4936 10444 4976
rect 10484 4936 10485 4976
rect 10443 4927 10485 4936
rect 10540 4976 10580 4987
rect 10540 4901 10580 4936
rect 10539 4892 10581 4901
rect 10539 4852 10540 4892
rect 10580 4852 10581 4892
rect 10539 4843 10581 4852
rect 10539 4136 10581 4145
rect 10539 4096 10540 4136
rect 10580 4096 10581 4136
rect 10539 4087 10581 4096
rect 10348 3415 10388 3424
rect 10347 2960 10389 2969
rect 10347 2920 10348 2960
rect 10388 2920 10389 2960
rect 10347 2911 10389 2920
rect 10348 2624 10388 2911
rect 10540 2876 10580 4087
rect 10540 2827 10580 2836
rect 10443 2792 10485 2801
rect 10443 2752 10444 2792
rect 10484 2752 10485 2792
rect 10443 2743 10485 2752
rect 10348 2540 10388 2584
rect 9388 2500 9524 2540
rect 8908 1903 8948 1912
rect 8524 1625 8564 1903
rect 9484 1877 9524 2500
rect 9580 2500 9812 2540
rect 10252 2500 10388 2540
rect 9483 1868 9525 1877
rect 9483 1828 9484 1868
rect 9524 1828 9525 1868
rect 9483 1819 9525 1828
rect 8716 1700 8756 1709
rect 7755 1616 7797 1625
rect 7755 1576 7756 1616
rect 7796 1576 7797 1616
rect 7755 1567 7797 1576
rect 8523 1616 8565 1625
rect 8523 1576 8524 1616
rect 8564 1576 8565 1616
rect 8523 1567 8565 1576
rect 7756 1112 7796 1567
rect 8139 1196 8181 1205
rect 8139 1156 8140 1196
rect 8180 1156 8181 1196
rect 8139 1147 8181 1156
rect 7756 1063 7796 1072
rect 8140 1112 8180 1147
rect 8716 1121 8756 1660
rect 9387 1280 9429 1289
rect 9387 1240 9388 1280
rect 9428 1240 9429 1280
rect 9387 1231 9429 1240
rect 9580 1280 9620 2500
rect 10155 1952 10197 1961
rect 10155 1912 10156 1952
rect 10196 1912 10197 1952
rect 10155 1903 10197 1912
rect 10156 1818 10196 1903
rect 10252 1289 10292 2500
rect 10444 1952 10484 2743
rect 10539 1952 10581 1961
rect 10444 1912 10540 1952
rect 10580 1912 10581 1952
rect 10539 1903 10581 1912
rect 10540 1818 10580 1903
rect 10636 1877 10676 5608
rect 10828 5564 10868 6271
rect 10924 5900 10964 7363
rect 11020 6497 11060 7531
rect 11116 7076 11156 7876
rect 11404 7832 11444 8674
rect 11499 8672 11541 8681
rect 11499 8632 11500 8672
rect 11540 8632 11541 8672
rect 11499 8623 11541 8632
rect 11500 8168 11540 8623
rect 11500 8119 11540 8128
rect 11404 7792 11540 7832
rect 11212 7748 11252 7757
rect 11252 7708 11396 7748
rect 11212 7699 11252 7708
rect 11356 7202 11396 7708
rect 11500 7421 11540 7792
rect 11499 7412 11541 7421
rect 11499 7372 11500 7412
rect 11540 7372 11541 7412
rect 11499 7363 11541 7372
rect 11499 7244 11541 7253
rect 11499 7204 11500 7244
rect 11540 7204 11541 7244
rect 11499 7195 11541 7204
rect 11356 7153 11396 7162
rect 11500 7076 11540 7195
rect 11116 7036 11348 7076
rect 11019 6488 11061 6497
rect 11019 6448 11020 6488
rect 11060 6448 11061 6488
rect 11019 6439 11061 6448
rect 10924 5851 10964 5860
rect 11019 5900 11061 5909
rect 11019 5860 11020 5900
rect 11060 5860 11061 5900
rect 11019 5851 11061 5860
rect 11020 5657 11060 5851
rect 11116 5732 11156 5741
rect 11156 5692 11252 5732
rect 11116 5683 11156 5692
rect 11019 5648 11061 5657
rect 11019 5608 11020 5648
rect 11060 5608 11061 5648
rect 11019 5599 11061 5608
rect 10828 5524 10964 5564
rect 10732 5480 10772 5489
rect 10772 5440 10868 5480
rect 10732 5431 10772 5440
rect 10828 5228 10868 5440
rect 10924 5312 10964 5524
rect 10924 5272 11156 5312
rect 10828 5188 11060 5228
rect 11020 4971 11060 5188
rect 11116 4976 11156 5272
rect 11212 5144 11252 5692
rect 11212 5095 11252 5104
rect 11116 4936 11252 4976
rect 11020 4922 11060 4931
rect 10827 4892 10869 4901
rect 10827 4852 10828 4892
rect 10868 4852 10869 4892
rect 10827 4843 10869 4852
rect 10828 3464 10868 4843
rect 11019 4640 11061 4649
rect 11019 4600 11020 4640
rect 11060 4600 11061 4640
rect 11019 4591 11061 4600
rect 11020 4229 11060 4591
rect 11019 4220 11061 4229
rect 11019 4180 11020 4220
rect 11060 4180 11061 4220
rect 11019 4171 11061 4180
rect 10923 4136 10965 4145
rect 10923 4096 10924 4136
rect 10964 4096 10965 4136
rect 10923 4087 10965 4096
rect 11020 4136 11060 4171
rect 10924 4002 10964 4087
rect 11020 4086 11060 4096
rect 10828 3415 10868 3424
rect 11019 3128 11061 3137
rect 11019 3088 11020 3128
rect 11060 3088 11061 3128
rect 11019 3079 11061 3088
rect 11020 2624 11060 3079
rect 11212 2969 11252 4936
rect 11308 4220 11348 7036
rect 11500 7027 11540 7036
rect 11499 6908 11541 6917
rect 11499 6868 11500 6908
rect 11540 6868 11541 6908
rect 11499 6859 11541 6868
rect 11404 4220 11444 4229
rect 11308 4180 11404 4220
rect 11308 4061 11348 4180
rect 11404 4171 11444 4180
rect 11500 4220 11540 6859
rect 11596 5060 11636 10672
rect 11691 9092 11733 9101
rect 11691 9052 11692 9092
rect 11732 9052 11733 9092
rect 11691 9043 11733 9052
rect 11692 8504 11732 9043
rect 11788 8849 11828 10672
rect 11787 8840 11829 8849
rect 11787 8800 11788 8840
rect 11828 8800 11829 8840
rect 11787 8791 11829 8800
rect 11884 8681 11924 8766
rect 11883 8672 11925 8681
rect 11883 8632 11884 8672
rect 11924 8632 11925 8672
rect 11883 8623 11925 8632
rect 11692 8464 11924 8504
rect 11884 8168 11924 8464
rect 11884 8119 11924 8128
rect 11787 8084 11829 8093
rect 11787 8044 11788 8084
rect 11828 8044 11829 8084
rect 11787 8035 11829 8044
rect 11691 7916 11733 7925
rect 11691 7876 11692 7916
rect 11732 7876 11733 7916
rect 11691 7867 11733 7876
rect 11692 7782 11732 7867
rect 11692 7412 11732 7421
rect 11788 7412 11828 8035
rect 11732 7372 11828 7412
rect 11883 7412 11925 7421
rect 11883 7372 11884 7412
rect 11924 7372 11925 7412
rect 11692 7363 11732 7372
rect 11883 7363 11925 7372
rect 11884 7244 11924 7363
rect 11884 7195 11924 7204
rect 11980 7076 12020 10672
rect 12172 9689 12212 10672
rect 12171 9680 12213 9689
rect 12171 9640 12172 9680
rect 12212 9640 12213 9680
rect 12171 9631 12213 9640
rect 12172 9512 12212 9521
rect 12172 9017 12212 9472
rect 12364 9428 12404 10672
rect 12364 9388 12500 9428
rect 12364 9260 12404 9269
rect 12171 9008 12213 9017
rect 12171 8968 12172 9008
rect 12212 8968 12213 9008
rect 12171 8959 12213 8968
rect 12364 8686 12404 9220
rect 12267 8672 12309 8681
rect 12267 8632 12268 8672
rect 12308 8632 12309 8672
rect 12364 8637 12404 8646
rect 12267 8623 12309 8632
rect 12076 7916 12116 7925
rect 12076 7589 12116 7876
rect 12075 7580 12117 7589
rect 12075 7540 12076 7580
rect 12116 7540 12117 7580
rect 12075 7531 12117 7540
rect 12075 7412 12117 7421
rect 12075 7372 12076 7412
rect 12116 7372 12117 7412
rect 12075 7363 12117 7372
rect 11884 7036 12020 7076
rect 11596 5020 11828 5060
rect 11692 4892 11732 4901
rect 11500 4145 11540 4180
rect 11596 4852 11692 4892
rect 11499 4136 11541 4145
rect 11499 4096 11500 4136
rect 11540 4096 11541 4136
rect 11499 4087 11541 4096
rect 11307 4052 11349 4061
rect 11500 4056 11540 4087
rect 11307 4012 11308 4052
rect 11348 4012 11349 4052
rect 11307 4003 11349 4012
rect 11500 3632 11540 3641
rect 11596 3632 11636 4852
rect 11692 4843 11732 4852
rect 11788 4733 11828 5020
rect 11884 4808 11924 7036
rect 11979 6488 12021 6497
rect 11979 6448 11980 6488
rect 12020 6448 12021 6488
rect 11979 6439 12021 6448
rect 11980 6354 12020 6439
rect 11979 6236 12021 6245
rect 11979 6196 11980 6236
rect 12020 6196 12021 6236
rect 11979 6187 12021 6196
rect 11884 4759 11924 4768
rect 11787 4724 11829 4733
rect 11980 4724 12020 6187
rect 12076 4892 12116 7363
rect 12171 6572 12213 6581
rect 12171 6532 12172 6572
rect 12212 6532 12213 6572
rect 12171 6523 12213 6532
rect 12172 6438 12212 6523
rect 12268 6329 12308 8623
rect 12363 8000 12405 8009
rect 12363 7960 12364 8000
rect 12404 7960 12405 8000
rect 12363 7951 12405 7960
rect 12267 6320 12309 6329
rect 12267 6280 12268 6320
rect 12308 6280 12309 6320
rect 12267 6271 12309 6280
rect 12267 5060 12309 5069
rect 12267 5020 12268 5060
rect 12308 5020 12309 5060
rect 12267 5011 12309 5020
rect 12268 4892 12308 5011
rect 12076 4852 12212 4892
rect 11787 4684 11788 4724
rect 11828 4684 11829 4724
rect 11787 4675 11829 4684
rect 11979 4684 12020 4724
rect 12075 4724 12117 4733
rect 12075 4684 12076 4724
rect 12116 4684 12117 4724
rect 11979 4640 12019 4684
rect 12075 4675 12117 4684
rect 11979 4600 12020 4640
rect 11980 4136 12020 4600
rect 12076 4590 12116 4675
rect 12172 4481 12212 4852
rect 12268 4843 12308 4852
rect 12171 4472 12213 4481
rect 12171 4432 12172 4472
rect 12212 4432 12213 4472
rect 12171 4423 12213 4432
rect 11980 4087 12020 4096
rect 12075 3884 12117 3893
rect 12075 3844 12076 3884
rect 12116 3844 12117 3884
rect 12075 3835 12117 3844
rect 11540 3592 11636 3632
rect 11500 3583 11540 3592
rect 11308 3450 11348 3459
rect 11211 2960 11253 2969
rect 11211 2920 11212 2960
rect 11252 2920 11253 2960
rect 11211 2911 11253 2920
rect 11212 2717 11252 2911
rect 11211 2708 11253 2717
rect 11211 2668 11212 2708
rect 11252 2668 11253 2708
rect 11211 2659 11253 2668
rect 11020 2129 11060 2584
rect 11019 2120 11061 2129
rect 11019 2080 11020 2120
rect 11060 2080 11061 2120
rect 11019 2071 11061 2080
rect 10635 1868 10677 1877
rect 10635 1828 10636 1868
rect 10676 1828 10677 1868
rect 10635 1819 10677 1828
rect 10348 1700 10388 1709
rect 9580 1231 9620 1240
rect 10251 1280 10293 1289
rect 10251 1240 10252 1280
rect 10292 1240 10293 1280
rect 10251 1231 10293 1240
rect 8140 1061 8180 1072
rect 8715 1112 8757 1121
rect 8715 1072 8716 1112
rect 8756 1072 8757 1112
rect 8715 1063 8757 1072
rect 9388 1112 9428 1231
rect 9388 1063 9428 1072
rect 9772 1112 9812 1121
rect 9772 953 9812 1072
rect 9867 1112 9909 1121
rect 9867 1072 9868 1112
rect 9908 1072 9909 1112
rect 9867 1063 9909 1072
rect 7947 944 7989 953
rect 7947 904 7948 944
rect 7988 904 7989 944
rect 7947 895 7989 904
rect 8715 944 8757 953
rect 8715 904 8716 944
rect 8756 904 8757 944
rect 8715 895 8757 904
rect 9771 944 9813 953
rect 9771 904 9772 944
rect 9812 904 9813 944
rect 9771 895 9813 904
rect 7948 810 7988 895
rect 8716 80 8756 895
rect 9868 80 9908 1063
rect 10348 113 10388 1660
rect 11019 1280 11061 1289
rect 11019 1240 11020 1280
rect 11060 1240 11061 1280
rect 11019 1231 11061 1240
rect 11212 1280 11252 1289
rect 11308 1280 11348 3410
rect 11403 2876 11445 2885
rect 11403 2836 11404 2876
rect 11444 2836 11445 2876
rect 11403 2827 11445 2836
rect 11404 2465 11444 2827
rect 11403 2456 11445 2465
rect 11403 2416 11404 2456
rect 11444 2416 11445 2456
rect 11403 2407 11445 2416
rect 11252 1240 11348 1280
rect 11212 1231 11252 1240
rect 11020 1112 11060 1231
rect 11020 1063 11060 1072
rect 11404 1112 11444 2407
rect 11788 1952 11828 1963
rect 12076 1952 12116 3835
rect 12267 3464 12309 3473
rect 12267 3424 12268 3464
rect 12308 3424 12309 3464
rect 12267 3415 12309 3424
rect 12268 3330 12308 3415
rect 12267 2708 12309 2717
rect 12267 2668 12268 2708
rect 12308 2668 12309 2708
rect 12267 2659 12309 2668
rect 12268 2624 12308 2659
rect 12268 2573 12308 2584
rect 12172 1952 12212 1961
rect 12076 1912 12172 1952
rect 11788 1877 11828 1912
rect 12172 1903 12212 1912
rect 11787 1868 11829 1877
rect 11787 1828 11788 1868
rect 11828 1828 11829 1868
rect 11787 1819 11829 1828
rect 11404 1063 11444 1072
rect 11980 1700 12020 1709
rect 11980 188 12020 1660
rect 12364 1121 12404 7951
rect 12460 7664 12500 9388
rect 12556 8849 12596 10672
rect 12555 8840 12597 8849
rect 12555 8800 12556 8840
rect 12596 8800 12597 8840
rect 12555 8791 12597 8800
rect 12556 8504 12596 8513
rect 12556 7925 12596 8464
rect 12748 8168 12788 10672
rect 12940 9185 12980 10672
rect 13132 10193 13172 10672
rect 13131 10184 13173 10193
rect 13131 10144 13132 10184
rect 13172 10144 13173 10184
rect 13131 10135 13173 10144
rect 13131 9512 13173 9521
rect 13131 9472 13132 9512
rect 13172 9472 13173 9512
rect 13131 9463 13173 9472
rect 12939 9176 12981 9185
rect 12939 9136 12940 9176
rect 12980 9136 12981 9176
rect 12939 9127 12981 9136
rect 12939 9008 12981 9017
rect 12939 8968 12940 9008
rect 12980 8968 12981 9008
rect 12939 8959 12981 8968
rect 12748 8128 12884 8168
rect 12747 8000 12789 8009
rect 12747 7960 12748 8000
rect 12788 7960 12789 8000
rect 12747 7951 12789 7960
rect 12555 7916 12597 7925
rect 12555 7876 12556 7916
rect 12596 7876 12597 7916
rect 12555 7867 12597 7876
rect 12748 7866 12788 7951
rect 12460 7624 12692 7664
rect 12555 6740 12597 6749
rect 12555 6700 12556 6740
rect 12596 6700 12597 6740
rect 12555 6691 12597 6700
rect 12459 6572 12501 6581
rect 12459 6532 12460 6572
rect 12500 6532 12501 6572
rect 12459 6523 12501 6532
rect 12460 6488 12500 6523
rect 12460 6437 12500 6448
rect 12556 6488 12596 6691
rect 12556 6439 12596 6448
rect 12459 5984 12501 5993
rect 12459 5944 12460 5984
rect 12500 5944 12501 5984
rect 12459 5935 12501 5944
rect 12460 4985 12500 5935
rect 12652 5900 12692 7624
rect 12747 7244 12789 7253
rect 12747 7204 12748 7244
rect 12788 7204 12789 7244
rect 12747 7195 12789 7204
rect 12748 7110 12788 7195
rect 12844 5900 12884 8128
rect 12940 7412 12980 8959
rect 13035 8672 13077 8681
rect 13035 8632 13036 8672
rect 13076 8632 13077 8672
rect 13035 8623 13077 8632
rect 13036 8538 13076 8623
rect 13132 7421 13172 9463
rect 13324 9101 13364 10672
rect 13323 9092 13365 9101
rect 13323 9052 13324 9092
rect 13364 9052 13365 9092
rect 13323 9043 13365 9052
rect 13516 8840 13556 10672
rect 13708 8924 13748 10672
rect 13900 9689 13940 10672
rect 13899 9680 13941 9689
rect 13899 9640 13900 9680
rect 13940 9640 13941 9680
rect 13899 9631 13941 9640
rect 13708 8884 13844 8924
rect 13516 8800 13748 8840
rect 12940 7363 12980 7372
rect 13131 7412 13173 7421
rect 13708 7412 13748 8800
rect 13804 8513 13844 8884
rect 14092 8849 14132 10672
rect 14187 9680 14229 9689
rect 14187 9640 14188 9680
rect 14228 9640 14229 9680
rect 14187 9631 14229 9640
rect 14188 9546 14228 9631
rect 14284 9017 14324 10672
rect 14380 9428 14420 9437
rect 14283 9008 14325 9017
rect 14283 8968 14284 9008
rect 14324 8968 14325 9008
rect 14283 8959 14325 8968
rect 14091 8840 14133 8849
rect 14091 8800 14092 8840
rect 14132 8800 14133 8840
rect 14091 8791 14133 8800
rect 14284 8672 14324 8681
rect 13803 8504 13845 8513
rect 13803 8464 13804 8504
rect 13844 8464 13845 8504
rect 13803 8455 13845 8464
rect 14284 8345 14324 8632
rect 13995 8336 14037 8345
rect 13995 8296 13996 8336
rect 14036 8296 14037 8336
rect 13995 8287 14037 8296
rect 14283 8336 14325 8345
rect 14283 8296 14284 8336
rect 14324 8296 14325 8336
rect 14283 8287 14325 8296
rect 13996 8000 14036 8287
rect 14091 8252 14133 8261
rect 14091 8212 14092 8252
rect 14132 8212 14133 8252
rect 14091 8203 14133 8212
rect 14092 8009 14132 8203
rect 14380 8168 14420 9388
rect 14476 8849 14516 10672
rect 14475 8840 14517 8849
rect 14475 8800 14476 8840
rect 14516 8800 14517 8840
rect 14668 8840 14708 10672
rect 14860 9605 14900 10672
rect 14859 9596 14901 9605
rect 14859 9556 14860 9596
rect 14900 9556 14901 9596
rect 14859 9547 14901 9556
rect 14955 9512 14997 9521
rect 14955 9472 14956 9512
rect 14996 9472 14997 9512
rect 14955 9463 14997 9472
rect 14956 9378 14996 9463
rect 15052 9185 15092 10672
rect 15244 9689 15284 10672
rect 15243 9680 15285 9689
rect 15243 9640 15244 9680
rect 15284 9640 15285 9680
rect 15243 9631 15285 9640
rect 15051 9176 15093 9185
rect 15051 9136 15052 9176
rect 15092 9136 15093 9176
rect 15051 9127 15093 9136
rect 15436 8849 15476 10672
rect 15628 8849 15668 10672
rect 15820 10109 15860 10672
rect 15819 10100 15861 10109
rect 15819 10060 15820 10100
rect 15860 10060 15861 10100
rect 15819 10051 15861 10060
rect 16012 8849 16052 10672
rect 16204 9857 16244 10672
rect 16203 9848 16245 9857
rect 16203 9808 16204 9848
rect 16244 9808 16245 9848
rect 16203 9799 16245 9808
rect 16396 9689 16436 10672
rect 16395 9680 16437 9689
rect 16395 9640 16396 9680
rect 16436 9640 16437 9680
rect 16395 9631 16437 9640
rect 16204 9512 16244 9521
rect 15435 8840 15477 8849
rect 14668 8800 14996 8840
rect 14475 8791 14517 8800
rect 14764 8672 14804 8681
rect 14476 8588 14516 8597
rect 14764 8588 14804 8632
rect 14859 8672 14901 8681
rect 14859 8632 14860 8672
rect 14900 8632 14901 8672
rect 14859 8623 14901 8632
rect 14516 8548 14804 8588
rect 14476 8539 14516 8548
rect 14860 8538 14900 8623
rect 14380 8128 14804 8168
rect 14188 8084 14228 8093
rect 14228 8044 14612 8084
rect 14188 8035 14228 8044
rect 13996 7951 14036 7960
rect 14091 8000 14133 8009
rect 14091 7960 14092 8000
rect 14132 7960 14133 8000
rect 14091 7951 14133 7960
rect 14572 8000 14612 8044
rect 14572 7951 14612 7960
rect 14667 8000 14709 8009
rect 14667 7960 14668 8000
rect 14708 7960 14709 8000
rect 14667 7951 14709 7960
rect 14668 7866 14708 7951
rect 13131 7372 13132 7412
rect 13172 7372 13364 7412
rect 13131 7363 13173 7372
rect 12939 7244 12981 7253
rect 12939 7204 12940 7244
rect 12980 7204 12981 7244
rect 12939 7195 12981 7204
rect 12940 6488 12980 7195
rect 13131 6992 13173 7001
rect 13131 6952 13132 6992
rect 13172 6952 13173 6992
rect 13131 6943 13173 6952
rect 12940 6439 12980 6448
rect 13035 6404 13077 6413
rect 13035 6364 13036 6404
rect 13076 6364 13077 6404
rect 13035 6355 13077 6364
rect 13036 6270 13076 6355
rect 12652 5860 12788 5900
rect 12652 5732 12692 5741
rect 12459 4976 12501 4985
rect 12459 4936 12460 4976
rect 12500 4936 12501 4976
rect 12459 4927 12501 4936
rect 12460 4842 12500 4927
rect 12555 4640 12597 4649
rect 12555 4600 12556 4640
rect 12596 4600 12597 4640
rect 12555 4591 12597 4600
rect 12460 4141 12500 4150
rect 12460 2876 12500 4101
rect 12556 3893 12596 4591
rect 12652 4052 12692 5692
rect 12652 4003 12692 4012
rect 12555 3884 12597 3893
rect 12555 3844 12556 3884
rect 12596 3844 12597 3884
rect 12555 3835 12597 3844
rect 12748 2876 12788 5860
rect 12844 5851 12884 5860
rect 13036 5648 13076 5657
rect 13132 5648 13172 6943
rect 13076 5608 13172 5648
rect 13036 5599 13076 5608
rect 13132 4136 13172 4145
rect 13132 3725 13172 4096
rect 13228 4136 13268 4147
rect 13228 4061 13268 4096
rect 13227 4052 13269 4061
rect 13227 4012 13228 4052
rect 13268 4012 13269 4052
rect 13227 4003 13269 4012
rect 13131 3716 13173 3725
rect 13131 3676 13132 3716
rect 13172 3676 13173 3716
rect 13131 3667 13173 3676
rect 12844 2876 12884 2885
rect 12748 2836 12844 2876
rect 12460 2827 12500 2836
rect 12844 2827 12884 2836
rect 13035 2708 13077 2717
rect 13035 2668 13036 2708
rect 13076 2668 13077 2708
rect 13035 2659 13077 2668
rect 13036 2574 13076 2659
rect 12651 1868 12693 1877
rect 12651 1828 12652 1868
rect 12692 1828 12693 1868
rect 12651 1819 12693 1828
rect 12363 1112 12405 1121
rect 12363 1072 12364 1112
rect 12404 1072 12405 1112
rect 12363 1063 12405 1072
rect 12652 1112 12692 1819
rect 12652 1063 12692 1072
rect 13036 1112 13076 1123
rect 13036 1037 13076 1072
rect 13324 1037 13364 7372
rect 13708 7363 13748 7372
rect 14379 7412 14421 7421
rect 14379 7372 14380 7412
rect 14420 7372 14421 7412
rect 14379 7363 14421 7372
rect 13900 7244 13940 7253
rect 13940 7204 14228 7244
rect 13900 7195 13940 7204
rect 13515 7160 13557 7169
rect 13515 7120 13516 7160
rect 13556 7120 13557 7160
rect 13515 7111 13557 7120
rect 13516 6581 13556 7111
rect 14188 6656 14228 7204
rect 14380 7160 14420 7363
rect 14380 7085 14420 7120
rect 14379 7076 14421 7085
rect 14379 7036 14380 7076
rect 14420 7036 14421 7076
rect 14379 7027 14421 7036
rect 14380 6996 14420 7027
rect 14188 6607 14228 6616
rect 14668 6656 14708 6665
rect 14764 6656 14804 8128
rect 14708 6616 14804 6656
rect 14668 6607 14708 6616
rect 13515 6572 13557 6581
rect 13515 6532 13516 6572
rect 13556 6532 13557 6572
rect 13515 6523 13557 6532
rect 13516 6488 13556 6523
rect 13516 6438 13556 6448
rect 13707 6488 13749 6497
rect 13707 6448 13708 6488
rect 13748 6448 13749 6488
rect 14187 6488 14229 6497
rect 13707 6439 13749 6448
rect 13996 6474 14036 6483
rect 13708 5657 13748 6439
rect 14187 6448 14188 6488
rect 14228 6448 14229 6488
rect 14187 6439 14229 6448
rect 14475 6488 14517 6497
rect 14475 6448 14476 6488
rect 14516 6448 14517 6488
rect 14475 6439 14517 6448
rect 14812 6446 14852 6455
rect 13803 6404 13845 6413
rect 13803 6364 13804 6404
rect 13844 6364 13845 6404
rect 13803 6355 13845 6364
rect 13707 5648 13749 5657
rect 13707 5608 13708 5648
rect 13748 5608 13749 5648
rect 13707 5599 13749 5608
rect 13708 4976 13748 5599
rect 13708 4927 13748 4936
rect 13804 4901 13844 6355
rect 13900 5060 13940 5069
rect 13996 5060 14036 6434
rect 13940 5020 14036 5060
rect 13900 5011 13940 5020
rect 13803 4892 13845 4901
rect 13803 4852 13804 4892
rect 13844 4852 13845 4892
rect 13803 4843 13845 4852
rect 13804 4724 13844 4843
rect 13708 4684 13844 4724
rect 13708 4220 13748 4684
rect 13803 4388 13845 4397
rect 13803 4348 13804 4388
rect 13844 4348 13845 4388
rect 13803 4339 13845 4348
rect 13708 4171 13748 4180
rect 13611 4136 13653 4145
rect 13611 4096 13612 4136
rect 13652 4096 13653 4136
rect 13611 4087 13653 4096
rect 13612 4002 13652 4087
rect 13707 3716 13749 3725
rect 13707 3676 13708 3716
rect 13748 3676 13749 3716
rect 13707 3667 13749 3676
rect 13708 3632 13748 3667
rect 13708 3581 13748 3592
rect 13515 3464 13557 3473
rect 13515 3424 13516 3464
rect 13556 3424 13557 3464
rect 13515 3415 13557 3424
rect 13516 3330 13556 3415
rect 13804 2801 13844 4339
rect 14188 4136 14228 6439
rect 14476 5900 14516 6439
rect 14812 6404 14852 6406
rect 14476 5851 14516 5860
rect 14668 6364 14852 6404
rect 14668 5900 14708 6364
rect 14859 5984 14901 5993
rect 14859 5944 14860 5984
rect 14900 5944 14901 5984
rect 14859 5935 14901 5944
rect 14668 5851 14708 5860
rect 14860 5657 14900 5935
rect 14283 5648 14325 5657
rect 14283 5608 14284 5648
rect 14324 5608 14325 5648
rect 14283 5599 14325 5608
rect 14859 5648 14901 5657
rect 14859 5608 14860 5648
rect 14900 5608 14901 5648
rect 14859 5599 14901 5608
rect 14284 5514 14324 5599
rect 14956 5480 14996 8800
rect 15435 8800 15436 8840
rect 15476 8800 15477 8840
rect 15435 8791 15477 8800
rect 15627 8840 15669 8849
rect 15627 8800 15628 8840
rect 15668 8800 15669 8840
rect 15627 8791 15669 8800
rect 16011 8840 16053 8849
rect 16011 8800 16012 8840
rect 16052 8800 16053 8840
rect 16011 8791 16053 8800
rect 15244 8672 15284 8681
rect 15244 8513 15284 8632
rect 15340 8672 15380 8681
rect 15243 8504 15285 8513
rect 15243 8464 15244 8504
rect 15284 8464 15285 8504
rect 15243 8455 15285 8464
rect 15147 8168 15189 8177
rect 15147 8128 15148 8168
rect 15188 8128 15189 8168
rect 15147 8119 15189 8128
rect 15148 8000 15188 8119
rect 15148 7951 15188 7960
rect 15052 7916 15092 7925
rect 15052 7757 15092 7876
rect 15051 7748 15093 7757
rect 15051 7708 15052 7748
rect 15092 7708 15093 7748
rect 15051 7699 15093 7708
rect 15244 7673 15284 8455
rect 15340 8261 15380 8632
rect 15819 8672 15861 8681
rect 15819 8632 15820 8672
rect 15860 8632 15861 8672
rect 15819 8623 15861 8632
rect 15820 8538 15860 8623
rect 16204 8345 16244 9472
rect 16491 9428 16533 9437
rect 16491 9388 16492 9428
rect 16532 9388 16533 9428
rect 16491 9379 16533 9388
rect 16396 9260 16436 9269
rect 16300 9220 16396 9260
rect 16300 8686 16340 9220
rect 16396 9211 16436 9220
rect 16300 8637 16340 8646
rect 16492 8588 16532 9379
rect 16492 8539 16532 8548
rect 15723 8336 15765 8345
rect 15723 8296 15724 8336
rect 15764 8296 15765 8336
rect 15723 8287 15765 8296
rect 16203 8336 16245 8345
rect 16203 8296 16204 8336
rect 16244 8296 16245 8336
rect 16203 8287 16245 8296
rect 15339 8252 15381 8261
rect 15339 8212 15340 8252
rect 15380 8212 15381 8252
rect 15339 8203 15381 8212
rect 15340 7841 15380 8203
rect 15628 7958 15668 7967
rect 15628 7841 15668 7918
rect 15339 7832 15381 7841
rect 15627 7832 15669 7841
rect 15339 7792 15340 7832
rect 15380 7792 15381 7832
rect 15339 7783 15381 7792
rect 15532 7792 15628 7832
rect 15668 7792 15669 7832
rect 15243 7664 15285 7673
rect 15243 7624 15244 7664
rect 15284 7624 15285 7664
rect 15243 7615 15285 7624
rect 15339 6572 15381 6581
rect 15339 6532 15340 6572
rect 15380 6532 15381 6572
rect 15339 6523 15381 6532
rect 15340 6488 15380 6523
rect 15340 6437 15380 6448
rect 15532 5909 15572 7792
rect 15627 7783 15669 7792
rect 15628 7698 15668 7783
rect 15628 7160 15668 7169
rect 15724 7160 15764 8287
rect 16300 8084 16340 8093
rect 16108 7986 16148 7995
rect 16108 7496 16148 7946
rect 16300 7925 16340 8044
rect 16299 7916 16341 7925
rect 16299 7876 16300 7916
rect 16340 7876 16341 7916
rect 16299 7867 16341 7876
rect 15820 7456 16148 7496
rect 15820 7412 15860 7456
rect 15820 7363 15860 7372
rect 15915 7244 15957 7253
rect 15915 7204 15916 7244
rect 15956 7204 15957 7244
rect 15915 7195 15957 7204
rect 15668 7120 15764 7160
rect 15531 5900 15573 5909
rect 15531 5860 15532 5900
rect 15572 5860 15573 5900
rect 15531 5851 15573 5860
rect 14668 5440 14996 5480
rect 14668 4808 14708 5440
rect 14668 4759 14708 4768
rect 14860 4892 14900 4901
rect 14188 4087 14228 4096
rect 14668 4141 14708 4150
rect 14283 3548 14325 3557
rect 14283 3508 14284 3548
rect 14324 3508 14325 3548
rect 14283 3499 14325 3508
rect 13899 3464 13941 3473
rect 13899 3424 13900 3464
rect 13940 3424 13941 3464
rect 13899 3415 13941 3424
rect 13900 3330 13940 3415
rect 13803 2792 13845 2801
rect 13803 2752 13804 2792
rect 13844 2752 13845 2792
rect 13803 2743 13845 2752
rect 13420 1952 13460 1963
rect 13420 1877 13460 1912
rect 13804 1952 13844 2743
rect 13804 1903 13844 1912
rect 13419 1868 13461 1877
rect 13419 1828 13420 1868
rect 13460 1828 13461 1868
rect 13419 1819 13461 1828
rect 13612 1700 13652 1709
rect 13035 1028 13077 1037
rect 13035 988 13036 1028
rect 13076 988 13077 1028
rect 13035 979 13077 988
rect 13323 1028 13365 1037
rect 13323 988 13324 1028
rect 13364 988 13365 1028
rect 13323 979 13365 988
rect 12844 944 12884 953
rect 11980 148 12212 188
rect 10347 104 10389 113
rect 6603 55 6645 64
rect 7544 0 7624 80
rect 8696 0 8776 80
rect 9848 0 9928 80
rect 10347 64 10348 104
rect 10388 64 10389 104
rect 11019 104 11061 113
rect 11019 80 11020 104
rect 10347 55 10389 64
rect 11000 64 11020 80
rect 11060 80 11061 104
rect 12172 80 12212 148
rect 12844 113 12884 904
rect 13036 701 13076 979
rect 13612 953 13652 1660
rect 14284 1112 14324 3499
rect 14380 2633 14420 2719
rect 14379 2624 14421 2633
rect 14379 2584 14380 2624
rect 14420 2584 14421 2624
rect 14379 2575 14421 2584
rect 14380 2213 14420 2575
rect 14668 2540 14708 4101
rect 14860 4052 14900 4852
rect 14860 4003 14900 4012
rect 15436 4136 15476 4145
rect 15340 3632 15380 3641
rect 15436 3632 15476 4096
rect 15532 4136 15572 4145
rect 15532 3809 15572 4096
rect 15531 3800 15573 3809
rect 15531 3760 15532 3800
rect 15572 3760 15573 3800
rect 15531 3751 15573 3760
rect 15380 3592 15476 3632
rect 15340 3583 15380 3592
rect 15628 3557 15668 7120
rect 15916 6488 15956 7195
rect 15820 6404 15860 6415
rect 15916 6413 15956 6448
rect 16012 7160 16052 7169
rect 15820 6329 15860 6364
rect 15915 6404 15957 6413
rect 15915 6364 15916 6404
rect 15956 6364 15957 6404
rect 15915 6355 15957 6364
rect 15819 6320 15861 6329
rect 15916 6324 15956 6355
rect 15819 6280 15820 6320
rect 15860 6280 15861 6320
rect 15819 6271 15861 6280
rect 16012 6245 16052 7120
rect 16491 6572 16533 6581
rect 16491 6532 16492 6572
rect 16532 6532 16533 6572
rect 16491 6523 16533 6532
rect 16300 6488 16340 6497
rect 16204 6448 16300 6488
rect 16011 6236 16053 6245
rect 16011 6196 16012 6236
rect 16052 6196 16053 6236
rect 16011 6187 16053 6196
rect 16012 5153 16052 6187
rect 16107 5648 16149 5657
rect 16107 5608 16108 5648
rect 16148 5608 16149 5648
rect 16107 5599 16149 5608
rect 16108 5405 16148 5599
rect 16107 5396 16149 5405
rect 16107 5356 16108 5396
rect 16148 5356 16149 5396
rect 16107 5347 16149 5356
rect 16011 5144 16053 5153
rect 16011 5104 16012 5144
rect 16052 5104 16053 5144
rect 16011 5095 16053 5104
rect 15916 4136 15956 4145
rect 15147 3548 15189 3557
rect 15147 3508 15148 3548
rect 15188 3508 15189 3548
rect 15147 3499 15189 3508
rect 15627 3548 15669 3557
rect 15627 3508 15628 3548
rect 15668 3508 15669 3548
rect 15627 3499 15669 3508
rect 15148 3464 15188 3499
rect 15148 3413 15188 3424
rect 15531 3464 15573 3473
rect 15531 3424 15532 3464
rect 15572 3424 15573 3464
rect 15531 3415 15573 3424
rect 15532 3330 15572 3415
rect 15916 3305 15956 4096
rect 16012 4136 16052 4145
rect 16204 4136 16244 6448
rect 16300 6439 16340 6448
rect 16395 6488 16437 6497
rect 16395 6448 16396 6488
rect 16436 6448 16437 6488
rect 16395 6439 16437 6448
rect 16396 6354 16436 6439
rect 16299 5732 16341 5741
rect 16299 5692 16300 5732
rect 16340 5692 16341 5732
rect 16299 5683 16341 5692
rect 16300 5648 16340 5683
rect 16300 5597 16340 5608
rect 16052 4096 16244 4136
rect 16492 4136 16532 6523
rect 16588 4808 16628 10672
rect 16780 8849 16820 10672
rect 16972 10529 17012 10672
rect 16971 10520 17013 10529
rect 16971 10480 16972 10520
rect 17012 10480 17013 10520
rect 16971 10471 17013 10480
rect 17164 9941 17204 10672
rect 17163 9932 17205 9941
rect 17163 9892 17164 9932
rect 17204 9892 17205 9932
rect 17163 9883 17205 9892
rect 17068 9680 17108 9689
rect 17356 9680 17396 10672
rect 17108 9640 17396 9680
rect 17068 9631 17108 9640
rect 16875 9428 16917 9437
rect 16875 9388 16876 9428
rect 16916 9388 16917 9428
rect 16875 9379 16917 9388
rect 16876 9294 16916 9379
rect 16971 9260 17013 9269
rect 17548 9260 17588 10672
rect 16971 9220 16972 9260
rect 17012 9220 17013 9260
rect 16971 9211 17013 9220
rect 17068 9220 17588 9260
rect 16779 8840 16821 8849
rect 16779 8800 16780 8840
rect 16820 8800 16821 8840
rect 16779 8791 16821 8800
rect 16972 8672 17012 9211
rect 16972 8429 17012 8632
rect 16971 8420 17013 8429
rect 16971 8380 16972 8420
rect 17012 8380 17013 8420
rect 16971 8371 17013 8380
rect 17068 8168 17108 9220
rect 17740 8849 17780 10672
rect 17355 8840 17397 8849
rect 17355 8800 17356 8840
rect 17396 8800 17397 8840
rect 17355 8791 17397 8800
rect 17739 8840 17781 8849
rect 17739 8800 17740 8840
rect 17780 8800 17781 8840
rect 17739 8791 17781 8800
rect 17068 8119 17108 8128
rect 16875 7916 16917 7925
rect 16875 7876 16876 7916
rect 16916 7876 16917 7916
rect 16875 7867 16917 7876
rect 16876 7782 16916 7867
rect 17260 7160 17300 7169
rect 17260 7001 17300 7120
rect 17259 6992 17301 7001
rect 17259 6952 17260 6992
rect 17300 6952 17301 6992
rect 17259 6943 17301 6952
rect 17260 5657 17300 6943
rect 17259 5648 17301 5657
rect 17259 5608 17260 5648
rect 17300 5608 17301 5648
rect 17259 5599 17301 5608
rect 16875 5228 16917 5237
rect 16875 5188 16876 5228
rect 16916 5188 16917 5228
rect 16875 5179 16917 5188
rect 16780 4808 16820 4817
rect 16588 4768 16780 4808
rect 16780 4759 16820 4768
rect 16876 4313 16916 5179
rect 16972 4892 17012 4901
rect 17164 4892 17204 4901
rect 17012 4852 17108 4892
rect 16972 4843 17012 4852
rect 16875 4304 16917 4313
rect 16875 4264 16876 4304
rect 16916 4264 16917 4304
rect 16875 4255 16917 4264
rect 16972 4141 17012 4150
rect 16532 4096 16916 4136
rect 15915 3296 15957 3305
rect 15915 3256 15916 3296
rect 15956 3256 15957 3296
rect 15915 3247 15957 3256
rect 16012 3137 16052 4096
rect 16492 4087 16532 4096
rect 16203 3800 16245 3809
rect 16203 3760 16204 3800
rect 16244 3760 16245 3800
rect 16203 3751 16245 3760
rect 15627 3128 15669 3137
rect 15627 3088 15628 3128
rect 15668 3088 15669 3128
rect 15627 3079 15669 3088
rect 16011 3128 16053 3137
rect 16011 3088 16012 3128
rect 16052 3088 16053 3128
rect 16011 3079 16053 3088
rect 15435 2960 15477 2969
rect 15435 2920 15436 2960
rect 15476 2920 15477 2960
rect 15435 2911 15477 2920
rect 14476 2500 14708 2540
rect 14379 2204 14421 2213
rect 14379 2164 14380 2204
rect 14420 2164 14421 2204
rect 14379 2155 14421 2164
rect 14476 1280 14516 2500
rect 15436 2129 15476 2911
rect 15628 2624 15668 3079
rect 16204 2885 16244 3751
rect 16779 3548 16821 3557
rect 16779 3508 16780 3548
rect 16820 3508 16821 3548
rect 16779 3499 16821 3508
rect 16780 3464 16820 3499
rect 16876 3464 16916 4096
rect 16972 3632 17012 4101
rect 17068 4052 17108 4852
rect 17204 4852 17300 4892
rect 17164 4843 17204 4852
rect 17164 4052 17204 4061
rect 17068 4012 17164 4052
rect 17164 4003 17204 4012
rect 17260 3977 17300 4852
rect 17356 4808 17396 8791
rect 17835 8756 17877 8765
rect 17835 8716 17836 8756
rect 17876 8716 17877 8756
rect 17835 8707 17877 8716
rect 17548 8000 17588 8009
rect 17452 7412 17492 7421
rect 17548 7412 17588 7960
rect 17643 8000 17685 8009
rect 17643 7960 17644 8000
rect 17684 7960 17685 8000
rect 17643 7951 17685 7960
rect 17644 7866 17684 7951
rect 17739 7664 17781 7673
rect 17739 7624 17740 7664
rect 17780 7624 17781 7664
rect 17739 7615 17781 7624
rect 17492 7372 17588 7412
rect 17452 7363 17492 7372
rect 17643 7160 17685 7169
rect 17643 7120 17644 7160
rect 17684 7120 17685 7160
rect 17643 7111 17685 7120
rect 17644 7026 17684 7111
rect 17740 6833 17780 7615
rect 17739 6824 17781 6833
rect 17739 6784 17740 6824
rect 17780 6784 17781 6824
rect 17739 6775 17781 6784
rect 17644 6488 17684 6497
rect 17644 5909 17684 6448
rect 17643 5900 17685 5909
rect 17643 5860 17644 5900
rect 17684 5860 17685 5900
rect 17643 5851 17685 5860
rect 17644 5741 17684 5851
rect 17643 5732 17685 5741
rect 17643 5692 17644 5732
rect 17684 5692 17685 5732
rect 17643 5683 17685 5692
rect 17547 5648 17589 5657
rect 17547 5608 17548 5648
rect 17588 5608 17589 5648
rect 17547 5599 17589 5608
rect 17548 5514 17588 5599
rect 17739 5564 17781 5573
rect 17739 5524 17740 5564
rect 17780 5524 17781 5564
rect 17739 5515 17781 5524
rect 17740 5430 17780 5515
rect 17356 4759 17396 4768
rect 17259 3968 17301 3977
rect 17259 3928 17260 3968
rect 17300 3928 17301 3968
rect 17259 3919 17301 3928
rect 16972 3583 17012 3592
rect 17740 3632 17780 3641
rect 17836 3632 17876 8707
rect 17780 3592 17876 3632
rect 17932 3632 17972 10672
rect 18124 8849 18164 10672
rect 18123 8840 18165 8849
rect 18123 8800 18124 8840
rect 18164 8800 18165 8840
rect 18123 8791 18165 8800
rect 18027 8672 18069 8681
rect 18027 8632 18028 8672
rect 18068 8632 18069 8672
rect 18027 8623 18069 8632
rect 18220 8672 18260 8681
rect 18028 7916 18068 8623
rect 18220 8345 18260 8632
rect 18219 8336 18261 8345
rect 18219 8296 18220 8336
rect 18260 8296 18261 8336
rect 18219 8287 18261 8296
rect 18123 8168 18165 8177
rect 18123 8128 18124 8168
rect 18164 8128 18165 8168
rect 18123 8119 18165 8128
rect 18124 8000 18164 8119
rect 18124 7951 18164 7960
rect 18028 7757 18068 7876
rect 18027 7748 18069 7757
rect 18027 7708 18028 7748
rect 18068 7708 18069 7748
rect 18316 7748 18356 10672
rect 18411 8840 18453 8849
rect 18411 8800 18412 8840
rect 18452 8800 18453 8840
rect 18411 8791 18453 8800
rect 18412 8706 18452 8791
rect 18508 8765 18548 10672
rect 18700 10529 18740 10672
rect 18699 10520 18741 10529
rect 18699 10480 18700 10520
rect 18740 10480 18741 10520
rect 18699 10471 18741 10480
rect 18892 10361 18932 10672
rect 18891 10352 18933 10361
rect 18891 10312 18892 10352
rect 18932 10312 18933 10352
rect 18891 10303 18933 10312
rect 18891 10016 18933 10025
rect 18891 9976 18892 10016
rect 18932 9976 18933 10016
rect 18891 9967 18933 9976
rect 18603 9512 18645 9521
rect 18603 9472 18604 9512
rect 18644 9472 18645 9512
rect 18603 9463 18645 9472
rect 18507 8756 18549 8765
rect 18507 8716 18508 8756
rect 18548 8716 18549 8756
rect 18507 8707 18549 8716
rect 18604 8672 18644 9463
rect 18795 9428 18837 9437
rect 18795 9388 18796 9428
rect 18836 9388 18837 9428
rect 18795 9379 18837 9388
rect 18796 9294 18836 9379
rect 18892 9353 18932 9967
rect 18988 9680 19028 9689
rect 19084 9680 19124 10672
rect 19179 9764 19221 9773
rect 19179 9724 19180 9764
rect 19220 9724 19221 9764
rect 19179 9715 19221 9724
rect 19028 9640 19124 9680
rect 18988 9631 19028 9640
rect 19180 9512 19220 9715
rect 19180 9353 19220 9472
rect 18891 9344 18933 9353
rect 18891 9304 18892 9344
rect 18932 9304 18933 9344
rect 18891 9295 18933 9304
rect 19179 9344 19221 9353
rect 19179 9304 19180 9344
rect 19220 9304 19221 9344
rect 19179 9295 19221 9304
rect 18808 9092 19176 9101
rect 18848 9052 18890 9092
rect 18930 9052 18972 9092
rect 19012 9052 19054 9092
rect 19094 9052 19136 9092
rect 18808 9043 19176 9052
rect 19276 8849 19316 10672
rect 19371 9428 19413 9437
rect 19371 9388 19372 9428
rect 19412 9388 19413 9428
rect 19371 9379 19413 9388
rect 18699 8840 18741 8849
rect 18699 8800 18700 8840
rect 18740 8800 18741 8840
rect 18699 8791 18741 8800
rect 19275 8840 19317 8849
rect 19275 8800 19276 8840
rect 19316 8800 19317 8840
rect 18603 8632 18644 8672
rect 18700 8672 18740 8791
rect 19180 8765 19220 8796
rect 19275 8791 19317 8800
rect 19179 8756 19221 8765
rect 19179 8716 19180 8756
rect 19220 8716 19221 8756
rect 19179 8707 19221 8716
rect 18603 8588 18643 8632
rect 18700 8623 18740 8632
rect 18796 8672 18836 8681
rect 18603 8548 18644 8588
rect 18604 8000 18644 8548
rect 18604 7841 18644 7960
rect 18603 7832 18645 7841
rect 18603 7792 18604 7832
rect 18644 7792 18645 7832
rect 18603 7783 18645 7792
rect 18796 7757 18836 8632
rect 19180 8672 19220 8707
rect 19180 8084 19220 8632
rect 19276 8672 19316 8683
rect 19276 8597 19316 8632
rect 19275 8588 19317 8597
rect 19275 8548 19276 8588
rect 19316 8548 19317 8588
rect 19275 8539 19317 8548
rect 19372 8420 19412 9379
rect 19276 8380 19412 8420
rect 19276 8210 19316 8380
rect 19276 8161 19316 8170
rect 19468 8168 19508 10672
rect 19563 8840 19605 8849
rect 19563 8800 19564 8840
rect 19604 8800 19605 8840
rect 19563 8791 19605 8800
rect 19468 8119 19508 8128
rect 19180 8044 19316 8084
rect 19276 8000 19316 8044
rect 19132 7958 19172 7967
rect 19276 7960 19412 8000
rect 19132 7916 19172 7918
rect 19132 7876 19316 7916
rect 18795 7748 18837 7757
rect 18316 7708 18452 7748
rect 18027 7699 18069 7708
rect 18315 7496 18357 7505
rect 18315 7456 18316 7496
rect 18356 7456 18357 7496
rect 18315 7447 18357 7456
rect 18316 6581 18356 7447
rect 18315 6572 18357 6581
rect 18315 6532 18316 6572
rect 18356 6532 18357 6572
rect 18315 6523 18357 6532
rect 18123 6152 18165 6161
rect 18123 6112 18124 6152
rect 18164 6112 18165 6152
rect 18123 6103 18165 6112
rect 18028 5648 18068 5659
rect 18124 5657 18164 6103
rect 18028 5573 18068 5608
rect 18123 5648 18165 5657
rect 18123 5608 18124 5648
rect 18164 5608 18165 5648
rect 18123 5599 18165 5608
rect 18027 5564 18069 5573
rect 18027 5524 18028 5564
rect 18068 5524 18069 5564
rect 18027 5515 18069 5524
rect 18124 5514 18164 5599
rect 18316 4976 18356 6523
rect 18316 4927 18356 4936
rect 18412 4817 18452 7708
rect 18795 7708 18796 7748
rect 18836 7708 18837 7748
rect 18795 7699 18837 7708
rect 18808 7580 19176 7589
rect 18848 7540 18890 7580
rect 18930 7540 18972 7580
rect 19012 7540 19054 7580
rect 19094 7540 19136 7580
rect 18808 7531 19176 7540
rect 19084 7412 19124 7421
rect 19276 7412 19316 7876
rect 19124 7372 19316 7412
rect 19084 7363 19124 7372
rect 18892 7160 18932 7169
rect 18892 7001 18932 7120
rect 18891 6992 18933 7001
rect 18891 6952 18892 6992
rect 18932 6952 18933 6992
rect 18891 6943 18933 6952
rect 19275 6992 19317 7001
rect 19275 6952 19276 6992
rect 19316 6952 19317 6992
rect 19275 6943 19317 6952
rect 18987 6908 19029 6917
rect 18987 6868 18988 6908
rect 19028 6868 19029 6908
rect 18987 6859 19029 6868
rect 18988 6665 19028 6859
rect 18987 6656 19029 6665
rect 18987 6616 18988 6656
rect 19028 6616 19029 6656
rect 18987 6607 19029 6616
rect 18891 6488 18933 6497
rect 18891 6448 18892 6488
rect 18932 6448 18933 6488
rect 18891 6439 18933 6448
rect 18892 6354 18932 6439
rect 19084 6329 19124 6414
rect 19083 6320 19125 6329
rect 19083 6280 19084 6320
rect 19124 6280 19125 6320
rect 19083 6271 19125 6280
rect 18808 6068 19176 6077
rect 18848 6028 18890 6068
rect 18930 6028 18972 6068
rect 19012 6028 19054 6068
rect 19094 6028 19136 6068
rect 18808 6019 19176 6028
rect 18604 5741 18644 5772
rect 18603 5732 18645 5741
rect 18603 5692 18604 5732
rect 18644 5692 18645 5732
rect 18603 5683 18645 5692
rect 18508 5648 18548 5657
rect 18508 5489 18548 5608
rect 18604 5648 18644 5683
rect 18507 5480 18549 5489
rect 18507 5440 18508 5480
rect 18548 5440 18549 5480
rect 18507 5431 18549 5440
rect 18604 5321 18644 5608
rect 19084 5648 19124 5657
rect 18603 5312 18645 5321
rect 18603 5272 18604 5312
rect 18644 5272 18645 5312
rect 18603 5263 18645 5272
rect 19084 5237 19124 5608
rect 19083 5228 19125 5237
rect 19083 5188 19084 5228
rect 19124 5188 19125 5228
rect 19083 5179 19125 5188
rect 19276 4985 19316 6943
rect 19372 6488 19412 7960
rect 19468 6656 19508 6665
rect 19564 6656 19604 8791
rect 19660 8504 19700 10672
rect 19755 10016 19797 10025
rect 19755 9976 19756 10016
rect 19796 9976 19797 10016
rect 19755 9967 19797 9976
rect 19756 8672 19796 9967
rect 19756 8623 19796 8632
rect 19660 8464 19796 8504
rect 19659 7160 19701 7169
rect 19659 7120 19660 7160
rect 19700 7120 19701 7160
rect 19659 7111 19701 7120
rect 19660 7026 19700 7111
rect 19756 6665 19796 8464
rect 19852 6917 19892 10672
rect 20044 10445 20084 10672
rect 20043 10436 20085 10445
rect 20043 10396 20044 10436
rect 20084 10396 20085 10436
rect 20043 10387 20085 10396
rect 20236 10016 20276 10672
rect 20428 10277 20468 10672
rect 20619 10648 20620 10672
rect 20660 10672 20680 10688
rect 20792 10672 20872 10752
rect 20984 10672 21064 10752
rect 21176 10672 21256 10752
rect 21368 10672 21448 10752
rect 21560 10672 21640 10752
rect 21752 10672 21832 10752
rect 21944 10672 22024 10752
rect 22136 10672 22216 10752
rect 22328 10672 22408 10752
rect 22520 10672 22600 10752
rect 22712 10672 22792 10752
rect 22904 10672 22984 10752
rect 23096 10672 23176 10752
rect 23288 10672 23368 10752
rect 23480 10672 23560 10752
rect 23672 10672 23752 10752
rect 23864 10672 23944 10752
rect 24056 10672 24136 10752
rect 24248 10672 24328 10752
rect 24440 10672 24520 10752
rect 24632 10672 24712 10752
rect 24824 10672 24904 10752
rect 25016 10672 25096 10752
rect 25208 10672 25288 10752
rect 25400 10672 25480 10752
rect 25592 10672 25672 10752
rect 25784 10672 25864 10752
rect 25976 10672 26056 10752
rect 26168 10672 26248 10752
rect 26360 10672 26440 10752
rect 26552 10672 26632 10752
rect 26744 10672 26824 10752
rect 26936 10672 27016 10752
rect 27128 10672 27208 10752
rect 27320 10672 27400 10752
rect 27512 10672 27592 10752
rect 27704 10672 27784 10752
rect 27896 10672 27976 10752
rect 28088 10672 28168 10752
rect 28280 10672 28360 10752
rect 28472 10672 28552 10752
rect 28664 10672 28744 10752
rect 28856 10672 28936 10752
rect 29048 10672 29128 10752
rect 29240 10672 29320 10752
rect 29432 10672 29512 10752
rect 29624 10672 29704 10752
rect 29816 10672 29896 10752
rect 30008 10672 30088 10752
rect 30200 10672 30280 10752
rect 30392 10672 30472 10752
rect 30584 10672 30664 10752
rect 30776 10672 30856 10752
rect 30968 10672 31048 10752
rect 31160 10672 31240 10752
rect 31352 10672 31432 10752
rect 31544 10672 31624 10752
rect 31736 10672 31816 10752
rect 31928 10672 32008 10752
rect 32120 10672 32200 10752
rect 32312 10672 32392 10752
rect 32504 10672 32584 10752
rect 32696 10688 32776 10752
rect 32631 10672 32776 10688
rect 32888 10672 32968 10752
rect 33080 10672 33160 10752
rect 33272 10672 33352 10752
rect 33464 10672 33544 10752
rect 20660 10648 20661 10672
rect 20619 10639 20661 10648
rect 20427 10268 20469 10277
rect 20427 10228 20428 10268
rect 20468 10228 20469 10268
rect 20427 10219 20469 10228
rect 20236 9976 20756 10016
rect 19947 9932 19989 9941
rect 19947 9892 19948 9932
rect 19988 9892 19989 9932
rect 19947 9883 19989 9892
rect 19948 8168 19988 9883
rect 20048 9848 20416 9857
rect 20088 9808 20130 9848
rect 20170 9808 20212 9848
rect 20252 9808 20294 9848
rect 20334 9808 20376 9848
rect 20048 9799 20416 9808
rect 20428 9512 20468 9521
rect 20236 9472 20428 9512
rect 20236 8840 20276 9472
rect 20428 9463 20468 9472
rect 20620 9260 20660 9269
rect 20140 8800 20276 8840
rect 20332 9220 20620 9260
rect 20140 8681 20180 8800
rect 20332 8756 20372 9220
rect 20620 9211 20660 9220
rect 20716 9092 20756 9976
rect 20284 8716 20372 8756
rect 20620 9052 20756 9092
rect 20284 8714 20324 8716
rect 20139 8672 20181 8681
rect 20139 8632 20140 8672
rect 20180 8632 20181 8672
rect 20284 8665 20324 8674
rect 20139 8623 20181 8632
rect 20428 8504 20468 8513
rect 20468 8464 20564 8504
rect 20428 8455 20468 8464
rect 20048 8336 20416 8345
rect 20088 8296 20130 8336
rect 20170 8296 20212 8336
rect 20252 8296 20294 8336
rect 20334 8296 20376 8336
rect 20048 8287 20416 8296
rect 20044 8168 20084 8177
rect 20524 8168 20564 8464
rect 19948 8128 20044 8168
rect 20044 8119 20084 8128
rect 20236 8128 20564 8168
rect 20236 7916 20276 8128
rect 20236 7867 20276 7876
rect 19851 6908 19893 6917
rect 19851 6868 19852 6908
rect 19892 6868 19893 6908
rect 19851 6859 19893 6868
rect 20048 6824 20416 6833
rect 20088 6784 20130 6824
rect 20170 6784 20212 6824
rect 20252 6784 20294 6824
rect 20334 6784 20376 6824
rect 20048 6775 20416 6784
rect 20620 6749 20660 9052
rect 20716 8672 20756 8681
rect 20716 7757 20756 8632
rect 20812 8177 20852 10672
rect 20907 10268 20949 10277
rect 20907 10228 20908 10268
rect 20948 10228 20949 10268
rect 21004 10268 21044 10672
rect 21099 10268 21141 10277
rect 21004 10228 21100 10268
rect 21140 10228 21141 10268
rect 20907 10219 20949 10228
rect 21099 10219 21141 10228
rect 20811 8168 20853 8177
rect 20811 8128 20812 8168
rect 20852 8128 20853 8168
rect 20811 8119 20853 8128
rect 20811 8000 20853 8009
rect 20811 7960 20812 8000
rect 20852 7960 20853 8000
rect 20811 7951 20853 7960
rect 20715 7748 20757 7757
rect 20715 7708 20716 7748
rect 20756 7708 20757 7748
rect 20812 7748 20852 7951
rect 20908 7925 20948 10219
rect 21003 8672 21045 8681
rect 21003 8632 21004 8672
rect 21044 8632 21045 8672
rect 21003 8623 21045 8632
rect 21004 8177 21044 8623
rect 21196 8513 21236 10672
rect 21195 8504 21237 8513
rect 21195 8464 21196 8504
rect 21236 8464 21237 8504
rect 21195 8455 21237 8464
rect 21003 8168 21045 8177
rect 21388 8168 21428 10672
rect 21580 9521 21620 10672
rect 21579 9512 21621 9521
rect 21579 9472 21580 9512
rect 21620 9472 21621 9512
rect 21579 9463 21621 9472
rect 21483 8924 21525 8933
rect 21483 8884 21484 8924
rect 21524 8884 21525 8924
rect 21483 8875 21525 8884
rect 21003 8128 21004 8168
rect 21044 8128 21045 8168
rect 21003 8119 21045 8128
rect 21292 8128 21428 8168
rect 21004 8000 21044 8009
rect 20907 7916 20949 7925
rect 20907 7876 20908 7916
rect 20948 7876 20949 7916
rect 20907 7867 20949 7876
rect 20812 7708 20948 7748
rect 20715 7699 20757 7708
rect 20811 7580 20853 7589
rect 20811 7540 20812 7580
rect 20852 7540 20853 7580
rect 20811 7531 20853 7540
rect 20619 6740 20661 6749
rect 20619 6700 20620 6740
rect 20660 6700 20661 6740
rect 20619 6691 20661 6700
rect 19508 6616 19604 6656
rect 19755 6656 19797 6665
rect 19755 6616 19756 6656
rect 19796 6616 19797 6656
rect 19468 6607 19508 6616
rect 19755 6607 19797 6616
rect 20331 6656 20373 6665
rect 20331 6616 20332 6656
rect 20372 6616 20373 6656
rect 20331 6607 20373 6616
rect 19851 6572 19893 6581
rect 19851 6532 19852 6572
rect 19892 6532 19893 6572
rect 19851 6523 19893 6532
rect 19852 6488 19892 6523
rect 19372 6448 19508 6488
rect 19371 6236 19413 6245
rect 19371 6196 19372 6236
rect 19412 6196 19413 6236
rect 19371 6187 19413 6196
rect 19372 5993 19412 6187
rect 19371 5984 19413 5993
rect 19371 5944 19372 5984
rect 19412 5944 19413 5984
rect 19371 5935 19413 5944
rect 19468 5816 19508 6448
rect 19372 5776 19508 5816
rect 19660 6404 19700 6413
rect 19275 4976 19317 4985
rect 19275 4936 19276 4976
rect 19316 4936 19317 4976
rect 19275 4927 19317 4936
rect 18411 4808 18453 4817
rect 18411 4768 18412 4808
rect 18452 4768 18453 4808
rect 18411 4759 18453 4768
rect 18808 4556 19176 4565
rect 18848 4516 18890 4556
rect 18930 4516 18972 4556
rect 19012 4516 19054 4556
rect 19094 4516 19136 4556
rect 18808 4507 19176 4516
rect 19372 4229 19412 5776
rect 19564 5653 19604 5662
rect 19467 5396 19509 5405
rect 19467 5356 19468 5396
rect 19508 5356 19509 5396
rect 19467 5347 19509 5356
rect 19371 4220 19413 4229
rect 19371 4180 19372 4220
rect 19412 4180 19413 4220
rect 19371 4171 19413 4180
rect 19275 3800 19317 3809
rect 19275 3760 19276 3800
rect 19316 3760 19317 3800
rect 19275 3751 19317 3760
rect 17740 3583 17780 3592
rect 17932 3583 17972 3592
rect 18315 3464 18357 3473
rect 16876 3424 17204 3464
rect 16780 3413 16820 3424
rect 16587 3296 16629 3305
rect 16587 3256 16588 3296
rect 16628 3256 16629 3296
rect 16587 3247 16629 3256
rect 16203 2876 16245 2885
rect 16203 2836 16204 2876
rect 16244 2836 16245 2876
rect 16203 2827 16245 2836
rect 15435 2120 15477 2129
rect 15435 2080 15436 2120
rect 15476 2080 15477 2120
rect 15052 2045 15092 2076
rect 15435 2071 15477 2080
rect 15051 2036 15093 2045
rect 15051 1996 15052 2036
rect 15092 1996 15093 2036
rect 15051 1987 15093 1996
rect 15052 1952 15092 1987
rect 15052 1877 15092 1912
rect 15436 1952 15476 2071
rect 15436 1903 15476 1912
rect 15051 1868 15093 1877
rect 15051 1828 15052 1868
rect 15092 1828 15093 1868
rect 15051 1819 15093 1828
rect 14476 1231 14516 1240
rect 15244 1700 15284 1709
rect 14284 1063 14324 1072
rect 14667 1112 14709 1121
rect 14667 1072 14668 1112
rect 14708 1072 14709 1112
rect 14667 1063 14709 1072
rect 14668 953 14708 1063
rect 13611 944 13653 953
rect 13611 904 13612 944
rect 13652 904 13653 944
rect 13611 895 13653 904
rect 14475 944 14517 953
rect 14475 904 14476 944
rect 14516 904 14517 944
rect 14475 895 14517 904
rect 14667 944 14709 953
rect 14667 904 14668 944
rect 14708 904 14709 944
rect 14667 895 14709 904
rect 13035 692 13077 701
rect 13035 652 13036 692
rect 13076 652 13077 692
rect 13035 643 13077 652
rect 12843 104 12885 113
rect 11060 64 11080 80
rect 11000 0 11080 64
rect 12152 0 12232 80
rect 12843 64 12844 104
rect 12884 64 12885 104
rect 13323 104 13365 113
rect 13323 80 13324 104
rect 12843 55 12885 64
rect 13304 64 13324 80
rect 13364 80 13365 104
rect 14476 80 14516 895
rect 13364 64 13384 80
rect 13304 0 13384 64
rect 14456 0 14536 80
rect 15244 60 15284 1660
rect 15628 1121 15668 2584
rect 16108 2624 16148 2633
rect 15820 2540 15860 2549
rect 16108 2540 16148 2584
rect 16204 2624 16244 2827
rect 16588 2708 16628 3247
rect 16683 3128 16725 3137
rect 16683 3088 16684 3128
rect 16724 3088 16725 3128
rect 16683 3079 16725 3088
rect 16588 2659 16628 2668
rect 16684 2708 16724 3079
rect 16684 2659 16724 2668
rect 16204 2575 16244 2584
rect 17164 2624 17204 3424
rect 18315 3424 18316 3464
rect 18356 3424 18357 3464
rect 18315 3415 18357 3424
rect 17548 3380 17588 3389
rect 18123 3380 18165 3389
rect 17588 3340 17876 3380
rect 17548 3331 17588 3340
rect 17692 2633 17732 2642
rect 17732 2593 17780 2624
rect 17692 2584 17780 2593
rect 15860 2500 16148 2540
rect 15820 2491 15860 2500
rect 16684 2045 16724 2076
rect 16683 2036 16725 2045
rect 16683 1996 16684 2036
rect 16724 1996 16725 2036
rect 16683 1987 16725 1996
rect 17164 2036 17204 2584
rect 17164 1987 17204 1996
rect 16299 1952 16341 1961
rect 16299 1912 16300 1952
rect 16340 1912 16341 1952
rect 16299 1903 16341 1912
rect 16684 1952 16724 1987
rect 15627 1112 15669 1121
rect 15627 1072 15628 1112
rect 15668 1072 15669 1112
rect 15627 1063 15669 1072
rect 16300 1112 16340 1903
rect 16684 1793 16724 1912
rect 17548 1952 17588 1961
rect 16683 1784 16725 1793
rect 16683 1744 16684 1784
rect 16724 1744 16725 1784
rect 16683 1735 16725 1744
rect 16876 1700 16916 1709
rect 16300 1063 16340 1072
rect 16780 1660 16876 1700
rect 15339 104 15381 113
rect 15339 64 15340 104
rect 15380 64 15381 104
rect 15627 104 15669 113
rect 15627 80 15628 104
rect 15339 60 15381 64
rect 15244 55 15381 60
rect 15608 64 15628 80
rect 15668 80 15669 104
rect 16780 80 16820 1660
rect 16876 1651 16916 1660
rect 17548 1289 17588 1912
rect 17547 1280 17589 1289
rect 17547 1240 17548 1280
rect 17588 1240 17589 1280
rect 17547 1231 17589 1240
rect 17740 1280 17780 2584
rect 17836 2540 17876 3340
rect 18123 3340 18124 3380
rect 18164 3340 18165 3380
rect 18123 3331 18165 3340
rect 18124 3246 18164 3331
rect 18316 3221 18356 3415
rect 18315 3212 18357 3221
rect 18315 3172 18316 3212
rect 18356 3172 18357 3212
rect 18315 3163 18357 3172
rect 18808 3044 19176 3053
rect 18848 3004 18890 3044
rect 18930 3004 18972 3044
rect 19012 3004 19054 3044
rect 19094 3004 19136 3044
rect 18808 2995 19176 3004
rect 18028 2633 18068 2718
rect 18027 2624 18069 2633
rect 18027 2584 18028 2624
rect 18068 2584 18069 2624
rect 18027 2575 18069 2584
rect 18411 2624 18453 2633
rect 18411 2584 18412 2624
rect 18452 2584 18453 2624
rect 18411 2575 18453 2584
rect 19276 2624 19316 3751
rect 19468 3296 19508 5347
rect 19564 5144 19604 5613
rect 19660 5564 19700 6364
rect 19852 5573 19892 6448
rect 19947 5816 19989 5825
rect 19947 5776 19948 5816
rect 19988 5776 19989 5816
rect 19947 5767 19989 5776
rect 19948 5682 19988 5767
rect 20332 5657 20372 6607
rect 20619 6320 20661 6329
rect 20619 6280 20620 6320
rect 20660 6280 20661 6320
rect 20619 6271 20661 6280
rect 20331 5648 20373 5657
rect 20331 5608 20332 5648
rect 20372 5608 20373 5648
rect 20331 5599 20373 5608
rect 20620 5648 20660 6271
rect 20620 5599 20660 5608
rect 19756 5564 19796 5573
rect 19660 5524 19756 5564
rect 19756 5515 19796 5524
rect 19851 5564 19893 5573
rect 20236 5564 20276 5573
rect 19851 5524 19852 5564
rect 19892 5524 19893 5564
rect 19851 5515 19893 5524
rect 19948 5524 20236 5564
rect 19948 5405 19988 5524
rect 20236 5515 20276 5524
rect 20332 5514 20372 5599
rect 19947 5396 19989 5405
rect 19947 5356 19948 5396
rect 19988 5356 19989 5396
rect 19947 5347 19989 5356
rect 20048 5312 20416 5321
rect 20088 5272 20130 5312
rect 20170 5272 20212 5312
rect 20252 5272 20294 5312
rect 20334 5272 20376 5312
rect 20048 5263 20416 5272
rect 19756 5144 19796 5153
rect 19564 5104 19756 5144
rect 19756 5095 19796 5104
rect 19563 4976 19605 4985
rect 19563 4936 19564 4976
rect 19604 4936 19605 4976
rect 19563 4927 19605 4936
rect 19564 4565 19604 4927
rect 19563 4556 19605 4565
rect 19563 4516 19564 4556
rect 19604 4516 19605 4556
rect 19563 4507 19605 4516
rect 19564 3809 19604 4507
rect 20331 4220 20373 4229
rect 20331 4180 20332 4220
rect 20372 4180 20373 4220
rect 20331 4171 20373 4180
rect 19852 4136 19892 4145
rect 19563 3800 19605 3809
rect 19563 3760 19564 3800
rect 19604 3760 19605 3800
rect 19563 3751 19605 3760
rect 19564 3464 19604 3751
rect 19756 3632 19796 3641
rect 19852 3632 19892 4096
rect 19947 4136 19989 4145
rect 19947 4096 19948 4136
rect 19988 4096 19989 4136
rect 19947 4087 19989 4096
rect 19948 4002 19988 4087
rect 20332 4086 20372 4171
rect 20428 4136 20468 4145
rect 20812 4136 20852 7531
rect 20908 7169 20948 7708
rect 21004 7412 21044 7960
rect 21100 8000 21140 8009
rect 21140 7960 21236 8000
rect 21100 7951 21140 7960
rect 21100 7412 21140 7421
rect 21004 7372 21100 7412
rect 21100 7363 21140 7372
rect 20907 7160 20949 7169
rect 20907 7120 20908 7160
rect 20948 7120 20949 7160
rect 20907 7111 20949 7120
rect 20908 7026 20948 7111
rect 21196 6581 21236 7960
rect 21292 6992 21332 8128
rect 21484 8084 21524 8875
rect 21675 8840 21717 8849
rect 21675 8800 21676 8840
rect 21716 8800 21717 8840
rect 21675 8791 21717 8800
rect 21579 8672 21621 8681
rect 21579 8632 21580 8672
rect 21620 8632 21621 8672
rect 21579 8623 21621 8632
rect 21388 8044 21524 8084
rect 21388 7748 21428 8044
rect 21580 8000 21620 8623
rect 21580 7951 21620 7960
rect 21484 7916 21524 7925
rect 21484 7832 21524 7876
rect 21579 7832 21621 7841
rect 21484 7792 21580 7832
rect 21620 7792 21621 7832
rect 21579 7783 21621 7792
rect 21388 7708 21524 7748
rect 21388 7160 21428 7169
rect 21484 7160 21524 7708
rect 21676 7673 21716 8791
rect 21772 8093 21812 10672
rect 21867 9344 21909 9353
rect 21867 9304 21868 9344
rect 21908 9304 21909 9344
rect 21867 9295 21909 9304
rect 21771 8084 21813 8093
rect 21771 8044 21772 8084
rect 21812 8044 21813 8084
rect 21771 8035 21813 8044
rect 21771 7916 21813 7925
rect 21771 7876 21772 7916
rect 21812 7876 21813 7916
rect 21771 7867 21813 7876
rect 21675 7664 21717 7673
rect 21675 7624 21676 7664
rect 21716 7624 21717 7664
rect 21675 7615 21717 7624
rect 21428 7120 21524 7160
rect 21388 7111 21428 7120
rect 21292 6952 21428 6992
rect 21291 6656 21333 6665
rect 21291 6616 21292 6656
rect 21332 6616 21333 6656
rect 21291 6607 21333 6616
rect 21195 6572 21237 6581
rect 21195 6532 21196 6572
rect 21236 6532 21237 6572
rect 21195 6523 21237 6532
rect 21292 6522 21332 6607
rect 21100 6488 21140 6497
rect 20907 6152 20949 6161
rect 20907 6112 20908 6152
rect 20948 6112 20949 6152
rect 20907 6103 20949 6112
rect 20908 5489 20948 6103
rect 21100 6077 21140 6448
rect 21388 6161 21428 6952
rect 21484 6917 21524 7120
rect 21483 6908 21525 6917
rect 21483 6868 21484 6908
rect 21524 6868 21525 6908
rect 21483 6859 21525 6868
rect 21483 6656 21525 6665
rect 21483 6616 21484 6656
rect 21524 6616 21525 6656
rect 21483 6607 21525 6616
rect 21484 6488 21524 6607
rect 21580 6488 21620 6497
rect 21484 6448 21580 6488
rect 21580 6439 21620 6448
rect 21676 6488 21716 7615
rect 21676 6439 21716 6448
rect 21772 6320 21812 7867
rect 21868 7841 21908 9295
rect 21964 8933 22004 10672
rect 22156 9092 22196 10672
rect 22251 9680 22293 9689
rect 22251 9640 22252 9680
rect 22292 9640 22293 9680
rect 22251 9631 22293 9640
rect 22252 9546 22292 9631
rect 22156 9052 22292 9092
rect 21963 8924 22005 8933
rect 21963 8884 21964 8924
rect 22004 8884 22005 8924
rect 21963 8875 22005 8884
rect 22155 8924 22197 8933
rect 22155 8884 22156 8924
rect 22196 8884 22197 8924
rect 22155 8875 22197 8884
rect 22156 8756 22196 8875
rect 22252 8849 22292 9052
rect 22251 8840 22293 8849
rect 22251 8800 22252 8840
rect 22292 8800 22293 8840
rect 22251 8791 22293 8800
rect 22348 8765 22388 10672
rect 22540 9605 22580 10672
rect 22732 10352 22772 10672
rect 22924 10436 22964 10672
rect 22924 10396 23060 10436
rect 22732 10312 22964 10352
rect 22827 10184 22869 10193
rect 22827 10144 22828 10184
rect 22868 10144 22869 10184
rect 22827 10135 22869 10144
rect 22539 9596 22581 9605
rect 22539 9556 22540 9596
rect 22580 9556 22581 9596
rect 22539 9547 22581 9556
rect 22731 9512 22773 9521
rect 22731 9472 22732 9512
rect 22772 9472 22773 9512
rect 22731 9463 22773 9472
rect 22444 9428 22484 9437
rect 22484 9388 22580 9428
rect 22444 9379 22484 9388
rect 22540 8840 22580 9388
rect 22732 9378 22772 9463
rect 22540 8800 22772 8840
rect 21964 8716 22196 8756
rect 22347 8756 22389 8765
rect 22347 8716 22348 8756
rect 22388 8716 22389 8756
rect 21964 8672 22004 8716
rect 22347 8707 22389 8716
rect 21867 7832 21909 7841
rect 21867 7792 21868 7832
rect 21908 7792 21909 7832
rect 21867 7783 21909 7792
rect 21484 6280 21812 6320
rect 21387 6152 21429 6161
rect 21387 6112 21388 6152
rect 21428 6112 21429 6152
rect 21387 6103 21429 6112
rect 21099 6068 21141 6077
rect 21099 6028 21100 6068
rect 21140 6028 21236 6068
rect 21099 6019 21141 6028
rect 20907 5480 20949 5489
rect 20907 5440 20908 5480
rect 20948 5440 20949 5480
rect 20907 5431 20949 5440
rect 21099 4892 21141 4901
rect 21099 4852 21100 4892
rect 21140 4852 21141 4892
rect 21099 4843 21141 4852
rect 20907 4808 20949 4817
rect 20907 4768 20908 4808
rect 20948 4768 20949 4808
rect 20907 4759 20949 4768
rect 20908 4674 20948 4759
rect 21100 4758 21140 4843
rect 20908 4136 20948 4145
rect 20468 4096 20564 4136
rect 20428 4087 20468 4096
rect 20048 3800 20416 3809
rect 20088 3760 20130 3800
rect 20170 3760 20212 3800
rect 20252 3760 20294 3800
rect 20334 3760 20376 3800
rect 20048 3751 20416 3760
rect 19796 3592 19892 3632
rect 19756 3583 19796 3592
rect 19564 3415 19604 3424
rect 20044 3464 20084 3475
rect 20044 3389 20084 3424
rect 19659 3380 19701 3389
rect 19659 3340 19660 3380
rect 19700 3340 19701 3380
rect 19659 3331 19701 3340
rect 20043 3380 20085 3389
rect 20043 3340 20044 3380
rect 20084 3340 20085 3380
rect 20043 3331 20085 3340
rect 19468 3256 19604 3296
rect 19467 2792 19509 2801
rect 19467 2752 19468 2792
rect 19508 2752 19509 2792
rect 19467 2743 19509 2752
rect 19468 2658 19508 2743
rect 17836 2491 17876 2500
rect 18412 1952 18452 2575
rect 18412 1903 18452 1912
rect 18808 1532 19176 1541
rect 18848 1492 18890 1532
rect 18930 1492 18972 1532
rect 19012 1492 19054 1532
rect 19094 1492 19136 1532
rect 18808 1483 19176 1492
rect 17932 1289 17972 1374
rect 19276 1289 19316 2584
rect 19564 2120 19604 3256
rect 19660 2540 19700 3331
rect 20331 3212 20373 3221
rect 20331 3172 20332 3212
rect 20372 3172 20373 3212
rect 20331 3163 20373 3172
rect 20043 2792 20085 2801
rect 20043 2752 20044 2792
rect 20084 2752 20085 2792
rect 20043 2743 20085 2752
rect 19660 2491 19700 2500
rect 19852 2629 19892 2638
rect 19564 2071 19604 2080
rect 17740 1231 17780 1240
rect 17931 1280 17973 1289
rect 17931 1240 17932 1280
rect 17972 1240 17973 1280
rect 17931 1231 17973 1240
rect 19083 1280 19125 1289
rect 19083 1240 19084 1280
rect 19124 1240 19125 1280
rect 19083 1231 19125 1240
rect 19275 1280 19317 1289
rect 19275 1240 19276 1280
rect 19316 1240 19317 1280
rect 19275 1231 19317 1240
rect 19659 1280 19701 1289
rect 19659 1240 19660 1280
rect 19700 1240 19701 1280
rect 19659 1231 19701 1240
rect 19852 1280 19892 2589
rect 20044 2549 20084 2743
rect 20332 2624 20372 3163
rect 20524 2885 20564 4096
rect 20812 4096 20908 4136
rect 20812 3641 20852 4096
rect 20908 4087 20948 4096
rect 20811 3632 20853 3641
rect 20811 3592 20812 3632
rect 20852 3592 20853 3632
rect 20811 3583 20853 3592
rect 21196 3464 21236 6028
rect 21291 5900 21333 5909
rect 21291 5860 21292 5900
rect 21332 5860 21333 5900
rect 21291 5851 21333 5860
rect 21292 5648 21332 5851
rect 21292 5237 21332 5608
rect 21291 5228 21333 5237
rect 21291 5188 21292 5228
rect 21332 5188 21333 5228
rect 21291 5179 21333 5188
rect 21388 4976 21428 4985
rect 21388 4304 21428 4936
rect 21484 4976 21524 6280
rect 21675 5900 21717 5909
rect 21675 5860 21676 5900
rect 21716 5860 21717 5900
rect 21675 5851 21717 5860
rect 21484 4927 21524 4936
rect 21579 4892 21621 4901
rect 21579 4852 21580 4892
rect 21620 4852 21621 4892
rect 21579 4843 21621 4852
rect 21388 4264 21524 4304
rect 21388 4141 21428 4150
rect 21292 3464 21332 3473
rect 21196 3424 21292 3464
rect 21388 3464 21428 4101
rect 21484 3632 21524 4264
rect 21580 4052 21620 4843
rect 21580 4003 21620 4012
rect 21484 3583 21524 3592
rect 21388 3424 21524 3464
rect 20907 3296 20949 3305
rect 20907 3256 20908 3296
rect 20948 3256 20949 3296
rect 20907 3247 20949 3256
rect 20715 3128 20757 3137
rect 20715 3088 20716 3128
rect 20756 3088 20757 3128
rect 20715 3079 20757 3088
rect 20523 2876 20565 2885
rect 20523 2836 20524 2876
rect 20564 2836 20565 2876
rect 20523 2827 20565 2836
rect 20332 2575 20372 2584
rect 20043 2540 20085 2549
rect 20043 2500 20044 2540
rect 20084 2500 20085 2540
rect 20043 2491 20085 2500
rect 20048 2288 20416 2297
rect 20088 2248 20130 2288
rect 20170 2248 20212 2288
rect 20252 2248 20294 2288
rect 20334 2248 20376 2288
rect 20048 2239 20416 2248
rect 20043 2120 20085 2129
rect 20043 2080 20044 2120
rect 20084 2080 20085 2120
rect 20043 2071 20085 2080
rect 20139 2120 20181 2129
rect 20139 2080 20140 2120
rect 20180 2080 20181 2120
rect 20139 2071 20181 2080
rect 20044 1709 20084 2071
rect 20140 1877 20180 2071
rect 20139 1868 20181 1877
rect 20139 1828 20140 1868
rect 20180 1828 20181 1868
rect 20139 1819 20181 1828
rect 20043 1700 20085 1709
rect 20043 1660 20044 1700
rect 20084 1660 20085 1700
rect 20043 1651 20085 1660
rect 19852 1231 19892 1240
rect 17547 1112 17589 1121
rect 17547 1072 17548 1112
rect 17588 1072 17589 1112
rect 17547 1063 17589 1072
rect 17931 1112 17973 1121
rect 17931 1072 17932 1112
rect 17972 1072 17973 1112
rect 17931 1063 17973 1072
rect 18412 1112 18452 1121
rect 17548 785 17588 1063
rect 17547 776 17589 785
rect 17547 736 17548 776
rect 17588 736 17589 776
rect 17547 727 17589 736
rect 17932 80 17972 1063
rect 18412 869 18452 1072
rect 18411 860 18453 869
rect 18411 820 18412 860
rect 18452 820 18453 860
rect 18411 811 18453 820
rect 18412 617 18452 811
rect 19084 785 19124 1231
rect 19660 1112 19700 1231
rect 19660 1063 19700 1072
rect 20044 1112 20084 1651
rect 20044 1063 20084 1072
rect 19083 776 19125 785
rect 19083 736 19084 776
rect 19124 736 19125 776
rect 19083 727 19125 736
rect 20048 776 20416 785
rect 20088 736 20130 776
rect 20170 736 20212 776
rect 20252 736 20294 776
rect 20334 736 20376 776
rect 20048 727 20416 736
rect 18411 608 18453 617
rect 18411 568 18412 608
rect 18452 568 18453 608
rect 18411 559 18453 568
rect 19084 80 19124 727
rect 20235 104 20277 113
rect 20235 80 20236 104
rect 15668 64 15688 80
rect 15244 20 15380 55
rect 15608 0 15688 64
rect 16760 0 16840 80
rect 17912 0 17992 80
rect 19064 0 19144 80
rect 20216 64 20236 80
rect 20276 80 20277 104
rect 20427 104 20469 113
rect 20276 64 20296 80
rect 20216 0 20296 64
rect 20427 64 20428 104
rect 20468 64 20469 104
rect 20427 60 20469 64
rect 20716 60 20756 3079
rect 20811 3044 20853 3053
rect 20811 3004 20812 3044
rect 20852 3004 20853 3044
rect 20811 2995 20853 3004
rect 20812 2801 20852 2995
rect 20811 2792 20853 2801
rect 20811 2752 20812 2792
rect 20852 2752 20853 2792
rect 20811 2743 20853 2752
rect 20812 2708 20852 2743
rect 20812 2658 20852 2668
rect 20908 2708 20948 3247
rect 20908 2659 20948 2668
rect 21196 2297 21236 3424
rect 21292 3415 21332 3424
rect 21291 2876 21333 2885
rect 21291 2836 21292 2876
rect 21332 2836 21333 2876
rect 21291 2827 21333 2836
rect 21292 2624 21332 2827
rect 21387 2792 21429 2801
rect 21387 2752 21388 2792
rect 21428 2752 21429 2792
rect 21387 2743 21429 2752
rect 21292 2575 21332 2584
rect 21388 2624 21428 2743
rect 21388 2575 21428 2584
rect 21195 2288 21237 2297
rect 21195 2248 21196 2288
rect 21236 2248 21237 2288
rect 21195 2239 21237 2248
rect 21387 2288 21429 2297
rect 21387 2248 21388 2288
rect 21428 2248 21429 2288
rect 21387 2239 21429 2248
rect 21291 2036 21333 2045
rect 21291 1996 21292 2036
rect 21332 1996 21333 2036
rect 21291 1987 21333 1996
rect 21292 1952 21332 1987
rect 21292 1901 21332 1912
rect 21291 1280 21333 1289
rect 21291 1240 21292 1280
rect 21332 1240 21333 1280
rect 21291 1231 21333 1240
rect 21292 1112 21332 1231
rect 21292 1063 21332 1072
rect 21388 80 21428 2239
rect 21484 1280 21524 3424
rect 21676 2540 21716 5851
rect 21868 5060 21908 7783
rect 21964 6665 22004 8632
rect 22444 8672 22484 8681
rect 22156 8588 22196 8597
rect 22444 8588 22484 8632
rect 22196 8548 22484 8588
rect 22540 8672 22580 8681
rect 22156 8539 22196 8548
rect 22540 8513 22580 8632
rect 22539 8504 22581 8513
rect 22539 8464 22540 8504
rect 22580 8464 22581 8504
rect 22539 8455 22581 8464
rect 22732 8168 22772 8800
rect 22828 8168 22868 10135
rect 22924 9848 22964 10312
rect 23020 10193 23060 10396
rect 23019 10184 23061 10193
rect 23019 10144 23020 10184
rect 23060 10144 23061 10184
rect 23019 10135 23061 10144
rect 23116 10025 23156 10672
rect 23211 10184 23253 10193
rect 23211 10144 23212 10184
rect 23252 10144 23253 10184
rect 23211 10135 23253 10144
rect 23115 10016 23157 10025
rect 23115 9976 23116 10016
rect 23156 9976 23157 10016
rect 23115 9967 23157 9976
rect 22924 9808 23156 9848
rect 23019 9512 23061 9521
rect 23019 9472 23020 9512
rect 23060 9472 23061 9512
rect 23019 9463 23061 9472
rect 22923 8756 22965 8765
rect 22923 8716 22924 8756
rect 22964 8716 22965 8756
rect 22923 8707 22965 8716
rect 23020 8756 23060 9463
rect 23020 8707 23060 8716
rect 22924 8622 22964 8707
rect 23116 8588 23156 9808
rect 23020 8548 23156 8588
rect 23020 8429 23060 8548
rect 23019 8420 23061 8429
rect 23019 8380 23020 8420
rect 23060 8380 23061 8420
rect 23019 8371 23061 8380
rect 22924 8168 22964 8177
rect 22828 8128 22924 8168
rect 22732 8119 22772 8128
rect 22924 8119 22964 8128
rect 22443 8084 22485 8093
rect 22443 8044 22444 8084
rect 22484 8044 22485 8084
rect 22443 8035 22485 8044
rect 22060 8000 22100 8009
rect 22060 7841 22100 7960
rect 22059 7832 22101 7841
rect 22059 7792 22060 7832
rect 22100 7792 22101 7832
rect 22059 7783 22101 7792
rect 22060 7589 22100 7783
rect 22059 7580 22101 7589
rect 22059 7540 22060 7580
rect 22100 7540 22101 7580
rect 22059 7531 22101 7540
rect 21963 6656 22005 6665
rect 21963 6616 21964 6656
rect 22004 6616 22005 6656
rect 21963 6607 22005 6616
rect 22059 6572 22101 6581
rect 22059 6532 22060 6572
rect 22100 6532 22101 6572
rect 22059 6523 22101 6532
rect 21963 6488 22005 6497
rect 21963 6448 21964 6488
rect 22004 6448 22005 6488
rect 21963 6439 22005 6448
rect 22060 6488 22100 6523
rect 21772 5020 21908 5060
rect 21772 4229 21812 5020
rect 21964 4976 22004 6439
rect 21964 4927 22004 4936
rect 22060 4901 22100 6448
rect 22155 6488 22197 6497
rect 22155 6448 22156 6488
rect 22196 6448 22197 6488
rect 22155 6439 22197 6448
rect 22156 6354 22196 6439
rect 22444 5909 22484 8035
rect 22588 7958 22628 7967
rect 22588 7916 22628 7918
rect 22588 7876 22868 7916
rect 22828 7412 22868 7876
rect 22828 7363 22868 7372
rect 23020 7244 23060 8371
rect 23212 8177 23252 10135
rect 23308 8261 23348 10672
rect 23500 8840 23540 10672
rect 23692 8849 23732 10672
rect 23787 9512 23829 9521
rect 23787 9472 23788 9512
rect 23828 9472 23829 9512
rect 23787 9463 23829 9472
rect 23691 8840 23733 8849
rect 23500 8800 23636 8840
rect 23500 8672 23540 8681
rect 23307 8252 23349 8261
rect 23307 8212 23308 8252
rect 23348 8212 23349 8252
rect 23307 8203 23349 8212
rect 23211 8168 23253 8177
rect 23211 8128 23212 8168
rect 23252 8128 23253 8168
rect 23211 8119 23253 8128
rect 23116 7916 23156 7925
rect 23156 7876 23348 7916
rect 23116 7867 23156 7876
rect 22828 7204 23060 7244
rect 22635 7160 22677 7169
rect 22635 7120 22636 7160
rect 22676 7120 22677 7160
rect 22635 7111 22677 7120
rect 22636 7026 22676 7111
rect 22636 6488 22676 6497
rect 22539 6068 22581 6077
rect 22539 6028 22540 6068
rect 22580 6028 22581 6068
rect 22539 6019 22581 6028
rect 22443 5900 22485 5909
rect 22443 5860 22444 5900
rect 22484 5860 22485 5900
rect 22443 5851 22485 5860
rect 22444 5321 22484 5851
rect 22540 5648 22580 6019
rect 22540 5599 22580 5608
rect 22443 5312 22485 5321
rect 22443 5272 22444 5312
rect 22484 5272 22485 5312
rect 22443 5263 22485 5272
rect 22636 4985 22676 6448
rect 22731 6068 22773 6077
rect 22731 6028 22732 6068
rect 22772 6028 22773 6068
rect 22731 6019 22773 6028
rect 22732 5900 22772 6019
rect 22732 5851 22772 5860
rect 22443 4976 22485 4985
rect 22443 4936 22444 4976
rect 22484 4936 22485 4976
rect 22443 4927 22485 4936
rect 22635 4976 22677 4985
rect 22635 4936 22636 4976
rect 22676 4936 22677 4976
rect 22635 4927 22677 4936
rect 21867 4892 21909 4901
rect 21867 4852 21868 4892
rect 21908 4852 21909 4892
rect 21867 4843 21909 4852
rect 22059 4892 22101 4901
rect 22059 4852 22060 4892
rect 22100 4852 22101 4892
rect 22059 4843 22101 4852
rect 21868 4313 21908 4843
rect 22444 4842 22484 4927
rect 22059 4724 22101 4733
rect 22059 4684 22060 4724
rect 22100 4684 22101 4724
rect 22059 4675 22101 4684
rect 21867 4304 21909 4313
rect 21867 4264 21868 4304
rect 21908 4264 21909 4304
rect 21867 4255 21909 4264
rect 21771 4220 21813 4229
rect 21771 4180 21772 4220
rect 21812 4180 21813 4220
rect 21771 4171 21813 4180
rect 22060 2969 22100 4675
rect 22732 3464 22772 3473
rect 22059 2960 22101 2969
rect 22059 2920 22060 2960
rect 22100 2920 22101 2960
rect 22059 2911 22101 2920
rect 22060 2624 22100 2911
rect 22060 2575 22100 2584
rect 21676 2500 21812 2540
rect 21772 1793 21812 2500
rect 22539 2120 22581 2129
rect 22539 2080 22540 2120
rect 22580 2080 22581 2120
rect 22539 2071 22581 2080
rect 22732 2120 22772 3424
rect 22828 3464 22868 7204
rect 23308 6656 23348 7876
rect 23500 7505 23540 8632
rect 23499 7496 23541 7505
rect 23499 7456 23500 7496
rect 23540 7456 23541 7496
rect 23499 7447 23541 7456
rect 23308 6607 23348 6616
rect 23596 6581 23636 8800
rect 23691 8800 23692 8840
rect 23732 8800 23733 8840
rect 23691 8791 23733 8800
rect 23595 6572 23637 6581
rect 23595 6532 23596 6572
rect 23636 6532 23637 6572
rect 23595 6523 23637 6532
rect 23116 6474 23156 6483
rect 23116 6077 23156 6434
rect 23115 6068 23157 6077
rect 23115 6028 23116 6068
rect 23156 6028 23157 6068
rect 23115 6019 23157 6028
rect 22924 5648 22964 5657
rect 22924 5573 22964 5608
rect 23499 5648 23541 5657
rect 23499 5608 23500 5648
rect 23540 5608 23541 5648
rect 23499 5599 23541 5608
rect 22923 5564 22965 5573
rect 22923 5524 22924 5564
rect 22964 5524 22965 5564
rect 22923 5515 22965 5524
rect 22924 5405 22964 5515
rect 22923 5396 22965 5405
rect 22923 5356 22924 5396
rect 22964 5356 22965 5396
rect 22923 5347 22965 5356
rect 23500 5069 23540 5599
rect 23115 5060 23157 5069
rect 23115 5020 23116 5060
rect 23156 5020 23157 5060
rect 23115 5011 23157 5020
rect 23499 5060 23541 5069
rect 23499 5020 23500 5060
rect 23540 5020 23541 5060
rect 23499 5011 23541 5020
rect 22972 4966 23012 4975
rect 23012 4926 23060 4957
rect 23116 4926 23156 5011
rect 22972 4917 23060 4926
rect 22828 3415 22868 3424
rect 23020 2540 23060 4917
rect 23307 4220 23349 4229
rect 23307 4180 23308 4220
rect 23348 4180 23349 4220
rect 23307 4171 23349 4180
rect 23211 3464 23253 3473
rect 23211 3424 23212 3464
rect 23252 3424 23253 3464
rect 23211 3415 23253 3424
rect 23308 3464 23348 4171
rect 23308 3415 23348 3424
rect 23404 4136 23444 4145
rect 23212 2885 23252 3415
rect 23307 3128 23349 3137
rect 23307 3088 23308 3128
rect 23348 3088 23349 3128
rect 23307 3079 23349 3088
rect 23211 2876 23253 2885
rect 23211 2836 23212 2876
rect 23252 2836 23253 2876
rect 23211 2827 23253 2836
rect 23308 2801 23348 3079
rect 23404 2876 23444 4096
rect 23500 4136 23540 5011
rect 23788 4229 23828 9463
rect 23884 9353 23924 10672
rect 24076 10193 24116 10672
rect 24075 10184 24117 10193
rect 24075 10144 24076 10184
rect 24116 10144 24117 10184
rect 24075 10135 24117 10144
rect 23980 9605 24020 9636
rect 23979 9596 24021 9605
rect 23979 9556 23980 9596
rect 24020 9556 24021 9596
rect 23979 9547 24021 9556
rect 23980 9512 24020 9547
rect 23883 9344 23925 9353
rect 23883 9304 23884 9344
rect 23924 9304 23925 9344
rect 23883 9295 23925 9304
rect 23980 8933 24020 9472
rect 24172 9260 24212 9269
rect 24076 9220 24172 9260
rect 23979 8924 24021 8933
rect 23979 8884 23980 8924
rect 24020 8884 24021 8924
rect 23979 8875 24021 8884
rect 23883 8756 23925 8765
rect 24076 8756 24116 9220
rect 24172 9211 24212 9220
rect 24171 9092 24213 9101
rect 24171 9052 24172 9092
rect 24212 9052 24213 9092
rect 24171 9043 24213 9052
rect 23883 8716 23884 8756
rect 23924 8716 23925 8756
rect 23883 8707 23925 8716
rect 24028 8716 24116 8756
rect 24028 8714 24068 8716
rect 23884 7580 23924 8707
rect 24028 8665 24068 8674
rect 24172 8588 24212 9043
rect 24268 8765 24308 10672
rect 24364 9512 24404 9521
rect 24267 8756 24309 8765
rect 24267 8716 24268 8756
rect 24308 8716 24309 8756
rect 24267 8707 24309 8716
rect 24172 8539 24212 8548
rect 24364 8093 24404 9472
rect 24460 8933 24500 10672
rect 24555 10100 24597 10109
rect 24555 10060 24556 10100
rect 24596 10060 24597 10100
rect 24555 10051 24597 10060
rect 24459 8924 24501 8933
rect 24459 8884 24460 8924
rect 24500 8884 24501 8924
rect 24459 8875 24501 8884
rect 24556 8840 24596 10051
rect 24556 8791 24596 8800
rect 24363 8084 24405 8093
rect 24363 8044 24364 8084
rect 24404 8044 24405 8084
rect 24363 8035 24405 8044
rect 24076 8000 24116 8011
rect 24076 7925 24116 7960
rect 24075 7916 24117 7925
rect 24075 7876 24076 7916
rect 24116 7876 24117 7916
rect 24075 7867 24117 7876
rect 23884 7540 24020 7580
rect 23980 6656 24020 7540
rect 24364 7421 24404 8035
rect 24555 7496 24597 7505
rect 24555 7456 24556 7496
rect 24596 7456 24597 7496
rect 24555 7447 24597 7456
rect 24363 7412 24405 7421
rect 24363 7372 24364 7412
rect 24404 7372 24405 7412
rect 24363 7363 24405 7372
rect 24171 7160 24213 7169
rect 24171 7120 24172 7160
rect 24212 7120 24213 7160
rect 24171 7111 24213 7120
rect 24364 7160 24404 7169
rect 23884 6616 24020 6656
rect 23884 5984 23924 6616
rect 24075 6572 24117 6581
rect 24075 6532 24076 6572
rect 24116 6532 24117 6572
rect 24075 6523 24117 6532
rect 23980 6488 24020 6497
rect 23980 6068 24020 6448
rect 24076 6488 24116 6523
rect 24076 6437 24116 6448
rect 23980 6028 24116 6068
rect 23884 5944 24020 5984
rect 23884 4976 23924 4987
rect 23884 4901 23924 4936
rect 23883 4892 23925 4901
rect 23883 4852 23884 4892
rect 23924 4852 23925 4892
rect 23883 4843 23925 4852
rect 23884 4397 23924 4843
rect 23883 4388 23925 4397
rect 23883 4348 23884 4388
rect 23924 4348 23925 4388
rect 23883 4339 23925 4348
rect 23787 4220 23829 4229
rect 23884 4220 23924 4229
rect 23787 4180 23788 4220
rect 23828 4180 23884 4220
rect 23787 4171 23829 4180
rect 23884 4171 23924 4180
rect 23980 4220 24020 5944
rect 24076 5825 24116 6028
rect 24075 5816 24117 5825
rect 24075 5776 24076 5816
rect 24116 5776 24117 5816
rect 24075 5767 24117 5776
rect 23500 4087 23540 4096
rect 23788 4086 23828 4171
rect 23787 3548 23829 3557
rect 23787 3508 23788 3548
rect 23828 3508 23829 3548
rect 23787 3499 23829 3508
rect 23788 3464 23828 3499
rect 23980 3473 24020 4180
rect 24172 5648 24212 7111
rect 24364 6152 24404 7120
rect 24459 6488 24501 6497
rect 24459 6448 24460 6488
rect 24500 6448 24501 6488
rect 24459 6439 24501 6448
rect 24556 6488 24596 7447
rect 24460 6354 24500 6439
rect 24556 6329 24596 6448
rect 24555 6320 24597 6329
rect 24555 6280 24556 6320
rect 24596 6280 24597 6320
rect 24555 6271 24597 6280
rect 24364 6112 24500 6152
rect 24363 5816 24405 5825
rect 24363 5776 24364 5816
rect 24404 5776 24405 5816
rect 24363 5767 24405 5776
rect 24364 5682 24404 5767
rect 23788 3413 23828 3424
rect 23979 3464 24021 3473
rect 23979 3424 23980 3464
rect 24020 3424 24021 3464
rect 23979 3415 24021 3424
rect 23500 2876 23540 2885
rect 23404 2836 23500 2876
rect 23500 2827 23540 2836
rect 24172 2801 24212 5608
rect 24363 5312 24405 5321
rect 24363 5272 24364 5312
rect 24404 5272 24405 5312
rect 24363 5263 24405 5272
rect 24364 4136 24404 5263
rect 24460 5237 24500 6112
rect 24459 5228 24501 5237
rect 24459 5188 24460 5228
rect 24500 5188 24501 5228
rect 24459 5179 24501 5188
rect 24459 4136 24501 4145
rect 24364 4096 24460 4136
rect 24500 4096 24501 4136
rect 24459 4087 24501 4096
rect 24460 4002 24500 4087
rect 24460 3548 24500 3557
rect 24316 3422 24356 3431
rect 24316 3380 24356 3382
rect 24316 3340 24404 3380
rect 23307 2792 23349 2801
rect 23307 2752 23308 2792
rect 23348 2752 23349 2792
rect 23307 2743 23349 2752
rect 24171 2792 24213 2801
rect 24171 2752 24172 2792
rect 24212 2752 24213 2792
rect 24171 2743 24213 2752
rect 23308 2624 23348 2743
rect 23692 2633 23732 2718
rect 23308 2575 23348 2584
rect 23691 2624 23733 2633
rect 23691 2584 23692 2624
rect 23732 2584 23733 2624
rect 23691 2575 23733 2584
rect 23020 2500 23156 2540
rect 22732 2071 22772 2080
rect 22827 2120 22869 2129
rect 22827 2080 22828 2120
rect 22868 2080 22869 2120
rect 22827 2071 22869 2080
rect 22540 1952 22580 2071
rect 22540 1903 22580 1912
rect 21771 1784 21813 1793
rect 21771 1744 21772 1784
rect 21812 1744 21813 1784
rect 21771 1735 21813 1744
rect 21675 1616 21717 1625
rect 21675 1576 21676 1616
rect 21716 1576 21717 1616
rect 21675 1567 21717 1576
rect 21484 1231 21524 1240
rect 21676 1112 21716 1567
rect 21772 1457 21812 1735
rect 21771 1448 21813 1457
rect 21771 1408 21772 1448
rect 21812 1408 21813 1448
rect 21771 1399 21813 1408
rect 22539 1448 22581 1457
rect 22539 1408 22540 1448
rect 22580 1408 22581 1448
rect 22539 1399 22581 1408
rect 21676 701 21716 1072
rect 21675 692 21717 701
rect 21675 652 21676 692
rect 21716 652 21717 692
rect 21675 643 21717 652
rect 22540 80 22580 1399
rect 22828 1112 22868 2071
rect 22923 1952 22965 1961
rect 22923 1912 22924 1952
rect 22964 1912 22965 1952
rect 22923 1903 22965 1912
rect 22924 1818 22964 1903
rect 23116 1280 23156 2500
rect 24171 2120 24213 2129
rect 24171 2080 24172 2120
rect 24212 2080 24213 2120
rect 24171 2071 24213 2080
rect 24364 2120 24404 3340
rect 24460 2717 24500 3508
rect 24652 3053 24692 10672
rect 24748 8756 24788 8765
rect 24748 4061 24788 8716
rect 24844 6833 24884 10672
rect 25036 9932 25076 10672
rect 24940 9892 25076 9932
rect 24843 6824 24885 6833
rect 24843 6784 24844 6824
rect 24884 6784 24885 6824
rect 24843 6775 24885 6784
rect 24940 4304 24980 9892
rect 25035 9764 25077 9773
rect 25035 9724 25036 9764
rect 25076 9724 25077 9764
rect 25035 9715 25077 9724
rect 25036 8840 25076 9715
rect 25228 8924 25268 10672
rect 25036 8791 25076 8800
rect 25132 8884 25268 8924
rect 25132 7421 25172 8884
rect 25228 8756 25268 8765
rect 25131 7412 25173 7421
rect 25131 7372 25132 7412
rect 25172 7372 25173 7412
rect 25131 7363 25173 7372
rect 25131 7160 25173 7169
rect 25131 7120 25132 7160
rect 25172 7120 25173 7160
rect 25131 7111 25173 7120
rect 25036 6488 25076 6497
rect 25036 5321 25076 6448
rect 25035 5312 25077 5321
rect 25035 5272 25036 5312
rect 25076 5272 25077 5312
rect 25035 5263 25077 5272
rect 25132 4976 25172 7111
rect 25228 6665 25268 8716
rect 25323 8336 25365 8345
rect 25323 8296 25324 8336
rect 25364 8296 25365 8336
rect 25420 8336 25460 10672
rect 25612 9680 25652 10672
rect 25516 9640 25652 9680
rect 25516 9344 25556 9640
rect 25707 9596 25749 9605
rect 25612 9556 25708 9596
rect 25748 9556 25749 9596
rect 25612 9512 25652 9556
rect 25707 9547 25749 9556
rect 25612 9463 25652 9472
rect 25804 9428 25844 10672
rect 25708 9388 25844 9428
rect 25516 9304 25652 9344
rect 25515 9176 25557 9185
rect 25515 9136 25516 9176
rect 25556 9136 25557 9176
rect 25515 9127 25557 9136
rect 25516 8840 25556 9127
rect 25516 8791 25556 8800
rect 25612 8513 25652 9304
rect 25708 8924 25748 9388
rect 25996 9344 26036 10672
rect 26188 9428 26228 10672
rect 26188 9388 26324 9428
rect 25996 9304 26228 9344
rect 25804 9260 25844 9269
rect 25844 9220 26036 9260
rect 25804 9211 25844 9220
rect 25708 8884 25940 8924
rect 25708 8756 25748 8765
rect 25611 8504 25653 8513
rect 25611 8464 25612 8504
rect 25652 8464 25653 8504
rect 25611 8455 25653 8464
rect 25420 8296 25652 8336
rect 25323 8287 25365 8296
rect 25324 8000 25364 8287
rect 25324 7951 25364 7960
rect 25516 7748 25556 7757
rect 25516 7589 25556 7708
rect 25515 7580 25557 7589
rect 25515 7540 25516 7580
rect 25556 7540 25557 7580
rect 25515 7531 25557 7540
rect 25612 7412 25652 8296
rect 25708 7673 25748 8716
rect 25900 8168 25940 8884
rect 25996 8672 26036 9220
rect 26092 8681 26132 8766
rect 25996 8623 26036 8632
rect 26091 8672 26133 8681
rect 26091 8632 26092 8672
rect 26132 8632 26133 8672
rect 26091 8623 26133 8632
rect 26091 8504 26133 8513
rect 26091 8464 26092 8504
rect 26132 8464 26133 8504
rect 26091 8455 26133 8464
rect 25900 8128 26036 8168
rect 25804 8000 25844 8009
rect 25707 7664 25749 7673
rect 25707 7624 25708 7664
rect 25748 7624 25749 7664
rect 25707 7615 25749 7624
rect 25804 7589 25844 7960
rect 25899 8000 25941 8009
rect 25899 7960 25900 8000
rect 25940 7960 25941 8000
rect 25899 7951 25941 7960
rect 25900 7866 25940 7951
rect 25803 7580 25845 7589
rect 25803 7540 25804 7580
rect 25844 7540 25845 7580
rect 25803 7531 25845 7540
rect 25996 7412 26036 8128
rect 25612 7372 25748 7412
rect 25611 7160 25653 7169
rect 25611 7120 25612 7160
rect 25652 7120 25653 7160
rect 25611 7111 25653 7120
rect 25612 7026 25652 7111
rect 25515 6992 25557 7001
rect 25515 6952 25516 6992
rect 25556 6952 25557 6992
rect 25515 6943 25557 6952
rect 25227 6656 25269 6665
rect 25227 6616 25228 6656
rect 25268 6616 25269 6656
rect 25227 6607 25269 6616
rect 25516 6483 25556 6943
rect 25708 6824 25748 7372
rect 25900 7372 26036 7412
rect 26092 7412 26132 8455
rect 26188 7589 26228 9304
rect 26284 9101 26324 9388
rect 26283 9092 26325 9101
rect 26283 9052 26284 9092
rect 26324 9052 26325 9092
rect 26283 9043 26325 9052
rect 26283 8840 26325 8849
rect 26283 8800 26284 8840
rect 26324 8800 26325 8840
rect 26283 8791 26325 8800
rect 26284 8000 26324 8791
rect 26380 8429 26420 10672
rect 26572 8924 26612 10672
rect 26572 8884 26708 8924
rect 26475 8840 26517 8849
rect 26475 8800 26476 8840
rect 26516 8800 26517 8840
rect 26475 8791 26517 8800
rect 26476 8756 26516 8791
rect 26476 8681 26516 8716
rect 26571 8756 26613 8765
rect 26571 8716 26572 8756
rect 26612 8716 26613 8756
rect 26571 8707 26613 8716
rect 26475 8672 26517 8681
rect 26475 8632 26476 8672
rect 26516 8632 26517 8672
rect 26475 8623 26517 8632
rect 26476 8592 26516 8623
rect 26379 8420 26421 8429
rect 26379 8380 26380 8420
rect 26420 8380 26421 8420
rect 26379 8371 26421 8380
rect 26284 7951 26324 7960
rect 26380 8000 26420 8009
rect 26572 8000 26612 8707
rect 26420 7960 26612 8000
rect 26380 7951 26420 7960
rect 26283 7832 26325 7841
rect 26283 7792 26284 7832
rect 26324 7792 26325 7832
rect 26283 7783 26325 7792
rect 26187 7580 26229 7589
rect 26187 7540 26188 7580
rect 26228 7540 26229 7580
rect 26187 7531 26229 7540
rect 26092 7372 26228 7412
rect 25804 7001 25844 7086
rect 25803 6992 25845 7001
rect 25803 6952 25804 6992
rect 25844 6952 25845 6992
rect 25803 6943 25845 6952
rect 25708 6784 25844 6824
rect 25707 6656 25749 6665
rect 25707 6616 25708 6656
rect 25748 6616 25749 6656
rect 25707 6607 25749 6616
rect 25708 6522 25748 6607
rect 25516 6434 25556 6443
rect 25804 5816 25844 6784
rect 25612 5776 25844 5816
rect 25515 5060 25557 5069
rect 25515 5020 25516 5060
rect 25556 5020 25557 5060
rect 25515 5011 25557 5020
rect 25132 4927 25172 4936
rect 25324 4724 25364 4733
rect 24844 4264 24980 4304
rect 25036 4684 25324 4724
rect 24747 4052 24789 4061
rect 24747 4012 24748 4052
rect 24788 4012 24789 4052
rect 24747 4003 24789 4012
rect 24844 3632 24884 4264
rect 25036 4220 25076 4684
rect 25324 4675 25364 4684
rect 24988 4180 25076 4220
rect 24988 4178 25028 4180
rect 24988 4129 25028 4138
rect 25420 4136 25460 4145
rect 25228 4096 25420 4136
rect 25131 4052 25173 4061
rect 25131 4012 25132 4052
rect 25172 4012 25173 4052
rect 25131 4003 25173 4012
rect 25132 3918 25172 4003
rect 25228 3800 25268 4096
rect 25420 4087 25460 4096
rect 25516 4136 25556 5011
rect 25516 4087 25556 4096
rect 25132 3760 25268 3800
rect 24844 3592 24980 3632
rect 24844 3464 24884 3473
rect 24651 3044 24693 3053
rect 24651 3004 24652 3044
rect 24692 3004 24693 3044
rect 24651 2995 24693 3004
rect 24459 2708 24501 2717
rect 24459 2668 24460 2708
rect 24500 2668 24501 2708
rect 24459 2659 24501 2668
rect 24652 2633 24692 2718
rect 24651 2624 24693 2633
rect 24651 2584 24652 2624
rect 24692 2584 24693 2624
rect 24651 2575 24693 2584
rect 24555 2372 24597 2381
rect 24555 2332 24556 2372
rect 24596 2332 24597 2372
rect 24555 2323 24597 2332
rect 24364 2071 24404 2080
rect 24172 1952 24212 2071
rect 24556 1961 24596 2323
rect 24172 1903 24212 1912
rect 24555 1952 24597 1961
rect 24555 1912 24556 1952
rect 24596 1912 24597 1952
rect 24555 1903 24597 1912
rect 24556 1818 24596 1903
rect 23787 1700 23829 1709
rect 23787 1660 23788 1700
rect 23828 1660 23829 1700
rect 23787 1651 23829 1660
rect 23116 1231 23156 1240
rect 23691 1280 23733 1289
rect 23691 1240 23692 1280
rect 23732 1240 23733 1280
rect 23691 1231 23733 1240
rect 22924 1112 22964 1121
rect 22828 1072 22924 1112
rect 22924 1063 22964 1072
rect 23692 1112 23732 1231
rect 23692 1063 23732 1072
rect 23788 860 23828 1651
rect 24844 1121 24884 3424
rect 24940 3305 24980 3592
rect 24939 3296 24981 3305
rect 24939 3256 24940 3296
rect 24980 3256 24981 3296
rect 24939 3247 24981 3256
rect 24940 2969 24980 3247
rect 24939 2960 24981 2969
rect 24939 2920 24940 2960
rect 24980 2920 24981 2960
rect 24939 2911 24981 2920
rect 24939 2792 24981 2801
rect 24939 2752 24940 2792
rect 24980 2752 24981 2792
rect 24939 2743 24981 2752
rect 24940 1961 24980 2743
rect 24939 1952 24981 1961
rect 24939 1912 24940 1952
rect 24980 1912 24981 1952
rect 24939 1903 24981 1912
rect 24843 1112 24885 1121
rect 24843 1072 24844 1112
rect 24884 1072 24885 1112
rect 24843 1063 24885 1072
rect 24940 1112 24980 1903
rect 25132 1280 25172 3760
rect 25612 3221 25652 5776
rect 25803 5648 25845 5657
rect 25803 5608 25804 5648
rect 25844 5608 25845 5648
rect 25803 5599 25845 5608
rect 25804 5514 25844 5599
rect 25900 4220 25940 7372
rect 26092 7160 26132 7169
rect 26092 6488 26132 7120
rect 26188 6665 26228 7372
rect 26187 6656 26229 6665
rect 26187 6616 26188 6656
rect 26228 6616 26229 6656
rect 26187 6607 26229 6616
rect 26284 6488 26324 7783
rect 26379 7664 26421 7673
rect 26379 7624 26380 7664
rect 26420 7624 26421 7664
rect 26379 7615 26421 7624
rect 26092 6448 26324 6488
rect 25995 6320 26037 6329
rect 25995 6280 25996 6320
rect 26036 6280 26037 6320
rect 25995 6271 26037 6280
rect 25900 4171 25940 4180
rect 25996 4220 26036 6271
rect 26092 5993 26132 6448
rect 26091 5984 26133 5993
rect 26091 5944 26092 5984
rect 26132 5944 26133 5984
rect 26091 5935 26133 5944
rect 26380 5489 26420 7615
rect 26668 6497 26708 8884
rect 26764 8765 26804 10672
rect 26956 10529 26996 10672
rect 26955 10520 26997 10529
rect 26955 10480 26956 10520
rect 26996 10480 26997 10520
rect 26955 10471 26997 10480
rect 27148 9680 27188 10672
rect 27148 9640 27284 9680
rect 26859 9596 26901 9605
rect 26859 9556 26860 9596
rect 26900 9556 26901 9596
rect 26859 9547 26901 9556
rect 27051 9596 27093 9605
rect 27051 9556 27052 9596
rect 27092 9556 27188 9596
rect 27051 9547 27093 9556
rect 26763 8756 26805 8765
rect 26763 8716 26764 8756
rect 26804 8716 26805 8756
rect 26763 8707 26805 8716
rect 26860 8261 26900 9547
rect 27148 9512 27188 9556
rect 27148 9463 27188 9472
rect 26956 9260 26996 9269
rect 26956 8849 26996 9220
rect 27147 8924 27189 8933
rect 27147 8884 27148 8924
rect 27188 8884 27189 8924
rect 27147 8875 27189 8884
rect 26955 8840 26997 8849
rect 26955 8800 26956 8840
rect 26996 8800 26997 8840
rect 26955 8791 26997 8800
rect 27052 8672 27092 8681
rect 26859 8252 26901 8261
rect 26859 8212 26860 8252
rect 26900 8212 26901 8252
rect 26859 8203 26901 8212
rect 26955 8168 26997 8177
rect 26955 8128 26956 8168
rect 26996 8128 26997 8168
rect 26955 8119 26997 8128
rect 26860 8000 26900 8009
rect 26860 7673 26900 7960
rect 26859 7664 26901 7673
rect 26859 7624 26860 7664
rect 26900 7624 26901 7664
rect 26859 7615 26901 7624
rect 26859 7328 26901 7337
rect 26859 7288 26860 7328
rect 26900 7288 26901 7328
rect 26859 7279 26901 7288
rect 26667 6488 26709 6497
rect 26667 6448 26668 6488
rect 26708 6448 26709 6488
rect 26667 6439 26709 6448
rect 26860 5648 26900 7279
rect 26956 5816 26996 8119
rect 27052 7673 27092 8632
rect 27051 7664 27093 7673
rect 27051 7624 27052 7664
rect 27092 7624 27093 7664
rect 27051 7615 27093 7624
rect 27148 6749 27188 8875
rect 27244 8261 27284 9640
rect 27340 9521 27380 10672
rect 27339 9512 27381 9521
rect 27339 9472 27340 9512
rect 27380 9472 27381 9512
rect 27339 9463 27381 9472
rect 27532 9344 27572 10672
rect 27724 10613 27764 10672
rect 27723 10604 27765 10613
rect 27723 10564 27724 10604
rect 27764 10564 27765 10604
rect 27723 10555 27765 10564
rect 27532 9304 27668 9344
rect 27339 9092 27381 9101
rect 27339 9052 27340 9092
rect 27380 9052 27381 9092
rect 27339 9043 27381 9052
rect 27340 8345 27380 9043
rect 27531 8840 27573 8849
rect 27531 8800 27532 8840
rect 27572 8800 27573 8840
rect 27531 8791 27573 8800
rect 27532 8686 27572 8791
rect 27532 8637 27572 8646
rect 27339 8336 27381 8345
rect 27339 8296 27340 8336
rect 27380 8296 27381 8336
rect 27339 8287 27381 8296
rect 27243 8252 27285 8261
rect 27243 8212 27244 8252
rect 27284 8212 27285 8252
rect 27243 8203 27285 8212
rect 27340 8084 27380 8287
rect 27531 8168 27573 8177
rect 27531 8128 27532 8168
rect 27572 8128 27573 8168
rect 27531 8119 27573 8128
rect 27244 8044 27380 8084
rect 27244 7160 27284 8044
rect 27532 8034 27572 8119
rect 27388 7958 27428 7967
rect 27388 7916 27428 7918
rect 27388 7876 27572 7916
rect 27532 7412 27572 7876
rect 27532 7363 27572 7372
rect 27340 7160 27380 7169
rect 27244 7120 27340 7160
rect 27380 7120 27476 7160
rect 27340 7111 27380 7120
rect 27147 6740 27189 6749
rect 27147 6700 27148 6740
rect 27188 6700 27189 6740
rect 27147 6691 27189 6700
rect 27148 6488 27188 6497
rect 27148 5900 27188 6448
rect 27244 6488 27284 6497
rect 27244 6161 27284 6448
rect 27243 6152 27285 6161
rect 27243 6112 27244 6152
rect 27284 6112 27285 6152
rect 27243 6103 27285 6112
rect 27244 5900 27284 5909
rect 27148 5860 27244 5900
rect 27244 5851 27284 5860
rect 26956 5776 27188 5816
rect 27148 5732 27188 5776
rect 27148 5692 27284 5732
rect 27052 5648 27092 5657
rect 26860 5608 27052 5648
rect 27052 5599 27092 5608
rect 26379 5480 26421 5489
rect 26379 5440 26380 5480
rect 26420 5440 26421 5480
rect 26379 5431 26421 5440
rect 27051 5480 27093 5489
rect 27051 5440 27052 5480
rect 27092 5440 27093 5480
rect 27051 5431 27093 5440
rect 26091 5060 26133 5069
rect 26091 5020 26092 5060
rect 26132 5020 26133 5060
rect 26091 5011 26133 5020
rect 25996 3557 26036 4180
rect 25995 3548 26037 3557
rect 25995 3508 25996 3548
rect 26036 3508 26037 3548
rect 25995 3499 26037 3508
rect 25707 3464 25749 3473
rect 25707 3424 25708 3464
rect 25748 3424 25749 3464
rect 25707 3415 25749 3424
rect 25900 3464 25940 3475
rect 25708 3330 25748 3415
rect 25900 3389 25940 3424
rect 25899 3380 25941 3389
rect 25899 3340 25900 3380
rect 25940 3340 25941 3380
rect 25899 3331 25941 3340
rect 25611 3212 25653 3221
rect 25611 3172 25612 3212
rect 25652 3172 25653 3212
rect 25611 3163 25653 3172
rect 25611 2960 25653 2969
rect 25611 2920 25612 2960
rect 25652 2920 25653 2960
rect 25611 2911 25653 2920
rect 25516 2624 25556 2633
rect 25516 2204 25556 2584
rect 25612 2624 25652 2911
rect 25900 2717 25940 3331
rect 25899 2708 25941 2717
rect 25899 2668 25900 2708
rect 25940 2668 25941 2708
rect 25899 2659 25941 2668
rect 25996 2708 26036 3499
rect 25996 2659 26036 2668
rect 26092 2708 26132 5011
rect 26571 4556 26613 4565
rect 26571 4516 26572 4556
rect 26612 4516 26613 4556
rect 26571 4507 26613 4516
rect 26475 4136 26517 4145
rect 26572 4136 26612 4507
rect 26475 4096 26476 4136
rect 26516 4096 26612 4136
rect 26475 4087 26517 4096
rect 26476 4002 26516 4087
rect 26475 3548 26517 3557
rect 26475 3508 26476 3548
rect 26516 3508 26517 3548
rect 26475 3499 26517 3508
rect 26092 2659 26132 2668
rect 25612 2575 25652 2584
rect 25516 2164 26036 2204
rect 25996 2120 26036 2164
rect 26476 2129 26516 3499
rect 26572 2624 26612 4096
rect 26572 2575 26612 2584
rect 26956 4141 26996 4150
rect 26956 2540 26996 4101
rect 27052 3968 27092 5431
rect 27148 4976 27188 4985
rect 27148 4136 27188 4936
rect 27244 4976 27284 5692
rect 27244 4927 27284 4936
rect 27148 4096 27380 4136
rect 27148 3968 27188 3977
rect 27052 3928 27148 3968
rect 27148 3919 27188 3928
rect 27340 3632 27380 4096
rect 27340 3583 27380 3592
rect 27436 3557 27476 7120
rect 27531 6740 27573 6749
rect 27531 6700 27532 6740
rect 27572 6700 27573 6740
rect 27628 6740 27668 9304
rect 27916 8672 27956 10672
rect 28108 8924 28148 10672
rect 27820 8632 27956 8672
rect 28012 8884 28148 8924
rect 27723 8504 27765 8513
rect 27723 8464 27724 8504
rect 27764 8464 27765 8504
rect 27723 8455 27765 8464
rect 27724 8370 27764 8455
rect 27723 7160 27765 7169
rect 27723 7120 27724 7160
rect 27764 7120 27765 7160
rect 27723 7111 27765 7120
rect 27724 7026 27764 7111
rect 27628 6700 27764 6740
rect 27531 6691 27573 6700
rect 27532 6488 27572 6691
rect 27628 6488 27668 6497
rect 27532 6448 27628 6488
rect 27628 4976 27668 6448
rect 27724 6488 27764 6700
rect 27724 4985 27764 6448
rect 27820 5657 27860 8632
rect 27915 8504 27957 8513
rect 27915 8464 27916 8504
rect 27956 8464 27957 8504
rect 27915 8455 27957 8464
rect 27916 8370 27956 8455
rect 28012 8168 28052 8884
rect 28108 8756 28148 8765
rect 28108 8177 28148 8716
rect 27916 8128 28052 8168
rect 28107 8168 28149 8177
rect 28107 8128 28108 8168
rect 28148 8128 28149 8168
rect 27819 5648 27861 5657
rect 27819 5608 27820 5648
rect 27860 5608 27861 5648
rect 27819 5599 27861 5608
rect 27916 5069 27956 8128
rect 28107 8119 28149 8128
rect 28011 8000 28053 8009
rect 28011 7960 28012 8000
rect 28052 7960 28053 8000
rect 28011 7951 28053 7960
rect 28203 8000 28245 8009
rect 28203 7960 28204 8000
rect 28244 7960 28245 8000
rect 28203 7951 28245 7960
rect 28012 6161 28052 7951
rect 28204 7757 28244 7951
rect 28203 7748 28245 7757
rect 28203 7708 28204 7748
rect 28244 7708 28245 7748
rect 28203 7699 28245 7708
rect 28300 7673 28340 10672
rect 28396 9512 28436 9521
rect 28396 9353 28436 9472
rect 28395 9344 28437 9353
rect 28395 9304 28396 9344
rect 28436 9304 28437 9344
rect 28395 9295 28437 9304
rect 28299 7664 28341 7673
rect 28299 7624 28300 7664
rect 28340 7624 28341 7664
rect 28299 7615 28341 7624
rect 28396 7160 28436 9295
rect 28108 7120 28436 7160
rect 28011 6152 28053 6161
rect 28011 6112 28012 6152
rect 28052 6112 28053 6152
rect 28011 6103 28053 6112
rect 28011 5984 28053 5993
rect 28011 5944 28012 5984
rect 28052 5944 28053 5984
rect 28011 5935 28053 5944
rect 27915 5060 27957 5069
rect 27915 5020 27916 5060
rect 27956 5020 27957 5060
rect 27915 5011 27957 5020
rect 27628 4817 27668 4936
rect 27723 4976 27765 4985
rect 27723 4936 27724 4976
rect 27764 4936 27765 4976
rect 27723 4927 27765 4936
rect 27724 4842 27764 4927
rect 27627 4808 27669 4817
rect 27627 4768 27628 4808
rect 27668 4768 27669 4808
rect 27627 4759 27669 4768
rect 27532 4136 27572 4145
rect 27532 3893 27572 4096
rect 28012 4061 28052 5935
rect 28011 4052 28053 4061
rect 28011 4012 28012 4052
rect 28052 4012 28053 4052
rect 28011 4003 28053 4012
rect 27531 3884 27573 3893
rect 27531 3844 27532 3884
rect 27572 3844 27573 3884
rect 27531 3835 27573 3844
rect 27147 3548 27189 3557
rect 27147 3508 27148 3548
rect 27188 3508 27189 3548
rect 27147 3499 27189 3508
rect 27435 3548 27477 3557
rect 27435 3508 27436 3548
rect 27476 3508 27477 3548
rect 27435 3499 27477 3508
rect 27148 3464 27188 3499
rect 27148 3413 27188 3424
rect 27627 3464 27669 3473
rect 27627 3424 27628 3464
rect 27668 3424 27669 3464
rect 27627 3415 27669 3424
rect 27243 3380 27285 3389
rect 27243 3340 27244 3380
rect 27284 3340 27285 3380
rect 27243 3331 27285 3340
rect 27100 2633 27140 2642
rect 27140 2593 27188 2624
rect 27100 2584 27188 2593
rect 26860 2500 26996 2540
rect 25996 2071 26036 2080
rect 26475 2120 26517 2129
rect 26475 2080 26476 2120
rect 26516 2080 26517 2120
rect 26475 2071 26517 2080
rect 26187 2036 26229 2045
rect 26187 1996 26188 2036
rect 26228 1996 26229 2036
rect 26187 1987 26229 1996
rect 25803 1952 25845 1961
rect 25803 1912 25804 1952
rect 25844 1912 25845 1952
rect 25803 1903 25845 1912
rect 26188 1952 26228 1987
rect 25804 1818 25844 1903
rect 26188 1901 26228 1912
rect 26667 1952 26709 1961
rect 26667 1912 26668 1952
rect 26708 1912 26709 1952
rect 26667 1903 26709 1912
rect 26475 1784 26517 1793
rect 26475 1744 26476 1784
rect 26516 1744 26517 1784
rect 26475 1735 26517 1744
rect 26476 1289 26516 1735
rect 25132 1231 25172 1240
rect 26475 1280 26517 1289
rect 26475 1240 26476 1280
rect 26516 1240 26517 1280
rect 26475 1231 26517 1240
rect 25419 1196 25461 1205
rect 25419 1156 25420 1196
rect 25460 1156 25461 1196
rect 25419 1147 25461 1156
rect 24940 1063 24980 1072
rect 25420 1112 25460 1147
rect 25420 1061 25460 1072
rect 26668 1112 26708 1903
rect 26860 1280 26900 2500
rect 27148 1700 27188 2584
rect 27244 2540 27284 3331
rect 27628 3330 27668 3415
rect 27916 3212 27956 3221
rect 27531 2960 27573 2969
rect 27531 2920 27532 2960
rect 27572 2920 27573 2960
rect 27531 2911 27573 2920
rect 27244 2491 27284 2500
rect 27532 2624 27572 2911
rect 27916 2633 27956 3172
rect 27435 1952 27477 1961
rect 27435 1912 27436 1952
rect 27476 1912 27477 1952
rect 27435 1903 27477 1912
rect 27436 1818 27476 1903
rect 27532 1877 27572 2584
rect 27915 2624 27957 2633
rect 27915 2584 27916 2624
rect 27956 2584 27957 2624
rect 27915 2575 27957 2584
rect 28108 2540 28148 7120
rect 28204 6581 28244 6612
rect 28203 6572 28245 6581
rect 28203 6532 28204 6572
rect 28244 6532 28245 6572
rect 28203 6523 28245 6532
rect 28204 6488 28244 6523
rect 28204 4976 28244 6448
rect 28492 6413 28532 10672
rect 28684 8345 28724 10672
rect 28683 8336 28725 8345
rect 28683 8296 28684 8336
rect 28724 8296 28725 8336
rect 28683 8287 28725 8296
rect 28876 7505 28916 10672
rect 29068 9185 29108 10672
rect 29067 9176 29109 9185
rect 29067 9136 29068 9176
rect 29108 9136 29109 9176
rect 29067 9127 29109 9136
rect 29260 9008 29300 10672
rect 29355 9596 29397 9605
rect 29355 9556 29356 9596
rect 29396 9556 29397 9596
rect 29355 9547 29397 9556
rect 28972 8968 29300 9008
rect 28875 7496 28917 7505
rect 28875 7456 28876 7496
rect 28916 7456 28917 7496
rect 28875 7447 28917 7456
rect 28972 7337 29012 8968
rect 29068 8672 29108 8681
rect 29068 8513 29108 8632
rect 29163 8672 29205 8681
rect 29163 8632 29164 8672
rect 29204 8632 29205 8672
rect 29163 8623 29205 8632
rect 29164 8538 29204 8623
rect 29067 8504 29109 8513
rect 29067 8464 29068 8504
rect 29108 8464 29109 8504
rect 29067 8455 29109 8464
rect 29356 8168 29396 9547
rect 29452 8849 29492 10672
rect 29644 9596 29684 10672
rect 29836 9680 29876 10672
rect 29836 9631 29876 9640
rect 30028 9680 30068 10672
rect 30220 9680 30260 10672
rect 30412 10025 30452 10672
rect 30411 10016 30453 10025
rect 30411 9976 30412 10016
rect 30452 9976 30453 10016
rect 30411 9967 30453 9976
rect 30507 9848 30549 9857
rect 30507 9808 30508 9848
rect 30548 9808 30549 9848
rect 30507 9799 30549 9808
rect 30412 9680 30452 9689
rect 30220 9640 30412 9680
rect 30028 9631 30068 9640
rect 30412 9631 30452 9640
rect 29644 9556 29780 9596
rect 29740 9512 29780 9556
rect 30411 9512 30453 9521
rect 29740 9472 29876 9512
rect 29644 9428 29684 9437
rect 29684 9388 29780 9428
rect 29644 9379 29684 9388
rect 29643 9176 29685 9185
rect 29643 9136 29644 9176
rect 29684 9136 29685 9176
rect 29643 9127 29685 9136
rect 29451 8840 29493 8849
rect 29451 8800 29452 8840
rect 29492 8800 29493 8840
rect 29451 8791 29493 8800
rect 29547 8756 29589 8765
rect 29547 8716 29548 8756
rect 29588 8716 29589 8756
rect 29547 8707 29589 8716
rect 29644 8756 29684 9127
rect 29548 8622 29588 8707
rect 29451 8504 29493 8513
rect 29451 8464 29452 8504
rect 29492 8464 29493 8504
rect 29451 8455 29493 8464
rect 29068 8128 29396 8168
rect 29452 8168 29492 8455
rect 28971 7328 29013 7337
rect 28971 7288 28972 7328
rect 29012 7288 29013 7328
rect 28971 7279 29013 7288
rect 28972 7160 29012 7169
rect 29068 7160 29108 8128
rect 29452 8119 29492 8128
rect 29547 8168 29589 8177
rect 29547 8128 29548 8168
rect 29588 8128 29589 8168
rect 29547 8119 29589 8128
rect 29260 8000 29300 8009
rect 29548 8000 29588 8119
rect 29300 7960 29588 8000
rect 29260 7951 29300 7960
rect 29355 7580 29397 7589
rect 29355 7540 29356 7580
rect 29396 7540 29397 7580
rect 29355 7531 29397 7540
rect 29547 7580 29589 7589
rect 29547 7540 29548 7580
rect 29588 7540 29589 7580
rect 29547 7531 29589 7540
rect 29259 7412 29301 7421
rect 29259 7372 29260 7412
rect 29300 7372 29301 7412
rect 29259 7363 29301 7372
rect 29012 7120 29108 7160
rect 28972 7111 29012 7120
rect 28683 6992 28725 7001
rect 28683 6952 28684 6992
rect 28724 6952 28725 6992
rect 28683 6943 28725 6952
rect 29163 6992 29205 7001
rect 29163 6952 29164 6992
rect 29204 6952 29205 6992
rect 29163 6943 29205 6952
rect 28684 6483 28724 6943
rect 29164 6858 29204 6943
rect 28876 6572 28916 6581
rect 28684 6434 28724 6443
rect 28780 6532 28876 6572
rect 28491 6404 28533 6413
rect 28491 6364 28492 6404
rect 28532 6364 28533 6404
rect 28491 6355 28533 6364
rect 28780 5900 28820 6532
rect 28876 6523 28916 6532
rect 29260 6497 29300 7363
rect 29164 6488 29204 6497
rect 28971 6404 29013 6413
rect 28971 6364 28972 6404
rect 29012 6364 29013 6404
rect 28971 6355 29013 6364
rect 28396 5860 28820 5900
rect 28299 5480 28341 5489
rect 28299 5440 28300 5480
rect 28340 5440 28341 5480
rect 28299 5431 28341 5440
rect 28300 5346 28340 5431
rect 28299 5060 28341 5069
rect 28299 5020 28300 5060
rect 28340 5020 28341 5060
rect 28299 5011 28341 5020
rect 28204 4927 28244 4936
rect 28300 4565 28340 5011
rect 28299 4556 28341 4565
rect 28299 4516 28300 4556
rect 28340 4516 28341 4556
rect 28299 4507 28341 4516
rect 28396 4481 28436 5860
rect 28492 5732 28532 5741
rect 28532 5692 28820 5732
rect 28492 5683 28532 5692
rect 28780 5144 28820 5692
rect 28876 5648 28916 5657
rect 28876 5312 28916 5608
rect 28972 5648 29012 6355
rect 29012 5608 29108 5648
rect 28972 5599 29012 5608
rect 28876 5272 29012 5312
rect 28876 5144 28916 5153
rect 28780 5104 28876 5144
rect 28876 5095 28916 5104
rect 28732 4966 28772 4975
rect 28772 4926 28916 4957
rect 28732 4917 28916 4926
rect 28395 4472 28437 4481
rect 28395 4432 28396 4472
rect 28436 4432 28437 4472
rect 28395 4423 28437 4432
rect 28780 4136 28820 4145
rect 28492 4096 28780 4136
rect 28299 2624 28341 2633
rect 28299 2584 28300 2624
rect 28340 2584 28341 2624
rect 28299 2575 28341 2584
rect 28012 2500 28148 2540
rect 27916 1952 27956 1963
rect 27916 1877 27956 1912
rect 27531 1868 27573 1877
rect 27531 1828 27532 1868
rect 27572 1828 27573 1868
rect 27531 1819 27573 1828
rect 27915 1868 27957 1877
rect 27915 1828 27916 1868
rect 27956 1828 27957 1868
rect 27915 1819 27957 1828
rect 27628 1700 27668 1709
rect 27148 1660 27628 1700
rect 27628 1651 27668 1660
rect 26860 1231 26900 1240
rect 27628 1205 27668 1236
rect 27627 1196 27669 1205
rect 27627 1156 27628 1196
rect 27668 1156 27669 1196
rect 27627 1147 27669 1156
rect 26668 1063 26708 1072
rect 27628 1112 27668 1147
rect 25995 944 26037 953
rect 25995 904 25996 944
rect 26036 904 26037 944
rect 25995 895 26037 904
rect 23692 820 23828 860
rect 23692 80 23732 820
rect 24843 524 24885 533
rect 24843 484 24844 524
rect 24884 484 24885 524
rect 24843 475 24885 484
rect 24844 80 24884 475
rect 25996 80 26036 895
rect 27147 692 27189 701
rect 27147 652 27148 692
rect 27188 652 27189 692
rect 27147 643 27189 652
rect 27148 80 27188 643
rect 27628 617 27668 1072
rect 28012 785 28052 2500
rect 28107 1868 28149 1877
rect 28107 1828 28108 1868
rect 28148 1828 28149 1868
rect 28107 1819 28149 1828
rect 28108 1625 28148 1819
rect 28107 1616 28149 1625
rect 28107 1576 28108 1616
rect 28148 1576 28149 1616
rect 28107 1567 28149 1576
rect 28011 776 28053 785
rect 28011 736 28012 776
rect 28052 736 28053 776
rect 28011 727 28053 736
rect 27627 608 27669 617
rect 27627 568 27628 608
rect 27668 568 27669 608
rect 27627 559 27669 568
rect 28300 80 28340 2575
rect 28492 1961 28532 4096
rect 28780 4087 28820 4096
rect 28683 3548 28725 3557
rect 28683 3508 28684 3548
rect 28724 3508 28725 3548
rect 28683 3499 28725 3508
rect 28587 3464 28629 3473
rect 28587 3424 28588 3464
rect 28628 3424 28629 3464
rect 28587 3415 28629 3424
rect 28588 3330 28628 3415
rect 28587 2876 28629 2885
rect 28587 2836 28588 2876
rect 28628 2836 28629 2876
rect 28587 2827 28629 2836
rect 28491 1952 28533 1961
rect 28491 1912 28492 1952
rect 28532 1912 28533 1952
rect 28491 1903 28533 1912
rect 28588 953 28628 2827
rect 28684 2624 28724 3499
rect 28779 3212 28821 3221
rect 28779 3172 28780 3212
rect 28820 3172 28821 3212
rect 28779 3163 28821 3172
rect 28780 3078 28820 3163
rect 28876 2876 28916 4917
rect 28972 4892 29012 5272
rect 29068 5060 29108 5608
rect 29164 5144 29204 6448
rect 29259 6488 29301 6497
rect 29259 6448 29260 6488
rect 29300 6448 29301 6488
rect 29259 6439 29301 6448
rect 29260 6354 29300 6439
rect 29356 5732 29396 7531
rect 29451 6572 29493 6581
rect 29451 6532 29452 6572
rect 29492 6532 29493 6572
rect 29451 6523 29493 6532
rect 29356 5683 29396 5692
rect 29452 5732 29492 6523
rect 29452 5683 29492 5692
rect 29164 5104 29396 5144
rect 29068 5020 29300 5060
rect 29260 4976 29300 5020
rect 29164 4957 29204 4966
rect 29260 4927 29300 4936
rect 28972 4852 29108 4892
rect 28971 4388 29013 4397
rect 28971 4348 28972 4388
rect 29012 4348 29013 4388
rect 28971 4339 29013 4348
rect 28972 4254 29012 4339
rect 28971 3380 29013 3389
rect 28971 3340 28972 3380
rect 29012 3340 29013 3380
rect 28971 3331 29013 3340
rect 28972 3246 29012 3331
rect 28972 2876 29012 2904
rect 28876 2836 28972 2876
rect 28972 2827 29012 2836
rect 28780 2624 28820 2633
rect 28684 2584 28780 2624
rect 28780 2575 28820 2584
rect 28875 1952 28917 1961
rect 28875 1912 28876 1952
rect 28916 1912 28917 1952
rect 28875 1903 28917 1912
rect 28876 1625 28916 1903
rect 28875 1616 28917 1625
rect 28875 1576 28876 1616
rect 28916 1576 28917 1616
rect 28875 1567 28917 1576
rect 28876 1112 28916 1567
rect 29068 1280 29108 4852
rect 29164 4397 29204 4917
rect 29356 4472 29396 5104
rect 29260 4432 29396 4472
rect 29163 4388 29205 4397
rect 29163 4348 29164 4388
rect 29204 4348 29205 4388
rect 29163 4339 29205 4348
rect 29260 2120 29300 4432
rect 29452 4304 29492 4313
rect 29356 3464 29396 3475
rect 29356 3389 29396 3424
rect 29355 3380 29397 3389
rect 29355 3340 29356 3380
rect 29396 3340 29397 3380
rect 29355 3331 29397 3340
rect 29356 2465 29396 3331
rect 29355 2456 29397 2465
rect 29355 2416 29356 2456
rect 29396 2416 29397 2456
rect 29355 2407 29397 2416
rect 29356 2120 29396 2129
rect 29260 2080 29356 2120
rect 29356 2071 29396 2080
rect 29164 1952 29204 1961
rect 29164 1625 29204 1912
rect 29163 1616 29205 1625
rect 29163 1576 29164 1616
rect 29204 1576 29205 1616
rect 29163 1567 29205 1576
rect 29068 1231 29108 1240
rect 29452 1196 29492 4264
rect 29548 3557 29588 7531
rect 29644 6581 29684 8716
rect 29740 8513 29780 9388
rect 29739 8504 29781 8513
rect 29739 8464 29740 8504
rect 29780 8464 29781 8504
rect 29739 8455 29781 8464
rect 29739 8000 29781 8009
rect 29739 7960 29740 8000
rect 29780 7960 29781 8000
rect 29739 7951 29781 7960
rect 29740 7866 29780 7951
rect 29739 7664 29781 7673
rect 29739 7624 29740 7664
rect 29780 7624 29781 7664
rect 29739 7615 29781 7624
rect 29643 6572 29685 6581
rect 29643 6532 29644 6572
rect 29684 6532 29685 6572
rect 29643 6523 29685 6532
rect 29644 6488 29684 6523
rect 29644 6438 29684 6448
rect 29740 6488 29780 7615
rect 29740 6439 29780 6448
rect 29643 4976 29685 4985
rect 29643 4936 29644 4976
rect 29684 4936 29685 4976
rect 29643 4927 29685 4936
rect 29644 4842 29684 4927
rect 29740 4892 29780 4903
rect 29740 4817 29780 4852
rect 29739 4808 29781 4817
rect 29739 4768 29740 4808
rect 29780 4768 29781 4808
rect 29739 4759 29781 4768
rect 29547 3548 29589 3557
rect 29547 3508 29548 3548
rect 29588 3508 29589 3548
rect 29547 3499 29589 3508
rect 29643 2708 29685 2717
rect 29643 2668 29644 2708
rect 29684 2668 29685 2708
rect 29643 2659 29685 2668
rect 29644 2624 29684 2659
rect 29644 2573 29684 2584
rect 29547 2204 29589 2213
rect 29547 2164 29548 2204
rect 29588 2164 29589 2204
rect 29547 2155 29589 2164
rect 29548 1961 29588 2155
rect 29547 1952 29589 1961
rect 29547 1912 29548 1952
rect 29588 1912 29589 1952
rect 29547 1903 29589 1912
rect 29548 1818 29588 1903
rect 29836 1364 29876 9472
rect 30411 9472 30412 9512
rect 30452 9472 30453 9512
rect 30411 9463 30453 9472
rect 30220 9428 30260 9437
rect 29931 8672 29973 8681
rect 29931 8632 29932 8672
rect 29972 8632 29973 8672
rect 29931 8623 29973 8632
rect 30123 8672 30165 8681
rect 30123 8632 30124 8672
rect 30164 8632 30165 8672
rect 30123 8623 30165 8632
rect 29932 7589 29972 8623
rect 30027 8504 30069 8513
rect 30027 8464 30028 8504
rect 30068 8464 30069 8504
rect 30027 8455 30069 8464
rect 29931 7580 29973 7589
rect 29931 7540 29932 7580
rect 29972 7540 29973 7580
rect 29931 7531 29973 7540
rect 29932 5639 29972 5659
rect 29932 5573 29972 5599
rect 29931 5564 29973 5573
rect 29931 5524 29932 5564
rect 29972 5524 29973 5564
rect 29931 5515 29973 5524
rect 30028 4649 30068 8455
rect 30124 6488 30164 8623
rect 30220 8177 30260 9388
rect 30219 8168 30261 8177
rect 30219 8128 30220 8168
rect 30260 8128 30261 8168
rect 30219 8119 30261 8128
rect 30219 7916 30261 7925
rect 30219 7876 30220 7916
rect 30260 7876 30261 7916
rect 30219 7867 30261 7876
rect 30220 7160 30260 7867
rect 30220 7111 30260 7120
rect 30220 6488 30260 6497
rect 30124 6448 30220 6488
rect 30220 5573 30260 6448
rect 30412 6077 30452 9463
rect 30411 6068 30453 6077
rect 30411 6028 30412 6068
rect 30452 6028 30453 6068
rect 30411 6019 30453 6028
rect 30508 5816 30548 9799
rect 30604 9596 30644 10672
rect 30796 10184 30836 10672
rect 30796 10144 30932 10184
rect 30795 10016 30837 10025
rect 30795 9976 30796 10016
rect 30836 9976 30837 10016
rect 30795 9967 30837 9976
rect 30796 9680 30836 9967
rect 30796 9631 30836 9640
rect 30604 9556 30740 9596
rect 30700 9512 30740 9556
rect 30892 9521 30932 10144
rect 30988 9689 31028 10672
rect 30987 9680 31029 9689
rect 31180 9680 31220 10672
rect 31372 9857 31412 10672
rect 31564 10529 31604 10672
rect 31563 10520 31605 10529
rect 31756 10520 31796 10672
rect 31563 10480 31564 10520
rect 31604 10480 31605 10520
rect 31563 10471 31605 10480
rect 31660 10480 31796 10520
rect 31851 10520 31893 10529
rect 31851 10480 31852 10520
rect 31892 10480 31893 10520
rect 31563 10268 31605 10277
rect 31563 10228 31564 10268
rect 31604 10228 31605 10268
rect 31563 10219 31605 10228
rect 31371 9848 31413 9857
rect 31371 9808 31372 9848
rect 31412 9808 31413 9848
rect 31371 9799 31413 9808
rect 30987 9640 30988 9680
rect 31028 9640 31029 9680
rect 30987 9631 31029 9640
rect 31084 9640 31220 9680
rect 31467 9680 31509 9689
rect 31467 9640 31468 9680
rect 31508 9640 31509 9680
rect 30891 9512 30933 9521
rect 30997 9512 31039 9521
rect 30700 9472 30836 9512
rect 30604 9428 30644 9437
rect 30604 9260 30644 9388
rect 30593 9220 30644 9260
rect 30593 9101 30633 9220
rect 30593 9092 30645 9101
rect 30593 9052 30604 9092
rect 30644 9052 30645 9092
rect 30603 9043 30645 9052
rect 30603 8924 30645 8933
rect 30603 8884 30604 8924
rect 30644 8884 30645 8924
rect 30603 8875 30645 8884
rect 30604 8686 30644 8875
rect 30604 8637 30644 8646
rect 30796 8597 30836 9472
rect 30891 9472 30892 9512
rect 30932 9472 30933 9512
rect 30891 9463 30933 9472
rect 30988 9472 30998 9512
rect 31038 9472 31039 9512
rect 30988 9463 31039 9472
rect 30988 9428 31028 9463
rect 30988 9379 31028 9388
rect 31084 9260 31124 9640
rect 31467 9631 31509 9640
rect 31179 9512 31221 9521
rect 31179 9472 31180 9512
rect 31220 9472 31221 9512
rect 31179 9463 31221 9472
rect 31180 9269 31220 9463
rect 30892 9220 31124 9260
rect 31179 9260 31221 9269
rect 31179 9220 31180 9260
rect 31220 9220 31221 9260
rect 30795 8588 30837 8597
rect 30795 8548 30796 8588
rect 30836 8548 30837 8588
rect 30795 8539 30837 8548
rect 30796 8462 30836 8471
rect 30796 7925 30836 8422
rect 30795 7916 30837 7925
rect 30795 7876 30796 7916
rect 30836 7876 30837 7916
rect 30795 7867 30837 7876
rect 30892 7748 30932 9220
rect 31179 9211 31221 9220
rect 31083 8924 31125 8933
rect 31083 8884 31084 8924
rect 31124 8884 31125 8924
rect 31083 8875 31125 8884
rect 30987 8504 31029 8513
rect 30987 8464 30988 8504
rect 31028 8464 31029 8504
rect 30987 8455 31029 8464
rect 30988 8370 31028 8455
rect 30987 8168 31029 8177
rect 30987 8128 30988 8168
rect 31028 8128 31029 8168
rect 31084 8168 31124 8875
rect 31180 8756 31220 8765
rect 31220 8716 31316 8756
rect 31180 8707 31220 8716
rect 31180 8168 31220 8177
rect 31084 8128 31180 8168
rect 30987 8119 31029 8128
rect 31180 8119 31220 8128
rect 30796 7708 30932 7748
rect 30988 8000 31028 8119
rect 30316 5776 30548 5816
rect 30700 6474 30740 6483
rect 30219 5564 30261 5573
rect 30219 5524 30220 5564
rect 30260 5524 30261 5564
rect 30219 5515 30261 5524
rect 30220 4976 30260 5515
rect 30027 4640 30069 4649
rect 30027 4600 30028 4640
rect 30068 4600 30069 4640
rect 30027 4591 30069 4600
rect 30124 4136 30164 4145
rect 29931 3464 29973 3473
rect 29931 3424 29932 3464
rect 29972 3424 29973 3464
rect 29931 3415 29973 3424
rect 29644 1324 29876 1364
rect 29644 1280 29684 1324
rect 29644 1231 29684 1240
rect 29452 1147 29492 1156
rect 28876 1063 28916 1072
rect 29932 1112 29972 3415
rect 30124 1289 30164 4096
rect 30220 3473 30260 4936
rect 30316 3809 30356 5776
rect 30460 5657 30500 5666
rect 30500 5617 30548 5648
rect 30460 5608 30548 5617
rect 30315 3800 30357 3809
rect 30315 3760 30316 3800
rect 30356 3760 30357 3800
rect 30315 3751 30357 3760
rect 30219 3464 30261 3473
rect 30219 3424 30220 3464
rect 30260 3424 30261 3464
rect 30219 3415 30261 3424
rect 30508 3305 30548 5608
rect 30603 5564 30645 5573
rect 30603 5524 30604 5564
rect 30644 5524 30645 5564
rect 30603 5515 30645 5524
rect 30604 5430 30644 5515
rect 30700 5060 30740 6434
rect 30796 6329 30836 7708
rect 30891 7496 30933 7505
rect 30891 7456 30892 7496
rect 30932 7456 30933 7496
rect 30891 7447 30933 7456
rect 30892 6656 30932 7447
rect 30988 7169 31028 7960
rect 30987 7160 31029 7169
rect 30987 7120 30988 7160
rect 31028 7120 31029 7160
rect 30987 7111 31029 7120
rect 30892 6607 30932 6616
rect 31276 6404 31316 8716
rect 31371 8504 31413 8513
rect 31371 8464 31372 8504
rect 31412 8464 31413 8504
rect 31371 8455 31413 8464
rect 31372 8370 31412 8455
rect 31371 7748 31413 7757
rect 31371 7708 31372 7748
rect 31412 7708 31413 7748
rect 31371 7699 31413 7708
rect 31372 7614 31412 7699
rect 31468 7328 31508 9631
rect 31564 9101 31604 10219
rect 31563 9092 31605 9101
rect 31563 9052 31564 9092
rect 31604 9052 31605 9092
rect 31563 9043 31605 9052
rect 31564 8756 31604 8765
rect 31564 8177 31604 8716
rect 31563 8168 31605 8177
rect 31563 8128 31564 8168
rect 31604 8128 31605 8168
rect 31563 8119 31605 8128
rect 31563 7916 31605 7925
rect 31563 7876 31564 7916
rect 31604 7876 31605 7916
rect 31563 7867 31605 7876
rect 31564 7782 31604 7867
rect 30892 6364 31316 6404
rect 31372 7288 31508 7328
rect 30795 6320 30837 6329
rect 30795 6280 30796 6320
rect 30836 6280 30837 6320
rect 30795 6271 30837 6280
rect 30604 5020 30740 5060
rect 30892 5060 30932 6364
rect 30987 6068 31029 6077
rect 30987 6028 30988 6068
rect 31028 6028 31029 6068
rect 30987 6019 31029 6028
rect 30604 4304 30644 5020
rect 30892 5011 30932 5020
rect 30700 4962 30740 4971
rect 30700 4388 30740 4922
rect 30891 4892 30933 4901
rect 30891 4852 30892 4892
rect 30932 4852 30933 4892
rect 30891 4843 30933 4852
rect 30892 4649 30932 4843
rect 30891 4640 30933 4649
rect 30891 4600 30892 4640
rect 30932 4600 30933 4640
rect 30891 4591 30933 4600
rect 30700 4348 30836 4388
rect 30604 4264 30740 4304
rect 30603 4136 30645 4145
rect 30603 4096 30604 4136
rect 30644 4096 30645 4136
rect 30603 4087 30645 4096
rect 30604 4002 30644 4087
rect 30603 3632 30645 3641
rect 30603 3592 30604 3632
rect 30644 3592 30645 3632
rect 30603 3583 30645 3592
rect 30604 3464 30644 3583
rect 30700 3464 30740 4264
rect 30796 3632 30836 4348
rect 30892 4145 30932 4591
rect 30891 4136 30933 4145
rect 30891 4096 30892 4136
rect 30932 4096 30933 4136
rect 30891 4087 30933 4096
rect 30988 3977 31028 6019
rect 30987 3968 31029 3977
rect 30987 3928 30988 3968
rect 31028 3928 31029 3968
rect 30987 3919 31029 3928
rect 31372 3716 31412 7288
rect 31660 7253 31700 10480
rect 31851 10471 31893 10480
rect 31755 8504 31797 8513
rect 31755 8464 31756 8504
rect 31796 8464 31797 8504
rect 31755 8455 31797 8464
rect 31756 8370 31796 8455
rect 31755 8168 31797 8177
rect 31755 8128 31756 8168
rect 31796 8128 31797 8168
rect 31755 8119 31797 8128
rect 31659 7244 31701 7253
rect 31659 7204 31660 7244
rect 31700 7204 31701 7244
rect 31659 7195 31701 7204
rect 31468 7160 31508 7169
rect 31563 7160 31605 7169
rect 31508 7120 31564 7160
rect 31604 7120 31605 7160
rect 31468 7111 31508 7120
rect 31563 7111 31605 7120
rect 31660 6992 31700 7001
rect 31468 6952 31660 6992
rect 31468 6488 31508 6952
rect 31660 6943 31700 6952
rect 31563 6824 31605 6833
rect 31563 6784 31564 6824
rect 31604 6784 31605 6824
rect 31563 6775 31605 6784
rect 31468 6439 31508 6448
rect 31564 6488 31604 6775
rect 31604 6448 31700 6488
rect 31564 6439 31604 6448
rect 31467 6320 31509 6329
rect 31467 6280 31468 6320
rect 31508 6280 31509 6320
rect 31467 6271 31509 6280
rect 30796 3583 30836 3592
rect 31276 3676 31412 3716
rect 30700 3424 31124 3464
rect 30507 3296 30549 3305
rect 30507 3256 30508 3296
rect 30548 3256 30549 3296
rect 30507 3247 30549 3256
rect 30604 2540 30644 3424
rect 30987 3296 31029 3305
rect 30987 3256 30988 3296
rect 31028 3256 31029 3296
rect 30987 3247 31029 3256
rect 30892 2624 30932 2633
rect 30796 2584 30892 2624
rect 30796 2540 30836 2584
rect 30892 2575 30932 2584
rect 30604 2500 30836 2540
rect 30796 1952 30836 2500
rect 30988 2120 31028 3247
rect 31084 2876 31124 3424
rect 31180 3296 31220 3305
rect 31276 3296 31316 3676
rect 31220 3256 31316 3296
rect 31372 3380 31412 3389
rect 31180 3247 31220 3256
rect 31372 2885 31412 3340
rect 31084 2827 31124 2836
rect 31371 2876 31413 2885
rect 31371 2836 31372 2876
rect 31412 2836 31413 2876
rect 31371 2827 31413 2836
rect 31468 2708 31508 6271
rect 31660 5993 31700 6448
rect 31659 5984 31701 5993
rect 31659 5944 31660 5984
rect 31700 5944 31701 5984
rect 31659 5935 31701 5944
rect 31564 5648 31604 5657
rect 31564 4397 31604 5608
rect 31660 5648 31700 5935
rect 31660 5599 31700 5608
rect 31756 5573 31796 8119
rect 31852 5648 31892 10471
rect 31948 8924 31988 10672
rect 31948 8884 32084 8924
rect 31948 8756 31988 8765
rect 31948 7505 31988 8716
rect 31947 7496 31989 7505
rect 31947 7456 31948 7496
rect 31988 7456 31989 7496
rect 31947 7447 31989 7456
rect 31947 7328 31989 7337
rect 31947 7288 31948 7328
rect 31988 7288 31989 7328
rect 31947 7279 31989 7288
rect 31948 7160 31988 7279
rect 31948 7111 31988 7120
rect 32044 6656 32084 8884
rect 32140 6824 32180 10672
rect 32235 10352 32277 10361
rect 32235 10312 32236 10352
rect 32276 10312 32277 10352
rect 32235 10303 32277 10312
rect 32236 8168 32276 10303
rect 32332 9773 32372 10672
rect 32331 9764 32373 9773
rect 32331 9724 32332 9764
rect 32372 9724 32373 9764
rect 32331 9715 32373 9724
rect 32427 9680 32469 9689
rect 32427 9640 32428 9680
rect 32468 9640 32469 9680
rect 32427 9631 32469 9640
rect 32428 9512 32468 9631
rect 32428 9463 32468 9472
rect 32427 9260 32469 9269
rect 32332 9220 32428 9260
rect 32468 9220 32469 9260
rect 32332 8672 32372 9220
rect 32427 9211 32469 9220
rect 32427 9092 32469 9101
rect 32427 9052 32428 9092
rect 32468 9052 32469 9092
rect 32427 9043 32469 9052
rect 32332 8623 32372 8632
rect 32428 8672 32468 9043
rect 32524 9008 32564 10672
rect 32631 10648 32756 10672
rect 32631 10604 32671 10648
rect 32620 10564 32671 10604
rect 32620 9605 32660 10564
rect 32811 10184 32853 10193
rect 32811 10144 32812 10184
rect 32852 10144 32853 10184
rect 32811 10135 32853 10144
rect 32715 9764 32757 9773
rect 32715 9724 32716 9764
rect 32756 9724 32757 9764
rect 32715 9715 32757 9724
rect 32619 9596 32661 9605
rect 32619 9556 32620 9596
rect 32660 9556 32661 9596
rect 32619 9547 32661 9556
rect 32619 9260 32661 9269
rect 32619 9220 32620 9260
rect 32660 9220 32661 9260
rect 32619 9211 32661 9220
rect 32620 9126 32660 9211
rect 32524 8968 32660 9008
rect 32428 8623 32468 8632
rect 32236 8119 32276 8128
rect 32620 8084 32660 8968
rect 32524 8044 32660 8084
rect 32428 7916 32468 7925
rect 32428 7673 32468 7876
rect 32427 7664 32469 7673
rect 32427 7624 32428 7664
rect 32468 7624 32469 7664
rect 32427 7615 32469 7624
rect 32524 7421 32564 8044
rect 32619 7748 32661 7757
rect 32619 7708 32620 7748
rect 32660 7708 32661 7748
rect 32619 7699 32661 7708
rect 32620 7614 32660 7699
rect 32523 7412 32565 7421
rect 32523 7372 32524 7412
rect 32564 7372 32565 7412
rect 32523 7363 32565 7372
rect 32140 6784 32468 6824
rect 32044 6616 32276 6656
rect 31947 6488 31989 6497
rect 31947 6448 31948 6488
rect 31988 6448 31989 6488
rect 31947 6439 31989 6448
rect 31948 5732 31988 6439
rect 32043 6404 32085 6413
rect 32043 6364 32044 6404
rect 32084 6364 32180 6404
rect 32043 6355 32085 6364
rect 32044 6270 32084 6355
rect 32044 5732 32084 5741
rect 31948 5692 32044 5732
rect 32044 5683 32084 5692
rect 32140 5732 32180 6364
rect 32140 5683 32180 5692
rect 31852 5608 31988 5648
rect 31755 5564 31797 5573
rect 31755 5524 31756 5564
rect 31796 5524 31797 5564
rect 31755 5515 31797 5524
rect 31659 5480 31701 5489
rect 31659 5440 31660 5480
rect 31700 5440 31701 5480
rect 31659 5431 31701 5440
rect 31563 4388 31605 4397
rect 31563 4348 31564 4388
rect 31604 4348 31605 4388
rect 31563 4339 31605 4348
rect 31563 3800 31605 3809
rect 31563 3760 31564 3800
rect 31604 3760 31605 3800
rect 31563 3751 31605 3760
rect 31564 3632 31604 3751
rect 31564 3583 31604 3592
rect 31382 2668 31508 2708
rect 31382 2540 31422 2668
rect 31660 2624 31700 5431
rect 31851 4556 31893 4565
rect 31851 4516 31852 4556
rect 31892 4516 31893 4556
rect 31851 4507 31893 4516
rect 31852 4136 31892 4507
rect 31852 4087 31892 4096
rect 31851 3968 31893 3977
rect 31851 3928 31852 3968
rect 31892 3928 31893 3968
rect 31851 3919 31893 3928
rect 31756 3380 31796 3389
rect 31756 2633 31796 3340
rect 31372 2500 31422 2540
rect 31468 2584 31700 2624
rect 31755 2624 31797 2633
rect 31755 2584 31756 2624
rect 31796 2584 31797 2624
rect 31468 2582 31508 2584
rect 31755 2575 31797 2584
rect 31468 2533 31508 2542
rect 30988 2071 31028 2080
rect 31179 2120 31221 2129
rect 31179 2080 31180 2120
rect 31220 2080 31221 2120
rect 31179 2071 31221 2080
rect 31180 1986 31220 2071
rect 31372 2036 31412 2500
rect 31852 2372 31892 3919
rect 31948 3809 31988 5608
rect 32139 5564 32181 5573
rect 32139 5524 32140 5564
rect 32180 5524 32181 5564
rect 32139 5515 32181 5524
rect 32044 4985 32084 5070
rect 32043 4976 32085 4985
rect 32043 4936 32044 4976
rect 32084 4936 32085 4976
rect 32043 4927 32085 4936
rect 32043 4388 32085 4397
rect 32043 4348 32044 4388
rect 32084 4348 32085 4388
rect 32043 4339 32085 4348
rect 32044 4254 32084 4339
rect 31947 3800 31989 3809
rect 31947 3760 31948 3800
rect 31988 3760 31989 3800
rect 31947 3751 31989 3760
rect 31564 2332 31892 2372
rect 31564 2120 31604 2332
rect 31564 2071 31604 2080
rect 31372 1996 31508 2036
rect 30796 1625 30836 1912
rect 30891 1952 30933 1961
rect 30891 1912 30892 1952
rect 30932 1912 30933 1952
rect 30891 1903 30933 1912
rect 30795 1616 30837 1625
rect 30795 1576 30796 1616
rect 30836 1576 30837 1616
rect 30795 1567 30837 1576
rect 30123 1280 30165 1289
rect 30123 1240 30124 1280
rect 30164 1240 30165 1280
rect 30123 1231 30165 1240
rect 29932 1063 29972 1072
rect 30892 1112 30932 1903
rect 31372 1868 31412 1877
rect 31372 1709 31412 1828
rect 31371 1700 31413 1709
rect 31371 1660 31372 1700
rect 31412 1660 31413 1700
rect 31371 1651 31413 1660
rect 30892 1063 30932 1072
rect 31179 1112 31221 1121
rect 31179 1072 31180 1112
rect 31220 1072 31221 1112
rect 31179 1063 31221 1072
rect 31180 978 31220 1063
rect 31468 953 31508 1996
rect 31756 1868 31796 1877
rect 31564 1828 31756 1868
rect 28587 944 28629 953
rect 28587 904 28588 944
rect 28628 904 28629 944
rect 28587 895 28629 904
rect 31467 944 31509 953
rect 31467 904 31468 944
rect 31508 904 31509 944
rect 31467 895 31509 904
rect 29451 776 29493 785
rect 29451 736 29452 776
rect 29492 736 29493 776
rect 29451 727 29493 736
rect 29452 80 29492 727
rect 30603 608 30645 617
rect 30603 568 30604 608
rect 30644 568 30645 608
rect 30603 559 30645 568
rect 30604 80 30644 559
rect 31564 533 31604 1828
rect 31756 1819 31796 1828
rect 31659 1280 31701 1289
rect 31659 1240 31660 1280
rect 31700 1240 31701 1280
rect 31659 1231 31701 1240
rect 31660 1146 31700 1231
rect 31755 1196 31797 1205
rect 31755 1156 31756 1196
rect 31796 1156 31797 1196
rect 31755 1147 31797 1156
rect 31563 524 31605 533
rect 31563 484 31564 524
rect 31604 484 31605 524
rect 31563 475 31605 484
rect 31756 80 31796 1147
rect 32140 869 32180 5515
rect 32236 5480 32276 6616
rect 32236 5440 32372 5480
rect 32235 4976 32277 4985
rect 32235 4936 32236 4976
rect 32276 4936 32277 4976
rect 32235 4927 32277 4936
rect 32236 4733 32276 4927
rect 32235 4724 32277 4733
rect 32235 4684 32236 4724
rect 32276 4684 32277 4724
rect 32235 4675 32277 4684
rect 32236 4481 32276 4675
rect 32235 4472 32277 4481
rect 32235 4432 32236 4472
rect 32276 4432 32277 4472
rect 32235 4423 32277 4432
rect 32235 3464 32277 3473
rect 32235 3424 32236 3464
rect 32276 3424 32277 3464
rect 32235 3415 32277 3424
rect 32236 2120 32276 3415
rect 32236 2071 32276 2080
rect 32332 1289 32372 5440
rect 32428 2372 32468 6784
rect 32524 6488 32564 6497
rect 32564 6448 32660 6488
rect 32524 6439 32564 6448
rect 32620 5648 32660 6448
rect 32620 5069 32660 5608
rect 32716 5573 32756 9715
rect 32812 8756 32852 10135
rect 32908 9680 32948 10672
rect 32908 9640 33044 9680
rect 32908 9512 32948 9523
rect 32908 9437 32948 9472
rect 32907 9428 32949 9437
rect 32907 9388 32908 9428
rect 32948 9388 32949 9428
rect 32907 9379 32949 9388
rect 32908 9269 32948 9379
rect 32907 9260 32949 9269
rect 32907 9220 32908 9260
rect 32948 9220 32949 9260
rect 32907 9211 32949 9220
rect 32812 8177 32852 8716
rect 32908 8672 32948 8683
rect 32908 8597 32948 8632
rect 32907 8588 32949 8597
rect 32907 8548 32908 8588
rect 32948 8548 32949 8588
rect 32907 8539 32949 8548
rect 32908 8261 32948 8539
rect 33004 8429 33044 9640
rect 33100 8765 33140 10672
rect 33292 8924 33332 10672
rect 33484 9437 33524 10672
rect 41451 10520 41493 10529
rect 41451 10480 41452 10520
rect 41492 10480 41493 10520
rect 41451 10471 41493 10480
rect 34731 10436 34773 10445
rect 34731 10396 34732 10436
rect 34772 10396 34773 10436
rect 34731 10387 34773 10396
rect 34155 9680 34197 9689
rect 34155 9640 34156 9680
rect 34196 9640 34197 9680
rect 34155 9631 34197 9640
rect 34156 9512 34196 9631
rect 33483 9428 33525 9437
rect 33483 9388 33484 9428
rect 33524 9388 33525 9428
rect 34156 9428 34196 9472
rect 34156 9388 34580 9428
rect 33483 9379 33525 9388
rect 34348 9260 34388 9269
rect 34388 9220 34484 9260
rect 34348 9211 34388 9220
rect 33928 9092 34296 9101
rect 33968 9052 34010 9092
rect 34050 9052 34092 9092
rect 34132 9052 34174 9092
rect 34214 9052 34256 9092
rect 33928 9043 34296 9052
rect 33292 8884 33812 8924
rect 33099 8756 33141 8765
rect 33099 8716 33100 8756
rect 33140 8716 33141 8756
rect 33099 8707 33141 8716
rect 33388 8672 33428 8681
rect 33196 8632 33388 8672
rect 33428 8632 33524 8672
rect 33003 8420 33045 8429
rect 33003 8380 33004 8420
rect 33044 8380 33045 8420
rect 33003 8371 33045 8380
rect 33099 8336 33141 8345
rect 33196 8336 33236 8632
rect 33388 8623 33428 8632
rect 33099 8296 33100 8336
rect 33140 8296 33236 8336
rect 33099 8287 33141 8296
rect 33484 8261 33524 8632
rect 32907 8252 32949 8261
rect 32907 8212 32908 8252
rect 32948 8212 32949 8252
rect 32907 8203 32949 8212
rect 33483 8252 33525 8261
rect 33483 8212 33484 8252
rect 33524 8212 33525 8252
rect 33483 8203 33525 8212
rect 32811 8168 32853 8177
rect 32811 8128 32812 8168
rect 32852 8128 32853 8168
rect 32811 8119 32853 8128
rect 33772 8084 33812 8884
rect 34347 8840 34389 8849
rect 34347 8800 34348 8840
rect 34388 8800 34389 8840
rect 34347 8791 34389 8800
rect 33867 8756 33909 8765
rect 33867 8716 33868 8756
rect 33908 8716 33909 8756
rect 33867 8707 33909 8716
rect 33868 8686 33908 8707
rect 34348 8706 34388 8791
rect 34444 8765 34484 9220
rect 34443 8756 34485 8765
rect 34443 8716 34444 8756
rect 34484 8716 34485 8756
rect 34443 8707 34485 8716
rect 33868 8621 33908 8646
rect 33676 8044 33812 8084
rect 34060 8504 34100 8513
rect 33291 8000 33333 8009
rect 33291 7960 33292 8000
rect 33332 7960 33333 8000
rect 33291 7951 33333 7960
rect 32812 7916 32852 7925
rect 32852 7876 33140 7916
rect 32812 7867 32852 7876
rect 32907 7664 32949 7673
rect 32907 7624 32908 7664
rect 32948 7624 32949 7664
rect 32907 7615 32949 7624
rect 32811 7244 32853 7253
rect 32811 7204 32812 7244
rect 32852 7204 32853 7244
rect 32811 7195 32853 7204
rect 32715 5564 32757 5573
rect 32715 5524 32716 5564
rect 32756 5524 32757 5564
rect 32715 5515 32757 5524
rect 32812 5396 32852 7195
rect 32908 5480 32948 7615
rect 33003 7160 33045 7169
rect 33003 7120 33004 7160
rect 33044 7120 33045 7160
rect 33003 7111 33045 7120
rect 33004 6665 33044 7111
rect 33003 6656 33045 6665
rect 33003 6616 33004 6656
rect 33044 6616 33045 6656
rect 33100 6656 33140 7876
rect 33292 7757 33332 7951
rect 33291 7748 33333 7757
rect 33291 7708 33292 7748
rect 33332 7708 33333 7748
rect 33291 7699 33333 7708
rect 33195 7160 33237 7169
rect 33195 7120 33196 7160
rect 33236 7120 33237 7160
rect 33676 7160 33716 8044
rect 34060 7748 34100 8464
rect 34540 8000 34580 9388
rect 34732 8849 34772 10387
rect 35168 9848 35536 9857
rect 35208 9808 35250 9848
rect 35290 9808 35332 9848
rect 35372 9808 35414 9848
rect 35454 9808 35496 9848
rect 35168 9799 35536 9808
rect 40299 9848 40341 9857
rect 40299 9808 40300 9848
rect 40340 9808 40341 9848
rect 40299 9799 40341 9808
rect 37131 9596 37173 9605
rect 37131 9556 37132 9596
rect 37172 9556 37173 9596
rect 37131 9547 37173 9556
rect 35020 9512 35060 9521
rect 35020 9269 35060 9472
rect 36268 9512 36308 9521
rect 35019 9260 35061 9269
rect 35019 9220 35020 9260
rect 35060 9220 35061 9260
rect 35019 9211 35061 9220
rect 36268 9101 36308 9472
rect 36460 9260 36500 9269
rect 36075 9092 36117 9101
rect 36075 9052 36076 9092
rect 36116 9052 36117 9092
rect 36075 9043 36117 9052
rect 36267 9092 36309 9101
rect 36267 9052 36268 9092
rect 36308 9052 36309 9092
rect 36267 9043 36309 9052
rect 34731 8840 34773 8849
rect 34731 8800 34732 8840
rect 34772 8800 34773 8840
rect 34731 8791 34773 8800
rect 35787 8840 35829 8849
rect 35787 8800 35788 8840
rect 35828 8800 35829 8840
rect 35787 8791 35829 8800
rect 34635 8672 34677 8681
rect 34635 8632 34636 8672
rect 34676 8632 34677 8672
rect 34635 8623 34677 8632
rect 34732 8672 34772 8791
rect 35595 8756 35637 8765
rect 35595 8716 35596 8756
rect 35636 8716 35637 8756
rect 35595 8707 35637 8716
rect 35020 8672 35060 8681
rect 34732 8623 34772 8632
rect 34828 8632 35020 8672
rect 34636 8538 34676 8623
rect 34732 8168 34772 8177
rect 34828 8168 34868 8632
rect 35020 8623 35060 8632
rect 35168 8336 35536 8345
rect 35208 8296 35250 8336
rect 35290 8296 35332 8336
rect 35372 8296 35414 8336
rect 35454 8296 35496 8336
rect 35168 8287 35536 8296
rect 34772 8128 34868 8168
rect 34732 8119 34772 8128
rect 34580 7960 34676 8000
rect 34540 7951 34580 7960
rect 33772 7708 34100 7748
rect 33772 7244 33812 7708
rect 33928 7580 34296 7589
rect 33968 7540 34010 7580
rect 34050 7540 34092 7580
rect 34132 7540 34174 7580
rect 34214 7540 34256 7580
rect 33928 7531 34296 7540
rect 33868 7244 33908 7253
rect 33772 7204 33868 7244
rect 33868 7195 33908 7204
rect 34540 7160 34580 7169
rect 33676 7120 33812 7160
rect 33195 7111 33237 7120
rect 33196 7026 33236 7111
rect 33388 6992 33428 7001
rect 33292 6952 33388 6992
rect 33196 6656 33236 6665
rect 33100 6616 33196 6656
rect 33003 6607 33045 6616
rect 33196 6607 33236 6616
rect 33052 6446 33092 6455
rect 33052 6404 33092 6406
rect 33292 6404 33332 6952
rect 33388 6943 33428 6952
rect 33675 6992 33717 7001
rect 33675 6952 33676 6992
rect 33716 6952 33717 6992
rect 33675 6943 33717 6952
rect 33676 6858 33716 6943
rect 33675 6656 33717 6665
rect 33675 6616 33676 6656
rect 33716 6616 33717 6656
rect 33675 6607 33717 6616
rect 33388 6497 33428 6582
rect 33387 6488 33429 6497
rect 33387 6448 33388 6488
rect 33428 6448 33429 6488
rect 33387 6439 33429 6448
rect 33052 6364 33332 6404
rect 33388 5692 33524 5732
rect 33148 5657 33188 5666
rect 33388 5657 33428 5692
rect 33188 5617 33428 5657
rect 33148 5608 33188 5617
rect 33292 5480 33332 5489
rect 32908 5440 33292 5480
rect 33292 5431 33332 5440
rect 32812 5356 33044 5396
rect 32619 5060 32661 5069
rect 32619 5020 32620 5060
rect 32660 5020 32661 5060
rect 32619 5011 32661 5020
rect 32524 4145 32564 4230
rect 32523 4136 32565 4145
rect 32523 4096 32524 4136
rect 32564 4096 32565 4136
rect 32523 4087 32565 4096
rect 32523 3800 32565 3809
rect 32523 3760 32524 3800
rect 32564 3760 32565 3800
rect 32523 3751 32565 3760
rect 32524 2456 32564 3751
rect 32811 3632 32853 3641
rect 32811 3592 32812 3632
rect 32852 3592 32853 3632
rect 32811 3583 32853 3592
rect 32715 3548 32757 3557
rect 32715 3508 32716 3548
rect 32756 3508 32757 3548
rect 32715 3499 32757 3508
rect 32620 3464 32660 3473
rect 32620 2885 32660 3424
rect 32716 3464 32756 3499
rect 32716 3413 32756 3424
rect 32619 2876 32661 2885
rect 32619 2836 32620 2876
rect 32660 2836 32661 2876
rect 32619 2827 32661 2836
rect 32716 2624 32756 2633
rect 32812 2624 32852 3583
rect 32907 2876 32949 2885
rect 32907 2836 32908 2876
rect 32948 2836 32949 2876
rect 32907 2827 32949 2836
rect 32908 2742 32948 2827
rect 32756 2584 32852 2624
rect 32716 2575 32756 2584
rect 32524 2416 32756 2456
rect 32428 2332 32660 2372
rect 32331 1280 32373 1289
rect 32331 1240 32332 1280
rect 32372 1240 32373 1280
rect 32331 1231 32373 1240
rect 32524 1196 32564 1205
rect 32331 944 32373 953
rect 32331 904 32332 944
rect 32372 904 32373 944
rect 32331 895 32373 904
rect 32139 860 32181 869
rect 32139 820 32140 860
rect 32180 820 32181 860
rect 32139 811 32181 820
rect 32332 810 32372 895
rect 32524 701 32564 1156
rect 32620 869 32660 2332
rect 32716 1280 32756 2416
rect 33004 1280 33044 5356
rect 33099 5312 33141 5321
rect 33099 5272 33100 5312
rect 33140 5272 33141 5312
rect 33099 5263 33141 5272
rect 33100 3725 33140 5263
rect 33484 5144 33524 5692
rect 33484 5095 33524 5104
rect 33292 4976 33332 4985
rect 33195 4808 33237 4817
rect 33195 4768 33196 4808
rect 33236 4768 33237 4808
rect 33195 4759 33237 4768
rect 33196 4145 33236 4759
rect 33292 4565 33332 4936
rect 33291 4556 33333 4565
rect 33291 4516 33292 4556
rect 33332 4516 33333 4556
rect 33291 4507 33333 4516
rect 33195 4136 33237 4145
rect 33195 4096 33196 4136
rect 33236 4096 33237 4136
rect 33195 4087 33237 4096
rect 33099 3716 33141 3725
rect 33099 3676 33100 3716
rect 33140 3676 33141 3716
rect 33099 3667 33141 3676
rect 33100 3464 33140 3667
rect 33100 3415 33140 3424
rect 33196 3464 33236 4087
rect 33196 3415 33236 3424
rect 33292 2633 33332 4507
rect 33676 4136 33716 6607
rect 33772 5153 33812 7120
rect 34444 7120 34540 7160
rect 34444 6497 34484 7120
rect 34540 7111 34580 7120
rect 34539 6908 34581 6917
rect 34539 6868 34540 6908
rect 34580 6868 34581 6908
rect 34539 6859 34581 6868
rect 34443 6488 34485 6497
rect 34443 6448 34444 6488
rect 34484 6448 34485 6488
rect 34443 6439 34485 6448
rect 34347 6236 34389 6245
rect 34347 6196 34348 6236
rect 34388 6196 34389 6236
rect 34347 6187 34389 6196
rect 33928 6068 34296 6077
rect 33968 6028 34010 6068
rect 34050 6028 34092 6068
rect 34132 6028 34174 6068
rect 34214 6028 34256 6068
rect 33928 6019 34296 6028
rect 34348 5648 34388 6187
rect 34443 5816 34485 5825
rect 34443 5776 34444 5816
rect 34484 5776 34485 5816
rect 34443 5767 34485 5776
rect 34348 5599 34388 5608
rect 34444 5648 34484 5767
rect 34444 5599 34484 5608
rect 33771 5144 33813 5153
rect 33771 5104 33772 5144
rect 33812 5104 33813 5144
rect 33771 5095 33813 5104
rect 34348 4976 34388 4985
rect 34540 4976 34580 6859
rect 34636 6497 34676 7960
rect 35168 6824 35536 6833
rect 35208 6784 35250 6824
rect 35290 6784 35332 6824
rect 35372 6784 35414 6824
rect 35454 6784 35496 6824
rect 35168 6775 35536 6784
rect 35596 6656 35636 8707
rect 35692 8672 35732 8681
rect 35692 7412 35732 8632
rect 35788 8672 35828 8791
rect 35788 8623 35828 8632
rect 35980 7412 36020 7421
rect 35692 7372 35980 7412
rect 35980 7363 36020 7372
rect 36076 7169 36116 9043
rect 36363 8840 36405 8849
rect 36363 8800 36364 8840
rect 36404 8800 36405 8840
rect 36363 8791 36405 8800
rect 36267 8756 36309 8765
rect 36267 8716 36268 8756
rect 36308 8716 36309 8756
rect 36267 8707 36309 8716
rect 36172 8672 36212 8681
rect 36172 8513 36212 8632
rect 36268 8622 36308 8707
rect 36171 8504 36213 8513
rect 36171 8464 36172 8504
rect 36212 8464 36213 8504
rect 36171 8455 36213 8464
rect 36268 8000 36308 8009
rect 36268 7832 36308 7960
rect 36364 8000 36404 8791
rect 36364 7951 36404 7960
rect 36460 7832 36500 9220
rect 37036 9260 37076 9269
rect 37036 9017 37076 9220
rect 37035 9008 37077 9017
rect 37035 8968 37036 9008
rect 37076 8968 37077 9008
rect 37035 8959 37077 8968
rect 36748 8672 36788 8681
rect 36652 8632 36748 8672
rect 36268 7792 36500 7832
rect 36555 7832 36597 7841
rect 36652 7832 36692 8632
rect 36748 8623 36788 8632
rect 36555 7792 36556 7832
rect 36596 7792 36692 7832
rect 36748 7916 36788 7925
rect 36555 7783 36597 7792
rect 36556 7673 36596 7783
rect 36555 7664 36597 7673
rect 36555 7624 36556 7664
rect 36596 7624 36597 7664
rect 36555 7615 36597 7624
rect 35788 7160 35828 7169
rect 36075 7160 36117 7169
rect 35828 7120 36076 7160
rect 36116 7120 36117 7160
rect 35788 7111 35828 7120
rect 36075 7111 36117 7120
rect 36268 7160 36308 7169
rect 36076 7026 36116 7111
rect 36268 6917 36308 7120
rect 36267 6908 36309 6917
rect 36267 6868 36268 6908
rect 36308 6868 36309 6908
rect 36267 6859 36309 6868
rect 35404 6616 35636 6656
rect 34635 6488 34677 6497
rect 34635 6448 34636 6488
rect 34676 6448 34677 6488
rect 34635 6439 34677 6448
rect 34636 6354 34676 6439
rect 34828 6245 34868 6330
rect 34827 6236 34869 6245
rect 34827 6196 34828 6236
rect 34868 6196 34869 6236
rect 34827 6187 34869 6196
rect 34827 5984 34869 5993
rect 34827 5944 34828 5984
rect 34868 5944 34869 5984
rect 34827 5935 34869 5944
rect 34828 5732 34868 5935
rect 35404 5825 35444 6616
rect 35595 6488 35637 6497
rect 35595 6448 35596 6488
rect 35636 6448 35637 6488
rect 35595 6439 35637 6448
rect 35403 5816 35445 5825
rect 35403 5776 35404 5816
rect 35444 5776 35445 5816
rect 35403 5767 35445 5776
rect 34828 5683 34868 5692
rect 34923 5648 34965 5657
rect 34923 5608 34924 5648
rect 34964 5608 34965 5648
rect 34923 5599 34965 5608
rect 35404 5648 35444 5767
rect 35404 5599 35444 5608
rect 34924 5514 34964 5599
rect 35168 5312 35536 5321
rect 35208 5272 35250 5312
rect 35290 5272 35332 5312
rect 35372 5272 35414 5312
rect 35454 5272 35496 5312
rect 35168 5263 35536 5272
rect 34388 4936 34580 4976
rect 35596 4976 35636 6439
rect 35884 6404 35924 6413
rect 36555 6404 36597 6413
rect 35924 6364 36020 6404
rect 35884 6355 35924 6364
rect 35691 6320 35733 6329
rect 35691 6280 35692 6320
rect 35732 6280 35733 6320
rect 35691 6271 35733 6280
rect 35692 6186 35732 6271
rect 35884 5653 35924 5662
rect 35788 5144 35828 5153
rect 35884 5144 35924 5613
rect 35980 5564 36020 6364
rect 36555 6364 36556 6404
rect 36596 6364 36597 6404
rect 36555 6355 36597 6364
rect 36267 5984 36309 5993
rect 36267 5944 36268 5984
rect 36308 5944 36309 5984
rect 36267 5935 36309 5944
rect 36076 5564 36116 5573
rect 35980 5524 36076 5564
rect 36076 5515 36116 5524
rect 35828 5104 35924 5144
rect 35788 5095 35828 5104
rect 34348 4927 34388 4936
rect 35596 4927 35636 4936
rect 33928 4556 34296 4565
rect 33968 4516 34010 4556
rect 34050 4516 34092 4556
rect 34132 4516 34174 4556
rect 34214 4516 34256 4556
rect 33928 4507 34296 4516
rect 35404 4264 35636 4304
rect 34348 4220 34388 4229
rect 33772 4136 33812 4145
rect 33676 4096 33772 4136
rect 33772 3641 33812 4096
rect 33964 3968 34004 3977
rect 34155 3968 34197 3977
rect 34004 3928 34100 3968
rect 33964 3919 34004 3928
rect 34060 3716 34100 3928
rect 34155 3928 34156 3968
rect 34196 3928 34197 3968
rect 34155 3919 34197 3928
rect 34156 3834 34196 3919
rect 34060 3676 34196 3716
rect 33771 3632 33813 3641
rect 33771 3592 33772 3632
rect 33812 3592 33813 3632
rect 33771 3583 33813 3592
rect 33676 3473 33716 3558
rect 33675 3464 33717 3473
rect 33675 3424 33676 3464
rect 33716 3424 33717 3464
rect 33675 3415 33717 3424
rect 34156 3459 34196 3676
rect 34348 3632 34388 4180
rect 35404 4220 35444 4264
rect 35596 4220 35636 4264
rect 35596 4180 35732 4220
rect 35404 4171 35444 4180
rect 34348 3583 34388 3592
rect 34924 4136 34964 4145
rect 34156 3410 34196 3419
rect 33675 3296 33717 3305
rect 33675 3256 33676 3296
rect 33716 3256 33717 3296
rect 33675 3247 33717 3256
rect 33291 2624 33333 2633
rect 33291 2584 33292 2624
rect 33332 2584 33333 2624
rect 33291 2575 33333 2584
rect 33676 2624 33716 3247
rect 33928 3044 34296 3053
rect 33968 3004 34010 3044
rect 34050 3004 34092 3044
rect 34132 3004 34174 3044
rect 34214 3004 34256 3044
rect 33928 2995 34296 3004
rect 34924 2876 34964 4096
rect 35020 4136 35060 4145
rect 35020 3557 35060 4096
rect 35499 4136 35541 4145
rect 35499 4096 35500 4136
rect 35540 4096 35541 4136
rect 35499 4087 35541 4096
rect 35500 4002 35540 4087
rect 35595 3884 35637 3893
rect 35595 3844 35596 3884
rect 35636 3844 35637 3884
rect 35595 3835 35637 3844
rect 35168 3800 35536 3809
rect 35208 3760 35250 3800
rect 35290 3760 35332 3800
rect 35372 3760 35414 3800
rect 35454 3760 35496 3800
rect 35168 3751 35536 3760
rect 35596 3641 35636 3835
rect 35692 3716 35732 4180
rect 35883 4136 35925 4145
rect 35883 4096 35884 4136
rect 35924 4096 35925 4136
rect 35883 4087 35925 4096
rect 35980 4136 36020 4145
rect 35787 3716 35829 3725
rect 35692 3676 35788 3716
rect 35828 3676 35829 3716
rect 35787 3667 35829 3676
rect 35595 3632 35637 3641
rect 35595 3592 35596 3632
rect 35636 3592 35637 3632
rect 35595 3583 35637 3592
rect 35019 3548 35061 3557
rect 35019 3508 35020 3548
rect 35060 3508 35061 3548
rect 35019 3499 35061 3508
rect 35403 3548 35445 3557
rect 35403 3508 35404 3548
rect 35444 3508 35445 3548
rect 35403 3499 35445 3508
rect 35308 3464 35348 3473
rect 35116 2876 35156 2885
rect 34924 2836 35116 2876
rect 35116 2827 35156 2836
rect 34924 2633 34964 2718
rect 33676 2575 33716 2584
rect 34923 2624 34965 2633
rect 34923 2584 34924 2624
rect 34964 2584 34965 2624
rect 34923 2575 34965 2584
rect 34827 2456 34869 2465
rect 34827 2416 34828 2456
rect 34868 2416 34869 2456
rect 34827 2407 34869 2416
rect 34828 2120 34868 2407
rect 34828 2071 34868 2080
rect 34635 2036 34677 2045
rect 34635 1996 34636 2036
rect 34676 1996 34677 2036
rect 34635 1987 34677 1996
rect 33387 1952 33429 1961
rect 33387 1912 33388 1952
rect 33428 1912 33429 1952
rect 33387 1903 33429 1912
rect 34252 1952 34292 1961
rect 34292 1912 34388 1952
rect 34252 1903 34292 1912
rect 33388 1818 33428 1903
rect 33928 1532 34296 1541
rect 33968 1492 34010 1532
rect 34050 1492 34092 1532
rect 34132 1492 34174 1532
rect 34214 1492 34256 1532
rect 33928 1483 34296 1492
rect 34348 1364 34388 1912
rect 34636 1902 34676 1987
rect 34924 1952 34964 2575
rect 35308 2465 35348 3424
rect 35404 3464 35444 3499
rect 35404 3413 35444 3424
rect 35500 2624 35540 2633
rect 35596 2624 35636 3583
rect 35788 3464 35828 3667
rect 35788 3415 35828 3424
rect 35884 3464 35924 4087
rect 35980 3473 36020 4096
rect 35884 3415 35924 3424
rect 35979 3464 36021 3473
rect 35979 3424 35980 3464
rect 36020 3424 36021 3464
rect 36268 3464 36308 5935
rect 36556 5741 36596 6355
rect 36555 5732 36597 5741
rect 36555 5692 36556 5732
rect 36596 5692 36597 5732
rect 36555 5683 36597 5692
rect 36364 5648 36404 5657
rect 36364 4052 36404 5608
rect 36459 5648 36501 5657
rect 36459 5608 36460 5648
rect 36500 5608 36501 5648
rect 36459 5599 36501 5608
rect 36460 5514 36500 5599
rect 36748 5573 36788 7876
rect 36844 7916 36884 7925
rect 36844 5993 36884 7876
rect 36843 5984 36885 5993
rect 36843 5944 36844 5984
rect 36884 5944 36885 5984
rect 36843 5935 36885 5944
rect 36844 5732 36884 5935
rect 36844 5683 36884 5692
rect 36940 5648 36980 5659
rect 36940 5573 36980 5608
rect 36747 5564 36789 5573
rect 36747 5524 36748 5564
rect 36788 5524 36789 5564
rect 36747 5515 36789 5524
rect 36939 5564 36981 5573
rect 36939 5524 36940 5564
rect 36980 5524 36981 5564
rect 36939 5515 36981 5524
rect 37132 5480 37172 9547
rect 38476 9512 38516 9521
rect 37228 9428 37268 9437
rect 37804 9428 37844 9437
rect 37268 9388 37364 9428
rect 37228 9379 37268 9388
rect 37228 8677 37268 8686
rect 37228 7832 37268 8637
rect 37324 8588 37364 9388
rect 37844 9388 38036 9428
rect 37804 9379 37844 9388
rect 37611 9260 37653 9269
rect 37611 9220 37612 9260
rect 37652 9220 37653 9260
rect 37611 9211 37653 9220
rect 37612 9126 37652 9211
rect 37803 8924 37845 8933
rect 37803 8884 37804 8924
rect 37844 8884 37845 8924
rect 37803 8875 37845 8884
rect 37804 8672 37844 8875
rect 37804 8623 37844 8632
rect 37420 8588 37460 8597
rect 37324 8548 37420 8588
rect 37420 8539 37460 8548
rect 37612 8504 37652 8513
rect 37324 8009 37364 8094
rect 37612 8009 37652 8464
rect 37996 8168 38036 9388
rect 38284 9260 38324 9269
rect 37996 8119 38036 8128
rect 38092 9220 38284 9260
rect 37323 8000 37365 8009
rect 37323 7960 37324 8000
rect 37364 7960 37365 8000
rect 37323 7951 37365 7960
rect 37611 8000 37653 8009
rect 38092 8000 38132 9220
rect 38284 9211 38324 9220
rect 38476 8933 38516 9472
rect 39723 9512 39765 9521
rect 39723 9472 39724 9512
rect 39764 9472 39765 9512
rect 39723 9463 39765 9472
rect 39724 9378 39764 9463
rect 38859 9344 38901 9353
rect 38859 9304 38860 9344
rect 38900 9304 38901 9344
rect 38859 9295 38901 9304
rect 38475 8924 38517 8933
rect 38475 8884 38476 8924
rect 38516 8884 38517 8924
rect 38475 8875 38517 8884
rect 38667 8504 38709 8513
rect 38667 8464 38668 8504
rect 38708 8464 38709 8504
rect 38667 8455 38709 8464
rect 38571 8252 38613 8261
rect 38571 8212 38572 8252
rect 38612 8212 38613 8252
rect 38571 8203 38613 8212
rect 37611 7960 37612 8000
rect 37652 7960 37653 8000
rect 37611 7951 37653 7960
rect 37852 7990 38132 8000
rect 37892 7960 38132 7990
rect 38283 8000 38325 8009
rect 38283 7960 38284 8000
rect 38324 7960 38325 8000
rect 38283 7951 38325 7960
rect 38380 8000 38420 8009
rect 38420 7960 38516 8000
rect 38380 7951 38420 7960
rect 37852 7941 37892 7950
rect 38284 7866 38324 7951
rect 37228 7792 37748 7832
rect 37708 7412 37748 7792
rect 37708 7363 37748 7372
rect 37515 7160 37557 7169
rect 37515 7120 37516 7160
rect 37556 7120 37557 7160
rect 37515 7111 37557 7120
rect 37419 6068 37461 6077
rect 37419 6028 37420 6068
rect 37460 6028 37461 6068
rect 37419 6019 37461 6028
rect 37420 5825 37460 6019
rect 37419 5816 37461 5825
rect 37419 5776 37420 5816
rect 37460 5776 37461 5816
rect 37419 5767 37461 5776
rect 37420 5648 37460 5767
rect 37420 5599 37460 5608
rect 37132 5440 37460 5480
rect 37227 4976 37269 4985
rect 37227 4936 37228 4976
rect 37268 4936 37269 4976
rect 37227 4927 37269 4936
rect 36844 4892 36884 4901
rect 36884 4852 37172 4892
rect 36844 4843 36884 4852
rect 36651 4808 36693 4817
rect 36651 4768 36652 4808
rect 36692 4768 36693 4808
rect 36651 4759 36693 4768
rect 36652 4674 36692 4759
rect 37036 4220 37076 4229
rect 36508 4145 36548 4154
rect 37036 4136 37076 4180
rect 36548 4105 36596 4136
rect 36508 4096 36596 4105
rect 36364 4012 36500 4052
rect 36364 3464 36404 3473
rect 36268 3424 36364 3464
rect 35979 3415 36021 3424
rect 36364 3415 36404 3424
rect 35540 2584 35636 2624
rect 35500 2575 35540 2584
rect 35307 2456 35349 2465
rect 35307 2416 35308 2456
rect 35348 2416 35349 2456
rect 35307 2407 35349 2416
rect 35168 2288 35536 2297
rect 35208 2248 35250 2288
rect 35290 2248 35332 2288
rect 35372 2248 35414 2288
rect 35454 2248 35496 2288
rect 35168 2239 35536 2248
rect 36460 2120 36500 4012
rect 36556 2885 36596 4096
rect 36748 4096 37076 4136
rect 36652 4052 36692 4061
rect 36748 4052 36788 4096
rect 36692 4012 36788 4052
rect 36652 4003 36692 4012
rect 36843 3968 36885 3977
rect 36843 3928 36844 3968
rect 36884 3928 36885 3968
rect 36843 3919 36885 3928
rect 36844 3834 36884 3919
rect 36651 3800 36693 3809
rect 36651 3760 36652 3800
rect 36692 3760 36693 3800
rect 36651 3751 36693 3760
rect 36555 2876 36597 2885
rect 36555 2836 36556 2876
rect 36596 2836 36597 2876
rect 36555 2827 36597 2836
rect 36460 2071 36500 2080
rect 35020 1952 35060 1961
rect 34924 1912 35020 1952
rect 35020 1903 35060 1912
rect 36268 1952 36308 1961
rect 36268 1793 36308 1912
rect 36652 1952 36692 3751
rect 37036 3632 37076 3641
rect 37132 3632 37172 4852
rect 37228 4061 37268 4927
rect 37323 4136 37365 4145
rect 37323 4096 37324 4136
rect 37364 4096 37365 4136
rect 37323 4087 37365 4096
rect 37227 4052 37269 4061
rect 37227 4012 37228 4052
rect 37268 4012 37269 4052
rect 37227 4003 37269 4012
rect 37076 3592 37172 3632
rect 37324 3632 37364 4087
rect 37036 3583 37076 3592
rect 37324 3583 37364 3592
rect 36892 3422 36932 3431
rect 36892 3380 36932 3382
rect 36892 3340 37076 3380
rect 36939 2876 36981 2885
rect 36939 2836 36940 2876
rect 36980 2836 36981 2876
rect 36939 2827 36981 2836
rect 36940 2742 36980 2827
rect 36748 2633 36788 2719
rect 36747 2624 36789 2633
rect 36747 2584 36748 2624
rect 36788 2584 36789 2624
rect 36747 2575 36789 2584
rect 36652 1903 36692 1912
rect 36267 1784 36309 1793
rect 36267 1744 36268 1784
rect 36308 1744 36309 1784
rect 36267 1735 36309 1744
rect 34060 1324 34388 1364
rect 33100 1280 33140 1289
rect 33004 1240 33100 1280
rect 32716 1231 32756 1240
rect 33100 1231 33140 1240
rect 33483 1280 33525 1289
rect 33483 1240 33484 1280
rect 33524 1240 33525 1280
rect 33483 1231 33525 1240
rect 34060 1280 34100 1324
rect 34060 1231 34100 1240
rect 35595 1280 35637 1289
rect 35595 1240 35596 1280
rect 35636 1240 35637 1280
rect 35595 1231 35637 1240
rect 32908 1196 32948 1205
rect 32812 1156 32908 1196
rect 32619 860 32661 869
rect 32619 820 32620 860
rect 32660 820 32661 860
rect 32619 811 32661 820
rect 32812 785 32852 1156
rect 32908 1147 32948 1156
rect 33292 1196 33332 1205
rect 32811 776 32853 785
rect 32811 736 32812 776
rect 32852 736 32853 776
rect 32811 727 32853 736
rect 32523 692 32565 701
rect 32523 652 32524 692
rect 32564 652 32565 692
rect 32523 643 32565 652
rect 32907 692 32949 701
rect 32907 652 32908 692
rect 32948 652 32949 692
rect 32907 643 32949 652
rect 32908 80 32948 643
rect 33292 617 33332 1156
rect 33484 1146 33524 1231
rect 33675 1196 33717 1205
rect 33675 1156 33676 1196
rect 33716 1156 33717 1196
rect 33675 1147 33717 1156
rect 34444 1196 34484 1205
rect 33676 1062 33716 1147
rect 34252 944 34292 953
rect 34155 860 34197 869
rect 34252 860 34292 904
rect 34155 820 34156 860
rect 34196 820 34292 860
rect 34155 811 34197 820
rect 34444 701 34484 1156
rect 34828 1196 34868 1205
rect 35212 1196 35252 1205
rect 34635 944 34677 953
rect 34635 904 34636 944
rect 34676 904 34677 944
rect 34635 895 34677 904
rect 34636 810 34676 895
rect 34443 692 34485 701
rect 34443 652 34444 692
rect 34484 652 34485 692
rect 34443 643 34485 652
rect 34828 617 34868 1156
rect 34924 1156 35212 1196
rect 33291 608 33333 617
rect 33291 568 33292 608
rect 33332 568 33333 608
rect 33291 559 33333 568
rect 34059 608 34101 617
rect 34059 568 34060 608
rect 34100 568 34101 608
rect 34059 559 34101 568
rect 34827 608 34869 617
rect 34827 568 34828 608
rect 34868 568 34869 608
rect 34827 559 34869 568
rect 34060 80 34100 559
rect 34924 113 34964 1156
rect 35212 1147 35252 1156
rect 35596 1112 35636 1231
rect 36363 1196 36405 1205
rect 36363 1156 36364 1196
rect 36404 1156 36405 1196
rect 36363 1147 36405 1156
rect 35596 1063 35636 1072
rect 35019 944 35061 953
rect 35019 904 35020 944
rect 35060 904 35061 944
rect 35019 895 35061 904
rect 35020 810 35060 895
rect 35168 776 35536 785
rect 35208 736 35250 776
rect 35290 736 35332 776
rect 35372 736 35414 776
rect 35454 736 35496 776
rect 35168 727 35536 736
rect 34923 104 34965 113
rect 20427 55 20756 60
rect 20428 20 20756 55
rect 21368 0 21448 80
rect 22520 0 22600 80
rect 23672 0 23752 80
rect 24824 0 24904 80
rect 25976 0 26056 80
rect 27128 0 27208 80
rect 28280 0 28360 80
rect 29432 0 29512 80
rect 30584 0 30664 80
rect 31736 0 31816 80
rect 32888 0 32968 80
rect 34040 0 34120 80
rect 34923 64 34924 104
rect 34964 64 34965 104
rect 35211 104 35253 113
rect 35211 80 35212 104
rect 34923 55 34965 64
rect 35192 64 35212 80
rect 35252 80 35253 104
rect 36364 80 36404 1147
rect 36748 1112 36788 2575
rect 37036 1280 37076 3340
rect 37132 2624 37172 2633
rect 37132 2213 37172 2584
rect 37420 2540 37460 5440
rect 37516 3809 37556 7111
rect 37611 6656 37653 6665
rect 37611 6616 37612 6656
rect 37652 6616 37653 6656
rect 37611 6607 37653 6616
rect 37612 6522 37652 6607
rect 38284 6488 38324 6497
rect 37804 6404 37844 6413
rect 37804 6320 37844 6364
rect 37804 6280 38132 6320
rect 37900 5653 37940 5662
rect 37900 4304 37940 5613
rect 38092 5564 38132 6280
rect 38092 5515 38132 5524
rect 38284 5069 38324 6448
rect 38379 6488 38421 6497
rect 38379 6448 38380 6488
rect 38420 6448 38421 6488
rect 38379 6439 38421 6448
rect 38380 6354 38420 6439
rect 38476 5144 38516 7960
rect 38572 6497 38612 8203
rect 38668 7916 38708 8455
rect 38860 8252 38900 9295
rect 40300 8840 40340 9799
rect 41452 9680 41492 10471
rect 41547 10184 41589 10193
rect 41547 10144 41548 10184
rect 41588 10144 41589 10184
rect 41547 10135 41589 10144
rect 41452 9631 41492 9640
rect 40491 9512 40533 9521
rect 40491 9472 40492 9512
rect 40532 9472 40533 9512
rect 40491 9463 40533 9472
rect 41067 9512 41109 9521
rect 41067 9472 41068 9512
rect 41108 9472 41109 9512
rect 41067 9463 41109 9472
rect 40300 8791 40340 8800
rect 39147 8756 39189 8765
rect 39147 8716 39148 8756
rect 39188 8716 39189 8756
rect 39147 8707 39189 8716
rect 39916 8756 39956 8765
rect 40108 8756 40148 8765
rect 39956 8716 40052 8756
rect 39916 8707 39956 8716
rect 39052 8672 39092 8681
rect 38956 8632 39052 8672
rect 38956 8429 38996 8632
rect 39052 8623 39092 8632
rect 38955 8420 38997 8429
rect 38955 8380 38956 8420
rect 38996 8380 38997 8420
rect 38955 8371 38997 8380
rect 38860 8212 38996 8252
rect 38764 7916 38804 7925
rect 38668 7876 38764 7916
rect 38571 6488 38613 6497
rect 38571 6448 38572 6488
rect 38612 6448 38613 6488
rect 38571 6439 38613 6448
rect 38668 6320 38708 7876
rect 38764 7867 38804 7876
rect 38860 7916 38900 7925
rect 38860 6908 38900 7876
rect 38956 7160 38996 8212
rect 39148 7337 39188 8707
rect 39723 8504 39765 8513
rect 39723 8464 39724 8504
rect 39764 8464 39765 8504
rect 39723 8455 39765 8464
rect 39724 8370 39764 8455
rect 40012 8168 40052 8716
rect 40012 8119 40052 8128
rect 39340 8000 39380 8009
rect 39340 7841 39380 7960
rect 39820 7986 39860 7995
rect 39339 7832 39381 7841
rect 39339 7792 39340 7832
rect 39380 7792 39381 7832
rect 39339 7783 39381 7792
rect 39147 7328 39189 7337
rect 39147 7288 39148 7328
rect 39188 7288 39189 7328
rect 39147 7279 39189 7288
rect 38956 7111 38996 7120
rect 38380 5104 38516 5144
rect 38572 6280 38708 6320
rect 38764 6868 38900 6908
rect 38764 6488 38804 6868
rect 38283 5060 38325 5069
rect 38283 5020 38284 5060
rect 38324 5020 38325 5060
rect 38283 5011 38325 5020
rect 37804 4264 37940 4304
rect 37515 3800 37557 3809
rect 37515 3760 37516 3800
rect 37556 3760 37557 3800
rect 37515 3751 37557 3760
rect 37516 3464 37556 3751
rect 37516 3415 37556 3424
rect 37804 2885 37844 4264
rect 38380 4220 38420 5104
rect 38476 4976 38516 4985
rect 38476 4817 38516 4936
rect 38475 4808 38517 4817
rect 38475 4768 38476 4808
rect 38516 4768 38517 4808
rect 38475 4759 38517 4768
rect 38284 4180 38380 4220
rect 37899 4136 37941 4145
rect 37899 4096 37900 4136
rect 37940 4096 37941 4136
rect 37899 4087 37941 4096
rect 37996 4136 38036 4145
rect 38091 4136 38133 4145
rect 38036 4096 38092 4136
rect 38132 4096 38133 4136
rect 37996 4087 38036 4096
rect 38091 4087 38133 4096
rect 37900 4002 37940 4087
rect 38284 3725 38324 4180
rect 38380 4171 38420 4180
rect 38476 4220 38516 4229
rect 38572 4220 38612 6280
rect 38764 6077 38804 6448
rect 38859 6488 38901 6497
rect 38859 6448 38860 6488
rect 38900 6448 38901 6488
rect 38859 6439 38901 6448
rect 39340 6488 39380 7783
rect 39820 7589 39860 7946
rect 39819 7580 39861 7589
rect 39819 7540 39820 7580
rect 39860 7540 39861 7580
rect 39819 7531 39861 7540
rect 40108 7496 40148 8716
rect 40492 8756 40532 9463
rect 40587 9428 40629 9437
rect 40587 9388 40588 9428
rect 40628 9388 40629 9428
rect 40587 9379 40629 9388
rect 40875 9428 40917 9437
rect 40875 9388 40876 9428
rect 40916 9388 40917 9428
rect 40875 9379 40917 9388
rect 40492 8707 40532 8716
rect 40491 8168 40533 8177
rect 40491 8128 40492 8168
rect 40532 8128 40533 8168
rect 40491 8119 40533 8128
rect 40492 7916 40532 8119
rect 40492 7867 40532 7876
rect 40395 7580 40437 7589
rect 40395 7540 40396 7580
rect 40436 7540 40437 7580
rect 40395 7531 40437 7540
rect 39916 7456 40148 7496
rect 39340 6439 39380 6448
rect 39820 6474 39860 6483
rect 38763 6068 38805 6077
rect 38763 6028 38764 6068
rect 38804 6028 38805 6068
rect 38763 6019 38805 6028
rect 38860 5228 38900 6439
rect 39820 6329 39860 6434
rect 39819 6320 39861 6329
rect 39819 6280 39820 6320
rect 39860 6280 39861 6320
rect 39819 6271 39861 6280
rect 38955 5648 38997 5657
rect 38955 5608 38956 5648
rect 38996 5608 38997 5648
rect 38955 5599 38997 5608
rect 38956 5489 38996 5599
rect 38955 5480 38997 5489
rect 38955 5440 38956 5480
rect 38996 5440 38997 5480
rect 38955 5431 38997 5440
rect 38860 5188 38996 5228
rect 38667 5060 38709 5069
rect 38667 5020 38668 5060
rect 38708 5020 38709 5060
rect 38667 5011 38709 5020
rect 38668 4926 38708 5011
rect 38667 4808 38709 4817
rect 38667 4768 38668 4808
rect 38708 4768 38709 4808
rect 38667 4759 38709 4768
rect 38516 4180 38612 4220
rect 38476 4171 38516 4180
rect 38668 3809 38708 4759
rect 38859 4724 38901 4733
rect 38859 4684 38860 4724
rect 38900 4684 38901 4724
rect 38859 4675 38901 4684
rect 38860 4590 38900 4675
rect 38956 4136 38996 5188
rect 39243 5144 39285 5153
rect 39243 5104 39244 5144
rect 39284 5104 39285 5144
rect 39243 5095 39285 5104
rect 39052 4976 39092 4985
rect 39052 4817 39092 4936
rect 39051 4808 39093 4817
rect 39051 4768 39052 4808
rect 39092 4768 39093 4808
rect 39051 4759 39093 4768
rect 38956 4087 38996 4096
rect 38379 3800 38421 3809
rect 38379 3760 38380 3800
rect 38420 3760 38421 3800
rect 38379 3751 38421 3760
rect 38667 3800 38709 3809
rect 38667 3760 38668 3800
rect 38708 3760 38709 3800
rect 38667 3751 38709 3760
rect 38283 3716 38325 3725
rect 38283 3676 38284 3716
rect 38324 3676 38325 3716
rect 38283 3667 38325 3676
rect 37803 2876 37845 2885
rect 37803 2836 37804 2876
rect 37844 2836 37845 2876
rect 37803 2827 37845 2836
rect 38380 2624 38420 3751
rect 38764 3464 38804 3475
rect 38764 3389 38804 3424
rect 38763 3380 38805 3389
rect 38763 3340 38764 3380
rect 38804 3340 38805 3380
rect 38763 3331 38805 3340
rect 38571 2876 38613 2885
rect 38571 2836 38572 2876
rect 38612 2836 38613 2876
rect 38571 2827 38613 2836
rect 38572 2742 38612 2827
rect 38380 2575 38420 2584
rect 37228 2500 37460 2540
rect 37131 2204 37173 2213
rect 37131 2164 37132 2204
rect 37172 2164 37173 2204
rect 37131 2155 37173 2164
rect 37132 1961 37172 2155
rect 37131 1952 37173 1961
rect 37131 1912 37132 1952
rect 37172 1912 37173 1952
rect 37131 1903 37173 1912
rect 37036 1231 37076 1240
rect 37228 1280 37268 2500
rect 39244 2120 39284 5095
rect 39627 4892 39669 4901
rect 39627 4852 39628 4892
rect 39668 4852 39669 4892
rect 39627 4843 39669 4852
rect 39435 4724 39477 4733
rect 39435 4684 39436 4724
rect 39476 4684 39477 4724
rect 39435 4675 39477 4684
rect 39436 4150 39476 4675
rect 39436 4101 39476 4110
rect 39628 4052 39668 4843
rect 39628 4003 39668 4012
rect 39244 2071 39284 2080
rect 37900 1952 37940 1961
rect 37611 1448 37653 1457
rect 37611 1408 37612 1448
rect 37652 1408 37653 1448
rect 37611 1399 37653 1408
rect 37228 1231 37268 1240
rect 37612 1280 37652 1399
rect 37612 1231 37652 1240
rect 37419 1196 37461 1205
rect 37419 1156 37420 1196
rect 37460 1156 37461 1196
rect 37419 1147 37461 1156
rect 37804 1196 37844 1205
rect 36844 1112 36884 1121
rect 36748 1072 36844 1112
rect 36844 1063 36884 1072
rect 37420 1062 37460 1147
rect 37804 113 37844 1156
rect 37900 1121 37940 1912
rect 38380 1868 38420 1877
rect 39436 1868 39476 1877
rect 38420 1828 38708 1868
rect 38380 1819 38420 1828
rect 38187 1700 38229 1709
rect 38187 1660 38188 1700
rect 38228 1660 38229 1700
rect 38187 1651 38229 1660
rect 38188 1566 38228 1651
rect 37899 1112 37941 1121
rect 37899 1072 37900 1112
rect 37940 1072 37941 1112
rect 37899 1063 37941 1072
rect 37515 104 37557 113
rect 37515 80 37516 104
rect 35252 64 35272 80
rect 35192 0 35272 64
rect 36344 0 36424 80
rect 37496 64 37516 80
rect 37556 80 37557 104
rect 37803 104 37845 113
rect 37556 64 37576 80
rect 37496 0 37576 64
rect 37803 64 37804 104
rect 37844 64 37845 104
rect 38668 80 38708 1828
rect 37803 55 37845 64
rect 38648 0 38728 80
rect 39436 60 39476 1828
rect 39628 1868 39668 1879
rect 39628 1793 39668 1828
rect 39627 1784 39669 1793
rect 39627 1744 39628 1784
rect 39668 1744 39669 1784
rect 39627 1735 39669 1744
rect 39820 1700 39860 1709
rect 39820 1457 39860 1660
rect 39819 1448 39861 1457
rect 39819 1408 39820 1448
rect 39860 1408 39861 1448
rect 39819 1399 39861 1408
rect 39916 953 39956 7456
rect 40396 7412 40436 7531
rect 40396 7363 40436 7372
rect 40204 7160 40244 7169
rect 40108 7120 40204 7160
rect 40012 6572 40052 6581
rect 40012 6413 40052 6532
rect 40011 6404 40053 6413
rect 40011 6364 40012 6404
rect 40052 6364 40053 6404
rect 40011 6355 40053 6364
rect 40108 5648 40148 7120
rect 40204 7111 40244 7120
rect 40204 6329 40244 6414
rect 40396 6413 40436 6498
rect 40395 6404 40437 6413
rect 40395 6364 40396 6404
rect 40436 6364 40437 6404
rect 40395 6355 40437 6364
rect 40203 6320 40245 6329
rect 40203 6280 40204 6320
rect 40244 6280 40245 6320
rect 40203 6271 40245 6280
rect 40299 6236 40341 6245
rect 40299 6196 40300 6236
rect 40340 6196 40341 6236
rect 40299 6187 40341 6196
rect 40300 5900 40340 6187
rect 40396 5900 40436 5909
rect 40300 5860 40396 5900
rect 40396 5851 40436 5860
rect 40204 5648 40244 5676
rect 40108 5608 40204 5648
rect 40108 4817 40148 5608
rect 40204 5599 40244 5608
rect 40300 4976 40340 4985
rect 40107 4808 40149 4817
rect 40107 4768 40108 4808
rect 40148 4768 40149 4808
rect 40107 4759 40149 4768
rect 40300 3641 40340 4936
rect 40492 4733 40532 4818
rect 40491 4724 40533 4733
rect 40491 4684 40492 4724
rect 40532 4684 40533 4724
rect 40491 4675 40533 4684
rect 40491 4472 40533 4481
rect 40491 4432 40492 4472
rect 40532 4432 40533 4472
rect 40491 4423 40533 4432
rect 40492 4220 40532 4423
rect 40492 4171 40532 4180
rect 40299 3632 40341 3641
rect 40299 3592 40300 3632
rect 40340 3592 40341 3632
rect 40299 3583 40341 3592
rect 40491 3380 40533 3389
rect 40491 3340 40492 3380
rect 40532 3340 40533 3380
rect 40491 3331 40533 3340
rect 40492 3246 40532 3331
rect 40492 2708 40532 2717
rect 40492 2297 40532 2668
rect 40491 2288 40533 2297
rect 40491 2248 40492 2288
rect 40532 2248 40533 2288
rect 40491 2239 40533 2248
rect 40396 2120 40436 2129
rect 40588 2120 40628 9379
rect 40876 9294 40916 9379
rect 41068 9344 41108 9463
rect 41260 9428 41300 9439
rect 41260 9353 41300 9388
rect 41068 9295 41108 9304
rect 41259 9344 41301 9353
rect 41259 9304 41260 9344
rect 41300 9304 41301 9344
rect 41259 9295 41301 9304
rect 41259 9176 41301 9185
rect 41259 9136 41260 9176
rect 41300 9136 41301 9176
rect 41259 9127 41301 9136
rect 40683 8924 40725 8933
rect 40683 8884 40684 8924
rect 40724 8884 40725 8924
rect 40683 8875 40725 8884
rect 40684 8840 40724 8875
rect 40684 8789 40724 8800
rect 40875 8756 40917 8765
rect 40875 8716 40876 8756
rect 40916 8716 40917 8756
rect 40875 8707 40917 8716
rect 41260 8756 41300 9127
rect 41451 9092 41493 9101
rect 41451 9052 41452 9092
rect 41492 9052 41493 9092
rect 41451 9043 41493 9052
rect 41452 8840 41492 9043
rect 41452 8791 41492 8800
rect 41260 8707 41300 8716
rect 40876 8622 40916 8707
rect 41067 8504 41109 8513
rect 41067 8464 41068 8504
rect 41108 8464 41109 8504
rect 41067 8455 41109 8464
rect 41068 8370 41108 8455
rect 41259 8420 41301 8429
rect 41259 8380 41260 8420
rect 41300 8380 41301 8420
rect 41259 8371 41301 8380
rect 40683 8168 40725 8177
rect 40683 8128 40684 8168
rect 40724 8128 40725 8168
rect 40683 8119 40725 8128
rect 40684 8034 40724 8119
rect 40876 7916 40916 7925
rect 41260 7916 41300 8371
rect 41452 8168 41492 8177
rect 41548 8168 41588 10135
rect 41492 8128 41588 8168
rect 41452 8119 41492 8128
rect 40916 7876 41012 7916
rect 40876 7867 40916 7876
rect 40875 7244 40917 7253
rect 40875 7204 40876 7244
rect 40916 7204 40917 7244
rect 40875 7195 40917 7204
rect 40876 7110 40916 7195
rect 40875 6992 40917 7001
rect 40875 6952 40876 6992
rect 40916 6952 40917 6992
rect 40875 6943 40917 6952
rect 40876 6404 40916 6943
rect 40876 6355 40916 6364
rect 40779 5900 40821 5909
rect 40779 5860 40780 5900
rect 40820 5860 40821 5900
rect 40779 5851 40821 5860
rect 40683 4892 40725 4901
rect 40683 4852 40684 4892
rect 40724 4852 40725 4892
rect 40683 4843 40725 4852
rect 40684 4758 40724 4843
rect 40683 4472 40725 4481
rect 40683 4432 40684 4472
rect 40724 4432 40725 4472
rect 40683 4423 40725 4432
rect 40684 4388 40724 4423
rect 40684 4337 40724 4348
rect 40780 4220 40820 5851
rect 40875 5732 40917 5741
rect 40875 5692 40876 5732
rect 40916 5692 40917 5732
rect 40875 5683 40917 5692
rect 40876 5598 40916 5683
rect 40875 5396 40917 5405
rect 40875 5356 40876 5396
rect 40916 5356 40917 5396
rect 40875 5347 40917 5356
rect 40876 4892 40916 5347
rect 40972 4985 41012 7876
rect 41260 7867 41300 7876
rect 41067 7832 41109 7841
rect 41067 7792 41068 7832
rect 41108 7792 41109 7832
rect 41067 7783 41109 7792
rect 41068 7698 41108 7783
rect 41355 7748 41397 7757
rect 41355 7708 41356 7748
rect 41396 7708 41397 7748
rect 41355 7699 41397 7708
rect 41260 7244 41300 7253
rect 41164 7204 41260 7244
rect 41067 7160 41109 7169
rect 41067 7120 41068 7160
rect 41108 7120 41109 7160
rect 41067 7111 41109 7120
rect 41068 6992 41108 7111
rect 41068 6943 41108 6952
rect 41067 6488 41109 6497
rect 41067 6448 41068 6488
rect 41108 6448 41109 6488
rect 41067 6439 41109 6448
rect 41068 6320 41108 6439
rect 41068 6271 41108 6280
rect 41067 6152 41109 6161
rect 41067 6112 41068 6152
rect 41108 6112 41109 6152
rect 41067 6103 41109 6112
rect 41068 5900 41108 6103
rect 41068 5851 41108 5860
rect 41164 5657 41204 7204
rect 41260 7195 41300 7204
rect 41260 6413 41300 6498
rect 41259 6404 41301 6413
rect 41259 6364 41260 6404
rect 41300 6364 41301 6404
rect 41259 6355 41301 6364
rect 41260 5732 41300 5741
rect 41163 5648 41205 5657
rect 41163 5608 41164 5648
rect 41204 5608 41205 5648
rect 41163 5599 41205 5608
rect 41067 5480 41109 5489
rect 41067 5440 41068 5480
rect 41108 5440 41109 5480
rect 41067 5431 41109 5440
rect 40971 4976 41013 4985
rect 40971 4936 40972 4976
rect 41012 4936 41013 4976
rect 40971 4927 41013 4936
rect 40876 4843 40916 4852
rect 41068 4808 41108 5431
rect 41260 5237 41300 5692
rect 41259 5228 41301 5237
rect 41259 5188 41260 5228
rect 41300 5188 41301 5228
rect 41259 5179 41301 5188
rect 41260 4892 41300 4901
rect 41356 4892 41396 7699
rect 41451 7496 41493 7505
rect 41451 7456 41452 7496
rect 41492 7456 41493 7496
rect 41451 7447 41493 7456
rect 41452 7412 41492 7447
rect 41452 7361 41492 7372
rect 41451 6824 41493 6833
rect 41451 6784 41452 6824
rect 41492 6784 41493 6824
rect 41451 6775 41493 6784
rect 41452 6656 41492 6775
rect 41452 6607 41492 6616
rect 41451 5816 41493 5825
rect 41451 5776 41452 5816
rect 41492 5776 41493 5816
rect 41451 5767 41493 5776
rect 41452 5682 41492 5767
rect 41451 5144 41493 5153
rect 41451 5104 41452 5144
rect 41492 5104 41493 5144
rect 41451 5095 41493 5104
rect 41300 4852 41396 4892
rect 41260 4843 41300 4852
rect 41068 4759 41108 4768
rect 41163 4808 41205 4817
rect 41163 4768 41164 4808
rect 41204 4768 41205 4808
rect 41163 4759 41205 4768
rect 41452 4808 41492 5095
rect 41452 4759 41492 4768
rect 41068 4388 41108 4397
rect 41164 4388 41204 4759
rect 41259 4640 41301 4649
rect 41259 4600 41260 4640
rect 41300 4600 41301 4640
rect 41259 4591 41301 4600
rect 41108 4348 41204 4388
rect 41068 4339 41108 4348
rect 40876 4220 40916 4229
rect 40780 4180 40876 4220
rect 40876 4171 40916 4180
rect 41260 4220 41300 4591
rect 41260 4171 41300 4180
rect 41451 4136 41493 4145
rect 41451 4096 41452 4136
rect 41492 4096 41493 4136
rect 41451 4087 41493 4096
rect 41452 3968 41492 4087
rect 41452 3919 41492 3928
rect 41067 3800 41109 3809
rect 41067 3760 41068 3800
rect 41108 3760 41109 3800
rect 41067 3751 41109 3760
rect 40875 3632 40917 3641
rect 40875 3592 40876 3632
rect 40916 3592 40917 3632
rect 40875 3583 40917 3592
rect 41068 3632 41108 3751
rect 41068 3583 41108 3592
rect 40683 3464 40725 3473
rect 40683 3424 40684 3464
rect 40724 3424 40725 3464
rect 40683 3415 40725 3424
rect 40684 3296 40724 3415
rect 40876 3380 40916 3583
rect 40876 3331 40916 3340
rect 40684 3247 40724 3256
rect 41067 3128 41109 3137
rect 41067 3088 41068 3128
rect 41108 3088 41109 3128
rect 41067 3079 41109 3088
rect 41068 2876 41108 3079
rect 41259 2960 41301 2969
rect 41259 2920 41260 2960
rect 41300 2920 41301 2960
rect 41259 2911 41301 2920
rect 41068 2827 41108 2836
rect 40683 2792 40725 2801
rect 40683 2752 40684 2792
rect 40724 2752 40725 2792
rect 40683 2743 40725 2752
rect 40684 2658 40724 2743
rect 40876 2708 40916 2717
rect 40779 2540 40821 2549
rect 40779 2500 40780 2540
rect 40820 2500 40821 2540
rect 40779 2491 40821 2500
rect 40436 2080 40628 2120
rect 40396 2071 40436 2080
rect 40491 1952 40533 1961
rect 40491 1912 40492 1952
rect 40532 1912 40533 1952
rect 40491 1903 40533 1912
rect 40011 1868 40053 1877
rect 40011 1828 40012 1868
rect 40052 1828 40053 1868
rect 40011 1819 40053 1828
rect 40012 1734 40052 1819
rect 40204 1700 40244 1709
rect 39915 944 39957 953
rect 39915 904 39916 944
rect 39956 904 39957 944
rect 39915 895 39957 904
rect 40204 449 40244 1660
rect 40492 1196 40532 1903
rect 40492 1147 40532 1156
rect 40588 1868 40628 1877
rect 40780 1868 40820 2491
rect 40876 2381 40916 2668
rect 41260 2708 41300 2911
rect 41260 2659 41300 2668
rect 41451 2456 41493 2465
rect 41451 2416 41452 2456
rect 41492 2416 41493 2456
rect 41451 2407 41493 2416
rect 40875 2372 40917 2381
rect 40875 2332 40876 2372
rect 40916 2332 40917 2372
rect 40875 2323 40917 2332
rect 41452 2322 41492 2407
rect 41067 2120 41109 2129
rect 41067 2080 41068 2120
rect 41108 2080 41109 2120
rect 41067 2071 41109 2080
rect 41068 1986 41108 2071
rect 40876 1868 40916 1877
rect 41260 1868 41300 1877
rect 40780 1828 40876 1868
rect 40203 440 40245 449
rect 40203 400 40204 440
rect 40244 400 40245 440
rect 40203 391 40245 400
rect 39627 104 39669 113
rect 39627 64 39628 104
rect 39668 64 39669 104
rect 39819 104 39861 113
rect 39819 80 39820 104
rect 39627 60 39669 64
rect 39436 55 39669 60
rect 39800 64 39820 80
rect 39860 80 39861 104
rect 39860 64 39880 80
rect 39436 20 39668 55
rect 39800 0 39880 64
rect 40588 60 40628 1828
rect 40876 1819 40916 1828
rect 41164 1828 41260 1868
rect 41164 1289 41204 1828
rect 41260 1819 41300 1828
rect 41451 1784 41493 1793
rect 41451 1744 41452 1784
rect 41492 1744 41493 1784
rect 41451 1735 41493 1744
rect 41452 1650 41492 1735
rect 41163 1280 41205 1289
rect 41163 1240 41164 1280
rect 41204 1240 41205 1280
rect 41163 1231 41205 1240
rect 40875 1196 40917 1205
rect 40875 1156 40876 1196
rect 40916 1156 40917 1196
rect 40875 1147 40917 1156
rect 41260 1196 41300 1205
rect 40683 1112 40725 1121
rect 40683 1072 40684 1112
rect 40724 1072 40725 1112
rect 40683 1063 40725 1072
rect 40684 944 40724 1063
rect 40876 1062 40916 1147
rect 41260 1037 41300 1156
rect 41259 1028 41301 1037
rect 41259 988 41260 1028
rect 41300 988 41301 1028
rect 41259 979 41301 988
rect 40684 895 40724 904
rect 41068 944 41108 953
rect 41068 197 41108 904
rect 41452 944 41492 953
rect 41452 785 41492 904
rect 41451 776 41493 785
rect 41451 736 41452 776
rect 41492 736 41493 776
rect 41451 727 41493 736
rect 41067 188 41109 197
rect 41067 148 41068 188
rect 41108 148 41109 188
rect 41067 139 41109 148
rect 40779 104 40821 113
rect 40779 64 40780 104
rect 40820 64 40821 104
rect 40971 104 41013 113
rect 40971 80 40972 104
rect 40779 60 40821 64
rect 40588 55 40821 60
rect 40952 64 40972 80
rect 41012 80 41013 104
rect 41012 64 41032 80
rect 40588 20 40820 55
rect 40952 0 41032 64
<< via2 >>
rect 8908 10648 8948 10688
rect 9484 10648 9524 10688
rect 2764 10144 2804 10184
rect 1900 9892 1940 9932
rect 1900 9136 1940 9176
rect 1804 8968 1844 9008
rect 1420 8128 1460 8168
rect 1228 6448 1268 6488
rect 1228 5440 1268 5480
rect 1516 6784 1556 6824
rect 1708 8128 1748 8168
rect 1900 8800 1940 8840
rect 2092 8716 2132 8756
rect 1900 8464 1940 8504
rect 2092 8380 2132 8420
rect 2476 7120 2516 7160
rect 1900 6868 1940 6908
rect 1708 6532 1748 6572
rect 1612 6280 1652 6320
rect 1516 5860 1556 5900
rect 1420 5356 1460 5396
rect 1900 6280 1940 6320
rect 1708 5944 1748 5984
rect 1804 5188 1844 5228
rect 1708 4936 1748 4976
rect 4928 9808 4968 9848
rect 5010 9808 5050 9848
rect 5092 9808 5132 9848
rect 5174 9808 5214 9848
rect 5256 9808 5296 9848
rect 3724 9640 3764 9680
rect 3532 9556 3572 9596
rect 3436 9472 3476 9512
rect 3340 9388 3380 9428
rect 3820 9472 3860 9512
rect 3628 9388 3668 9428
rect 3532 9304 3572 9344
rect 3688 9052 3728 9092
rect 3770 9052 3810 9092
rect 3852 9052 3892 9092
rect 3934 9052 3974 9092
rect 4016 9052 4056 9092
rect 3724 8632 3764 8672
rect 3244 8548 3284 8588
rect 3340 8128 3380 8168
rect 3532 8212 3572 8252
rect 3820 8464 3860 8504
rect 3916 8128 3956 8168
rect 5740 9640 5780 9680
rect 5356 9556 5396 9596
rect 4204 8632 4244 8672
rect 4396 9472 4436 9512
rect 4300 8296 4340 8336
rect 3688 7540 3728 7580
rect 3770 7540 3810 7580
rect 3852 7540 3892 7580
rect 3934 7540 3974 7580
rect 4016 7540 4056 7580
rect 4492 9388 4532 9428
rect 4876 9304 4916 9344
rect 5164 8968 5204 9008
rect 4684 8800 4724 8840
rect 4588 8212 4628 8252
rect 4492 7960 4532 8000
rect 4972 8548 5012 8588
rect 5932 9556 5972 9596
rect 5452 8968 5492 9008
rect 5548 8800 5588 8840
rect 5836 9304 5876 9344
rect 5932 8632 5972 8672
rect 5260 8464 5300 8504
rect 4928 8296 4968 8336
rect 5010 8296 5050 8336
rect 5092 8296 5132 8336
rect 5174 8296 5214 8336
rect 5256 8296 5296 8336
rect 5356 7960 5396 8000
rect 5836 8296 5876 8336
rect 5644 7960 5684 8000
rect 5452 7792 5492 7832
rect 5356 7708 5396 7748
rect 4684 7624 4724 7664
rect 2764 6952 2804 6992
rect 3820 7120 3860 7160
rect 2860 6448 2900 6488
rect 2476 5440 2516 5480
rect 2476 5188 2516 5228
rect 3052 5188 3092 5228
rect 4108 7120 4148 7160
rect 4396 7120 4436 7160
rect 4012 7036 4052 7076
rect 3916 6700 3956 6740
rect 4588 7204 4628 7244
rect 4588 6700 4628 6740
rect 4012 6448 4052 6488
rect 4204 6280 4244 6320
rect 3688 6028 3728 6068
rect 3770 6028 3810 6068
rect 3852 6028 3892 6068
rect 3934 6028 3974 6068
rect 4016 6028 4056 6068
rect 4492 6532 4532 6572
rect 4204 5944 4244 5984
rect 4396 5944 4436 5984
rect 4780 7120 4820 7160
rect 4928 6784 4968 6824
rect 5010 6784 5050 6824
rect 5092 6784 5132 6824
rect 5174 6784 5214 6824
rect 5256 6784 5296 6824
rect 4684 6280 4724 6320
rect 4780 6196 4820 6236
rect 4780 6028 4820 6068
rect 4300 5776 4340 5816
rect 4780 5608 4820 5648
rect 5164 6448 5204 6488
rect 5164 6280 5204 6320
rect 5164 5608 5204 5648
rect 5932 8212 5972 8252
rect 6988 9472 7028 9512
rect 7852 9472 7892 9512
rect 7180 9388 7220 9428
rect 7564 9388 7604 9428
rect 7468 9304 7508 9344
rect 6604 8800 6644 8840
rect 6124 8632 6164 8672
rect 6220 8296 6260 8336
rect 6028 8128 6068 8168
rect 6892 8800 6932 8840
rect 6700 8632 6740 8672
rect 6604 8212 6644 8252
rect 6316 7792 6356 7832
rect 6028 7708 6068 7748
rect 5644 6784 5684 6824
rect 5836 7036 5876 7076
rect 5740 6364 5780 6404
rect 5644 6196 5684 6236
rect 6220 6952 6260 6992
rect 6028 6448 6068 6488
rect 6220 6364 6260 6404
rect 6124 6280 6164 6320
rect 6316 6280 6356 6320
rect 5836 5944 5876 5984
rect 5740 5776 5780 5816
rect 5548 5608 5588 5648
rect 3532 5020 3572 5060
rect 2764 4348 2804 4388
rect 2668 3928 2708 3968
rect 3148 4936 3188 4976
rect 3340 4852 3380 4892
rect 3148 4768 3188 4808
rect 3436 4684 3476 4724
rect 3340 4180 3380 4220
rect 2764 3760 2804 3800
rect 3052 3760 3092 3800
rect 3724 4852 3764 4892
rect 4108 4936 4148 4976
rect 4396 4768 4436 4808
rect 3628 4684 3668 4724
rect 3916 4684 3956 4724
rect 3688 4516 3728 4556
rect 3770 4516 3810 4556
rect 3852 4516 3892 4556
rect 3934 4516 3974 4556
rect 4016 4516 4056 4556
rect 3532 4180 3572 4220
rect 4012 4180 4052 4220
rect 3052 3424 3092 3464
rect 3436 3424 3476 3464
rect 4108 4096 4148 4136
rect 4012 3844 4052 3884
rect 4108 3760 4148 3800
rect 3820 3592 3860 3632
rect 3724 3508 3764 3548
rect 3820 3424 3860 3464
rect 4108 3424 4148 3464
rect 4396 4600 4436 4640
rect 4300 4516 4340 4556
rect 5260 5440 5300 5480
rect 4928 5272 4968 5312
rect 5010 5272 5050 5312
rect 5092 5272 5132 5312
rect 5174 5272 5214 5312
rect 5256 5272 5296 5312
rect 5164 5020 5204 5060
rect 5260 4936 5300 4976
rect 5836 5608 5876 5648
rect 5452 5440 5492 5480
rect 6124 5944 6164 5984
rect 4588 4768 4628 4808
rect 5068 4768 5108 4808
rect 4492 4516 4532 4556
rect 4492 4264 4532 4304
rect 4588 4096 4628 4136
rect 4492 3760 4532 3800
rect 4588 3676 4628 3716
rect 5068 4180 5108 4220
rect 4876 4096 4916 4136
rect 5644 5188 5684 5228
rect 5932 5188 5972 5228
rect 5740 5020 5780 5060
rect 6316 5272 6356 5312
rect 6220 5188 6260 5228
rect 6508 7120 6548 7160
rect 6700 6952 6740 6992
rect 6604 6532 6644 6572
rect 6508 6448 6548 6488
rect 6796 6280 6836 6320
rect 6604 6196 6644 6236
rect 6508 6112 6548 6152
rect 6412 5020 6452 5060
rect 6028 4768 6068 4808
rect 6124 4684 6164 4724
rect 5356 4432 5396 4472
rect 5452 4096 5492 4136
rect 4928 3760 4968 3800
rect 5010 3760 5050 3800
rect 5092 3760 5132 3800
rect 5174 3760 5214 3800
rect 5256 3760 5296 3800
rect 4876 3592 4916 3632
rect 5068 3592 5108 3632
rect 5932 3676 5972 3716
rect 5740 3508 5780 3548
rect 3916 3340 3956 3380
rect 3340 3256 3380 3296
rect 4108 3172 4148 3212
rect 3688 3004 3728 3044
rect 3770 3004 3810 3044
rect 3852 3004 3892 3044
rect 3934 3004 3974 3044
rect 4016 3004 4056 3044
rect 4396 2920 4436 2960
rect 3340 2752 3380 2792
rect 3436 2668 3476 2708
rect 1804 1828 1844 1868
rect 2476 1072 2516 1112
rect 3724 2584 3764 2624
rect 3148 2164 3188 2204
rect 3532 2164 3572 2204
rect 3340 1660 3380 1700
rect 3916 1912 3956 1952
rect 4204 2248 4244 2288
rect 3820 1660 3860 1700
rect 3688 1492 3728 1532
rect 3770 1492 3810 1532
rect 3852 1492 3892 1532
rect 3934 1492 3974 1532
rect 4016 1492 4056 1532
rect 4108 1072 4148 1112
rect 4972 2668 5012 2708
rect 4492 2584 4532 2624
rect 4876 2584 4916 2624
rect 5644 3424 5684 3464
rect 6796 5608 6836 5648
rect 6988 7876 7028 7916
rect 7372 8632 7412 8672
rect 7276 7120 7316 7160
rect 7180 6700 7220 6740
rect 6988 6364 7028 6404
rect 6988 5944 7028 5984
rect 6988 5776 7028 5816
rect 6892 5188 6932 5228
rect 7180 6448 7220 6488
rect 7564 8800 7604 8840
rect 8812 9052 8852 9092
rect 9676 9808 9716 9848
rect 8428 8716 8468 8756
rect 9196 8716 9236 8756
rect 8812 8632 8852 8672
rect 7468 7456 7508 7496
rect 8044 7120 8084 7160
rect 7468 6616 7508 6656
rect 9292 7540 9332 7580
rect 8812 6448 8852 6488
rect 7564 6280 7604 6320
rect 8716 6280 8756 6320
rect 7372 6196 7412 6236
rect 7084 5440 7124 5480
rect 7276 5440 7316 5480
rect 6700 4852 6740 4892
rect 6508 4096 6548 4136
rect 6220 3928 6260 3968
rect 6028 3340 6068 3380
rect 6604 3340 6644 3380
rect 5164 3172 5204 3212
rect 5548 2668 5588 2708
rect 4588 2248 4628 2288
rect 4928 2248 4968 2288
rect 5010 2248 5050 2288
rect 5092 2248 5132 2288
rect 5174 2248 5214 2288
rect 5256 2248 5296 2288
rect 5068 1996 5108 2036
rect 5452 2164 5492 2204
rect 4300 1660 4340 1700
rect 4396 1576 4436 1616
rect 4396 1156 4436 1196
rect 4780 1072 4820 1112
rect 5068 1156 5108 1196
rect 3916 988 3956 1028
rect 4684 988 4724 1028
rect 5356 1912 5396 1952
rect 5356 988 5396 1028
rect 4108 904 4148 944
rect 4972 904 5012 944
rect 4928 736 4968 776
rect 5010 736 5050 776
rect 5092 736 5132 776
rect 5174 736 5214 776
rect 5256 736 5296 776
rect 5356 400 5396 440
rect 5644 2584 5684 2624
rect 7084 4264 7124 4304
rect 5740 2248 5780 2288
rect 6412 2080 6452 2120
rect 5548 1996 5588 2036
rect 5740 1996 5780 2036
rect 6508 1912 6548 1952
rect 6412 904 6452 944
rect 6988 4096 7028 4136
rect 7276 5188 7316 5228
rect 7468 5440 7508 5480
rect 7660 5860 7700 5900
rect 7948 5608 7988 5648
rect 7660 5440 7700 5480
rect 7660 5188 7700 5228
rect 7468 4264 7508 4304
rect 7564 4180 7604 4220
rect 7084 3760 7124 3800
rect 7372 3424 7412 3464
rect 7468 3172 7508 3212
rect 7276 2416 7316 2456
rect 7948 4264 7988 4304
rect 7756 3760 7796 3800
rect 7756 3004 7796 3044
rect 8620 3928 8660 3968
rect 7468 2080 7508 2120
rect 7276 1660 7316 1700
rect 6604 64 6644 104
rect 7852 2584 7892 2624
rect 8908 6280 8948 6320
rect 10156 9808 10196 9848
rect 10060 9136 10100 9176
rect 9964 9052 10004 9092
rect 10348 9388 10388 9428
rect 10348 8968 10388 9008
rect 10252 8800 10292 8840
rect 9772 8632 9812 8672
rect 10252 8674 10292 8714
rect 10540 9976 10580 10016
rect 10540 9136 10580 9176
rect 10444 7372 10484 7412
rect 9484 7204 9524 7244
rect 9868 7204 9908 7244
rect 9868 6700 9908 6740
rect 9484 6616 9524 6656
rect 9580 6448 9620 6488
rect 9964 6280 10004 6320
rect 9292 5944 9332 5984
rect 9292 5608 9332 5648
rect 9100 4936 9140 4976
rect 9100 4012 9140 4052
rect 8908 3256 8948 3296
rect 9772 5776 9812 5816
rect 9580 5608 9620 5648
rect 9580 5272 9620 5312
rect 9772 5272 9812 5312
rect 9484 4936 9524 4976
rect 10348 6952 10388 6992
rect 9964 4936 10004 4976
rect 10252 4936 10292 4976
rect 9868 4432 9908 4472
rect 9388 3592 9428 3632
rect 9100 2668 9140 2708
rect 8908 2584 8948 2624
rect 8812 2164 8852 2204
rect 7756 1912 7796 1952
rect 8524 1912 8564 1952
rect 10252 3760 10292 3800
rect 10636 8716 10676 8756
rect 11116 10564 11156 10604
rect 11116 8968 11156 9008
rect 11500 10396 11540 10436
rect 11404 9052 11444 9092
rect 11020 8800 11060 8840
rect 11212 8800 11252 8840
rect 10828 8632 10868 8672
rect 10924 8548 10964 8588
rect 10924 8212 10964 8252
rect 11020 7540 11060 7580
rect 10924 7372 10964 7412
rect 10732 7288 10772 7328
rect 10828 7120 10868 7160
rect 10540 6952 10580 6992
rect 10828 6448 10868 6488
rect 10732 6364 10772 6404
rect 10636 6280 10676 6320
rect 10540 5776 10580 5816
rect 10828 6280 10868 6320
rect 10732 5860 10772 5900
rect 10444 4936 10484 4976
rect 10540 4852 10580 4892
rect 10540 4096 10580 4136
rect 10348 2920 10388 2960
rect 10444 2752 10484 2792
rect 9484 1828 9524 1868
rect 7756 1576 7796 1616
rect 8524 1576 8564 1616
rect 8140 1156 8180 1196
rect 9388 1240 9428 1280
rect 10156 1912 10196 1952
rect 10540 1912 10580 1952
rect 11500 8632 11540 8672
rect 11500 7372 11540 7412
rect 11500 7204 11540 7244
rect 11020 6448 11060 6488
rect 11020 5860 11060 5900
rect 11020 5608 11060 5648
rect 10828 4852 10868 4892
rect 11020 4600 11060 4640
rect 11020 4180 11060 4220
rect 10924 4096 10964 4136
rect 11020 3088 11060 3128
rect 11500 6868 11540 6908
rect 11692 9052 11732 9092
rect 11788 8800 11828 8840
rect 11884 8632 11924 8672
rect 11788 8044 11828 8084
rect 11692 7876 11732 7916
rect 11884 7372 11924 7412
rect 12172 9640 12212 9680
rect 12172 8968 12212 9008
rect 12268 8632 12308 8672
rect 12076 7540 12116 7580
rect 12076 7372 12116 7412
rect 11500 4096 11540 4136
rect 11308 4012 11348 4052
rect 11980 6448 12020 6488
rect 11980 6196 12020 6236
rect 12172 6532 12212 6572
rect 12364 7960 12404 8000
rect 12268 6280 12308 6320
rect 12268 5020 12308 5060
rect 11788 4684 11828 4724
rect 12076 4684 12116 4724
rect 12172 4432 12212 4472
rect 12076 3844 12116 3884
rect 11212 2920 11252 2960
rect 11212 2668 11252 2708
rect 11020 2080 11060 2120
rect 10636 1828 10676 1868
rect 10252 1240 10292 1280
rect 8716 1072 8756 1112
rect 9868 1072 9908 1112
rect 7948 904 7988 944
rect 8716 904 8756 944
rect 9772 904 9812 944
rect 11020 1240 11060 1280
rect 11404 2836 11444 2876
rect 11404 2416 11444 2456
rect 12268 3424 12308 3464
rect 12268 2668 12308 2708
rect 11788 1828 11828 1868
rect 12556 8800 12596 8840
rect 13132 10144 13172 10184
rect 13132 9472 13172 9512
rect 12940 9136 12980 9176
rect 12940 8968 12980 9008
rect 12748 7960 12788 8000
rect 12556 7876 12596 7916
rect 12556 6700 12596 6740
rect 12460 6532 12500 6572
rect 12460 5944 12500 5984
rect 12748 7204 12788 7244
rect 13036 8632 13076 8672
rect 13324 9052 13364 9092
rect 13900 9640 13940 9680
rect 14188 9640 14228 9680
rect 14284 8968 14324 9008
rect 14092 8800 14132 8840
rect 13804 8464 13844 8504
rect 13996 8296 14036 8336
rect 14284 8296 14324 8336
rect 14092 8212 14132 8252
rect 14476 8800 14516 8840
rect 14860 9556 14900 9596
rect 14956 9472 14996 9512
rect 15244 9640 15284 9680
rect 15052 9136 15092 9176
rect 15820 10060 15860 10100
rect 16204 9808 16244 9848
rect 16396 9640 16436 9680
rect 14860 8632 14900 8672
rect 14092 7960 14132 8000
rect 14668 7960 14708 8000
rect 13132 7372 13172 7412
rect 12940 7204 12980 7244
rect 13132 6952 13172 6992
rect 13036 6364 13076 6404
rect 12460 4936 12500 4976
rect 12556 4600 12596 4640
rect 12556 3844 12596 3884
rect 13228 4012 13268 4052
rect 13132 3676 13172 3716
rect 13036 2668 13076 2708
rect 12652 1828 12692 1868
rect 12364 1072 12404 1112
rect 14380 7372 14420 7412
rect 13516 7120 13556 7160
rect 14380 7036 14420 7076
rect 13516 6532 13556 6572
rect 13708 6448 13748 6488
rect 14188 6448 14228 6488
rect 14476 6448 14516 6488
rect 13804 6364 13844 6404
rect 13708 5608 13748 5648
rect 13804 4852 13844 4892
rect 13804 4348 13844 4388
rect 13612 4096 13652 4136
rect 13708 3676 13748 3716
rect 13516 3424 13556 3464
rect 14860 5944 14900 5984
rect 14284 5608 14324 5648
rect 14860 5608 14900 5648
rect 15436 8800 15476 8840
rect 15628 8800 15668 8840
rect 16012 8800 16052 8840
rect 15244 8464 15284 8504
rect 15148 8128 15188 8168
rect 15052 7708 15092 7748
rect 15820 8632 15860 8672
rect 16492 9388 16532 9428
rect 15724 8296 15764 8336
rect 16204 8296 16244 8336
rect 15340 8212 15380 8252
rect 15340 7792 15380 7832
rect 15628 7792 15668 7832
rect 15244 7624 15284 7664
rect 15340 6532 15380 6572
rect 16300 7876 16340 7916
rect 15916 7204 15956 7244
rect 15532 5860 15572 5900
rect 14284 3508 14324 3548
rect 13900 3424 13940 3464
rect 13804 2752 13844 2792
rect 13420 1828 13460 1868
rect 13036 988 13076 1028
rect 13324 988 13364 1028
rect 10348 64 10388 104
rect 11020 64 11060 104
rect 14380 2584 14420 2624
rect 15532 3760 15572 3800
rect 15916 6364 15956 6404
rect 15820 6280 15860 6320
rect 16492 6532 16532 6572
rect 16012 6196 16052 6236
rect 16108 5608 16148 5648
rect 16108 5356 16148 5396
rect 16012 5104 16052 5144
rect 15148 3508 15188 3548
rect 15628 3508 15668 3548
rect 15532 3424 15572 3464
rect 16396 6448 16436 6488
rect 16300 5692 16340 5732
rect 16972 10480 17012 10520
rect 17164 9892 17204 9932
rect 16876 9388 16916 9428
rect 16972 9220 17012 9260
rect 16780 8800 16820 8840
rect 16972 8380 17012 8420
rect 17356 8800 17396 8840
rect 17740 8800 17780 8840
rect 16876 7876 16916 7916
rect 17260 6952 17300 6992
rect 17260 5608 17300 5648
rect 16876 5188 16916 5228
rect 16876 4264 16916 4304
rect 15916 3256 15956 3296
rect 16204 3760 16244 3800
rect 15628 3088 15668 3128
rect 16012 3088 16052 3128
rect 15436 2920 15476 2960
rect 14380 2164 14420 2204
rect 16780 3508 16820 3548
rect 17836 8716 17876 8756
rect 17644 7960 17684 8000
rect 17740 7624 17780 7664
rect 17644 7120 17684 7160
rect 17740 6784 17780 6824
rect 17644 5860 17684 5900
rect 17644 5692 17684 5732
rect 17548 5608 17588 5648
rect 17740 5524 17780 5564
rect 17260 3928 17300 3968
rect 18124 8800 18164 8840
rect 18028 8632 18068 8672
rect 18220 8296 18260 8336
rect 18124 8128 18164 8168
rect 18028 7708 18068 7748
rect 18412 8800 18452 8840
rect 18700 10480 18740 10520
rect 18892 10312 18932 10352
rect 18892 9976 18932 10016
rect 18604 9472 18644 9512
rect 18508 8716 18548 8756
rect 18796 9388 18836 9428
rect 19180 9724 19220 9764
rect 18892 9304 18932 9344
rect 19180 9304 19220 9344
rect 18808 9052 18848 9092
rect 18890 9052 18930 9092
rect 18972 9052 19012 9092
rect 19054 9052 19094 9092
rect 19136 9052 19176 9092
rect 19372 9388 19412 9428
rect 18700 8800 18740 8840
rect 19276 8800 19316 8840
rect 19180 8716 19220 8756
rect 18604 7792 18644 7832
rect 19276 8548 19316 8588
rect 19564 8800 19604 8840
rect 18316 7456 18356 7496
rect 18316 6532 18356 6572
rect 18124 6112 18164 6152
rect 18124 5608 18164 5648
rect 18028 5524 18068 5564
rect 18796 7708 18836 7748
rect 18808 7540 18848 7580
rect 18890 7540 18930 7580
rect 18972 7540 19012 7580
rect 19054 7540 19094 7580
rect 19136 7540 19176 7580
rect 18892 6952 18932 6992
rect 19276 6952 19316 6992
rect 18988 6868 19028 6908
rect 18988 6616 19028 6656
rect 18892 6448 18932 6488
rect 19084 6280 19124 6320
rect 18808 6028 18848 6068
rect 18890 6028 18930 6068
rect 18972 6028 19012 6068
rect 19054 6028 19094 6068
rect 19136 6028 19176 6068
rect 18604 5692 18644 5732
rect 18508 5440 18548 5480
rect 18604 5272 18644 5312
rect 19084 5188 19124 5228
rect 19756 9976 19796 10016
rect 19660 7120 19700 7160
rect 20044 10396 20084 10436
rect 20620 10648 20660 10688
rect 20428 10228 20468 10268
rect 19948 9892 19988 9932
rect 20048 9808 20088 9848
rect 20130 9808 20170 9848
rect 20212 9808 20252 9848
rect 20294 9808 20334 9848
rect 20376 9808 20416 9848
rect 20140 8632 20180 8672
rect 20048 8296 20088 8336
rect 20130 8296 20170 8336
rect 20212 8296 20252 8336
rect 20294 8296 20334 8336
rect 20376 8296 20416 8336
rect 19852 6868 19892 6908
rect 20048 6784 20088 6824
rect 20130 6784 20170 6824
rect 20212 6784 20252 6824
rect 20294 6784 20334 6824
rect 20376 6784 20416 6824
rect 20908 10228 20948 10268
rect 21100 10228 21140 10268
rect 20812 8128 20852 8168
rect 20812 7960 20852 8000
rect 20716 7708 20756 7748
rect 21004 8632 21044 8672
rect 21196 8464 21236 8504
rect 21580 9472 21620 9512
rect 21484 8884 21524 8924
rect 21004 8128 21044 8168
rect 20908 7876 20948 7916
rect 20812 7540 20852 7580
rect 20620 6700 20660 6740
rect 19756 6616 19796 6656
rect 20332 6616 20372 6656
rect 19852 6532 19892 6572
rect 19372 6196 19412 6236
rect 19372 5944 19412 5984
rect 19276 4936 19316 4976
rect 18412 4768 18452 4808
rect 18808 4516 18848 4556
rect 18890 4516 18930 4556
rect 18972 4516 19012 4556
rect 19054 4516 19094 4556
rect 19136 4516 19176 4556
rect 19468 5356 19508 5396
rect 19372 4180 19412 4220
rect 19276 3760 19316 3800
rect 16588 3256 16628 3296
rect 16204 2836 16244 2876
rect 15436 2080 15476 2120
rect 15052 1996 15092 2036
rect 15052 1828 15092 1868
rect 14668 1072 14708 1112
rect 13612 904 13652 944
rect 14476 904 14516 944
rect 14668 904 14708 944
rect 13036 652 13076 692
rect 12844 64 12884 104
rect 13324 64 13364 104
rect 16684 3088 16724 3128
rect 18316 3424 18356 3464
rect 16684 1996 16724 2036
rect 16300 1912 16340 1952
rect 15628 1072 15668 1112
rect 16684 1744 16724 1784
rect 15340 64 15380 104
rect 15628 64 15668 104
rect 17548 1240 17588 1280
rect 18124 3340 18164 3380
rect 18316 3172 18356 3212
rect 18808 3004 18848 3044
rect 18890 3004 18930 3044
rect 18972 3004 19012 3044
rect 19054 3004 19094 3044
rect 19136 3004 19176 3044
rect 18028 2584 18068 2624
rect 18412 2584 18452 2624
rect 19948 5776 19988 5816
rect 20620 6280 20660 6320
rect 20332 5608 20372 5648
rect 19852 5524 19892 5564
rect 19948 5356 19988 5396
rect 20048 5272 20088 5312
rect 20130 5272 20170 5312
rect 20212 5272 20252 5312
rect 20294 5272 20334 5312
rect 20376 5272 20416 5312
rect 19564 4936 19604 4976
rect 19564 4516 19604 4556
rect 20332 4180 20372 4220
rect 19564 3760 19604 3800
rect 19948 4096 19988 4136
rect 20908 7120 20948 7160
rect 21676 8800 21716 8840
rect 21580 8632 21620 8672
rect 21580 7792 21620 7832
rect 21868 9304 21908 9344
rect 21772 8044 21812 8084
rect 21772 7876 21812 7916
rect 21676 7624 21716 7664
rect 21292 6616 21332 6656
rect 21196 6532 21236 6572
rect 20908 6112 20948 6152
rect 21484 6868 21524 6908
rect 21484 6616 21524 6656
rect 22252 9640 22292 9680
rect 21964 8884 22004 8924
rect 22156 8884 22196 8924
rect 22252 8800 22292 8840
rect 22828 10144 22868 10184
rect 22540 9556 22580 9596
rect 22732 9472 22772 9512
rect 22348 8716 22388 8756
rect 21868 7792 21908 7832
rect 21388 6112 21428 6152
rect 21100 6028 21140 6068
rect 20908 5440 20948 5480
rect 21100 4852 21140 4892
rect 20908 4768 20948 4808
rect 20048 3760 20088 3800
rect 20130 3760 20170 3800
rect 20212 3760 20252 3800
rect 20294 3760 20334 3800
rect 20376 3760 20416 3800
rect 19660 3340 19700 3380
rect 20044 3340 20084 3380
rect 19468 2752 19508 2792
rect 18808 1492 18848 1532
rect 18890 1492 18930 1532
rect 18972 1492 19012 1532
rect 19054 1492 19094 1532
rect 19136 1492 19176 1532
rect 20332 3172 20372 3212
rect 20044 2752 20084 2792
rect 17932 1240 17972 1280
rect 19084 1240 19124 1280
rect 19276 1240 19316 1280
rect 19660 1240 19700 1280
rect 20812 3592 20852 3632
rect 21292 5860 21332 5900
rect 21292 5188 21332 5228
rect 21676 5860 21716 5900
rect 21580 4852 21620 4892
rect 20908 3256 20948 3296
rect 20716 3088 20756 3128
rect 20524 2836 20564 2876
rect 20044 2500 20084 2540
rect 20048 2248 20088 2288
rect 20130 2248 20170 2288
rect 20212 2248 20252 2288
rect 20294 2248 20334 2288
rect 20376 2248 20416 2288
rect 20044 2080 20084 2120
rect 20140 2080 20180 2120
rect 20140 1828 20180 1868
rect 20044 1660 20084 1700
rect 17548 1072 17588 1112
rect 17932 1072 17972 1112
rect 17548 736 17588 776
rect 18412 820 18452 860
rect 19084 736 19124 776
rect 20048 736 20088 776
rect 20130 736 20170 776
rect 20212 736 20252 776
rect 20294 736 20334 776
rect 20376 736 20416 776
rect 18412 568 18452 608
rect 20236 64 20276 104
rect 20428 64 20468 104
rect 20812 3004 20852 3044
rect 20812 2752 20852 2792
rect 21292 2836 21332 2876
rect 21388 2752 21428 2792
rect 21196 2248 21236 2288
rect 21388 2248 21428 2288
rect 21292 1996 21332 2036
rect 21292 1240 21332 1280
rect 22540 8464 22580 8504
rect 23020 10144 23060 10184
rect 23212 10144 23252 10184
rect 23116 9976 23156 10016
rect 23020 9472 23060 9512
rect 22924 8716 22964 8756
rect 23020 8380 23060 8420
rect 22444 8044 22484 8084
rect 22060 7792 22100 7832
rect 22060 7540 22100 7580
rect 21964 6616 22004 6656
rect 22060 6532 22100 6572
rect 21964 6448 22004 6488
rect 22156 6448 22196 6488
rect 23788 9472 23828 9512
rect 23308 8212 23348 8252
rect 23212 8128 23252 8168
rect 22636 7120 22676 7160
rect 22540 6028 22580 6068
rect 22444 5860 22484 5900
rect 22444 5272 22484 5312
rect 22732 6028 22772 6068
rect 22444 4936 22484 4976
rect 22636 4936 22676 4976
rect 21868 4852 21908 4892
rect 22060 4852 22100 4892
rect 22060 4684 22100 4724
rect 21868 4264 21908 4304
rect 21772 4180 21812 4220
rect 22060 2920 22100 2960
rect 22540 2080 22580 2120
rect 23500 7456 23540 7496
rect 23692 8800 23732 8840
rect 23596 6532 23636 6572
rect 23116 6028 23156 6068
rect 23500 5608 23540 5648
rect 22924 5524 22964 5564
rect 22924 5356 22964 5396
rect 23116 5020 23156 5060
rect 23500 5020 23540 5060
rect 23308 4180 23348 4220
rect 23212 3424 23252 3464
rect 23308 3088 23348 3128
rect 23212 2836 23252 2876
rect 24076 10144 24116 10184
rect 23980 9556 24020 9596
rect 23884 9304 23924 9344
rect 23980 8884 24020 8924
rect 24172 9052 24212 9092
rect 23884 8716 23924 8756
rect 24268 8716 24308 8756
rect 24556 10060 24596 10100
rect 24460 8884 24500 8924
rect 24364 8044 24404 8084
rect 24076 7876 24116 7916
rect 24556 7456 24596 7496
rect 24364 7372 24404 7412
rect 24172 7120 24212 7160
rect 24076 6532 24116 6572
rect 23884 4852 23924 4892
rect 23884 4348 23924 4388
rect 23788 4180 23828 4220
rect 24076 5776 24116 5816
rect 23788 3508 23828 3548
rect 24460 6448 24500 6488
rect 24556 6280 24596 6320
rect 24364 5776 24404 5816
rect 23980 3424 24020 3464
rect 24364 5272 24404 5312
rect 24460 5188 24500 5228
rect 24460 4096 24500 4136
rect 23308 2752 23348 2792
rect 24172 2752 24212 2792
rect 23692 2584 23732 2624
rect 22828 2080 22868 2120
rect 21772 1744 21812 1784
rect 21676 1576 21716 1616
rect 21772 1408 21812 1448
rect 22540 1408 22580 1448
rect 21676 652 21716 692
rect 22924 1912 22964 1952
rect 24172 2080 24212 2120
rect 24844 6784 24884 6824
rect 25036 9724 25076 9764
rect 25132 7372 25172 7412
rect 25132 7120 25172 7160
rect 25036 5272 25076 5312
rect 25324 8296 25364 8336
rect 25708 9556 25748 9596
rect 25516 9136 25556 9176
rect 25612 8464 25652 8504
rect 25516 7540 25556 7580
rect 26092 8632 26132 8672
rect 26092 8464 26132 8504
rect 25708 7624 25748 7664
rect 25900 7960 25940 8000
rect 25804 7540 25844 7580
rect 25612 7120 25652 7160
rect 25516 6952 25556 6992
rect 25228 6616 25268 6656
rect 26284 9052 26324 9092
rect 26284 8800 26324 8840
rect 26476 8800 26516 8840
rect 26572 8716 26612 8756
rect 26476 8632 26516 8672
rect 26380 8380 26420 8420
rect 26284 7792 26324 7832
rect 26188 7540 26228 7580
rect 25804 6952 25844 6992
rect 25708 6616 25748 6656
rect 25516 5020 25556 5060
rect 24748 4012 24788 4052
rect 25132 4012 25172 4052
rect 24652 3004 24692 3044
rect 24460 2668 24500 2708
rect 24652 2584 24692 2624
rect 24556 2332 24596 2372
rect 24556 1912 24596 1952
rect 23788 1660 23828 1700
rect 23692 1240 23732 1280
rect 24940 3256 24980 3296
rect 24940 2920 24980 2960
rect 24940 2752 24980 2792
rect 24940 1912 24980 1952
rect 24844 1072 24884 1112
rect 25804 5608 25844 5648
rect 26188 6616 26228 6656
rect 26380 7624 26420 7664
rect 25996 6280 26036 6320
rect 26092 5944 26132 5984
rect 26956 10480 26996 10520
rect 26860 9556 26900 9596
rect 27052 9556 27092 9596
rect 26764 8716 26804 8756
rect 27148 8884 27188 8924
rect 26956 8800 26996 8840
rect 26860 8212 26900 8252
rect 26956 8128 26996 8168
rect 26860 7624 26900 7664
rect 26860 7288 26900 7328
rect 26668 6448 26708 6488
rect 27052 7624 27092 7664
rect 27340 9472 27380 9512
rect 27724 10564 27764 10604
rect 27340 9052 27380 9092
rect 27532 8800 27572 8840
rect 27340 8296 27380 8336
rect 27244 8212 27284 8252
rect 27532 8128 27572 8168
rect 27148 6700 27188 6740
rect 27244 6112 27284 6152
rect 26380 5440 26420 5480
rect 27052 5440 27092 5480
rect 26092 5020 26132 5060
rect 25996 3508 26036 3548
rect 25708 3424 25748 3464
rect 25900 3340 25940 3380
rect 25612 3172 25652 3212
rect 25612 2920 25652 2960
rect 25900 2668 25940 2708
rect 26572 4516 26612 4556
rect 26476 4096 26516 4136
rect 26476 3508 26516 3548
rect 27532 6700 27572 6740
rect 27724 8464 27764 8504
rect 27724 7120 27764 7160
rect 27916 8464 27956 8504
rect 28108 8128 28148 8168
rect 27820 5608 27860 5648
rect 28012 7960 28052 8000
rect 28204 7960 28244 8000
rect 28204 7708 28244 7748
rect 28396 9304 28436 9344
rect 28300 7624 28340 7664
rect 28012 6112 28052 6152
rect 28012 5944 28052 5984
rect 27916 5020 27956 5060
rect 27724 4936 27764 4976
rect 27628 4768 27668 4808
rect 28012 4012 28052 4052
rect 27532 3844 27572 3884
rect 27148 3508 27188 3548
rect 27436 3508 27476 3548
rect 27628 3424 27668 3464
rect 27244 3340 27284 3380
rect 26476 2080 26516 2120
rect 26188 1996 26228 2036
rect 25804 1912 25844 1952
rect 26668 1912 26708 1952
rect 26476 1744 26516 1784
rect 26476 1240 26516 1280
rect 25420 1156 25460 1196
rect 27532 2920 27572 2960
rect 27436 1912 27476 1952
rect 27916 2584 27956 2624
rect 28204 6532 28244 6572
rect 28684 8296 28724 8336
rect 29068 9136 29108 9176
rect 29356 9556 29396 9596
rect 28876 7456 28916 7496
rect 29164 8632 29204 8672
rect 29068 8464 29108 8504
rect 30412 9976 30452 10016
rect 30508 9808 30548 9848
rect 29644 9136 29684 9176
rect 29452 8800 29492 8840
rect 29548 8716 29588 8756
rect 29452 8464 29492 8504
rect 28972 7288 29012 7328
rect 29548 8128 29588 8168
rect 29356 7540 29396 7580
rect 29548 7540 29588 7580
rect 29260 7372 29300 7412
rect 28684 6952 28724 6992
rect 29164 6952 29204 6992
rect 28492 6364 28532 6404
rect 28972 6364 29012 6404
rect 28300 5440 28340 5480
rect 28300 5020 28340 5060
rect 28300 4516 28340 4556
rect 28396 4432 28436 4472
rect 28300 2584 28340 2624
rect 27532 1828 27572 1868
rect 27916 1828 27956 1868
rect 27628 1156 27668 1196
rect 25996 904 26036 944
rect 24844 484 24884 524
rect 27148 652 27188 692
rect 28108 1828 28148 1868
rect 28108 1576 28148 1616
rect 28012 736 28052 776
rect 27628 568 27668 608
rect 28684 3508 28724 3548
rect 28588 3424 28628 3464
rect 28588 2836 28628 2876
rect 28492 1912 28532 1952
rect 28780 3172 28820 3212
rect 29260 6448 29300 6488
rect 29452 6532 29492 6572
rect 28972 4348 29012 4388
rect 28972 3340 29012 3380
rect 28876 1912 28916 1952
rect 28876 1576 28916 1616
rect 29164 4348 29204 4388
rect 29356 3340 29396 3380
rect 29356 2416 29396 2456
rect 29164 1576 29204 1616
rect 29740 8464 29780 8504
rect 29740 7960 29780 8000
rect 29740 7624 29780 7664
rect 29644 6532 29684 6572
rect 29644 4936 29684 4976
rect 29740 4768 29780 4808
rect 29548 3508 29588 3548
rect 29644 2668 29684 2708
rect 29548 2164 29588 2204
rect 29548 1912 29588 1952
rect 30412 9472 30452 9512
rect 29932 8632 29972 8672
rect 30124 8632 30164 8672
rect 30028 8464 30068 8504
rect 29932 7540 29972 7580
rect 29932 5524 29972 5564
rect 30220 8128 30260 8168
rect 30220 7876 30260 7916
rect 30412 6028 30452 6068
rect 30796 9976 30836 10016
rect 31564 10480 31604 10520
rect 31852 10480 31892 10520
rect 31564 10228 31604 10268
rect 31372 9808 31412 9848
rect 30988 9640 31028 9680
rect 31468 9640 31508 9680
rect 30604 9052 30644 9092
rect 30604 8884 30644 8924
rect 30892 9472 30932 9512
rect 30998 9472 31038 9512
rect 31180 9472 31220 9512
rect 31180 9220 31220 9260
rect 30796 8548 30836 8588
rect 30796 7876 30836 7916
rect 31084 8884 31124 8924
rect 30988 8464 31028 8504
rect 30988 8128 31028 8168
rect 30220 5524 30260 5564
rect 30028 4600 30068 4640
rect 29932 3424 29972 3464
rect 30316 3760 30356 3800
rect 30220 3424 30260 3464
rect 30604 5524 30644 5564
rect 30892 7456 30932 7496
rect 30988 7120 31028 7160
rect 31372 8464 31412 8504
rect 31372 7708 31412 7748
rect 31564 9052 31604 9092
rect 31564 8128 31604 8168
rect 31564 7876 31604 7916
rect 30796 6280 30836 6320
rect 30988 6028 31028 6068
rect 30892 4852 30932 4892
rect 30892 4600 30932 4640
rect 30604 4096 30644 4136
rect 30604 3592 30644 3632
rect 30892 4096 30932 4136
rect 30988 3928 31028 3968
rect 31756 8464 31796 8504
rect 31756 8128 31796 8168
rect 31660 7204 31700 7244
rect 31564 7120 31604 7160
rect 31564 6784 31604 6824
rect 31468 6280 31508 6320
rect 30508 3256 30548 3296
rect 30988 3256 31028 3296
rect 31372 2836 31412 2876
rect 31660 5944 31700 5984
rect 31948 7456 31988 7496
rect 31948 7288 31988 7328
rect 32236 10312 32276 10352
rect 32332 9724 32372 9764
rect 32428 9640 32468 9680
rect 32428 9220 32468 9260
rect 32428 9052 32468 9092
rect 32812 10144 32852 10184
rect 32716 9724 32756 9764
rect 32620 9556 32660 9596
rect 32620 9220 32660 9260
rect 32428 7624 32468 7664
rect 32620 7708 32660 7748
rect 32524 7372 32564 7412
rect 31948 6448 31988 6488
rect 32044 6364 32084 6404
rect 31756 5524 31796 5564
rect 31660 5440 31700 5480
rect 31564 4348 31604 4388
rect 31564 3760 31604 3800
rect 31852 4516 31892 4556
rect 31852 3928 31892 3968
rect 31756 2584 31796 2624
rect 31180 2080 31220 2120
rect 32140 5524 32180 5564
rect 32044 4936 32084 4976
rect 32044 4348 32084 4388
rect 31948 3760 31988 3800
rect 30892 1912 30932 1952
rect 30796 1576 30836 1616
rect 30124 1240 30164 1280
rect 31372 1660 31412 1700
rect 31180 1072 31220 1112
rect 28588 904 28628 944
rect 31468 904 31508 944
rect 29452 736 29492 776
rect 30604 568 30644 608
rect 31660 1240 31700 1280
rect 31756 1156 31796 1196
rect 31564 484 31604 524
rect 32236 4936 32276 4976
rect 32236 4684 32276 4724
rect 32236 4432 32276 4472
rect 32236 3424 32276 3464
rect 32908 9388 32948 9428
rect 32908 9220 32948 9260
rect 32908 8548 32948 8588
rect 41452 10480 41492 10520
rect 34732 10396 34772 10436
rect 34156 9640 34196 9680
rect 33484 9388 33524 9428
rect 33928 9052 33968 9092
rect 34010 9052 34050 9092
rect 34092 9052 34132 9092
rect 34174 9052 34214 9092
rect 34256 9052 34296 9092
rect 33100 8716 33140 8756
rect 33004 8380 33044 8420
rect 33100 8296 33140 8336
rect 32908 8212 32948 8252
rect 33484 8212 33524 8252
rect 32812 8128 32852 8168
rect 34348 8800 34388 8840
rect 33868 8716 33908 8756
rect 34444 8716 34484 8756
rect 33292 7960 33332 8000
rect 32908 7624 32948 7664
rect 32812 7204 32852 7244
rect 32716 5524 32756 5564
rect 33004 7120 33044 7160
rect 33004 6616 33044 6656
rect 33292 7708 33332 7748
rect 33196 7120 33236 7160
rect 35168 9808 35208 9848
rect 35250 9808 35290 9848
rect 35332 9808 35372 9848
rect 35414 9808 35454 9848
rect 35496 9808 35536 9848
rect 40300 9808 40340 9848
rect 37132 9556 37172 9596
rect 35020 9220 35060 9260
rect 36076 9052 36116 9092
rect 36268 9052 36308 9092
rect 34732 8800 34772 8840
rect 35788 8800 35828 8840
rect 34636 8632 34676 8672
rect 35596 8716 35636 8756
rect 35168 8296 35208 8336
rect 35250 8296 35290 8336
rect 35332 8296 35372 8336
rect 35414 8296 35454 8336
rect 35496 8296 35536 8336
rect 33928 7540 33968 7580
rect 34010 7540 34050 7580
rect 34092 7540 34132 7580
rect 34174 7540 34214 7580
rect 34256 7540 34296 7580
rect 33676 6952 33716 6992
rect 33676 6616 33716 6656
rect 33388 6448 33428 6488
rect 32620 5020 32660 5060
rect 32524 4096 32564 4136
rect 32524 3760 32564 3800
rect 32812 3592 32852 3632
rect 32716 3508 32756 3548
rect 32620 2836 32660 2876
rect 32908 2836 32948 2876
rect 32332 1240 32372 1280
rect 32332 904 32372 944
rect 32140 820 32180 860
rect 33100 5272 33140 5312
rect 33196 4768 33236 4808
rect 33292 4516 33332 4556
rect 33196 4096 33236 4136
rect 33100 3676 33140 3716
rect 34540 6868 34580 6908
rect 34444 6448 34484 6488
rect 34348 6196 34388 6236
rect 33928 6028 33968 6068
rect 34010 6028 34050 6068
rect 34092 6028 34132 6068
rect 34174 6028 34214 6068
rect 34256 6028 34296 6068
rect 34444 5776 34484 5816
rect 33772 5104 33812 5144
rect 35168 6784 35208 6824
rect 35250 6784 35290 6824
rect 35332 6784 35372 6824
rect 35414 6784 35454 6824
rect 35496 6784 35536 6824
rect 36364 8800 36404 8840
rect 36268 8716 36308 8756
rect 36172 8464 36212 8504
rect 37036 8968 37076 9008
rect 36556 7792 36596 7832
rect 36556 7624 36596 7664
rect 36076 7120 36116 7160
rect 36268 6868 36308 6908
rect 34636 6448 34676 6488
rect 34828 6196 34868 6236
rect 34828 5944 34868 5984
rect 35596 6448 35636 6488
rect 35404 5776 35444 5816
rect 34924 5608 34964 5648
rect 35168 5272 35208 5312
rect 35250 5272 35290 5312
rect 35332 5272 35372 5312
rect 35414 5272 35454 5312
rect 35496 5272 35536 5312
rect 35692 6280 35732 6320
rect 36556 6364 36596 6404
rect 36268 5944 36308 5984
rect 33928 4516 33968 4556
rect 34010 4516 34050 4556
rect 34092 4516 34132 4556
rect 34174 4516 34214 4556
rect 34256 4516 34296 4556
rect 34156 3928 34196 3968
rect 33772 3592 33812 3632
rect 33676 3424 33716 3464
rect 33676 3256 33716 3296
rect 33292 2584 33332 2624
rect 33928 3004 33968 3044
rect 34010 3004 34050 3044
rect 34092 3004 34132 3044
rect 34174 3004 34214 3044
rect 34256 3004 34296 3044
rect 35500 4096 35540 4136
rect 35596 3844 35636 3884
rect 35168 3760 35208 3800
rect 35250 3760 35290 3800
rect 35332 3760 35372 3800
rect 35414 3760 35454 3800
rect 35496 3760 35536 3800
rect 35884 4096 35924 4136
rect 35788 3676 35828 3716
rect 35596 3592 35636 3632
rect 35020 3508 35060 3548
rect 35404 3508 35444 3548
rect 34924 2584 34964 2624
rect 34828 2416 34868 2456
rect 34636 1996 34676 2036
rect 33388 1912 33428 1952
rect 33928 1492 33968 1532
rect 34010 1492 34050 1532
rect 34092 1492 34132 1532
rect 34174 1492 34214 1532
rect 34256 1492 34296 1532
rect 35980 3424 36020 3464
rect 36556 5692 36596 5732
rect 36460 5608 36500 5648
rect 36844 5944 36884 5984
rect 36748 5524 36788 5564
rect 36940 5524 36980 5564
rect 37612 9220 37652 9260
rect 37804 8884 37844 8924
rect 37324 7960 37364 8000
rect 39724 9472 39764 9512
rect 38860 9304 38900 9344
rect 38476 8884 38516 8924
rect 38668 8464 38708 8504
rect 38572 8212 38612 8252
rect 37612 7960 37652 8000
rect 38284 7960 38324 8000
rect 37516 7120 37556 7160
rect 37420 6028 37460 6068
rect 37420 5776 37460 5816
rect 37228 4936 37268 4976
rect 36652 4768 36692 4808
rect 35308 2416 35348 2456
rect 35168 2248 35208 2288
rect 35250 2248 35290 2288
rect 35332 2248 35372 2288
rect 35414 2248 35454 2288
rect 35496 2248 35536 2288
rect 36844 3928 36884 3968
rect 36652 3760 36692 3800
rect 36556 2836 36596 2876
rect 37324 4096 37364 4136
rect 37228 4012 37268 4052
rect 36940 2836 36980 2876
rect 36748 2584 36788 2624
rect 36268 1744 36308 1784
rect 33484 1240 33524 1280
rect 35596 1240 35636 1280
rect 32620 820 32660 860
rect 32812 736 32852 776
rect 32524 652 32564 692
rect 32908 652 32948 692
rect 33676 1156 33716 1196
rect 34156 820 34196 860
rect 34636 904 34676 944
rect 34444 652 34484 692
rect 33292 568 33332 608
rect 34060 568 34100 608
rect 34828 568 34868 608
rect 36364 1156 36404 1196
rect 35020 904 35060 944
rect 35168 736 35208 776
rect 35250 736 35290 776
rect 35332 736 35372 776
rect 35414 736 35454 776
rect 35496 736 35536 776
rect 34924 64 34964 104
rect 35212 64 35252 104
rect 37612 6616 37652 6656
rect 38380 6448 38420 6488
rect 41548 10144 41588 10184
rect 40492 9472 40532 9512
rect 41068 9472 41108 9512
rect 39148 8716 39188 8756
rect 38956 8380 38996 8420
rect 38572 6448 38612 6488
rect 39724 8464 39764 8504
rect 39340 7792 39380 7832
rect 39148 7288 39188 7328
rect 38284 5020 38324 5060
rect 37516 3760 37556 3800
rect 38476 4768 38516 4808
rect 37900 4096 37940 4136
rect 38092 4096 38132 4136
rect 38860 6448 38900 6488
rect 39820 7540 39860 7580
rect 40588 9388 40628 9428
rect 40876 9388 40916 9428
rect 40492 8128 40532 8168
rect 40396 7540 40436 7580
rect 38764 6028 38804 6068
rect 39820 6280 39860 6320
rect 38956 5608 38996 5648
rect 38956 5440 38996 5480
rect 38668 5020 38708 5060
rect 38668 4768 38708 4808
rect 38860 4684 38900 4724
rect 39244 5104 39284 5144
rect 39052 4768 39092 4808
rect 38380 3760 38420 3800
rect 38668 3760 38708 3800
rect 38284 3676 38324 3716
rect 37804 2836 37844 2876
rect 38764 3340 38804 3380
rect 38572 2836 38612 2876
rect 37132 2164 37172 2204
rect 37132 1912 37172 1952
rect 39628 4852 39668 4892
rect 39436 4684 39476 4724
rect 37612 1408 37652 1448
rect 37420 1156 37460 1196
rect 38188 1660 38228 1700
rect 37900 1072 37940 1112
rect 37516 64 37556 104
rect 37804 64 37844 104
rect 39628 1744 39668 1784
rect 39820 1408 39860 1448
rect 40012 6364 40052 6404
rect 40396 6364 40436 6404
rect 40204 6280 40244 6320
rect 40300 6196 40340 6236
rect 40108 4768 40148 4808
rect 40492 4684 40532 4724
rect 40492 4432 40532 4472
rect 40300 3592 40340 3632
rect 40492 3340 40532 3380
rect 40492 2248 40532 2288
rect 41260 9304 41300 9344
rect 41260 9136 41300 9176
rect 40684 8884 40724 8924
rect 40876 8716 40916 8756
rect 41452 9052 41492 9092
rect 41068 8464 41108 8504
rect 41260 8380 41300 8420
rect 40684 8128 40724 8168
rect 40876 7204 40916 7244
rect 40876 6952 40916 6992
rect 40780 5860 40820 5900
rect 40684 4852 40724 4892
rect 40684 4432 40724 4472
rect 40876 5692 40916 5732
rect 40876 5356 40916 5396
rect 41068 7792 41108 7832
rect 41356 7708 41396 7748
rect 41068 7120 41108 7160
rect 41068 6448 41108 6488
rect 41068 6112 41108 6152
rect 41260 6364 41300 6404
rect 41164 5608 41204 5648
rect 41068 5440 41108 5480
rect 40972 4936 41012 4976
rect 41260 5188 41300 5228
rect 41452 7456 41492 7496
rect 41452 6784 41492 6824
rect 41452 5776 41492 5816
rect 41452 5104 41492 5144
rect 41164 4768 41204 4808
rect 41260 4600 41300 4640
rect 41452 4096 41492 4136
rect 41068 3760 41108 3800
rect 40876 3592 40916 3632
rect 40684 3424 40724 3464
rect 41068 3088 41108 3128
rect 41260 2920 41300 2960
rect 40684 2752 40724 2792
rect 40780 2500 40820 2540
rect 40492 1912 40532 1952
rect 40012 1828 40052 1868
rect 39916 904 39956 944
rect 41452 2416 41492 2456
rect 40876 2332 40916 2372
rect 41068 2080 41108 2120
rect 40204 400 40244 440
rect 39628 64 39668 104
rect 39820 64 39860 104
rect 41452 1744 41492 1784
rect 41164 1240 41204 1280
rect 40876 1156 40916 1196
rect 40684 1072 40724 1112
rect 41260 988 41300 1028
rect 41452 736 41492 776
rect 41068 148 41108 188
rect 40780 64 40820 104
rect 40972 64 41012 104
<< metal3 >>
rect 20611 10688 20669 10689
rect 8899 10648 8908 10688
rect 8948 10648 9484 10688
rect 9524 10648 9533 10688
rect 20526 10648 20620 10688
rect 20660 10648 20669 10688
rect 20611 10647 20669 10648
rect 11107 10564 11116 10604
rect 11156 10564 27724 10604
rect 27764 10564 27773 10604
rect 0 10520 80 10540
rect 4579 10520 4637 10521
rect 16963 10520 17021 10521
rect 18691 10520 18749 10521
rect 42928 10520 43008 10540
rect 0 10480 4588 10520
rect 4628 10480 4637 10520
rect 16878 10480 16972 10520
rect 17012 10480 17021 10520
rect 18606 10480 18700 10520
rect 18740 10480 18749 10520
rect 0 10460 80 10480
rect 4579 10479 4637 10480
rect 16963 10479 17021 10480
rect 18691 10479 18749 10480
rect 18796 10480 26956 10520
rect 26996 10480 27005 10520
rect 31555 10480 31564 10520
rect 31604 10480 31852 10520
rect 31892 10480 31901 10520
rect 41443 10480 41452 10520
rect 41492 10480 43008 10520
rect 18796 10436 18836 10480
rect 42928 10460 43008 10480
rect 11491 10396 11500 10436
rect 11540 10396 18836 10436
rect 20035 10396 20044 10436
rect 20084 10396 34732 10436
rect 34772 10396 34781 10436
rect 18883 10312 18892 10352
rect 18932 10312 32236 10352
rect 32276 10312 32285 10352
rect 21091 10268 21149 10269
rect 20419 10228 20428 10268
rect 20468 10228 20908 10268
rect 20948 10228 20957 10268
rect 21091 10228 21100 10268
rect 21140 10228 31564 10268
rect 31604 10228 31613 10268
rect 21091 10227 21149 10228
rect 0 10184 80 10204
rect 42928 10184 43008 10204
rect 0 10144 2764 10184
rect 2804 10144 2813 10184
rect 13123 10144 13132 10184
rect 13172 10144 22828 10184
rect 22868 10144 22877 10184
rect 23011 10144 23020 10184
rect 23060 10144 23212 10184
rect 23252 10144 23261 10184
rect 24067 10144 24076 10184
rect 24116 10144 32812 10184
rect 32852 10144 32861 10184
rect 41539 10144 41548 10184
rect 41588 10144 43008 10184
rect 0 10124 80 10144
rect 42928 10124 43008 10144
rect 15811 10060 15820 10100
rect 15860 10060 24556 10100
rect 24596 10060 24605 10100
rect 16387 10016 16445 10017
rect 10531 9976 10540 10016
rect 10580 9976 16396 10016
rect 16436 9976 16445 10016
rect 18883 9976 18892 10016
rect 18932 9976 19756 10016
rect 19796 9976 23116 10016
rect 23156 9976 23165 10016
rect 30403 9976 30412 10016
rect 30452 9976 30796 10016
rect 30836 9976 30845 10016
rect 16387 9975 16445 9976
rect 1891 9892 1900 9932
rect 1940 9892 2540 9932
rect 17155 9892 17164 9932
rect 17204 9892 19948 9932
rect 19988 9892 19997 9932
rect 0 9848 80 9868
rect 1603 9848 1661 9849
rect 0 9808 1612 9848
rect 1652 9808 1661 9848
rect 0 9788 80 9808
rect 1603 9807 1661 9808
rect 2500 9764 2540 9892
rect 42928 9848 43008 9868
rect 4919 9808 4928 9848
rect 4968 9808 5010 9848
rect 5050 9808 5092 9848
rect 5132 9808 5174 9848
rect 5214 9808 5256 9848
rect 5296 9808 5305 9848
rect 9667 9808 9676 9848
rect 9716 9808 10156 9848
rect 10196 9808 10205 9848
rect 16195 9808 16204 9848
rect 16244 9808 19316 9848
rect 20039 9808 20048 9848
rect 20088 9808 20130 9848
rect 20170 9808 20212 9848
rect 20252 9808 20294 9848
rect 20334 9808 20376 9848
rect 20416 9808 20425 9848
rect 30499 9808 30508 9848
rect 30548 9808 31372 9848
rect 31412 9808 31421 9848
rect 35159 9808 35168 9848
rect 35208 9808 35250 9848
rect 35290 9808 35332 9848
rect 35372 9808 35414 9848
rect 35454 9808 35496 9848
rect 35536 9808 35545 9848
rect 40291 9808 40300 9848
rect 40340 9808 43008 9848
rect 19276 9764 19316 9808
rect 42928 9788 43008 9808
rect 2500 9724 19180 9764
rect 19220 9724 19229 9764
rect 19276 9724 25036 9764
rect 25076 9724 25085 9764
rect 32323 9724 32332 9764
rect 32372 9724 32716 9764
rect 32756 9724 32765 9764
rect 12643 9680 12701 9681
rect 15235 9680 15293 9681
rect 3715 9640 3724 9680
rect 3764 9640 5740 9680
rect 5780 9640 5789 9680
rect 12163 9640 12172 9680
rect 12212 9640 12652 9680
rect 12692 9640 12701 9680
rect 13891 9640 13900 9680
rect 13940 9640 14188 9680
rect 14228 9640 14237 9680
rect 15150 9640 15244 9680
rect 15284 9640 15293 9680
rect 16387 9640 16396 9680
rect 16436 9640 22252 9680
rect 22292 9640 22301 9680
rect 30979 9640 30988 9680
rect 31028 9640 31468 9680
rect 31508 9640 31517 9680
rect 32419 9640 32428 9680
rect 32468 9640 34156 9680
rect 34196 9640 34205 9680
rect 12643 9639 12701 9640
rect 15235 9639 15293 9640
rect 16387 9596 16445 9597
rect 22627 9596 22685 9597
rect 32428 9596 32468 9640
rect 3523 9556 3532 9596
rect 3572 9556 5356 9596
rect 5396 9556 5405 9596
rect 5452 9556 5932 9596
rect 5972 9556 11360 9596
rect 14851 9556 14860 9596
rect 14900 9556 16396 9596
rect 16436 9556 16445 9596
rect 22531 9556 22540 9596
rect 22580 9556 22636 9596
rect 22676 9556 22685 9596
rect 23971 9556 23980 9596
rect 24020 9556 25708 9596
rect 25748 9556 26860 9596
rect 26900 9556 27052 9596
rect 27092 9556 29356 9596
rect 29396 9556 32468 9596
rect 32611 9556 32620 9596
rect 32660 9556 37132 9596
rect 37172 9556 37181 9596
rect 0 9512 80 9532
rect 5452 9513 5492 9556
rect 5443 9512 5501 9513
rect 0 9472 3436 9512
rect 3476 9472 3485 9512
rect 3811 9472 3820 9512
rect 3860 9472 4396 9512
rect 4436 9472 4445 9512
rect 5443 9472 5452 9512
rect 5492 9472 5501 9512
rect 6979 9472 6988 9512
rect 7028 9472 7852 9512
rect 7892 9472 7901 9512
rect 0 9452 80 9472
rect 5443 9471 5501 9472
rect 7555 9428 7613 9429
rect 10339 9428 10397 9429
rect 3331 9388 3340 9428
rect 3380 9388 3628 9428
rect 3668 9388 4492 9428
rect 4532 9388 7180 9428
rect 7220 9388 7229 9428
rect 7470 9388 7564 9428
rect 7604 9388 7613 9428
rect 10254 9388 10348 9428
rect 10388 9388 10397 9428
rect 7555 9387 7613 9388
rect 10339 9387 10397 9388
rect 11320 9344 11360 9556
rect 16387 9555 16445 9556
rect 22627 9555 22685 9556
rect 22819 9512 22877 9513
rect 31084 9512 31124 9556
rect 42928 9512 43008 9532
rect 13123 9472 13132 9512
rect 13172 9472 14956 9512
rect 14996 9472 15005 9512
rect 18595 9472 18604 9512
rect 18644 9472 21580 9512
rect 21620 9472 21629 9512
rect 22723 9472 22732 9512
rect 22772 9472 22828 9512
rect 22868 9472 22877 9512
rect 23011 9472 23020 9512
rect 23060 9472 23788 9512
rect 23828 9472 27340 9512
rect 27380 9472 27389 9512
rect 30403 9472 30412 9512
rect 30452 9472 30892 9512
rect 30932 9472 30941 9512
rect 30989 9472 30998 9512
rect 31038 9472 31124 9512
rect 31171 9472 31180 9512
rect 31220 9472 39724 9512
rect 39764 9472 40492 9512
rect 40532 9472 40541 9512
rect 41059 9472 41068 9512
rect 41108 9472 43008 9512
rect 22819 9471 22877 9472
rect 42928 9452 43008 9472
rect 40867 9428 40925 9429
rect 16483 9388 16492 9428
rect 16532 9388 16876 9428
rect 16916 9388 16925 9428
rect 18787 9388 18796 9428
rect 18836 9388 19372 9428
rect 19412 9388 19421 9428
rect 20140 9388 32908 9428
rect 32948 9388 32957 9428
rect 33475 9388 33484 9428
rect 33524 9388 40588 9428
rect 40628 9388 40637 9428
rect 40782 9388 40876 9428
rect 40916 9388 40925 9428
rect 20140 9344 20180 9388
rect 40867 9387 40925 9388
rect 3523 9304 3532 9344
rect 3572 9304 4876 9344
rect 4916 9304 5836 9344
rect 5876 9304 7468 9344
rect 7508 9304 7517 9344
rect 11320 9304 18892 9344
rect 18932 9304 18941 9344
rect 19171 9304 19180 9344
rect 19220 9304 20180 9344
rect 21859 9304 21868 9344
rect 21908 9304 23884 9344
rect 23924 9304 23933 9344
rect 28387 9304 28396 9344
rect 28436 9304 38860 9344
rect 38900 9304 41260 9344
rect 41300 9304 41309 9344
rect 37603 9260 37661 9261
rect 16963 9220 16972 9260
rect 17012 9220 31180 9260
rect 31220 9220 31229 9260
rect 32419 9220 32428 9260
rect 32468 9220 32620 9260
rect 32660 9220 32669 9260
rect 32899 9220 32908 9260
rect 32948 9220 35020 9260
rect 35060 9220 35069 9260
rect 37518 9220 37612 9260
rect 37652 9220 37661 9260
rect 0 9176 80 9196
rect 14179 9176 14237 9177
rect 35020 9176 35060 9220
rect 37603 9219 37661 9220
rect 42928 9176 43008 9196
rect 0 9136 1900 9176
rect 1940 9136 1949 9176
rect 10051 9136 10060 9176
rect 10100 9136 10540 9176
rect 10580 9136 10589 9176
rect 12931 9136 12940 9176
rect 12980 9136 14188 9176
rect 14228 9136 14237 9176
rect 15043 9136 15052 9176
rect 15092 9136 25516 9176
rect 25556 9136 25565 9176
rect 29059 9136 29068 9176
rect 29108 9136 29644 9176
rect 29684 9136 29693 9176
rect 30604 9136 34964 9176
rect 35020 9136 41260 9176
rect 41300 9136 41309 9176
rect 41452 9136 43008 9176
rect 0 9116 80 9136
rect 14179 9135 14237 9136
rect 22723 9092 22781 9093
rect 26275 9092 26333 9093
rect 30604 9092 30644 9136
rect 34924 9092 34964 9136
rect 41452 9092 41492 9136
rect 42928 9116 43008 9136
rect 3679 9052 3688 9092
rect 3728 9052 3770 9092
rect 3810 9052 3852 9092
rect 3892 9052 3934 9092
rect 3974 9052 4016 9092
rect 4056 9052 4065 9092
rect 8803 9052 8812 9092
rect 8852 9052 9964 9092
rect 10004 9052 11252 9092
rect 11395 9052 11404 9092
rect 11444 9052 11692 9092
rect 11732 9052 11741 9092
rect 13315 9052 13324 9092
rect 13364 9052 14420 9092
rect 18799 9052 18808 9092
rect 18848 9052 18890 9092
rect 18930 9052 18972 9092
rect 19012 9052 19054 9092
rect 19094 9052 19136 9092
rect 19176 9052 19185 9092
rect 22723 9052 22732 9092
rect 22772 9052 24172 9092
rect 24212 9052 24221 9092
rect 26190 9052 26284 9092
rect 26324 9052 26333 9092
rect 27331 9052 27340 9092
rect 27380 9052 30604 9092
rect 30644 9052 30653 9092
rect 31555 9052 31564 9092
rect 31604 9052 32428 9092
rect 32468 9052 32477 9092
rect 33919 9052 33928 9092
rect 33968 9052 34010 9092
rect 34050 9052 34092 9092
rect 34132 9052 34174 9092
rect 34214 9052 34256 9092
rect 34296 9052 34305 9092
rect 34924 9052 36076 9092
rect 36116 9052 36268 9092
rect 36308 9052 37820 9092
rect 41443 9052 41452 9092
rect 41492 9052 41501 9092
rect 11212 9008 11252 9052
rect 14380 9008 14420 9052
rect 22723 9051 22781 9052
rect 26275 9051 26333 9052
rect 1795 8968 1804 9008
rect 1844 8968 2540 9008
rect 5155 8968 5164 9008
rect 5204 8968 5452 9008
rect 5492 8968 5501 9008
rect 10339 8968 10348 9008
rect 10388 8968 11116 9008
rect 11156 8968 11165 9008
rect 11212 8968 12172 9008
rect 12212 8968 12221 9008
rect 12931 8968 12940 9008
rect 12980 8968 14284 9008
rect 14324 8968 14333 9008
rect 14380 8968 37036 9008
rect 37076 8968 37085 9008
rect 2500 8924 2540 8968
rect 37780 8924 37820 9052
rect 2500 8884 21484 8924
rect 21524 8884 21533 8924
rect 21955 8884 21964 8924
rect 22004 8884 22013 8924
rect 22147 8884 22156 8924
rect 22196 8884 23980 8924
rect 24020 8884 24029 8924
rect 24451 8884 24460 8924
rect 24500 8884 27148 8924
rect 27188 8884 27197 8924
rect 30595 8884 30604 8924
rect 30644 8884 31084 8924
rect 31124 8884 31133 8924
rect 31660 8884 32660 8924
rect 0 8840 80 8860
rect 10243 8840 10301 8841
rect 11011 8840 11069 8841
rect 11779 8840 11837 8841
rect 12547 8840 12605 8841
rect 14083 8840 14141 8841
rect 14467 8840 14525 8841
rect 15427 8840 15485 8841
rect 15619 8840 15677 8841
rect 16003 8840 16061 8841
rect 16771 8840 16829 8841
rect 18115 8840 18173 8841
rect 21964 8840 22004 8884
rect 22243 8840 22301 8841
rect 31660 8840 31700 8884
rect 0 8800 1844 8840
rect 1891 8800 1900 8840
rect 1940 8800 4684 8840
rect 4724 8800 4733 8840
rect 5539 8800 5548 8840
rect 5588 8800 6604 8840
rect 6644 8800 6653 8840
rect 6883 8800 6892 8840
rect 6932 8800 7564 8840
rect 7604 8800 7613 8840
rect 10158 8800 10252 8840
rect 10292 8800 10301 8840
rect 10926 8800 11020 8840
rect 11060 8800 11069 8840
rect 11203 8800 11212 8840
rect 11252 8800 11540 8840
rect 11694 8800 11788 8840
rect 11828 8800 11837 8840
rect 12462 8800 12556 8840
rect 12596 8800 12605 8840
rect 13998 8800 14092 8840
rect 14132 8800 14141 8840
rect 14382 8800 14476 8840
rect 14516 8800 14525 8840
rect 15342 8800 15436 8840
rect 15476 8800 15485 8840
rect 15534 8800 15628 8840
rect 15668 8800 15677 8840
rect 15918 8800 16012 8840
rect 16052 8800 16061 8840
rect 16686 8800 16780 8840
rect 16820 8800 16829 8840
rect 17347 8800 17356 8840
rect 17396 8800 17740 8840
rect 17780 8800 17789 8840
rect 18030 8800 18124 8840
rect 18164 8800 18173 8840
rect 18403 8800 18412 8840
rect 18452 8800 18700 8840
rect 18740 8800 18749 8840
rect 19267 8800 19276 8840
rect 19316 8800 19564 8840
rect 19604 8800 19613 8840
rect 21667 8800 21676 8840
rect 21716 8800 22004 8840
rect 22158 8800 22252 8840
rect 22292 8800 22301 8840
rect 23683 8800 23692 8840
rect 23732 8800 26284 8840
rect 26324 8800 26476 8840
rect 26516 8800 26525 8840
rect 26947 8800 26956 8840
rect 26996 8800 27532 8840
rect 27572 8800 27581 8840
rect 29443 8800 29452 8840
rect 29492 8800 31700 8840
rect 32620 8840 32660 8884
rect 33676 8884 34484 8924
rect 37780 8884 37804 8924
rect 37844 8884 38476 8924
rect 38516 8884 38525 8924
rect 40675 8884 40684 8924
rect 40724 8884 41600 8924
rect 33676 8840 33716 8884
rect 32620 8800 33716 8840
rect 33763 8840 33821 8841
rect 34444 8840 34484 8884
rect 41560 8840 41600 8884
rect 42928 8840 43008 8860
rect 33763 8800 33772 8840
rect 33812 8800 34348 8840
rect 34388 8800 34397 8840
rect 34444 8800 34676 8840
rect 34723 8800 34732 8840
rect 34772 8800 35788 8840
rect 35828 8800 36364 8840
rect 36404 8800 36413 8840
rect 41560 8800 43008 8840
rect 0 8780 80 8800
rect 1804 8756 1844 8800
rect 10243 8799 10301 8800
rect 11011 8799 11069 8800
rect 11395 8756 11453 8757
rect 1804 8716 2092 8756
rect 2132 8716 2141 8756
rect 8419 8716 8428 8756
rect 8468 8716 9196 8756
rect 9236 8716 9245 8756
rect 10627 8716 10636 8756
rect 10676 8716 11404 8756
rect 11444 8716 11453 8756
rect 11395 8715 11453 8716
rect 10243 8674 10252 8714
rect 10292 8674 10388 8714
rect 3715 8672 3773 8673
rect 8803 8672 8861 8673
rect 9763 8672 9821 8673
rect 3630 8632 3724 8672
rect 3764 8632 3773 8672
rect 4195 8632 4204 8672
rect 4244 8632 5396 8672
rect 5923 8632 5932 8672
rect 5972 8632 6124 8672
rect 6164 8632 6173 8672
rect 6691 8632 6700 8672
rect 6740 8632 7372 8672
rect 7412 8632 7421 8672
rect 8718 8632 8812 8672
rect 8852 8632 9772 8672
rect 9812 8632 9821 8672
rect 10348 8672 10388 8674
rect 11500 8672 11540 8800
rect 11779 8799 11837 8800
rect 12547 8799 12605 8800
rect 14083 8799 14141 8800
rect 14467 8799 14525 8800
rect 15427 8799 15485 8800
rect 15619 8799 15677 8800
rect 16003 8799 16061 8800
rect 16771 8799 16829 8800
rect 18115 8799 18173 8800
rect 22243 8799 22301 8800
rect 33763 8799 33821 8800
rect 33187 8756 33245 8757
rect 34636 8756 34676 8800
rect 42928 8780 43008 8800
rect 17827 8716 17836 8756
rect 17876 8716 18508 8756
rect 18548 8716 18557 8756
rect 19171 8716 19180 8756
rect 19220 8716 22348 8756
rect 22388 8716 22397 8756
rect 22915 8716 22924 8756
rect 22964 8716 23884 8756
rect 23924 8716 24268 8756
rect 24308 8716 24317 8756
rect 26563 8716 26572 8756
rect 26612 8716 26764 8756
rect 26804 8716 29548 8756
rect 29588 8716 29597 8756
rect 33091 8716 33100 8756
rect 33140 8716 33196 8756
rect 33236 8716 33245 8756
rect 33859 8716 33868 8756
rect 33908 8716 34444 8756
rect 34484 8716 34493 8756
rect 34636 8716 35596 8756
rect 35636 8716 36268 8756
rect 36308 8716 36317 8756
rect 39139 8716 39148 8756
rect 39188 8716 40876 8756
rect 40916 8716 40925 8756
rect 13027 8672 13085 8673
rect 14851 8672 14909 8673
rect 15811 8672 15869 8673
rect 19459 8672 19517 8673
rect 22924 8672 22964 8716
rect 33187 8715 33245 8716
rect 10348 8632 10828 8672
rect 10868 8632 10877 8672
rect 11491 8632 11500 8672
rect 11540 8632 11549 8672
rect 11875 8632 11884 8672
rect 11924 8632 12268 8672
rect 12308 8632 12317 8672
rect 12942 8632 13036 8672
rect 13076 8632 13085 8672
rect 14766 8632 14860 8672
rect 14900 8632 14909 8672
rect 15726 8632 15820 8672
rect 15860 8632 15869 8672
rect 18019 8632 18028 8672
rect 18068 8632 19412 8672
rect 3715 8631 3773 8632
rect 3235 8548 3244 8588
rect 3284 8548 4972 8588
rect 5012 8548 5021 8588
rect 0 8504 80 8524
rect 5356 8504 5396 8632
rect 7372 8588 7412 8632
rect 8803 8631 8861 8632
rect 9763 8631 9821 8632
rect 13027 8631 13085 8632
rect 14851 8631 14909 8632
rect 15811 8631 15869 8632
rect 7372 8548 10924 8588
rect 10964 8548 10973 8588
rect 11320 8548 19276 8588
rect 19316 8548 19325 8588
rect 5539 8504 5597 8505
rect 11320 8504 11360 8548
rect 13987 8504 14045 8505
rect 18883 8504 18941 8505
rect 0 8464 1900 8504
rect 1940 8464 1949 8504
rect 3811 8464 3820 8504
rect 3860 8464 5260 8504
rect 5300 8464 5309 8504
rect 5356 8464 5548 8504
rect 5588 8464 11360 8504
rect 13795 8464 13804 8504
rect 13844 8464 13996 8504
rect 14036 8464 14045 8504
rect 15235 8464 15244 8504
rect 15284 8464 18892 8504
rect 18932 8464 18941 8504
rect 0 8444 80 8464
rect 5539 8463 5597 8464
rect 13987 8463 14045 8464
rect 18883 8463 18941 8464
rect 19276 8420 19316 8548
rect 19372 8504 19412 8632
rect 19459 8632 19468 8672
rect 19508 8632 20140 8672
rect 20180 8632 21004 8672
rect 21044 8632 21053 8672
rect 21571 8632 21580 8672
rect 21620 8632 22964 8672
rect 23116 8632 26092 8672
rect 26132 8632 26141 8672
rect 26467 8632 26476 8672
rect 26516 8632 29164 8672
rect 29204 8632 29932 8672
rect 29972 8632 29981 8672
rect 30115 8632 30124 8672
rect 30164 8632 34636 8672
rect 34676 8632 34685 8672
rect 19459 8631 19517 8632
rect 19372 8464 21196 8504
rect 21236 8464 22540 8504
rect 22580 8464 22589 8504
rect 2083 8380 2092 8420
rect 2132 8380 16972 8420
rect 17012 8380 17021 8420
rect 19276 8380 23020 8420
rect 23060 8380 23069 8420
rect 4099 8336 4157 8337
rect 19459 8336 19517 8337
rect 20611 8336 20669 8337
rect 23116 8336 23156 8632
rect 30787 8588 30845 8589
rect 30702 8548 30796 8588
rect 30836 8548 30845 8588
rect 32899 8548 32908 8588
rect 32948 8548 37820 8588
rect 30787 8547 30845 8548
rect 27715 8504 27773 8505
rect 25603 8464 25612 8504
rect 25652 8464 26092 8504
rect 26132 8464 26141 8504
rect 27630 8464 27724 8504
rect 27764 8464 27773 8504
rect 27715 8463 27773 8464
rect 27907 8504 27965 8505
rect 30979 8504 31037 8505
rect 31363 8504 31421 8505
rect 31747 8504 31805 8505
rect 37780 8504 37820 8548
rect 39715 8504 39773 8505
rect 42928 8504 43008 8524
rect 27907 8464 27916 8504
rect 27956 8464 28050 8504
rect 29059 8464 29068 8504
rect 29108 8464 29452 8504
rect 29492 8464 29501 8504
rect 29731 8464 29740 8504
rect 29780 8464 30028 8504
rect 30068 8464 30077 8504
rect 30894 8464 30988 8504
rect 31028 8464 31037 8504
rect 31278 8464 31372 8504
rect 31412 8464 31421 8504
rect 31662 8464 31756 8504
rect 31796 8464 31805 8504
rect 27907 8463 27965 8464
rect 30979 8463 31037 8464
rect 31363 8463 31421 8464
rect 31747 8463 31805 8464
rect 32524 8464 36172 8504
rect 36212 8464 36221 8504
rect 37780 8464 38668 8504
rect 38708 8464 38717 8504
rect 39630 8464 39724 8504
rect 39764 8464 39773 8504
rect 41059 8464 41068 8504
rect 41108 8464 43008 8504
rect 32524 8420 32564 8464
rect 39715 8463 39773 8464
rect 42928 8444 43008 8464
rect 32995 8420 33053 8421
rect 26371 8380 26380 8420
rect 26420 8380 32564 8420
rect 32910 8380 33004 8420
rect 33044 8380 33053 8420
rect 32995 8379 33053 8380
rect 33196 8380 38956 8420
rect 38996 8380 41260 8420
rect 41300 8380 41309 8420
rect 3340 8296 4108 8336
rect 4148 8296 4300 8336
rect 4340 8296 4820 8336
rect 4919 8296 4928 8336
rect 4968 8296 5010 8336
rect 5050 8296 5092 8336
rect 5132 8296 5174 8336
rect 5214 8296 5256 8336
rect 5296 8296 5305 8336
rect 5827 8296 5836 8336
rect 5876 8296 6220 8336
rect 6260 8296 11360 8336
rect 13987 8296 13996 8336
rect 14036 8296 14284 8336
rect 14324 8296 15724 8336
rect 15764 8296 16204 8336
rect 16244 8296 18220 8336
rect 18260 8296 19468 8336
rect 19508 8296 19517 8336
rect 20039 8296 20048 8336
rect 20088 8296 20130 8336
rect 20170 8296 20212 8336
rect 20252 8296 20294 8336
rect 20334 8296 20376 8336
rect 20416 8296 20425 8336
rect 20611 8296 20620 8336
rect 20660 8296 23156 8336
rect 25315 8296 25324 8336
rect 25364 8296 27340 8336
rect 27380 8296 27389 8336
rect 28675 8296 28684 8336
rect 28724 8296 33100 8336
rect 33140 8296 33149 8336
rect 0 8168 80 8188
rect 3340 8168 3380 8296
rect 4099 8295 4157 8296
rect 4780 8252 4820 8296
rect 6595 8252 6653 8253
rect 11320 8252 11360 8296
rect 19459 8295 19517 8296
rect 20611 8295 20669 8296
rect 23299 8252 23357 8253
rect 26851 8252 26909 8253
rect 3523 8212 3532 8252
rect 3572 8212 4588 8252
rect 4628 8212 4637 8252
rect 4780 8212 5932 8252
rect 5972 8212 5981 8252
rect 6510 8212 6604 8252
rect 6644 8212 6653 8252
rect 10915 8212 10924 8252
rect 10964 8212 10973 8252
rect 11320 8212 14092 8252
rect 14132 8212 14141 8252
rect 15331 8212 15340 8252
rect 15380 8212 23252 8252
rect 6595 8211 6653 8212
rect 10924 8168 10964 8212
rect 23212 8168 23252 8212
rect 23299 8212 23308 8252
rect 23348 8212 23442 8252
rect 26766 8212 26860 8252
rect 26900 8212 26909 8252
rect 27235 8212 27244 8252
rect 27284 8212 32908 8252
rect 32948 8212 32957 8252
rect 23299 8211 23357 8212
rect 26851 8211 26909 8212
rect 33091 8168 33149 8169
rect 0 8128 1420 8168
rect 1460 8128 1469 8168
rect 1699 8128 1708 8168
rect 1748 8128 3340 8168
rect 3380 8128 3389 8168
rect 3907 8128 3916 8168
rect 3956 8128 6028 8168
rect 6068 8128 6077 8168
rect 10924 8128 15148 8168
rect 15188 8128 18124 8168
rect 18164 8128 20812 8168
rect 20852 8128 20861 8168
rect 20995 8128 21004 8168
rect 21044 8128 21053 8168
rect 23203 8128 23212 8168
rect 23252 8128 26956 8168
rect 26996 8128 27005 8168
rect 27523 8128 27532 8168
rect 27572 8128 28108 8168
rect 28148 8128 28157 8168
rect 28780 8128 29000 8168
rect 29539 8128 29548 8168
rect 29588 8128 30220 8168
rect 30260 8128 30988 8168
rect 31028 8128 31037 8168
rect 31555 8128 31564 8168
rect 31604 8128 31756 8168
rect 31796 8128 31805 8168
rect 32803 8128 32812 8168
rect 32852 8128 33100 8168
rect 33140 8128 33149 8168
rect 0 8108 80 8128
rect 11395 8084 11453 8085
rect 11395 8044 11404 8084
rect 11444 8044 11788 8084
rect 11828 8044 11837 8084
rect 11395 8043 11453 8044
rect 6403 8000 6461 8001
rect 12355 8000 12413 8001
rect 21004 8000 21044 8128
rect 28780 8084 28820 8128
rect 21763 8044 21772 8084
rect 21812 8044 22444 8084
rect 22484 8044 22493 8084
rect 24355 8044 24364 8084
rect 24404 8044 28820 8084
rect 28960 8084 29000 8128
rect 33091 8127 33149 8128
rect 33196 8084 33236 8380
rect 35159 8296 35168 8336
rect 35208 8296 35250 8336
rect 35290 8296 35332 8336
rect 35372 8296 35414 8336
rect 35454 8296 35496 8336
rect 35536 8296 35545 8336
rect 33475 8212 33484 8252
rect 33524 8212 38572 8252
rect 38612 8212 38621 8252
rect 42928 8168 43008 8188
rect 28960 8044 33236 8084
rect 33484 8128 40492 8168
rect 40532 8128 40541 8168
rect 40675 8128 40684 8168
rect 40724 8128 43008 8168
rect 4483 7960 4492 8000
rect 4532 7960 5356 8000
rect 5396 7960 5405 8000
rect 5635 7960 5644 8000
rect 5684 7960 6412 8000
rect 6452 7960 6461 8000
rect 12270 7960 12364 8000
rect 12404 7960 12748 8000
rect 12788 7960 12797 8000
rect 14083 7960 14092 8000
rect 14132 7960 14668 8000
rect 14708 7960 17644 8000
rect 17684 7960 17693 8000
rect 20803 7960 20812 8000
rect 20852 7960 21044 8000
rect 22243 8000 22301 8001
rect 28003 8000 28061 8001
rect 28867 8000 28925 8001
rect 22243 7960 22252 8000
rect 22292 7960 25900 8000
rect 25940 7960 25949 8000
rect 27918 7960 28012 8000
rect 28052 7960 28061 8000
rect 28195 7960 28204 8000
rect 28244 7960 28820 8000
rect 6403 7959 6461 7960
rect 12355 7959 12413 7960
rect 6019 7916 6077 7917
rect 17644 7916 17684 7960
rect 22243 7959 22301 7960
rect 28003 7959 28061 7960
rect 23875 7916 23933 7917
rect 24067 7916 24125 7917
rect 28780 7916 28820 7960
rect 28867 7960 28876 8000
rect 28916 7960 29740 8000
rect 29780 7960 33292 8000
rect 33332 7960 33341 8000
rect 28867 7959 28925 7960
rect 6019 7876 6028 7916
rect 6068 7876 6988 7916
rect 7028 7876 7037 7916
rect 11683 7876 11692 7916
rect 11732 7876 12556 7916
rect 12596 7876 12605 7916
rect 16291 7876 16300 7916
rect 16340 7876 16876 7916
rect 16916 7876 16925 7916
rect 17644 7876 20908 7916
rect 20948 7876 21772 7916
rect 21812 7876 21821 7916
rect 23875 7876 23884 7916
rect 23924 7876 24076 7916
rect 24116 7876 24125 7916
rect 6019 7875 6077 7876
rect 23875 7875 23933 7876
rect 24067 7875 24125 7876
rect 26092 7876 28724 7916
rect 28780 7876 30220 7916
rect 30260 7876 30740 7916
rect 30787 7876 30796 7916
rect 30836 7876 31564 7916
rect 31604 7876 31613 7916
rect 0 7832 80 7852
rect 1891 7832 1949 7833
rect 5443 7832 5501 7833
rect 26092 7832 26132 7876
rect 28579 7832 28637 7833
rect 0 7792 1900 7832
rect 1940 7792 1949 7832
rect 5358 7792 5452 7832
rect 5492 7792 5501 7832
rect 0 7772 80 7792
rect 1891 7791 1949 7792
rect 5443 7791 5501 7792
rect 5548 7792 6316 7832
rect 6356 7792 15340 7832
rect 15380 7792 15389 7832
rect 15619 7792 15628 7832
rect 15668 7792 18604 7832
rect 18644 7792 18653 7832
rect 21571 7792 21580 7832
rect 21620 7792 21868 7832
rect 21908 7792 21917 7832
rect 22051 7792 22060 7832
rect 22100 7792 26132 7832
rect 26275 7792 26284 7832
rect 26324 7792 28588 7832
rect 28628 7792 28637 7832
rect 5548 7748 5588 7792
rect 28579 7791 28637 7792
rect 5347 7708 5356 7748
rect 5396 7708 5588 7748
rect 5731 7748 5789 7749
rect 20707 7748 20765 7749
rect 28684 7748 28724 7876
rect 30700 7832 30740 7876
rect 33484 7832 33524 8128
rect 42928 8108 43008 8128
rect 37315 7960 37324 8000
rect 37364 7960 37373 8000
rect 37603 7960 37612 8000
rect 37652 7960 38284 8000
rect 38324 7960 38333 8000
rect 37324 7832 37364 7960
rect 42928 7832 43008 7852
rect 30700 7792 33524 7832
rect 36547 7792 36556 7832
rect 36596 7792 39340 7832
rect 39380 7792 39389 7832
rect 41059 7792 41068 7832
rect 41108 7792 43008 7832
rect 42928 7772 43008 7792
rect 31363 7748 31421 7749
rect 32611 7748 32669 7749
rect 5731 7708 5740 7748
rect 5780 7708 6028 7748
rect 6068 7708 15052 7748
rect 15092 7708 18028 7748
rect 18068 7708 18077 7748
rect 18787 7708 18796 7748
rect 18836 7708 18876 7748
rect 20622 7708 20716 7748
rect 20756 7708 28204 7748
rect 28244 7708 28253 7748
rect 28684 7708 31220 7748
rect 31278 7708 31372 7748
rect 31412 7708 31421 7748
rect 32526 7708 32620 7748
rect 32660 7708 32669 7748
rect 33283 7708 33292 7748
rect 33332 7708 41356 7748
rect 41396 7708 41405 7748
rect 5731 7707 5789 7708
rect 18796 7664 18836 7708
rect 20707 7707 20765 7708
rect 4675 7624 4684 7664
rect 4724 7624 15244 7664
rect 15284 7624 15293 7664
rect 17731 7624 17740 7664
rect 17780 7624 21676 7664
rect 21716 7624 21725 7664
rect 25699 7624 25708 7664
rect 25748 7624 26380 7664
rect 26420 7624 26429 7664
rect 26851 7624 26860 7664
rect 26900 7624 27052 7664
rect 27092 7624 28300 7664
rect 28340 7624 29740 7664
rect 29780 7624 29789 7664
rect 12067 7580 12125 7581
rect 31180 7580 31220 7708
rect 31363 7707 31421 7708
rect 32611 7707 32669 7708
rect 34627 7664 34685 7665
rect 32419 7624 32428 7664
rect 32468 7624 32908 7664
rect 32948 7624 32957 7664
rect 33772 7624 34636 7664
rect 34676 7624 36556 7664
rect 36596 7624 36605 7664
rect 33772 7580 33812 7624
rect 34627 7623 34685 7624
rect 3679 7540 3688 7580
rect 3728 7540 3770 7580
rect 3810 7540 3852 7580
rect 3892 7540 3934 7580
rect 3974 7540 4016 7580
rect 4056 7540 4065 7580
rect 9283 7540 9292 7580
rect 9332 7540 11020 7580
rect 11060 7540 11069 7580
rect 11982 7540 12076 7580
rect 12116 7540 12125 7580
rect 18799 7540 18808 7580
rect 18848 7540 18890 7580
rect 18930 7540 18972 7580
rect 19012 7540 19054 7580
rect 19094 7540 19136 7580
rect 19176 7540 19185 7580
rect 20803 7540 20812 7580
rect 20852 7540 22060 7580
rect 22100 7540 22109 7580
rect 25507 7540 25516 7580
rect 25556 7540 25804 7580
rect 25844 7540 25853 7580
rect 26179 7540 26188 7580
rect 26228 7540 29356 7580
rect 29396 7540 29405 7580
rect 29539 7540 29548 7580
rect 29588 7540 29932 7580
rect 29972 7540 29981 7580
rect 31180 7540 33812 7580
rect 33919 7540 33928 7580
rect 33968 7540 34010 7580
rect 34050 7540 34092 7580
rect 34132 7540 34174 7580
rect 34214 7540 34256 7580
rect 34296 7540 34305 7580
rect 39811 7540 39820 7580
rect 39860 7540 40396 7580
rect 40436 7540 40445 7580
rect 12067 7539 12125 7540
rect 0 7496 80 7516
rect 2467 7496 2525 7497
rect 42928 7496 43008 7516
rect 0 7456 2476 7496
rect 2516 7456 2525 7496
rect 7459 7456 7468 7496
rect 7508 7456 18316 7496
rect 18356 7456 18365 7496
rect 23491 7456 23500 7496
rect 23540 7456 24556 7496
rect 24596 7456 28876 7496
rect 28916 7456 28925 7496
rect 30883 7456 30892 7496
rect 30932 7456 31948 7496
rect 31988 7456 31997 7496
rect 41443 7456 41452 7496
rect 41492 7456 43008 7496
rect 0 7436 80 7456
rect 2467 7455 2525 7456
rect 42928 7436 43008 7456
rect 11491 7412 11549 7413
rect 35011 7412 35069 7413
rect 10435 7372 10444 7412
rect 10484 7372 10924 7412
rect 10964 7372 10973 7412
rect 11491 7372 11500 7412
rect 11540 7372 11634 7412
rect 11875 7372 11884 7412
rect 11924 7372 12076 7412
rect 12116 7372 12125 7412
rect 12268 7372 13132 7412
rect 13172 7372 13181 7412
rect 14371 7372 14380 7412
rect 14420 7372 24364 7412
rect 24404 7372 24413 7412
rect 25123 7372 25132 7412
rect 25172 7372 29260 7412
rect 29300 7372 29309 7412
rect 32515 7372 32524 7412
rect 32564 7372 35020 7412
rect 35060 7372 35069 7412
rect 11491 7371 11549 7372
rect 12268 7328 12308 7372
rect 35011 7371 35069 7372
rect 26275 7328 26333 7329
rect 26851 7328 26909 7329
rect 31939 7328 31997 7329
rect 8044 7288 10732 7328
rect 10772 7288 12308 7328
rect 12940 7288 26284 7328
rect 26324 7288 26333 7328
rect 26766 7288 26860 7328
rect 26900 7288 26909 7328
rect 4579 7244 4637 7245
rect 4494 7204 4588 7244
rect 4628 7204 4637 7244
rect 4579 7203 4637 7204
rect 0 7160 80 7180
rect 8044 7161 8084 7288
rect 12940 7244 12980 7288
rect 26275 7287 26333 7288
rect 26851 7287 26909 7288
rect 28960 7288 28972 7328
rect 29012 7288 29021 7328
rect 31854 7288 31948 7328
rect 31988 7288 39148 7328
rect 39188 7288 39197 7328
rect 28960 7244 29000 7288
rect 31939 7287 31997 7288
rect 40291 7244 40349 7245
rect 9475 7204 9484 7244
rect 9524 7204 9868 7244
rect 9908 7204 9917 7244
rect 11491 7204 11500 7244
rect 11540 7204 12748 7244
rect 12788 7204 12797 7244
rect 12931 7204 12940 7244
rect 12980 7204 12989 7244
rect 15907 7204 15916 7244
rect 15956 7204 29000 7244
rect 31651 7204 31660 7244
rect 31700 7204 32812 7244
rect 32852 7204 32861 7244
rect 40291 7204 40300 7244
rect 40340 7204 40876 7244
rect 40916 7204 40925 7244
rect 40291 7203 40349 7204
rect 4099 7160 4157 7161
rect 5347 7160 5405 7161
rect 8035 7160 8093 7161
rect 17635 7160 17693 7161
rect 0 7120 2476 7160
rect 2516 7120 2525 7160
rect 3811 7120 3820 7160
rect 3860 7120 4108 7160
rect 4148 7120 4157 7160
rect 4387 7120 4396 7160
rect 4436 7120 4780 7160
rect 4820 7120 5356 7160
rect 5396 7120 5405 7160
rect 6499 7120 6508 7160
rect 6548 7120 7276 7160
rect 7316 7120 7325 7160
rect 7950 7120 8044 7160
rect 8084 7120 8093 7160
rect 10819 7120 10828 7160
rect 10868 7120 13516 7160
rect 13556 7120 13565 7160
rect 17550 7120 17644 7160
rect 17684 7120 17693 7160
rect 0 7100 80 7120
rect 4099 7119 4157 7120
rect 5347 7119 5405 7120
rect 8035 7119 8093 7120
rect 17635 7119 17693 7120
rect 19363 7160 19421 7161
rect 27811 7160 27869 7161
rect 42928 7160 43008 7180
rect 19363 7120 19372 7160
rect 19412 7120 19660 7160
rect 19700 7120 19709 7160
rect 20899 7120 20908 7160
rect 20948 7120 22636 7160
rect 22676 7120 24172 7160
rect 24212 7120 25132 7160
rect 25172 7120 25612 7160
rect 25652 7120 25661 7160
rect 27715 7120 27724 7160
rect 27764 7120 27820 7160
rect 27860 7120 27869 7160
rect 30979 7120 30988 7160
rect 31028 7120 31564 7160
rect 31604 7120 33004 7160
rect 33044 7120 33196 7160
rect 33236 7120 33245 7160
rect 36067 7120 36076 7160
rect 36116 7120 37516 7160
rect 37556 7120 37565 7160
rect 41059 7120 41068 7160
rect 41108 7120 43008 7160
rect 19363 7119 19421 7120
rect 27811 7119 27869 7120
rect 42928 7100 43008 7120
rect 28963 7076 29021 7077
rect 4003 7036 4012 7076
rect 4052 7036 5836 7076
rect 5876 7036 5885 7076
rect 5932 7036 14380 7076
rect 14420 7036 14429 7076
rect 20140 7036 28972 7076
rect 29012 7036 29021 7076
rect 5932 6992 5972 7036
rect 13795 6992 13853 6993
rect 2755 6952 2764 6992
rect 2804 6952 5972 6992
rect 6211 6952 6220 6992
rect 6260 6952 6700 6992
rect 6740 6952 6749 6992
rect 10339 6952 10348 6992
rect 10388 6952 10540 6992
rect 10580 6952 10589 6992
rect 11320 6952 13132 6992
rect 13172 6952 13804 6992
rect 13844 6952 13853 6992
rect 17251 6952 17260 6992
rect 17300 6952 18892 6992
rect 18932 6952 19276 6992
rect 19316 6952 19325 6992
rect 11320 6908 11360 6952
rect 13795 6951 13853 6952
rect 11491 6908 11549 6909
rect 20140 6908 20180 7036
rect 28963 7035 29021 7036
rect 29539 6992 29597 6993
rect 25507 6952 25516 6992
rect 25556 6952 25804 6992
rect 25844 6952 25853 6992
rect 28675 6952 28684 6992
rect 28724 6952 29164 6992
rect 29204 6952 29213 6992
rect 29539 6952 29548 6992
rect 29588 6952 33676 6992
rect 33716 6952 33725 6992
rect 37780 6952 40876 6992
rect 40916 6952 40925 6992
rect 29539 6951 29597 6952
rect 37780 6908 37820 6952
rect 1891 6868 1900 6908
rect 1940 6868 11360 6908
rect 11406 6868 11500 6908
rect 11540 6868 11549 6908
rect 18979 6868 18988 6908
rect 19028 6868 19852 6908
rect 19892 6868 20180 6908
rect 21475 6868 21484 6908
rect 21524 6868 34540 6908
rect 34580 6868 36268 6908
rect 36308 6868 37820 6908
rect 11491 6867 11549 6868
rect 0 6824 80 6844
rect 42928 6824 43008 6844
rect 0 6784 1516 6824
rect 1556 6784 1565 6824
rect 4919 6784 4928 6824
rect 4968 6784 5010 6824
rect 5050 6784 5092 6824
rect 5132 6784 5174 6824
rect 5214 6784 5256 6824
rect 5296 6784 5305 6824
rect 5635 6784 5644 6824
rect 5684 6784 17740 6824
rect 17780 6784 17789 6824
rect 20039 6784 20048 6824
rect 20088 6784 20130 6824
rect 20170 6784 20212 6824
rect 20252 6784 20294 6824
rect 20334 6784 20376 6824
rect 20416 6784 20425 6824
rect 24835 6784 24844 6824
rect 24884 6784 31564 6824
rect 31604 6784 31613 6824
rect 35159 6784 35168 6824
rect 35208 6784 35250 6824
rect 35290 6784 35332 6824
rect 35372 6784 35414 6824
rect 35454 6784 35496 6824
rect 35536 6784 35545 6824
rect 41443 6784 41452 6824
rect 41492 6784 43008 6824
rect 0 6764 80 6784
rect 42928 6764 43008 6784
rect 7171 6740 7229 6741
rect 30211 6740 30269 6741
rect 3907 6700 3916 6740
rect 3956 6700 4588 6740
rect 4628 6700 4637 6740
rect 7171 6700 7180 6740
rect 7220 6700 7314 6740
rect 9859 6700 9868 6740
rect 9908 6700 12556 6740
rect 12596 6700 20620 6740
rect 20660 6700 20669 6740
rect 27139 6700 27148 6740
rect 27188 6700 27532 6740
rect 27572 6700 27581 6740
rect 30211 6700 30220 6740
rect 30260 6700 37652 6740
rect 7171 6699 7229 6700
rect 30211 6699 30269 6700
rect 21667 6656 21725 6657
rect 37612 6656 37652 6700
rect 2500 6616 7468 6656
rect 7508 6616 7517 6656
rect 9475 6616 9484 6656
rect 9524 6616 18988 6656
rect 19028 6616 19037 6656
rect 19747 6616 19756 6656
rect 19796 6616 20332 6656
rect 20372 6616 20381 6656
rect 21283 6616 21292 6656
rect 21332 6616 21484 6656
rect 21524 6616 21533 6656
rect 21667 6616 21676 6656
rect 21716 6616 21964 6656
rect 22004 6616 22013 6656
rect 25219 6616 25228 6656
rect 25268 6616 25708 6656
rect 25748 6616 25757 6656
rect 26179 6616 26188 6656
rect 26228 6616 32084 6656
rect 32995 6616 33004 6656
rect 33044 6616 33676 6656
rect 33716 6616 33725 6656
rect 37603 6616 37612 6656
rect 37652 6616 37661 6656
rect 1132 6532 1708 6572
rect 1748 6532 1757 6572
rect 0 6488 80 6508
rect 1132 6488 1172 6532
rect 2500 6488 2540 6616
rect 21667 6615 21725 6616
rect 32044 6572 32084 6616
rect 4483 6532 4492 6572
rect 4532 6532 6604 6572
rect 6644 6532 6653 6572
rect 12163 6532 12172 6572
rect 12212 6532 12460 6572
rect 12500 6532 12509 6572
rect 13507 6532 13516 6572
rect 13556 6532 15340 6572
rect 15380 6532 16492 6572
rect 16532 6532 16541 6572
rect 18307 6532 18316 6572
rect 18356 6532 19852 6572
rect 19892 6532 19901 6572
rect 21187 6532 21196 6572
rect 21236 6532 22060 6572
rect 22100 6532 23596 6572
rect 23636 6532 24076 6572
rect 24116 6532 24125 6572
rect 28195 6532 28204 6572
rect 28244 6532 29452 6572
rect 29492 6532 29644 6572
rect 29684 6532 29693 6572
rect 32044 6532 38420 6572
rect 5539 6488 5597 6489
rect 14188 6488 14228 6532
rect 21667 6488 21725 6489
rect 0 6448 1172 6488
rect 1219 6448 1228 6488
rect 1268 6448 2540 6488
rect 2851 6448 2860 6488
rect 2900 6448 4012 6488
rect 4052 6448 4061 6488
rect 5155 6448 5164 6488
rect 5204 6448 5548 6488
rect 5588 6448 5597 6488
rect 6019 6448 6028 6488
rect 6068 6448 6508 6488
rect 6548 6448 7180 6488
rect 7220 6448 7229 6488
rect 8803 6448 8812 6488
rect 8852 6448 9580 6488
rect 9620 6448 10828 6488
rect 10868 6448 10877 6488
rect 10924 6448 11020 6488
rect 11060 6448 11980 6488
rect 12020 6448 13708 6488
rect 13748 6448 13757 6488
rect 14179 6448 14188 6488
rect 14228 6448 14268 6488
rect 14467 6448 14476 6488
rect 14516 6448 16396 6488
rect 16436 6448 16445 6488
rect 18883 6448 18892 6488
rect 18932 6448 21676 6488
rect 21716 6448 21725 6488
rect 21955 6448 21964 6488
rect 22004 6448 22156 6488
rect 22196 6448 24460 6488
rect 24500 6448 26668 6488
rect 26708 6448 26717 6488
rect 29251 6448 29260 6488
rect 29300 6448 31948 6488
rect 31988 6448 31997 6488
rect 0 6428 80 6448
rect 5539 6447 5597 6448
rect 6019 6404 6077 6405
rect 10723 6404 10781 6405
rect 5731 6364 5740 6404
rect 5780 6364 6028 6404
rect 6068 6364 6077 6404
rect 6211 6364 6220 6404
rect 6260 6364 6988 6404
rect 7028 6364 7037 6404
rect 10638 6364 10732 6404
rect 10772 6364 10781 6404
rect 6019 6363 6077 6364
rect 10723 6363 10781 6364
rect 1603 6320 1661 6321
rect 1891 6320 1949 6321
rect 10924 6320 10964 6448
rect 21667 6447 21725 6448
rect 28963 6404 29021 6405
rect 32044 6404 32084 6532
rect 33379 6488 33437 6489
rect 38380 6488 38420 6532
rect 42928 6488 43008 6508
rect 33294 6448 33388 6488
rect 33428 6448 34444 6488
rect 34484 6448 34493 6488
rect 34627 6448 34636 6488
rect 34676 6448 35596 6488
rect 35636 6448 35645 6488
rect 38371 6448 38380 6488
rect 38420 6448 38429 6488
rect 38563 6448 38572 6488
rect 38612 6448 38860 6488
rect 38900 6448 38909 6488
rect 41059 6448 41068 6488
rect 41108 6448 43008 6488
rect 33379 6447 33437 6448
rect 34444 6404 34484 6448
rect 42928 6428 43008 6448
rect 41251 6404 41309 6405
rect 13027 6364 13036 6404
rect 13076 6364 13804 6404
rect 13844 6364 15916 6404
rect 15956 6364 15965 6404
rect 16012 6364 28492 6404
rect 28532 6364 28541 6404
rect 28963 6364 28972 6404
rect 29012 6364 29106 6404
rect 32035 6364 32044 6404
rect 32084 6364 32093 6404
rect 34444 6364 36556 6404
rect 36596 6364 36605 6404
rect 40003 6364 40012 6404
rect 40052 6364 40396 6404
rect 40436 6364 40445 6404
rect 41166 6364 41260 6404
rect 41300 6364 41309 6404
rect 16012 6320 16052 6364
rect 28963 6363 29021 6364
rect 41251 6363 41309 6364
rect 35683 6320 35741 6321
rect 40195 6320 40253 6321
rect 1518 6280 1612 6320
rect 1652 6280 1661 6320
rect 1806 6280 1900 6320
rect 1940 6280 1949 6320
rect 4195 6280 4204 6320
rect 4244 6280 4684 6320
rect 4724 6280 5164 6320
rect 5204 6280 5213 6320
rect 6115 6280 6124 6320
rect 6164 6280 6316 6320
rect 6356 6280 6365 6320
rect 6787 6280 6796 6320
rect 6836 6280 7564 6320
rect 7604 6280 7613 6320
rect 8707 6280 8716 6320
rect 8756 6280 8908 6320
rect 8948 6280 9964 6320
rect 10004 6280 10636 6320
rect 10676 6280 10685 6320
rect 10819 6280 10828 6320
rect 10868 6280 10964 6320
rect 11980 6280 12268 6320
rect 12308 6280 15820 6320
rect 15860 6280 16052 6320
rect 19075 6280 19084 6320
rect 19124 6280 20620 6320
rect 20660 6280 20669 6320
rect 24547 6280 24556 6320
rect 24596 6280 25996 6320
rect 26036 6280 26045 6320
rect 30787 6280 30796 6320
rect 30836 6280 31468 6320
rect 31508 6280 31517 6320
rect 35598 6280 35692 6320
rect 35732 6280 35741 6320
rect 39780 6280 39820 6320
rect 39860 6280 39869 6320
rect 40110 6280 40204 6320
rect 40244 6280 40253 6320
rect 1603 6279 1661 6280
rect 1891 6279 1949 6280
rect 4675 6236 4733 6237
rect 11980 6236 12020 6280
rect 35683 6279 35741 6280
rect 39820 6236 39860 6280
rect 40195 6279 40253 6280
rect 4675 6196 4684 6236
rect 4724 6196 4780 6236
rect 4820 6196 4829 6236
rect 5164 6196 5644 6236
rect 5684 6196 5693 6236
rect 6595 6196 6604 6236
rect 6644 6196 7372 6236
rect 7412 6196 7421 6236
rect 11971 6196 11980 6236
rect 12020 6196 12029 6236
rect 16003 6196 16012 6236
rect 16052 6196 19372 6236
rect 19412 6196 19421 6236
rect 34339 6196 34348 6236
rect 34388 6196 34828 6236
rect 34868 6196 34877 6236
rect 39820 6196 40300 6236
rect 40340 6196 40349 6236
rect 4675 6195 4733 6196
rect 0 6152 80 6172
rect 1699 6152 1757 6153
rect 4291 6152 4349 6153
rect 5164 6152 5204 6196
rect 6595 6152 6653 6153
rect 42928 6152 43008 6172
rect 0 6112 1708 6152
rect 1748 6112 1757 6152
rect 0 6092 80 6112
rect 1699 6111 1757 6112
rect 4204 6112 4300 6152
rect 4340 6112 5204 6152
rect 6499 6112 6508 6152
rect 6548 6112 6604 6152
rect 6644 6112 18124 6152
rect 18164 6112 18173 6152
rect 20899 6112 20908 6152
rect 20948 6112 21388 6152
rect 21428 6112 27244 6152
rect 27284 6112 27293 6152
rect 28003 6112 28012 6152
rect 28052 6112 29108 6152
rect 41059 6112 41068 6152
rect 41108 6112 43008 6152
rect 3679 6028 3688 6068
rect 3728 6028 3770 6068
rect 3810 6028 3852 6068
rect 3892 6028 3934 6068
rect 3974 6028 4016 6068
rect 4056 6028 4065 6068
rect 4204 5984 4244 6112
rect 4291 6111 4349 6112
rect 6595 6111 6653 6112
rect 14851 6068 14909 6069
rect 4771 6028 4780 6068
rect 4820 6028 14860 6068
rect 14900 6028 14909 6068
rect 18799 6028 18808 6068
rect 18848 6028 18890 6068
rect 18930 6028 18972 6068
rect 19012 6028 19054 6068
rect 19094 6028 19136 6068
rect 19176 6028 19185 6068
rect 19276 6028 21100 6068
rect 21140 6028 22540 6068
rect 22580 6028 22589 6068
rect 22723 6028 22732 6068
rect 22772 6028 23116 6068
rect 23156 6028 23165 6068
rect 14851 6027 14909 6028
rect 4387 5984 4445 5985
rect 7171 5984 7229 5985
rect 19276 5984 19316 6028
rect 27811 5984 27869 5985
rect 28963 5984 29021 5985
rect 1699 5944 1708 5984
rect 1748 5944 4204 5984
rect 4244 5944 4253 5984
rect 4302 5944 4396 5984
rect 4436 5944 4445 5984
rect 5827 5944 5836 5984
rect 5876 5944 6124 5984
rect 6164 5944 6173 5984
rect 6979 5944 6988 5984
rect 7028 5944 7180 5984
rect 7220 5944 7229 5984
rect 9283 5944 9292 5984
rect 9332 5944 12460 5984
rect 12500 5944 12509 5984
rect 14851 5944 14860 5984
rect 14900 5944 19316 5984
rect 19363 5944 19372 5984
rect 19412 5944 26092 5984
rect 26132 5944 26141 5984
rect 27811 5944 27820 5984
rect 27860 5944 28012 5984
rect 28052 5944 28061 5984
rect 28960 5944 28972 5984
rect 29012 5944 29021 5984
rect 4387 5943 4445 5944
rect 7171 5943 7229 5944
rect 27811 5943 27869 5944
rect 28960 5943 29021 5944
rect 21667 5900 21725 5901
rect 28960 5900 29000 5943
rect 1507 5860 1516 5900
rect 1556 5860 7660 5900
rect 7700 5860 10732 5900
rect 10772 5860 10781 5900
rect 11011 5860 11020 5900
rect 11060 5860 15532 5900
rect 15572 5860 15581 5900
rect 17635 5860 17644 5900
rect 17684 5860 21292 5900
rect 21332 5860 21341 5900
rect 21582 5860 21676 5900
rect 21716 5860 21725 5900
rect 22435 5860 22444 5900
rect 22484 5860 29000 5900
rect 29068 5900 29108 6112
rect 42928 6092 43008 6112
rect 30403 6028 30412 6068
rect 30452 6028 30988 6068
rect 31028 6028 31037 6068
rect 33919 6028 33928 6068
rect 33968 6028 34010 6068
rect 34050 6028 34092 6068
rect 34132 6028 34174 6068
rect 34214 6028 34256 6068
rect 34296 6028 34305 6068
rect 37411 6028 37420 6068
rect 37460 6028 38764 6068
rect 38804 6028 38813 6068
rect 31651 5944 31660 5984
rect 31700 5944 34828 5984
rect 34868 5944 36268 5984
rect 36308 5944 36844 5984
rect 36884 5944 36893 5984
rect 29068 5860 40780 5900
rect 40820 5860 40829 5900
rect 21667 5859 21725 5860
rect 0 5816 80 5836
rect 4195 5816 4253 5817
rect 21091 5816 21149 5817
rect 29059 5816 29117 5817
rect 42928 5816 43008 5836
rect 0 5776 2420 5816
rect 0 5756 80 5776
rect 2380 5648 2420 5776
rect 4195 5776 4204 5816
rect 4244 5776 4300 5816
rect 4340 5776 5740 5816
rect 5780 5776 5789 5816
rect 6979 5776 6988 5816
rect 7028 5776 9772 5816
rect 9812 5776 9821 5816
rect 10531 5776 10540 5816
rect 10580 5776 19948 5816
rect 19988 5776 19997 5816
rect 20140 5776 21100 5816
rect 21140 5776 21149 5816
rect 24067 5776 24076 5816
rect 24116 5776 24364 5816
rect 24404 5776 24413 5816
rect 29059 5776 29068 5816
rect 29108 5776 34444 5816
rect 34484 5776 34493 5816
rect 35395 5776 35404 5816
rect 35444 5776 37420 5816
rect 37460 5776 37469 5816
rect 41443 5776 41452 5816
rect 41492 5776 43008 5816
rect 4195 5775 4253 5776
rect 20140 5732 20180 5776
rect 21091 5775 21149 5776
rect 29059 5775 29117 5776
rect 42928 5756 43008 5776
rect 20611 5732 20669 5733
rect 2500 5692 16300 5732
rect 16340 5692 17644 5732
rect 17684 5692 17693 5732
rect 18595 5692 18604 5732
rect 18644 5692 20180 5732
rect 20236 5692 20620 5732
rect 20660 5692 20669 5732
rect 2500 5648 2540 5692
rect 2380 5608 2540 5648
rect 4099 5648 4157 5649
rect 5731 5648 5789 5649
rect 6019 5648 6077 5649
rect 16099 5648 16157 5649
rect 20236 5648 20276 5692
rect 20611 5691 20669 5692
rect 23299 5732 23357 5733
rect 23299 5692 23308 5732
rect 23348 5692 36500 5732
rect 36547 5692 36556 5732
rect 36596 5692 40876 5732
rect 40916 5692 40925 5732
rect 23299 5691 23357 5692
rect 25795 5648 25853 5649
rect 36460 5648 36500 5692
rect 4099 5608 4108 5648
rect 4148 5608 4780 5648
rect 4820 5608 4829 5648
rect 5155 5608 5164 5648
rect 5204 5608 5548 5648
rect 5588 5608 5597 5648
rect 5731 5608 5740 5648
rect 5780 5608 5836 5648
rect 5876 5608 5885 5648
rect 6019 5608 6028 5648
rect 6068 5608 6796 5648
rect 6836 5608 7948 5648
rect 7988 5608 7997 5648
rect 9283 5608 9292 5648
rect 9332 5608 9341 5648
rect 9571 5608 9580 5648
rect 9620 5608 11020 5648
rect 11060 5608 11069 5648
rect 13699 5608 13708 5648
rect 13748 5608 14284 5648
rect 14324 5608 14860 5648
rect 14900 5608 14909 5648
rect 16014 5608 16108 5648
rect 16148 5608 16157 5648
rect 17251 5608 17260 5648
rect 17300 5608 17548 5648
rect 17588 5608 17597 5648
rect 18115 5608 18124 5648
rect 18164 5608 20276 5648
rect 20323 5608 20332 5648
rect 20372 5608 23500 5648
rect 23540 5608 23549 5648
rect 25710 5608 25804 5648
rect 25844 5608 25853 5648
rect 27811 5608 27820 5648
rect 27860 5608 34924 5648
rect 34964 5608 34973 5648
rect 36451 5608 36460 5648
rect 36500 5608 36509 5648
rect 38947 5608 38956 5648
rect 38996 5608 41164 5648
rect 41204 5608 41213 5648
rect 4099 5607 4157 5608
rect 5731 5607 5789 5608
rect 6019 5607 6077 5608
rect 9292 5564 9332 5608
rect 16099 5607 16157 5608
rect 25795 5607 25853 5608
rect 25804 5564 25844 5607
rect 34924 5564 34964 5608
rect 2500 5524 9332 5564
rect 17731 5524 17740 5564
rect 17780 5524 18028 5564
rect 18068 5524 18077 5564
rect 19843 5524 19852 5564
rect 19892 5524 22924 5564
rect 22964 5524 22973 5564
rect 25804 5524 29000 5564
rect 29923 5524 29932 5564
rect 29972 5524 30220 5564
rect 30260 5524 30269 5564
rect 30595 5524 30604 5564
rect 30644 5524 31756 5564
rect 31796 5524 31805 5564
rect 32131 5524 32140 5564
rect 32180 5524 32716 5564
rect 32756 5524 32765 5564
rect 34924 5524 36748 5564
rect 36788 5524 36940 5564
rect 36980 5524 36989 5564
rect 0 5480 80 5500
rect 2500 5480 2540 5524
rect 5251 5480 5309 5481
rect 28291 5480 28349 5481
rect 0 5440 1228 5480
rect 1268 5440 1277 5480
rect 2467 5440 2476 5480
rect 2516 5440 2540 5480
rect 5166 5440 5260 5480
rect 5300 5440 5309 5480
rect 5443 5440 5452 5480
rect 5492 5440 7084 5480
rect 7124 5440 7133 5480
rect 7267 5440 7276 5480
rect 7316 5440 7468 5480
rect 7508 5440 7517 5480
rect 7651 5440 7660 5480
rect 7700 5440 18508 5480
rect 18548 5440 20908 5480
rect 20948 5440 20957 5480
rect 26371 5440 26380 5480
rect 26420 5440 27052 5480
rect 27092 5440 27101 5480
rect 28206 5440 28300 5480
rect 28340 5440 28349 5480
rect 28960 5480 29000 5524
rect 42928 5480 43008 5500
rect 28960 5440 31660 5480
rect 31700 5440 38956 5480
rect 38996 5440 39005 5480
rect 41059 5440 41068 5480
rect 41108 5440 43008 5480
rect 0 5420 80 5440
rect 5251 5439 5309 5440
rect 28291 5439 28349 5440
rect 42928 5420 43008 5440
rect 1411 5356 1420 5396
rect 1460 5356 16108 5396
rect 16148 5356 16157 5396
rect 19459 5356 19468 5396
rect 19508 5356 19948 5396
rect 19988 5356 22868 5396
rect 22915 5356 22924 5396
rect 22964 5356 40876 5396
rect 40916 5356 40925 5396
rect 22828 5312 22868 5356
rect 33091 5312 33149 5313
rect 4919 5272 4928 5312
rect 4968 5272 5010 5312
rect 5050 5272 5092 5312
rect 5132 5272 5174 5312
rect 5214 5272 5256 5312
rect 5296 5272 5305 5312
rect 6307 5272 6316 5312
rect 6356 5272 9580 5312
rect 9620 5272 9629 5312
rect 9763 5272 9772 5312
rect 9812 5272 18604 5312
rect 18644 5272 18653 5312
rect 20039 5272 20048 5312
rect 20088 5272 20130 5312
rect 20170 5272 20212 5312
rect 20252 5272 20294 5312
rect 20334 5272 20376 5312
rect 20416 5272 20425 5312
rect 21196 5272 22444 5312
rect 22484 5272 22493 5312
rect 22828 5272 24364 5312
rect 24404 5272 25036 5312
rect 25076 5272 25085 5312
rect 33006 5272 33100 5312
rect 33140 5272 33149 5312
rect 35159 5272 35168 5312
rect 35208 5272 35250 5312
rect 35290 5272 35332 5312
rect 35372 5272 35414 5312
rect 35454 5272 35496 5312
rect 35536 5272 35545 5312
rect 21196 5228 21236 5272
rect 33091 5271 33149 5272
rect 1795 5188 1804 5228
rect 1844 5188 2476 5228
rect 2516 5188 2525 5228
rect 3043 5188 3052 5228
rect 3092 5188 5644 5228
rect 5684 5188 5932 5228
rect 5972 5188 5981 5228
rect 6211 5188 6220 5228
rect 6260 5188 6892 5228
rect 6932 5188 7276 5228
rect 7316 5188 7660 5228
rect 7700 5188 7709 5228
rect 16867 5188 16876 5228
rect 16916 5188 19084 5228
rect 19124 5188 21236 5228
rect 21283 5188 21292 5228
rect 21332 5188 24460 5228
rect 24500 5188 41260 5228
rect 41300 5188 41309 5228
rect 0 5144 80 5164
rect 42928 5144 43008 5164
rect 0 5104 16012 5144
rect 16052 5104 16061 5144
rect 33763 5104 33772 5144
rect 33812 5104 39244 5144
rect 39284 5104 39293 5144
rect 41443 5104 41452 5144
rect 41492 5104 43008 5144
rect 0 5084 80 5104
rect 42928 5084 43008 5104
rect 3523 5020 3532 5060
rect 3572 5020 5164 5060
rect 5204 5020 5213 5060
rect 5731 5020 5740 5060
rect 5780 5020 6412 5060
rect 6452 5020 6461 5060
rect 12259 5020 12268 5060
rect 12308 5020 23116 5060
rect 23156 5020 23165 5060
rect 23491 5020 23500 5060
rect 23540 5020 25516 5060
rect 25556 5020 25565 5060
rect 25612 5020 26092 5060
rect 26132 5020 27916 5060
rect 27956 5020 27965 5060
rect 28291 5020 28300 5060
rect 28340 5020 32620 5060
rect 32660 5020 32669 5060
rect 38275 5020 38284 5060
rect 38324 5020 38668 5060
rect 38708 5020 38717 5060
rect 1699 4976 1757 4977
rect 5347 4976 5405 4977
rect 15523 4976 15581 4977
rect 25612 4976 25652 5020
rect 1614 4936 1708 4976
rect 1748 4936 1757 4976
rect 3139 4936 3148 4976
rect 3188 4936 3197 4976
rect 3628 4936 4108 4976
rect 4148 4936 4157 4976
rect 5251 4936 5260 4976
rect 5300 4936 5356 4976
rect 5396 4936 5405 4976
rect 9091 4936 9100 4976
rect 9140 4936 9484 4976
rect 9524 4936 9533 4976
rect 9955 4936 9964 4976
rect 10004 4936 10252 4976
rect 10292 4936 10444 4976
rect 10484 4936 10493 4976
rect 12451 4936 12460 4976
rect 12500 4936 15532 4976
rect 15572 4936 15581 4976
rect 19267 4936 19276 4976
rect 19316 4936 19564 4976
rect 19604 4936 19613 4976
rect 22435 4936 22444 4976
rect 22484 4936 22636 4976
rect 22676 4936 25652 4976
rect 27715 4936 27724 4976
rect 27764 4936 29644 4976
rect 29684 4936 29693 4976
rect 32035 4936 32044 4976
rect 32084 4936 32236 4976
rect 32276 4936 32285 4976
rect 37219 4936 37228 4976
rect 37268 4936 40972 4976
rect 41012 4936 41021 4976
rect 1699 4935 1757 4936
rect 3148 4892 3188 4936
rect 3628 4892 3668 4936
rect 5347 4935 5405 4936
rect 15523 4935 15581 4936
rect 3148 4852 3340 4892
rect 3380 4852 3668 4892
rect 3715 4852 3724 4892
rect 3764 4852 6700 4892
rect 6740 4852 6749 4892
rect 10531 4852 10540 4892
rect 10580 4852 10828 4892
rect 10868 4852 13804 4892
rect 13844 4852 13853 4892
rect 21091 4852 21100 4892
rect 21140 4852 21580 4892
rect 21620 4852 21629 4892
rect 21859 4852 21868 4892
rect 21908 4852 22060 4892
rect 22100 4852 22109 4892
rect 23875 4852 23884 4892
rect 23924 4852 30892 4892
rect 30932 4852 30941 4892
rect 39619 4852 39628 4892
rect 39668 4852 40684 4892
rect 40724 4852 40733 4892
rect 0 4808 80 4828
rect 1219 4808 1277 4809
rect 4195 4808 4253 4809
rect 36643 4808 36701 4809
rect 42928 4808 43008 4828
rect 0 4768 1228 4808
rect 1268 4768 1277 4808
rect 3139 4768 3148 4808
rect 3188 4768 4204 4808
rect 4244 4768 4396 4808
rect 4436 4768 4588 4808
rect 4628 4768 5068 4808
rect 5108 4768 6028 4808
rect 6068 4768 6077 4808
rect 18403 4768 18412 4808
rect 18452 4768 20908 4808
rect 20948 4768 20957 4808
rect 27619 4768 27628 4808
rect 27668 4768 29740 4808
rect 29780 4768 33196 4808
rect 33236 4768 33245 4808
rect 36558 4768 36652 4808
rect 36692 4768 36701 4808
rect 38467 4768 38476 4808
rect 38516 4768 38668 4808
rect 38708 4768 39052 4808
rect 39092 4768 40108 4808
rect 40148 4768 40157 4808
rect 41155 4768 41164 4808
rect 41204 4768 43008 4808
rect 0 4748 80 4768
rect 1219 4767 1277 4768
rect 4195 4767 4253 4768
rect 36643 4767 36701 4768
rect 42928 4748 43008 4768
rect 40483 4724 40541 4725
rect 3427 4684 3436 4724
rect 3476 4684 3628 4724
rect 3668 4684 3677 4724
rect 3907 4684 3916 4724
rect 3956 4684 6124 4724
rect 6164 4684 6173 4724
rect 11779 4684 11788 4724
rect 11828 4684 12076 4724
rect 12116 4684 12125 4724
rect 22051 4684 22060 4724
rect 22100 4684 32236 4724
rect 32276 4684 32285 4724
rect 38851 4684 38860 4724
rect 38900 4684 39436 4724
rect 39476 4684 39485 4724
rect 40398 4684 40492 4724
rect 40532 4684 40541 4724
rect 40483 4683 40541 4684
rect 4387 4640 4445 4641
rect 4302 4600 4396 4640
rect 4436 4600 11020 4640
rect 11060 4600 11069 4640
rect 11320 4600 12556 4640
rect 12596 4600 12605 4640
rect 20140 4600 30028 4640
rect 30068 4600 30077 4640
rect 30883 4600 30892 4640
rect 30932 4600 41260 4640
rect 41300 4600 41309 4640
rect 4387 4599 4445 4600
rect 3679 4516 3688 4556
rect 3728 4516 3770 4556
rect 3810 4516 3852 4556
rect 3892 4516 3934 4556
rect 3974 4516 4016 4556
rect 4056 4516 4065 4556
rect 4291 4516 4300 4556
rect 4340 4516 4492 4556
rect 4532 4516 4541 4556
rect 0 4472 80 4492
rect 4771 4472 4829 4473
rect 0 4432 4780 4472
rect 4820 4432 4829 4472
rect 5347 4432 5356 4472
rect 5396 4432 9868 4472
rect 9908 4432 9917 4472
rect 0 4412 80 4432
rect 4771 4431 4829 4432
rect 11320 4388 11360 4600
rect 20140 4556 20180 4600
rect 30028 4556 30068 4600
rect 18799 4516 18808 4556
rect 18848 4516 18890 4556
rect 18930 4516 18972 4556
rect 19012 4516 19054 4556
rect 19094 4516 19136 4556
rect 19176 4516 19185 4556
rect 19555 4516 19564 4556
rect 19604 4516 20180 4556
rect 26563 4516 26572 4556
rect 26612 4516 28300 4556
rect 28340 4516 28349 4556
rect 30028 4516 31852 4556
rect 31892 4516 33292 4556
rect 33332 4516 33341 4556
rect 33919 4516 33928 4556
rect 33968 4516 34010 4556
rect 34050 4516 34092 4556
rect 34132 4516 34174 4556
rect 34214 4516 34256 4556
rect 34296 4516 34305 4556
rect 42928 4472 43008 4492
rect 12163 4432 12172 4472
rect 12212 4432 28396 4472
rect 28436 4432 28445 4472
rect 32227 4432 32236 4472
rect 32276 4432 40492 4472
rect 40532 4432 40541 4472
rect 40675 4432 40684 4472
rect 40724 4432 43008 4472
rect 42928 4412 43008 4432
rect 2755 4348 2764 4388
rect 2804 4348 11360 4388
rect 13795 4348 13804 4388
rect 13844 4348 23884 4388
rect 23924 4348 23933 4388
rect 28963 4348 28972 4388
rect 29012 4348 29164 4388
rect 29204 4348 29213 4388
rect 31555 4348 31564 4388
rect 31604 4348 32044 4388
rect 32084 4348 32093 4388
rect 4675 4304 4733 4305
rect 22627 4304 22685 4305
rect 4483 4264 4492 4304
rect 4532 4264 4684 4304
rect 4724 4264 4733 4304
rect 7075 4264 7084 4304
rect 7124 4264 7468 4304
rect 7508 4264 7517 4304
rect 7939 4264 7948 4304
rect 7988 4264 16876 4304
rect 16916 4264 16925 4304
rect 20140 4264 21868 4304
rect 21908 4264 21917 4304
rect 22627 4264 22636 4304
rect 22676 4264 38132 4304
rect 4675 4263 4733 4264
rect 3331 4180 3340 4220
rect 3380 4180 3532 4220
rect 3572 4180 4012 4220
rect 4052 4180 5068 4220
rect 5108 4180 7564 4220
rect 7604 4180 7613 4220
rect 11011 4180 11020 4220
rect 11060 4180 19372 4220
rect 19412 4180 19421 4220
rect 0 4136 80 4156
rect 4579 4136 4637 4137
rect 20140 4136 20180 4264
rect 22627 4263 22685 4264
rect 20323 4180 20332 4220
rect 20372 4180 21772 4220
rect 21812 4180 21821 4220
rect 23299 4180 23308 4220
rect 23348 4180 23788 4220
rect 23828 4180 23837 4220
rect 0 4096 4052 4136
rect 4099 4096 4108 4136
rect 4148 4096 4588 4136
rect 4628 4096 4637 4136
rect 4867 4096 4876 4136
rect 4916 4096 5452 4136
rect 5492 4096 5501 4136
rect 6499 4096 6508 4136
rect 6548 4096 6988 4136
rect 7028 4096 7037 4136
rect 10531 4096 10540 4136
rect 10580 4096 10924 4136
rect 10964 4096 10973 4136
rect 11491 4096 11500 4136
rect 11540 4096 13612 4136
rect 13652 4096 13661 4136
rect 19939 4096 19948 4136
rect 19988 4096 20180 4136
rect 0 4076 80 4096
rect 4012 4052 4052 4096
rect 4579 4095 4637 4096
rect 20332 4052 20372 4180
rect 38092 4136 38132 4264
rect 42928 4136 43008 4156
rect 24451 4096 24460 4136
rect 24500 4096 26476 4136
rect 26516 4096 26525 4136
rect 30595 4096 30604 4136
rect 30644 4096 30892 4136
rect 30932 4096 30941 4136
rect 32515 4096 32524 4136
rect 32564 4096 32573 4136
rect 33187 4096 33196 4136
rect 33236 4096 35500 4136
rect 35540 4096 35884 4136
rect 35924 4096 35933 4136
rect 37315 4096 37324 4136
rect 37364 4096 37900 4136
rect 37940 4096 37949 4136
rect 38083 4096 38092 4136
rect 38132 4096 38141 4136
rect 41443 4096 41452 4136
rect 41492 4096 43008 4136
rect 32524 4052 32564 4096
rect 42928 4076 43008 4096
rect 4012 4012 9100 4052
rect 9140 4012 9149 4052
rect 11299 4012 11308 4052
rect 11348 4012 13228 4052
rect 13268 4012 20372 4052
rect 24739 4012 24748 4052
rect 24788 4012 25132 4052
rect 25172 4012 25181 4052
rect 28003 4012 28012 4052
rect 28052 4012 37228 4052
rect 37268 4012 37277 4052
rect 34051 3968 34109 3969
rect 36835 3968 36893 3969
rect 2659 3928 2668 3968
rect 2708 3928 6220 3968
rect 6260 3928 6269 3968
rect 8611 3928 8620 3968
rect 8660 3928 17260 3968
rect 17300 3928 17309 3968
rect 30979 3928 30988 3968
rect 31028 3928 31852 3968
rect 31892 3928 31901 3968
rect 34051 3928 34060 3968
rect 34100 3928 34156 3968
rect 34196 3928 34205 3968
rect 36750 3928 36844 3968
rect 36884 3928 36893 3968
rect 34051 3927 34109 3928
rect 36835 3927 36893 3928
rect 4003 3844 4012 3884
rect 4052 3844 4532 3884
rect 12067 3844 12076 3884
rect 12116 3844 12556 3884
rect 12596 3844 27532 3884
rect 27572 3844 35596 3884
rect 35636 3844 35645 3884
rect 0 3800 80 3820
rect 4492 3800 4532 3844
rect 42928 3800 43008 3820
rect 0 3760 2764 3800
rect 2804 3760 2813 3800
rect 3043 3760 3052 3800
rect 3092 3760 4108 3800
rect 4148 3760 4157 3800
rect 4483 3760 4492 3800
rect 4532 3760 4541 3800
rect 4919 3760 4928 3800
rect 4968 3760 5010 3800
rect 5050 3760 5092 3800
rect 5132 3760 5174 3800
rect 5214 3760 5256 3800
rect 5296 3760 5305 3800
rect 7075 3760 7084 3800
rect 7124 3760 7756 3800
rect 7796 3760 7805 3800
rect 10243 3760 10252 3800
rect 10292 3760 15532 3800
rect 15572 3760 16204 3800
rect 16244 3760 16253 3800
rect 19267 3760 19276 3800
rect 19316 3760 19564 3800
rect 19604 3760 19613 3800
rect 20039 3760 20048 3800
rect 20088 3760 20130 3800
rect 20170 3760 20212 3800
rect 20252 3760 20294 3800
rect 20334 3760 20376 3800
rect 20416 3760 20425 3800
rect 30307 3760 30316 3800
rect 30356 3760 31564 3800
rect 31604 3760 31613 3800
rect 31939 3760 31948 3800
rect 31988 3760 32524 3800
rect 32564 3760 32573 3800
rect 35159 3760 35168 3800
rect 35208 3760 35250 3800
rect 35290 3760 35332 3800
rect 35372 3760 35414 3800
rect 35454 3760 35496 3800
rect 35536 3760 35545 3800
rect 36643 3760 36652 3800
rect 36692 3760 37516 3800
rect 37556 3760 38380 3800
rect 38420 3760 38668 3800
rect 38708 3760 38717 3800
rect 41059 3760 41068 3800
rect 41108 3760 43008 3800
rect 0 3740 80 3760
rect 42928 3740 43008 3760
rect 4579 3676 4588 3716
rect 4628 3676 5932 3716
rect 5972 3676 5981 3716
rect 13123 3676 13132 3716
rect 13172 3676 13708 3716
rect 13748 3676 13757 3716
rect 33091 3676 33100 3716
rect 33140 3676 35788 3716
rect 35828 3676 38284 3716
rect 38324 3676 38333 3716
rect 5539 3632 5597 3633
rect 3811 3592 3820 3632
rect 3860 3592 4876 3632
rect 4916 3592 4925 3632
rect 5059 3592 5068 3632
rect 5108 3592 5548 3632
rect 5588 3592 5597 3632
rect 9379 3592 9388 3632
rect 9428 3592 20812 3632
rect 20852 3592 20861 3632
rect 30595 3592 30604 3632
rect 30644 3592 32812 3632
rect 32852 3592 33772 3632
rect 33812 3592 33821 3632
rect 35587 3592 35596 3632
rect 35636 3592 40300 3632
rect 40340 3592 40876 3632
rect 40916 3592 40925 3632
rect 5539 3591 5597 3592
rect 3715 3508 3724 3548
rect 3764 3508 5740 3548
rect 5780 3508 5789 3548
rect 13516 3508 14284 3548
rect 14324 3508 15148 3548
rect 15188 3508 15628 3548
rect 15668 3508 16780 3548
rect 16820 3508 16829 3548
rect 23779 3508 23788 3548
rect 23828 3508 25996 3548
rect 26036 3508 26045 3548
rect 26467 3508 26476 3548
rect 26516 3508 27148 3548
rect 27188 3508 27436 3548
rect 27476 3508 28684 3548
rect 28724 3508 28733 3548
rect 29539 3508 29548 3548
rect 29588 3508 32716 3548
rect 32756 3508 35020 3548
rect 35060 3508 35404 3548
rect 35444 3508 35453 3548
rect 0 3464 80 3484
rect 12259 3464 12317 3465
rect 13516 3464 13556 3508
rect 13891 3464 13949 3465
rect 15523 3464 15581 3465
rect 42928 3464 43008 3484
rect 0 3424 2540 3464
rect 3043 3424 3052 3464
rect 3092 3424 3436 3464
rect 3476 3424 3820 3464
rect 3860 3424 3869 3464
rect 4099 3424 4108 3464
rect 4148 3424 5644 3464
rect 5684 3424 7372 3464
rect 7412 3424 7421 3464
rect 12174 3424 12268 3464
rect 12308 3424 12317 3464
rect 13507 3424 13516 3464
rect 13556 3424 13565 3464
rect 13806 3424 13900 3464
rect 13940 3424 13949 3464
rect 15438 3424 15532 3464
rect 15572 3424 15581 3464
rect 18307 3424 18316 3464
rect 18356 3424 20180 3464
rect 23203 3424 23212 3464
rect 23252 3424 23980 3464
rect 24020 3424 24029 3464
rect 25699 3424 25708 3464
rect 25748 3424 27628 3464
rect 27668 3424 27677 3464
rect 28579 3424 28588 3464
rect 28628 3424 29932 3464
rect 29972 3424 29981 3464
rect 30211 3424 30220 3464
rect 30260 3424 32236 3464
rect 32276 3424 33676 3464
rect 33716 3424 35980 3464
rect 36020 3424 36029 3464
rect 40675 3424 40684 3464
rect 40724 3424 43008 3464
rect 0 3404 80 3424
rect 2500 3212 2540 3424
rect 12259 3423 12317 3424
rect 13891 3423 13949 3424
rect 15523 3423 15581 3424
rect 12268 3380 12308 3423
rect 19939 3380 19997 3381
rect 20140 3380 20180 3424
rect 42928 3404 43008 3424
rect 3907 3340 3916 3380
rect 3956 3340 6028 3380
rect 6068 3340 6077 3380
rect 6595 3340 6604 3380
rect 6644 3340 12308 3380
rect 18115 3340 18124 3380
rect 18164 3340 19660 3380
rect 19700 3340 19709 3380
rect 19939 3340 19948 3380
rect 19988 3340 20044 3380
rect 20084 3340 20093 3380
rect 20140 3340 25900 3380
rect 25940 3340 25949 3380
rect 27235 3340 27244 3380
rect 27284 3340 28972 3380
rect 29012 3340 29021 3380
rect 29347 3340 29356 3380
rect 29396 3340 38764 3380
rect 38804 3340 40492 3380
rect 40532 3340 40541 3380
rect 19939 3339 19997 3340
rect 33676 3296 33716 3340
rect 3331 3256 3340 3296
rect 3380 3256 8908 3296
rect 8948 3256 8957 3296
rect 15907 3256 15916 3296
rect 15956 3256 16588 3296
rect 16628 3256 20908 3296
rect 20948 3256 24940 3296
rect 24980 3256 24989 3296
rect 30499 3256 30508 3296
rect 30548 3256 30988 3296
rect 31028 3256 31037 3296
rect 33667 3256 33676 3296
rect 33716 3256 33725 3296
rect 4099 3212 4157 3213
rect 2500 3172 3572 3212
rect 4014 3172 4108 3212
rect 4148 3172 4157 3212
rect 0 3128 80 3148
rect 0 3088 3476 3128
rect 0 3068 80 3088
rect 0 2792 80 2812
rect 3436 2792 3476 3088
rect 3532 2876 3572 3172
rect 4099 3171 4157 3172
rect 4579 3212 4637 3213
rect 28771 3212 28829 3213
rect 4579 3172 4588 3212
rect 4628 3172 5164 3212
rect 5204 3172 5213 3212
rect 7459 3172 7468 3212
rect 7508 3172 18316 3212
rect 18356 3172 18365 3212
rect 20140 3172 20332 3212
rect 20372 3172 25612 3212
rect 25652 3172 25661 3212
rect 28686 3172 28780 3212
rect 28820 3172 28829 3212
rect 4579 3171 4637 3172
rect 4771 3128 4829 3129
rect 20140 3128 20180 3172
rect 28771 3171 28829 3172
rect 42928 3128 43008 3148
rect 4771 3088 4780 3128
rect 4820 3088 11020 3128
rect 11060 3088 11069 3128
rect 11212 3088 15628 3128
rect 15668 3088 15677 3128
rect 16003 3088 16012 3128
rect 16052 3088 16684 3128
rect 16724 3088 20180 3128
rect 20707 3088 20716 3128
rect 20756 3088 23308 3128
rect 23348 3088 23357 3128
rect 41059 3088 41068 3128
rect 41108 3088 43008 3128
rect 4771 3087 4829 3088
rect 11212 3044 11252 3088
rect 42928 3068 43008 3088
rect 3679 3004 3688 3044
rect 3728 3004 3770 3044
rect 3810 3004 3852 3044
rect 3892 3004 3934 3044
rect 3974 3004 4016 3044
rect 4056 3004 4065 3044
rect 7747 3004 7756 3044
rect 7796 3004 11252 3044
rect 18799 3004 18808 3044
rect 18848 3004 18890 3044
rect 18930 3004 18972 3044
rect 19012 3004 19054 3044
rect 19094 3004 19136 3044
rect 19176 3004 19185 3044
rect 20803 3004 20812 3044
rect 20852 3004 24652 3044
rect 24692 3004 24701 3044
rect 33919 3004 33928 3044
rect 33968 3004 34010 3044
rect 34050 3004 34092 3044
rect 34132 3004 34174 3044
rect 34214 3004 34256 3044
rect 34296 3004 34305 3044
rect 4291 2960 4349 2961
rect 4291 2920 4300 2960
rect 4340 2920 4396 2960
rect 4436 2920 4445 2960
rect 10339 2920 10348 2960
rect 10388 2920 11212 2960
rect 11252 2920 11261 2960
rect 15427 2920 15436 2960
rect 15476 2920 22060 2960
rect 22100 2920 22109 2960
rect 24931 2920 24940 2960
rect 24980 2920 25612 2960
rect 25652 2920 25661 2960
rect 27523 2920 27532 2960
rect 27572 2920 41260 2960
rect 41300 2920 41309 2960
rect 4291 2919 4349 2920
rect 3532 2836 11404 2876
rect 11444 2836 11453 2876
rect 16195 2836 16204 2876
rect 16244 2836 20180 2876
rect 20515 2836 20524 2876
rect 20564 2836 21292 2876
rect 21332 2836 23212 2876
rect 23252 2836 23261 2876
rect 28579 2836 28588 2876
rect 28628 2836 31372 2876
rect 31412 2836 31421 2876
rect 32611 2836 32620 2876
rect 32660 2836 32908 2876
rect 32948 2836 32957 2876
rect 36547 2836 36556 2876
rect 36596 2836 36940 2876
rect 36980 2836 36989 2876
rect 37795 2836 37804 2876
rect 37844 2836 38572 2876
rect 38612 2836 38621 2876
rect 20140 2792 20180 2836
rect 21379 2792 21437 2793
rect 42928 2792 43008 2812
rect 0 2752 3340 2792
rect 3380 2752 3389 2792
rect 3436 2752 10444 2792
rect 10484 2752 10493 2792
rect 10540 2752 13804 2792
rect 13844 2752 13853 2792
rect 19459 2752 19468 2792
rect 19508 2752 20044 2792
rect 20084 2752 20093 2792
rect 20140 2752 20812 2792
rect 20852 2752 20861 2792
rect 21294 2752 21388 2792
rect 21428 2752 21437 2792
rect 23299 2752 23308 2792
rect 23348 2752 24172 2792
rect 24212 2752 24940 2792
rect 24980 2752 24989 2792
rect 40675 2752 40684 2792
rect 40724 2752 43008 2792
rect 0 2732 80 2752
rect 10540 2708 10580 2752
rect 21379 2751 21437 2752
rect 42928 2732 43008 2752
rect 3427 2668 3436 2708
rect 3476 2668 4972 2708
rect 5012 2668 5548 2708
rect 5588 2668 5597 2708
rect 9091 2668 9100 2708
rect 9140 2668 10580 2708
rect 11203 2668 11212 2708
rect 11252 2668 12268 2708
rect 12308 2668 12317 2708
rect 13027 2668 13036 2708
rect 13076 2668 24460 2708
rect 24500 2668 24509 2708
rect 25891 2668 25900 2708
rect 25940 2668 29644 2708
rect 29684 2668 37820 2708
rect 4675 2624 4733 2625
rect 3715 2584 3724 2624
rect 3764 2584 4492 2624
rect 4532 2584 4541 2624
rect 4675 2584 4684 2624
rect 4724 2584 4876 2624
rect 4916 2584 4925 2624
rect 5635 2584 5644 2624
rect 5684 2584 7852 2624
rect 7892 2584 7901 2624
rect 8899 2584 8908 2624
rect 8948 2584 14380 2624
rect 14420 2584 14429 2624
rect 18019 2584 18028 2624
rect 18068 2584 18077 2624
rect 18403 2584 18412 2624
rect 18452 2584 23692 2624
rect 23732 2584 23741 2624
rect 24643 2584 24652 2624
rect 24692 2584 27916 2624
rect 27956 2584 27965 2624
rect 28291 2584 28300 2624
rect 28340 2584 31756 2624
rect 31796 2584 31805 2624
rect 33283 2584 33292 2624
rect 33332 2584 34924 2624
rect 34964 2584 36748 2624
rect 36788 2584 36797 2624
rect 4675 2583 4733 2584
rect 18028 2541 18068 2584
rect 18019 2540 18077 2541
rect 21379 2540 21437 2541
rect 18019 2500 18028 2540
rect 18068 2500 18079 2540
rect 20035 2500 20044 2540
rect 20084 2500 20276 2540
rect 21348 2500 21388 2540
rect 21428 2500 21437 2540
rect 37780 2540 37820 2668
rect 37780 2500 40780 2540
rect 40820 2500 40829 2540
rect 18019 2499 18077 2500
rect 0 2456 80 2476
rect 20236 2456 20276 2500
rect 21379 2499 21437 2500
rect 21388 2456 21428 2499
rect 42928 2456 43008 2476
rect 0 2416 7276 2456
rect 7316 2416 7325 2456
rect 11395 2416 11404 2456
rect 11444 2416 20180 2456
rect 20236 2416 21428 2456
rect 23212 2416 29356 2456
rect 29396 2416 29405 2456
rect 34819 2416 34828 2456
rect 34868 2416 35308 2456
rect 35348 2416 35357 2456
rect 41443 2416 41452 2456
rect 41492 2416 43008 2456
rect 0 2396 80 2416
rect 20140 2372 20180 2416
rect 23212 2372 23252 2416
rect 42928 2396 43008 2416
rect 20140 2332 23252 2372
rect 24547 2332 24556 2372
rect 24596 2332 40876 2372
rect 40916 2332 40925 2372
rect 4195 2248 4204 2288
rect 4244 2248 4588 2288
rect 4628 2248 4637 2288
rect 4919 2248 4928 2288
rect 4968 2248 5010 2288
rect 5050 2248 5092 2288
rect 5132 2248 5174 2288
rect 5214 2248 5256 2288
rect 5296 2248 5305 2288
rect 5356 2248 5740 2288
rect 5780 2248 5789 2288
rect 20039 2248 20048 2288
rect 20088 2248 20130 2288
rect 20170 2248 20212 2288
rect 20252 2248 20294 2288
rect 20334 2248 20376 2288
rect 20416 2248 20425 2288
rect 21187 2248 21196 2288
rect 21236 2248 21388 2288
rect 21428 2248 22580 2288
rect 35159 2248 35168 2288
rect 35208 2248 35250 2288
rect 35290 2248 35332 2288
rect 35372 2248 35414 2288
rect 35454 2248 35496 2288
rect 35536 2248 35545 2288
rect 40483 2248 40492 2288
rect 40532 2248 40541 2288
rect 5356 2204 5396 2248
rect 3139 2164 3148 2204
rect 3188 2164 3532 2204
rect 3572 2164 5396 2204
rect 5443 2164 5452 2204
rect 5492 2164 8812 2204
rect 8852 2164 8861 2204
rect 14371 2164 14380 2204
rect 14420 2164 21332 2204
rect 0 2120 80 2140
rect 0 2080 6412 2120
rect 6452 2080 7468 2120
rect 7508 2080 7517 2120
rect 11011 2080 11020 2120
rect 11060 2080 15436 2120
rect 15476 2080 15485 2120
rect 20035 2080 20044 2120
rect 20084 2080 20140 2120
rect 20180 2080 20208 2120
rect 0 2060 80 2080
rect 21292 2036 21332 2164
rect 22540 2120 22580 2248
rect 29539 2164 29548 2204
rect 29588 2164 37132 2204
rect 37172 2164 37181 2204
rect 30787 2120 30845 2121
rect 40492 2120 40532 2248
rect 42928 2120 43008 2140
rect 22531 2080 22540 2120
rect 22580 2080 22828 2120
rect 22868 2080 24172 2120
rect 24212 2080 26476 2120
rect 26516 2080 26525 2120
rect 30787 2080 30796 2120
rect 30836 2080 31180 2120
rect 31220 2080 31229 2120
rect 34444 2080 40532 2120
rect 41059 2080 41068 2120
rect 41108 2080 43008 2120
rect 30787 2079 30845 2080
rect 34444 2036 34484 2080
rect 42928 2060 43008 2080
rect 34627 2036 34685 2037
rect 5059 1996 5068 2036
rect 5108 1996 5548 2036
rect 5588 1996 5597 2036
rect 5731 1996 5740 2036
rect 5780 1996 6320 2036
rect 15043 1996 15052 2036
rect 15092 1996 16684 2036
rect 16724 1996 16733 2036
rect 21283 1996 21292 2036
rect 21332 1996 26188 2036
rect 26228 1996 34484 2036
rect 34542 1996 34636 2036
rect 34676 1996 34685 2036
rect 6280 1952 6320 1996
rect 34627 1995 34685 1996
rect 29539 1952 29597 1953
rect 3907 1912 3916 1952
rect 3956 1912 5356 1952
rect 5396 1912 5405 1952
rect 6280 1912 6508 1952
rect 6548 1912 7756 1952
rect 7796 1912 7805 1952
rect 8515 1912 8524 1952
rect 8564 1912 10156 1952
rect 10196 1912 10205 1952
rect 10531 1912 10540 1952
rect 10580 1912 16300 1952
rect 16340 1912 22924 1952
rect 22964 1912 24556 1952
rect 24596 1912 24605 1952
rect 24931 1912 24940 1952
rect 24980 1912 25804 1952
rect 25844 1912 26668 1952
rect 26708 1912 27436 1952
rect 27476 1912 28492 1952
rect 28532 1912 28876 1952
rect 28916 1912 28925 1952
rect 29454 1912 29548 1952
rect 29588 1912 29597 1952
rect 30883 1912 30892 1952
rect 30932 1912 33388 1952
rect 33428 1912 33437 1952
rect 37123 1912 37132 1952
rect 37172 1912 40492 1952
rect 40532 1912 40541 1952
rect 10156 1868 10196 1912
rect 29539 1911 29597 1912
rect 1795 1828 1804 1868
rect 1844 1828 9484 1868
rect 9524 1828 9533 1868
rect 10156 1828 10636 1868
rect 10676 1828 11788 1868
rect 11828 1828 12652 1868
rect 12692 1828 13420 1868
rect 13460 1828 15052 1868
rect 15092 1828 15101 1868
rect 20131 1828 20140 1868
rect 20180 1828 27532 1868
rect 27572 1828 27916 1868
rect 27956 1828 27965 1868
rect 28099 1828 28108 1868
rect 28148 1828 40012 1868
rect 40052 1828 40061 1868
rect 0 1784 80 1804
rect 9763 1784 9821 1785
rect 42928 1784 43008 1804
rect 0 1744 9772 1784
rect 9812 1744 9821 1784
rect 16675 1744 16684 1784
rect 16724 1744 21772 1784
rect 21812 1744 21821 1784
rect 26467 1744 26476 1784
rect 26516 1744 36268 1784
rect 36308 1744 39628 1784
rect 39668 1744 39677 1784
rect 41443 1744 41452 1784
rect 41492 1744 43008 1784
rect 0 1724 80 1744
rect 9763 1743 9821 1744
rect 42928 1724 43008 1744
rect 33187 1700 33245 1701
rect 3331 1660 3340 1700
rect 3380 1660 3820 1700
rect 3860 1660 4300 1700
rect 4340 1660 4349 1700
rect 7267 1660 7276 1700
rect 7316 1660 20044 1700
rect 20084 1660 20093 1700
rect 23779 1660 23788 1700
rect 23828 1660 31372 1700
rect 31412 1660 31421 1700
rect 33187 1660 33196 1700
rect 33236 1660 38188 1700
rect 38228 1660 38237 1700
rect 33187 1659 33245 1660
rect 4483 1616 4541 1617
rect 4387 1576 4396 1616
rect 4436 1576 4492 1616
rect 4532 1576 4541 1616
rect 7747 1576 7756 1616
rect 7796 1576 8524 1616
rect 8564 1576 8573 1616
rect 21667 1576 21676 1616
rect 21716 1576 28108 1616
rect 28148 1576 28157 1616
rect 28867 1576 28876 1616
rect 28916 1576 29164 1616
rect 29204 1576 30796 1616
rect 30836 1576 30845 1616
rect 4483 1575 4541 1576
rect 3679 1492 3688 1532
rect 3728 1492 3770 1532
rect 3810 1492 3852 1532
rect 3892 1492 3934 1532
rect 3974 1492 4016 1532
rect 4056 1492 4065 1532
rect 18799 1492 18808 1532
rect 18848 1492 18890 1532
rect 18930 1492 18972 1532
rect 19012 1492 19054 1532
rect 19094 1492 19136 1532
rect 19176 1492 19185 1532
rect 33919 1492 33928 1532
rect 33968 1492 34010 1532
rect 34050 1492 34092 1532
rect 34132 1492 34174 1532
rect 34214 1492 34256 1532
rect 34296 1492 34305 1532
rect 0 1448 80 1468
rect 32995 1448 33053 1449
rect 42928 1448 43008 1468
rect 0 1408 212 1448
rect 21763 1408 21772 1448
rect 21812 1408 22540 1448
rect 22580 1408 22589 1448
rect 32995 1408 33004 1448
rect 33044 1408 37612 1448
rect 37652 1408 37661 1448
rect 39811 1408 39820 1448
rect 39860 1408 43008 1448
rect 0 1388 80 1408
rect 172 1280 212 1408
rect 32995 1407 33053 1408
rect 42928 1388 43008 1408
rect 35587 1280 35645 1281
rect 172 1240 8180 1280
rect 9379 1240 9388 1280
rect 9428 1240 10252 1280
rect 10292 1240 11020 1280
rect 11060 1240 11069 1280
rect 17539 1240 17548 1280
rect 17588 1240 17932 1280
rect 17972 1240 17981 1280
rect 19075 1240 19084 1280
rect 19124 1240 19276 1280
rect 19316 1240 19660 1280
rect 19700 1240 21292 1280
rect 21332 1240 21341 1280
rect 23683 1240 23692 1280
rect 23732 1240 26476 1280
rect 26516 1240 26525 1280
rect 30115 1240 30124 1280
rect 30164 1240 31660 1280
rect 31700 1240 31709 1280
rect 32323 1240 32332 1280
rect 32372 1240 33484 1280
rect 33524 1240 33533 1280
rect 35502 1240 35596 1280
rect 35636 1240 41164 1280
rect 41204 1240 41213 1280
rect 8140 1196 8180 1240
rect 23692 1196 23732 1240
rect 35587 1239 35645 1240
rect 25411 1196 25469 1197
rect 40867 1196 40925 1197
rect 76 1156 212 1196
rect 4387 1156 4396 1196
rect 4436 1156 5068 1196
rect 5108 1156 5117 1196
rect 8131 1156 8140 1196
rect 8180 1156 23732 1196
rect 25326 1156 25420 1196
rect 25460 1156 25469 1196
rect 27619 1156 27628 1196
rect 27668 1156 31316 1196
rect 31747 1156 31756 1196
rect 31796 1156 33676 1196
rect 33716 1156 33725 1196
rect 36355 1156 36364 1196
rect 36404 1156 37420 1196
rect 37460 1156 37469 1196
rect 40782 1156 40876 1196
rect 40916 1156 40925 1196
rect 76 1132 116 1156
rect 0 1072 116 1132
rect 0 1052 80 1072
rect 172 860 212 1156
rect 25411 1155 25469 1156
rect 2467 1112 2525 1113
rect 31276 1112 31316 1156
rect 40867 1155 40925 1156
rect 42928 1112 43008 1132
rect 2382 1072 2476 1112
rect 2516 1072 2525 1112
rect 4099 1072 4108 1112
rect 4148 1072 4780 1112
rect 4820 1072 4829 1112
rect 8707 1072 8716 1112
rect 8756 1072 9868 1112
rect 9908 1072 9917 1112
rect 12355 1072 12364 1112
rect 12404 1072 14668 1112
rect 14708 1072 14717 1112
rect 15619 1072 15628 1112
rect 15668 1072 17548 1112
rect 17588 1072 17597 1112
rect 17923 1072 17932 1112
rect 17972 1072 24844 1112
rect 24884 1072 31180 1112
rect 31220 1072 31229 1112
rect 31276 1072 37900 1112
rect 37940 1072 37949 1112
rect 40675 1072 40684 1112
rect 40724 1072 43008 1112
rect 2467 1071 2525 1072
rect 37900 1028 37940 1072
rect 42928 1052 43008 1072
rect 3907 988 3916 1028
rect 3956 988 4684 1028
rect 4724 988 4733 1028
rect 5347 988 5356 1028
rect 5396 988 13036 1028
rect 13076 988 13085 1028
rect 13315 988 13324 1028
rect 13364 988 36404 1028
rect 37900 988 41260 1028
rect 41300 988 41309 1028
rect 6403 944 6461 945
rect 9763 944 9821 945
rect 35011 944 35069 945
rect 4099 904 4108 944
rect 4148 904 4972 944
rect 5012 904 5021 944
rect 6318 904 6412 944
rect 6452 904 6461 944
rect 7939 904 7948 944
rect 7988 904 8716 944
rect 8756 904 8765 944
rect 9678 904 9772 944
rect 9812 904 9821 944
rect 13603 904 13612 944
rect 13652 904 14476 944
rect 14516 904 14525 944
rect 14659 904 14668 944
rect 14708 904 24116 944
rect 25987 904 25996 944
rect 26036 904 28588 944
rect 28628 904 28637 944
rect 31459 904 31468 944
rect 31508 904 32332 944
rect 32372 904 32381 944
rect 32428 904 34636 944
rect 34676 904 34685 944
rect 34926 904 35020 944
rect 35060 904 35069 944
rect 36364 944 36404 988
rect 36364 904 39916 944
rect 39956 904 39965 944
rect 6403 903 6461 904
rect 9763 903 9821 904
rect 18019 860 18077 861
rect 172 820 18028 860
rect 18068 820 18077 860
rect 18403 820 18412 860
rect 18452 820 23924 860
rect 18019 819 18077 820
rect 0 776 80 796
rect 0 736 212 776
rect 4919 736 4928 776
rect 4968 736 5010 776
rect 5050 736 5092 776
rect 5132 736 5174 776
rect 5214 736 5256 776
rect 5296 736 5305 776
rect 17539 736 17548 776
rect 17588 736 19084 776
rect 19124 736 19133 776
rect 20039 736 20048 776
rect 20088 736 20130 776
rect 20170 736 20212 776
rect 20252 736 20294 776
rect 20334 736 20376 776
rect 20416 736 20425 776
rect 0 716 80 736
rect 172 608 212 736
rect 13027 652 13036 692
rect 13076 652 21676 692
rect 21716 652 21725 692
rect 23884 608 23924 820
rect 24076 776 24116 904
rect 32428 860 32468 904
rect 35011 903 35069 904
rect 32131 820 32140 860
rect 32180 820 32468 860
rect 32611 820 32620 860
rect 32660 820 34156 860
rect 34196 820 34205 860
rect 42928 776 43008 796
rect 24076 736 28012 776
rect 28052 736 28061 776
rect 29443 736 29452 776
rect 29492 736 32812 776
rect 32852 736 32861 776
rect 35159 736 35168 776
rect 35208 736 35250 776
rect 35290 736 35332 776
rect 35372 736 35414 776
rect 35454 736 35496 776
rect 35536 736 35545 776
rect 41443 736 41452 776
rect 41492 736 43008 776
rect 42928 716 43008 736
rect 27139 652 27148 692
rect 27188 652 32524 692
rect 32564 652 32573 692
rect 32899 652 32908 692
rect 32948 652 34444 692
rect 34484 652 34493 692
rect 172 568 18412 608
rect 18452 568 18461 608
rect 23884 568 27628 608
rect 27668 568 27677 608
rect 30595 568 30604 608
rect 30644 568 33292 608
rect 33332 568 33341 608
rect 34051 568 34060 608
rect 34100 568 34828 608
rect 34868 568 34877 608
rect 24835 484 24844 524
rect 24884 484 31564 524
rect 31604 484 31613 524
rect 0 440 80 460
rect 42928 440 43008 460
rect 0 400 5356 440
rect 5396 400 5405 440
rect 40195 400 40204 440
rect 40244 400 43008 440
rect 0 380 80 400
rect 42928 380 43008 400
rect 41059 148 41068 188
rect 41108 148 41600 188
rect 0 104 80 124
rect 41560 104 41600 148
rect 42928 104 43008 124
rect 0 64 6604 104
rect 6644 64 6653 104
rect 10339 64 10348 104
rect 10388 64 11020 104
rect 11060 64 11069 104
rect 12835 64 12844 104
rect 12884 64 13324 104
rect 13364 64 13373 104
rect 15331 64 15340 104
rect 15380 64 15628 104
rect 15668 64 15677 104
rect 20227 64 20236 104
rect 20276 64 20428 104
rect 20468 64 20477 104
rect 34915 64 34924 104
rect 34964 64 35212 104
rect 35252 64 35261 104
rect 37507 64 37516 104
rect 37556 64 37804 104
rect 37844 64 37853 104
rect 39619 64 39628 104
rect 39668 64 39820 104
rect 39860 64 39869 104
rect 40771 64 40780 104
rect 40820 64 40972 104
rect 41012 64 41021 104
rect 41560 64 43008 104
rect 0 44 80 64
rect 42928 44 43008 64
<< via3 >>
rect 20620 10648 20660 10688
rect 4588 10480 4628 10520
rect 16972 10480 17012 10520
rect 18700 10480 18740 10520
rect 21100 10228 21140 10268
rect 16396 9976 16436 10016
rect 1612 9808 1652 9848
rect 4928 9808 4968 9848
rect 5010 9808 5050 9848
rect 5092 9808 5132 9848
rect 5174 9808 5214 9848
rect 5256 9808 5296 9848
rect 20048 9808 20088 9848
rect 20130 9808 20170 9848
rect 20212 9808 20252 9848
rect 20294 9808 20334 9848
rect 20376 9808 20416 9848
rect 35168 9808 35208 9848
rect 35250 9808 35290 9848
rect 35332 9808 35372 9848
rect 35414 9808 35454 9848
rect 35496 9808 35536 9848
rect 12652 9640 12692 9680
rect 15244 9640 15284 9680
rect 16396 9556 16436 9596
rect 22636 9556 22676 9596
rect 5452 9472 5492 9512
rect 7564 9388 7604 9428
rect 10348 9388 10388 9428
rect 22828 9472 22868 9512
rect 40876 9388 40916 9428
rect 37612 9220 37652 9260
rect 14188 9136 14228 9176
rect 3688 9052 3728 9092
rect 3770 9052 3810 9092
rect 3852 9052 3892 9092
rect 3934 9052 3974 9092
rect 4016 9052 4056 9092
rect 18808 9052 18848 9092
rect 18890 9052 18930 9092
rect 18972 9052 19012 9092
rect 19054 9052 19094 9092
rect 19136 9052 19176 9092
rect 22732 9052 22772 9092
rect 26284 9052 26324 9092
rect 33928 9052 33968 9092
rect 34010 9052 34050 9092
rect 34092 9052 34132 9092
rect 34174 9052 34214 9092
rect 34256 9052 34296 9092
rect 10252 8800 10292 8840
rect 11020 8800 11060 8840
rect 11788 8800 11828 8840
rect 12556 8800 12596 8840
rect 14092 8800 14132 8840
rect 14476 8800 14516 8840
rect 15436 8800 15476 8840
rect 15628 8800 15668 8840
rect 16012 8800 16052 8840
rect 16780 8800 16820 8840
rect 18124 8800 18164 8840
rect 22252 8800 22292 8840
rect 33772 8800 33812 8840
rect 11404 8716 11444 8756
rect 3724 8632 3764 8672
rect 8812 8632 8852 8672
rect 9772 8632 9812 8672
rect 33196 8716 33236 8756
rect 13036 8632 13076 8672
rect 14860 8632 14900 8672
rect 15820 8632 15860 8672
rect 5548 8464 5588 8504
rect 13996 8464 14036 8504
rect 18892 8464 18932 8504
rect 19468 8632 19508 8672
rect 30796 8548 30836 8588
rect 27724 8464 27764 8504
rect 27916 8464 27956 8504
rect 30988 8464 31028 8504
rect 31372 8464 31412 8504
rect 31756 8464 31796 8504
rect 39724 8464 39764 8504
rect 33004 8380 33044 8420
rect 4108 8296 4148 8336
rect 4928 8296 4968 8336
rect 5010 8296 5050 8336
rect 5092 8296 5132 8336
rect 5174 8296 5214 8336
rect 5256 8296 5296 8336
rect 19468 8296 19508 8336
rect 20048 8296 20088 8336
rect 20130 8296 20170 8336
rect 20212 8296 20252 8336
rect 20294 8296 20334 8336
rect 20376 8296 20416 8336
rect 20620 8296 20660 8336
rect 6604 8212 6644 8252
rect 23308 8212 23348 8252
rect 26860 8212 26900 8252
rect 33100 8128 33140 8168
rect 11404 8044 11444 8084
rect 35168 8296 35208 8336
rect 35250 8296 35290 8336
rect 35332 8296 35372 8336
rect 35414 8296 35454 8336
rect 35496 8296 35536 8336
rect 6412 7960 6452 8000
rect 12364 7960 12404 8000
rect 22252 7960 22292 8000
rect 28012 7960 28052 8000
rect 28876 7960 28916 8000
rect 6028 7876 6068 7916
rect 23884 7876 23924 7916
rect 24076 7876 24116 7916
rect 1900 7792 1940 7832
rect 5452 7792 5492 7832
rect 28588 7792 28628 7832
rect 5740 7708 5780 7748
rect 20716 7708 20756 7748
rect 31372 7708 31412 7748
rect 32620 7708 32660 7748
rect 34636 7624 34676 7664
rect 3688 7540 3728 7580
rect 3770 7540 3810 7580
rect 3852 7540 3892 7580
rect 3934 7540 3974 7580
rect 4016 7540 4056 7580
rect 12076 7540 12116 7580
rect 18808 7540 18848 7580
rect 18890 7540 18930 7580
rect 18972 7540 19012 7580
rect 19054 7540 19094 7580
rect 19136 7540 19176 7580
rect 33928 7540 33968 7580
rect 34010 7540 34050 7580
rect 34092 7540 34132 7580
rect 34174 7540 34214 7580
rect 34256 7540 34296 7580
rect 2476 7456 2516 7496
rect 11500 7372 11540 7412
rect 35020 7372 35060 7412
rect 26284 7288 26324 7328
rect 26860 7288 26900 7328
rect 4588 7204 4628 7244
rect 31948 7288 31988 7328
rect 40300 7204 40340 7244
rect 4108 7120 4148 7160
rect 5356 7120 5396 7160
rect 8044 7120 8084 7160
rect 17644 7120 17684 7160
rect 19372 7120 19412 7160
rect 27820 7120 27860 7160
rect 28972 7036 29012 7076
rect 13804 6952 13844 6992
rect 29548 6952 29588 6992
rect 11500 6868 11540 6908
rect 4928 6784 4968 6824
rect 5010 6784 5050 6824
rect 5092 6784 5132 6824
rect 5174 6784 5214 6824
rect 5256 6784 5296 6824
rect 20048 6784 20088 6824
rect 20130 6784 20170 6824
rect 20212 6784 20252 6824
rect 20294 6784 20334 6824
rect 20376 6784 20416 6824
rect 35168 6784 35208 6824
rect 35250 6784 35290 6824
rect 35332 6784 35372 6824
rect 35414 6784 35454 6824
rect 35496 6784 35536 6824
rect 7180 6700 7220 6740
rect 30220 6700 30260 6740
rect 21676 6616 21716 6656
rect 5548 6448 5588 6488
rect 21676 6448 21716 6488
rect 6028 6364 6068 6404
rect 10732 6364 10772 6404
rect 33388 6448 33428 6488
rect 28972 6364 29012 6404
rect 41260 6364 41300 6404
rect 1612 6280 1652 6320
rect 1900 6280 1940 6320
rect 35692 6280 35732 6320
rect 40204 6280 40244 6320
rect 4684 6196 4724 6236
rect 1708 6112 1748 6152
rect 4300 6112 4340 6152
rect 6604 6112 6644 6152
rect 3688 6028 3728 6068
rect 3770 6028 3810 6068
rect 3852 6028 3892 6068
rect 3934 6028 3974 6068
rect 4016 6028 4056 6068
rect 14860 6028 14900 6068
rect 18808 6028 18848 6068
rect 18890 6028 18930 6068
rect 18972 6028 19012 6068
rect 19054 6028 19094 6068
rect 19136 6028 19176 6068
rect 4396 5944 4436 5984
rect 7180 5944 7220 5984
rect 27820 5944 27860 5984
rect 28972 5944 29012 5984
rect 21676 5860 21716 5900
rect 33928 6028 33968 6068
rect 34010 6028 34050 6068
rect 34092 6028 34132 6068
rect 34174 6028 34214 6068
rect 34256 6028 34296 6068
rect 4204 5776 4244 5816
rect 21100 5776 21140 5816
rect 29068 5776 29108 5816
rect 20620 5692 20660 5732
rect 23308 5692 23348 5732
rect 4108 5608 4148 5648
rect 5740 5608 5780 5648
rect 6028 5608 6068 5648
rect 16108 5608 16148 5648
rect 25804 5608 25844 5648
rect 5260 5440 5300 5480
rect 28300 5440 28340 5480
rect 4928 5272 4968 5312
rect 5010 5272 5050 5312
rect 5092 5272 5132 5312
rect 5174 5272 5214 5312
rect 5256 5272 5296 5312
rect 20048 5272 20088 5312
rect 20130 5272 20170 5312
rect 20212 5272 20252 5312
rect 20294 5272 20334 5312
rect 20376 5272 20416 5312
rect 33100 5272 33140 5312
rect 35168 5272 35208 5312
rect 35250 5272 35290 5312
rect 35332 5272 35372 5312
rect 35414 5272 35454 5312
rect 35496 5272 35536 5312
rect 1708 4936 1748 4976
rect 5356 4936 5396 4976
rect 15532 4936 15572 4976
rect 1228 4768 1268 4808
rect 4204 4768 4244 4808
rect 36652 4768 36692 4808
rect 40492 4684 40532 4724
rect 4396 4600 4436 4640
rect 3688 4516 3728 4556
rect 3770 4516 3810 4556
rect 3852 4516 3892 4556
rect 3934 4516 3974 4556
rect 4016 4516 4056 4556
rect 4780 4432 4820 4472
rect 18808 4516 18848 4556
rect 18890 4516 18930 4556
rect 18972 4516 19012 4556
rect 19054 4516 19094 4556
rect 19136 4516 19176 4556
rect 33928 4516 33968 4556
rect 34010 4516 34050 4556
rect 34092 4516 34132 4556
rect 34174 4516 34214 4556
rect 34256 4516 34296 4556
rect 4684 4264 4724 4304
rect 22636 4264 22676 4304
rect 4588 4096 4628 4136
rect 34060 3928 34100 3968
rect 36844 3928 36884 3968
rect 4928 3760 4968 3800
rect 5010 3760 5050 3800
rect 5092 3760 5132 3800
rect 5174 3760 5214 3800
rect 5256 3760 5296 3800
rect 20048 3760 20088 3800
rect 20130 3760 20170 3800
rect 20212 3760 20252 3800
rect 20294 3760 20334 3800
rect 20376 3760 20416 3800
rect 35168 3760 35208 3800
rect 35250 3760 35290 3800
rect 35332 3760 35372 3800
rect 35414 3760 35454 3800
rect 35496 3760 35536 3800
rect 5548 3592 5588 3632
rect 12268 3424 12308 3464
rect 13900 3424 13940 3464
rect 15532 3424 15572 3464
rect 19948 3340 19988 3380
rect 4108 3172 4148 3212
rect 4588 3172 4628 3212
rect 28780 3172 28820 3212
rect 4780 3088 4820 3128
rect 3688 3004 3728 3044
rect 3770 3004 3810 3044
rect 3852 3004 3892 3044
rect 3934 3004 3974 3044
rect 4016 3004 4056 3044
rect 18808 3004 18848 3044
rect 18890 3004 18930 3044
rect 18972 3004 19012 3044
rect 19054 3004 19094 3044
rect 19136 3004 19176 3044
rect 33928 3004 33968 3044
rect 34010 3004 34050 3044
rect 34092 3004 34132 3044
rect 34174 3004 34214 3044
rect 34256 3004 34296 3044
rect 4300 2920 4340 2960
rect 21388 2752 21428 2792
rect 4684 2584 4724 2624
rect 18028 2500 18068 2540
rect 21388 2500 21428 2540
rect 4928 2248 4968 2288
rect 5010 2248 5050 2288
rect 5092 2248 5132 2288
rect 5174 2248 5214 2288
rect 5256 2248 5296 2288
rect 20048 2248 20088 2288
rect 20130 2248 20170 2288
rect 20212 2248 20252 2288
rect 20294 2248 20334 2288
rect 20376 2248 20416 2288
rect 35168 2248 35208 2288
rect 35250 2248 35290 2288
rect 35332 2248 35372 2288
rect 35414 2248 35454 2288
rect 35496 2248 35536 2288
rect 30796 2080 30836 2120
rect 34636 1996 34676 2036
rect 29548 1912 29588 1952
rect 9772 1744 9812 1784
rect 33196 1660 33236 1700
rect 4492 1576 4532 1616
rect 3688 1492 3728 1532
rect 3770 1492 3810 1532
rect 3852 1492 3892 1532
rect 3934 1492 3974 1532
rect 4016 1492 4056 1532
rect 18808 1492 18848 1532
rect 18890 1492 18930 1532
rect 18972 1492 19012 1532
rect 19054 1492 19094 1532
rect 19136 1492 19176 1532
rect 33928 1492 33968 1532
rect 34010 1492 34050 1532
rect 34092 1492 34132 1532
rect 34174 1492 34214 1532
rect 34256 1492 34296 1532
rect 33004 1408 33044 1448
rect 35596 1240 35636 1280
rect 25420 1156 25460 1196
rect 40876 1156 40916 1196
rect 2476 1072 2516 1112
rect 6412 904 6452 944
rect 9772 904 9812 944
rect 35020 904 35060 944
rect 18028 820 18068 860
rect 4928 736 4968 776
rect 5010 736 5050 776
rect 5092 736 5132 776
rect 5174 736 5214 776
rect 5256 736 5296 776
rect 20048 736 20088 776
rect 20130 736 20170 776
rect 20212 736 20252 776
rect 20294 736 20334 776
rect 20376 736 20416 776
rect 35168 736 35208 776
rect 35250 736 35290 776
rect 35332 736 35372 776
rect 35414 736 35454 776
rect 35496 736 35536 776
<< metal4 >>
rect 20620 10688 20660 10697
rect 4588 10520 4628 10529
rect 1612 9848 1652 9857
rect 1612 7169 1652 9808
rect 3688 9092 4056 9101
rect 3728 9052 3770 9092
rect 3810 9052 3852 9092
rect 3892 9052 3934 9092
rect 3974 9052 4016 9092
rect 3688 9043 4056 9052
rect 3723 8672 3765 8681
rect 3723 8632 3724 8672
rect 3764 8632 3765 8672
rect 3723 8623 3765 8632
rect 3724 8538 3764 8623
rect 4108 8336 4148 8345
rect 1900 7832 1940 7841
rect 1900 7337 1940 7792
rect 3688 7580 4056 7589
rect 3728 7540 3770 7580
rect 3810 7540 3852 7580
rect 3892 7540 3934 7580
rect 3974 7540 4016 7580
rect 3688 7531 4056 7540
rect 2476 7496 2516 7505
rect 1899 7328 1941 7337
rect 1899 7288 1900 7328
rect 1940 7288 1941 7328
rect 1899 7279 1941 7288
rect 1611 7160 1653 7169
rect 1611 7120 1612 7160
rect 1652 7120 1653 7160
rect 1611 7111 1653 7120
rect 1612 6320 1652 7111
rect 1612 6271 1652 6280
rect 1900 6320 1940 7279
rect 1900 6271 1940 6280
rect 1708 6152 1748 6161
rect 1708 4985 1748 6112
rect 1707 4976 1749 4985
rect 1707 4936 1708 4976
rect 1748 4936 1749 4976
rect 1707 4927 1749 4936
rect 1708 4842 1748 4927
rect 1227 4808 1269 4817
rect 1227 4768 1228 4808
rect 1268 4768 1269 4808
rect 1227 4759 1269 4768
rect 1228 4674 1268 4759
rect 2476 1112 2516 7456
rect 4108 7160 4148 8296
rect 4588 8177 4628 10480
rect 16972 10520 17012 10529
rect 16395 10016 16437 10025
rect 16395 9976 16396 10016
rect 16436 9976 16437 10016
rect 16395 9967 16437 9976
rect 16396 9882 16436 9967
rect 4928 9848 5296 9857
rect 4968 9808 5010 9848
rect 5050 9808 5092 9848
rect 5132 9808 5174 9848
rect 5214 9808 5256 9848
rect 4928 9799 5296 9808
rect 12652 9680 12692 9689
rect 5452 9512 5492 9521
rect 5355 8504 5397 8513
rect 5355 8464 5356 8504
rect 5396 8464 5397 8504
rect 5355 8455 5397 8464
rect 4928 8336 5296 8345
rect 4968 8296 5010 8336
rect 5050 8296 5092 8336
rect 5132 8296 5174 8336
rect 5214 8296 5256 8336
rect 4928 8287 5296 8296
rect 4587 8168 4629 8177
rect 4587 8128 4588 8168
rect 4628 8128 4629 8168
rect 4587 8119 4629 8128
rect 4588 7244 4628 8119
rect 4588 7195 4628 7204
rect 4108 7111 4148 7120
rect 5356 7160 5396 8455
rect 5452 7832 5492 9472
rect 7564 9428 7604 9437
rect 5452 7783 5492 7792
rect 5548 8504 5588 8513
rect 5356 7111 5396 7120
rect 4928 6824 5296 6833
rect 4968 6784 5010 6824
rect 5050 6784 5092 6824
rect 5132 6784 5174 6824
rect 5214 6784 5256 6824
rect 4928 6775 5296 6784
rect 5548 6488 5588 8464
rect 6604 8252 6644 8261
rect 6412 8000 6452 8009
rect 6028 7916 6068 7925
rect 4684 6236 4724 6245
rect 4300 6152 4340 6161
rect 3688 6068 4056 6077
rect 3728 6028 3770 6068
rect 3810 6028 3852 6068
rect 3892 6028 3934 6068
rect 3974 6028 4016 6068
rect 3688 6019 4056 6028
rect 4204 5816 4244 5825
rect 4108 5648 4148 5657
rect 3688 4556 4056 4565
rect 3728 4516 3770 4556
rect 3810 4516 3852 4556
rect 3892 4516 3934 4556
rect 3974 4516 4016 4556
rect 3688 4507 4056 4516
rect 4108 3212 4148 5608
rect 4204 4808 4244 5776
rect 4204 4759 4244 4768
rect 4108 3163 4148 3172
rect 3688 3044 4056 3053
rect 3728 3004 3770 3044
rect 3810 3004 3852 3044
rect 3892 3004 3934 3044
rect 3974 3004 4016 3044
rect 3688 2995 4056 3004
rect 4300 2960 4340 6112
rect 4396 5984 4436 5993
rect 4396 4640 4436 5944
rect 4436 4600 4532 4640
rect 4396 4591 4436 4600
rect 4300 2911 4340 2920
rect 4492 1616 4532 4600
rect 4684 4304 4724 6196
rect 5260 5480 5300 5489
rect 5300 5440 5396 5480
rect 5260 5431 5300 5440
rect 4928 5312 5296 5321
rect 4968 5272 5010 5312
rect 5050 5272 5092 5312
rect 5132 5272 5174 5312
rect 5214 5272 5256 5312
rect 4928 5263 5296 5272
rect 5356 4976 5396 5440
rect 5356 4927 5396 4936
rect 4588 4136 4628 4145
rect 4588 3212 4628 4096
rect 4588 3163 4628 3172
rect 4684 2624 4724 4264
rect 4780 4472 4820 4481
rect 4780 3128 4820 4432
rect 4928 3800 5296 3809
rect 4968 3760 5010 3800
rect 5050 3760 5092 3800
rect 5132 3760 5174 3800
rect 5214 3760 5256 3800
rect 4928 3751 5296 3760
rect 5548 3632 5588 6448
rect 5740 7748 5780 7757
rect 5740 5648 5780 7708
rect 5740 5599 5780 5608
rect 6028 6404 6068 7876
rect 6028 5648 6068 6364
rect 6028 5599 6068 5608
rect 5548 3583 5588 3592
rect 4780 3079 4820 3088
rect 4684 2575 4724 2584
rect 4928 2288 5296 2297
rect 4968 2248 5010 2288
rect 5050 2248 5092 2288
rect 5132 2248 5174 2288
rect 5214 2248 5256 2288
rect 4928 2239 5296 2248
rect 4492 1567 4532 1576
rect 3688 1532 4056 1541
rect 3728 1492 3770 1532
rect 3810 1492 3852 1532
rect 3892 1492 3934 1532
rect 3974 1492 4016 1532
rect 3688 1483 4056 1492
rect 2476 617 2516 1072
rect 6412 944 6452 7960
rect 6604 6152 6644 8212
rect 7564 7085 7604 9388
rect 10348 9428 10388 9437
rect 10252 8840 10292 8849
rect 8811 8672 8853 8681
rect 8811 8632 8812 8672
rect 8852 8632 8853 8672
rect 8811 8623 8853 8632
rect 9771 8672 9813 8681
rect 9771 8632 9772 8672
rect 9812 8632 9813 8672
rect 9771 8623 9813 8632
rect 8812 8538 8852 8623
rect 9772 8538 9812 8623
rect 8043 7160 8085 7169
rect 8043 7120 8044 7160
rect 8084 7120 8085 7160
rect 8043 7111 8085 7120
rect 7563 7076 7605 7085
rect 7563 7036 7564 7076
rect 7604 7036 7605 7076
rect 7563 7027 7605 7036
rect 6604 6103 6644 6112
rect 7180 6740 7220 6749
rect 7180 5984 7220 6700
rect 7180 5935 7220 5944
rect 7564 4817 7604 7027
rect 8044 7026 8084 7111
rect 7563 4808 7605 4817
rect 7563 4768 7564 4808
rect 7604 4768 7605 4808
rect 7563 4759 7605 4768
rect 10252 2465 10292 8800
rect 10348 4901 10388 9388
rect 11020 8840 11060 8849
rect 10731 6404 10773 6413
rect 10731 6364 10732 6404
rect 10772 6364 10773 6404
rect 10731 6355 10773 6364
rect 10732 6270 10772 6355
rect 10347 4892 10389 4901
rect 10347 4852 10348 4892
rect 10388 4852 10389 4892
rect 10347 4843 10389 4852
rect 11020 3305 11060 8800
rect 11788 8840 11828 8849
rect 11404 8756 11444 8765
rect 11404 8084 11444 8716
rect 11404 8035 11444 8044
rect 11500 7412 11540 7421
rect 11500 6908 11540 7372
rect 11500 6859 11540 6868
rect 11019 3296 11061 3305
rect 11019 3256 11020 3296
rect 11060 3256 11061 3296
rect 11019 3247 11061 3256
rect 10251 2456 10293 2465
rect 10251 2416 10252 2456
rect 10292 2416 10293 2456
rect 10251 2407 10293 2416
rect 11788 2045 11828 8800
rect 12556 8840 12596 8849
rect 12363 8168 12405 8177
rect 12363 8128 12364 8168
rect 12404 8128 12405 8168
rect 12363 8119 12405 8128
rect 12364 8000 12404 8119
rect 12364 7951 12404 7960
rect 12076 7580 12116 7589
rect 11787 2036 11829 2045
rect 11787 1996 11788 2036
rect 11828 1996 11829 2036
rect 11787 1987 11829 1996
rect 12076 1877 12116 7540
rect 12556 5312 12596 8800
rect 12652 5489 12692 9640
rect 15244 9680 15284 9689
rect 14188 9176 14228 9185
rect 14092 8840 14132 8849
rect 13035 8672 13077 8681
rect 13035 8632 13036 8672
rect 13076 8632 13077 8672
rect 13035 8623 13077 8632
rect 13036 6245 13076 8623
rect 13996 8504 14036 8513
rect 13803 7244 13845 7253
rect 13803 7204 13804 7244
rect 13844 7204 13845 7244
rect 13803 7195 13845 7204
rect 13804 6992 13844 7195
rect 13804 6943 13844 6952
rect 13899 6404 13941 6413
rect 13899 6364 13900 6404
rect 13940 6364 13941 6404
rect 13899 6355 13941 6364
rect 13035 6236 13077 6245
rect 13035 6196 13036 6236
rect 13076 6196 13077 6236
rect 13035 6187 13077 6196
rect 12651 5480 12693 5489
rect 12651 5440 12652 5480
rect 12692 5440 12693 5480
rect 12651 5431 12693 5440
rect 12556 5272 12692 5312
rect 12652 4733 12692 5272
rect 12651 4724 12693 4733
rect 12651 4684 12652 4724
rect 12692 4684 12693 4724
rect 12651 4675 12693 4684
rect 12267 3464 12309 3473
rect 12267 3424 12268 3464
rect 12308 3424 12309 3464
rect 12267 3415 12309 3424
rect 13900 3464 13940 6355
rect 13996 6329 14036 8464
rect 13995 6320 14037 6329
rect 13995 6280 13996 6320
rect 14036 6280 14037 6320
rect 13995 6271 14037 6280
rect 13900 3415 13940 3424
rect 12268 3330 12308 3415
rect 14092 2129 14132 8800
rect 14188 5909 14228 9136
rect 14476 8840 14516 8849
rect 14187 5900 14229 5909
rect 14187 5860 14188 5900
rect 14228 5860 14229 5900
rect 14187 5851 14229 5860
rect 14091 2120 14133 2129
rect 14091 2080 14092 2120
rect 14132 2080 14133 2120
rect 14091 2071 14133 2080
rect 12075 1868 12117 1877
rect 12075 1828 12076 1868
rect 12116 1828 12117 1868
rect 12075 1819 12117 1828
rect 9772 1784 9812 1793
rect 9772 1037 9812 1744
rect 14476 1121 14516 8800
rect 14860 8672 14900 8683
rect 14860 8597 14900 8632
rect 14859 8588 14901 8597
rect 14859 8548 14860 8588
rect 14900 8548 14901 8588
rect 14859 8539 14901 8548
rect 14860 6068 14900 8539
rect 14860 6019 14900 6028
rect 15244 3641 15284 9640
rect 16396 9596 16436 9605
rect 15436 8840 15476 8849
rect 15243 3632 15285 3641
rect 15243 3592 15244 3632
rect 15284 3592 15285 3632
rect 15243 3583 15285 3592
rect 15436 3221 15476 8800
rect 15628 8840 15668 8849
rect 15628 5825 15668 8800
rect 16012 8840 16052 8849
rect 15820 8672 15860 8681
rect 15820 8513 15860 8632
rect 15819 8504 15861 8513
rect 15819 8464 15820 8504
rect 15860 8464 15861 8504
rect 15819 8455 15861 8464
rect 15820 8177 15860 8455
rect 15819 8168 15861 8177
rect 15819 8128 15820 8168
rect 15860 8128 15861 8168
rect 15819 8119 15861 8128
rect 15627 5816 15669 5825
rect 15627 5776 15628 5816
rect 15668 5776 15669 5816
rect 15627 5767 15669 5776
rect 15532 4976 15572 4985
rect 15532 3464 15572 4936
rect 16012 3557 16052 8800
rect 16396 8513 16436 9556
rect 16780 8840 16820 8849
rect 16395 8504 16437 8513
rect 16395 8464 16396 8504
rect 16436 8464 16437 8504
rect 16395 8455 16437 8464
rect 16107 5648 16149 5657
rect 16107 5608 16108 5648
rect 16148 5608 16149 5648
rect 16107 5599 16149 5608
rect 16108 5514 16148 5599
rect 16780 4061 16820 8800
rect 16972 7757 17012 10480
rect 18700 10520 18740 10529
rect 18124 8840 18164 8849
rect 16971 7748 17013 7757
rect 16971 7708 16972 7748
rect 17012 7708 17013 7748
rect 16971 7699 17013 7708
rect 17643 7412 17685 7421
rect 17643 7372 17644 7412
rect 17684 7372 17685 7412
rect 17643 7363 17685 7372
rect 17644 7160 17684 7363
rect 17644 7085 17684 7120
rect 17643 7076 17685 7085
rect 17643 7036 17644 7076
rect 17684 7036 17685 7076
rect 17643 7027 17685 7036
rect 18124 4817 18164 8800
rect 18123 4808 18165 4817
rect 18123 4768 18124 4808
rect 18164 4768 18165 4808
rect 18123 4759 18165 4768
rect 16779 4052 16821 4061
rect 16779 4012 16780 4052
rect 16820 4012 16821 4052
rect 16779 4003 16821 4012
rect 18700 3977 18740 10480
rect 20048 9848 20416 9857
rect 20088 9808 20130 9848
rect 20170 9808 20212 9848
rect 20252 9808 20294 9848
rect 20334 9808 20376 9848
rect 20048 9799 20416 9808
rect 18808 9092 19176 9101
rect 18848 9052 18890 9092
rect 18930 9052 18972 9092
rect 19012 9052 19054 9092
rect 19094 9052 19136 9092
rect 18808 9043 19176 9052
rect 19468 8672 19508 8681
rect 18892 8504 18932 8513
rect 18892 7841 18932 8464
rect 19468 8336 19508 8632
rect 19468 8287 19508 8296
rect 20048 8336 20416 8345
rect 20088 8296 20130 8336
rect 20170 8296 20212 8336
rect 20252 8296 20294 8336
rect 20334 8296 20376 8336
rect 20048 8287 20416 8296
rect 20620 8336 20660 10648
rect 18891 7832 18933 7841
rect 18891 7792 18892 7832
rect 18932 7792 18933 7832
rect 18891 7783 18933 7792
rect 18808 7580 19176 7589
rect 18848 7540 18890 7580
rect 18930 7540 18972 7580
rect 19012 7540 19054 7580
rect 19094 7540 19136 7580
rect 18808 7531 19176 7540
rect 19372 7160 19412 7169
rect 18808 6068 19176 6077
rect 18848 6028 18890 6068
rect 18930 6028 18972 6068
rect 19012 6028 19054 6068
rect 19094 6028 19136 6068
rect 18808 6019 19176 6028
rect 19372 4985 19412 7120
rect 20048 6824 20416 6833
rect 20088 6784 20130 6824
rect 20170 6784 20212 6824
rect 20252 6784 20294 6824
rect 20334 6784 20376 6824
rect 20048 6775 20416 6784
rect 20043 6320 20085 6329
rect 20043 6280 20044 6320
rect 20084 6280 20085 6320
rect 20043 6271 20085 6280
rect 20044 6161 20084 6271
rect 20235 6236 20277 6245
rect 20235 6196 20236 6236
rect 20276 6196 20277 6236
rect 20235 6187 20277 6196
rect 20043 6152 20085 6161
rect 20043 6112 20044 6152
rect 20084 6112 20085 6152
rect 20043 6103 20085 6112
rect 20236 5993 20276 6187
rect 20235 5984 20277 5993
rect 20235 5944 20236 5984
rect 20276 5944 20277 5984
rect 20235 5935 20277 5944
rect 20620 5732 20660 8296
rect 21100 10268 21140 10277
rect 20620 5683 20660 5692
rect 20716 7748 20756 7757
rect 20716 5657 20756 7708
rect 21100 5816 21140 10228
rect 22731 10016 22773 10025
rect 22731 9976 22732 10016
rect 22772 9976 22773 10016
rect 22731 9967 22773 9976
rect 22636 9596 22676 9605
rect 22252 8840 22292 8849
rect 22252 8597 22292 8800
rect 22251 8588 22293 8597
rect 22251 8548 22252 8588
rect 22292 8548 22293 8588
rect 22251 8539 22293 8548
rect 22252 8000 22292 8539
rect 22252 7951 22292 7960
rect 22636 7841 22676 9556
rect 22732 9092 22772 9967
rect 35168 9848 35536 9857
rect 35208 9808 35250 9848
rect 35290 9808 35332 9848
rect 35372 9808 35414 9848
rect 35454 9808 35496 9848
rect 35168 9799 35536 9808
rect 22732 9043 22772 9052
rect 22828 9512 22868 9521
rect 22635 7832 22677 7841
rect 22635 7792 22636 7832
rect 22676 7792 22677 7832
rect 22635 7783 22677 7792
rect 21676 6656 21716 6665
rect 21676 6488 21716 6616
rect 21676 5900 21716 6448
rect 21676 5851 21716 5860
rect 21100 5767 21140 5776
rect 20715 5648 20757 5657
rect 20715 5608 20716 5648
rect 20756 5608 20757 5648
rect 20715 5599 20757 5608
rect 20048 5312 20416 5321
rect 20088 5272 20130 5312
rect 20170 5272 20212 5312
rect 20252 5272 20294 5312
rect 20334 5272 20376 5312
rect 20048 5263 20416 5272
rect 19371 4976 19413 4985
rect 19371 4936 19372 4976
rect 19412 4936 19413 4976
rect 19371 4927 19413 4936
rect 18808 4556 19176 4565
rect 18848 4516 18890 4556
rect 18930 4516 18972 4556
rect 19012 4516 19054 4556
rect 19094 4516 19136 4556
rect 18808 4507 19176 4516
rect 18699 3968 18741 3977
rect 18699 3928 18700 3968
rect 18740 3928 18741 3968
rect 18699 3919 18741 3928
rect 16011 3548 16053 3557
rect 16011 3508 16012 3548
rect 16052 3508 16053 3548
rect 16011 3499 16053 3508
rect 15435 3212 15477 3221
rect 15435 3172 15436 3212
rect 15476 3172 15477 3212
rect 15435 3163 15477 3172
rect 14475 1112 14517 1121
rect 14475 1072 14476 1112
rect 14516 1072 14517 1112
rect 14475 1063 14517 1072
rect 9771 1028 9813 1037
rect 9771 988 9772 1028
rect 9812 988 9813 1028
rect 9771 979 9813 988
rect 6412 895 6452 904
rect 9772 944 9812 979
rect 15532 953 15572 3424
rect 19372 3389 19412 4927
rect 22636 4304 22676 7783
rect 22828 7253 22868 9472
rect 40876 9428 40916 9437
rect 37612 9260 37652 9269
rect 26284 9092 26324 9101
rect 23308 8252 23348 8261
rect 23308 8177 23348 8212
rect 23307 8168 23349 8177
rect 23307 8128 23308 8168
rect 23348 8128 23349 8168
rect 23307 8119 23349 8128
rect 22827 7244 22869 7253
rect 22827 7204 22828 7244
rect 22868 7204 22869 7244
rect 22827 7195 22869 7204
rect 23308 5732 23348 8119
rect 23884 7916 23924 7925
rect 23884 7421 23924 7876
rect 24075 7916 24117 7925
rect 24075 7876 24076 7916
rect 24116 7876 24117 7916
rect 24075 7867 24117 7876
rect 24076 7782 24116 7867
rect 23883 7412 23925 7421
rect 23883 7372 23884 7412
rect 23924 7372 23925 7412
rect 23883 7363 23925 7372
rect 26284 7328 26324 9052
rect 33928 9092 34296 9101
rect 33968 9052 34010 9092
rect 34050 9052 34092 9092
rect 34132 9052 34174 9092
rect 34214 9052 34256 9092
rect 33928 9043 34296 9052
rect 33772 8840 33812 8849
rect 33196 8756 33236 8765
rect 30796 8588 30836 8597
rect 27724 8504 27764 8513
rect 26284 7279 26324 7288
rect 26860 8252 26900 8261
rect 26860 7328 26900 8212
rect 26860 7279 26900 7288
rect 23308 5683 23348 5692
rect 22636 4255 22676 4264
rect 25804 5648 25844 5657
rect 20048 3800 20416 3809
rect 20088 3760 20130 3800
rect 20170 3760 20212 3800
rect 20252 3760 20294 3800
rect 20334 3760 20376 3800
rect 20048 3751 20416 3760
rect 19948 3473 19988 3504
rect 19947 3464 19989 3473
rect 19947 3424 19948 3464
rect 19988 3424 19989 3464
rect 19947 3415 19989 3424
rect 19371 3380 19413 3389
rect 19371 3340 19372 3380
rect 19412 3340 19413 3380
rect 19371 3331 19413 3340
rect 19948 3380 19988 3415
rect 18808 3044 19176 3053
rect 18848 3004 18890 3044
rect 18930 3004 18972 3044
rect 19012 3004 19054 3044
rect 19094 3004 19136 3044
rect 18808 2995 19176 3004
rect 18028 2540 18068 2549
rect 18028 1961 18068 2500
rect 18027 1952 18069 1961
rect 18027 1912 18028 1952
rect 18068 1912 18069 1952
rect 18027 1903 18069 1912
rect 9772 893 9812 904
rect 15531 944 15573 953
rect 15531 904 15532 944
rect 15572 904 15573 944
rect 15531 895 15573 904
rect 18028 860 18068 1903
rect 18808 1532 19176 1541
rect 18848 1492 18890 1532
rect 18930 1492 18972 1532
rect 19012 1492 19054 1532
rect 19094 1492 19136 1532
rect 18808 1483 19176 1492
rect 19948 1205 19988 3340
rect 21388 2792 21428 2801
rect 21388 2540 21428 2752
rect 21388 2491 21428 2500
rect 20048 2288 20416 2297
rect 20088 2248 20130 2288
rect 20170 2248 20212 2288
rect 20252 2248 20294 2288
rect 20334 2248 20376 2288
rect 20048 2239 20416 2248
rect 19947 1196 19989 1205
rect 19947 1156 19948 1196
rect 19988 1156 19989 1196
rect 19947 1147 19989 1156
rect 25420 1196 25460 1205
rect 25420 1037 25460 1156
rect 25419 1028 25461 1037
rect 25419 988 25420 1028
rect 25460 988 25461 1028
rect 25419 979 25461 988
rect 18028 811 18068 820
rect 4928 776 5296 785
rect 4968 736 5010 776
rect 5050 736 5092 776
rect 5132 736 5174 776
rect 5214 736 5256 776
rect 4928 727 5296 736
rect 20048 776 20416 785
rect 20088 736 20130 776
rect 20170 736 20212 776
rect 20252 736 20294 776
rect 20334 736 20376 776
rect 20048 727 20416 736
rect 25804 617 25844 5608
rect 27724 1877 27764 8464
rect 27916 8504 27956 8513
rect 27819 7328 27861 7337
rect 27819 7288 27820 7328
rect 27860 7288 27861 7328
rect 27819 7279 27861 7288
rect 27820 7160 27860 7279
rect 27820 5984 27860 7120
rect 27820 5935 27860 5944
rect 27916 5909 27956 8464
rect 28012 8000 28052 8011
rect 28012 7925 28052 7960
rect 28876 8000 28916 8009
rect 28011 7916 28053 7925
rect 28011 7876 28012 7916
rect 28052 7876 28053 7916
rect 28011 7867 28053 7876
rect 28588 7832 28628 7841
rect 28876 7832 28916 7960
rect 28628 7792 28916 7832
rect 28588 7783 28628 7792
rect 28972 7076 29012 7085
rect 28972 6404 29012 7036
rect 28972 6355 29012 6364
rect 29548 6992 29588 7001
rect 28972 5984 29012 5993
rect 29012 5944 29108 5984
rect 28972 5935 29012 5944
rect 27915 5900 27957 5909
rect 27915 5860 27916 5900
rect 27956 5860 27957 5900
rect 27915 5851 27957 5860
rect 29068 5816 29108 5944
rect 29068 5767 29108 5776
rect 28299 5480 28341 5489
rect 28299 5440 28300 5480
rect 28340 5440 28341 5480
rect 28299 5431 28341 5440
rect 28300 5346 28340 5431
rect 29548 3305 29588 6952
rect 30220 6740 30260 6749
rect 29547 3296 29589 3305
rect 29547 3256 29548 3296
rect 29588 3256 29589 3296
rect 29547 3247 29589 3256
rect 28779 3212 28821 3221
rect 28779 3172 28780 3212
rect 28820 3172 28821 3212
rect 28779 3163 28821 3172
rect 28780 3078 28820 3163
rect 30220 2045 30260 6700
rect 30796 2120 30836 8548
rect 30988 8504 31028 8513
rect 30988 5825 31028 8464
rect 31371 8504 31413 8513
rect 31371 8464 31372 8504
rect 31412 8464 31413 8504
rect 31371 8455 31413 8464
rect 31756 8504 31796 8513
rect 31372 8370 31412 8455
rect 31372 7748 31412 7757
rect 30987 5816 31029 5825
rect 30987 5776 30988 5816
rect 31028 5776 31029 5816
rect 30987 5767 31029 5776
rect 31372 3557 31412 7708
rect 31756 3641 31796 8464
rect 33004 8420 33044 8429
rect 32619 7748 32661 7757
rect 32619 7708 32620 7748
rect 32660 7708 32661 7748
rect 32619 7699 32661 7708
rect 32620 7614 32660 7699
rect 31947 7328 31989 7337
rect 31947 7288 31948 7328
rect 31988 7288 31989 7328
rect 31947 7279 31989 7288
rect 31948 7194 31988 7279
rect 31755 3632 31797 3641
rect 31755 3592 31756 3632
rect 31796 3592 31797 3632
rect 31755 3583 31797 3592
rect 31371 3548 31413 3557
rect 31371 3508 31372 3548
rect 31412 3508 31413 3548
rect 31371 3499 31413 3508
rect 30796 2071 30836 2080
rect 30219 2036 30261 2045
rect 30219 1996 30220 2036
rect 30260 1996 30261 2036
rect 30219 1987 30261 1996
rect 29547 1952 29589 1961
rect 29547 1912 29548 1952
rect 29588 1912 29589 1952
rect 29547 1903 29589 1912
rect 27723 1868 27765 1877
rect 27723 1828 27724 1868
rect 27764 1828 27765 1868
rect 27723 1819 27765 1828
rect 29548 1818 29588 1903
rect 33004 1448 33044 8380
rect 33100 8168 33140 8177
rect 33100 5312 33140 8128
rect 33100 5263 33140 5272
rect 33196 1700 33236 8716
rect 33388 6488 33428 6497
rect 33388 3389 33428 6448
rect 33772 4901 33812 8800
rect 35168 8336 35536 8345
rect 35208 8296 35250 8336
rect 35290 8296 35332 8336
rect 35372 8296 35414 8336
rect 35454 8296 35496 8336
rect 35168 8287 35536 8296
rect 34636 7664 34676 7673
rect 33928 7580 34296 7589
rect 33968 7540 34010 7580
rect 34050 7540 34092 7580
rect 34132 7540 34174 7580
rect 34214 7540 34256 7580
rect 33928 7531 34296 7540
rect 33928 6068 34296 6077
rect 33968 6028 34010 6068
rect 34050 6028 34092 6068
rect 34132 6028 34174 6068
rect 34214 6028 34256 6068
rect 33928 6019 34296 6028
rect 33771 4892 33813 4901
rect 33771 4852 33772 4892
rect 33812 4852 33813 4892
rect 33771 4843 33813 4852
rect 33928 4556 34296 4565
rect 33968 4516 34010 4556
rect 34050 4516 34092 4556
rect 34132 4516 34174 4556
rect 34214 4516 34256 4556
rect 33928 4507 34296 4516
rect 33963 4052 34005 4061
rect 33963 4012 33964 4052
rect 34004 4012 34100 4052
rect 33963 4003 34005 4012
rect 34060 3968 34100 4012
rect 34060 3919 34100 3928
rect 33387 3380 33429 3389
rect 33387 3340 33388 3380
rect 33428 3340 33429 3380
rect 33387 3331 33429 3340
rect 33928 3044 34296 3053
rect 33968 3004 34010 3044
rect 34050 3004 34092 3044
rect 34132 3004 34174 3044
rect 34214 3004 34256 3044
rect 33928 2995 34296 3004
rect 34636 2036 34676 7624
rect 34636 1987 34676 1996
rect 35020 7412 35060 7421
rect 33196 1651 33236 1660
rect 33928 1532 34296 1541
rect 33968 1492 34010 1532
rect 34050 1492 34092 1532
rect 34132 1492 34174 1532
rect 34214 1492 34256 1532
rect 33928 1483 34296 1492
rect 33004 1399 33044 1408
rect 35020 944 35060 7372
rect 35168 6824 35536 6833
rect 35208 6784 35250 6824
rect 35290 6784 35332 6824
rect 35372 6784 35414 6824
rect 35454 6784 35496 6824
rect 35168 6775 35536 6784
rect 35692 6320 35732 6329
rect 35168 5312 35536 5321
rect 35208 5272 35250 5312
rect 35290 5272 35332 5312
rect 35372 5272 35414 5312
rect 35454 5272 35496 5312
rect 35168 5263 35536 5272
rect 35168 3800 35536 3809
rect 35208 3760 35250 3800
rect 35290 3760 35332 3800
rect 35372 3760 35414 3800
rect 35454 3760 35496 3800
rect 35168 3751 35536 3760
rect 35692 2465 35732 6280
rect 36651 4808 36693 4817
rect 36651 4768 36652 4808
rect 36692 4768 36693 4808
rect 36651 4759 36693 4768
rect 36652 4674 36692 4759
rect 36843 3968 36885 3977
rect 36843 3928 36844 3968
rect 36884 3928 36885 3968
rect 36843 3919 36885 3928
rect 36844 3834 36884 3919
rect 35691 2456 35733 2465
rect 35691 2416 35692 2456
rect 35732 2416 35733 2456
rect 35691 2407 35733 2416
rect 35168 2288 35536 2297
rect 35208 2248 35250 2288
rect 35290 2248 35332 2288
rect 35372 2248 35414 2288
rect 35454 2248 35496 2288
rect 35168 2239 35536 2248
rect 37612 2129 37652 9220
rect 39724 8504 39764 8513
rect 37611 2120 37653 2129
rect 37611 2080 37612 2120
rect 37652 2080 37653 2120
rect 37611 2071 37653 2080
rect 35596 1280 35636 1289
rect 35596 1037 35636 1240
rect 39724 1121 39764 8464
rect 40300 7244 40340 7253
rect 40204 6320 40244 6360
rect 40204 6245 40244 6280
rect 40203 6236 40245 6245
rect 40203 6196 40204 6236
rect 40244 6196 40245 6236
rect 40203 6187 40245 6196
rect 39723 1112 39765 1121
rect 39723 1072 39724 1112
rect 39764 1072 39765 1112
rect 39723 1063 39765 1072
rect 35595 1028 35637 1037
rect 35595 988 35596 1028
rect 35636 988 35637 1028
rect 35595 979 35637 988
rect 40300 953 40340 7204
rect 40876 5909 40916 9388
rect 41260 6413 41300 6498
rect 41259 6404 41301 6413
rect 41259 6364 41260 6404
rect 41300 6364 41301 6404
rect 41259 6355 41301 6364
rect 40875 5900 40917 5909
rect 40875 5860 40876 5900
rect 40916 5860 40917 5900
rect 40875 5851 40917 5860
rect 40491 4724 40533 4733
rect 40491 4684 40492 4724
rect 40532 4684 40533 4724
rect 40491 4675 40533 4684
rect 40492 4590 40532 4675
rect 40875 1196 40917 1205
rect 40875 1156 40876 1196
rect 40916 1156 40917 1196
rect 40875 1147 40917 1156
rect 40876 1062 40916 1147
rect 35020 895 35060 904
rect 40299 944 40341 953
rect 40299 904 40300 944
rect 40340 904 40341 944
rect 40299 895 40341 904
rect 35168 776 35536 785
rect 35208 736 35250 776
rect 35290 736 35332 776
rect 35372 736 35414 776
rect 35454 736 35496 776
rect 35168 727 35536 736
rect 2475 608 2517 617
rect 2475 568 2476 608
rect 2516 568 2517 608
rect 2475 559 2517 568
rect 25803 608 25845 617
rect 25803 568 25804 608
rect 25844 568 25845 608
rect 25803 559 25845 568
<< via4 >>
rect 3688 9052 3728 9092
rect 3770 9052 3810 9092
rect 3852 9052 3892 9092
rect 3934 9052 3974 9092
rect 4016 9052 4056 9092
rect 3724 8632 3764 8672
rect 3688 7540 3728 7580
rect 3770 7540 3810 7580
rect 3852 7540 3892 7580
rect 3934 7540 3974 7580
rect 4016 7540 4056 7580
rect 1900 7288 1940 7328
rect 1612 7120 1652 7160
rect 1708 4936 1748 4976
rect 1228 4768 1268 4808
rect 16396 9976 16436 10016
rect 4928 9808 4968 9848
rect 5010 9808 5050 9848
rect 5092 9808 5132 9848
rect 5174 9808 5214 9848
rect 5256 9808 5296 9848
rect 5356 8464 5396 8504
rect 4928 8296 4968 8336
rect 5010 8296 5050 8336
rect 5092 8296 5132 8336
rect 5174 8296 5214 8336
rect 5256 8296 5296 8336
rect 4588 8128 4628 8168
rect 4928 6784 4968 6824
rect 5010 6784 5050 6824
rect 5092 6784 5132 6824
rect 5174 6784 5214 6824
rect 5256 6784 5296 6824
rect 3688 6028 3728 6068
rect 3770 6028 3810 6068
rect 3852 6028 3892 6068
rect 3934 6028 3974 6068
rect 4016 6028 4056 6068
rect 3688 4516 3728 4556
rect 3770 4516 3810 4556
rect 3852 4516 3892 4556
rect 3934 4516 3974 4556
rect 4016 4516 4056 4556
rect 3688 3004 3728 3044
rect 3770 3004 3810 3044
rect 3852 3004 3892 3044
rect 3934 3004 3974 3044
rect 4016 3004 4056 3044
rect 4928 5272 4968 5312
rect 5010 5272 5050 5312
rect 5092 5272 5132 5312
rect 5174 5272 5214 5312
rect 5256 5272 5296 5312
rect 4928 3760 4968 3800
rect 5010 3760 5050 3800
rect 5092 3760 5132 3800
rect 5174 3760 5214 3800
rect 5256 3760 5296 3800
rect 4928 2248 4968 2288
rect 5010 2248 5050 2288
rect 5092 2248 5132 2288
rect 5174 2248 5214 2288
rect 5256 2248 5296 2288
rect 3688 1492 3728 1532
rect 3770 1492 3810 1532
rect 3852 1492 3892 1532
rect 3934 1492 3974 1532
rect 4016 1492 4056 1532
rect 8812 8632 8852 8672
rect 9772 8632 9812 8672
rect 8044 7120 8084 7160
rect 7564 7036 7604 7076
rect 7564 4768 7604 4808
rect 10732 6364 10772 6404
rect 10348 4852 10388 4892
rect 11020 3256 11060 3296
rect 10252 2416 10292 2456
rect 12364 8128 12404 8168
rect 11788 1996 11828 2036
rect 13036 8632 13076 8672
rect 13804 7204 13844 7244
rect 13900 6364 13940 6404
rect 13036 6196 13076 6236
rect 12652 5440 12692 5480
rect 12652 4684 12692 4724
rect 12268 3424 12308 3464
rect 13996 6280 14036 6320
rect 14188 5860 14228 5900
rect 14092 2080 14132 2120
rect 12076 1828 12116 1868
rect 14860 8548 14900 8588
rect 15244 3592 15284 3632
rect 15820 8464 15860 8504
rect 15820 8128 15860 8168
rect 15628 5776 15668 5816
rect 16396 8464 16436 8504
rect 16108 5608 16148 5648
rect 16972 7708 17012 7748
rect 17644 7372 17684 7412
rect 17644 7036 17684 7076
rect 18124 4768 18164 4808
rect 16780 4012 16820 4052
rect 20048 9808 20088 9848
rect 20130 9808 20170 9848
rect 20212 9808 20252 9848
rect 20294 9808 20334 9848
rect 20376 9808 20416 9848
rect 18808 9052 18848 9092
rect 18890 9052 18930 9092
rect 18972 9052 19012 9092
rect 19054 9052 19094 9092
rect 19136 9052 19176 9092
rect 20048 8296 20088 8336
rect 20130 8296 20170 8336
rect 20212 8296 20252 8336
rect 20294 8296 20334 8336
rect 20376 8296 20416 8336
rect 18892 7792 18932 7832
rect 18808 7540 18848 7580
rect 18890 7540 18930 7580
rect 18972 7540 19012 7580
rect 19054 7540 19094 7580
rect 19136 7540 19176 7580
rect 18808 6028 18848 6068
rect 18890 6028 18930 6068
rect 18972 6028 19012 6068
rect 19054 6028 19094 6068
rect 19136 6028 19176 6068
rect 20048 6784 20088 6824
rect 20130 6784 20170 6824
rect 20212 6784 20252 6824
rect 20294 6784 20334 6824
rect 20376 6784 20416 6824
rect 20044 6280 20084 6320
rect 20236 6196 20276 6236
rect 20044 6112 20084 6152
rect 20236 5944 20276 5984
rect 22732 9976 22772 10016
rect 22252 8548 22292 8588
rect 35168 9808 35208 9848
rect 35250 9808 35290 9848
rect 35332 9808 35372 9848
rect 35414 9808 35454 9848
rect 35496 9808 35536 9848
rect 22636 7792 22676 7832
rect 20716 5608 20756 5648
rect 20048 5272 20088 5312
rect 20130 5272 20170 5312
rect 20212 5272 20252 5312
rect 20294 5272 20334 5312
rect 20376 5272 20416 5312
rect 19372 4936 19412 4976
rect 18808 4516 18848 4556
rect 18890 4516 18930 4556
rect 18972 4516 19012 4556
rect 19054 4516 19094 4556
rect 19136 4516 19176 4556
rect 18700 3928 18740 3968
rect 16012 3508 16052 3548
rect 15436 3172 15476 3212
rect 14476 1072 14516 1112
rect 9772 988 9812 1028
rect 23308 8128 23348 8168
rect 22828 7204 22868 7244
rect 24076 7876 24116 7916
rect 23884 7372 23924 7412
rect 33928 9052 33968 9092
rect 34010 9052 34050 9092
rect 34092 9052 34132 9092
rect 34174 9052 34214 9092
rect 34256 9052 34296 9092
rect 20048 3760 20088 3800
rect 20130 3760 20170 3800
rect 20212 3760 20252 3800
rect 20294 3760 20334 3800
rect 20376 3760 20416 3800
rect 19948 3424 19988 3464
rect 19372 3340 19412 3380
rect 18808 3004 18848 3044
rect 18890 3004 18930 3044
rect 18972 3004 19012 3044
rect 19054 3004 19094 3044
rect 19136 3004 19176 3044
rect 18028 1912 18068 1952
rect 15532 904 15572 944
rect 18808 1492 18848 1532
rect 18890 1492 18930 1532
rect 18972 1492 19012 1532
rect 19054 1492 19094 1532
rect 19136 1492 19176 1532
rect 20048 2248 20088 2288
rect 20130 2248 20170 2288
rect 20212 2248 20252 2288
rect 20294 2248 20334 2288
rect 20376 2248 20416 2288
rect 19948 1156 19988 1196
rect 25420 988 25460 1028
rect 4928 736 4968 776
rect 5010 736 5050 776
rect 5092 736 5132 776
rect 5174 736 5214 776
rect 5256 736 5296 776
rect 20048 736 20088 776
rect 20130 736 20170 776
rect 20212 736 20252 776
rect 20294 736 20334 776
rect 20376 736 20416 776
rect 27820 7288 27860 7328
rect 28012 7876 28052 7916
rect 27916 5860 27956 5900
rect 28300 5440 28340 5480
rect 29548 3256 29588 3296
rect 28780 3172 28820 3212
rect 31372 8464 31412 8504
rect 30988 5776 31028 5816
rect 32620 7708 32660 7748
rect 31948 7288 31988 7328
rect 31756 3592 31796 3632
rect 31372 3508 31412 3548
rect 30220 1996 30260 2036
rect 29548 1912 29588 1952
rect 27724 1828 27764 1868
rect 35168 8296 35208 8336
rect 35250 8296 35290 8336
rect 35332 8296 35372 8336
rect 35414 8296 35454 8336
rect 35496 8296 35536 8336
rect 33928 7540 33968 7580
rect 34010 7540 34050 7580
rect 34092 7540 34132 7580
rect 34174 7540 34214 7580
rect 34256 7540 34296 7580
rect 33928 6028 33968 6068
rect 34010 6028 34050 6068
rect 34092 6028 34132 6068
rect 34174 6028 34214 6068
rect 34256 6028 34296 6068
rect 33772 4852 33812 4892
rect 33928 4516 33968 4556
rect 34010 4516 34050 4556
rect 34092 4516 34132 4556
rect 34174 4516 34214 4556
rect 34256 4516 34296 4556
rect 33964 4012 34004 4052
rect 33388 3340 33428 3380
rect 33928 3004 33968 3044
rect 34010 3004 34050 3044
rect 34092 3004 34132 3044
rect 34174 3004 34214 3044
rect 34256 3004 34296 3044
rect 33928 1492 33968 1532
rect 34010 1492 34050 1532
rect 34092 1492 34132 1532
rect 34174 1492 34214 1532
rect 34256 1492 34296 1532
rect 35168 6784 35208 6824
rect 35250 6784 35290 6824
rect 35332 6784 35372 6824
rect 35414 6784 35454 6824
rect 35496 6784 35536 6824
rect 35168 5272 35208 5312
rect 35250 5272 35290 5312
rect 35332 5272 35372 5312
rect 35414 5272 35454 5312
rect 35496 5272 35536 5312
rect 35168 3760 35208 3800
rect 35250 3760 35290 3800
rect 35332 3760 35372 3800
rect 35414 3760 35454 3800
rect 35496 3760 35536 3800
rect 36652 4768 36692 4808
rect 36844 3928 36884 3968
rect 35692 2416 35732 2456
rect 35168 2248 35208 2288
rect 35250 2248 35290 2288
rect 35332 2248 35372 2288
rect 35414 2248 35454 2288
rect 35496 2248 35536 2288
rect 37612 2080 37652 2120
rect 40204 6196 40244 6236
rect 39724 1072 39764 1112
rect 35596 988 35636 1028
rect 41260 6364 41300 6404
rect 40876 5860 40916 5900
rect 40492 4684 40532 4724
rect 40876 1156 40916 1196
rect 40300 904 40340 944
rect 35168 736 35208 776
rect 35250 736 35290 776
rect 35332 736 35372 776
rect 35414 736 35454 776
rect 35496 736 35536 776
rect 2476 568 2516 608
rect 25804 568 25844 608
<< metal5 >>
rect 16387 9976 16396 10016
rect 16436 9976 22732 10016
rect 22772 9976 22781 10016
rect 4919 9871 5305 9890
rect 4919 9848 4985 9871
rect 5071 9848 5153 9871
rect 5239 9848 5305 9871
rect 4919 9808 4928 9848
rect 4968 9808 4985 9848
rect 5071 9808 5092 9848
rect 5132 9808 5153 9848
rect 5239 9808 5256 9848
rect 5296 9808 5305 9848
rect 4919 9785 4985 9808
rect 5071 9785 5153 9808
rect 5239 9785 5305 9808
rect 4919 9766 5305 9785
rect 20039 9871 20425 9890
rect 20039 9848 20105 9871
rect 20191 9848 20273 9871
rect 20359 9848 20425 9871
rect 20039 9808 20048 9848
rect 20088 9808 20105 9848
rect 20191 9808 20212 9848
rect 20252 9808 20273 9848
rect 20359 9808 20376 9848
rect 20416 9808 20425 9848
rect 20039 9785 20105 9808
rect 20191 9785 20273 9808
rect 20359 9785 20425 9808
rect 20039 9766 20425 9785
rect 35159 9871 35545 9890
rect 35159 9848 35225 9871
rect 35311 9848 35393 9871
rect 35479 9848 35545 9871
rect 35159 9808 35168 9848
rect 35208 9808 35225 9848
rect 35311 9808 35332 9848
rect 35372 9808 35393 9848
rect 35479 9808 35496 9848
rect 35536 9808 35545 9848
rect 35159 9785 35225 9808
rect 35311 9785 35393 9808
rect 35479 9785 35545 9808
rect 35159 9766 35545 9785
rect 3679 9115 4065 9134
rect 3679 9092 3745 9115
rect 3831 9092 3913 9115
rect 3999 9092 4065 9115
rect 3679 9052 3688 9092
rect 3728 9052 3745 9092
rect 3831 9052 3852 9092
rect 3892 9052 3913 9092
rect 3999 9052 4016 9092
rect 4056 9052 4065 9092
rect 3679 9029 3745 9052
rect 3831 9029 3913 9052
rect 3999 9029 4065 9052
rect 3679 9010 4065 9029
rect 18799 9115 19185 9134
rect 18799 9092 18865 9115
rect 18951 9092 19033 9115
rect 19119 9092 19185 9115
rect 18799 9052 18808 9092
rect 18848 9052 18865 9092
rect 18951 9052 18972 9092
rect 19012 9052 19033 9092
rect 19119 9052 19136 9092
rect 19176 9052 19185 9092
rect 18799 9029 18865 9052
rect 18951 9029 19033 9052
rect 19119 9029 19185 9052
rect 18799 9010 19185 9029
rect 33919 9115 34305 9134
rect 33919 9092 33985 9115
rect 34071 9092 34153 9115
rect 34239 9092 34305 9115
rect 33919 9052 33928 9092
rect 33968 9052 33985 9092
rect 34071 9052 34092 9092
rect 34132 9052 34153 9092
rect 34239 9052 34256 9092
rect 34296 9052 34305 9092
rect 33919 9029 33985 9052
rect 34071 9029 34153 9052
rect 34239 9029 34305 9052
rect 33919 9010 34305 9029
rect 3715 8632 3724 8672
rect 3764 8632 8812 8672
rect 8852 8632 8861 8672
rect 9763 8632 9772 8672
rect 9812 8632 13036 8672
rect 13076 8632 13085 8672
rect 14851 8548 14860 8588
rect 14900 8548 22252 8588
rect 22292 8548 22301 8588
rect 5347 8464 5356 8504
rect 5396 8464 15820 8504
rect 15860 8464 15869 8504
rect 16387 8464 16396 8504
rect 16436 8464 31372 8504
rect 31412 8464 31421 8504
rect 4919 8359 5305 8378
rect 4919 8336 4985 8359
rect 5071 8336 5153 8359
rect 5239 8336 5305 8359
rect 4919 8296 4928 8336
rect 4968 8296 4985 8336
rect 5071 8296 5092 8336
rect 5132 8296 5153 8336
rect 5239 8296 5256 8336
rect 5296 8296 5305 8336
rect 4919 8273 4985 8296
rect 5071 8273 5153 8296
rect 5239 8273 5305 8296
rect 4919 8254 5305 8273
rect 20039 8359 20425 8378
rect 20039 8336 20105 8359
rect 20191 8336 20273 8359
rect 20359 8336 20425 8359
rect 20039 8296 20048 8336
rect 20088 8296 20105 8336
rect 20191 8296 20212 8336
rect 20252 8296 20273 8336
rect 20359 8296 20376 8336
rect 20416 8296 20425 8336
rect 20039 8273 20105 8296
rect 20191 8273 20273 8296
rect 20359 8273 20425 8296
rect 20039 8254 20425 8273
rect 35159 8359 35545 8378
rect 35159 8336 35225 8359
rect 35311 8336 35393 8359
rect 35479 8336 35545 8359
rect 35159 8296 35168 8336
rect 35208 8296 35225 8336
rect 35311 8296 35332 8336
rect 35372 8296 35393 8336
rect 35479 8296 35496 8336
rect 35536 8296 35545 8336
rect 35159 8273 35225 8296
rect 35311 8273 35393 8296
rect 35479 8273 35545 8296
rect 35159 8254 35545 8273
rect 4579 8128 4588 8168
rect 4628 8128 12364 8168
rect 12404 8128 12413 8168
rect 15811 8128 15820 8168
rect 15860 8128 23308 8168
rect 23348 8128 23357 8168
rect 24067 7876 24076 7916
rect 24116 7876 28012 7916
rect 28052 7876 28061 7916
rect 18883 7792 18892 7832
rect 18932 7792 22636 7832
rect 22676 7792 22685 7832
rect 16963 7708 16972 7748
rect 17012 7708 32620 7748
rect 32660 7708 32669 7748
rect 3679 7603 4065 7622
rect 3679 7580 3745 7603
rect 3831 7580 3913 7603
rect 3999 7580 4065 7603
rect 3679 7540 3688 7580
rect 3728 7540 3745 7580
rect 3831 7540 3852 7580
rect 3892 7540 3913 7580
rect 3999 7540 4016 7580
rect 4056 7540 4065 7580
rect 3679 7517 3745 7540
rect 3831 7517 3913 7540
rect 3999 7517 4065 7540
rect 3679 7498 4065 7517
rect 18799 7603 19185 7622
rect 18799 7580 18865 7603
rect 18951 7580 19033 7603
rect 19119 7580 19185 7603
rect 18799 7540 18808 7580
rect 18848 7540 18865 7580
rect 18951 7540 18972 7580
rect 19012 7540 19033 7580
rect 19119 7540 19136 7580
rect 19176 7540 19185 7580
rect 18799 7517 18865 7540
rect 18951 7517 19033 7540
rect 19119 7517 19185 7540
rect 18799 7498 19185 7517
rect 33919 7603 34305 7622
rect 33919 7580 33985 7603
rect 34071 7580 34153 7603
rect 34239 7580 34305 7603
rect 33919 7540 33928 7580
rect 33968 7540 33985 7580
rect 34071 7540 34092 7580
rect 34132 7540 34153 7580
rect 34239 7540 34256 7580
rect 34296 7540 34305 7580
rect 33919 7517 33985 7540
rect 34071 7517 34153 7540
rect 34239 7517 34305 7540
rect 33919 7498 34305 7517
rect 17635 7372 17644 7412
rect 17684 7372 23884 7412
rect 23924 7372 23933 7412
rect 1891 7288 1900 7328
rect 1940 7288 27820 7328
rect 27860 7288 27869 7328
rect 28960 7288 31948 7328
rect 31988 7288 31997 7328
rect 28960 7244 29000 7288
rect 13795 7204 13804 7244
rect 13844 7204 22828 7244
rect 22868 7204 29000 7244
rect 1603 7120 1612 7160
rect 1652 7120 8044 7160
rect 8084 7120 8093 7160
rect 7555 7036 7564 7076
rect 7604 7036 17644 7076
rect 17684 7036 17693 7076
rect 4919 6847 5305 6866
rect 4919 6824 4985 6847
rect 5071 6824 5153 6847
rect 5239 6824 5305 6847
rect 4919 6784 4928 6824
rect 4968 6784 4985 6824
rect 5071 6784 5092 6824
rect 5132 6784 5153 6824
rect 5239 6784 5256 6824
rect 5296 6784 5305 6824
rect 4919 6761 4985 6784
rect 5071 6761 5153 6784
rect 5239 6761 5305 6784
rect 4919 6742 5305 6761
rect 20039 6847 20425 6866
rect 20039 6824 20105 6847
rect 20191 6824 20273 6847
rect 20359 6824 20425 6847
rect 20039 6784 20048 6824
rect 20088 6784 20105 6824
rect 20191 6784 20212 6824
rect 20252 6784 20273 6824
rect 20359 6784 20376 6824
rect 20416 6784 20425 6824
rect 20039 6761 20105 6784
rect 20191 6761 20273 6784
rect 20359 6761 20425 6784
rect 20039 6742 20425 6761
rect 35159 6847 35545 6866
rect 35159 6824 35225 6847
rect 35311 6824 35393 6847
rect 35479 6824 35545 6847
rect 35159 6784 35168 6824
rect 35208 6784 35225 6824
rect 35311 6784 35332 6824
rect 35372 6784 35393 6824
rect 35479 6784 35496 6824
rect 35536 6784 35545 6824
rect 35159 6761 35225 6784
rect 35311 6761 35393 6784
rect 35479 6761 35545 6784
rect 35159 6742 35545 6761
rect 10723 6364 10732 6404
rect 10772 6364 13900 6404
rect 13940 6364 41260 6404
rect 41300 6364 41309 6404
rect 13987 6280 13996 6320
rect 14036 6280 20044 6320
rect 20084 6280 20093 6320
rect 20372 6280 37820 6320
rect 13027 6196 13036 6236
rect 13076 6196 20236 6236
rect 20276 6196 20285 6236
rect 20372 6152 20412 6280
rect 37780 6236 37820 6280
rect 37780 6196 40204 6236
rect 40244 6196 40253 6236
rect 20035 6112 20044 6152
rect 20084 6112 20412 6152
rect 3679 6091 4065 6110
rect 3679 6068 3745 6091
rect 3831 6068 3913 6091
rect 3999 6068 4065 6091
rect 3679 6028 3688 6068
rect 3728 6028 3745 6068
rect 3831 6028 3852 6068
rect 3892 6028 3913 6068
rect 3999 6028 4016 6068
rect 4056 6028 4065 6068
rect 3679 6005 3745 6028
rect 3831 6005 3913 6028
rect 3999 6005 4065 6028
rect 3679 5986 4065 6005
rect 18799 6091 19185 6110
rect 18799 6068 18865 6091
rect 18951 6068 19033 6091
rect 19119 6068 19185 6091
rect 18799 6028 18808 6068
rect 18848 6028 18865 6068
rect 18951 6028 18972 6068
rect 19012 6028 19033 6068
rect 19119 6028 19136 6068
rect 19176 6028 19185 6068
rect 18799 6005 18865 6028
rect 18951 6005 19033 6028
rect 19119 6005 19185 6028
rect 18799 5986 19185 6005
rect 33919 6091 34305 6110
rect 33919 6068 33985 6091
rect 34071 6068 34153 6091
rect 34239 6068 34305 6091
rect 33919 6028 33928 6068
rect 33968 6028 33985 6068
rect 34071 6028 34092 6068
rect 34132 6028 34153 6068
rect 34239 6028 34256 6068
rect 34296 6028 34305 6068
rect 33919 6005 33985 6028
rect 34071 6005 34153 6028
rect 34239 6005 34305 6028
rect 33919 5986 34305 6005
rect 20227 5944 20236 5984
rect 20276 5944 29000 5984
rect 28960 5900 29000 5944
rect 14179 5860 14188 5900
rect 14228 5860 27916 5900
rect 27956 5860 27965 5900
rect 28960 5860 40876 5900
rect 40916 5860 40925 5900
rect 15619 5776 15628 5816
rect 15668 5776 30988 5816
rect 31028 5776 31037 5816
rect 16099 5608 16108 5648
rect 16148 5608 20716 5648
rect 20756 5608 20765 5648
rect 12643 5440 12652 5480
rect 12692 5440 28300 5480
rect 28340 5440 28349 5480
rect 4919 5335 5305 5354
rect 4919 5312 4985 5335
rect 5071 5312 5153 5335
rect 5239 5312 5305 5335
rect 4919 5272 4928 5312
rect 4968 5272 4985 5312
rect 5071 5272 5092 5312
rect 5132 5272 5153 5312
rect 5239 5272 5256 5312
rect 5296 5272 5305 5312
rect 4919 5249 4985 5272
rect 5071 5249 5153 5272
rect 5239 5249 5305 5272
rect 4919 5230 5305 5249
rect 20039 5335 20425 5354
rect 20039 5312 20105 5335
rect 20191 5312 20273 5335
rect 20359 5312 20425 5335
rect 20039 5272 20048 5312
rect 20088 5272 20105 5312
rect 20191 5272 20212 5312
rect 20252 5272 20273 5312
rect 20359 5272 20376 5312
rect 20416 5272 20425 5312
rect 20039 5249 20105 5272
rect 20191 5249 20273 5272
rect 20359 5249 20425 5272
rect 20039 5230 20425 5249
rect 35159 5335 35545 5354
rect 35159 5312 35225 5335
rect 35311 5312 35393 5335
rect 35479 5312 35545 5335
rect 35159 5272 35168 5312
rect 35208 5272 35225 5312
rect 35311 5272 35332 5312
rect 35372 5272 35393 5312
rect 35479 5272 35496 5312
rect 35536 5272 35545 5312
rect 35159 5249 35225 5272
rect 35311 5249 35393 5272
rect 35479 5249 35545 5272
rect 35159 5230 35545 5249
rect 1699 4936 1708 4976
rect 1748 4936 19372 4976
rect 19412 4936 19421 4976
rect 10339 4852 10348 4892
rect 10388 4852 33772 4892
rect 33812 4852 33821 4892
rect 1219 4768 1228 4808
rect 1268 4768 7564 4808
rect 7604 4768 7613 4808
rect 18115 4768 18124 4808
rect 18164 4768 36652 4808
rect 36692 4768 36701 4808
rect 12643 4684 12652 4724
rect 12692 4684 40492 4724
rect 40532 4684 40541 4724
rect 3679 4579 4065 4598
rect 3679 4556 3745 4579
rect 3831 4556 3913 4579
rect 3999 4556 4065 4579
rect 3679 4516 3688 4556
rect 3728 4516 3745 4556
rect 3831 4516 3852 4556
rect 3892 4516 3913 4556
rect 3999 4516 4016 4556
rect 4056 4516 4065 4556
rect 3679 4493 3745 4516
rect 3831 4493 3913 4516
rect 3999 4493 4065 4516
rect 3679 4474 4065 4493
rect 18799 4579 19185 4598
rect 18799 4556 18865 4579
rect 18951 4556 19033 4579
rect 19119 4556 19185 4579
rect 18799 4516 18808 4556
rect 18848 4516 18865 4556
rect 18951 4516 18972 4556
rect 19012 4516 19033 4556
rect 19119 4516 19136 4556
rect 19176 4516 19185 4556
rect 18799 4493 18865 4516
rect 18951 4493 19033 4516
rect 19119 4493 19185 4516
rect 18799 4474 19185 4493
rect 33919 4579 34305 4598
rect 33919 4556 33985 4579
rect 34071 4556 34153 4579
rect 34239 4556 34305 4579
rect 33919 4516 33928 4556
rect 33968 4516 33985 4556
rect 34071 4516 34092 4556
rect 34132 4516 34153 4556
rect 34239 4516 34256 4556
rect 34296 4516 34305 4556
rect 33919 4493 33985 4516
rect 34071 4493 34153 4516
rect 34239 4493 34305 4516
rect 33919 4474 34305 4493
rect 16771 4012 16780 4052
rect 16820 4012 33964 4052
rect 34004 4012 34013 4052
rect 18691 3928 18700 3968
rect 18740 3928 36844 3968
rect 36884 3928 36893 3968
rect 4919 3823 5305 3842
rect 4919 3800 4985 3823
rect 5071 3800 5153 3823
rect 5239 3800 5305 3823
rect 4919 3760 4928 3800
rect 4968 3760 4985 3800
rect 5071 3760 5092 3800
rect 5132 3760 5153 3800
rect 5239 3760 5256 3800
rect 5296 3760 5305 3800
rect 4919 3737 4985 3760
rect 5071 3737 5153 3760
rect 5239 3737 5305 3760
rect 4919 3718 5305 3737
rect 20039 3823 20425 3842
rect 20039 3800 20105 3823
rect 20191 3800 20273 3823
rect 20359 3800 20425 3823
rect 20039 3760 20048 3800
rect 20088 3760 20105 3800
rect 20191 3760 20212 3800
rect 20252 3760 20273 3800
rect 20359 3760 20376 3800
rect 20416 3760 20425 3800
rect 20039 3737 20105 3760
rect 20191 3737 20273 3760
rect 20359 3737 20425 3760
rect 20039 3718 20425 3737
rect 35159 3823 35545 3842
rect 35159 3800 35225 3823
rect 35311 3800 35393 3823
rect 35479 3800 35545 3823
rect 35159 3760 35168 3800
rect 35208 3760 35225 3800
rect 35311 3760 35332 3800
rect 35372 3760 35393 3800
rect 35479 3760 35496 3800
rect 35536 3760 35545 3800
rect 35159 3737 35225 3760
rect 35311 3737 35393 3760
rect 35479 3737 35545 3760
rect 35159 3718 35545 3737
rect 15235 3592 15244 3632
rect 15284 3592 31756 3632
rect 31796 3592 31805 3632
rect 16003 3508 16012 3548
rect 16052 3508 31372 3548
rect 31412 3508 31421 3548
rect 12259 3424 12268 3464
rect 12308 3424 19948 3464
rect 19988 3424 19997 3464
rect 19363 3340 19372 3380
rect 19412 3340 33388 3380
rect 33428 3340 33437 3380
rect 11011 3256 11020 3296
rect 11060 3256 29548 3296
rect 29588 3256 29597 3296
rect 15427 3172 15436 3212
rect 15476 3172 28780 3212
rect 28820 3172 28829 3212
rect 3679 3067 4065 3086
rect 3679 3044 3745 3067
rect 3831 3044 3913 3067
rect 3999 3044 4065 3067
rect 3679 3004 3688 3044
rect 3728 3004 3745 3044
rect 3831 3004 3852 3044
rect 3892 3004 3913 3044
rect 3999 3004 4016 3044
rect 4056 3004 4065 3044
rect 3679 2981 3745 3004
rect 3831 2981 3913 3004
rect 3999 2981 4065 3004
rect 3679 2962 4065 2981
rect 18799 3067 19185 3086
rect 18799 3044 18865 3067
rect 18951 3044 19033 3067
rect 19119 3044 19185 3067
rect 18799 3004 18808 3044
rect 18848 3004 18865 3044
rect 18951 3004 18972 3044
rect 19012 3004 19033 3044
rect 19119 3004 19136 3044
rect 19176 3004 19185 3044
rect 18799 2981 18865 3004
rect 18951 2981 19033 3004
rect 19119 2981 19185 3004
rect 18799 2962 19185 2981
rect 33919 3067 34305 3086
rect 33919 3044 33985 3067
rect 34071 3044 34153 3067
rect 34239 3044 34305 3067
rect 33919 3004 33928 3044
rect 33968 3004 33985 3044
rect 34071 3004 34092 3044
rect 34132 3004 34153 3044
rect 34239 3004 34256 3044
rect 34296 3004 34305 3044
rect 33919 2981 33985 3004
rect 34071 2981 34153 3004
rect 34239 2981 34305 3004
rect 33919 2962 34305 2981
rect 10243 2416 10252 2456
rect 10292 2416 35692 2456
rect 35732 2416 35741 2456
rect 4919 2311 5305 2330
rect 4919 2288 4985 2311
rect 5071 2288 5153 2311
rect 5239 2288 5305 2311
rect 4919 2248 4928 2288
rect 4968 2248 4985 2288
rect 5071 2248 5092 2288
rect 5132 2248 5153 2288
rect 5239 2248 5256 2288
rect 5296 2248 5305 2288
rect 4919 2225 4985 2248
rect 5071 2225 5153 2248
rect 5239 2225 5305 2248
rect 4919 2206 5305 2225
rect 20039 2311 20425 2330
rect 20039 2288 20105 2311
rect 20191 2288 20273 2311
rect 20359 2288 20425 2311
rect 20039 2248 20048 2288
rect 20088 2248 20105 2288
rect 20191 2248 20212 2288
rect 20252 2248 20273 2288
rect 20359 2248 20376 2288
rect 20416 2248 20425 2288
rect 20039 2225 20105 2248
rect 20191 2225 20273 2248
rect 20359 2225 20425 2248
rect 20039 2206 20425 2225
rect 35159 2311 35545 2330
rect 35159 2288 35225 2311
rect 35311 2288 35393 2311
rect 35479 2288 35545 2311
rect 35159 2248 35168 2288
rect 35208 2248 35225 2288
rect 35311 2248 35332 2288
rect 35372 2248 35393 2288
rect 35479 2248 35496 2288
rect 35536 2248 35545 2288
rect 35159 2225 35225 2248
rect 35311 2225 35393 2248
rect 35479 2225 35545 2248
rect 35159 2206 35545 2225
rect 14083 2080 14092 2120
rect 14132 2080 37612 2120
rect 37652 2080 37661 2120
rect 11779 1996 11788 2036
rect 11828 1996 30220 2036
rect 30260 1996 30269 2036
rect 18019 1912 18028 1952
rect 18068 1912 29548 1952
rect 29588 1912 29597 1952
rect 12067 1828 12076 1868
rect 12116 1828 27724 1868
rect 27764 1828 27773 1868
rect 3679 1555 4065 1574
rect 3679 1532 3745 1555
rect 3831 1532 3913 1555
rect 3999 1532 4065 1555
rect 3679 1492 3688 1532
rect 3728 1492 3745 1532
rect 3831 1492 3852 1532
rect 3892 1492 3913 1532
rect 3999 1492 4016 1532
rect 4056 1492 4065 1532
rect 3679 1469 3745 1492
rect 3831 1469 3913 1492
rect 3999 1469 4065 1492
rect 3679 1450 4065 1469
rect 18799 1555 19185 1574
rect 18799 1532 18865 1555
rect 18951 1532 19033 1555
rect 19119 1532 19185 1555
rect 18799 1492 18808 1532
rect 18848 1492 18865 1532
rect 18951 1492 18972 1532
rect 19012 1492 19033 1532
rect 19119 1492 19136 1532
rect 19176 1492 19185 1532
rect 18799 1469 18865 1492
rect 18951 1469 19033 1492
rect 19119 1469 19185 1492
rect 18799 1450 19185 1469
rect 33919 1555 34305 1574
rect 33919 1532 33985 1555
rect 34071 1532 34153 1555
rect 34239 1532 34305 1555
rect 33919 1492 33928 1532
rect 33968 1492 33985 1532
rect 34071 1492 34092 1532
rect 34132 1492 34153 1532
rect 34239 1492 34256 1532
rect 34296 1492 34305 1532
rect 33919 1469 33985 1492
rect 34071 1469 34153 1492
rect 34239 1469 34305 1492
rect 33919 1450 34305 1469
rect 19939 1156 19948 1196
rect 19988 1156 40876 1196
rect 40916 1156 40925 1196
rect 14467 1072 14476 1112
rect 14516 1072 39724 1112
rect 39764 1072 39773 1112
rect 9763 988 9772 1028
rect 9812 988 25420 1028
rect 25460 988 35596 1028
rect 35636 988 35645 1028
rect 15523 904 15532 944
rect 15572 904 40300 944
rect 40340 904 40349 944
rect 4919 799 5305 818
rect 4919 776 4985 799
rect 5071 776 5153 799
rect 5239 776 5305 799
rect 4919 736 4928 776
rect 4968 736 4985 776
rect 5071 736 5092 776
rect 5132 736 5153 776
rect 5239 736 5256 776
rect 5296 736 5305 776
rect 4919 713 4985 736
rect 5071 713 5153 736
rect 5239 713 5305 736
rect 4919 694 5305 713
rect 20039 799 20425 818
rect 20039 776 20105 799
rect 20191 776 20273 799
rect 20359 776 20425 799
rect 20039 736 20048 776
rect 20088 736 20105 776
rect 20191 736 20212 776
rect 20252 736 20273 776
rect 20359 736 20376 776
rect 20416 736 20425 776
rect 20039 713 20105 736
rect 20191 713 20273 736
rect 20359 713 20425 736
rect 20039 694 20425 713
rect 35159 799 35545 818
rect 35159 776 35225 799
rect 35311 776 35393 799
rect 35479 776 35545 799
rect 35159 736 35168 776
rect 35208 736 35225 776
rect 35311 736 35332 776
rect 35372 736 35393 776
rect 35479 736 35496 776
rect 35536 736 35545 776
rect 35159 713 35225 736
rect 35311 713 35393 736
rect 35479 713 35545 736
rect 35159 694 35545 713
rect 2467 568 2476 608
rect 2516 568 25804 608
rect 25844 568 25853 608
<< via5 >>
rect 4985 9848 5071 9871
rect 5153 9848 5239 9871
rect 4985 9808 5010 9848
rect 5010 9808 5050 9848
rect 5050 9808 5071 9848
rect 5153 9808 5174 9848
rect 5174 9808 5214 9848
rect 5214 9808 5239 9848
rect 4985 9785 5071 9808
rect 5153 9785 5239 9808
rect 20105 9848 20191 9871
rect 20273 9848 20359 9871
rect 20105 9808 20130 9848
rect 20130 9808 20170 9848
rect 20170 9808 20191 9848
rect 20273 9808 20294 9848
rect 20294 9808 20334 9848
rect 20334 9808 20359 9848
rect 20105 9785 20191 9808
rect 20273 9785 20359 9808
rect 35225 9848 35311 9871
rect 35393 9848 35479 9871
rect 35225 9808 35250 9848
rect 35250 9808 35290 9848
rect 35290 9808 35311 9848
rect 35393 9808 35414 9848
rect 35414 9808 35454 9848
rect 35454 9808 35479 9848
rect 35225 9785 35311 9808
rect 35393 9785 35479 9808
rect 3745 9092 3831 9115
rect 3913 9092 3999 9115
rect 3745 9052 3770 9092
rect 3770 9052 3810 9092
rect 3810 9052 3831 9092
rect 3913 9052 3934 9092
rect 3934 9052 3974 9092
rect 3974 9052 3999 9092
rect 3745 9029 3831 9052
rect 3913 9029 3999 9052
rect 18865 9092 18951 9115
rect 19033 9092 19119 9115
rect 18865 9052 18890 9092
rect 18890 9052 18930 9092
rect 18930 9052 18951 9092
rect 19033 9052 19054 9092
rect 19054 9052 19094 9092
rect 19094 9052 19119 9092
rect 18865 9029 18951 9052
rect 19033 9029 19119 9052
rect 33985 9092 34071 9115
rect 34153 9092 34239 9115
rect 33985 9052 34010 9092
rect 34010 9052 34050 9092
rect 34050 9052 34071 9092
rect 34153 9052 34174 9092
rect 34174 9052 34214 9092
rect 34214 9052 34239 9092
rect 33985 9029 34071 9052
rect 34153 9029 34239 9052
rect 4985 8336 5071 8359
rect 5153 8336 5239 8359
rect 4985 8296 5010 8336
rect 5010 8296 5050 8336
rect 5050 8296 5071 8336
rect 5153 8296 5174 8336
rect 5174 8296 5214 8336
rect 5214 8296 5239 8336
rect 4985 8273 5071 8296
rect 5153 8273 5239 8296
rect 20105 8336 20191 8359
rect 20273 8336 20359 8359
rect 20105 8296 20130 8336
rect 20130 8296 20170 8336
rect 20170 8296 20191 8336
rect 20273 8296 20294 8336
rect 20294 8296 20334 8336
rect 20334 8296 20359 8336
rect 20105 8273 20191 8296
rect 20273 8273 20359 8296
rect 35225 8336 35311 8359
rect 35393 8336 35479 8359
rect 35225 8296 35250 8336
rect 35250 8296 35290 8336
rect 35290 8296 35311 8336
rect 35393 8296 35414 8336
rect 35414 8296 35454 8336
rect 35454 8296 35479 8336
rect 35225 8273 35311 8296
rect 35393 8273 35479 8296
rect 3745 7580 3831 7603
rect 3913 7580 3999 7603
rect 3745 7540 3770 7580
rect 3770 7540 3810 7580
rect 3810 7540 3831 7580
rect 3913 7540 3934 7580
rect 3934 7540 3974 7580
rect 3974 7540 3999 7580
rect 3745 7517 3831 7540
rect 3913 7517 3999 7540
rect 18865 7580 18951 7603
rect 19033 7580 19119 7603
rect 18865 7540 18890 7580
rect 18890 7540 18930 7580
rect 18930 7540 18951 7580
rect 19033 7540 19054 7580
rect 19054 7540 19094 7580
rect 19094 7540 19119 7580
rect 18865 7517 18951 7540
rect 19033 7517 19119 7540
rect 33985 7580 34071 7603
rect 34153 7580 34239 7603
rect 33985 7540 34010 7580
rect 34010 7540 34050 7580
rect 34050 7540 34071 7580
rect 34153 7540 34174 7580
rect 34174 7540 34214 7580
rect 34214 7540 34239 7580
rect 33985 7517 34071 7540
rect 34153 7517 34239 7540
rect 4985 6824 5071 6847
rect 5153 6824 5239 6847
rect 4985 6784 5010 6824
rect 5010 6784 5050 6824
rect 5050 6784 5071 6824
rect 5153 6784 5174 6824
rect 5174 6784 5214 6824
rect 5214 6784 5239 6824
rect 4985 6761 5071 6784
rect 5153 6761 5239 6784
rect 20105 6824 20191 6847
rect 20273 6824 20359 6847
rect 20105 6784 20130 6824
rect 20130 6784 20170 6824
rect 20170 6784 20191 6824
rect 20273 6784 20294 6824
rect 20294 6784 20334 6824
rect 20334 6784 20359 6824
rect 20105 6761 20191 6784
rect 20273 6761 20359 6784
rect 35225 6824 35311 6847
rect 35393 6824 35479 6847
rect 35225 6784 35250 6824
rect 35250 6784 35290 6824
rect 35290 6784 35311 6824
rect 35393 6784 35414 6824
rect 35414 6784 35454 6824
rect 35454 6784 35479 6824
rect 35225 6761 35311 6784
rect 35393 6761 35479 6784
rect 3745 6068 3831 6091
rect 3913 6068 3999 6091
rect 3745 6028 3770 6068
rect 3770 6028 3810 6068
rect 3810 6028 3831 6068
rect 3913 6028 3934 6068
rect 3934 6028 3974 6068
rect 3974 6028 3999 6068
rect 3745 6005 3831 6028
rect 3913 6005 3999 6028
rect 18865 6068 18951 6091
rect 19033 6068 19119 6091
rect 18865 6028 18890 6068
rect 18890 6028 18930 6068
rect 18930 6028 18951 6068
rect 19033 6028 19054 6068
rect 19054 6028 19094 6068
rect 19094 6028 19119 6068
rect 18865 6005 18951 6028
rect 19033 6005 19119 6028
rect 33985 6068 34071 6091
rect 34153 6068 34239 6091
rect 33985 6028 34010 6068
rect 34010 6028 34050 6068
rect 34050 6028 34071 6068
rect 34153 6028 34174 6068
rect 34174 6028 34214 6068
rect 34214 6028 34239 6068
rect 33985 6005 34071 6028
rect 34153 6005 34239 6028
rect 4985 5312 5071 5335
rect 5153 5312 5239 5335
rect 4985 5272 5010 5312
rect 5010 5272 5050 5312
rect 5050 5272 5071 5312
rect 5153 5272 5174 5312
rect 5174 5272 5214 5312
rect 5214 5272 5239 5312
rect 4985 5249 5071 5272
rect 5153 5249 5239 5272
rect 20105 5312 20191 5335
rect 20273 5312 20359 5335
rect 20105 5272 20130 5312
rect 20130 5272 20170 5312
rect 20170 5272 20191 5312
rect 20273 5272 20294 5312
rect 20294 5272 20334 5312
rect 20334 5272 20359 5312
rect 20105 5249 20191 5272
rect 20273 5249 20359 5272
rect 35225 5312 35311 5335
rect 35393 5312 35479 5335
rect 35225 5272 35250 5312
rect 35250 5272 35290 5312
rect 35290 5272 35311 5312
rect 35393 5272 35414 5312
rect 35414 5272 35454 5312
rect 35454 5272 35479 5312
rect 35225 5249 35311 5272
rect 35393 5249 35479 5272
rect 3745 4556 3831 4579
rect 3913 4556 3999 4579
rect 3745 4516 3770 4556
rect 3770 4516 3810 4556
rect 3810 4516 3831 4556
rect 3913 4516 3934 4556
rect 3934 4516 3974 4556
rect 3974 4516 3999 4556
rect 3745 4493 3831 4516
rect 3913 4493 3999 4516
rect 18865 4556 18951 4579
rect 19033 4556 19119 4579
rect 18865 4516 18890 4556
rect 18890 4516 18930 4556
rect 18930 4516 18951 4556
rect 19033 4516 19054 4556
rect 19054 4516 19094 4556
rect 19094 4516 19119 4556
rect 18865 4493 18951 4516
rect 19033 4493 19119 4516
rect 33985 4556 34071 4579
rect 34153 4556 34239 4579
rect 33985 4516 34010 4556
rect 34010 4516 34050 4556
rect 34050 4516 34071 4556
rect 34153 4516 34174 4556
rect 34174 4516 34214 4556
rect 34214 4516 34239 4556
rect 33985 4493 34071 4516
rect 34153 4493 34239 4516
rect 4985 3800 5071 3823
rect 5153 3800 5239 3823
rect 4985 3760 5010 3800
rect 5010 3760 5050 3800
rect 5050 3760 5071 3800
rect 5153 3760 5174 3800
rect 5174 3760 5214 3800
rect 5214 3760 5239 3800
rect 4985 3737 5071 3760
rect 5153 3737 5239 3760
rect 20105 3800 20191 3823
rect 20273 3800 20359 3823
rect 20105 3760 20130 3800
rect 20130 3760 20170 3800
rect 20170 3760 20191 3800
rect 20273 3760 20294 3800
rect 20294 3760 20334 3800
rect 20334 3760 20359 3800
rect 20105 3737 20191 3760
rect 20273 3737 20359 3760
rect 35225 3800 35311 3823
rect 35393 3800 35479 3823
rect 35225 3760 35250 3800
rect 35250 3760 35290 3800
rect 35290 3760 35311 3800
rect 35393 3760 35414 3800
rect 35414 3760 35454 3800
rect 35454 3760 35479 3800
rect 35225 3737 35311 3760
rect 35393 3737 35479 3760
rect 3745 3044 3831 3067
rect 3913 3044 3999 3067
rect 3745 3004 3770 3044
rect 3770 3004 3810 3044
rect 3810 3004 3831 3044
rect 3913 3004 3934 3044
rect 3934 3004 3974 3044
rect 3974 3004 3999 3044
rect 3745 2981 3831 3004
rect 3913 2981 3999 3004
rect 18865 3044 18951 3067
rect 19033 3044 19119 3067
rect 18865 3004 18890 3044
rect 18890 3004 18930 3044
rect 18930 3004 18951 3044
rect 19033 3004 19054 3044
rect 19054 3004 19094 3044
rect 19094 3004 19119 3044
rect 18865 2981 18951 3004
rect 19033 2981 19119 3004
rect 33985 3044 34071 3067
rect 34153 3044 34239 3067
rect 33985 3004 34010 3044
rect 34010 3004 34050 3044
rect 34050 3004 34071 3044
rect 34153 3004 34174 3044
rect 34174 3004 34214 3044
rect 34214 3004 34239 3044
rect 33985 2981 34071 3004
rect 34153 2981 34239 3004
rect 4985 2288 5071 2311
rect 5153 2288 5239 2311
rect 4985 2248 5010 2288
rect 5010 2248 5050 2288
rect 5050 2248 5071 2288
rect 5153 2248 5174 2288
rect 5174 2248 5214 2288
rect 5214 2248 5239 2288
rect 4985 2225 5071 2248
rect 5153 2225 5239 2248
rect 20105 2288 20191 2311
rect 20273 2288 20359 2311
rect 20105 2248 20130 2288
rect 20130 2248 20170 2288
rect 20170 2248 20191 2288
rect 20273 2248 20294 2288
rect 20294 2248 20334 2288
rect 20334 2248 20359 2288
rect 20105 2225 20191 2248
rect 20273 2225 20359 2248
rect 35225 2288 35311 2311
rect 35393 2288 35479 2311
rect 35225 2248 35250 2288
rect 35250 2248 35290 2288
rect 35290 2248 35311 2288
rect 35393 2248 35414 2288
rect 35414 2248 35454 2288
rect 35454 2248 35479 2288
rect 35225 2225 35311 2248
rect 35393 2225 35479 2248
rect 3745 1532 3831 1555
rect 3913 1532 3999 1555
rect 3745 1492 3770 1532
rect 3770 1492 3810 1532
rect 3810 1492 3831 1532
rect 3913 1492 3934 1532
rect 3934 1492 3974 1532
rect 3974 1492 3999 1532
rect 3745 1469 3831 1492
rect 3913 1469 3999 1492
rect 18865 1532 18951 1555
rect 19033 1532 19119 1555
rect 18865 1492 18890 1532
rect 18890 1492 18930 1532
rect 18930 1492 18951 1532
rect 19033 1492 19054 1532
rect 19054 1492 19094 1532
rect 19094 1492 19119 1532
rect 18865 1469 18951 1492
rect 19033 1469 19119 1492
rect 33985 1532 34071 1555
rect 34153 1532 34239 1555
rect 33985 1492 34010 1532
rect 34010 1492 34050 1532
rect 34050 1492 34071 1532
rect 34153 1492 34174 1532
rect 34174 1492 34214 1532
rect 34214 1492 34239 1532
rect 33985 1469 34071 1492
rect 34153 1469 34239 1492
rect 4985 776 5071 799
rect 5153 776 5239 799
rect 4985 736 5010 776
rect 5010 736 5050 776
rect 5050 736 5071 776
rect 5153 736 5174 776
rect 5174 736 5214 776
rect 5214 736 5239 776
rect 4985 713 5071 736
rect 5153 713 5239 736
rect 20105 776 20191 799
rect 20273 776 20359 799
rect 20105 736 20130 776
rect 20130 736 20170 776
rect 20170 736 20191 776
rect 20273 736 20294 776
rect 20294 736 20334 776
rect 20334 736 20359 776
rect 20105 713 20191 736
rect 20273 713 20359 736
rect 35225 776 35311 799
rect 35393 776 35479 799
rect 35225 736 35250 776
rect 35250 736 35290 776
rect 35290 736 35311 776
rect 35393 736 35414 776
rect 35414 736 35454 776
rect 35454 736 35479 776
rect 35225 713 35311 736
rect 35393 713 35479 736
<< metal6 >>
rect 3652 9115 4092 10752
rect 3652 9029 3745 9115
rect 3831 9029 3913 9115
rect 3999 9029 4092 9115
rect 3652 7603 4092 9029
rect 3652 7517 3745 7603
rect 3831 7517 3913 7603
rect 3999 7517 4092 7603
rect 3652 6091 4092 7517
rect 3652 6005 3745 6091
rect 3831 6005 3913 6091
rect 3999 6005 4092 6091
rect 3652 4579 4092 6005
rect 3652 4493 3745 4579
rect 3831 4493 3913 4579
rect 3999 4493 4092 4579
rect 3652 3067 4092 4493
rect 3652 2981 3745 3067
rect 3831 2981 3913 3067
rect 3999 2981 4092 3067
rect 3652 1555 4092 2981
rect 3652 1469 3745 1555
rect 3831 1469 3913 1555
rect 3999 1469 4092 1555
rect 3652 0 4092 1469
rect 4892 9871 5332 10752
rect 4892 9785 4985 9871
rect 5071 9785 5153 9871
rect 5239 9785 5332 9871
rect 4892 8359 5332 9785
rect 4892 8273 4985 8359
rect 5071 8273 5153 8359
rect 5239 8273 5332 8359
rect 4892 6847 5332 8273
rect 4892 6761 4985 6847
rect 5071 6761 5153 6847
rect 5239 6761 5332 6847
rect 4892 5335 5332 6761
rect 4892 5249 4985 5335
rect 5071 5249 5153 5335
rect 5239 5249 5332 5335
rect 4892 3823 5332 5249
rect 4892 3737 4985 3823
rect 5071 3737 5153 3823
rect 5239 3737 5332 3823
rect 4892 2311 5332 3737
rect 4892 2225 4985 2311
rect 5071 2225 5153 2311
rect 5239 2225 5332 2311
rect 4892 799 5332 2225
rect 4892 713 4985 799
rect 5071 713 5153 799
rect 5239 713 5332 799
rect 4892 0 5332 713
rect 18772 9115 19212 10752
rect 18772 9029 18865 9115
rect 18951 9029 19033 9115
rect 19119 9029 19212 9115
rect 18772 7603 19212 9029
rect 18772 7517 18865 7603
rect 18951 7517 19033 7603
rect 19119 7517 19212 7603
rect 18772 6091 19212 7517
rect 18772 6005 18865 6091
rect 18951 6005 19033 6091
rect 19119 6005 19212 6091
rect 18772 4579 19212 6005
rect 18772 4493 18865 4579
rect 18951 4493 19033 4579
rect 19119 4493 19212 4579
rect 18772 3067 19212 4493
rect 18772 2981 18865 3067
rect 18951 2981 19033 3067
rect 19119 2981 19212 3067
rect 18772 1555 19212 2981
rect 18772 1469 18865 1555
rect 18951 1469 19033 1555
rect 19119 1469 19212 1555
rect 18772 0 19212 1469
rect 20012 9871 20452 10752
rect 20012 9785 20105 9871
rect 20191 9785 20273 9871
rect 20359 9785 20452 9871
rect 20012 8359 20452 9785
rect 20012 8273 20105 8359
rect 20191 8273 20273 8359
rect 20359 8273 20452 8359
rect 20012 6847 20452 8273
rect 20012 6761 20105 6847
rect 20191 6761 20273 6847
rect 20359 6761 20452 6847
rect 20012 5335 20452 6761
rect 20012 5249 20105 5335
rect 20191 5249 20273 5335
rect 20359 5249 20452 5335
rect 20012 3823 20452 5249
rect 20012 3737 20105 3823
rect 20191 3737 20273 3823
rect 20359 3737 20452 3823
rect 20012 2311 20452 3737
rect 20012 2225 20105 2311
rect 20191 2225 20273 2311
rect 20359 2225 20452 2311
rect 20012 799 20452 2225
rect 20012 713 20105 799
rect 20191 713 20273 799
rect 20359 713 20452 799
rect 20012 0 20452 713
rect 33892 9115 34332 10752
rect 33892 9029 33985 9115
rect 34071 9029 34153 9115
rect 34239 9029 34332 9115
rect 33892 7603 34332 9029
rect 33892 7517 33985 7603
rect 34071 7517 34153 7603
rect 34239 7517 34332 7603
rect 33892 6091 34332 7517
rect 33892 6005 33985 6091
rect 34071 6005 34153 6091
rect 34239 6005 34332 6091
rect 33892 4579 34332 6005
rect 33892 4493 33985 4579
rect 34071 4493 34153 4579
rect 34239 4493 34332 4579
rect 33892 3067 34332 4493
rect 33892 2981 33985 3067
rect 34071 2981 34153 3067
rect 34239 2981 34332 3067
rect 33892 1555 34332 2981
rect 33892 1469 33985 1555
rect 34071 1469 34153 1555
rect 34239 1469 34332 1555
rect 33892 0 34332 1469
rect 35132 9871 35572 10752
rect 35132 9785 35225 9871
rect 35311 9785 35393 9871
rect 35479 9785 35572 9871
rect 35132 8359 35572 9785
rect 35132 8273 35225 8359
rect 35311 8273 35393 8359
rect 35479 8273 35572 8359
rect 35132 6847 35572 8273
rect 35132 6761 35225 6847
rect 35311 6761 35393 6847
rect 35479 6761 35572 6847
rect 35132 5335 35572 6761
rect 35132 5249 35225 5335
rect 35311 5249 35393 5335
rect 35479 5249 35572 5335
rect 35132 3823 35572 5249
rect 35132 3737 35225 3823
rect 35311 3737 35393 3823
rect 35479 3737 35572 3823
rect 35132 2311 35572 3737
rect 35132 2225 35225 2311
rect 35311 2225 35393 2311
rect 35479 2225 35572 2311
rect 35132 799 35572 2225
rect 35132 713 35225 799
rect 35311 713 35393 799
rect 35479 713 35572 799
rect 35132 0 35572 713
use sg13g2_mux4_1  _047_
timestamp 1677257233
transform 1 0 35520 0 1 8316
box -48 -56 2064 834
use sg13g2_mux4_1  _048_
timestamp 1677257233
transform 1 0 21408 0 -1 6804
box -48 -56 2064 834
use sg13g2_mux4_1  _049_
timestamp 1677257233
transform 1 0 25632 0 -1 8316
box -48 -56 2064 834
use sg13g2_mux4_1  _050_
timestamp 1677257233
transform 1 0 10752 0 1 3780
box -48 -56 2064 834
use sg13g2_mux4_1  _051_
timestamp 1677257233
transform 1 0 37728 0 1 3780
box -48 -56 2064 834
use sg13g2_mux4_1  _052_
timestamp 1677257233
transform 1 0 22560 0 -1 3780
box -48 -56 2064 834
use sg13g2_mux4_1  _053_
timestamp 1677257233
transform 1 0 26976 0 -1 5292
box -48 -56 2064 834
use sg13g2_mux4_1  _054_
timestamp 1677257233
transform 1 0 9600 0 -1 3780
box -48 -56 2064 834
use sg13g2_mux4_1  _055_
timestamp 1677257233
transform 1 0 36192 0 1 5292
box -48 -56 2064 834
use sg13g2_mux4_1  _056_
timestamp 1677257233
transform 1 0 21216 0 -1 5292
box -48 -56 2064 834
use sg13g2_mux4_1  _057_
timestamp 1677257233
transform 1 0 25824 0 1 8316
box -48 -56 2064 834
use sg13g2_mux4_1  _058_
timestamp 1677257233
transform 1 0 10656 0 1 8316
box -48 -56 2064 834
use sg13g2_mux4_1  _059_
timestamp 1677257233
transform 1 0 32160 0 1 8316
box -48 -56 2064 834
use sg13g2_mux4_1  _060_
timestamp 1677257233
transform 1 0 22272 0 1 8316
box -48 -56 2064 834
use sg13g2_mux4_1  _061_
timestamp 1677257233
transform 1 0 26976 0 -1 6804
box -48 -56 2064 834
use sg13g2_mux4_1  _062_
timestamp 1677257233
transform 1 0 9312 0 -1 5292
box -48 -56 2064 834
use sg13g2_mux4_1  _063_
timestamp 1677257233
transform 1 0 34176 0 1 5292
box -48 -56 2064 834
use sg13g2_mux2_1  _064_
timestamp 1677247768
transform -1 0 20832 0 1 5292
box -48 -56 1008 834
use sg13g2_mux2_1  _065_
timestamp 1677247768
transform 1 0 9024 0 -1 6804
box -48 -56 1008 834
use sg13g2_mux2_1  _066_
timestamp 1677247768
transform -1 0 35232 0 1 8316
box -48 -56 1008 834
use sg13g2_mux2_1  _067_
timestamp 1677247768
transform -1 0 10080 0 -1 9828
box -48 -56 1008 834
use sg13g2_nand2b_1  _068_
timestamp 1676567195
transform 1 0 4800 0 1 2268
box -48 -56 528 834
use sg13g2_o21ai_1  _069_
timestamp 1685175443
transform -1 0 5760 0 1 2268
box -48 -56 538 834
use sg13g2_nand3_1  _070_
timestamp 1683988354
transform 1 0 3648 0 1 2268
box -48 -56 528 834
use sg13g2_o21ai_1  _071_
timestamp 1685175443
transform 1 0 3744 0 -1 2268
box -48 -56 538 834
use sg13g2_nand3b_1  _072_
timestamp 1676573470
transform 1 0 4128 0 1 2268
box -48 -56 720 834
use sg13g2_o21ai_1  _073_
timestamp 1685175443
transform -1 0 4608 0 1 756
box -48 -56 538 834
use sg13g2_nand2_1  _074_
timestamp 1676557249
transform -1 0 5184 0 -1 2268
box -48 -56 432 834
use sg13g2_nand4_1  _075_
timestamp 1685201930
transform -1 0 4800 0 -1 2268
box -48 -56 624 834
use sg13g2_o21ai_1  _076_
timestamp 1685175443
transform 1 0 4608 0 1 756
box -48 -56 538 834
use sg13g2_nand2b_1  _077_
timestamp 1676567195
transform 1 0 5088 0 1 5292
box -48 -56 528 834
use sg13g2_mux4_1  _078_
timestamp 1677257233
transform -1 0 6432 0 -1 6804
box -48 -56 2064 834
use sg13g2_o21ai_1  _079_
timestamp 1685175443
transform 1 0 5376 0 -1 5292
box -48 -56 538 834
use sg13g2_o21ai_1  _080_
timestamp 1685175443
transform 1 0 6912 0 -1 6804
box -48 -56 538 834
use sg13g2_nand2b_1  _081_
timestamp 1676567195
transform -1 0 6624 0 1 6804
box -48 -56 528 834
use sg13g2_o21ai_1  _082_
timestamp 1685175443
transform 1 0 6432 0 -1 6804
box -48 -56 538 834
use sg13g2_inv_1  _083_
timestamp 1676382929
transform -1 0 4896 0 1 5292
box -48 -56 336 834
use sg13g2_inv_1  _084_
timestamp 1676382929
transform 1 0 3360 0 1 2268
box -48 -56 336 834
use sg13g2_mux2_1  _085_
timestamp 1677247768
transform 1 0 4128 0 -1 8316
box -48 -56 1008 834
use sg13g2_or2_1  _086_
timestamp 1684236171
transform 1 0 1536 0 1 8316
box -48 -56 528 834
use sg13g2_a21oi_1  _087_
timestamp 1683973020
transform 1 0 3552 0 1 6804
box -48 -56 528 834
use sg13g2_a221oi_1  _088_
timestamp 1685197497
transform 1 0 4416 0 -1 9828
box -48 -56 816 834
use sg13g2_nand2_1  _089_
timestamp 1676557249
transform -1 0 6528 0 -1 9828
box -48 -56 432 834
use sg13g2_nand2b_1  _090_
timestamp 1676567195
transform -1 0 4416 0 -1 9828
box -48 -56 528 834
use sg13g2_a21oi_1  _091_
timestamp 1683973020
transform 1 0 3648 0 -1 8316
box -48 -56 528 834
use sg13g2_nor2b_1  _092_
timestamp 1685181386
transform 1 0 4032 0 1 6804
box -54 -56 528 834
use sg13g2_o21ai_1  _093_
timestamp 1685175443
transform -1 0 6144 0 -1 9828
box -48 -56 538 834
use sg13g2_o21ai_1  _094_
timestamp 1685175443
transform -1 0 3936 0 -1 9828
box -48 -56 538 834
use sg13g2_o21ai_1  _095_
timestamp 1685175443
transform 1 0 5184 0 -1 9828
box -48 -56 538 834
use sg13g2_mux4_1  _096_
timestamp 1677257233
transform 1 0 5760 0 -1 8316
box -48 -56 2064 834
use sg13g2_mux4_1  _097_
timestamp 1677257233
transform 1 0 5952 0 1 8316
box -48 -56 2064 834
use sg13g2_mux2_1  _098_
timestamp 1677247768
transform -1 0 7488 0 -1 9828
box -48 -56 1008 834
use sg13g2_nand2b_1  _099_
timestamp 1676567195
transform 1 0 5376 0 1 8316
box -48 -56 528 834
use sg13g2_o21ai_1  _100_
timestamp 1685175443
transform 1 0 5280 0 -1 8316
box -48 -56 538 834
use sg13g2_mux2_1  _101_
timestamp 1677247768
transform 1 0 3936 0 1 3780
box -48 -56 1008 834
use sg13g2_or2_1  _102_
timestamp 1684236171
transform 1 0 4128 0 1 5292
box -48 -56 528 834
use sg13g2_a21oi_1  _103_
timestamp 1683973020
transform 1 0 4032 0 -1 5292
box -48 -56 528 834
use sg13g2_a221oi_1  _104_
timestamp 1685197497
transform 1 0 4032 0 -1 3780
box -48 -56 816 834
use sg13g2_nand2_1  _105_
timestamp 1676557249
transform 1 0 4992 0 -1 5292
box -48 -56 432 834
use sg13g2_nand2b_1  _106_
timestamp 1676567195
transform -1 0 5280 0 -1 3780
box -48 -56 528 834
use sg13g2_a21oi_1  _107_
timestamp 1683973020
transform 1 0 3456 0 1 3780
box -48 -56 528 834
use sg13g2_nor2b_1  _108_
timestamp 1685181386
transform 1 0 4512 0 -1 5292
box -54 -56 528 834
use sg13g2_o21ai_1  _109_
timestamp 1685175443
transform -1 0 5376 0 1 3780
box -48 -56 538 834
use sg13g2_o21ai_1  _110_
timestamp 1685175443
transform 1 0 5376 0 1 3780
box -48 -56 538 834
use sg13g2_o21ai_1  _111_
timestamp 1685175443
transform 1 0 3552 0 -1 3780
box -48 -56 538 834
use sg13g2_mux4_1  _112_
timestamp 1677257233
transform 1 0 5856 0 -1 5292
box -48 -56 2064 834
use sg13g2_mux4_1  _113_
timestamp 1677257233
transform 1 0 5568 0 1 5292
box -48 -56 2064 834
use sg13g2_mux2_1  _114_
timestamp 1677247768
transform -1 0 7584 0 -1 3780
box -48 -56 1008 834
use sg13g2_nand2b_1  _115_
timestamp 1676567195
transform 1 0 3552 0 -1 5292
box -48 -56 528 834
use sg13g2_o21ai_1  _116_
timestamp 1685175443
transform 1 0 5856 0 1 3780
box -48 -56 538 834
use sg13g2_mux4_1  _117_
timestamp 1677257233
transform 1 0 17856 0 1 5292
box -48 -56 2064 834
use sg13g2_mux4_1  _118_
timestamp 1677257233
transform 1 0 17376 0 -1 8316
box -48 -56 2064 834
use sg13g2_mux4_1  _119_
timestamp 1677257233
transform 1 0 31392 0 1 5292
box -48 -56 2064 834
use sg13g2_mux4_1  _120_
timestamp 1677257233
transform 1 0 34752 0 1 3780
box -48 -56 2064 834
use sg13g2_mux4_1  _121_
timestamp 1677257233
transform 1 0 15936 0 1 2268
box -48 -56 2064 834
use sg13g2_mux4_1  _122_
timestamp 1677257233
transform 1 0 19680 0 1 3780
box -48 -56 2064 834
use sg13g2_mux4_1  _123_
timestamp 1677257233
transform 1 0 35136 0 -1 3780
box -48 -56 2064 834
use sg13g2_mux4_1  _124_
timestamp 1677257233
transform -1 0 21600 0 1 2268
box -48 -56 2064 834
use sg13g2_mux4_1  _125_
timestamp 1677257233
transform 1 0 6720 0 1 3780
box -48 -56 2064 834
use sg13g2_mux4_1  _126_
timestamp 1677257233
transform 1 0 14400 0 -1 8316
box -48 -56 2064 834
use sg13g2_mux4_1  _127_
timestamp 1677257233
transform 1 0 14592 0 1 8316
box -48 -56 2064 834
use sg13g2_mux4_1  _128_
timestamp 1677257233
transform 1 0 18528 0 1 8316
box -48 -56 2064 834
use sg13g2_mux4_1  _129_
timestamp 1677257233
transform 1 0 31296 0 -1 6804
box -48 -56 2064 834
use sg13g2_mux4_1  _130_
timestamp 1677257233
transform 1 0 32448 0 -1 3780
box -48 -56 2064 834
use sg13g2_mux4_1  _131_
timestamp 1677257233
transform 1 0 15264 0 1 3780
box -48 -56 2064 834
use sg13g2_mux4_1  _132_
timestamp 1677257233
transform 1 0 20832 0 -1 8316
box -48 -56 2064 834
use sg13g2_mux4_1  _133_
timestamp 1677257233
transform 1 0 23808 0 -1 6804
box -48 -56 2064 834
use sg13g2_mux4_1  _134_
timestamp 1677257233
transform 1 0 28896 0 1 8316
box -48 -56 2064 834
use sg13g2_mux4_1  _135_
timestamp 1677257233
transform 1 0 23232 0 1 3780
box -48 -56 2064 834
use sg13g2_mux4_1  _136_
timestamp 1677257233
transform 1 0 28992 0 -1 5292
box -48 -56 2064 834
use sg13g2_mux4_1  _137_
timestamp 1677257233
transform 1 0 25344 0 1 2268
box -48 -56 2064 834
use sg13g2_mux4_1  _138_
timestamp 1677257233
transform 1 0 28992 0 -1 6804
box -48 -56 2064 834
use sg13g2_mux4_1  _139_
timestamp 1677257233
transform 1 0 25248 0 1 3780
box -48 -56 2064 834
use sg13g2_mux4_1  _140_
timestamp 1677257233
transform 1 0 28704 0 1 5292
box -48 -56 2064 834
use sg13g2_mux4_1  _141_
timestamp 1677257233
transform 1 0 12960 0 1 3780
box -48 -56 2064 834
use sg13g2_mux4_1  _142_
timestamp 1677257233
transform 1 0 38112 0 -1 8316
box -48 -56 2064 834
use sg13g2_mux4_1  _143_
timestamp 1677257233
transform 1 0 9600 0 1 6804
box -48 -56 2064 834
use sg13g2_mux4_1  _144_
timestamp 1677257233
transform 1 0 36096 0 -1 8316
box -48 -56 2064 834
use sg13g2_mux4_1  _145_
timestamp 1677257233
transform -1 0 16608 0 -1 6804
box -48 -56 2064 834
use sg13g2_mux4_1  _146_
timestamp 1677257233
transform 1 0 38112 0 -1 6804
box -48 -56 2064 834
use sg13g2_mux4_1  _147_
timestamp 1677257233
transform 1 0 12288 0 -1 6804
box -48 -56 2064 834
use sg13g2_dlhq_1  _148_
timestamp 1678805552
transform 1 0 6432 0 1 756
box -50 -56 1692 834
use sg13g2_dlhq_1  _149_
timestamp 1678805552
transform 1 0 7200 0 -1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _150_
timestamp 1678805552
transform 1 0 8832 0 -1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _151_
timestamp 1678805552
transform 1 0 10464 0 -1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _152_
timestamp 1678805552
transform 1 0 11328 0 1 756
box -50 -56 1692 834
use sg13g2_dlhq_1  _153_
timestamp 1678805552
transform 1 0 12096 0 -1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _154_
timestamp 1678805552
transform 1 0 13728 0 -1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _155_
timestamp 1678805552
transform 1 0 15360 0 -1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _156_
timestamp 1678805552
transform 1 0 7488 0 -1 9828
box -50 -56 1692 834
use sg13g2_dlhq_1  _157_
timestamp 1678805552
transform 1 0 33216 0 -1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _158_
timestamp 1678805552
transform 1 0 7392 0 -1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _159_
timestamp 1678805552
transform 1 0 17568 0 -1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _160_
timestamp 1678805552
transform 1 0 33312 0 -1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _161_
timestamp 1678805552
transform 1 0 34272 0 -1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _162_
timestamp 1678805552
transform 1 0 7584 0 1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _163_
timestamp 1678805552
transform 1 0 9216 0 1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _164_
timestamp 1678805552
transform 1 0 25728 0 1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _165_
timestamp 1678805552
transform 1 0 27648 0 1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _166_
timestamp 1678805552
transform 1 0 20640 0 1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _167_
timestamp 1678805552
transform 1 0 22656 0 -1 9828
box -50 -56 1692 834
use sg13g2_dlhq_1  _168_
timestamp 1678805552
transform 1 0 31104 0 -1 9828
box -50 -56 1692 834
use sg13g2_dlhq_1  _169_
timestamp 1678805552
transform 1 0 32832 0 -1 9828
box -50 -56 1692 834
use sg13g2_dlhq_1  _170_
timestamp 1678805552
transform 1 0 8736 0 1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _171_
timestamp 1678805552
transform 1 0 10848 0 -1 9828
box -50 -56 1692 834
use sg13g2_dlhq_1  _172_
timestamp 1678805552
transform 1 0 24288 0 -1 9828
box -50 -56 1692 834
use sg13g2_dlhq_1  _173_
timestamp 1678805552
transform -1 0 28512 0 -1 9828
box -50 -56 1692 834
use sg13g2_dlhq_1  _174_
timestamp 1678805552
transform 1 0 19968 0 -1 3780
box -50 -56 1692 834
use sg13g2_dlhq_1  _175_
timestamp 1678805552
transform 1 0 21600 0 1 756
box -50 -56 1692 834
use sg13g2_dlhq_1  _176_
timestamp 1678805552
transform -1 0 38016 0 -1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _177_
timestamp 1678805552
transform 1 0 37056 0 1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _178_
timestamp 1678805552
transform 1 0 8064 0 1 756
box -50 -56 1692 834
use sg13g2_dlhq_1  _179_
timestamp 1678805552
transform 1 0 9696 0 1 756
box -50 -56 1692 834
use sg13g2_dlhq_1  _180_
timestamp 1678805552
transform 1 0 25824 0 -1 3780
box -50 -56 1692 834
use sg13g2_dlhq_1  _181_
timestamp 1678805552
transform 1 0 27456 0 1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _182_
timestamp 1678805552
transform 1 0 21216 0 -1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _183_
timestamp 1678805552
transform 1 0 22848 0 -1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _184_
timestamp 1678805552
transform -1 0 38880 0 -1 3780
box -50 -56 1692 834
use sg13g2_dlhq_1  _185_
timestamp 1678805552
transform -1 0 40416 0 -1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _186_
timestamp 1678805552
transform 1 0 9024 0 1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _187_
timestamp 1678805552
transform 1 0 10944 0 1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _188_
timestamp 1678805552
transform 1 0 24000 0 -1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _189_
timestamp 1678805552
transform 1 0 26016 0 1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _190_
timestamp 1678805552
transform 1 0 19776 0 -1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _191_
timestamp 1678805552
transform 1 0 21216 0 1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _192_
timestamp 1678805552
transform 1 0 34464 0 1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _193_
timestamp 1678805552
transform 1 0 36192 0 1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _194_
timestamp 1678805552
transform 1 0 10656 0 -1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _195_
timestamp 1678805552
transform 1 0 12384 0 -1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _196_
timestamp 1678805552
transform 1 0 38880 0 1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _197_
timestamp 1678805552
transform 1 0 37152 0 -1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _198_
timestamp 1678805552
transform -1 0 16224 0 1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _199_
timestamp 1678805552
transform 1 0 12960 0 1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _200_
timestamp 1678805552
transform -1 0 39840 0 -1 9828
box -50 -56 1692 834
use sg13g2_dlhq_1  _201_
timestamp 1678805552
transform 1 0 34944 0 -1 9828
box -50 -56 1692 834
use sg13g2_dlhq_1  _202_
timestamp 1678805552
transform 1 0 9696 0 -1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _203_
timestamp 1678805552
transform 1 0 7968 0 1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _204_
timestamp 1678805552
transform -1 0 39168 0 1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _205_
timestamp 1678805552
transform 1 0 38880 0 1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _206_
timestamp 1678805552
transform 1 0 12192 0 -1 3780
box -50 -56 1692 834
use sg13g2_dlhq_1  _207_
timestamp 1678805552
transform 1 0 12960 0 1 756
box -50 -56 1692 834
use sg13g2_dlhq_1  _208_
timestamp 1678805552
transform 1 0 27552 0 1 756
box -50 -56 1692 834
use sg13g2_dlhq_1  _209_
timestamp 1678805552
transform 1 0 29472 0 -1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _210_
timestamp 1678805552
transform 1 0 23616 0 1 756
box -50 -56 1692 834
use sg13g2_dlhq_1  _211_
timestamp 1678805552
transform 1 0 25344 0 1 756
box -50 -56 1692 834
use sg13g2_dlhq_1  _212_
timestamp 1678805552
transform 1 0 29568 0 1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _213_
timestamp 1678805552
transform 1 0 27840 0 -1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _214_
timestamp 1678805552
transform 1 0 26112 0 -1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _215_
timestamp 1678805552
transform 1 0 24480 0 -1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _216_
timestamp 1678805552
transform 1 0 29280 0 -1 3780
box -50 -56 1692 834
use sg13g2_dlhq_1  _217_
timestamp 1678805552
transform 1 0 27456 0 1 3780
box -50 -56 1692 834
use sg13g2_dlhq_1  _218_
timestamp 1678805552
transform 1 0 23808 0 -1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _219_
timestamp 1678805552
transform 1 0 21984 0 1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _220_
timestamp 1678805552
transform 1 0 27936 0 -1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _221_
timestamp 1678805552
transform 1 0 29664 0 -1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _222_
timestamp 1678805552
transform 1 0 22848 0 1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _223_
timestamp 1678805552
transform 1 0 24288 0 1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _224_
timestamp 1678805552
transform 1 0 19584 0 1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _225_
timestamp 1678805552
transform 1 0 21312 0 1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _226_
timestamp 1678805552
transform 1 0 13824 0 -1 3780
box -50 -56 1692 834
use sg13g2_dlhq_1  _227_
timestamp 1678805552
transform 1 0 15456 0 -1 3780
box -50 -56 1692 834
use sg13g2_dlhq_1  _228_
timestamp 1678805552
transform 1 0 31392 0 1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _229_
timestamp 1678805552
transform 1 0 32448 0 1 3780
box -50 -56 1692 834
use sg13g2_dlhq_1  _230_
timestamp 1678805552
transform 1 0 30144 0 1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _231_
timestamp 1678805552
transform 1 0 31872 0 1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _232_
timestamp 1678805552
transform 1 0 16896 0 1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _233_
timestamp 1678805552
transform 1 0 19104 0 -1 9828
box -50 -56 1692 834
use sg13g2_dlhq_1  _234_
timestamp 1678805552
transform 1 0 12960 0 1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _235_
timestamp 1678805552
transform 1 0 14880 0 -1 9828
box -50 -56 1692 834
use sg13g2_dlhq_1  _236_
timestamp 1678805552
transform 1 0 14304 0 1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _237_
timestamp 1678805552
transform 1 0 12672 0 -1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _238_
timestamp 1678805552
transform 1 0 6432 0 1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _239_
timestamp 1678805552
transform 1 0 5184 0 -1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _240_
timestamp 1678805552
transform 1 0 18336 0 1 756
box -50 -56 1692 834
use sg13g2_dlhq_1  _241_
timestamp 1678805552
transform 1 0 17952 0 1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _242_
timestamp 1678805552
transform -1 0 36384 0 -1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _243_
timestamp 1678805552
transform 1 0 35520 0 1 756
box -50 -56 1692 834
use sg13g2_dlhq_1  _244_
timestamp 1678805552
transform 1 0 18240 0 -1 3780
box -50 -56 1692 834
use sg13g2_dlhq_1  _245_
timestamp 1678805552
transform 1 0 19968 0 1 756
box -50 -56 1692 834
use sg13g2_dlhq_1  _246_
timestamp 1678805552
transform 1 0 14304 0 1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _247_
timestamp 1678805552
transform 1 0 16224 0 1 756
box -50 -56 1692 834
use sg13g2_dlhq_1  _248_
timestamp 1678805552
transform 1 0 33600 0 1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _249_
timestamp 1678805552
transform 1 0 35424 0 1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _250_
timestamp 1678805552
transform 1 0 30528 0 1 3780
box -50 -56 1692 834
use sg13g2_dlhq_1  _251_
timestamp 1678805552
transform 1 0 31968 0 -1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _252_
timestamp 1678805552
transform 1 0 17568 0 1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _253_
timestamp 1678805552
transform 1 0 15936 0 1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _254_
timestamp 1678805552
transform 1 0 18240 0 -1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _255_
timestamp 1678805552
transform 1 0 16224 0 1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _256_
timestamp 1678805552
transform 1 0 1632 0 -1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _257_
timestamp 1678805552
transform 1 0 1632 0 1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _258_
timestamp 1678805552
transform 1 0 1536 0 1 3780
box -50 -56 1692 834
use sg13g2_dlhq_1  _259_
timestamp 1678805552
transform 1 0 1536 0 -1 3780
box -50 -56 1692 834
use sg13g2_dlhq_1  _260_
timestamp 1678805552
transform 1 0 2400 0 1 756
box -50 -56 1692 834
use sg13g2_dlhq_1  _261_
timestamp 1678805552
transform 1 0 1824 0 -1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _262_
timestamp 1678805552
transform 1 0 1728 0 1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _263_
timestamp 1678805552
transform 1 0 1824 0 -1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _264_
timestamp 1678805552
transform 1 0 2016 0 1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _265_
timestamp 1678805552
transform 1 0 1824 0 -1 9828
box -50 -56 1692 834
use sg13g2_dlhq_1  _266_
timestamp 1678805552
transform 1 0 3648 0 1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _267_
timestamp 1678805552
transform 1 0 1536 0 1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _268_
timestamp 1678805552
transform 1 0 2688 0 -1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _269_
timestamp 1678805552
transform 1 0 4512 0 1 6804
box -50 -56 1692 834
use sg13g2_dfrbpq_1  _270_
timestamp 1746535128
transform -1 0 34752 0 -1 2268
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _271_
timestamp 1746535128
transform 1 0 17088 0 -1 2268
box -48 -56 2640 834
use sg13g2_tiehi  _272_
timestamp 1680000651
transform 1 0 33792 0 1 756
box -48 -56 432 834
use sg13g2_tiehi  _273_
timestamp 1680000651
transform -1 0 18240 0 1 756
box -48 -56 432 834
use sg13g2_tielo  _274_
timestamp 1680000637
transform -1 0 19776 0 -1 8316
box -48 -56 432 834
use sg13g2_buf_1  _275_
timestamp 1676381911
transform 1 0 40800 0 1 756
box -48 -56 432 834
use sg13g2_buf_1  _276_
timestamp 1676381911
transform 1 0 39936 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _277_
timestamp 1676381911
transform 1 0 41184 0 1 756
box -48 -56 432 834
use sg13g2_buf_1  _278_
timestamp 1676381911
transform 1 0 40416 0 1 756
box -48 -56 432 834
use sg13g2_buf_1  _279_
timestamp 1676381911
transform 1 0 39552 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _280_
timestamp 1676381911
transform 1 0 41184 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _281_
timestamp 1676381911
transform 1 0 40800 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _282_
timestamp 1676381911
transform 1 0 41184 0 1 2268
box -48 -56 432 834
use sg13g2_buf_1  _283_
timestamp 1676381911
transform 1 0 40416 0 1 2268
box -48 -56 432 834
use sg13g2_buf_1  _284_
timestamp 1676381911
transform 1 0 40800 0 1 2268
box -48 -56 432 834
use sg13g2_buf_1  _285_
timestamp 1676381911
transform 1 0 40416 0 -1 3780
box -48 -56 432 834
use sg13g2_buf_1  _286_
timestamp 1676381911
transform 1 0 40800 0 -1 3780
box -48 -56 432 834
use sg13g2_buf_1  _287_
timestamp 1676381911
transform 1 0 41184 0 1 3780
box -48 -56 432 834
use sg13g2_buf_1  _288_
timestamp 1676381911
transform 1 0 40416 0 1 3780
box -48 -56 432 834
use sg13g2_buf_1  _289_
timestamp 1676381911
transform 1 0 40800 0 1 3780
box -48 -56 432 834
use sg13g2_buf_1  _290_
timestamp 1676381911
transform 1 0 41184 0 -1 5292
box -48 -56 432 834
use sg13g2_buf_1  _291_
timestamp 1676381911
transform 1 0 40800 0 -1 5292
box -48 -56 432 834
use sg13g2_buf_1  _292_
timestamp 1676381911
transform 1 0 41184 0 1 5292
box -48 -56 432 834
use sg13g2_buf_1  _293_
timestamp 1676381911
transform 1 0 40800 0 1 5292
box -48 -56 432 834
use sg13g2_buf_1  _294_
timestamp 1676381911
transform 1 0 40800 0 -1 6804
box -48 -56 432 834
use sg13g2_buf_1  _295_
timestamp 1676381911
transform 1 0 41184 0 -1 6804
box -48 -56 432 834
use sg13g2_buf_1  _296_
timestamp 1676381911
transform 1 0 40800 0 1 6804
box -48 -56 432 834
use sg13g2_buf_1  _297_
timestamp 1676381911
transform 1 0 41184 0 1 6804
box -48 -56 432 834
use sg13g2_buf_1  _298_
timestamp 1676381911
transform 1 0 40800 0 -1 8316
box -48 -56 432 834
use sg13g2_buf_1  _299_
timestamp 1676381911
transform 1 0 40416 0 -1 8316
box -48 -56 432 834
use sg13g2_buf_1  _300_
timestamp 1676381911
transform 1 0 40800 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  _301_
timestamp 1676381911
transform 1 0 40416 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  _302_
timestamp 1676381911
transform 1 0 41184 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  _303_
timestamp 1676381911
transform 1 0 40800 0 -1 9828
box -48 -56 432 834
use sg13g2_buf_1  _304_
timestamp 1676381911
transform 1 0 40032 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  _305_
timestamp 1676381911
transform 1 0 41184 0 -1 8316
box -48 -56 432 834
use sg13g2_buf_1  _306_
timestamp 1676381911
transform 1 0 41184 0 -1 9828
box -48 -56 432 834
use sg13g2_buf_1  _307_
timestamp 1676381911
transform 1 0 29568 0 -1 9828
box -48 -56 432 834
use sg13g2_buf_1  _308_
timestamp 1676381911
transform -1 0 30336 0 -1 9828
box -48 -56 432 834
use sg13g2_buf_1  _309_
timestamp 1676381911
transform -1 0 30720 0 -1 9828
box -48 -56 432 834
use sg13g2_buf_1  _310_
timestamp 1676381911
transform -1 0 31104 0 -1 9828
box -48 -56 432 834
use sg13g2_buf_1  _311_
timestamp 1676381911
transform -1 0 31488 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _312_
timestamp 1676381911
transform -1 0 31872 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _313_
timestamp 1676381911
transform -1 0 31488 0 -1 3780
box -48 -56 432 834
use sg13g2_buf_1  _314_
timestamp 1676381911
transform -1 0 32640 0 1 756
box -48 -56 432 834
use sg13g2_buf_1  _315_
timestamp 1676381911
transform -1 0 31872 0 -1 3780
box -48 -56 432 834
use sg13g2_buf_1  _316_
timestamp 1676381911
transform -1 0 33024 0 1 756
box -48 -56 432 834
use sg13g2_buf_1  _317_
timestamp 1676381911
transform -1 0 33408 0 1 756
box -48 -56 432 834
use sg13g2_buf_1  _318_
timestamp 1676381911
transform -1 0 33792 0 1 756
box -48 -56 432 834
use sg13g2_buf_1  _319_
timestamp 1676381911
transform -1 0 34560 0 1 756
box -48 -56 432 834
use sg13g2_buf_1  _320_
timestamp 1676381911
transform -1 0 34944 0 1 756
box -48 -56 432 834
use sg13g2_buf_1  _321_
timestamp 1676381911
transform -1 0 35328 0 1 756
box -48 -56 432 834
use sg13g2_buf_1  _322_
timestamp 1676381911
transform -1 0 37536 0 1 756
box -48 -56 432 834
use sg13g2_buf_1  _323_
timestamp 1676381911
transform -1 0 37920 0 1 756
box -48 -56 432 834
use sg13g2_buf_1  _324_
timestamp 1676381911
transform -1 0 38496 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _325_
timestamp 1676381911
transform -1 0 39552 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _326_
timestamp 1676381911
transform -1 0 40704 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _327_
timestamp 1676381911
transform 1 0 8352 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  _328_
timestamp 1676381911
transform -1 0 10464 0 -1 9828
box -48 -56 432 834
use sg13g2_buf_1  _329_
timestamp 1676381911
transform 1 0 9312 0 -1 8316
box -48 -56 432 834
use sg13g2_buf_1  _330_
timestamp 1676381911
transform -1 0 10656 0 -1 6804
box -48 -56 432 834
use sg13g2_buf_1  _331_
timestamp 1676381911
transform -1 0 36000 0 -1 6804
box -48 -56 432 834
use sg13g2_buf_1  _332_
timestamp 1676381911
transform -1 0 11232 0 1 5292
box -48 -56 432 834
use sg13g2_buf_1  _333_
timestamp 1676381911
transform -1 0 12000 0 1 6804
box -48 -56 432 834
use sg13g2_buf_1  _334_
timestamp 1676381911
transform 1 0 10464 0 -1 9828
box -48 -56 432 834
use sg13g2_buf_1  _335_
timestamp 1676381911
transform -1 0 33984 0 1 6804
box -48 -56 432 834
use sg13g2_buf_1  _336_
timestamp 1676381911
transform -1 0 11808 0 -1 8316
box -48 -56 432 834
use sg13g2_buf_1  _337_
timestamp 1676381911
transform -1 0 12192 0 -1 8316
box -48 -56 432 834
use sg13g2_buf_1  _338_
timestamp 1676381911
transform -1 0 12384 0 -1 5292
box -48 -56 432 834
use sg13g2_buf_1  _339_
timestamp 1676381911
transform -1 0 37920 0 -1 6804
box -48 -56 432 834
use sg13g2_buf_1  _340_
timestamp 1676381911
transform 1 0 11616 0 -1 5292
box -48 -56 432 834
use sg13g2_buf_1  _341_
timestamp 1676381911
transform -1 0 28608 0 1 5292
box -48 -56 432 834
use sg13g2_buf_1  _342_
timestamp 1676381911
transform -1 0 13152 0 1 2268
box -48 -56 432 834
use sg13g2_buf_1  _343_
timestamp 1676381911
transform -1 0 40800 0 -1 5292
box -48 -56 432 834
use sg13g2_buf_1  _344_
timestamp 1676381911
transform 1 0 12576 0 1 5292
box -48 -56 432 834
use sg13g2_buf_1  _345_
timestamp 1676381911
transform -1 0 28224 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  _346_
timestamp 1676381911
transform -1 0 23232 0 -1 8316
box -48 -56 432 834
use sg13g2_buf_1  _347_
timestamp 1676381911
transform -1 0 37344 0 -1 9828
box -48 -56 432 834
use sg13g2_buf_1  _348_
timestamp 1676381911
transform -1 0 14016 0 1 6804
box -48 -56 432 834
use sg13g2_buf_1  _349_
timestamp 1676381911
transform -1 0 40512 0 -1 6804
box -48 -56 432 834
use sg13g2_buf_1  _350_
timestamp 1676381911
transform -1 0 14496 0 -1 9828
box -48 -56 432 834
use sg13g2_buf_1  _351_
timestamp 1676381911
transform -1 0 37920 0 -1 9828
box -48 -56 432 834
use sg13g2_buf_1  _352_
timestamp 1676381911
transform 1 0 12672 0 1 6804
box -48 -56 432 834
use sg13g2_buf_1  _353_
timestamp 1676381911
transform -1 0 40032 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  _354_
timestamp 1676381911
transform -1 0 14976 0 -1 5292
box -48 -56 432 834
use sg13g2_buf_1  _355_
timestamp 1676381911
transform -1 0 31680 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  _356_
timestamp 1676381911
transform -1 0 25824 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  _357_
timestamp 1676381911
transform -1 0 32064 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  _358_
timestamp 1676381911
transform -1 0 29088 0 -1 3780
box -48 -56 432 834
use sg13g2_buf_1  _359_
timestamp 1676381911
transform -1 0 31296 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  _360_
timestamp 1676381911
transform -1 0 24864 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  _361_
timestamp 1676381911
transform -1 0 31680 0 -1 8316
box -48 -56 432 834
use sg13g2_buf_1  _362_
timestamp 1676381911
transform -1 0 25344 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  _363_
timestamp 1676381911
transform -1 0 22560 0 -1 9828
box -48 -56 432 834
use sg13g2_buf_1  _364_
timestamp 1676381911
transform -1 0 17088 0 -1 5292
box -48 -56 432 834
use sg13g2_buf_1  _365_
timestamp 1676381911
transform -1 0 34464 0 1 3780
box -48 -56 432 834
use sg13g2_buf_1  _366_
timestamp 1676381911
transform -1 0 32928 0 -1 8316
box -48 -56 432 834
use sg13g2_buf_1  _367_
timestamp 1676381911
transform -1 0 20352 0 -1 8316
box -48 -56 432 834
use sg13g2_buf_1  _368_
timestamp 1676381911
transform 1 0 16800 0 -1 9828
box -48 -56 432 834
use sg13g2_buf_1  _369_
timestamp 1676381911
transform 1 0 16800 0 -1 8316
box -48 -56 432 834
use sg13g2_buf_1  _370_
timestamp 1676381911
transform 1 0 17088 0 -1 5292
box -48 -56 432 834
use sg13g2_buf_1  _371_
timestamp 1676381911
transform -1 0 18240 0 -1 3780
box -48 -56 432 834
use sg13g2_buf_1  _372_
timestamp 1676381911
transform -1 0 36960 0 -1 5292
box -48 -56 432 834
use sg13g2_buf_1  _373_
timestamp 1676381911
transform -1 0 21216 0 -1 5292
box -48 -56 432 834
use sg13g2_buf_1  _374_
timestamp 1676381911
transform 1 0 17472 0 -1 3780
box -48 -56 432 834
use sg13g2_buf_1  _375_
timestamp 1676381911
transform -1 0 37152 0 1 3780
box -48 -56 432 834
use sg13g2_buf_1  _376_
timestamp 1676381911
transform -1 0 32544 0 -1 8316
box -48 -56 432 834
use sg13g2_buf_1  _377_
timestamp 1676381911
transform 1 0 18720 0 -1 9828
box -48 -56 432 834
use sg13g2_buf_1  _378_
timestamp 1676381911
transform -1 0 19776 0 -1 6804
box -48 -56 432 834
use sg13g2_buf_1  _379_
timestamp 1676381911
transform 1 0 29376 0 1 756
box -48 -56 432 834
use sg13g2_buf_8  clkbuf_0_UserCLK_regs
timestamp 1676451365
transform 1 0 27456 0 -1 3780
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_0_UserCLK
timestamp 1676451365
transform 1 0 31008 0 1 756
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_1_0__f_UserCLK
timestamp 1676451365
transform -1 0 30336 0 1 3780
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_1_0__f_UserCLK_regs
timestamp 1676451365
transform -1 0 24864 0 1 2268
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_1_1__f_UserCLK_regs
timestamp 1676451365
transform 1 0 29760 0 1 756
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_regs_0_UserCLK
timestamp 1676451365
transform 1 0 24576 0 -1 3780
box -48 -56 1296 834
use sg13g2_decap_8  FILLER_0_0
timestamp 1679581782
transform 1 0 1152 0 1 756
box -48 -56 720 834
use sg13g2_decap_4  FILLER_0_7
timestamp 1679577901
transform 1 0 1824 0 1 756
box -48 -56 432 834
use sg13g2_fill_2  FILLER_0_11
timestamp 1677580104
transform 1 0 2208 0 1 756
box -48 -56 240 834
use sg13g2_fill_1  FILLER_0_30
timestamp 1677579658
transform 1 0 4032 0 1 756
box -48 -56 144 834
use sg13g2_decap_8  FILLER_0_41
timestamp 1679581782
transform 1 0 5088 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_48
timestamp 1679581782
transform 1 0 5760 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_140
timestamp 1679581782
transform 1 0 14592 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_147
timestamp 1679581782
transform 1 0 15264 0 1 756
box -48 -56 720 834
use sg13g2_fill_2  FILLER_0_154
timestamp 1677580104
transform 1 0 15936 0 1 756
box -48 -56 240 834
use sg13g2_fill_1  FILLER_0_156
timestamp 1677579658
transform 1 0 16128 0 1 756
box -48 -56 144 834
use sg13g2_fill_1  FILLER_0_178
timestamp 1677579658
transform 1 0 18240 0 1 756
box -48 -56 144 834
use sg13g2_decap_4  FILLER_0_230
timestamp 1679577901
transform 1 0 23232 0 1 756
box -48 -56 432 834
use sg13g2_fill_1  FILLER_0_251
timestamp 1677579658
transform 1 0 25248 0 1 756
box -48 -56 144 834
use sg13g2_decap_4  FILLER_0_269
timestamp 1679577901
transform 1 0 26976 0 1 756
box -48 -56 432 834
use sg13g2_fill_2  FILLER_0_273
timestamp 1677580104
transform 1 0 27360 0 1 756
box -48 -56 240 834
use sg13g2_fill_2  FILLER_0_292
timestamp 1677580104
transform 1 0 29184 0 1 756
box -48 -56 240 834
use sg13g2_fill_2  FILLER_0_356
timestamp 1677580104
transform 1 0 35328 0 1 756
box -48 -56 240 834
use sg13g2_decap_8  FILLER_0_383
timestamp 1679581782
transform 1 0 37920 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_390
timestamp 1679581782
transform 1 0 38592 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_397
timestamp 1679581782
transform 1 0 39264 0 1 756
box -48 -56 720 834
use sg13g2_decap_4  FILLER_0_404
timestamp 1679577901
transform 1 0 39936 0 1 756
box -48 -56 432 834
use sg13g2_fill_1  FILLER_0_408
timestamp 1677579658
transform 1 0 40320 0 1 756
box -48 -56 144 834
use sg13g2_fill_2  FILLER_0_421
timestamp 1677580104
transform 1 0 41568 0 1 756
box -48 -56 240 834
use sg13g2_fill_1  FILLER_0_423
timestamp 1677579658
transform 1 0 41760 0 1 756
box -48 -56 144 834
use sg13g2_decap_8  FILLER_1_0
timestamp 1679581782
transform 1 0 1152 0 -1 2268
box -48 -56 720 834
use sg13g2_fill_2  FILLER_1_24
timestamp 1677580104
transform 1 0 3456 0 -1 2268
box -48 -56 240 834
use sg13g2_fill_1  FILLER_1_26
timestamp 1677579658
transform 1 0 3648 0 -1 2268
box -48 -56 144 834
use sg13g2_decap_4  FILLER_1_59
timestamp 1679577901
transform 1 0 6816 0 -1 2268
box -48 -56 432 834
use sg13g2_fill_1  FILLER_1_165
timestamp 1677579658
transform 1 0 16992 0 -1 2268
box -48 -56 144 834
use sg13g2_decap_8  FILLER_1_193
timestamp 1679581782
transform 1 0 19680 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_200
timestamp 1679581782
transform 1 0 20352 0 -1 2268
box -48 -56 720 834
use sg13g2_fill_2  FILLER_1_207
timestamp 1677580104
transform 1 0 21024 0 -1 2268
box -48 -56 240 834
use sg13g2_fill_1  FILLER_1_277
timestamp 1677579658
transform 1 0 27744 0 -1 2268
box -48 -56 144 834
use sg13g2_fill_2  FILLER_1_320
timestamp 1677580104
transform 1 0 31872 0 -1 2268
box -48 -56 240 834
use sg13g2_fill_1  FILLER_1_322
timestamp 1677579658
transform 1 0 32064 0 -1 2268
box -48 -56 144 834
use sg13g2_fill_1  FILLER_1_384
timestamp 1677579658
transform 1 0 38016 0 -1 2268
box -48 -56 144 834
use sg13g2_decap_8  FILLER_1_389
timestamp 1679581782
transform 1 0 38496 0 -1 2268
box -48 -56 720 834
use sg13g2_fill_1  FILLER_1_412
timestamp 1677579658
transform 1 0 40704 0 -1 2268
box -48 -56 144 834
use sg13g2_fill_2  FILLER_1_421
timestamp 1677580104
transform 1 0 41568 0 -1 2268
box -48 -56 240 834
use sg13g2_fill_1  FILLER_1_423
timestamp 1677579658
transform 1 0 41760 0 -1 2268
box -48 -56 144 834
use sg13g2_decap_4  FILLER_2_0
timestamp 1679577901
transform 1 0 1152 0 1 2268
box -48 -56 432 834
use sg13g2_fill_2  FILLER_2_4
timestamp 1677580104
transform 1 0 1536 0 1 2268
box -48 -56 240 834
use sg13g2_decap_8  FILLER_2_48
timestamp 1679581782
transform 1 0 5760 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_72
timestamp 1679581782
transform 1 0 8064 0 1 2268
box -48 -56 720 834
use sg13g2_fill_2  FILLER_2_79
timestamp 1677580104
transform 1 0 8736 0 1 2268
box -48 -56 240 834
use sg13g2_fill_1  FILLER_2_81
timestamp 1677579658
transform 1 0 8928 0 1 2268
box -48 -56 144 834
use sg13g2_fill_2  FILLER_2_99
timestamp 1677580104
transform 1 0 10656 0 1 2268
box -48 -56 240 834
use sg13g2_fill_1  FILLER_2_101
timestamp 1677579658
transform 1 0 10848 0 1 2268
box -48 -56 144 834
use sg13g2_fill_2  FILLER_2_119
timestamp 1677580104
transform 1 0 12576 0 1 2268
box -48 -56 240 834
use sg13g2_decap_8  FILLER_2_125
timestamp 1679581782
transform 1 0 13152 0 1 2268
box -48 -56 720 834
use sg13g2_decap_4  FILLER_2_132
timestamp 1679577901
transform 1 0 13824 0 1 2268
box -48 -56 432 834
use sg13g2_fill_1  FILLER_2_136
timestamp 1677579658
transform 1 0 14208 0 1 2268
box -48 -56 144 834
use sg13g2_decap_4  FILLER_2_213
timestamp 1679577901
transform 1 0 21600 0 1 2268
box -48 -56 432 834
use sg13g2_decap_4  FILLER_2_247
timestamp 1679577901
transform 1 0 24864 0 1 2268
box -48 -56 432 834
use sg13g2_fill_1  FILLER_2_251
timestamp 1677579658
transform 1 0 25248 0 1 2268
box -48 -56 144 834
use sg13g2_fill_1  FILLER_2_273
timestamp 1677579658
transform 1 0 27360 0 1 2268
box -48 -56 144 834
use sg13g2_decap_4  FILLER_2_291
timestamp 1679577901
transform 1 0 29088 0 1 2268
box -48 -56 432 834
use sg13g2_fill_1  FILLER_2_295
timestamp 1677579658
transform 1 0 29472 0 1 2268
box -48 -56 144 834
use sg13g2_fill_2  FILLER_2_313
timestamp 1677580104
transform 1 0 31200 0 1 2268
box -48 -56 240 834
use sg13g2_decap_4  FILLER_2_332
timestamp 1679577901
transform 1 0 33024 0 1 2268
box -48 -56 432 834
use sg13g2_fill_2  FILLER_2_336
timestamp 1677580104
transform 1 0 33408 0 1 2268
box -48 -56 240 834
use sg13g2_fill_2  FILLER_2_355
timestamp 1677580104
transform 1 0 35232 0 1 2268
box -48 -56 240 834
use sg13g2_decap_8  FILLER_2_391
timestamp 1679581782
transform 1 0 38688 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_398
timestamp 1679581782
transform 1 0 39360 0 1 2268
box -48 -56 720 834
use sg13g2_decap_4  FILLER_2_405
timestamp 1679577901
transform 1 0 40032 0 1 2268
box -48 -56 432 834
use sg13g2_fill_2  FILLER_2_421
timestamp 1677580104
transform 1 0 41568 0 1 2268
box -48 -56 240 834
use sg13g2_fill_1  FILLER_2_423
timestamp 1677579658
transform 1 0 41760 0 1 2268
box -48 -56 144 834
use sg13g2_decap_4  FILLER_3_0
timestamp 1679577901
transform 1 0 1152 0 -1 3780
box -48 -56 432 834
use sg13g2_decap_4  FILLER_3_21
timestamp 1679577901
transform 1 0 3168 0 -1 3780
box -48 -56 432 834
use sg13g2_decap_8  FILLER_3_43
timestamp 1679581782
transform 1 0 5280 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_50
timestamp 1679581782
transform 1 0 5952 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_67
timestamp 1679581782
transform 1 0 7584 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_74
timestamp 1679581782
transform 1 0 8256 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_81
timestamp 1679581782
transform 1 0 8928 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_4  FILLER_3_109
timestamp 1679577901
transform 1 0 11616 0 -1 3780
box -48 -56 432 834
use sg13g2_fill_2  FILLER_3_113
timestamp 1677580104
transform 1 0 12000 0 -1 3780
box -48 -56 240 834
use sg13g2_decap_4  FILLER_3_166
timestamp 1679577901
transform 1 0 17088 0 -1 3780
box -48 -56 432 834
use sg13g2_fill_1  FILLER_3_195
timestamp 1677579658
transform 1 0 19872 0 -1 3780
box -48 -56 144 834
use sg13g2_decap_8  FILLER_3_213
timestamp 1679581782
transform 1 0 21600 0 -1 3780
box -48 -56 720 834
use sg13g2_fill_2  FILLER_3_220
timestamp 1677580104
transform 1 0 22272 0 -1 3780
box -48 -56 240 834
use sg13g2_fill_1  FILLER_3_222
timestamp 1677579658
transform 1 0 22464 0 -1 3780
box -48 -56 144 834
use sg13g2_fill_2  FILLER_3_291
timestamp 1677580104
transform 1 0 29088 0 -1 3780
box -48 -56 240 834
use sg13g2_fill_2  FILLER_3_310
timestamp 1677580104
transform 1 0 30912 0 -1 3780
box -48 -56 240 834
use sg13g2_decap_4  FILLER_3_320
timestamp 1679577901
transform 1 0 31872 0 -1 3780
box -48 -56 432 834
use sg13g2_fill_2  FILLER_3_324
timestamp 1677580104
transform 1 0 32256 0 -1 3780
box -48 -56 240 834
use sg13g2_decap_8  FILLER_3_347
timestamp 1679581782
transform 1 0 34464 0 -1 3780
box -48 -56 720 834
use sg13g2_fill_1  FILLER_3_375
timestamp 1677579658
transform 1 0 37152 0 -1 3780
box -48 -56 144 834
use sg13g2_decap_8  FILLER_3_393
timestamp 1679581782
transform 1 0 38880 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_400
timestamp 1679581782
transform 1 0 39552 0 -1 3780
box -48 -56 720 834
use sg13g2_fill_2  FILLER_3_407
timestamp 1677580104
transform 1 0 40224 0 -1 3780
box -48 -56 240 834
use sg13g2_decap_8  FILLER_3_417
timestamp 1679581782
transform 1 0 41184 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_4  FILLER_4_0
timestamp 1679577901
transform 1 0 1152 0 1 3780
box -48 -56 432 834
use sg13g2_fill_2  FILLER_4_21
timestamp 1677580104
transform 1 0 3168 0 1 3780
box -48 -56 240 834
use sg13g2_fill_1  FILLER_4_23
timestamp 1677579658
transform 1 0 3360 0 1 3780
box -48 -56 144 834
use sg13g2_decap_4  FILLER_4_54
timestamp 1679577901
transform 1 0 6336 0 1 3780
box -48 -56 432 834
use sg13g2_decap_8  FILLER_4_79
timestamp 1679581782
transform 1 0 8736 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_86
timestamp 1679581782
transform 1 0 9408 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_93
timestamp 1679581782
transform 1 0 10080 0 1 3780
box -48 -56 720 834
use sg13g2_fill_2  FILLER_4_121
timestamp 1677580104
transform 1 0 12768 0 1 3780
box -48 -56 240 834
use sg13g2_fill_2  FILLER_4_144
timestamp 1677580104
transform 1 0 14976 0 1 3780
box -48 -56 240 834
use sg13g2_fill_1  FILLER_4_146
timestamp 1677579658
transform 1 0 15168 0 1 3780
box -48 -56 144 834
use sg13g2_decap_8  FILLER_4_168
timestamp 1679581782
transform 1 0 17280 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_175
timestamp 1679581782
transform 1 0 17952 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_182
timestamp 1679581782
transform 1 0 18624 0 1 3780
box -48 -56 720 834
use sg13g2_decap_4  FILLER_4_189
timestamp 1679577901
transform 1 0 19296 0 1 3780
box -48 -56 432 834
use sg13g2_decap_8  FILLER_4_214
timestamp 1679581782
transform 1 0 21696 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_221
timestamp 1679581782
transform 1 0 22368 0 1 3780
box -48 -56 720 834
use sg13g2_fill_2  FILLER_4_228
timestamp 1677580104
transform 1 0 23040 0 1 3780
box -48 -56 240 834
use sg13g2_fill_2  FILLER_4_272
timestamp 1677580104
transform 1 0 27264 0 1 3780
box -48 -56 240 834
use sg13g2_fill_2  FILLER_4_304
timestamp 1677580104
transform 1 0 30336 0 1 3780
box -48 -56 240 834
use sg13g2_fill_2  FILLER_4_323
timestamp 1677580104
transform 1 0 32160 0 1 3780
box -48 -56 240 834
use sg13g2_fill_1  FILLER_4_325
timestamp 1677579658
transform 1 0 32352 0 1 3780
box -48 -56 144 834
use sg13g2_fill_2  FILLER_4_347
timestamp 1677580104
transform 1 0 34464 0 1 3780
box -48 -56 240 834
use sg13g2_fill_1  FILLER_4_349
timestamp 1677579658
transform 1 0 34656 0 1 3780
box -48 -56 144 834
use sg13g2_decap_4  FILLER_4_375
timestamp 1679577901
transform 1 0 37152 0 1 3780
box -48 -56 432 834
use sg13g2_fill_2  FILLER_4_379
timestamp 1677580104
transform 1 0 37536 0 1 3780
box -48 -56 240 834
use sg13g2_decap_8  FILLER_4_402
timestamp 1679581782
transform 1 0 39744 0 1 3780
box -48 -56 720 834
use sg13g2_fill_2  FILLER_4_421
timestamp 1677580104
transform 1 0 41568 0 1 3780
box -48 -56 240 834
use sg13g2_fill_1  FILLER_4_423
timestamp 1677579658
transform 1 0 41760 0 1 3780
box -48 -56 144 834
use sg13g2_decap_4  FILLER_5_0
timestamp 1679577901
transform 1 0 1152 0 -1 5292
box -48 -56 432 834
use sg13g2_fill_1  FILLER_5_4
timestamp 1677579658
transform 1 0 1536 0 -1 5292
box -48 -56 144 834
use sg13g2_fill_2  FILLER_5_22
timestamp 1677580104
transform 1 0 3264 0 -1 5292
box -48 -56 240 834
use sg13g2_fill_1  FILLER_5_24
timestamp 1677579658
transform 1 0 3456 0 -1 5292
box -48 -56 144 834
use sg13g2_decap_8  FILLER_5_70
timestamp 1679581782
transform 1 0 7872 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_77
timestamp 1679581782
transform 1 0 8544 0 -1 5292
box -48 -56 720 834
use sg13g2_fill_1  FILLER_5_84
timestamp 1677579658
transform 1 0 9216 0 -1 5292
box -48 -56 144 834
use sg13g2_fill_2  FILLER_5_106
timestamp 1677580104
transform 1 0 11328 0 -1 5292
box -48 -56 240 834
use sg13g2_fill_1  FILLER_5_108
timestamp 1677579658
transform 1 0 11520 0 -1 5292
box -48 -56 144 834
use sg13g2_decap_4  FILLER_5_134
timestamp 1679577901
transform 1 0 14016 0 -1 5292
box -48 -56 432 834
use sg13g2_fill_2  FILLER_5_138
timestamp 1677580104
transform 1 0 14400 0 -1 5292
box -48 -56 240 834
use sg13g2_decap_8  FILLER_5_144
timestamp 1679581782
transform 1 0 14976 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_151
timestamp 1679581782
transform 1 0 15648 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_4  FILLER_5_158
timestamp 1679577901
transform 1 0 16320 0 -1 5292
box -48 -56 432 834
use sg13g2_decap_8  FILLER_5_170
timestamp 1679581782
transform 1 0 17472 0 -1 5292
box -48 -56 720 834
use sg13g2_fill_1  FILLER_5_177
timestamp 1677579658
transform 1 0 18144 0 -1 5292
box -48 -56 144 834
use sg13g2_decap_8  FILLER_5_195
timestamp 1679581782
transform 1 0 19872 0 -1 5292
box -48 -56 720 834
use sg13g2_fill_2  FILLER_5_202
timestamp 1677580104
transform 1 0 20544 0 -1 5292
box -48 -56 240 834
use sg13g2_fill_1  FILLER_5_204
timestamp 1677579658
transform 1 0 20736 0 -1 5292
box -48 -56 144 834
use sg13g2_decap_4  FILLER_5_230
timestamp 1679577901
transform 1 0 23232 0 -1 5292
box -48 -56 432 834
use sg13g2_fill_2  FILLER_5_234
timestamp 1677580104
transform 1 0 23616 0 -1 5292
box -48 -56 240 834
use sg13g2_decap_8  FILLER_5_253
timestamp 1679581782
transform 1 0 25440 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_260
timestamp 1679581782
transform 1 0 26112 0 -1 5292
box -48 -56 720 834
use sg13g2_fill_2  FILLER_5_267
timestamp 1677580104
transform 1 0 26784 0 -1 5292
box -48 -56 240 834
use sg13g2_decap_8  FILLER_5_311
timestamp 1679581782
transform 1 0 31008 0 -1 5292
box -48 -56 720 834
use sg13g2_fill_2  FILLER_5_318
timestamp 1677580104
transform 1 0 31680 0 -1 5292
box -48 -56 240 834
use sg13g2_fill_1  FILLER_5_320
timestamp 1677579658
transform 1 0 31872 0 -1 5292
box -48 -56 144 834
use sg13g2_decap_8  FILLER_5_338
timestamp 1679581782
transform 1 0 33600 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_362
timestamp 1679581782
transform 1 0 35904 0 -1 5292
box -48 -56 720 834
use sg13g2_fill_2  FILLER_5_373
timestamp 1677580104
transform 1 0 36960 0 -1 5292
box -48 -56 240 834
use sg13g2_fill_2  FILLER_5_421
timestamp 1677580104
transform 1 0 41568 0 -1 5292
box -48 -56 240 834
use sg13g2_fill_1  FILLER_5_423
timestamp 1677579658
transform 1 0 41760 0 -1 5292
box -48 -56 144 834
use sg13g2_decap_4  FILLER_6_0
timestamp 1679577901
transform 1 0 1152 0 1 5292
box -48 -56 432 834
use sg13g2_decap_8  FILLER_6_21
timestamp 1679581782
transform 1 0 3168 0 1 5292
box -48 -56 720 834
use sg13g2_fill_2  FILLER_6_28
timestamp 1677580104
transform 1 0 3840 0 1 5292
box -48 -56 240 834
use sg13g2_fill_1  FILLER_6_30
timestamp 1677579658
transform 1 0 4032 0 1 5292
box -48 -56 144 834
use sg13g2_fill_2  FILLER_6_39
timestamp 1677580104
transform 1 0 4896 0 1 5292
box -48 -56 240 834
use sg13g2_decap_8  FILLER_6_105
timestamp 1679581782
transform 1 0 11232 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_112
timestamp 1679581782
transform 1 0 11904 0 1 5292
box -48 -56 720 834
use sg13g2_decap_4  FILLER_6_205
timestamp 1679577901
transform 1 0 20832 0 1 5292
box -48 -56 432 834
use sg13g2_decap_8  FILLER_6_243
timestamp 1679581782
transform 1 0 24480 0 1 5292
box -48 -56 720 834
use sg13g2_decap_4  FILLER_6_250
timestamp 1679577901
transform 1 0 25152 0 1 5292
box -48 -56 432 834
use sg13g2_fill_2  FILLER_6_254
timestamp 1677580104
transform 1 0 25536 0 1 5292
box -48 -56 240 834
use sg13g2_decap_8  FILLER_6_273
timestamp 1679581782
transform 1 0 27360 0 1 5292
box -48 -56 720 834
use sg13g2_fill_2  FILLER_6_280
timestamp 1677580104
transform 1 0 28032 0 1 5292
box -48 -56 240 834
use sg13g2_fill_1  FILLER_6_286
timestamp 1677579658
transform 1 0 28608 0 1 5292
box -48 -56 144 834
use sg13g2_decap_8  FILLER_6_308
timestamp 1679581782
transform 1 0 30720 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_336
timestamp 1679581782
transform 1 0 33408 0 1 5292
box -48 -56 720 834
use sg13g2_fill_1  FILLER_6_343
timestamp 1677579658
transform 1 0 34080 0 1 5292
box -48 -56 144 834
use sg13g2_decap_8  FILLER_6_386
timestamp 1679581782
transform 1 0 38208 0 1 5292
box -48 -56 720 834
use sg13g2_fill_2  FILLER_6_410
timestamp 1677580104
transform 1 0 40512 0 1 5292
box -48 -56 240 834
use sg13g2_fill_1  FILLER_6_412
timestamp 1677579658
transform 1 0 40704 0 1 5292
box -48 -56 144 834
use sg13g2_fill_2  FILLER_6_421
timestamp 1677580104
transform 1 0 41568 0 1 5292
box -48 -56 240 834
use sg13g2_fill_1  FILLER_6_423
timestamp 1677579658
transform 1 0 41760 0 1 5292
box -48 -56 144 834
use sg13g2_decap_8  FILLER_7_0
timestamp 1679581782
transform 1 0 1152 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_7
timestamp 1679581782
transform 1 0 1824 0 -1 6804
box -48 -56 720 834
use sg13g2_fill_2  FILLER_7_14
timestamp 1677580104
transform 1 0 2496 0 -1 6804
box -48 -56 240 834
use sg13g2_fill_1  FILLER_7_33
timestamp 1677579658
transform 1 0 4320 0 -1 6804
box -48 -56 144 834
use sg13g2_fill_2  FILLER_7_92
timestamp 1677580104
transform 1 0 9984 0 -1 6804
box -48 -56 240 834
use sg13g2_fill_1  FILLER_7_94
timestamp 1677579658
transform 1 0 10176 0 -1 6804
box -48 -56 144 834
use sg13g2_fill_2  FILLER_7_137
timestamp 1677580104
transform 1 0 14304 0 -1 6804
box -48 -56 240 834
use sg13g2_fill_1  FILLER_7_139
timestamp 1677579658
transform 1 0 14496 0 -1 6804
box -48 -56 144 834
use sg13g2_decap_8  FILLER_7_161
timestamp 1679581782
transform 1 0 16608 0 -1 6804
box -48 -56 720 834
use sg13g2_fill_2  FILLER_7_168
timestamp 1677580104
transform 1 0 17280 0 -1 6804
box -48 -56 240 834
use sg13g2_fill_1  FILLER_7_170
timestamp 1677579658
transform 1 0 17472 0 -1 6804
box -48 -56 144 834
use sg13g2_fill_2  FILLER_7_188
timestamp 1677580104
transform 1 0 19200 0 -1 6804
box -48 -56 240 834
use sg13g2_decap_4  FILLER_7_232
timestamp 1679577901
transform 1 0 23424 0 -1 6804
box -48 -56 432 834
use sg13g2_decap_8  FILLER_7_257
timestamp 1679581782
transform 1 0 25824 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_4  FILLER_7_264
timestamp 1679577901
transform 1 0 26496 0 -1 6804
box -48 -56 432 834
use sg13g2_fill_1  FILLER_7_268
timestamp 1677579658
transform 1 0 26880 0 -1 6804
box -48 -56 144 834
use sg13g2_fill_2  FILLER_7_311
timestamp 1677580104
transform 1 0 31008 0 -1 6804
box -48 -56 240 834
use sg13g2_fill_1  FILLER_7_313
timestamp 1677579658
transform 1 0 31200 0 -1 6804
box -48 -56 144 834
use sg13g2_decap_8  FILLER_7_352
timestamp 1679581782
transform 1 0 34944 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_363
timestamp 1679581782
transform 1 0 36000 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_370
timestamp 1679581782
transform 1 0 36672 0 -1 6804
box -48 -56 720 834
use sg13g2_fill_2  FILLER_7_377
timestamp 1677580104
transform 1 0 37344 0 -1 6804
box -48 -56 240 834
use sg13g2_fill_2  FILLER_7_383
timestamp 1677580104
transform 1 0 37920 0 -1 6804
box -48 -56 240 834
use sg13g2_fill_2  FILLER_7_410
timestamp 1677580104
transform 1 0 40512 0 -1 6804
box -48 -56 240 834
use sg13g2_fill_1  FILLER_7_412
timestamp 1677579658
transform 1 0 40704 0 -1 6804
box -48 -56 144 834
use sg13g2_fill_2  FILLER_7_421
timestamp 1677580104
transform 1 0 41568 0 -1 6804
box -48 -56 240 834
use sg13g2_fill_1  FILLER_7_423
timestamp 1677579658
transform 1 0 41760 0 -1 6804
box -48 -56 144 834
use sg13g2_decap_4  FILLER_8_0
timestamp 1679577901
transform 1 0 1152 0 1 6804
box -48 -56 432 834
use sg13g2_fill_1  FILLER_8_4
timestamp 1677579658
transform 1 0 1536 0 1 6804
box -48 -56 144 834
use sg13g2_fill_2  FILLER_8_22
timestamp 1677580104
transform 1 0 3264 0 1 6804
box -48 -56 240 834
use sg13g2_fill_1  FILLER_8_24
timestamp 1677579658
transform 1 0 3456 0 1 6804
box -48 -56 144 834
use sg13g2_decap_8  FILLER_8_57
timestamp 1679581782
transform 1 0 6624 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_64
timestamp 1679581782
transform 1 0 7296 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_113
timestamp 1679581782
transform 1 0 12000 0 1 6804
box -48 -56 720 834
use sg13g2_decap_4  FILLER_8_124
timestamp 1679577901
transform 1 0 13056 0 1 6804
box -48 -56 432 834
use sg13g2_fill_2  FILLER_8_128
timestamp 1677580104
transform 1 0 13440 0 1 6804
box -48 -56 240 834
use sg13g2_fill_2  FILLER_8_134
timestamp 1677580104
transform 1 0 14016 0 1 6804
box -48 -56 240 834
use sg13g2_fill_1  FILLER_8_136
timestamp 1677579658
transform 1 0 14208 0 1 6804
box -48 -56 144 834
use sg13g2_decap_4  FILLER_8_188
timestamp 1679577901
transform 1 0 19200 0 1 6804
box -48 -56 432 834
use sg13g2_fill_1  FILLER_8_209
timestamp 1677579658
transform 1 0 21216 0 1 6804
box -48 -56 144 834
use sg13g2_decap_8  FILLER_8_227
timestamp 1679581782
transform 1 0 22944 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_234
timestamp 1679581782
transform 1 0 23616 0 1 6804
box -48 -56 720 834
use sg13g2_fill_1  FILLER_8_258
timestamp 1677579658
transform 1 0 25920 0 1 6804
box -48 -56 144 834
use sg13g2_decap_8  FILLER_8_293
timestamp 1679581782
transform 1 0 29280 0 1 6804
box -48 -56 720 834
use sg13g2_fill_2  FILLER_8_300
timestamp 1677580104
transform 1 0 29952 0 1 6804
box -48 -56 240 834
use sg13g2_fill_1  FILLER_8_319
timestamp 1677579658
transform 1 0 31776 0 1 6804
box -48 -56 144 834
use sg13g2_fill_1  FILLER_8_337
timestamp 1677579658
transform 1 0 33504 0 1 6804
box -48 -56 144 834
use sg13g2_decap_4  FILLER_8_342
timestamp 1679577901
transform 1 0 33984 0 1 6804
box -48 -56 432 834
use sg13g2_fill_1  FILLER_8_346
timestamp 1677579658
transform 1 0 34368 0 1 6804
box -48 -56 144 834
use sg13g2_fill_1  FILLER_8_364
timestamp 1677579658
transform 1 0 36096 0 1 6804
box -48 -56 144 834
use sg13g2_decap_8  FILLER_8_382
timestamp 1679581782
transform 1 0 37824 0 1 6804
box -48 -56 720 834
use sg13g2_decap_4  FILLER_8_389
timestamp 1679577901
transform 1 0 38496 0 1 6804
box -48 -56 432 834
use sg13g2_fill_2  FILLER_8_410
timestamp 1677580104
transform 1 0 40512 0 1 6804
box -48 -56 240 834
use sg13g2_fill_1  FILLER_8_412
timestamp 1677579658
transform 1 0 40704 0 1 6804
box -48 -56 144 834
use sg13g2_fill_2  FILLER_8_421
timestamp 1677580104
transform 1 0 41568 0 1 6804
box -48 -56 240 834
use sg13g2_fill_1  FILLER_8_423
timestamp 1677579658
transform 1 0 41760 0 1 6804
box -48 -56 144 834
use sg13g2_decap_8  FILLER_9_0
timestamp 1679581782
transform 1 0 1152 0 -1 8316
box -48 -56 720 834
use sg13g2_fill_2  FILLER_9_24
timestamp 1677580104
transform 1 0 3456 0 -1 8316
box -48 -56 240 834
use sg13g2_fill_2  FILLER_9_41
timestamp 1677580104
transform 1 0 5088 0 -1 8316
box -48 -56 240 834
use sg13g2_decap_8  FILLER_9_69
timestamp 1679581782
transform 1 0 7776 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_76
timestamp 1679581782
transform 1 0 8448 0 -1 8316
box -48 -56 720 834
use sg13g2_fill_2  FILLER_9_83
timestamp 1677580104
transform 1 0 9120 0 -1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_9_106
timestamp 1677579658
transform 1 0 11328 0 -1 8316
box -48 -56 144 834
use sg13g2_decap_4  FILLER_9_115
timestamp 1679577901
transform 1 0 12192 0 -1 8316
box -48 -56 432 834
use sg13g2_fill_1  FILLER_9_119
timestamp 1677579658
transform 1 0 12576 0 -1 8316
box -48 -56 144 834
use sg13g2_fill_1  FILLER_9_137
timestamp 1677579658
transform 1 0 14304 0 -1 8316
box -48 -56 144 834
use sg13g2_decap_4  FILLER_9_159
timestamp 1679577901
transform 1 0 16416 0 -1 8316
box -48 -56 432 834
use sg13g2_fill_2  FILLER_9_167
timestamp 1677580104
transform 1 0 17184 0 -1 8316
box -48 -56 240 834
use sg13g2_fill_2  FILLER_9_194
timestamp 1677580104
transform 1 0 19776 0 -1 8316
box -48 -56 240 834
use sg13g2_decap_4  FILLER_9_200
timestamp 1679577901
transform 1 0 20352 0 -1 8316
box -48 -56 432 834
use sg13g2_fill_1  FILLER_9_204
timestamp 1677579658
transform 1 0 20736 0 -1 8316
box -48 -56 144 834
use sg13g2_decap_8  FILLER_9_230
timestamp 1679581782
transform 1 0 23232 0 -1 8316
box -48 -56 720 834
use sg13g2_fill_1  FILLER_9_237
timestamp 1677579658
transform 1 0 23904 0 -1 8316
box -48 -56 144 834
use sg13g2_fill_2  FILLER_9_276
timestamp 1677580104
transform 1 0 27648 0 -1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_9_278
timestamp 1677579658
transform 1 0 27840 0 -1 8316
box -48 -56 144 834
use sg13g2_fill_1  FILLER_9_296
timestamp 1677579658
transform 1 0 29568 0 -1 8316
box -48 -56 144 834
use sg13g2_decap_4  FILLER_9_318
timestamp 1679577901
transform 1 0 31680 0 -1 8316
box -48 -56 432 834
use sg13g2_fill_1  FILLER_9_322
timestamp 1677579658
transform 1 0 32064 0 -1 8316
box -48 -56 144 834
use sg13g2_fill_2  FILLER_9_331
timestamp 1677580104
transform 1 0 32928 0 -1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_9_333
timestamp 1677579658
transform 1 0 33120 0 -1 8316
box -48 -56 144 834
use sg13g2_decap_8  FILLER_9_351
timestamp 1679581782
transform 1 0 34848 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_4  FILLER_9_358
timestamp 1679577901
transform 1 0 35520 0 -1 8316
box -48 -56 432 834
use sg13g2_fill_2  FILLER_9_362
timestamp 1677580104
transform 1 0 35904 0 -1 8316
box -48 -56 240 834
use sg13g2_fill_2  FILLER_9_406
timestamp 1677580104
transform 1 0 40128 0 -1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_9_408
timestamp 1677579658
transform 1 0 40320 0 -1 8316
box -48 -56 144 834
use sg13g2_fill_2  FILLER_9_421
timestamp 1677580104
transform 1 0 41568 0 -1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_9_423
timestamp 1677579658
transform 1 0 41760 0 -1 8316
box -48 -56 144 834
use sg13g2_decap_4  FILLER_10_0
timestamp 1679577901
transform 1 0 1152 0 1 8316
box -48 -56 432 834
use sg13g2_fill_1  FILLER_10_43
timestamp 1677579658
transform 1 0 5280 0 1 8316
box -48 -56 144 834
use sg13g2_fill_1  FILLER_10_49
timestamp 1677579658
transform 1 0 5856 0 1 8316
box -48 -56 144 834
use sg13g2_decap_4  FILLER_10_71
timestamp 1679577901
transform 1 0 7968 0 1 8316
box -48 -56 432 834
use sg13g2_fill_2  FILLER_10_96
timestamp 1677580104
transform 1 0 10368 0 1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_10_98
timestamp 1677579658
transform 1 0 10560 0 1 8316
box -48 -56 144 834
use sg13g2_fill_2  FILLER_10_120
timestamp 1677580104
transform 1 0 12672 0 1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_10_122
timestamp 1677579658
transform 1 0 12864 0 1 8316
box -48 -56 144 834
use sg13g2_fill_2  FILLER_10_161
timestamp 1677580104
transform 1 0 16608 0 1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_10_163
timestamp 1677579658
transform 1 0 16800 0 1 8316
box -48 -56 144 834
use sg13g2_fill_1  FILLER_10_202
timestamp 1677579658
transform 1 0 20544 0 1 8316
box -48 -56 144 834
use sg13g2_fill_2  FILLER_10_241
timestamp 1677580104
transform 1 0 24288 0 1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_10_247
timestamp 1677579658
transform 1 0 24864 0 1 8316
box -48 -56 144 834
use sg13g2_fill_1  FILLER_10_252
timestamp 1677579658
transform 1 0 25344 0 1 8316
box -48 -56 144 834
use sg13g2_decap_8  FILLER_10_282
timestamp 1679581782
transform 1 0 28224 0 1 8316
box -48 -56 720 834
use sg13g2_fill_1  FILLER_10_322
timestamp 1677579658
transform 1 0 32064 0 1 8316
box -48 -56 144 834
use sg13g2_fill_1  FILLER_10_344
timestamp 1677579658
transform 1 0 34176 0 1 8316
box -48 -56 144 834
use sg13g2_fill_2  FILLER_10_355
timestamp 1677580104
transform 1 0 35232 0 1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_10_357
timestamp 1677579658
transform 1 0 35424 0 1 8316
box -48 -56 144 834
use sg13g2_decap_4  FILLER_10_396
timestamp 1679577901
transform 1 0 39168 0 1 8316
box -48 -56 432 834
use sg13g2_fill_1  FILLER_10_400
timestamp 1677579658
transform 1 0 39552 0 1 8316
box -48 -56 144 834
use sg13g2_fill_2  FILLER_10_421
timestamp 1677580104
transform 1 0 41568 0 1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_10_423
timestamp 1677579658
transform 1 0 41760 0 1 8316
box -48 -56 144 834
use sg13g2_decap_8  FILLER_11_0
timestamp 1679581782
transform 1 0 1152 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_118
timestamp 1679581782
transform 1 0 12480 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_125
timestamp 1679581782
transform 1 0 13152 0 -1 9828
box -48 -56 720 834
use sg13g2_fill_2  FILLER_11_132
timestamp 1677580104
transform 1 0 13824 0 -1 9828
box -48 -56 240 834
use sg13g2_fill_1  FILLER_11_134
timestamp 1677579658
transform 1 0 14016 0 -1 9828
box -48 -56 144 834
use sg13g2_decap_4  FILLER_11_139
timestamp 1679577901
transform 1 0 14496 0 -1 9828
box -48 -56 432 834
use sg13g2_fill_2  FILLER_11_160
timestamp 1677580104
transform 1 0 16512 0 -1 9828
box -48 -56 240 834
use sg13g2_fill_1  FILLER_11_162
timestamp 1677579658
transform 1 0 16704 0 -1 9828
box -48 -56 144 834
use sg13g2_decap_8  FILLER_11_167
timestamp 1679581782
transform 1 0 17184 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_174
timestamp 1679581782
transform 1 0 17856 0 -1 9828
box -48 -56 720 834
use sg13g2_fill_2  FILLER_11_181
timestamp 1677580104
transform 1 0 18528 0 -1 9828
box -48 -56 240 834
use sg13g2_decap_8  FILLER_11_204
timestamp 1679581782
transform 1 0 20736 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_211
timestamp 1679581782
transform 1 0 21408 0 -1 9828
box -48 -56 720 834
use sg13g2_fill_1  FILLER_11_218
timestamp 1677579658
transform 1 0 22080 0 -1 9828
box -48 -56 144 834
use sg13g2_fill_1  FILLER_11_223
timestamp 1677579658
transform 1 0 22560 0 -1 9828
box -48 -56 144 834
use sg13g2_decap_8  FILLER_11_258
timestamp 1679581782
transform 1 0 25920 0 -1 9828
box -48 -56 720 834
use sg13g2_fill_2  FILLER_11_265
timestamp 1677580104
transform 1 0 26592 0 -1 9828
box -48 -56 240 834
use sg13g2_fill_1  FILLER_11_267
timestamp 1677579658
transform 1 0 26784 0 -1 9828
box -48 -56 144 834
use sg13g2_decap_8  FILLER_11_285
timestamp 1679581782
transform 1 0 28512 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_4  FILLER_11_292
timestamp 1679577901
transform 1 0 29184 0 -1 9828
box -48 -56 432 834
use sg13g2_fill_1  FILLER_11_329
timestamp 1677579658
transform 1 0 32736 0 -1 9828
box -48 -56 144 834
use sg13g2_decap_4  FILLER_11_347
timestamp 1679577901
transform 1 0 34464 0 -1 9828
box -48 -56 432 834
use sg13g2_fill_1  FILLER_11_351
timestamp 1677579658
transform 1 0 34848 0 -1 9828
box -48 -56 144 834
use sg13g2_decap_4  FILLER_11_369
timestamp 1679577901
transform 1 0 36576 0 -1 9828
box -48 -56 432 834
use sg13g2_fill_2  FILLER_11_377
timestamp 1677580104
transform 1 0 37344 0 -1 9828
box -48 -56 240 834
use sg13g2_fill_2  FILLER_11_383
timestamp 1677580104
transform 1 0 37920 0 -1 9828
box -48 -56 240 834
use sg13g2_fill_1  FILLER_11_385
timestamp 1677579658
transform 1 0 38112 0 -1 9828
box -48 -56 144 834
use sg13g2_decap_8  FILLER_11_403
timestamp 1679581782
transform 1 0 39840 0 -1 9828
box -48 -56 720 834
use sg13g2_fill_2  FILLER_11_410
timestamp 1677580104
transform 1 0 40512 0 -1 9828
box -48 -56 240 834
use sg13g2_fill_1  FILLER_11_412
timestamp 1677579658
transform 1 0 40704 0 -1 9828
box -48 -56 144 834
use sg13g2_fill_2  FILLER_11_421
timestamp 1677580104
transform 1 0 41568 0 -1 9828
box -48 -56 240 834
use sg13g2_fill_1  FILLER_11_423
timestamp 1677579658
transform 1 0 41760 0 -1 9828
box -48 -56 144 834
<< labels >>
flabel metal2 s 2936 0 3016 80 0 FreeSans 320 0 0 0 A_I_top
port 0 nsew signal output
flabel metal2 s 1784 0 1864 80 0 FreeSans 320 0 0 0 A_O_top
port 1 nsew signal input
flabel metal2 s 4088 0 4168 80 0 FreeSans 320 0 0 0 A_T_top
port 2 nsew signal output
flabel metal2 s 8696 0 8776 80 0 FreeSans 320 0 0 0 A_config_C_bit0
port 3 nsew signal output
flabel metal2 s 9848 0 9928 80 0 FreeSans 320 0 0 0 A_config_C_bit1
port 4 nsew signal output
flabel metal2 s 11000 0 11080 80 0 FreeSans 320 0 0 0 A_config_C_bit2
port 5 nsew signal output
flabel metal2 s 12152 0 12232 80 0 FreeSans 320 0 0 0 A_config_C_bit3
port 6 nsew signal output
flabel metal2 s 6392 0 6472 80 0 FreeSans 320 0 0 0 B_I_top
port 7 nsew signal output
flabel metal2 s 5240 0 5320 80 0 FreeSans 320 0 0 0 B_O_top
port 8 nsew signal input
flabel metal2 s 7544 0 7624 80 0 FreeSans 320 0 0 0 B_T_top
port 9 nsew signal output
flabel metal2 s 13304 0 13384 80 0 FreeSans 320 0 0 0 B_config_C_bit0
port 10 nsew signal output
flabel metal2 s 14456 0 14536 80 0 FreeSans 320 0 0 0 B_config_C_bit1
port 11 nsew signal output
flabel metal2 s 15608 0 15688 80 0 FreeSans 320 0 0 0 B_config_C_bit2
port 12 nsew signal output
flabel metal2 s 16760 0 16840 80 0 FreeSans 320 0 0 0 B_config_C_bit3
port 13 nsew signal output
flabel metal2 s 19448 10672 19528 10752 0 FreeSans 320 0 0 0 Co
port 14 nsew signal output
flabel metal3 s 0 44 80 124 0 FreeSans 320 0 0 0 FrameData[0]
port 15 nsew signal input
flabel metal3 s 0 3404 80 3484 0 FreeSans 320 0 0 0 FrameData[10]
port 16 nsew signal input
flabel metal3 s 0 3740 80 3820 0 FreeSans 320 0 0 0 FrameData[11]
port 17 nsew signal input
flabel metal3 s 0 4076 80 4156 0 FreeSans 320 0 0 0 FrameData[12]
port 18 nsew signal input
flabel metal3 s 0 4412 80 4492 0 FreeSans 320 0 0 0 FrameData[13]
port 19 nsew signal input
flabel metal3 s 0 4748 80 4828 0 FreeSans 320 0 0 0 FrameData[14]
port 20 nsew signal input
flabel metal3 s 0 5084 80 5164 0 FreeSans 320 0 0 0 FrameData[15]
port 21 nsew signal input
flabel metal3 s 0 5420 80 5500 0 FreeSans 320 0 0 0 FrameData[16]
port 22 nsew signal input
flabel metal3 s 0 5756 80 5836 0 FreeSans 320 0 0 0 FrameData[17]
port 23 nsew signal input
flabel metal3 s 0 6092 80 6172 0 FreeSans 320 0 0 0 FrameData[18]
port 24 nsew signal input
flabel metal3 s 0 6428 80 6508 0 FreeSans 320 0 0 0 FrameData[19]
port 25 nsew signal input
flabel metal3 s 0 380 80 460 0 FreeSans 320 0 0 0 FrameData[1]
port 26 nsew signal input
flabel metal3 s 0 6764 80 6844 0 FreeSans 320 0 0 0 FrameData[20]
port 27 nsew signal input
flabel metal3 s 0 7100 80 7180 0 FreeSans 320 0 0 0 FrameData[21]
port 28 nsew signal input
flabel metal3 s 0 7436 80 7516 0 FreeSans 320 0 0 0 FrameData[22]
port 29 nsew signal input
flabel metal3 s 0 7772 80 7852 0 FreeSans 320 0 0 0 FrameData[23]
port 30 nsew signal input
flabel metal3 s 0 8108 80 8188 0 FreeSans 320 0 0 0 FrameData[24]
port 31 nsew signal input
flabel metal3 s 0 8444 80 8524 0 FreeSans 320 0 0 0 FrameData[25]
port 32 nsew signal input
flabel metal3 s 0 8780 80 8860 0 FreeSans 320 0 0 0 FrameData[26]
port 33 nsew signal input
flabel metal3 s 0 9116 80 9196 0 FreeSans 320 0 0 0 FrameData[27]
port 34 nsew signal input
flabel metal3 s 0 9452 80 9532 0 FreeSans 320 0 0 0 FrameData[28]
port 35 nsew signal input
flabel metal3 s 0 9788 80 9868 0 FreeSans 320 0 0 0 FrameData[29]
port 36 nsew signal input
flabel metal3 s 0 716 80 796 0 FreeSans 320 0 0 0 FrameData[2]
port 37 nsew signal input
flabel metal3 s 0 10124 80 10204 0 FreeSans 320 0 0 0 FrameData[30]
port 38 nsew signal input
flabel metal3 s 0 10460 80 10540 0 FreeSans 320 0 0 0 FrameData[31]
port 39 nsew signal input
flabel metal3 s 0 1052 80 1132 0 FreeSans 320 0 0 0 FrameData[3]
port 40 nsew signal input
flabel metal3 s 0 1388 80 1468 0 FreeSans 320 0 0 0 FrameData[4]
port 41 nsew signal input
flabel metal3 s 0 1724 80 1804 0 FreeSans 320 0 0 0 FrameData[5]
port 42 nsew signal input
flabel metal3 s 0 2060 80 2140 0 FreeSans 320 0 0 0 FrameData[6]
port 43 nsew signal input
flabel metal3 s 0 2396 80 2476 0 FreeSans 320 0 0 0 FrameData[7]
port 44 nsew signal input
flabel metal3 s 0 2732 80 2812 0 FreeSans 320 0 0 0 FrameData[8]
port 45 nsew signal input
flabel metal3 s 0 3068 80 3148 0 FreeSans 320 0 0 0 FrameData[9]
port 46 nsew signal input
flabel metal3 s 42928 44 43008 124 0 FreeSans 320 0 0 0 FrameData_O[0]
port 47 nsew signal output
flabel metal3 s 42928 3404 43008 3484 0 FreeSans 320 0 0 0 FrameData_O[10]
port 48 nsew signal output
flabel metal3 s 42928 3740 43008 3820 0 FreeSans 320 0 0 0 FrameData_O[11]
port 49 nsew signal output
flabel metal3 s 42928 4076 43008 4156 0 FreeSans 320 0 0 0 FrameData_O[12]
port 50 nsew signal output
flabel metal3 s 42928 4412 43008 4492 0 FreeSans 320 0 0 0 FrameData_O[13]
port 51 nsew signal output
flabel metal3 s 42928 4748 43008 4828 0 FreeSans 320 0 0 0 FrameData_O[14]
port 52 nsew signal output
flabel metal3 s 42928 5084 43008 5164 0 FreeSans 320 0 0 0 FrameData_O[15]
port 53 nsew signal output
flabel metal3 s 42928 5420 43008 5500 0 FreeSans 320 0 0 0 FrameData_O[16]
port 54 nsew signal output
flabel metal3 s 42928 5756 43008 5836 0 FreeSans 320 0 0 0 FrameData_O[17]
port 55 nsew signal output
flabel metal3 s 42928 6092 43008 6172 0 FreeSans 320 0 0 0 FrameData_O[18]
port 56 nsew signal output
flabel metal3 s 42928 6428 43008 6508 0 FreeSans 320 0 0 0 FrameData_O[19]
port 57 nsew signal output
flabel metal3 s 42928 380 43008 460 0 FreeSans 320 0 0 0 FrameData_O[1]
port 58 nsew signal output
flabel metal3 s 42928 6764 43008 6844 0 FreeSans 320 0 0 0 FrameData_O[20]
port 59 nsew signal output
flabel metal3 s 42928 7100 43008 7180 0 FreeSans 320 0 0 0 FrameData_O[21]
port 60 nsew signal output
flabel metal3 s 42928 7436 43008 7516 0 FreeSans 320 0 0 0 FrameData_O[22]
port 61 nsew signal output
flabel metal3 s 42928 7772 43008 7852 0 FreeSans 320 0 0 0 FrameData_O[23]
port 62 nsew signal output
flabel metal3 s 42928 8108 43008 8188 0 FreeSans 320 0 0 0 FrameData_O[24]
port 63 nsew signal output
flabel metal3 s 42928 8444 43008 8524 0 FreeSans 320 0 0 0 FrameData_O[25]
port 64 nsew signal output
flabel metal3 s 42928 8780 43008 8860 0 FreeSans 320 0 0 0 FrameData_O[26]
port 65 nsew signal output
flabel metal3 s 42928 9116 43008 9196 0 FreeSans 320 0 0 0 FrameData_O[27]
port 66 nsew signal output
flabel metal3 s 42928 9452 43008 9532 0 FreeSans 320 0 0 0 FrameData_O[28]
port 67 nsew signal output
flabel metal3 s 42928 9788 43008 9868 0 FreeSans 320 0 0 0 FrameData_O[29]
port 68 nsew signal output
flabel metal3 s 42928 716 43008 796 0 FreeSans 320 0 0 0 FrameData_O[2]
port 69 nsew signal output
flabel metal3 s 42928 10124 43008 10204 0 FreeSans 320 0 0 0 FrameData_O[30]
port 70 nsew signal output
flabel metal3 s 42928 10460 43008 10540 0 FreeSans 320 0 0 0 FrameData_O[31]
port 71 nsew signal output
flabel metal3 s 42928 1052 43008 1132 0 FreeSans 320 0 0 0 FrameData_O[3]
port 72 nsew signal output
flabel metal3 s 42928 1388 43008 1468 0 FreeSans 320 0 0 0 FrameData_O[4]
port 73 nsew signal output
flabel metal3 s 42928 1724 43008 1804 0 FreeSans 320 0 0 0 FrameData_O[5]
port 74 nsew signal output
flabel metal3 s 42928 2060 43008 2140 0 FreeSans 320 0 0 0 FrameData_O[6]
port 75 nsew signal output
flabel metal3 s 42928 2396 43008 2476 0 FreeSans 320 0 0 0 FrameData_O[7]
port 76 nsew signal output
flabel metal3 s 42928 2732 43008 2812 0 FreeSans 320 0 0 0 FrameData_O[8]
port 77 nsew signal output
flabel metal3 s 42928 3068 43008 3148 0 FreeSans 320 0 0 0 FrameData_O[9]
port 78 nsew signal output
flabel metal2 s 19064 0 19144 80 0 FreeSans 320 0 0 0 FrameStrobe[0]
port 79 nsew signal input
flabel metal2 s 30584 0 30664 80 0 FreeSans 320 0 0 0 FrameStrobe[10]
port 80 nsew signal input
flabel metal2 s 31736 0 31816 80 0 FreeSans 320 0 0 0 FrameStrobe[11]
port 81 nsew signal input
flabel metal2 s 32888 0 32968 80 0 FreeSans 320 0 0 0 FrameStrobe[12]
port 82 nsew signal input
flabel metal2 s 34040 0 34120 80 0 FreeSans 320 0 0 0 FrameStrobe[13]
port 83 nsew signal input
flabel metal2 s 35192 0 35272 80 0 FreeSans 320 0 0 0 FrameStrobe[14]
port 84 nsew signal input
flabel metal2 s 36344 0 36424 80 0 FreeSans 320 0 0 0 FrameStrobe[15]
port 85 nsew signal input
flabel metal2 s 37496 0 37576 80 0 FreeSans 320 0 0 0 FrameStrobe[16]
port 86 nsew signal input
flabel metal2 s 38648 0 38728 80 0 FreeSans 320 0 0 0 FrameStrobe[17]
port 87 nsew signal input
flabel metal2 s 39800 0 39880 80 0 FreeSans 320 0 0 0 FrameStrobe[18]
port 88 nsew signal input
flabel metal2 s 40952 0 41032 80 0 FreeSans 320 0 0 0 FrameStrobe[19]
port 89 nsew signal input
flabel metal2 s 20216 0 20296 80 0 FreeSans 320 0 0 0 FrameStrobe[1]
port 90 nsew signal input
flabel metal2 s 21368 0 21448 80 0 FreeSans 320 0 0 0 FrameStrobe[2]
port 91 nsew signal input
flabel metal2 s 22520 0 22600 80 0 FreeSans 320 0 0 0 FrameStrobe[3]
port 92 nsew signal input
flabel metal2 s 23672 0 23752 80 0 FreeSans 320 0 0 0 FrameStrobe[4]
port 93 nsew signal input
flabel metal2 s 24824 0 24904 80 0 FreeSans 320 0 0 0 FrameStrobe[5]
port 94 nsew signal input
flabel metal2 s 25976 0 26056 80 0 FreeSans 320 0 0 0 FrameStrobe[6]
port 95 nsew signal input
flabel metal2 s 27128 0 27208 80 0 FreeSans 320 0 0 0 FrameStrobe[7]
port 96 nsew signal input
flabel metal2 s 28280 0 28360 80 0 FreeSans 320 0 0 0 FrameStrobe[8]
port 97 nsew signal input
flabel metal2 s 29432 0 29512 80 0 FreeSans 320 0 0 0 FrameStrobe[9]
port 98 nsew signal input
flabel metal2 s 29816 10672 29896 10752 0 FreeSans 320 0 0 0 FrameStrobe_O[0]
port 99 nsew signal output
flabel metal2 s 31736 10672 31816 10752 0 FreeSans 320 0 0 0 FrameStrobe_O[10]
port 100 nsew signal output
flabel metal2 s 31928 10672 32008 10752 0 FreeSans 320 0 0 0 FrameStrobe_O[11]
port 101 nsew signal output
flabel metal2 s 32120 10672 32200 10752 0 FreeSans 320 0 0 0 FrameStrobe_O[12]
port 102 nsew signal output
flabel metal2 s 32312 10672 32392 10752 0 FreeSans 320 0 0 0 FrameStrobe_O[13]
port 103 nsew signal output
flabel metal2 s 32504 10672 32584 10752 0 FreeSans 320 0 0 0 FrameStrobe_O[14]
port 104 nsew signal output
flabel metal2 s 32696 10672 32776 10752 0 FreeSans 320 0 0 0 FrameStrobe_O[15]
port 105 nsew signal output
flabel metal2 s 32888 10672 32968 10752 0 FreeSans 320 0 0 0 FrameStrobe_O[16]
port 106 nsew signal output
flabel metal2 s 33080 10672 33160 10752 0 FreeSans 320 0 0 0 FrameStrobe_O[17]
port 107 nsew signal output
flabel metal2 s 33272 10672 33352 10752 0 FreeSans 320 0 0 0 FrameStrobe_O[18]
port 108 nsew signal output
flabel metal2 s 33464 10672 33544 10752 0 FreeSans 320 0 0 0 FrameStrobe_O[19]
port 109 nsew signal output
flabel metal2 s 30008 10672 30088 10752 0 FreeSans 320 0 0 0 FrameStrobe_O[1]
port 110 nsew signal output
flabel metal2 s 30200 10672 30280 10752 0 FreeSans 320 0 0 0 FrameStrobe_O[2]
port 111 nsew signal output
flabel metal2 s 30392 10672 30472 10752 0 FreeSans 320 0 0 0 FrameStrobe_O[3]
port 112 nsew signal output
flabel metal2 s 30584 10672 30664 10752 0 FreeSans 320 0 0 0 FrameStrobe_O[4]
port 113 nsew signal output
flabel metal2 s 30776 10672 30856 10752 0 FreeSans 320 0 0 0 FrameStrobe_O[5]
port 114 nsew signal output
flabel metal2 s 30968 10672 31048 10752 0 FreeSans 320 0 0 0 FrameStrobe_O[6]
port 115 nsew signal output
flabel metal2 s 31160 10672 31240 10752 0 FreeSans 320 0 0 0 FrameStrobe_O[7]
port 116 nsew signal output
flabel metal2 s 31352 10672 31432 10752 0 FreeSans 320 0 0 0 FrameStrobe_O[8]
port 117 nsew signal output
flabel metal2 s 31544 10672 31624 10752 0 FreeSans 320 0 0 0 FrameStrobe_O[9]
port 118 nsew signal output
flabel metal2 s 9464 10672 9544 10752 0 FreeSans 320 0 0 0 N1BEG[0]
port 119 nsew signal output
flabel metal2 s 9656 10672 9736 10752 0 FreeSans 320 0 0 0 N1BEG[1]
port 120 nsew signal output
flabel metal2 s 9848 10672 9928 10752 0 FreeSans 320 0 0 0 N1BEG[2]
port 121 nsew signal output
flabel metal2 s 10040 10672 10120 10752 0 FreeSans 320 0 0 0 N1BEG[3]
port 122 nsew signal output
flabel metal2 s 10232 10672 10312 10752 0 FreeSans 320 0 0 0 N2BEG[0]
port 123 nsew signal output
flabel metal2 s 10424 10672 10504 10752 0 FreeSans 320 0 0 0 N2BEG[1]
port 124 nsew signal output
flabel metal2 s 10616 10672 10696 10752 0 FreeSans 320 0 0 0 N2BEG[2]
port 125 nsew signal output
flabel metal2 s 10808 10672 10888 10752 0 FreeSans 320 0 0 0 N2BEG[3]
port 126 nsew signal output
flabel metal2 s 11000 10672 11080 10752 0 FreeSans 320 0 0 0 N2BEG[4]
port 127 nsew signal output
flabel metal2 s 11192 10672 11272 10752 0 FreeSans 320 0 0 0 N2BEG[5]
port 128 nsew signal output
flabel metal2 s 11384 10672 11464 10752 0 FreeSans 320 0 0 0 N2BEG[6]
port 129 nsew signal output
flabel metal2 s 11576 10672 11656 10752 0 FreeSans 320 0 0 0 N2BEG[7]
port 130 nsew signal output
flabel metal2 s 11768 10672 11848 10752 0 FreeSans 320 0 0 0 N2BEGb[0]
port 131 nsew signal output
flabel metal2 s 11960 10672 12040 10752 0 FreeSans 320 0 0 0 N2BEGb[1]
port 132 nsew signal output
flabel metal2 s 12152 10672 12232 10752 0 FreeSans 320 0 0 0 N2BEGb[2]
port 133 nsew signal output
flabel metal2 s 12344 10672 12424 10752 0 FreeSans 320 0 0 0 N2BEGb[3]
port 134 nsew signal output
flabel metal2 s 12536 10672 12616 10752 0 FreeSans 320 0 0 0 N2BEGb[4]
port 135 nsew signal output
flabel metal2 s 12728 10672 12808 10752 0 FreeSans 320 0 0 0 N2BEGb[5]
port 136 nsew signal output
flabel metal2 s 12920 10672 13000 10752 0 FreeSans 320 0 0 0 N2BEGb[6]
port 137 nsew signal output
flabel metal2 s 13112 10672 13192 10752 0 FreeSans 320 0 0 0 N2BEGb[7]
port 138 nsew signal output
flabel metal2 s 13304 10672 13384 10752 0 FreeSans 320 0 0 0 N4BEG[0]
port 139 nsew signal output
flabel metal2 s 15224 10672 15304 10752 0 FreeSans 320 0 0 0 N4BEG[10]
port 140 nsew signal output
flabel metal2 s 15416 10672 15496 10752 0 FreeSans 320 0 0 0 N4BEG[11]
port 141 nsew signal output
flabel metal2 s 15608 10672 15688 10752 0 FreeSans 320 0 0 0 N4BEG[12]
port 142 nsew signal output
flabel metal2 s 15800 10672 15880 10752 0 FreeSans 320 0 0 0 N4BEG[13]
port 143 nsew signal output
flabel metal2 s 15992 10672 16072 10752 0 FreeSans 320 0 0 0 N4BEG[14]
port 144 nsew signal output
flabel metal2 s 16184 10672 16264 10752 0 FreeSans 320 0 0 0 N4BEG[15]
port 145 nsew signal output
flabel metal2 s 13496 10672 13576 10752 0 FreeSans 320 0 0 0 N4BEG[1]
port 146 nsew signal output
flabel metal2 s 13688 10672 13768 10752 0 FreeSans 320 0 0 0 N4BEG[2]
port 147 nsew signal output
flabel metal2 s 13880 10672 13960 10752 0 FreeSans 320 0 0 0 N4BEG[3]
port 148 nsew signal output
flabel metal2 s 14072 10672 14152 10752 0 FreeSans 320 0 0 0 N4BEG[4]
port 149 nsew signal output
flabel metal2 s 14264 10672 14344 10752 0 FreeSans 320 0 0 0 N4BEG[5]
port 150 nsew signal output
flabel metal2 s 14456 10672 14536 10752 0 FreeSans 320 0 0 0 N4BEG[6]
port 151 nsew signal output
flabel metal2 s 14648 10672 14728 10752 0 FreeSans 320 0 0 0 N4BEG[7]
port 152 nsew signal output
flabel metal2 s 14840 10672 14920 10752 0 FreeSans 320 0 0 0 N4BEG[8]
port 153 nsew signal output
flabel metal2 s 15032 10672 15112 10752 0 FreeSans 320 0 0 0 N4BEG[9]
port 154 nsew signal output
flabel metal2 s 16376 10672 16456 10752 0 FreeSans 320 0 0 0 NN4BEG[0]
port 155 nsew signal output
flabel metal2 s 18296 10672 18376 10752 0 FreeSans 320 0 0 0 NN4BEG[10]
port 156 nsew signal output
flabel metal2 s 18488 10672 18568 10752 0 FreeSans 320 0 0 0 NN4BEG[11]
port 157 nsew signal output
flabel metal2 s 18680 10672 18760 10752 0 FreeSans 320 0 0 0 NN4BEG[12]
port 158 nsew signal output
flabel metal2 s 18872 10672 18952 10752 0 FreeSans 320 0 0 0 NN4BEG[13]
port 159 nsew signal output
flabel metal2 s 19064 10672 19144 10752 0 FreeSans 320 0 0 0 NN4BEG[14]
port 160 nsew signal output
flabel metal2 s 19256 10672 19336 10752 0 FreeSans 320 0 0 0 NN4BEG[15]
port 161 nsew signal output
flabel metal2 s 16568 10672 16648 10752 0 FreeSans 320 0 0 0 NN4BEG[1]
port 162 nsew signal output
flabel metal2 s 16760 10672 16840 10752 0 FreeSans 320 0 0 0 NN4BEG[2]
port 163 nsew signal output
flabel metal2 s 16952 10672 17032 10752 0 FreeSans 320 0 0 0 NN4BEG[3]
port 164 nsew signal output
flabel metal2 s 17144 10672 17224 10752 0 FreeSans 320 0 0 0 NN4BEG[4]
port 165 nsew signal output
flabel metal2 s 17336 10672 17416 10752 0 FreeSans 320 0 0 0 NN4BEG[5]
port 166 nsew signal output
flabel metal2 s 17528 10672 17608 10752 0 FreeSans 320 0 0 0 NN4BEG[6]
port 167 nsew signal output
flabel metal2 s 17720 10672 17800 10752 0 FreeSans 320 0 0 0 NN4BEG[7]
port 168 nsew signal output
flabel metal2 s 17912 10672 17992 10752 0 FreeSans 320 0 0 0 NN4BEG[8]
port 169 nsew signal output
flabel metal2 s 18104 10672 18184 10752 0 FreeSans 320 0 0 0 NN4BEG[9]
port 170 nsew signal output
flabel metal2 s 19640 10672 19720 10752 0 FreeSans 320 0 0 0 S1END[0]
port 171 nsew signal input
flabel metal2 s 19832 10672 19912 10752 0 FreeSans 320 0 0 0 S1END[1]
port 172 nsew signal input
flabel metal2 s 20024 10672 20104 10752 0 FreeSans 320 0 0 0 S1END[2]
port 173 nsew signal input
flabel metal2 s 20216 10672 20296 10752 0 FreeSans 320 0 0 0 S1END[3]
port 174 nsew signal input
flabel metal2 s 21944 10672 22024 10752 0 FreeSans 320 0 0 0 S2END[0]
port 175 nsew signal input
flabel metal2 s 22136 10672 22216 10752 0 FreeSans 320 0 0 0 S2END[1]
port 176 nsew signal input
flabel metal2 s 22328 10672 22408 10752 0 FreeSans 320 0 0 0 S2END[2]
port 177 nsew signal input
flabel metal2 s 22520 10672 22600 10752 0 FreeSans 320 0 0 0 S2END[3]
port 178 nsew signal input
flabel metal2 s 22712 10672 22792 10752 0 FreeSans 320 0 0 0 S2END[4]
port 179 nsew signal input
flabel metal2 s 22904 10672 22984 10752 0 FreeSans 320 0 0 0 S2END[5]
port 180 nsew signal input
flabel metal2 s 23096 10672 23176 10752 0 FreeSans 320 0 0 0 S2END[6]
port 181 nsew signal input
flabel metal2 s 23288 10672 23368 10752 0 FreeSans 320 0 0 0 S2END[7]
port 182 nsew signal input
flabel metal2 s 20408 10672 20488 10752 0 FreeSans 320 0 0 0 S2MID[0]
port 183 nsew signal input
flabel metal2 s 20600 10672 20680 10752 0 FreeSans 320 0 0 0 S2MID[1]
port 184 nsew signal input
flabel metal2 s 20792 10672 20872 10752 0 FreeSans 320 0 0 0 S2MID[2]
port 185 nsew signal input
flabel metal2 s 20984 10672 21064 10752 0 FreeSans 320 0 0 0 S2MID[3]
port 186 nsew signal input
flabel metal2 s 21176 10672 21256 10752 0 FreeSans 320 0 0 0 S2MID[4]
port 187 nsew signal input
flabel metal2 s 21368 10672 21448 10752 0 FreeSans 320 0 0 0 S2MID[5]
port 188 nsew signal input
flabel metal2 s 21560 10672 21640 10752 0 FreeSans 320 0 0 0 S2MID[6]
port 189 nsew signal input
flabel metal2 s 21752 10672 21832 10752 0 FreeSans 320 0 0 0 S2MID[7]
port 190 nsew signal input
flabel metal2 s 23480 10672 23560 10752 0 FreeSans 320 0 0 0 S4END[0]
port 191 nsew signal input
flabel metal2 s 25400 10672 25480 10752 0 FreeSans 320 0 0 0 S4END[10]
port 192 nsew signal input
flabel metal2 s 25592 10672 25672 10752 0 FreeSans 320 0 0 0 S4END[11]
port 193 nsew signal input
flabel metal2 s 25784 10672 25864 10752 0 FreeSans 320 0 0 0 S4END[12]
port 194 nsew signal input
flabel metal2 s 25976 10672 26056 10752 0 FreeSans 320 0 0 0 S4END[13]
port 195 nsew signal input
flabel metal2 s 26168 10672 26248 10752 0 FreeSans 320 0 0 0 S4END[14]
port 196 nsew signal input
flabel metal2 s 26360 10672 26440 10752 0 FreeSans 320 0 0 0 S4END[15]
port 197 nsew signal input
flabel metal2 s 23672 10672 23752 10752 0 FreeSans 320 0 0 0 S4END[1]
port 198 nsew signal input
flabel metal2 s 23864 10672 23944 10752 0 FreeSans 320 0 0 0 S4END[2]
port 199 nsew signal input
flabel metal2 s 24056 10672 24136 10752 0 FreeSans 320 0 0 0 S4END[3]
port 200 nsew signal input
flabel metal2 s 24248 10672 24328 10752 0 FreeSans 320 0 0 0 S4END[4]
port 201 nsew signal input
flabel metal2 s 24440 10672 24520 10752 0 FreeSans 320 0 0 0 S4END[5]
port 202 nsew signal input
flabel metal2 s 24632 10672 24712 10752 0 FreeSans 320 0 0 0 S4END[6]
port 203 nsew signal input
flabel metal2 s 24824 10672 24904 10752 0 FreeSans 320 0 0 0 S4END[7]
port 204 nsew signal input
flabel metal2 s 25016 10672 25096 10752 0 FreeSans 320 0 0 0 S4END[8]
port 205 nsew signal input
flabel metal2 s 25208 10672 25288 10752 0 FreeSans 320 0 0 0 S4END[9]
port 206 nsew signal input
flabel metal2 s 26552 10672 26632 10752 0 FreeSans 320 0 0 0 SS4END[0]
port 207 nsew signal input
flabel metal2 s 28472 10672 28552 10752 0 FreeSans 320 0 0 0 SS4END[10]
port 208 nsew signal input
flabel metal2 s 28664 10672 28744 10752 0 FreeSans 320 0 0 0 SS4END[11]
port 209 nsew signal input
flabel metal2 s 28856 10672 28936 10752 0 FreeSans 320 0 0 0 SS4END[12]
port 210 nsew signal input
flabel metal2 s 29048 10672 29128 10752 0 FreeSans 320 0 0 0 SS4END[13]
port 211 nsew signal input
flabel metal2 s 29240 10672 29320 10752 0 FreeSans 320 0 0 0 SS4END[14]
port 212 nsew signal input
flabel metal2 s 29432 10672 29512 10752 0 FreeSans 320 0 0 0 SS4END[15]
port 213 nsew signal input
flabel metal2 s 26744 10672 26824 10752 0 FreeSans 320 0 0 0 SS4END[1]
port 214 nsew signal input
flabel metal2 s 26936 10672 27016 10752 0 FreeSans 320 0 0 0 SS4END[2]
port 215 nsew signal input
flabel metal2 s 27128 10672 27208 10752 0 FreeSans 320 0 0 0 SS4END[3]
port 216 nsew signal input
flabel metal2 s 27320 10672 27400 10752 0 FreeSans 320 0 0 0 SS4END[4]
port 217 nsew signal input
flabel metal2 s 27512 10672 27592 10752 0 FreeSans 320 0 0 0 SS4END[5]
port 218 nsew signal input
flabel metal2 s 27704 10672 27784 10752 0 FreeSans 320 0 0 0 SS4END[6]
port 219 nsew signal input
flabel metal2 s 27896 10672 27976 10752 0 FreeSans 320 0 0 0 SS4END[7]
port 220 nsew signal input
flabel metal2 s 28088 10672 28168 10752 0 FreeSans 320 0 0 0 SS4END[8]
port 221 nsew signal input
flabel metal2 s 28280 10672 28360 10752 0 FreeSans 320 0 0 0 SS4END[9]
port 222 nsew signal input
flabel metal2 s 17912 0 17992 80 0 FreeSans 320 0 0 0 UserCLK
port 223 nsew signal input
flabel metal2 s 29624 10672 29704 10752 0 FreeSans 320 0 0 0 UserCLKo
port 224 nsew signal output
flabel metal6 s 4892 0 5332 10752 0 FreeSans 2624 90 0 0 VGND
port 225 nsew ground bidirectional
flabel metal6 s 4892 0 5332 328 0 FreeSans 2624 0 0 0 VGND
port 225 nsew ground bidirectional
flabel metal6 s 4892 10424 5332 10752 0 FreeSans 2624 0 0 0 VGND
port 225 nsew ground bidirectional
flabel metal6 s 20012 0 20452 10752 0 FreeSans 2624 90 0 0 VGND
port 225 nsew ground bidirectional
flabel metal6 s 20012 0 20452 328 0 FreeSans 2624 0 0 0 VGND
port 225 nsew ground bidirectional
flabel metal6 s 20012 10424 20452 10752 0 FreeSans 2624 0 0 0 VGND
port 225 nsew ground bidirectional
flabel metal6 s 35132 0 35572 10752 0 FreeSans 2624 90 0 0 VGND
port 225 nsew ground bidirectional
flabel metal6 s 35132 0 35572 328 0 FreeSans 2624 0 0 0 VGND
port 225 nsew ground bidirectional
flabel metal6 s 35132 10424 35572 10752 0 FreeSans 2624 0 0 0 VGND
port 225 nsew ground bidirectional
flabel metal6 s 3652 0 4092 10752 0 FreeSans 2624 90 0 0 VPWR
port 226 nsew power bidirectional
flabel metal6 s 3652 0 4092 328 0 FreeSans 2624 0 0 0 VPWR
port 226 nsew power bidirectional
flabel metal6 s 3652 10424 4092 10752 0 FreeSans 2624 0 0 0 VPWR
port 226 nsew power bidirectional
flabel metal6 s 18772 0 19212 10752 0 FreeSans 2624 90 0 0 VPWR
port 226 nsew power bidirectional
flabel metal6 s 18772 0 19212 328 0 FreeSans 2624 0 0 0 VPWR
port 226 nsew power bidirectional
flabel metal6 s 18772 10424 19212 10752 0 FreeSans 2624 0 0 0 VPWR
port 226 nsew power bidirectional
flabel metal6 s 33892 0 34332 10752 0 FreeSans 2624 90 0 0 VPWR
port 226 nsew power bidirectional
flabel metal6 s 33892 0 34332 328 0 FreeSans 2624 0 0 0 VPWR
port 226 nsew power bidirectional
flabel metal6 s 33892 10424 34332 10752 0 FreeSans 2624 0 0 0 VPWR
port 226 nsew power bidirectional
rlabel metal1 21504 9828 21504 9828 0 VGND
rlabel metal1 21504 9072 21504 9072 0 VPWR
rlabel metal2 2976 1290 2976 1290 0 A_I_top
rlabel metal2 1824 954 1824 954 0 A_O_top
rlabel metal2 4128 492 4128 492 0 A_T_top
rlabel metal2 8736 492 8736 492 0 A_config_C_bit0
rlabel metal2 9888 576 9888 576 0 A_config_C_bit1
rlabel via2 11040 72 11040 72 0 A_config_C_bit2
rlabel metal2 12192 114 12192 114 0 A_config_C_bit3
rlabel metal2 6432 492 6432 492 0 B_I_top
rlabel metal2 5280 72 5280 72 0 B_O_top
rlabel metal2 7584 1290 7584 1290 0 B_T_top
rlabel via2 13344 72 13344 72 0 B_config_C_bit0
rlabel metal2 14496 492 14496 492 0 B_config_C_bit1
rlabel via2 15648 72 15648 72 0 B_config_C_bit2
rlabel metal2 16800 870 16800 870 0 B_config_C_bit3
rlabel metal2 19488 9420 19488 9420 0 Co
rlabel metal3 3342 84 3342 84 0 FrameData[0]
rlabel metal2 38784 3402 38784 3402 0 FrameData[10]
rlabel metal2 40896 3486 40896 3486 0 FrameData[11]
rlabel metal2 41280 4410 41280 4410 0 FrameData[12]
rlabel metal2 40512 4326 40512 4326 0 FrameData[13]
rlabel metal3 654 4788 654 4788 0 FrameData[14]
rlabel metal2 41328 4872 41328 4872 0 FrameData[15]
rlabel metal3 654 5460 654 5460 0 FrameData[16]
rlabel metal3 1230 5796 1230 5796 0 FrameData[17]
rlabel metal3 894 6132 894 6132 0 FrameData[18]
rlabel metal2 1776 7140 1776 7140 0 FrameData[19]
rlabel metal2 5376 714 5376 714 0 FrameData[1]
rlabel metal2 1584 4116 1584 4116 0 FrameData[20]
rlabel metal3 2160 5208 2160 5208 0 FrameData[21]
rlabel metal4 2496 840 2496 840 0 FrameData[22]
rlabel metal2 1920 4116 1920 4116 0 FrameData[23]
rlabel metal2 1632 2604 1632 2604 0 FrameData[24]
rlabel metal2 1920 7434 1920 7434 0 FrameData[25]
rlabel metal2 2112 8526 2112 8526 0 FrameData[26]
rlabel metal2 1920 9702 1920 9702 0 FrameData[27]
rlabel metal4 40896 7644 40896 7644 0 FrameData[28]
rlabel metal3 36384 966 36384 966 0 FrameData[29]
rlabel metal3 126 756 126 756 0 FrameData[2]
rlabel metal2 39024 8652 39024 8652 0 FrameData[30]
rlabel metal2 38976 7686 38976 7686 0 FrameData[31]
rlabel metal3 78 1092 78 1092 0 FrameData[3]
rlabel metal3 126 1428 126 1428 0 FrameData[4]
rlabel metal2 35616 1176 35616 1176 0 FrameData[5]
rlabel metal2 40800 2184 40800 2184 0 FrameData[6]
rlabel metal2 20064 1596 20064 1596 0 FrameData[7]
rlabel metal3 34464 2058 34464 2058 0 FrameData[8]
rlabel metal2 16320 1512 16320 1512 0 FrameData[9]
rlabel metal2 41088 546 41088 546 0 FrameData_O[0]
rlabel metal2 40704 3360 40704 3360 0 FrameData_O[10]
rlabel metal2 41088 3696 41088 3696 0 FrameData_O[11]
rlabel metal2 41472 4032 41472 4032 0 FrameData_O[12]
rlabel metal2 40704 4410 40704 4410 0 FrameData_O[13]
rlabel metal2 41136 4368 41136 4368 0 FrameData_O[14]
rlabel metal2 41472 4956 41472 4956 0 FrameData_O[15]
rlabel metal2 41088 5124 41088 5124 0 FrameData_O[16]
rlabel metal3 42210 5796 42210 5796 0 FrameData_O[17]
rlabel metal2 41088 6006 41088 6006 0 FrameData_O[18]
rlabel metal2 41088 6384 41088 6384 0 FrameData_O[19]
rlabel metal2 40224 1050 40224 1050 0 FrameData_O[1]
rlabel metal2 41472 6720 41472 6720 0 FrameData_O[20]
rlabel metal2 41088 7056 41088 7056 0 FrameData_O[21]
rlabel metal2 41472 7434 41472 7434 0 FrameData_O[22]
rlabel metal3 42018 7812 42018 7812 0 FrameData_O[23]
rlabel metal3 41826 8148 41826 8148 0 FrameData_O[24]
rlabel metal3 42018 8484 42018 8484 0 FrameData_O[25]
rlabel metal2 40704 8862 40704 8862 0 FrameData_O[26]
rlabel metal2 41472 8946 41472 8946 0 FrameData_O[27]
rlabel metal2 41088 9408 41088 9408 0 FrameData_O[28]
rlabel metal2 40320 9324 40320 9324 0 FrameData_O[29]
rlabel metal2 41472 840 41472 840 0 FrameData_O[2]
rlabel metal2 41520 8148 41520 8148 0 FrameData_O[30]
rlabel metal2 41472 10080 41472 10080 0 FrameData_O[31]
rlabel metal2 40704 1008 40704 1008 0 FrameData_O[3]
rlabel metal2 39840 1554 39840 1554 0 FrameData_O[4]
rlabel metal3 42210 1764 42210 1764 0 FrameData_O[5]
rlabel metal3 42018 2100 42018 2100 0 FrameData_O[6]
rlabel metal3 42210 2436 42210 2436 0 FrameData_O[7]
rlabel metal3 41826 2772 41826 2772 0 FrameData_O[8]
rlabel metal2 41088 2982 41088 2982 0 FrameData_O[9]
rlabel metal2 3168 2058 3168 2058 0 FrameStrobe[0]
rlabel metal2 33312 882 33312 882 0 FrameStrobe[10]
rlabel metal2 31776 618 31776 618 0 FrameStrobe[11]
rlabel metal2 32928 366 32928 366 0 FrameStrobe[12]
rlabel metal2 34080 324 34080 324 0 FrameStrobe[13]
rlabel via2 35232 72 35232 72 0 FrameStrobe[14]
rlabel metal2 36384 618 36384 618 0 FrameStrobe[15]
rlabel via2 37536 72 37536 72 0 FrameStrobe[16]
rlabel metal2 38688 954 38688 954 0 FrameStrobe[17]
rlabel via2 39840 72 39840 72 0 FrameStrobe[18]
rlabel via2 40992 72 40992 72 0 FrameStrobe[19]
rlabel metal2 29184 1764 29184 1764 0 FrameStrobe[1]
rlabel metal2 38400 3192 38400 3192 0 FrameStrobe[2]
rlabel metal2 16704 1848 16704 1848 0 FrameStrobe[3]
rlabel metal2 31392 1764 31392 1764 0 FrameStrobe[4]
rlabel metal2 31584 1176 31584 1176 0 FrameStrobe[5]
rlabel metal2 26016 492 26016 492 0 FrameStrobe[6]
rlabel metal2 32544 924 32544 924 0 FrameStrobe[7]
rlabel metal2 31776 2982 31776 2982 0 FrameStrobe[8]
rlabel metal2 32832 966 32832 966 0 FrameStrobe[9]
rlabel metal2 29856 10176 29856 10176 0 FrameStrobe_O[0]
rlabel metal2 33072 1260 33072 1260 0 FrameStrobe_O[10]
rlabel metal3 32928 1260 32928 1260 0 FrameStrobe_O[11]
rlabel metal2 34224 840 34224 840 0 FrameStrobe_O[12]
rlabel metal3 32304 840 32304 840 0 FrameStrobe_O[13]
rlabel metal2 32544 9840 32544 9840 0 FrameStrobe_O[14]
rlabel metal2 37248 1890 37248 1890 0 FrameStrobe_O[15]
rlabel metal2 37632 1344 37632 1344 0 FrameStrobe_O[16]
rlabel metal3 33168 8736 33168 8736 0 FrameStrobe_O[17]
rlabel metal2 39264 3612 39264 3612 0 FrameStrobe_O[18]
rlabel metal2 40512 2100 40512 2100 0 FrameStrobe_O[19]
rlabel metal2 30048 10176 30048 10176 0 FrameStrobe_O[1]
rlabel metal2 30336 9660 30336 9660 0 FrameStrobe_O[2]
rlabel metal2 30816 9828 30816 9828 0 FrameStrobe_O[3]
rlabel metal2 30624 10134 30624 10134 0 FrameStrobe_O[4]
rlabel metal2 31584 2226 31584 2226 0 FrameStrobe_O[5]
rlabel metal3 31248 9660 31248 9660 0 FrameStrobe_O[6]
rlabel metal3 31920 924 31920 924 0 FrameStrobe_O[7]
rlabel metal2 31584 3696 31584 3696 0 FrameStrobe_O[8]
rlabel metal2 32736 1848 32736 1848 0 FrameStrobe_O[9]
rlabel metal2 36000 3780 36000 3780 0 Inst_A_IO_1_bidirectional_frame_config_pass.Q
rlabel metal2 19488 4326 19488 4326 0 Inst_B_IO_1_bidirectional_frame_config_pass.Q
rlabel metal2 7968 3108 7968 3108 0 Inst_S_IO_ConfigMem.Inst_frame0_bit0.Q
rlabel metal2 6816 2100 6816 2100 0 Inst_S_IO_ConfigMem.Inst_frame0_bit1.Q
rlabel metal2 35040 2856 35040 2856 0 Inst_S_IO_ConfigMem.Inst_frame0_bit10.Q
rlabel metal3 36768 2856 36768 2856 0 Inst_S_IO_ConfigMem.Inst_frame0_bit11.Q
rlabel metal3 31824 4368 31824 4368 0 Inst_S_IO_ConfigMem.Inst_frame0_bit12.Q
rlabel metal2 33504 5418 33504 5418 0 Inst_S_IO_ConfigMem.Inst_frame0_bit13.Q
rlabel metal2 19200 7392 19200 7392 0 Inst_S_IO_ConfigMem.Inst_frame0_bit14.Q
rlabel metal2 17520 7392 17520 7392 0 Inst_S_IO_ConfigMem.Inst_frame0_bit15.Q
rlabel metal2 19680 5124 19680 5124 0 Inst_S_IO_ConfigMem.Inst_frame0_bit16.Q
rlabel metal2 18048 5586 18048 5586 0 Inst_S_IO_ConfigMem.Inst_frame0_bit17.Q
rlabel metal2 4416 4872 4416 4872 0 Inst_S_IO_ConfigMem.Inst_frame0_bit18.Q
rlabel metal3 3888 4956 3888 4956 0 Inst_S_IO_ConfigMem.Inst_frame0_bit19.Q
rlabel metal2 19872 1934 19872 1934 0 Inst_S_IO_ConfigMem.Inst_frame0_bit2.Q
rlabel metal2 5664 3780 5664 3780 0 Inst_S_IO_ConfigMem.Inst_frame0_bit20.Q
rlabel metal3 3648 3444 3648 3444 0 Inst_S_IO_ConfigMem.Inst_frame0_bit21.Q
rlabel metal2 4704 1050 4704 1050 0 Inst_S_IO_ConfigMem.Inst_frame0_bit22.Q
rlabel metal2 3840 1806 3840 1806 0 Inst_S_IO_ConfigMem.Inst_frame0_bit23.Q
rlabel metal2 5088 1974 5088 1974 0 Inst_S_IO_ConfigMem.Inst_frame0_bit24.Q
rlabel metal2 6048 9408 6048 9408 0 Inst_S_IO_ConfigMem.Inst_frame0_bit25.Q
rlabel metal2 3504 8484 3504 8484 0 Inst_S_IO_ConfigMem.Inst_frame0_bit26.Q
rlabel metal2 4512 9450 4512 9450 0 Inst_S_IO_ConfigMem.Inst_frame0_bit27.Q
rlabel metal2 5472 9072 5472 9072 0 Inst_S_IO_ConfigMem.Inst_frame0_bit28.Q
rlabel metal2 5664 5082 5664 5082 0 Inst_S_IO_ConfigMem.Inst_frame0_bit29.Q
rlabel metal2 20064 2646 20064 2646 0 Inst_S_IO_ConfigMem.Inst_frame0_bit3.Q
rlabel metal3 5376 5628 5376 5628 0 Inst_S_IO_ConfigMem.Inst_frame0_bit30.Q
rlabel metal3 6288 6468 6288 6468 0 Inst_S_IO_ConfigMem.Inst_frame0_bit31.Q
rlabel metal2 34848 2268 34848 2268 0 Inst_S_IO_ConfigMem.Inst_frame0_bit4.Q
rlabel metal2 36984 3360 36984 3360 0 Inst_S_IO_ConfigMem.Inst_frame0_bit5.Q
rlabel metal2 19824 3612 19824 3612 0 Inst_S_IO_ConfigMem.Inst_frame0_bit6.Q
rlabel metal2 21456 3444 21456 3444 0 Inst_S_IO_ConfigMem.Inst_frame0_bit7.Q
rlabel metal2 16128 2562 16128 2562 0 Inst_S_IO_ConfigMem.Inst_frame0_bit8.Q
rlabel metal2 17736 2604 17736 2604 0 Inst_S_IO_ConfigMem.Inst_frame0_bit9.Q
rlabel metal2 13728 3654 13728 3654 0 Inst_S_IO_ConfigMem.Inst_frame1_bit0.Q
rlabel metal2 14496 1890 14496 1890 0 Inst_S_IO_ConfigMem.Inst_frame1_bit1.Q
rlabel metal2 30816 3990 30816 3990 0 Inst_S_IO_ConfigMem.Inst_frame1_bit10.Q
rlabel metal3 29088 4368 29088 4368 0 Inst_S_IO_ConfigMem.Inst_frame1_bit11.Q
rlabel metal2 25008 4179 25008 4179 0 Inst_S_IO_ConfigMem.Inst_frame1_bit12.Q
rlabel metal2 23472 2856 23472 2856 0 Inst_S_IO_ConfigMem.Inst_frame1_bit13.Q
rlabel metal2 29472 8316 29472 8316 0 Inst_S_IO_ConfigMem.Inst_frame1_bit14.Q
rlabel metal2 31152 8148 31152 8148 0 Inst_S_IO_ConfigMem.Inst_frame1_bit15.Q
rlabel metal3 24240 5796 24240 5796 0 Inst_S_IO_ConfigMem.Inst_frame1_bit16.Q
rlabel metal2 25536 6717 25536 6717 0 Inst_S_IO_ConfigMem.Inst_frame1_bit17.Q
rlabel metal2 21072 7392 21072 7392 0 Inst_S_IO_ConfigMem.Inst_frame1_bit18.Q
rlabel metal2 22848 7644 22848 7644 0 Inst_S_IO_ConfigMem.Inst_frame1_bit19.Q
rlabel metal2 28992 5082 28992 5082 0 Inst_S_IO_ConfigMem.Inst_frame1_bit2.Q
rlabel metal2 15408 3612 15408 3612 0 Inst_S_IO_ConfigMem.Inst_frame1_bit20.Q
rlabel metal2 16992 3866 16992 3866 0 Inst_S_IO_ConfigMem.Inst_frame1_bit21.Q
rlabel metal3 32784 2856 32784 2856 0 Inst_S_IO_ConfigMem.Inst_frame1_bit22.Q
rlabel metal2 34176 3567 34176 3567 0 Inst_S_IO_ConfigMem.Inst_frame1_bit23.Q
rlabel metal2 31488 6720 31488 6720 0 Inst_S_IO_ConfigMem.Inst_frame1_bit24.Q
rlabel metal2 33072 6405 33072 6405 0 Inst_S_IO_ConfigMem.Inst_frame1_bit25.Q
rlabel metal2 18720 8736 18720 8736 0 Inst_S_IO_ConfigMem.Inst_frame1_bit26.Q
rlabel metal2 20496 9240 20496 9240 0 Inst_S_IO_ConfigMem.Inst_frame1_bit27.Q
rlabel metal2 14784 8610 14784 8610 0 Inst_S_IO_ConfigMem.Inst_frame1_bit28.Q
rlabel metal2 16320 8953 16320 8953 0 Inst_S_IO_ConfigMem.Inst_frame1_bit29.Q
rlabel metal3 30768 3276 30768 3276 0 Inst_S_IO_ConfigMem.Inst_frame1_bit3.Q
rlabel metal2 15840 7434 15840 7434 0 Inst_S_IO_ConfigMem.Inst_frame1_bit30.Q
rlabel metal2 14592 8022 14592 8022 0 Inst_S_IO_ConfigMem.Inst_frame1_bit31.Q
rlabel metal2 25200 3780 25200 3780 0 Inst_S_IO_ConfigMem.Inst_frame1_bit4.Q
rlabel metal2 26880 1890 26880 1890 0 Inst_S_IO_ConfigMem.Inst_frame1_bit5.Q
rlabel metal2 31104 3150 31104 3150 0 Inst_S_IO_ConfigMem.Inst_frame1_bit6.Q
rlabel metal2 29328 2100 29328 2100 0 Inst_S_IO_ConfigMem.Inst_frame1_bit7.Q
rlabel metal2 27408 1680 27408 1680 0 Inst_S_IO_ConfigMem.Inst_frame1_bit8.Q
rlabel metal2 26016 2142 26016 2142 0 Inst_S_IO_ConfigMem.Inst_frame1_bit9.Q
rlabel metal2 21504 3948 21504 3948 0 Inst_S_IO_ConfigMem.Inst_frame2_bit0.Q
rlabel metal2 23136 1890 23136 1890 0 Inst_S_IO_ConfigMem.Inst_frame2_bit1.Q
rlabel metal2 37344 3864 37344 3864 0 Inst_S_IO_ConfigMem.Inst_frame2_bit10.Q
rlabel metal2 39456 4417 39456 4417 0 Inst_S_IO_ConfigMem.Inst_frame2_bit11.Q
rlabel metal2 10560 3486 10560 3486 0 Inst_S_IO_ConfigMem.Inst_frame2_bit12.Q
rlabel metal2 12480 3488 12480 3488 0 Inst_S_IO_ConfigMem.Inst_frame2_bit13.Q
rlabel metal2 25824 7770 25824 7770 0 Inst_S_IO_ConfigMem.Inst_frame2_bit14.Q
rlabel metal2 27552 7644 27552 7644 0 Inst_S_IO_ConfigMem.Inst_frame2_bit15.Q
rlabel metal2 21552 6468 21552 6468 0 Inst_S_IO_ConfigMem.Inst_frame2_bit16.Q
rlabel metal2 22752 5964 22752 5964 0 Inst_S_IO_ConfigMem.Inst_frame2_bit17.Q
rlabel metal2 35856 7392 35856 7392 0 Inst_S_IO_ConfigMem.Inst_frame2_bit18.Q
rlabel metal2 37728 7602 37728 7602 0 Inst_S_IO_ConfigMem.Inst_frame2_bit19.Q
rlabel metal2 36432 4032 36432 4032 0 Inst_S_IO_ConfigMem.Inst_frame2_bit2.Q
rlabel metal2 12480 6510 12480 6510 0 Inst_S_IO_ConfigMem.Inst_frame2_bit20.Q
rlabel metal2 13968 5040 13968 5040 0 Inst_S_IO_ConfigMem.Inst_frame2_bit21.Q
rlabel metal2 40368 5880 40368 5880 0 Inst_S_IO_ConfigMem.Inst_frame2_bit22.Q
rlabel metal3 38496 5040 38496 5040 0 Inst_S_IO_ConfigMem.Inst_frame2_bit23.Q
rlabel metal2 14688 6132 14688 6132 0 Inst_S_IO_ConfigMem.Inst_frame2_bit24.Q
rlabel metal2 14496 6174 14496 6174 0 Inst_S_IO_ConfigMem.Inst_frame2_bit25.Q
rlabel via1 37872 7975 37872 7975 0 Inst_S_IO_ConfigMem.Inst_frame2_bit26.Q
rlabel metal2 36288 7896 36288 7896 0 Inst_S_IO_ConfigMem.Inst_frame2_bit27.Q
rlabel metal2 11376 7455 11376 7455 0 Inst_S_IO_ConfigMem.Inst_frame2_bit28.Q
rlabel metal2 9792 7098 9792 7098 0 Inst_S_IO_ConfigMem.Inst_frame2_bit29.Q
rlabel metal3 38208 2856 38208 2856 0 Inst_S_IO_ConfigMem.Inst_frame2_bit3.Q
rlabel metal2 37632 8232 37632 8232 0 Inst_S_IO_ConfigMem.Inst_frame2_bit30.Q
rlabel metal2 40416 7476 40416 7476 0 Inst_S_IO_ConfigMem.Inst_frame2_bit31.Q
rlabel metal2 9600 1890 9600 1890 0 Inst_S_IO_ConfigMem.Inst_frame2_bit4.Q
rlabel metal2 11280 1260 11280 1260 0 Inst_S_IO_ConfigMem.Inst_frame2_bit5.Q
rlabel metal2 27360 3864 27360 3864 0 Inst_S_IO_ConfigMem.Inst_frame2_bit6.Q
rlabel metal2 28896 3896 28896 3896 0 Inst_S_IO_ConfigMem.Inst_frame2_bit7.Q
rlabel metal2 22752 2772 22752 2772 0 Inst_S_IO_ConfigMem.Inst_frame2_bit8.Q
rlabel metal2 24384 2730 24384 2730 0 Inst_S_IO_ConfigMem.Inst_frame2_bit9.Q
rlabel metal2 34368 5922 34368 5922 0 Inst_S_IO_ConfigMem.Inst_frame3_bit18.Q
rlabel metal2 35856 5124 35856 5124 0 Inst_S_IO_ConfigMem.Inst_frame3_bit19.Q
rlabel metal3 9312 4956 9312 4956 0 Inst_S_IO_ConfigMem.Inst_frame3_bit20.Q
rlabel metal2 11040 5079 11040 5079 0 Inst_S_IO_ConfigMem.Inst_frame3_bit21.Q
rlabel metal2 27216 5880 27216 5880 0 Inst_S_IO_ConfigMem.Inst_frame3_bit22.Q
rlabel metal2 28704 6717 28704 6717 0 Inst_S_IO_ConfigMem.Inst_frame3_bit23.Q
rlabel metal2 22464 8610 22464 8610 0 Inst_S_IO_ConfigMem.Inst_frame3_bit24.Q
rlabel metal2 24144 9240 24144 9240 0 Inst_S_IO_ConfigMem.Inst_frame3_bit25.Q
rlabel metal2 32352 8946 32352 8946 0 Inst_S_IO_ConfigMem.Inst_frame3_bit26.Q
rlabel metal2 33888 8701 33888 8701 0 Inst_S_IO_ConfigMem.Inst_frame3_bit27.Q
rlabel metal3 10608 8652 10608 8652 0 Inst_S_IO_ConfigMem.Inst_frame3_bit28.Q
rlabel metal2 12384 8953 12384 8953 0 Inst_S_IO_ConfigMem.Inst_frame3_bit29.Q
rlabel metal2 26016 8946 26016 8946 0 Inst_S_IO_ConfigMem.Inst_frame3_bit30.Q
rlabel metal2 27552 8743 27552 8743 0 Inst_S_IO_ConfigMem.Inst_frame3_bit31.Q
rlabel metal2 9888 9576 9888 9576 0 Inst_S_IO_switch_matrix.DEBUG_select_N1BEG0[0]
rlabel metal2 34800 8148 34800 8148 0 Inst_S_IO_switch_matrix.DEBUG_select_N1BEG1[0]
rlabel metal2 9216 6510 9216 6510 0 Inst_S_IO_switch_matrix.DEBUG_select_N1BEG2[0]
rlabel metal2 20640 5964 20640 5964 0 Inst_S_IO_switch_matrix.DEBUG_select_N1BEG3[0]
rlabel metal3 8832 8736 8832 8736 0 Inst_S_IO_switch_matrix.N1BEG0
rlabel metal4 33792 6846 33792 6846 0 Inst_S_IO_switch_matrix.N1BEG1
rlabel metal2 9408 7098 9408 7098 0 Inst_S_IO_switch_matrix.N1BEG2
rlabel metal2 10560 6090 10560 6090 0 Inst_S_IO_switch_matrix.N1BEG3
rlabel metal2 35952 6384 35952 6384 0 Inst_S_IO_switch_matrix.N2BEG0
rlabel metal2 11232 5418 11232 5418 0 Inst_S_IO_switch_matrix.N2BEG1
rlabel metal2 12192 4662 12192 4662 0 Inst_S_IO_switch_matrix.N2BEG2
rlabel metal2 10560 9702 10560 9702 0 Inst_S_IO_switch_matrix.N2BEG3
rlabel metal2 33840 7224 33840 7224 0 Inst_S_IO_switch_matrix.N2BEG4
rlabel metal3 12144 7896 12144 7896 0 Inst_S_IO_switch_matrix.N2BEG5
rlabel metal2 12096 7728 12096 7728 0 Inst_S_IO_switch_matrix.N2BEG6
rlabel metal2 12288 4956 12288 4956 0 Inst_S_IO_switch_matrix.N2BEG7
rlabel metal2 38112 5922 38112 5922 0 Inst_S_IO_switch_matrix.N2BEGb0
rlabel metal2 11568 3612 11568 3612 0 Inst_S_IO_switch_matrix.N2BEGb1
rlabel metal2 28848 5124 28848 5124 0 Inst_S_IO_switch_matrix.N2BEGb2
rlabel metal2 24480 3108 24480 3108 0 Inst_S_IO_switch_matrix.N2BEGb3
rlabel metal3 40176 4872 40176 4872 0 Inst_S_IO_switch_matrix.N2BEGb4
rlabel metal2 12672 4872 12672 4872 0 Inst_S_IO_switch_matrix.N2BEGb5
rlabel metal3 27840 8148 27840 8148 0 Inst_S_IO_switch_matrix.N2BEGb6
rlabel metal2 23328 7266 23328 7266 0 Inst_S_IO_switch_matrix.N2BEGb7
rlabel metal2 37296 9408 37296 9408 0 Inst_S_IO_switch_matrix.N4BEG0
rlabel metal2 14208 6930 14208 6930 0 Inst_S_IO_switch_matrix.N4BEG1
rlabel metal2 30912 7056 30912 7056 0 Inst_S_IO_switch_matrix.N4BEG10
rlabel metal2 27264 2940 27264 2940 0 Inst_S_IO_switch_matrix.N4BEG11
rlabel metal2 30912 5712 30912 5712 0 Inst_S_IO_switch_matrix.N4BEG12
rlabel metal2 24768 6384 24768 6384 0 Inst_S_IO_switch_matrix.N4BEG13
rlabel metal3 31200 7896 31200 7896 0 Inst_S_IO_switch_matrix.N4BEG14
rlabel metal3 25488 6636 25488 6636 0 Inst_S_IO_switch_matrix.N4BEG15
rlabel metal3 40224 6384 40224 6384 0 Inst_S_IO_switch_matrix.N4BEG2
rlabel metal2 14736 6636 14736 6636 0 Inst_S_IO_switch_matrix.N4BEG3
rlabel metal2 38016 8778 38016 8778 0 Inst_S_IO_switch_matrix.N4BEG4
rlabel metal3 12144 7224 12144 7224 0 Inst_S_IO_switch_matrix.N4BEG5
rlabel metal2 40032 8442 40032 8442 0 Inst_S_IO_switch_matrix.N4BEG6
rlabel metal2 14880 4452 14880 4452 0 Inst_S_IO_switch_matrix.N4BEG7
rlabel metal2 31584 8442 31584 8442 0 Inst_S_IO_switch_matrix.N4BEG8
rlabel metal2 25728 8190 25728 8190 0 Inst_S_IO_switch_matrix.N4BEG9
rlabel metal2 22752 8484 22752 8484 0 Inst_S_IO_switch_matrix.NN4BEG0
rlabel metal2 17040 4872 17040 4872 0 Inst_S_IO_switch_matrix.NN4BEG1
rlabel metal3 21360 4872 21360 4872 0 Inst_S_IO_switch_matrix.NN4BEG10
rlabel metal2 17856 2940 17856 2940 0 Inst_S_IO_switch_matrix.NN4BEG11
rlabel metal2 37056 4158 37056 4158 0 Inst_S_IO_switch_matrix.NN4BEG12
rlabel metal2 32448 7770 32448 7770 0 Inst_S_IO_switch_matrix.NN4BEG13
rlabel metal2 19296 8295 19296 8295 0 Inst_S_IO_switch_matrix.NN4BEG14
rlabel metal2 19680 5964 19680 5964 0 Inst_S_IO_switch_matrix.NN4BEG15
rlabel metal2 34368 3906 34368 3906 0 Inst_S_IO_switch_matrix.NN4BEG2
rlabel metal2 33168 6636 33168 6636 0 Inst_S_IO_switch_matrix.NN4BEG3
rlabel metal2 20256 8022 20256 8022 0 Inst_S_IO_switch_matrix.NN4BEG4
rlabel metal3 16704 9408 16704 9408 0 Inst_S_IO_switch_matrix.NN4BEG5
rlabel metal3 16608 7896 16608 7896 0 Inst_S_IO_switch_matrix.NN4BEG6
rlabel metal2 17280 4410 17280 4410 0 Inst_S_IO_switch_matrix.NN4BEG7
rlabel metal2 19680 2940 19680 2940 0 Inst_S_IO_switch_matrix.NN4BEG8
rlabel metal2 37104 3612 37104 3612 0 Inst_S_IO_switch_matrix.NN4BEG9
rlabel via2 9504 10680 9504 10680 0 N1BEG[0]
rlabel metal2 10176 9744 10176 9744 0 N1BEG[1]
rlabel metal2 9600 8694 9600 8694 0 N1BEG[2]
rlabel metal2 10368 6804 10368 6804 0 N1BEG[3]
rlabel metal4 35712 4368 35712 4368 0 N2BEG[0]
rlabel metal2 10944 6636 10944 6636 0 N2BEG[1]
rlabel metal2 11760 7392 11760 7392 0 N2BEG[2]
rlabel metal2 10800 9660 10800 9660 0 N2BEG[3]
rlabel metal4 29568 5124 29568 5124 0 N2BEG[4]
rlabel metal2 11520 8400 11520 8400 0 N2BEG[5]
rlabel metal2 11904 8316 11904 8316 0 N2BEG[6]
rlabel metal3 11952 4704 11952 4704 0 N2BEG[7]
rlabel metal2 11808 9756 11808 9756 0 N2BEGb[0]
rlabel metal2 11904 5922 11904 5922 0 N2BEGb[1]
rlabel metal2 12192 10176 12192 10176 0 N2BEGb[2]
rlabel metal2 12816 2856 12816 2856 0 N2BEGb[3]
rlabel metal2 12576 9756 12576 9756 0 N2BEGb[4]
rlabel metal2 12864 7014 12864 7014 0 N2BEGb[5]
rlabel metal2 12960 9924 12960 9924 0 N2BEGb[6]
rlabel metal2 13152 10428 13152 10428 0 N2BEGb[7]
rlabel metal2 13344 9882 13344 9882 0 N4BEG[0]
rlabel metal2 15264 10176 15264 10176 0 N4BEG[10]
rlabel metal2 15456 9756 15456 9756 0 N4BEG[11]
rlabel metal2 15648 9756 15648 9756 0 N4BEG[12]
rlabel metal2 15840 10386 15840 10386 0 N4BEG[13]
rlabel metal2 16032 9756 16032 9756 0 N4BEG[14]
rlabel metal2 16224 10260 16224 10260 0 N4BEG[15]
rlabel metal2 13728 8106 13728 8106 0 N4BEG[1]
rlabel metal4 40224 6258 40224 6258 0 N4BEG[2]
rlabel metal3 14064 9660 14064 9660 0 N4BEG[3]
rlabel metal2 14112 9756 14112 9756 0 N4BEG[4]
rlabel metal2 12960 8190 12960 8190 0 N4BEG[5]
rlabel metal4 39744 4788 39744 4788 0 N4BEG[6]
rlabel metal2 14688 5124 14688 5124 0 N4BEG[7]
rlabel metal2 14880 10134 14880 10134 0 N4BEG[8]
rlabel metal2 15072 9924 15072 9924 0 N4BEG[9]
rlabel metal2 16416 10176 16416 10176 0 NN4BEG[0]
rlabel metal2 18336 9210 18336 9210 0 NN4BEG[10]
rlabel metal2 17808 3612 17808 3612 0 NN4BEG[11]
rlabel metal2 18720 10596 18720 10596 0 NN4BEG[12]
rlabel metal2 18912 10512 18912 10512 0 NN4BEG[13]
rlabel metal2 19056 9660 19056 9660 0 NN4BEG[14]
rlabel metal2 19536 6636 19536 6636 0 NN4BEG[15]
rlabel metal2 16704 4788 16704 4788 0 NN4BEG[1]
rlabel metal2 16800 9756 16800 9756 0 NN4BEG[2]
rlabel metal2 16992 10596 16992 10596 0 NN4BEG[3]
rlabel metal2 20016 8148 20016 8148 0 NN4BEG[4]
rlabel metal2 17232 9660 17232 9660 0 NN4BEG[5]
rlabel metal2 17088 8694 17088 8694 0 NN4BEG[6]
rlabel metal2 17376 6804 17376 6804 0 NN4BEG[7]
rlabel metal2 17952 7152 17952 7152 0 NN4BEG[8]
rlabel metal2 18144 9756 18144 9756 0 NN4BEG[9]
rlabel metal2 19680 9588 19680 9588 0 S1END[0]
rlabel metal2 19008 6762 19008 6762 0 S1END[1]
rlabel metal2 20064 10554 20064 10554 0 S1END[2]
rlabel metal2 12576 6594 12576 6594 0 S1END[3]
rlabel metal2 17760 7224 17760 7224 0 S2END[0]
rlabel metal4 14880 8610 14880 8610 0 S2END[1]
rlabel metal3 4464 1596 4464 1596 0 S2END[2]
rlabel metal3 38112 4200 38112 4200 0 S2END[3]
rlabel metal2 19296 8610 19296 8610 0 S2END[4]
rlabel via2 15360 8232 15360 8232 0 S2END[5]
rlabel metal2 18912 9660 18912 9660 0 S2END[6]
rlabel metal4 15840 8400 15840 8400 0 S2END[7]
rlabel metal3 14400 7980 14400 7980 0 S2MID[0]
rlabel metal2 18144 5880 18144 5880 0 S2MID[1]
rlabel metal2 15168 8064 15168 8064 0 S2MID[2]
rlabel metal2 18624 5460 18624 5460 0 S2MID[3]
rlabel metal2 15072 7812 15072 7812 0 S2MID[4]
rlabel metal2 18528 5544 18528 5544 0 S2MID[5]
rlabel metal2 15648 7875 15648 7875 0 S2MID[6]
rlabel metal2 16896 4746 16896 4746 0 S2MID[7]
rlabel metal3 20064 4116 20064 4116 0 S4END[0]
rlabel metal2 16704 2898 16704 2898 0 S4END[10]
rlabel metal3 38400 6510 38400 6510 0 S4END[11]
rlabel metal2 25920 5796 25920 5796 0 S4END[12]
rlabel metal2 29376 6636 29376 6636 0 S4END[13]
rlabel metal2 12960 6846 12960 6846 0 S4END[14]
rlabel metal3 32544 8442 32544 8442 0 S4END[15]
rlabel metal2 32736 3486 32736 3486 0 S4END[1]
rlabel metal2 21504 7854 21504 7854 0 S4END[2]
rlabel metal2 38400 4662 38400 4662 0 S4END[3]
rlabel metal3 23616 8736 23616 8736 0 S4END[4]
rlabel metal2 29760 4830 29760 4830 0 S4END[5]
rlabel metal2 15552 3948 15552 3948 0 S4END[6]
rlabel metal2 31584 6636 31584 6636 0 S4END[7]
rlabel metal2 16608 2982 16608 2982 0 S4END[8]
rlabel metal2 29280 6930 29280 6930 0 S4END[9]
rlabel metal3 25584 6468 25584 6468 0 SS4END[0]
rlabel metal2 15840 6342 15840 6342 0 SS4END[10]
rlabel metal2 38928 5208 38928 5208 0 SS4END[11]
rlabel metal2 23520 8064 23520 8064 0 SS4END[12]
rlabel metal2 29664 8946 29664 8946 0 SS4END[13]
rlabel metal2 15936 6846 15936 6846 0 SS4END[14]
rlabel metal2 38784 6678 38784 6678 0 SS4END[15]
rlabel metal2 26496 7980 26496 7980 0 SS4END[1]
rlabel metal2 11424 8757 11424 8757 0 SS4END[2]
rlabel metal2 38544 4200 38544 4200 0 SS4END[3]
rlabel metal2 23040 9114 23040 9114 0 SS4END[4]
rlabel metal2 27744 6594 27744 6594 0 SS4END[5]
rlabel metal2 10272 7266 10272 7266 0 SS4END[6]
rlabel metal2 36960 5586 36960 5586 0 SS4END[7]
rlabel metal2 22656 5712 22656 5712 0 SS4END[8]
rlabel metal2 29760 7056 29760 7056 0 SS4END[9]
rlabel metal2 17952 576 17952 576 0 UserCLK
rlabel metal3 26688 3444 26688 3444 0 UserCLK_regs
rlabel metal2 29664 1302 29664 1302 0 UserCLKo
rlabel metal2 4656 5880 4656 5880 0 _000_
rlabel metal2 3648 2604 3648 2604 0 _001_
rlabel metal2 5053 9316 5053 9316 0 _002_
rlabel metal2 4752 9492 4752 9492 0 _003_
rlabel metal2 3600 7392 3600 7392 0 _004_
rlabel metal3 4944 7980 4944 7980 0 _005_
rlabel metal2 3936 8064 3936 8064 0 _006_
rlabel metal2 4080 7980 4080 7980 0 _007_
rlabel metal2 3840 8316 3840 8316 0 _008_
rlabel metal2 4416 8442 4416 8442 0 _009_
rlabel metal2 3744 9576 3744 9576 0 _010_
rlabel metal2 5376 9534 5376 9534 0 _011_
rlabel metal2 5472 8232 5472 8232 0 _012_
rlabel metal2 7632 8148 7632 8148 0 _013_
rlabel metal3 7440 9492 7440 9492 0 _014_
rlabel metal2 5568 8736 5568 8736 0 _015_
rlabel metal2 5760 8358 5760 8358 0 _016_
rlabel via1 4685 3444 4685 3444 0 _017_
rlabel metal2 4368 3444 4368 3444 0 _018_
rlabel metal2 4224 4074 4224 4074 0 _019_
rlabel metal2 4608 3654 4608 3654 0 _020_
rlabel metal2 3744 4242 3744 4242 0 _021_
rlabel metal2 3840 3864 3840 3864 0 _022_
rlabel metal2 3648 3696 3648 3696 0 _023_
rlabel metal3 5184 4116 5184 4116 0 _024_
rlabel metal2 5280 3948 5280 3948 0 _025_
rlabel metal2 3744 3486 3744 3486 0 _026_
rlabel metal2 3936 3402 3936 3402 0 _027_
rlabel metal2 7104 3612 7104 3612 0 _028_
rlabel metal2 7008 3738 7008 3738 0 _029_
rlabel metal2 3744 4914 3744 4914 0 _030_
rlabel metal2 6144 4410 6144 4410 0 _031_
rlabel metal2 5328 2604 5328 2604 0 _032_
rlabel metal3 4656 1932 4656 1932 0 _033_
rlabel metal2 4032 2184 4032 2184 0 _034_
rlabel metal3 4464 1092 4464 1092 0 _035_
rlabel metal2 4512 2226 4512 2226 0 _036_
rlabel metal2 4224 1680 4224 1680 0 _037_
rlabel metal2 4704 1848 4704 1848 0 _038_
rlabel metal2 4896 1386 4896 1386 0 _039_
rlabel metal2 7104 5964 7104 5964 0 _040_
rlabel metal2 6624 6510 6624 6510 0 _041_
rlabel metal3 6096 5040 6096 5040 0 _042_
rlabel metal2 7296 6888 7296 6888 0 _043_
rlabel metal3 6480 6972 6480 6972 0 _044_
rlabel metal2 34080 1302 34080 1302 0 _045_
rlabel metal3 17760 1260 17760 1260 0 _046_
rlabel metal3 30912 1260 30912 1260 0 clknet_0_UserCLK
rlabel metal2 29952 2268 29952 2268 0 clknet_0_UserCLK_regs
rlabel metal2 29472 2730 29472 2730 0 clknet_1_0__leaf_UserCLK
rlabel metal2 18432 2268 18432 2268 0 clknet_1_0__leaf_UserCLK_regs
rlabel metal2 30912 1512 30912 1512 0 clknet_1_1__leaf_UserCLK_regs
<< properties >>
string FIXED_BBOX 0 0 43008 10752
<< end >>
