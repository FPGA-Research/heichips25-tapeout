magic
tech ihp-sg13g2
magscale 1 2
timestamp 1752758680
<< metal1 >>
rect 1152 41600 20452 41624
rect 1152 41560 4928 41600
rect 4968 41560 5010 41600
rect 5050 41560 5092 41600
rect 5132 41560 5174 41600
rect 5214 41560 5256 41600
rect 5296 41560 20048 41600
rect 20088 41560 20130 41600
rect 20170 41560 20212 41600
rect 20252 41560 20294 41600
rect 20334 41560 20376 41600
rect 20416 41560 20452 41600
rect 1152 41536 20452 41560
rect 8235 41432 8277 41441
rect 8235 41392 8236 41432
rect 8276 41392 8277 41432
rect 8235 41383 8277 41392
rect 18603 41432 18645 41441
rect 18603 41392 18604 41432
rect 18644 41392 18645 41432
rect 18603 41383 18645 41392
rect 18987 41432 19029 41441
rect 18987 41392 18988 41432
rect 19028 41392 19029 41432
rect 18987 41383 19029 41392
rect 19371 41432 19413 41441
rect 19371 41392 19372 41432
rect 19412 41392 19413 41432
rect 19371 41383 19413 41392
rect 1795 41264 1853 41265
rect 1795 41224 1804 41264
rect 1844 41224 1853 41264
rect 1795 41223 1853 41224
rect 3043 41264 3101 41265
rect 3043 41224 3052 41264
rect 3092 41224 3101 41264
rect 3043 41223 3101 41224
rect 3427 41264 3485 41265
rect 3427 41224 3436 41264
rect 3476 41224 3485 41264
rect 3427 41223 3485 41224
rect 4675 41264 4733 41265
rect 4675 41224 4684 41264
rect 4724 41224 4733 41264
rect 4675 41223 4733 41224
rect 6307 41264 6365 41265
rect 6307 41224 6316 41264
rect 6356 41224 6365 41264
rect 6307 41223 6365 41224
rect 7555 41264 7613 41265
rect 7555 41224 7564 41264
rect 7604 41224 7613 41264
rect 7555 41223 7613 41224
rect 8707 41264 8765 41265
rect 8707 41224 8716 41264
rect 8756 41224 8765 41264
rect 8707 41223 8765 41224
rect 9955 41264 10013 41265
rect 9955 41224 9964 41264
rect 10004 41224 10013 41264
rect 9955 41223 10013 41224
rect 10339 41264 10397 41265
rect 10339 41224 10348 41264
rect 10388 41224 10397 41264
rect 10339 41223 10397 41224
rect 11587 41264 11645 41265
rect 11587 41224 11596 41264
rect 11636 41224 11645 41264
rect 11587 41223 11645 41224
rect 12163 41264 12221 41265
rect 12163 41224 12172 41264
rect 12212 41224 12221 41264
rect 12163 41223 12221 41224
rect 13411 41264 13469 41265
rect 13411 41224 13420 41264
rect 13460 41224 13469 41264
rect 13411 41223 13469 41224
rect 13795 41264 13853 41265
rect 13795 41224 13804 41264
rect 13844 41224 13853 41264
rect 13795 41223 13853 41224
rect 15043 41264 15101 41265
rect 15043 41224 15052 41264
rect 15092 41224 15101 41264
rect 15043 41223 15101 41224
rect 16675 41264 16733 41265
rect 16675 41224 16684 41264
rect 16724 41224 16733 41264
rect 16675 41223 16733 41224
rect 17923 41264 17981 41265
rect 17923 41224 17932 41264
rect 17972 41224 17981 41264
rect 17923 41223 17981 41224
rect 8035 41180 8093 41181
rect 8035 41140 8044 41180
rect 8084 41140 8093 41180
rect 8035 41139 8093 41140
rect 15427 41180 15485 41181
rect 15427 41140 15436 41180
rect 15476 41140 15485 41180
rect 15427 41139 15485 41140
rect 15811 41180 15869 41181
rect 15811 41140 15820 41180
rect 15860 41140 15869 41180
rect 15811 41139 15869 41140
rect 16195 41180 16253 41181
rect 16195 41140 16204 41180
rect 16244 41140 16253 41180
rect 16195 41139 16253 41140
rect 18787 41180 18845 41181
rect 18787 41140 18796 41180
rect 18836 41140 18845 41180
rect 18787 41139 18845 41140
rect 19171 41180 19229 41181
rect 19171 41140 19180 41180
rect 19220 41140 19229 41180
rect 19171 41139 19229 41140
rect 19555 41180 19613 41181
rect 19555 41140 19564 41180
rect 19604 41140 19613 41180
rect 19555 41139 19613 41140
rect 19747 41180 19805 41181
rect 19747 41140 19756 41180
rect 19796 41140 19805 41180
rect 19747 41139 19805 41140
rect 1323 41096 1365 41105
rect 1323 41056 1324 41096
rect 1364 41056 1365 41096
rect 1323 41047 1365 41056
rect 18315 41096 18357 41105
rect 18315 41056 18316 41096
rect 18356 41056 18357 41096
rect 18315 41047 18357 41056
rect 3243 41012 3285 41021
rect 3243 40972 3244 41012
rect 3284 40972 3285 41012
rect 3243 40963 3285 40972
rect 4875 41012 4917 41021
rect 4875 40972 4876 41012
rect 4916 40972 4917 41012
rect 4875 40963 4917 40972
rect 6123 41012 6165 41021
rect 6123 40972 6124 41012
rect 6164 40972 6165 41012
rect 6123 40963 6165 40972
rect 10155 41012 10197 41021
rect 10155 40972 10156 41012
rect 10196 40972 10197 41012
rect 10155 40963 10197 40972
rect 11787 41012 11829 41021
rect 11787 40972 11788 41012
rect 11828 40972 11829 41012
rect 11787 40963 11829 40972
rect 11979 41012 12021 41021
rect 11979 40972 11980 41012
rect 12020 40972 12021 41012
rect 11979 40963 12021 40972
rect 13611 41012 13653 41021
rect 13611 40972 13612 41012
rect 13652 40972 13653 41012
rect 13611 40963 13653 40972
rect 15243 41012 15285 41021
rect 15243 40972 15244 41012
rect 15284 40972 15285 41012
rect 15243 40963 15285 40972
rect 15627 41012 15669 41021
rect 15627 40972 15628 41012
rect 15668 40972 15669 41012
rect 15627 40963 15669 40972
rect 16011 41012 16053 41021
rect 16011 40972 16012 41012
rect 16052 40972 16053 41012
rect 16011 40963 16053 40972
rect 18123 41012 18165 41021
rect 18123 40972 18124 41012
rect 18164 40972 18165 41012
rect 18123 40963 18165 40972
rect 19947 41012 19989 41021
rect 19947 40972 19948 41012
rect 19988 40972 19989 41012
rect 19947 40963 19989 40972
rect 1152 40844 20352 40868
rect 1152 40804 3688 40844
rect 3728 40804 3770 40844
rect 3810 40804 3852 40844
rect 3892 40804 3934 40844
rect 3974 40804 4016 40844
rect 4056 40804 18808 40844
rect 18848 40804 18890 40844
rect 18930 40804 18972 40844
rect 19012 40804 19054 40844
rect 19094 40804 19136 40844
rect 19176 40804 20352 40844
rect 1152 40780 20352 40804
rect 1707 40676 1749 40685
rect 1707 40636 1708 40676
rect 1748 40636 1749 40676
rect 1707 40627 1749 40636
rect 3915 40676 3957 40685
rect 3915 40636 3916 40676
rect 3956 40636 3957 40676
rect 3915 40627 3957 40636
rect 6219 40676 6261 40685
rect 6219 40636 6220 40676
rect 6260 40636 6261 40676
rect 6219 40627 6261 40636
rect 13707 40676 13749 40685
rect 13707 40636 13708 40676
rect 13748 40636 13749 40676
rect 13707 40627 13749 40636
rect 17451 40676 17493 40685
rect 17451 40636 17452 40676
rect 17492 40636 17493 40676
rect 17451 40627 17493 40636
rect 18315 40676 18357 40685
rect 18315 40636 18316 40676
rect 18356 40636 18357 40676
rect 18315 40627 18357 40636
rect 19083 40676 19125 40685
rect 19083 40636 19084 40676
rect 19124 40636 19125 40676
rect 19083 40627 19125 40636
rect 19467 40676 19509 40685
rect 19467 40636 19468 40676
rect 19508 40636 19509 40676
rect 19467 40627 19509 40636
rect 19851 40676 19893 40685
rect 19851 40636 19852 40676
rect 19892 40636 19893 40676
rect 19851 40627 19893 40636
rect 1323 40592 1365 40601
rect 1323 40552 1324 40592
rect 1364 40552 1365 40592
rect 1323 40543 1365 40552
rect 3531 40592 3573 40601
rect 3531 40552 3532 40592
rect 3572 40552 3573 40592
rect 3531 40543 3573 40552
rect 14091 40592 14133 40601
rect 14091 40552 14092 40592
rect 14132 40552 14133 40592
rect 14091 40543 14133 40552
rect 14475 40592 14517 40601
rect 14475 40552 14476 40592
rect 14516 40552 14517 40592
rect 14475 40543 14517 40552
rect 14859 40592 14901 40601
rect 14859 40552 14860 40592
rect 14900 40552 14901 40592
rect 14859 40543 14901 40552
rect 15243 40592 15285 40601
rect 15243 40552 15244 40592
rect 15284 40552 15285 40592
rect 15243 40543 15285 40552
rect 15627 40592 15669 40601
rect 15627 40552 15628 40592
rect 15668 40552 15669 40592
rect 15627 40543 15669 40552
rect 16011 40592 16053 40601
rect 16011 40552 16012 40592
rect 16052 40552 16053 40592
rect 16011 40543 16053 40552
rect 16395 40592 16437 40601
rect 16395 40552 16396 40592
rect 16436 40552 16437 40592
rect 16395 40543 16437 40552
rect 17643 40592 17685 40601
rect 17643 40552 17644 40592
rect 17684 40552 17685 40592
rect 17643 40543 17685 40552
rect 18699 40592 18741 40601
rect 18699 40552 18700 40592
rect 18740 40552 18741 40592
rect 18699 40543 18741 40552
rect 16579 40519 16637 40520
rect 1507 40508 1565 40509
rect 1507 40468 1516 40508
rect 1556 40468 1565 40508
rect 1507 40467 1565 40468
rect 3715 40508 3773 40509
rect 3715 40468 3724 40508
rect 3764 40468 3773 40508
rect 3715 40467 3773 40468
rect 6019 40508 6077 40509
rect 6019 40468 6028 40508
rect 6068 40468 6077 40508
rect 13891 40508 13949 40509
rect 6019 40467 6077 40468
rect 11739 40466 11781 40475
rect 13891 40468 13900 40508
rect 13940 40468 13949 40508
rect 13891 40467 13949 40468
rect 14275 40508 14333 40509
rect 14275 40468 14284 40508
rect 14324 40468 14333 40508
rect 14275 40467 14333 40468
rect 14659 40508 14717 40509
rect 14659 40468 14668 40508
rect 14708 40468 14717 40508
rect 14659 40467 14717 40468
rect 15043 40508 15101 40509
rect 15043 40468 15052 40508
rect 15092 40468 15101 40508
rect 15043 40467 15101 40468
rect 15427 40508 15485 40509
rect 15427 40468 15436 40508
rect 15476 40468 15485 40508
rect 15427 40467 15485 40468
rect 15811 40508 15869 40509
rect 15811 40468 15820 40508
rect 15860 40468 15869 40508
rect 15811 40467 15869 40468
rect 16195 40508 16253 40509
rect 16195 40468 16204 40508
rect 16244 40468 16253 40508
rect 16579 40479 16588 40519
rect 16628 40479 16637 40519
rect 16579 40478 16637 40479
rect 16963 40508 17021 40509
rect 16195 40467 16253 40468
rect 16963 40468 16972 40508
rect 17012 40468 17021 40508
rect 16963 40467 17021 40468
rect 17251 40508 17309 40509
rect 17251 40468 17260 40508
rect 17300 40468 17309 40508
rect 17251 40467 17309 40468
rect 17827 40508 17885 40509
rect 17827 40468 17836 40508
rect 17876 40468 17885 40508
rect 17827 40467 17885 40468
rect 18027 40508 18069 40517
rect 18027 40468 18028 40508
rect 18068 40468 18069 40508
rect 2083 40424 2141 40425
rect 2083 40384 2092 40424
rect 2132 40384 2141 40424
rect 2083 40383 2141 40384
rect 3331 40424 3389 40425
rect 3331 40384 3340 40424
rect 3380 40384 3389 40424
rect 3331 40383 3389 40384
rect 4099 40424 4157 40425
rect 4099 40384 4108 40424
rect 4148 40384 4157 40424
rect 4099 40383 4157 40384
rect 5347 40424 5405 40425
rect 5347 40384 5356 40424
rect 5396 40384 5405 40424
rect 5347 40383 5405 40384
rect 6403 40424 6461 40425
rect 6403 40384 6412 40424
rect 6452 40384 6461 40424
rect 6403 40383 6461 40384
rect 7651 40424 7709 40425
rect 7651 40384 7660 40424
rect 7700 40384 7709 40424
rect 7651 40383 7709 40384
rect 8131 40424 8189 40425
rect 8131 40384 8140 40424
rect 8180 40384 8189 40424
rect 8131 40383 8189 40384
rect 9379 40424 9437 40425
rect 9379 40384 9388 40424
rect 9428 40384 9437 40424
rect 9379 40383 9437 40384
rect 10155 40424 10197 40433
rect 10155 40384 10156 40424
rect 10196 40384 10197 40424
rect 10155 40375 10197 40384
rect 10251 40424 10293 40433
rect 10251 40384 10252 40424
rect 10292 40384 10293 40424
rect 10251 40375 10293 40384
rect 10635 40424 10677 40433
rect 10635 40384 10636 40424
rect 10676 40384 10677 40424
rect 10635 40375 10677 40384
rect 10731 40424 10773 40433
rect 11739 40426 11740 40466
rect 11780 40426 11781 40466
rect 18027 40459 18069 40468
rect 18499 40508 18557 40509
rect 18499 40468 18508 40508
rect 18548 40468 18557 40508
rect 18499 40467 18557 40468
rect 18883 40508 18941 40509
rect 18883 40468 18892 40508
rect 18932 40468 18941 40508
rect 18883 40467 18941 40468
rect 19267 40508 19325 40509
rect 19267 40468 19276 40508
rect 19316 40468 19325 40508
rect 19267 40467 19325 40468
rect 19651 40508 19709 40509
rect 19651 40468 19660 40508
rect 19700 40468 19709 40508
rect 19651 40467 19709 40468
rect 20035 40508 20093 40509
rect 20035 40468 20044 40508
rect 20084 40468 20093 40508
rect 20035 40467 20093 40468
rect 10731 40384 10732 40424
rect 10772 40384 10773 40424
rect 10731 40375 10773 40384
rect 11203 40424 11261 40425
rect 11203 40384 11212 40424
rect 11252 40384 11261 40424
rect 11739 40417 11781 40426
rect 12259 40424 12317 40425
rect 11203 40383 11261 40384
rect 12259 40384 12268 40424
rect 12308 40384 12317 40424
rect 12259 40383 12317 40384
rect 13507 40424 13565 40425
rect 13507 40384 13516 40424
rect 13556 40384 13565 40424
rect 13507 40383 13565 40384
rect 5547 40340 5589 40349
rect 5547 40300 5548 40340
rect 5588 40300 5589 40340
rect 5547 40291 5589 40300
rect 9771 40340 9813 40349
rect 9771 40300 9772 40340
rect 9812 40300 9813 40340
rect 9771 40291 9813 40300
rect 7851 40256 7893 40265
rect 7851 40216 7852 40256
rect 7892 40216 7893 40256
rect 7851 40207 7893 40216
rect 9579 40256 9621 40265
rect 9579 40216 9580 40256
rect 9620 40216 9621 40256
rect 12075 40256 12117 40265
rect 9579 40207 9621 40216
rect 11883 40214 11925 40223
rect 11883 40174 11884 40214
rect 11924 40174 11925 40214
rect 12075 40216 12076 40256
rect 12116 40216 12117 40256
rect 12075 40207 12117 40216
rect 16779 40256 16821 40265
rect 16779 40216 16780 40256
rect 16820 40216 16821 40256
rect 16779 40207 16821 40216
rect 11883 40165 11925 40174
rect 1152 40088 20452 40112
rect 1152 40048 4928 40088
rect 4968 40048 5010 40088
rect 5050 40048 5092 40088
rect 5132 40048 5174 40088
rect 5214 40048 5256 40088
rect 5296 40048 20048 40088
rect 20088 40048 20130 40088
rect 20170 40048 20212 40088
rect 20252 40048 20294 40088
rect 20334 40048 20376 40088
rect 20416 40048 20452 40088
rect 1152 40024 20452 40048
rect 1419 39920 1461 39929
rect 1419 39880 1420 39920
rect 1460 39880 1461 39920
rect 1419 39871 1461 39880
rect 3531 39920 3573 39929
rect 3531 39880 3532 39920
rect 3572 39880 3573 39920
rect 3531 39871 3573 39880
rect 10251 39920 10293 39929
rect 10251 39880 10252 39920
rect 10292 39880 10293 39920
rect 10251 39871 10293 39880
rect 13131 39920 13173 39929
rect 13131 39880 13132 39920
rect 13172 39880 13173 39920
rect 13131 39871 13173 39880
rect 17547 39920 17589 39929
rect 17547 39880 17548 39920
rect 17588 39880 17589 39920
rect 17547 39871 17589 39880
rect 18411 39920 18453 39929
rect 18411 39880 18412 39920
rect 18452 39880 18453 39920
rect 18411 39871 18453 39880
rect 18603 39920 18645 39929
rect 18603 39880 18604 39920
rect 18644 39880 18645 39920
rect 18603 39871 18645 39880
rect 18987 39920 19029 39929
rect 18987 39880 18988 39920
rect 19028 39880 19029 39920
rect 18987 39871 19029 39880
rect 12747 39836 12789 39845
rect 12747 39796 12748 39836
rect 12788 39796 12789 39836
rect 12747 39787 12789 39796
rect 1699 39752 1757 39753
rect 1699 39712 1708 39752
rect 1748 39712 1757 39752
rect 1699 39711 1757 39712
rect 2947 39752 3005 39753
rect 2947 39712 2956 39752
rect 2996 39712 3005 39752
rect 2947 39711 3005 39712
rect 4387 39752 4445 39753
rect 4387 39712 4396 39752
rect 4436 39712 4445 39752
rect 4387 39711 4445 39712
rect 5635 39752 5693 39753
rect 5635 39712 5644 39752
rect 5684 39712 5693 39752
rect 5635 39711 5693 39712
rect 6979 39752 7037 39753
rect 6979 39712 6988 39752
rect 7028 39712 7037 39752
rect 6979 39711 7037 39712
rect 8227 39752 8285 39753
rect 8227 39712 8236 39752
rect 8276 39712 8285 39752
rect 8227 39711 8285 39712
rect 8611 39752 8669 39753
rect 8611 39712 8620 39752
rect 8660 39712 8669 39752
rect 8611 39711 8669 39712
rect 9859 39752 9917 39753
rect 9859 39712 9868 39752
rect 9908 39712 9917 39752
rect 9859 39711 9917 39712
rect 11019 39752 11061 39761
rect 11019 39712 11020 39752
rect 11060 39712 11061 39752
rect 11019 39703 11061 39712
rect 11115 39752 11157 39761
rect 11115 39712 11116 39752
rect 11156 39712 11157 39752
rect 11115 39703 11157 39712
rect 12067 39752 12125 39753
rect 12067 39712 12076 39752
rect 12116 39712 12125 39752
rect 12067 39711 12125 39712
rect 12555 39747 12597 39756
rect 12555 39707 12556 39747
rect 12596 39707 12597 39747
rect 13315 39752 13373 39753
rect 13315 39712 13324 39752
rect 13364 39712 13373 39752
rect 13315 39711 13373 39712
rect 14563 39752 14621 39753
rect 14563 39712 14572 39752
rect 14612 39712 14621 39752
rect 14563 39711 14621 39712
rect 15235 39752 15293 39753
rect 15235 39712 15244 39752
rect 15284 39712 15293 39752
rect 15235 39711 15293 39712
rect 16483 39752 16541 39753
rect 16483 39712 16492 39752
rect 16532 39712 16541 39752
rect 16483 39711 16541 39712
rect 12555 39698 12597 39707
rect 1219 39668 1277 39669
rect 1219 39628 1228 39668
rect 1268 39628 1277 39668
rect 1219 39627 1277 39628
rect 3331 39668 3389 39669
rect 3331 39628 3340 39668
rect 3380 39628 3389 39668
rect 3331 39627 3389 39628
rect 10435 39668 10493 39669
rect 10435 39628 10444 39668
rect 10484 39628 10493 39668
rect 10435 39627 10493 39628
rect 11499 39668 11541 39677
rect 11499 39628 11500 39668
rect 11540 39628 11541 39668
rect 11499 39619 11541 39628
rect 11595 39668 11637 39677
rect 11595 39628 11596 39668
rect 11636 39628 11637 39668
rect 11595 39619 11637 39628
rect 12931 39668 12989 39669
rect 12931 39628 12940 39668
rect 12980 39628 12989 39668
rect 12931 39627 12989 39628
rect 17059 39668 17117 39669
rect 17059 39628 17068 39668
rect 17108 39628 17117 39668
rect 17059 39627 17117 39628
rect 17731 39668 17789 39669
rect 17731 39628 17740 39668
rect 17780 39628 17789 39668
rect 17731 39627 17789 39628
rect 18211 39668 18269 39669
rect 18211 39628 18220 39668
rect 18260 39628 18269 39668
rect 18211 39627 18269 39628
rect 18787 39668 18845 39669
rect 18787 39628 18796 39668
rect 18836 39628 18845 39668
rect 18787 39627 18845 39628
rect 19171 39668 19229 39669
rect 19171 39628 19180 39668
rect 19220 39628 19229 39668
rect 19171 39627 19229 39628
rect 19363 39668 19421 39669
rect 19363 39628 19372 39668
rect 19412 39628 19421 39668
rect 19363 39627 19421 39628
rect 19747 39668 19805 39669
rect 19747 39628 19756 39668
rect 19796 39628 19805 39668
rect 19747 39627 19805 39628
rect 3819 39584 3861 39593
rect 3819 39544 3820 39584
rect 3860 39544 3861 39584
rect 3819 39535 3861 39544
rect 6027 39584 6069 39593
rect 6027 39544 6028 39584
rect 6068 39544 6069 39584
rect 6027 39535 6069 39544
rect 10635 39584 10677 39593
rect 10635 39544 10636 39584
rect 10676 39544 10677 39584
rect 10635 39535 10677 39544
rect 17259 39584 17301 39593
rect 17259 39544 17260 39584
rect 17300 39544 17301 39584
rect 17259 39535 17301 39544
rect 18027 39584 18069 39593
rect 18027 39544 18028 39584
rect 18068 39544 18069 39584
rect 18027 39535 18069 39544
rect 20139 39584 20181 39593
rect 20139 39544 20140 39584
rect 20180 39544 20181 39584
rect 20139 39535 20181 39544
rect 3147 39500 3189 39509
rect 3147 39460 3148 39500
rect 3188 39460 3189 39500
rect 3147 39451 3189 39460
rect 5835 39500 5877 39509
rect 5835 39460 5836 39500
rect 5876 39460 5877 39500
rect 5835 39451 5877 39460
rect 8427 39500 8469 39509
rect 8427 39460 8428 39500
rect 8468 39460 8469 39500
rect 8427 39451 8469 39460
rect 10059 39500 10101 39509
rect 10059 39460 10060 39500
rect 10100 39460 10101 39500
rect 10059 39451 10101 39460
rect 14763 39500 14805 39509
rect 14763 39460 14764 39500
rect 14804 39460 14805 39500
rect 14763 39451 14805 39460
rect 16683 39500 16725 39509
rect 16683 39460 16684 39500
rect 16724 39460 16725 39500
rect 16683 39451 16725 39460
rect 16875 39500 16917 39509
rect 16875 39460 16876 39500
rect 16916 39460 16917 39500
rect 16875 39451 16917 39460
rect 19563 39500 19605 39509
rect 19563 39460 19564 39500
rect 19604 39460 19605 39500
rect 19563 39451 19605 39460
rect 19947 39500 19989 39509
rect 19947 39460 19948 39500
rect 19988 39460 19989 39500
rect 19947 39451 19989 39460
rect 1152 39332 20352 39356
rect 1152 39292 3688 39332
rect 3728 39292 3770 39332
rect 3810 39292 3852 39332
rect 3892 39292 3934 39332
rect 3974 39292 4016 39332
rect 4056 39292 18808 39332
rect 18848 39292 18890 39332
rect 18930 39292 18972 39332
rect 19012 39292 19054 39332
rect 19094 39292 19136 39332
rect 19176 39292 20352 39332
rect 1152 39268 20352 39292
rect 17451 39164 17493 39173
rect 17451 39124 17452 39164
rect 17492 39124 17493 39164
rect 17451 39115 17493 39124
rect 1515 39080 1557 39089
rect 1515 39040 1516 39080
rect 1556 39040 1557 39080
rect 1515 39031 1557 39040
rect 4395 39080 4437 39089
rect 4395 39040 4396 39080
rect 4436 39040 4437 39080
rect 4395 39031 4437 39040
rect 14667 39080 14709 39089
rect 14667 39040 14668 39080
rect 14708 39040 14709 39080
rect 14667 39031 14709 39040
rect 17643 39080 17685 39089
rect 17643 39040 17644 39080
rect 17684 39040 17685 39080
rect 17643 39031 17685 39040
rect 18507 39080 18549 39089
rect 18507 39040 18508 39080
rect 18548 39040 18549 39080
rect 18507 39031 18549 39040
rect 1315 38996 1373 38997
rect 1315 38956 1324 38996
rect 1364 38956 1373 38996
rect 1315 38955 1373 38956
rect 4195 38996 4253 38997
rect 4195 38956 4204 38996
rect 4244 38956 4253 38996
rect 4195 38955 4253 38956
rect 6315 38996 6357 39005
rect 6315 38956 6316 38996
rect 6356 38956 6357 38996
rect 6315 38947 6357 38956
rect 8331 38996 8373 39005
rect 8331 38956 8332 38996
rect 8372 38956 8373 38996
rect 8331 38947 8373 38956
rect 12067 38996 12125 38997
rect 12067 38956 12076 38996
rect 12116 38956 12125 38996
rect 12067 38955 12125 38956
rect 14467 38996 14525 38997
rect 14467 38956 14476 38996
rect 14516 38956 14525 38996
rect 14467 38955 14525 38956
rect 15531 38996 15573 39005
rect 15531 38956 15532 38996
rect 15572 38956 15573 38996
rect 15531 38947 15573 38956
rect 16867 38996 16925 38997
rect 16867 38956 16876 38996
rect 16916 38956 16925 38996
rect 16867 38955 16925 38956
rect 17251 38996 17309 38997
rect 17251 38956 17260 38996
rect 17300 38956 17309 38996
rect 17251 38955 17309 38956
rect 17827 38996 17885 38997
rect 17827 38956 17836 38996
rect 17876 38956 17885 38996
rect 17827 38955 17885 38956
rect 18691 38996 18749 38997
rect 18691 38956 18700 38996
rect 18740 38956 18749 38996
rect 18691 38955 18749 38956
rect 19267 38996 19325 38997
rect 19267 38956 19276 38996
rect 19316 38956 19325 38996
rect 19267 38955 19325 38956
rect 19651 38996 19709 38997
rect 19651 38956 19660 38996
rect 19700 38956 19709 38996
rect 19651 38955 19709 38956
rect 20035 38996 20093 38997
rect 20035 38956 20044 38996
rect 20084 38956 20093 38996
rect 20035 38955 20093 38956
rect 7371 38926 7413 38935
rect 1699 38912 1757 38913
rect 1699 38872 1708 38912
rect 1748 38872 1757 38912
rect 1699 38871 1757 38872
rect 2947 38912 3005 38913
rect 2947 38872 2956 38912
rect 2996 38872 3005 38912
rect 2947 38871 3005 38872
rect 5835 38912 5877 38921
rect 5835 38872 5836 38912
rect 5876 38872 5877 38912
rect 5835 38863 5877 38872
rect 5931 38912 5973 38921
rect 5931 38872 5932 38912
rect 5972 38872 5973 38912
rect 5931 38863 5973 38872
rect 6411 38912 6453 38921
rect 6411 38872 6412 38912
rect 6452 38872 6453 38912
rect 6411 38863 6453 38872
rect 6883 38912 6941 38913
rect 6883 38872 6892 38912
rect 6932 38872 6941 38912
rect 7371 38886 7372 38926
rect 7412 38886 7413 38926
rect 9387 38926 9429 38935
rect 7371 38877 7413 38886
rect 7851 38912 7893 38921
rect 6883 38871 6941 38872
rect 7851 38872 7852 38912
rect 7892 38872 7893 38912
rect 7851 38863 7893 38872
rect 7947 38912 7989 38921
rect 7947 38872 7948 38912
rect 7988 38872 7989 38912
rect 7947 38863 7989 38872
rect 8427 38912 8469 38921
rect 8427 38872 8428 38912
rect 8468 38872 8469 38912
rect 8427 38863 8469 38872
rect 8899 38912 8957 38913
rect 8899 38872 8908 38912
rect 8948 38872 8957 38912
rect 9387 38886 9388 38926
rect 9428 38886 9429 38926
rect 16539 38921 16581 38930
rect 9387 38877 9429 38886
rect 10243 38912 10301 38913
rect 8899 38871 8957 38872
rect 10243 38872 10252 38912
rect 10292 38872 10301 38912
rect 10243 38871 10301 38872
rect 11491 38912 11549 38913
rect 11491 38872 11500 38912
rect 11540 38872 11549 38912
rect 11491 38871 11549 38872
rect 12547 38912 12605 38913
rect 12547 38872 12556 38912
rect 12596 38872 12605 38912
rect 12547 38871 12605 38872
rect 13795 38912 13853 38913
rect 13795 38872 13804 38912
rect 13844 38872 13853 38912
rect 13795 38871 13853 38872
rect 14955 38912 14997 38921
rect 14955 38872 14956 38912
rect 14996 38872 14997 38912
rect 14955 38863 14997 38872
rect 15051 38912 15093 38921
rect 15051 38872 15052 38912
rect 15092 38872 15093 38912
rect 15051 38863 15093 38872
rect 15435 38912 15477 38921
rect 15435 38872 15436 38912
rect 15476 38872 15477 38912
rect 15435 38863 15477 38872
rect 16003 38912 16061 38913
rect 16003 38872 16012 38912
rect 16052 38872 16061 38912
rect 16539 38881 16540 38921
rect 16580 38881 16581 38921
rect 16539 38872 16581 38881
rect 16003 38871 16061 38872
rect 3147 38744 3189 38753
rect 3147 38704 3148 38744
rect 3188 38704 3189 38744
rect 3147 38695 3189 38704
rect 3331 38744 3389 38745
rect 3331 38704 3340 38744
rect 3380 38704 3389 38744
rect 3331 38703 3389 38704
rect 7563 38744 7605 38753
rect 7563 38704 7564 38744
rect 7604 38704 7605 38744
rect 7563 38695 7605 38704
rect 9579 38744 9621 38753
rect 9579 38704 9580 38744
rect 9620 38704 9621 38744
rect 9579 38695 9621 38704
rect 11691 38744 11733 38753
rect 11691 38704 11692 38744
rect 11732 38704 11733 38744
rect 11691 38695 11733 38704
rect 12267 38744 12309 38753
rect 12267 38704 12268 38744
rect 12308 38704 12309 38744
rect 12267 38695 12309 38704
rect 13995 38744 14037 38753
rect 13995 38704 13996 38744
rect 14036 38704 14037 38744
rect 13995 38695 14037 38704
rect 16683 38744 16725 38753
rect 16683 38704 16684 38744
rect 16724 38704 16725 38744
rect 16683 38695 16725 38704
rect 17067 38744 17109 38753
rect 17067 38704 17068 38744
rect 17108 38704 17109 38744
rect 17067 38695 17109 38704
rect 18211 38744 18269 38745
rect 18211 38704 18220 38744
rect 18260 38704 18269 38744
rect 18211 38703 18269 38704
rect 18979 38744 19037 38745
rect 18979 38704 18988 38744
rect 19028 38704 19037 38744
rect 18979 38703 19037 38704
rect 19467 38744 19509 38753
rect 19467 38704 19468 38744
rect 19508 38704 19509 38744
rect 19467 38695 19509 38704
rect 19851 38744 19893 38753
rect 19851 38704 19852 38744
rect 19892 38704 19893 38744
rect 19851 38695 19893 38704
rect 20235 38744 20277 38753
rect 20235 38704 20236 38744
rect 20276 38704 20277 38744
rect 20235 38695 20277 38704
rect 1152 38576 20452 38600
rect 1152 38536 4928 38576
rect 4968 38536 5010 38576
rect 5050 38536 5092 38576
rect 5132 38536 5174 38576
rect 5214 38536 5256 38576
rect 5296 38536 20048 38576
rect 20088 38536 20130 38576
rect 20170 38536 20212 38576
rect 20252 38536 20294 38576
rect 20334 38536 20376 38576
rect 20416 38536 20452 38576
rect 1152 38512 20452 38536
rect 1419 38408 1461 38417
rect 1419 38368 1420 38408
rect 1460 38368 1461 38408
rect 1419 38359 1461 38368
rect 1803 38408 1845 38417
rect 1803 38368 1804 38408
rect 1844 38368 1845 38408
rect 1803 38359 1845 38368
rect 6891 38408 6933 38417
rect 6891 38368 6892 38408
rect 6932 38368 6933 38408
rect 6891 38359 6933 38368
rect 7275 38408 7317 38417
rect 7275 38368 7276 38408
rect 7316 38368 7317 38408
rect 7275 38359 7317 38368
rect 12267 38408 12309 38417
rect 12267 38368 12268 38408
rect 12308 38368 12309 38408
rect 12267 38359 12309 38368
rect 12651 38408 12693 38417
rect 12651 38368 12652 38408
rect 12692 38368 12693 38408
rect 12651 38359 12693 38368
rect 13035 38408 13077 38417
rect 13035 38368 13036 38408
rect 13076 38368 13077 38408
rect 13035 38359 13077 38368
rect 13419 38408 13461 38417
rect 13419 38368 13420 38408
rect 13460 38368 13461 38408
rect 13419 38359 13461 38368
rect 17067 38408 17109 38417
rect 17067 38368 17068 38408
rect 17108 38368 17109 38408
rect 17067 38359 17109 38368
rect 19179 38408 19221 38417
rect 19179 38368 19180 38408
rect 19220 38368 19221 38408
rect 19179 38359 19221 38368
rect 4203 38324 4245 38333
rect 4203 38284 4204 38324
rect 4244 38284 4245 38324
rect 4203 38275 4245 38284
rect 6507 38324 6549 38333
rect 6507 38284 6508 38324
rect 6548 38284 6549 38324
rect 6507 38275 6549 38284
rect 11691 38324 11733 38333
rect 11691 38284 11692 38324
rect 11732 38284 11733 38324
rect 11691 38275 11733 38284
rect 20139 38324 20181 38333
rect 20139 38284 20140 38324
rect 20180 38284 20181 38324
rect 20139 38275 20181 38284
rect 2475 38240 2517 38249
rect 2475 38200 2476 38240
rect 2516 38200 2517 38240
rect 2475 38191 2517 38200
rect 2571 38240 2613 38249
rect 2571 38200 2572 38240
rect 2612 38200 2613 38240
rect 2571 38191 2613 38200
rect 3523 38240 3581 38241
rect 3523 38200 3532 38240
rect 3572 38200 3581 38240
rect 3523 38199 3581 38200
rect 4011 38235 4053 38244
rect 4011 38195 4012 38235
rect 4052 38195 4053 38235
rect 4011 38186 4053 38195
rect 4779 38240 4821 38249
rect 4779 38200 4780 38240
rect 4820 38200 4821 38240
rect 4779 38191 4821 38200
rect 4875 38240 4917 38249
rect 4875 38200 4876 38240
rect 4916 38200 4917 38240
rect 4875 38191 4917 38200
rect 5827 38240 5885 38241
rect 5827 38200 5836 38240
rect 5876 38200 5885 38240
rect 7843 38240 7901 38241
rect 5827 38199 5885 38200
rect 6363 38198 6405 38207
rect 7843 38200 7852 38240
rect 7892 38200 7901 38240
rect 7843 38199 7901 38200
rect 9091 38240 9149 38241
rect 9091 38200 9100 38240
rect 9140 38200 9149 38240
rect 9091 38199 9149 38200
rect 9579 38240 9621 38249
rect 9579 38200 9580 38240
rect 9620 38200 9621 38240
rect 1219 38156 1277 38157
rect 1219 38116 1228 38156
rect 1268 38116 1277 38156
rect 1219 38115 1277 38116
rect 1603 38156 1661 38157
rect 1603 38116 1612 38156
rect 1652 38116 1661 38156
rect 1603 38115 1661 38116
rect 1987 38156 2045 38157
rect 1987 38116 1996 38156
rect 2036 38116 2045 38156
rect 1987 38115 2045 38116
rect 2955 38156 2997 38165
rect 2955 38116 2956 38156
rect 2996 38116 2997 38156
rect 2955 38107 2997 38116
rect 3051 38156 3093 38165
rect 3051 38116 3052 38156
rect 3092 38116 3093 38156
rect 3051 38107 3093 38116
rect 5259 38156 5301 38165
rect 5259 38116 5260 38156
rect 5300 38116 5301 38156
rect 5259 38107 5301 38116
rect 5355 38156 5397 38165
rect 5355 38116 5356 38156
rect 5396 38116 5397 38156
rect 6363 38158 6364 38198
rect 6404 38158 6405 38198
rect 9579 38191 9621 38200
rect 9963 38240 10005 38249
rect 9963 38200 9964 38240
rect 10004 38200 10005 38240
rect 9963 38191 10005 38200
rect 10059 38240 10101 38249
rect 10059 38200 10060 38240
rect 10100 38200 10101 38240
rect 10059 38191 10101 38200
rect 10539 38240 10581 38249
rect 10539 38200 10540 38240
rect 10580 38200 10581 38240
rect 10539 38191 10581 38200
rect 11011 38240 11069 38241
rect 11011 38200 11020 38240
rect 11060 38200 11069 38240
rect 13603 38240 13661 38241
rect 11011 38199 11069 38200
rect 11547 38230 11589 38239
rect 11547 38190 11548 38230
rect 11588 38190 11589 38230
rect 13603 38200 13612 38240
rect 13652 38200 13661 38240
rect 13603 38199 13661 38200
rect 14851 38240 14909 38241
rect 14851 38200 14860 38240
rect 14900 38200 14909 38240
rect 14851 38199 14909 38200
rect 15339 38240 15381 38249
rect 15339 38200 15340 38240
rect 15380 38200 15381 38240
rect 15339 38191 15381 38200
rect 15435 38240 15477 38249
rect 15435 38200 15436 38240
rect 15476 38200 15477 38240
rect 15435 38191 15477 38200
rect 15819 38240 15861 38249
rect 15819 38200 15820 38240
rect 15860 38200 15861 38240
rect 15819 38191 15861 38200
rect 15915 38240 15957 38249
rect 15915 38200 15916 38240
rect 15956 38200 15957 38240
rect 15915 38191 15957 38200
rect 16387 38240 16445 38241
rect 16387 38200 16396 38240
rect 16436 38200 16445 38240
rect 17443 38240 17501 38241
rect 16387 38199 16445 38200
rect 16875 38226 16917 38235
rect 11547 38181 11589 38190
rect 16875 38186 16876 38226
rect 16916 38186 16917 38226
rect 17443 38200 17452 38240
rect 17492 38200 17501 38240
rect 17443 38199 17501 38200
rect 18691 38240 18749 38241
rect 18691 38200 18700 38240
rect 18740 38200 18749 38240
rect 18691 38199 18749 38200
rect 16875 38177 16917 38186
rect 6363 38149 6405 38158
rect 7075 38156 7133 38157
rect 5355 38107 5397 38116
rect 7075 38116 7084 38156
rect 7124 38116 7133 38156
rect 7075 38115 7133 38116
rect 7459 38156 7517 38157
rect 7459 38116 7468 38156
rect 7508 38116 7517 38156
rect 7459 38115 7517 38116
rect 10443 38156 10485 38165
rect 10443 38116 10444 38156
rect 10484 38116 10485 38156
rect 10443 38107 10485 38116
rect 12067 38156 12125 38157
rect 12067 38116 12076 38156
rect 12116 38116 12125 38156
rect 12067 38115 12125 38116
rect 12451 38156 12509 38157
rect 12451 38116 12460 38156
rect 12500 38116 12509 38156
rect 12451 38115 12509 38116
rect 12835 38156 12893 38157
rect 12835 38116 12844 38156
rect 12884 38116 12893 38156
rect 12835 38115 12893 38116
rect 13219 38156 13277 38157
rect 13219 38116 13228 38156
rect 13268 38116 13277 38156
rect 13219 38115 13277 38116
rect 18979 38156 19037 38157
rect 18979 38116 18988 38156
rect 19028 38116 19037 38156
rect 18979 38115 19037 38116
rect 19363 38156 19421 38157
rect 19363 38116 19372 38156
rect 19412 38116 19421 38156
rect 19363 38115 19421 38116
rect 19747 38156 19805 38157
rect 19747 38116 19756 38156
rect 19796 38116 19805 38156
rect 19747 38115 19805 38116
rect 15051 38072 15093 38081
rect 15051 38032 15052 38072
rect 15092 38032 15093 38072
rect 15051 38023 15093 38032
rect 2187 37988 2229 37997
rect 2187 37948 2188 37988
rect 2228 37948 2229 37988
rect 2187 37939 2229 37948
rect 9291 37988 9333 37997
rect 9291 37948 9292 37988
rect 9332 37948 9333 37988
rect 9291 37939 9333 37948
rect 17259 37988 17301 37997
rect 17259 37948 17260 37988
rect 17300 37948 17301 37988
rect 17259 37939 17301 37948
rect 19563 37988 19605 37997
rect 19563 37948 19564 37988
rect 19604 37948 19605 37988
rect 19563 37939 19605 37948
rect 19947 37988 19989 37997
rect 19947 37948 19948 37988
rect 19988 37948 19989 37988
rect 19947 37939 19989 37948
rect 1152 37820 20352 37844
rect 1152 37780 3688 37820
rect 3728 37780 3770 37820
rect 3810 37780 3852 37820
rect 3892 37780 3934 37820
rect 3974 37780 4016 37820
rect 4056 37780 18808 37820
rect 18848 37780 18890 37820
rect 18930 37780 18972 37820
rect 19012 37780 19054 37820
rect 19094 37780 19136 37820
rect 19176 37780 20352 37820
rect 1152 37756 20352 37780
rect 1803 37652 1845 37661
rect 1803 37612 1804 37652
rect 1844 37612 1845 37652
rect 1803 37603 1845 37612
rect 4683 37652 4725 37661
rect 4683 37612 4684 37652
rect 4724 37612 4725 37652
rect 4683 37603 4725 37612
rect 5067 37652 5109 37661
rect 5067 37612 5068 37652
rect 5108 37612 5109 37652
rect 5067 37603 5109 37612
rect 5451 37652 5493 37661
rect 5451 37612 5452 37652
rect 5492 37612 5493 37652
rect 5451 37603 5493 37612
rect 15435 37652 15477 37661
rect 15435 37612 15436 37652
rect 15476 37612 15477 37652
rect 15435 37603 15477 37612
rect 17067 37652 17109 37661
rect 17067 37612 17068 37652
rect 17108 37612 17109 37652
rect 17067 37603 17109 37612
rect 1419 37568 1461 37577
rect 1419 37528 1420 37568
rect 1460 37528 1461 37568
rect 1419 37519 1461 37528
rect 7371 37568 7413 37577
rect 7371 37528 7372 37568
rect 7412 37528 7413 37568
rect 7371 37519 7413 37528
rect 17451 37568 17493 37577
rect 17451 37528 17452 37568
rect 17492 37528 17493 37568
rect 17451 37519 17493 37528
rect 1219 37484 1277 37485
rect 1219 37444 1228 37484
rect 1268 37444 1277 37484
rect 1219 37443 1277 37444
rect 1603 37484 1661 37485
rect 1603 37444 1612 37484
rect 1652 37444 1661 37484
rect 4483 37484 4541 37485
rect 1603 37443 1661 37444
rect 4059 37442 4101 37451
rect 4483 37444 4492 37484
rect 4532 37444 4541 37484
rect 4483 37443 4541 37444
rect 4867 37484 4925 37485
rect 4867 37444 4876 37484
rect 4916 37444 4925 37484
rect 4867 37443 4925 37444
rect 5251 37484 5309 37485
rect 5251 37444 5260 37484
rect 5300 37444 5309 37484
rect 15235 37484 15293 37485
rect 5251 37443 5309 37444
rect 2475 37400 2517 37409
rect 2475 37360 2476 37400
rect 2516 37360 2517 37400
rect 2475 37351 2517 37360
rect 2571 37400 2613 37409
rect 2571 37360 2572 37400
rect 2612 37360 2613 37400
rect 2571 37351 2613 37360
rect 2955 37400 2997 37409
rect 2955 37360 2956 37400
rect 2996 37360 2997 37400
rect 2955 37351 2997 37360
rect 3051 37400 3093 37409
rect 4059 37402 4060 37442
rect 4100 37402 4101 37442
rect 9243 37442 9285 37451
rect 15235 37444 15244 37484
rect 15284 37444 15293 37484
rect 15235 37443 15293 37444
rect 17251 37484 17309 37485
rect 17251 37444 17260 37484
rect 17300 37444 17309 37484
rect 17251 37443 17309 37444
rect 18219 37484 18261 37493
rect 18219 37444 18220 37484
rect 18260 37444 18261 37484
rect 3051 37360 3052 37400
rect 3092 37360 3093 37400
rect 3051 37351 3093 37360
rect 3523 37400 3581 37401
rect 3523 37360 3532 37400
rect 3572 37360 3581 37400
rect 4059 37393 4101 37402
rect 5635 37400 5693 37401
rect 3523 37359 3581 37360
rect 5635 37360 5644 37400
rect 5684 37360 5693 37400
rect 5635 37359 5693 37360
rect 6883 37400 6941 37401
rect 6883 37360 6892 37400
rect 6932 37360 6941 37400
rect 6883 37359 6941 37360
rect 7659 37400 7701 37409
rect 7659 37360 7660 37400
rect 7700 37360 7701 37400
rect 7659 37351 7701 37360
rect 7755 37400 7797 37409
rect 7755 37360 7756 37400
rect 7796 37360 7797 37400
rect 7755 37351 7797 37360
rect 8139 37400 8181 37409
rect 8139 37360 8140 37400
rect 8180 37360 8181 37400
rect 8139 37351 8181 37360
rect 8235 37400 8277 37409
rect 9243 37402 9244 37442
rect 9284 37402 9285 37442
rect 18219 37435 18261 37444
rect 19651 37484 19709 37485
rect 19651 37444 19660 37484
rect 19700 37444 19709 37484
rect 19651 37443 19709 37444
rect 20035 37484 20093 37485
rect 20035 37444 20044 37484
rect 20084 37444 20093 37484
rect 20035 37443 20093 37444
rect 19275 37414 19317 37423
rect 8235 37360 8236 37400
rect 8276 37360 8277 37400
rect 8235 37351 8277 37360
rect 8707 37400 8765 37401
rect 8707 37360 8716 37400
rect 8756 37360 8765 37400
rect 9243 37393 9285 37402
rect 9763 37400 9821 37401
rect 8707 37359 8765 37360
rect 9763 37360 9772 37400
rect 9812 37360 9821 37400
rect 9763 37359 9821 37360
rect 11011 37400 11069 37401
rect 11011 37360 11020 37400
rect 11060 37360 11069 37400
rect 11011 37359 11069 37360
rect 11491 37400 11549 37401
rect 11491 37360 11500 37400
rect 11540 37360 11549 37400
rect 11491 37359 11549 37360
rect 12739 37400 12797 37401
rect 12739 37360 12748 37400
rect 12788 37360 12797 37400
rect 12739 37359 12797 37360
rect 13315 37400 13373 37401
rect 13315 37360 13324 37400
rect 13364 37360 13373 37400
rect 13315 37359 13373 37360
rect 14563 37400 14621 37401
rect 14563 37360 14572 37400
rect 14612 37360 14621 37400
rect 14563 37359 14621 37360
rect 15619 37400 15677 37401
rect 15619 37360 15628 37400
rect 15668 37360 15677 37400
rect 15619 37359 15677 37360
rect 16867 37400 16925 37401
rect 16867 37360 16876 37400
rect 16916 37360 16925 37400
rect 16867 37359 16925 37360
rect 17739 37400 17781 37409
rect 17739 37360 17740 37400
rect 17780 37360 17781 37400
rect 17739 37351 17781 37360
rect 17835 37400 17877 37409
rect 17835 37360 17836 37400
rect 17876 37360 17877 37400
rect 17835 37351 17877 37360
rect 18315 37400 18357 37409
rect 18315 37360 18316 37400
rect 18356 37360 18357 37400
rect 18315 37351 18357 37360
rect 18787 37400 18845 37401
rect 18787 37360 18796 37400
rect 18836 37360 18845 37400
rect 19275 37374 19276 37414
rect 19316 37374 19317 37414
rect 19275 37365 19317 37374
rect 18787 37359 18845 37360
rect 7083 37316 7125 37325
rect 7083 37276 7084 37316
rect 7124 37276 7125 37316
rect 7083 37267 7125 37276
rect 19467 37316 19509 37325
rect 19467 37276 19468 37316
rect 19508 37276 19509 37316
rect 19467 37267 19509 37276
rect 1987 37232 2045 37233
rect 1987 37192 1996 37232
rect 2036 37192 2045 37232
rect 1987 37191 2045 37192
rect 4203 37232 4245 37241
rect 4203 37192 4204 37232
rect 4244 37192 4245 37232
rect 4203 37183 4245 37192
rect 7267 37232 7325 37233
rect 7267 37192 7276 37232
rect 7316 37192 7325 37232
rect 9579 37232 9621 37241
rect 7267 37191 7325 37192
rect 9387 37190 9429 37199
rect 9387 37150 9388 37190
rect 9428 37150 9429 37190
rect 9579 37192 9580 37232
rect 9620 37192 9621 37232
rect 9579 37183 9621 37192
rect 12939 37232 12981 37241
rect 12939 37192 12940 37232
rect 12980 37192 12981 37232
rect 12939 37183 12981 37192
rect 14763 37232 14805 37241
rect 14763 37192 14764 37232
rect 14804 37192 14805 37232
rect 14763 37183 14805 37192
rect 19851 37232 19893 37241
rect 19851 37192 19852 37232
rect 19892 37192 19893 37232
rect 19851 37183 19893 37192
rect 20235 37232 20277 37241
rect 20235 37192 20236 37232
rect 20276 37192 20277 37232
rect 20235 37183 20277 37192
rect 9387 37141 9429 37150
rect 1152 37064 20452 37088
rect 1152 37024 4928 37064
rect 4968 37024 5010 37064
rect 5050 37024 5092 37064
rect 5132 37024 5174 37064
rect 5214 37024 5256 37064
rect 5296 37024 20048 37064
rect 20088 37024 20130 37064
rect 20170 37024 20212 37064
rect 20252 37024 20294 37064
rect 20334 37024 20376 37064
rect 20416 37024 20452 37064
rect 1152 37000 20452 37024
rect 1515 36896 1557 36905
rect 1515 36856 1516 36896
rect 1556 36856 1557 36896
rect 1515 36847 1557 36856
rect 1899 36896 1941 36905
rect 1899 36856 1900 36896
rect 1940 36856 1941 36896
rect 1899 36847 1941 36856
rect 3819 36896 3861 36905
rect 3819 36856 3820 36896
rect 3860 36856 3861 36896
rect 3819 36847 3861 36856
rect 4683 36896 4725 36905
rect 4683 36856 4684 36896
rect 4724 36856 4725 36896
rect 4683 36847 4725 36856
rect 7083 36896 7125 36905
rect 7083 36856 7084 36896
rect 7124 36856 7125 36896
rect 7083 36847 7125 36856
rect 14667 36896 14709 36905
rect 14667 36856 14668 36896
rect 14708 36856 14709 36896
rect 14667 36847 14709 36856
rect 15051 36896 15093 36905
rect 15051 36856 15052 36896
rect 15092 36856 15093 36896
rect 15051 36847 15093 36856
rect 17067 36896 17109 36905
rect 17067 36856 17068 36896
rect 17108 36856 17109 36896
rect 17067 36847 17109 36856
rect 19179 36896 19221 36905
rect 19179 36856 19180 36896
rect 19220 36856 19221 36896
rect 19179 36847 19221 36856
rect 19563 36896 19605 36905
rect 19563 36856 19564 36896
rect 19604 36856 19605 36896
rect 19563 36847 19605 36856
rect 12171 36812 12213 36821
rect 12171 36772 12172 36812
rect 12212 36772 12213 36812
rect 12171 36763 12213 36772
rect 14187 36812 14229 36821
rect 14187 36772 14188 36812
rect 14228 36772 14229 36812
rect 14187 36763 14229 36772
rect 4963 36728 5021 36729
rect 4963 36688 4972 36728
rect 5012 36688 5021 36728
rect 4963 36687 5021 36688
rect 6211 36728 6269 36729
rect 6211 36688 6220 36728
rect 6260 36688 6269 36728
rect 6211 36687 6269 36688
rect 7459 36728 7517 36729
rect 7459 36688 7468 36728
rect 7508 36688 7517 36728
rect 7459 36687 7517 36688
rect 8707 36728 8765 36729
rect 8707 36688 8716 36728
rect 8756 36688 8765 36728
rect 8707 36687 8765 36688
rect 9091 36728 9149 36729
rect 9091 36688 9100 36728
rect 9140 36688 9149 36728
rect 9091 36687 9149 36688
rect 10339 36728 10397 36729
rect 10339 36688 10348 36728
rect 10388 36688 10397 36728
rect 10339 36687 10397 36688
rect 10723 36728 10781 36729
rect 10723 36688 10732 36728
rect 10772 36688 10781 36728
rect 10723 36687 10781 36688
rect 12459 36728 12501 36737
rect 12459 36688 12460 36728
rect 12500 36688 12501 36728
rect 11971 36686 12029 36687
rect 1315 36644 1373 36645
rect 1315 36604 1324 36644
rect 1364 36604 1373 36644
rect 1315 36603 1373 36604
rect 1699 36644 1757 36645
rect 1699 36604 1708 36644
rect 1748 36604 1757 36644
rect 1699 36603 1757 36604
rect 2179 36644 2237 36645
rect 2179 36604 2188 36644
rect 2228 36604 2237 36644
rect 2179 36603 2237 36604
rect 4299 36644 4341 36653
rect 11971 36646 11980 36686
rect 12020 36646 12029 36686
rect 12459 36679 12501 36688
rect 12555 36728 12597 36737
rect 12555 36688 12556 36728
rect 12596 36688 12597 36728
rect 12555 36679 12597 36688
rect 13507 36728 13565 36729
rect 13507 36688 13516 36728
rect 13556 36688 13565 36728
rect 13507 36687 13565 36688
rect 13995 36723 14037 36732
rect 13995 36683 13996 36723
rect 14036 36683 14037 36723
rect 13995 36674 14037 36683
rect 15339 36728 15381 36737
rect 15339 36688 15340 36728
rect 15380 36688 15381 36728
rect 15339 36679 15381 36688
rect 15435 36728 15477 36737
rect 15435 36688 15436 36728
rect 15476 36688 15477 36728
rect 15435 36679 15477 36688
rect 16387 36728 16445 36729
rect 16387 36688 16396 36728
rect 16436 36688 16445 36728
rect 17443 36728 17501 36729
rect 16387 36687 16445 36688
rect 16875 36714 16917 36723
rect 16875 36674 16876 36714
rect 16916 36674 16917 36714
rect 17443 36688 17452 36728
rect 17492 36688 17501 36728
rect 17443 36687 17501 36688
rect 18691 36728 18749 36729
rect 18691 36688 18700 36728
rect 18740 36688 18749 36728
rect 18691 36687 18749 36688
rect 16875 36665 16917 36674
rect 11971 36645 12029 36646
rect 4299 36604 4300 36644
rect 4340 36604 4341 36644
rect 4299 36595 4341 36604
rect 4483 36644 4541 36645
rect 4483 36604 4492 36644
rect 4532 36604 4541 36644
rect 4483 36603 4541 36604
rect 6883 36644 6941 36645
rect 6883 36604 6892 36644
rect 6932 36604 6941 36644
rect 6883 36603 6941 36604
rect 12939 36644 12981 36653
rect 12939 36604 12940 36644
rect 12980 36604 12981 36644
rect 12939 36595 12981 36604
rect 13035 36644 13077 36653
rect 13035 36604 13036 36644
rect 13076 36604 13077 36644
rect 13035 36595 13077 36604
rect 14467 36644 14525 36645
rect 14467 36604 14476 36644
rect 14516 36604 14525 36644
rect 14467 36603 14525 36604
rect 14851 36644 14909 36645
rect 14851 36604 14860 36644
rect 14900 36604 14909 36644
rect 14851 36603 14909 36604
rect 15819 36644 15861 36653
rect 15819 36604 15820 36644
rect 15860 36604 15861 36644
rect 15819 36595 15861 36604
rect 15915 36644 15957 36653
rect 15915 36604 15916 36644
rect 15956 36604 15957 36644
rect 15915 36595 15957 36604
rect 18979 36644 19037 36645
rect 18979 36604 18988 36644
rect 19028 36604 19037 36644
rect 18979 36603 19037 36604
rect 19363 36644 19421 36645
rect 19363 36604 19372 36644
rect 19412 36604 19421 36644
rect 19363 36603 19421 36604
rect 19747 36644 19805 36645
rect 19747 36604 19756 36644
rect 19796 36604 19805 36644
rect 19747 36603 19805 36604
rect 2379 36560 2421 36569
rect 2379 36520 2380 36560
rect 2420 36520 2421 36560
rect 2379 36511 2421 36520
rect 6699 36560 6741 36569
rect 6699 36520 6700 36560
rect 6740 36520 6741 36560
rect 6699 36511 6741 36520
rect 19947 36560 19989 36569
rect 19947 36520 19948 36560
rect 19988 36520 19989 36560
rect 19947 36511 19989 36520
rect 6411 36476 6453 36485
rect 6411 36436 6412 36476
rect 6452 36436 6453 36476
rect 6411 36427 6453 36436
rect 8907 36476 8949 36485
rect 8907 36436 8908 36476
rect 8948 36436 8949 36476
rect 8907 36427 8949 36436
rect 10539 36476 10581 36485
rect 10539 36436 10540 36476
rect 10580 36436 10581 36476
rect 10539 36427 10581 36436
rect 17259 36476 17301 36485
rect 17259 36436 17260 36476
rect 17300 36436 17301 36476
rect 17259 36427 17301 36436
rect 1152 36308 20352 36332
rect 1152 36268 3688 36308
rect 3728 36268 3770 36308
rect 3810 36268 3852 36308
rect 3892 36268 3934 36308
rect 3974 36268 4016 36308
rect 4056 36268 18808 36308
rect 18848 36268 18890 36308
rect 18930 36268 18972 36308
rect 19012 36268 19054 36308
rect 19094 36268 19136 36308
rect 19176 36268 20352 36308
rect 1152 36244 20352 36268
rect 1515 36140 1557 36149
rect 1515 36100 1516 36140
rect 1556 36100 1557 36140
rect 1515 36091 1557 36100
rect 3435 36140 3477 36149
rect 3435 36100 3436 36140
rect 3476 36100 3477 36140
rect 3435 36091 3477 36100
rect 4011 36140 4053 36149
rect 4011 36100 4012 36140
rect 4052 36100 4053 36140
rect 4011 36091 4053 36100
rect 11595 36140 11637 36149
rect 11595 36100 11596 36140
rect 11636 36100 11637 36140
rect 11595 36091 11637 36100
rect 12363 36140 12405 36149
rect 12363 36100 12364 36140
rect 12404 36100 12405 36140
rect 12363 36091 12405 36100
rect 15051 36140 15093 36149
rect 15051 36100 15052 36140
rect 15092 36100 15093 36140
rect 15051 36091 15093 36100
rect 16683 36140 16725 36149
rect 16683 36100 16684 36140
rect 16724 36100 16725 36140
rect 16683 36091 16725 36100
rect 1315 35972 1373 35973
rect 1315 35932 1324 35972
rect 1364 35932 1373 35972
rect 1315 35931 1373 35932
rect 3619 35972 3677 35973
rect 3619 35932 3628 35972
rect 3668 35932 3677 35972
rect 3619 35931 3677 35932
rect 3811 35972 3869 35973
rect 3811 35932 3820 35972
rect 3860 35932 3869 35972
rect 3811 35931 3869 35932
rect 6987 35972 7029 35981
rect 6987 35932 6988 35972
rect 7028 35932 7029 35972
rect 6987 35923 7029 35932
rect 7083 35972 7125 35981
rect 7083 35932 7084 35972
rect 7124 35932 7125 35972
rect 7083 35923 7125 35932
rect 11395 35972 11453 35973
rect 11395 35932 11404 35972
rect 11444 35932 11453 35972
rect 19939 35972 19997 35973
rect 11395 35931 11453 35932
rect 14715 35930 14757 35939
rect 19939 35932 19948 35972
rect 19988 35932 19997 35972
rect 19939 35931 19997 35932
rect 11019 35902 11061 35911
rect 4963 35888 5021 35889
rect 4963 35848 4972 35888
rect 5012 35848 5021 35888
rect 4963 35847 5021 35848
rect 6211 35888 6269 35889
rect 6211 35848 6220 35888
rect 6260 35848 6269 35888
rect 6211 35847 6269 35848
rect 6507 35888 6549 35897
rect 6507 35848 6508 35888
rect 6548 35848 6549 35888
rect 6507 35839 6549 35848
rect 6603 35888 6645 35897
rect 8043 35893 8085 35902
rect 6603 35848 6604 35888
rect 6644 35848 6645 35888
rect 6603 35839 6645 35848
rect 7555 35888 7613 35889
rect 7555 35848 7564 35888
rect 7604 35848 7613 35888
rect 7555 35847 7613 35848
rect 8043 35853 8044 35893
rect 8084 35853 8085 35893
rect 8043 35844 8085 35853
rect 9483 35888 9525 35897
rect 9483 35848 9484 35888
rect 9524 35848 9525 35888
rect 9483 35839 9525 35848
rect 9579 35888 9621 35897
rect 9579 35848 9580 35888
rect 9620 35848 9621 35888
rect 9579 35839 9621 35848
rect 9963 35888 10005 35897
rect 9963 35848 9964 35888
rect 10004 35848 10005 35888
rect 9963 35839 10005 35848
rect 10059 35888 10101 35897
rect 10059 35848 10060 35888
rect 10100 35848 10101 35888
rect 10059 35839 10101 35848
rect 10531 35888 10589 35889
rect 10531 35848 10540 35888
rect 10580 35848 10589 35888
rect 11019 35862 11020 35902
rect 11060 35862 11061 35902
rect 11019 35853 11061 35862
rect 11875 35888 11933 35889
rect 10531 35847 10589 35848
rect 11875 35848 11884 35888
rect 11924 35848 11933 35888
rect 11875 35847 11933 35848
rect 13131 35888 13173 35897
rect 13131 35848 13132 35888
rect 13172 35848 13173 35888
rect 13131 35839 13173 35848
rect 13227 35888 13269 35897
rect 13227 35848 13228 35888
rect 13268 35848 13269 35888
rect 13227 35839 13269 35848
rect 13611 35888 13653 35897
rect 13611 35848 13612 35888
rect 13652 35848 13653 35888
rect 13611 35839 13653 35848
rect 13707 35888 13749 35897
rect 14715 35890 14716 35930
rect 14756 35890 14757 35930
rect 13707 35848 13708 35888
rect 13748 35848 13749 35888
rect 13707 35839 13749 35848
rect 14179 35888 14237 35889
rect 14179 35848 14188 35888
rect 14228 35848 14237 35888
rect 14715 35881 14757 35890
rect 15235 35888 15293 35889
rect 14179 35847 14237 35848
rect 15235 35848 15244 35888
rect 15284 35848 15293 35888
rect 15235 35847 15293 35848
rect 16483 35888 16541 35889
rect 16483 35848 16492 35888
rect 16532 35848 16541 35888
rect 16483 35847 16541 35848
rect 16867 35888 16925 35889
rect 16867 35848 16876 35888
rect 16916 35848 16925 35888
rect 16867 35847 16925 35848
rect 18115 35888 18173 35889
rect 18115 35848 18124 35888
rect 18164 35848 18173 35888
rect 18115 35847 18173 35848
rect 18307 35888 18365 35889
rect 18307 35848 18316 35888
rect 18356 35848 18365 35888
rect 18307 35847 18365 35848
rect 19555 35888 19613 35889
rect 19555 35848 19564 35888
rect 19604 35848 19613 35888
rect 19555 35847 19613 35848
rect 8235 35804 8277 35813
rect 8235 35764 8236 35804
rect 8276 35764 8277 35804
rect 8235 35755 8277 35764
rect 2179 35720 2237 35721
rect 2179 35680 2188 35720
rect 2228 35680 2237 35720
rect 2179 35679 2237 35680
rect 4483 35720 4541 35721
rect 4483 35680 4492 35720
rect 4532 35680 4541 35720
rect 4483 35679 4541 35680
rect 4779 35720 4821 35729
rect 4779 35680 4780 35720
rect 4820 35680 4821 35720
rect 4779 35671 4821 35680
rect 11211 35720 11253 35729
rect 11211 35680 11212 35720
rect 11252 35680 11253 35720
rect 11211 35671 11253 35680
rect 14859 35720 14901 35729
rect 14859 35680 14860 35720
rect 14900 35680 14901 35720
rect 14859 35671 14901 35680
rect 19755 35720 19797 35729
rect 19755 35680 19756 35720
rect 19796 35680 19797 35720
rect 19755 35671 19797 35680
rect 20139 35720 20181 35729
rect 20139 35680 20140 35720
rect 20180 35680 20181 35720
rect 20139 35671 20181 35680
rect 1152 35552 20452 35576
rect 1152 35512 4928 35552
rect 4968 35512 5010 35552
rect 5050 35512 5092 35552
rect 5132 35512 5174 35552
rect 5214 35512 5256 35552
rect 5296 35512 20048 35552
rect 20088 35512 20130 35552
rect 20170 35512 20212 35552
rect 20252 35512 20294 35552
rect 20334 35512 20376 35552
rect 20416 35512 20452 35552
rect 1152 35488 20452 35512
rect 7563 35384 7605 35393
rect 7563 35344 7564 35384
rect 7604 35344 7605 35384
rect 7563 35335 7605 35344
rect 3627 35300 3669 35309
rect 3627 35260 3628 35300
rect 3668 35260 3669 35300
rect 3627 35251 3669 35260
rect 5643 35300 5685 35309
rect 5643 35260 5644 35300
rect 5684 35260 5685 35300
rect 5643 35251 5685 35260
rect 19275 35300 19317 35309
rect 19275 35260 19276 35300
rect 19316 35260 19317 35300
rect 19275 35251 19317 35260
rect 1899 35216 1941 35225
rect 1899 35176 1900 35216
rect 1940 35176 1941 35216
rect 1899 35167 1941 35176
rect 1995 35216 2037 35225
rect 1995 35176 1996 35216
rect 2036 35176 2037 35216
rect 1995 35167 2037 35176
rect 2475 35216 2517 35225
rect 2475 35176 2476 35216
rect 2516 35176 2517 35216
rect 2475 35167 2517 35176
rect 2947 35216 3005 35217
rect 2947 35176 2956 35216
rect 2996 35176 3005 35216
rect 3915 35216 3957 35225
rect 2947 35175 3005 35176
rect 3435 35202 3477 35211
rect 3435 35162 3436 35202
rect 3476 35162 3477 35202
rect 3915 35176 3916 35216
rect 3956 35176 3957 35216
rect 3915 35167 3957 35176
rect 4011 35216 4053 35225
rect 4011 35176 4012 35216
rect 4052 35176 4053 35216
rect 4011 35167 4053 35176
rect 4963 35216 5021 35217
rect 4963 35176 4972 35216
rect 5012 35176 5021 35216
rect 4963 35175 5021 35176
rect 5451 35211 5493 35220
rect 5451 35171 5452 35211
rect 5492 35171 5493 35211
rect 6115 35216 6173 35217
rect 6115 35176 6124 35216
rect 6164 35176 6173 35216
rect 6115 35175 6173 35176
rect 7363 35216 7421 35217
rect 7363 35176 7372 35216
rect 7412 35176 7421 35216
rect 7363 35175 7421 35176
rect 7747 35216 7805 35217
rect 7747 35176 7756 35216
rect 7796 35176 7805 35216
rect 7747 35175 7805 35176
rect 8995 35216 9053 35217
rect 8995 35176 9004 35216
rect 9044 35176 9053 35216
rect 8995 35175 9053 35176
rect 9379 35216 9437 35217
rect 9379 35176 9388 35216
rect 9428 35176 9437 35216
rect 9379 35175 9437 35176
rect 10627 35216 10685 35217
rect 10627 35176 10636 35216
rect 10676 35176 10685 35216
rect 10627 35175 10685 35176
rect 11011 35216 11069 35217
rect 11011 35176 11020 35216
rect 11060 35176 11069 35216
rect 11011 35175 11069 35176
rect 12259 35216 12317 35217
rect 12259 35176 12268 35216
rect 12308 35176 12317 35216
rect 12259 35175 12317 35176
rect 12643 35216 12701 35217
rect 12643 35176 12652 35216
rect 12692 35176 12701 35216
rect 12643 35175 12701 35176
rect 13891 35216 13949 35217
rect 13891 35176 13900 35216
rect 13940 35176 13949 35216
rect 13891 35175 13949 35176
rect 15715 35216 15773 35217
rect 15715 35176 15724 35216
rect 15764 35176 15773 35216
rect 15715 35175 15773 35176
rect 17547 35216 17589 35225
rect 17547 35176 17548 35216
rect 17588 35176 17589 35216
rect 5451 35162 5493 35171
rect 14467 35174 14525 35175
rect 3435 35153 3477 35162
rect 1411 35132 1469 35133
rect 1411 35092 1420 35132
rect 1460 35092 1469 35132
rect 1411 35091 1469 35092
rect 2379 35132 2421 35141
rect 2379 35092 2380 35132
rect 2420 35092 2421 35132
rect 2379 35083 2421 35092
rect 4395 35132 4437 35141
rect 4395 35092 4396 35132
rect 4436 35092 4437 35132
rect 4395 35083 4437 35092
rect 4491 35132 4533 35141
rect 14467 35134 14476 35174
rect 14516 35134 14525 35174
rect 17547 35167 17589 35176
rect 17643 35216 17685 35225
rect 17643 35176 17644 35216
rect 17684 35176 17685 35216
rect 17643 35167 17685 35176
rect 18027 35216 18069 35225
rect 18027 35176 18028 35216
rect 18068 35176 18069 35216
rect 18027 35167 18069 35176
rect 18123 35216 18165 35225
rect 18123 35176 18124 35216
rect 18164 35176 18165 35216
rect 18123 35167 18165 35176
rect 18595 35216 18653 35217
rect 18595 35176 18604 35216
rect 18644 35176 18653 35216
rect 18595 35175 18653 35176
rect 19083 35211 19125 35220
rect 19083 35171 19084 35211
rect 19124 35171 19125 35211
rect 19083 35162 19125 35171
rect 14467 35133 14525 35134
rect 4491 35092 4492 35132
rect 4532 35092 4533 35132
rect 4491 35083 4533 35092
rect 15907 35132 15965 35133
rect 15907 35092 15916 35132
rect 15956 35092 15965 35132
rect 15907 35091 15965 35092
rect 16291 35132 16349 35133
rect 16291 35092 16300 35132
rect 16340 35092 16349 35132
rect 16291 35091 16349 35092
rect 16675 35132 16733 35133
rect 16675 35092 16684 35132
rect 16724 35092 16733 35132
rect 16675 35091 16733 35092
rect 17059 35132 17117 35133
rect 17059 35092 17068 35132
rect 17108 35092 17117 35132
rect 17059 35091 17117 35092
rect 19459 35132 19517 35133
rect 19459 35092 19468 35132
rect 19508 35092 19517 35132
rect 19459 35091 19517 35092
rect 19843 35132 19901 35133
rect 19843 35092 19852 35132
rect 19892 35092 19901 35132
rect 19843 35091 19901 35092
rect 1611 35048 1653 35057
rect 1611 35008 1612 35048
rect 1652 35008 1653 35048
rect 1611 34999 1653 35008
rect 16107 35048 16149 35057
rect 16107 35008 16108 35048
rect 16148 35008 16149 35048
rect 16107 34999 16149 35008
rect 16491 35048 16533 35057
rect 16491 35008 16492 35048
rect 16532 35008 16533 35048
rect 16491 34999 16533 35008
rect 16875 35048 16917 35057
rect 16875 35008 16876 35048
rect 16916 35008 16917 35048
rect 16875 34999 16917 35008
rect 17259 35048 17301 35057
rect 17259 35008 17260 35048
rect 17300 35008 17301 35048
rect 17259 34999 17301 35008
rect 9195 34964 9237 34973
rect 9195 34924 9196 34964
rect 9236 34924 9237 34964
rect 9195 34915 9237 34924
rect 10827 34964 10869 34973
rect 10827 34924 10828 34964
rect 10868 34924 10869 34964
rect 10827 34915 10869 34924
rect 12459 34964 12501 34973
rect 12459 34924 12460 34964
rect 12500 34924 12501 34964
rect 12459 34915 12501 34924
rect 14091 34964 14133 34973
rect 14091 34924 14092 34964
rect 14132 34924 14133 34964
rect 14091 34915 14133 34924
rect 14283 34964 14325 34973
rect 14283 34924 14284 34964
rect 14324 34924 14325 34964
rect 14283 34915 14325 34924
rect 19659 34964 19701 34973
rect 19659 34924 19660 34964
rect 19700 34924 19701 34964
rect 19659 34915 19701 34924
rect 20043 34964 20085 34973
rect 20043 34924 20044 34964
rect 20084 34924 20085 34964
rect 20043 34915 20085 34924
rect 1152 34796 20352 34820
rect 1152 34756 3688 34796
rect 3728 34756 3770 34796
rect 3810 34756 3852 34796
rect 3892 34756 3934 34796
rect 3974 34756 4016 34796
rect 4056 34756 18808 34796
rect 18848 34756 18890 34796
rect 18930 34756 18972 34796
rect 19012 34756 19054 34796
rect 19094 34756 19136 34796
rect 19176 34756 20352 34796
rect 1152 34732 20352 34756
rect 2955 34628 2997 34637
rect 2955 34588 2956 34628
rect 2996 34588 2997 34628
rect 2955 34579 2997 34588
rect 3139 34460 3197 34461
rect 3139 34420 3148 34460
rect 3188 34420 3197 34460
rect 3139 34419 3197 34420
rect 3915 34460 3957 34469
rect 3915 34420 3916 34460
rect 3956 34420 3957 34460
rect 3915 34411 3957 34420
rect 8427 34460 8469 34469
rect 8427 34420 8428 34460
rect 8468 34420 8469 34460
rect 8427 34411 8469 34420
rect 13803 34460 13845 34469
rect 13803 34420 13804 34460
rect 13844 34420 13845 34460
rect 13803 34411 13845 34420
rect 18595 34460 18653 34461
rect 18595 34420 18604 34460
rect 18644 34420 18653 34460
rect 18595 34419 18653 34420
rect 18979 34460 19037 34461
rect 18979 34420 18988 34460
rect 19028 34420 19037 34460
rect 18979 34419 19037 34420
rect 19363 34460 19421 34461
rect 19363 34420 19372 34460
rect 19412 34420 19421 34460
rect 19363 34419 19421 34420
rect 19747 34460 19805 34461
rect 19747 34420 19756 34460
rect 19796 34420 19805 34460
rect 19747 34419 19805 34420
rect 9483 34390 9525 34399
rect 1219 34376 1277 34377
rect 1219 34336 1228 34376
rect 1268 34336 1277 34376
rect 1219 34335 1277 34336
rect 2467 34376 2525 34377
rect 2467 34336 2476 34376
rect 2516 34336 2525 34376
rect 2467 34335 2525 34336
rect 3331 34376 3389 34377
rect 3331 34336 3340 34376
rect 3380 34336 3389 34376
rect 3331 34335 3389 34336
rect 3435 34376 3477 34385
rect 3435 34336 3436 34376
rect 3476 34336 3477 34376
rect 3435 34327 3477 34336
rect 3627 34376 3669 34385
rect 3627 34336 3628 34376
rect 3668 34336 3669 34376
rect 3627 34327 3669 34336
rect 4195 34376 4253 34377
rect 4195 34336 4204 34376
rect 4244 34336 4253 34376
rect 4195 34335 4253 34336
rect 5443 34376 5501 34377
rect 5443 34336 5452 34376
rect 5492 34336 5501 34376
rect 5443 34335 5501 34336
rect 6019 34376 6077 34377
rect 6019 34336 6028 34376
rect 6068 34336 6077 34376
rect 6019 34335 6077 34336
rect 6211 34376 6269 34377
rect 6211 34336 6220 34376
rect 6260 34336 6269 34376
rect 6211 34335 6269 34336
rect 7459 34376 7517 34377
rect 7459 34336 7468 34376
rect 7508 34336 7517 34376
rect 7459 34335 7517 34336
rect 7947 34376 7989 34385
rect 7947 34336 7948 34376
rect 7988 34336 7989 34376
rect 7947 34327 7989 34336
rect 8043 34376 8085 34385
rect 8043 34336 8044 34376
rect 8084 34336 8085 34376
rect 8043 34327 8085 34336
rect 8523 34376 8565 34385
rect 8523 34336 8524 34376
rect 8564 34336 8565 34376
rect 8523 34327 8565 34336
rect 8995 34376 9053 34377
rect 8995 34336 9004 34376
rect 9044 34336 9053 34376
rect 9483 34350 9484 34390
rect 9524 34350 9525 34390
rect 14859 34390 14901 34399
rect 9483 34341 9525 34350
rect 11011 34376 11069 34377
rect 8995 34335 9053 34336
rect 11011 34336 11020 34376
rect 11060 34336 11069 34376
rect 11011 34335 11069 34336
rect 12259 34376 12317 34377
rect 12259 34336 12268 34376
rect 12308 34336 12317 34376
rect 12259 34335 12317 34336
rect 13323 34376 13365 34385
rect 13323 34336 13324 34376
rect 13364 34336 13365 34376
rect 13323 34327 13365 34336
rect 13419 34376 13461 34385
rect 13419 34336 13420 34376
rect 13460 34336 13461 34376
rect 13419 34327 13461 34336
rect 13899 34376 13941 34385
rect 13899 34336 13900 34376
rect 13940 34336 13941 34376
rect 13899 34327 13941 34336
rect 14371 34376 14429 34377
rect 14371 34336 14380 34376
rect 14420 34336 14429 34376
rect 14859 34350 14860 34390
rect 14900 34350 14901 34390
rect 14859 34341 14901 34350
rect 15235 34376 15293 34377
rect 14371 34335 14429 34336
rect 15235 34336 15244 34376
rect 15284 34336 15293 34376
rect 15235 34335 15293 34336
rect 16483 34376 16541 34377
rect 16483 34336 16492 34376
rect 16532 34336 16541 34376
rect 16483 34335 16541 34336
rect 16867 34376 16925 34377
rect 16867 34336 16876 34376
rect 16916 34336 16925 34376
rect 16867 34335 16925 34336
rect 18115 34376 18173 34377
rect 18115 34336 18124 34376
rect 18164 34336 18173 34376
rect 18115 34335 18173 34336
rect 5643 34292 5685 34301
rect 5643 34252 5644 34292
rect 5684 34252 5685 34292
rect 5643 34243 5685 34252
rect 7659 34292 7701 34301
rect 7659 34252 7660 34292
rect 7700 34252 7701 34292
rect 7659 34243 7701 34252
rect 2667 34208 2709 34217
rect 2667 34168 2668 34208
rect 2708 34168 2709 34208
rect 2667 34159 2709 34168
rect 3523 34208 3581 34209
rect 3523 34168 3532 34208
rect 3572 34168 3581 34208
rect 3523 34167 3581 34168
rect 5931 34208 5973 34217
rect 5931 34168 5932 34208
rect 5972 34168 5973 34208
rect 5931 34159 5973 34168
rect 9675 34208 9717 34217
rect 9675 34168 9676 34208
rect 9716 34168 9717 34208
rect 9675 34159 9717 34168
rect 12459 34208 12501 34217
rect 12459 34168 12460 34208
rect 12500 34168 12501 34208
rect 12459 34159 12501 34168
rect 15051 34208 15093 34217
rect 15051 34168 15052 34208
rect 15092 34168 15093 34208
rect 15051 34159 15093 34168
rect 16683 34208 16725 34217
rect 16683 34168 16684 34208
rect 16724 34168 16725 34208
rect 16683 34159 16725 34168
rect 18315 34208 18357 34217
rect 18315 34168 18316 34208
rect 18356 34168 18357 34208
rect 18315 34159 18357 34168
rect 18795 34208 18837 34217
rect 18795 34168 18796 34208
rect 18836 34168 18837 34208
rect 18795 34159 18837 34168
rect 19179 34208 19221 34217
rect 19179 34168 19180 34208
rect 19220 34168 19221 34208
rect 19179 34159 19221 34168
rect 19563 34208 19605 34217
rect 19563 34168 19564 34208
rect 19604 34168 19605 34208
rect 19563 34159 19605 34168
rect 19947 34208 19989 34217
rect 19947 34168 19948 34208
rect 19988 34168 19989 34208
rect 19947 34159 19989 34168
rect 1152 34040 20452 34064
rect 1152 34000 4928 34040
rect 4968 34000 5010 34040
rect 5050 34000 5092 34040
rect 5132 34000 5174 34040
rect 5214 34000 5256 34040
rect 5296 34000 20048 34040
rect 20088 34000 20130 34040
rect 20170 34000 20212 34040
rect 20252 34000 20294 34040
rect 20334 34000 20376 34040
rect 20416 34000 20452 34040
rect 1152 33976 20452 34000
rect 1611 33872 1653 33881
rect 1611 33832 1612 33872
rect 1652 33832 1653 33872
rect 1611 33823 1653 33832
rect 3907 33872 3965 33873
rect 3907 33832 3916 33872
rect 3956 33832 3965 33872
rect 3907 33831 3965 33832
rect 5643 33872 5685 33881
rect 5643 33832 5644 33872
rect 5684 33832 5685 33872
rect 5643 33823 5685 33832
rect 5835 33872 5877 33881
rect 5835 33832 5836 33872
rect 5876 33832 5877 33872
rect 5835 33823 5877 33832
rect 15723 33872 15765 33881
rect 15723 33832 15724 33872
rect 15764 33832 15765 33872
rect 15723 33823 15765 33832
rect 17739 33872 17781 33881
rect 17739 33832 17740 33872
rect 17780 33832 17781 33872
rect 17739 33823 17781 33832
rect 3627 33788 3669 33797
rect 3627 33748 3628 33788
rect 3668 33748 3669 33788
rect 3627 33739 3669 33748
rect 9675 33788 9717 33797
rect 9675 33748 9676 33788
rect 9716 33748 9717 33788
rect 9675 33739 9717 33748
rect 11691 33788 11733 33797
rect 11691 33748 11692 33788
rect 11732 33748 11733 33788
rect 11691 33739 11733 33748
rect 14187 33788 14229 33797
rect 14187 33748 14188 33788
rect 14228 33748 14229 33788
rect 14187 33739 14229 33748
rect 1899 33704 1941 33713
rect 1899 33664 1900 33704
rect 1940 33664 1941 33704
rect 1899 33655 1941 33664
rect 1995 33704 2037 33713
rect 1995 33664 1996 33704
rect 2036 33664 2037 33704
rect 1995 33655 2037 33664
rect 2475 33704 2517 33713
rect 2475 33664 2476 33704
rect 2516 33664 2517 33704
rect 2475 33655 2517 33664
rect 2966 33691 3008 33700
rect 2966 33651 2967 33691
rect 3007 33651 3008 33691
rect 2966 33642 3008 33651
rect 3435 33699 3477 33708
rect 3435 33659 3436 33699
rect 3476 33659 3477 33699
rect 4195 33704 4253 33705
rect 4195 33664 4204 33704
rect 4244 33664 4253 33704
rect 4195 33663 4253 33664
rect 5443 33704 5501 33705
rect 5443 33664 5452 33704
rect 5492 33664 5501 33704
rect 5443 33663 5501 33664
rect 6019 33704 6077 33705
rect 6019 33664 6028 33704
rect 6068 33664 6077 33704
rect 6019 33663 6077 33664
rect 7267 33704 7325 33705
rect 7267 33664 7276 33704
rect 7316 33664 7325 33704
rect 7267 33663 7325 33664
rect 7467 33704 7509 33713
rect 7467 33664 7468 33704
rect 7508 33664 7509 33704
rect 3435 33650 3477 33659
rect 7467 33655 7509 33664
rect 7843 33704 7901 33705
rect 7843 33664 7852 33704
rect 7892 33664 7901 33704
rect 7843 33663 7901 33664
rect 8227 33704 8285 33705
rect 8227 33664 8236 33704
rect 8276 33664 8285 33704
rect 8227 33663 8285 33664
rect 9475 33704 9533 33705
rect 9475 33664 9484 33704
rect 9524 33664 9533 33704
rect 9475 33663 9533 33664
rect 9963 33704 10005 33713
rect 9963 33664 9964 33704
rect 10004 33664 10005 33704
rect 9963 33655 10005 33664
rect 10059 33704 10101 33713
rect 10059 33664 10060 33704
rect 10100 33664 10101 33704
rect 10059 33655 10101 33664
rect 10443 33704 10485 33713
rect 10443 33664 10444 33704
rect 10484 33664 10485 33704
rect 10443 33655 10485 33664
rect 10539 33704 10581 33713
rect 10539 33664 10540 33704
rect 10580 33664 10581 33704
rect 10539 33655 10581 33664
rect 11011 33704 11069 33705
rect 11011 33664 11020 33704
rect 11060 33664 11069 33704
rect 11011 33663 11069 33664
rect 11499 33699 11541 33708
rect 11499 33659 11500 33699
rect 11540 33659 11541 33699
rect 11499 33650 11541 33659
rect 12459 33704 12501 33713
rect 12459 33664 12460 33704
rect 12500 33664 12501 33704
rect 12459 33655 12501 33664
rect 12555 33704 12597 33713
rect 12555 33664 12556 33704
rect 12596 33664 12597 33704
rect 12555 33655 12597 33664
rect 13507 33704 13565 33705
rect 13507 33664 13516 33704
rect 13556 33664 13565 33704
rect 16011 33704 16053 33713
rect 13507 33663 13565 33664
rect 14043 33694 14085 33703
rect 14043 33654 14044 33694
rect 14084 33654 14085 33694
rect 16011 33664 16012 33704
rect 16052 33664 16053 33704
rect 16011 33655 16053 33664
rect 16107 33704 16149 33713
rect 16107 33664 16108 33704
rect 16148 33664 16149 33704
rect 16107 33655 16149 33664
rect 17059 33704 17117 33705
rect 17059 33664 17068 33704
rect 17108 33664 17117 33704
rect 17059 33663 17117 33664
rect 17547 33699 17589 33708
rect 17547 33659 17548 33699
rect 17588 33659 17589 33699
rect 14043 33645 14085 33654
rect 17547 33650 17589 33659
rect 1411 33620 1469 33621
rect 1411 33580 1420 33620
rect 1460 33580 1469 33620
rect 1411 33579 1469 33580
rect 2379 33620 2421 33629
rect 2379 33580 2380 33620
rect 2420 33580 2421 33620
rect 2379 33571 2421 33580
rect 7563 33620 7605 33629
rect 7563 33580 7564 33620
rect 7604 33580 7605 33620
rect 7563 33571 7605 33580
rect 7755 33620 7797 33629
rect 7755 33580 7756 33620
rect 7796 33580 7797 33620
rect 7755 33571 7797 33580
rect 12939 33620 12981 33629
rect 12939 33580 12940 33620
rect 12980 33580 12981 33620
rect 12939 33571 12981 33580
rect 13035 33620 13077 33629
rect 13035 33580 13036 33620
rect 13076 33580 13077 33620
rect 13035 33571 13077 33580
rect 15523 33620 15581 33621
rect 15523 33580 15532 33620
rect 15572 33580 15581 33620
rect 15523 33579 15581 33580
rect 16491 33620 16533 33629
rect 16491 33580 16492 33620
rect 16532 33580 16533 33620
rect 16491 33571 16533 33580
rect 16587 33620 16629 33629
rect 16587 33580 16588 33620
rect 16628 33580 16629 33620
rect 16587 33571 16629 33580
rect 18211 33620 18269 33621
rect 18211 33580 18220 33620
rect 18260 33580 18269 33620
rect 18211 33579 18269 33580
rect 18595 33620 18653 33621
rect 18595 33580 18604 33620
rect 18644 33580 18653 33620
rect 18595 33579 18653 33580
rect 18979 33620 19037 33621
rect 18979 33580 18988 33620
rect 19028 33580 19037 33620
rect 18979 33579 19037 33580
rect 19363 33620 19421 33621
rect 19363 33580 19372 33620
rect 19412 33580 19421 33620
rect 19363 33579 19421 33580
rect 19747 33620 19805 33621
rect 19747 33580 19756 33620
rect 19796 33580 19805 33620
rect 19747 33579 19805 33580
rect 7659 33536 7701 33545
rect 7659 33496 7660 33536
rect 7700 33496 7701 33536
rect 7659 33487 7701 33496
rect 15339 33536 15381 33545
rect 15339 33496 15340 33536
rect 15380 33496 15381 33536
rect 15339 33487 15381 33496
rect 19179 33536 19221 33545
rect 19179 33496 19180 33536
rect 19220 33496 19221 33536
rect 19179 33487 19221 33496
rect 5643 33452 5685 33461
rect 5643 33412 5644 33452
rect 5684 33412 5685 33452
rect 5643 33403 5685 33412
rect 18411 33452 18453 33461
rect 18411 33412 18412 33452
rect 18452 33412 18453 33452
rect 18411 33403 18453 33412
rect 18795 33452 18837 33461
rect 18795 33412 18796 33452
rect 18836 33412 18837 33452
rect 18795 33403 18837 33412
rect 19563 33452 19605 33461
rect 19563 33412 19564 33452
rect 19604 33412 19605 33452
rect 19563 33403 19605 33412
rect 19947 33452 19989 33461
rect 19947 33412 19948 33452
rect 19988 33412 19989 33452
rect 19947 33403 19989 33412
rect 1152 33284 20352 33308
rect 1152 33244 3688 33284
rect 3728 33244 3770 33284
rect 3810 33244 3852 33284
rect 3892 33244 3934 33284
rect 3974 33244 4016 33284
rect 4056 33244 18808 33284
rect 18848 33244 18890 33284
rect 18930 33244 18972 33284
rect 19012 33244 19054 33284
rect 19094 33244 19136 33284
rect 19176 33244 20352 33284
rect 1152 33220 20352 33244
rect 1515 33116 1557 33125
rect 1515 33076 1516 33116
rect 1556 33076 1557 33116
rect 1515 33067 1557 33076
rect 1899 33116 1941 33125
rect 1899 33076 1900 33116
rect 1940 33076 1941 33116
rect 1899 33067 1941 33076
rect 5451 33116 5493 33125
rect 5451 33076 5452 33116
rect 5492 33076 5493 33116
rect 5451 33067 5493 33076
rect 5827 33116 5885 33117
rect 5827 33076 5836 33116
rect 5876 33076 5885 33116
rect 5827 33075 5885 33076
rect 7083 33116 7125 33125
rect 7083 33076 7084 33116
rect 7124 33076 7125 33116
rect 7083 33067 7125 33076
rect 19563 33116 19605 33125
rect 19563 33076 19564 33116
rect 19604 33076 19605 33116
rect 19563 33067 19605 33076
rect 2283 33032 2325 33041
rect 2283 32992 2284 33032
rect 2324 32992 2325 33032
rect 2283 32983 2325 32992
rect 19947 33032 19989 33041
rect 19947 32992 19948 33032
rect 19988 32992 19989 33032
rect 19947 32983 19989 32992
rect 1315 32948 1373 32949
rect 1315 32908 1324 32948
rect 1364 32908 1373 32948
rect 1315 32907 1373 32908
rect 1699 32948 1757 32949
rect 1699 32908 1708 32948
rect 1748 32908 1757 32948
rect 1699 32907 1757 32908
rect 11883 32948 11925 32957
rect 11883 32908 11884 32948
rect 11924 32908 11925 32948
rect 11883 32899 11925 32908
rect 17739 32948 17781 32957
rect 17739 32908 17740 32948
rect 17780 32908 17781 32948
rect 17739 32899 17781 32908
rect 19363 32948 19421 32949
rect 19363 32908 19372 32948
rect 19412 32908 19421 32948
rect 19363 32907 19421 32908
rect 19747 32948 19805 32949
rect 19747 32908 19756 32948
rect 19796 32908 19805 32948
rect 19747 32907 19805 32908
rect 18747 32873 18789 32882
rect 2467 32864 2525 32865
rect 2467 32824 2476 32864
rect 2516 32824 2525 32864
rect 2467 32823 2525 32824
rect 3715 32864 3773 32865
rect 3715 32824 3724 32864
rect 3764 32824 3773 32864
rect 3715 32823 3773 32824
rect 4003 32864 4061 32865
rect 4003 32824 4012 32864
rect 4052 32824 4061 32864
rect 4003 32823 4061 32824
rect 5251 32864 5309 32865
rect 5251 32824 5260 32864
rect 5300 32824 5309 32864
rect 5251 32823 5309 32824
rect 6219 32864 6261 32873
rect 6219 32824 6220 32864
rect 6260 32824 6261 32864
rect 6219 32815 6261 32824
rect 6499 32864 6557 32865
rect 6499 32824 6508 32864
rect 6548 32824 6557 32864
rect 6499 32823 6557 32824
rect 6787 32864 6845 32865
rect 6787 32824 6796 32864
rect 6836 32824 6845 32864
rect 6787 32823 6845 32824
rect 6891 32864 6933 32873
rect 6891 32824 6892 32864
rect 6932 32824 6933 32864
rect 6891 32815 6933 32824
rect 7083 32864 7125 32873
rect 7083 32824 7084 32864
rect 7124 32824 7125 32864
rect 7083 32815 7125 32824
rect 7275 32864 7317 32873
rect 7275 32824 7276 32864
rect 7316 32824 7317 32864
rect 7275 32815 7317 32824
rect 7467 32864 7509 32873
rect 7467 32824 7468 32864
rect 7508 32824 7509 32864
rect 7467 32815 7509 32824
rect 7555 32864 7613 32865
rect 7555 32824 7564 32864
rect 7604 32824 7613 32864
rect 7555 32823 7613 32824
rect 7747 32864 7805 32865
rect 7747 32824 7756 32864
rect 7796 32824 7805 32864
rect 7747 32823 7805 32824
rect 7851 32864 7893 32873
rect 7851 32824 7852 32864
rect 7892 32824 7893 32864
rect 7851 32815 7893 32824
rect 8035 32864 8093 32865
rect 8035 32824 8044 32864
rect 8084 32824 8093 32864
rect 8035 32823 8093 32824
rect 9283 32864 9341 32865
rect 9283 32824 9292 32864
rect 9332 32824 9341 32864
rect 9283 32823 9341 32824
rect 10147 32864 10205 32865
rect 10147 32824 10156 32864
rect 10196 32824 10205 32864
rect 10147 32823 10205 32824
rect 11395 32864 11453 32865
rect 11395 32824 11404 32864
rect 11444 32824 11453 32864
rect 11395 32823 11453 32824
rect 12651 32864 12693 32873
rect 12651 32824 12652 32864
rect 12692 32824 12693 32864
rect 12651 32815 12693 32824
rect 13315 32864 13373 32865
rect 13315 32824 13324 32864
rect 13364 32824 13373 32864
rect 13315 32823 13373 32824
rect 14563 32864 14621 32865
rect 14563 32824 14572 32864
rect 14612 32824 14621 32864
rect 14563 32823 14621 32824
rect 15427 32864 15485 32865
rect 15427 32824 15436 32864
rect 15476 32824 15485 32864
rect 15427 32823 15485 32824
rect 16675 32864 16733 32865
rect 16675 32824 16684 32864
rect 16724 32824 16733 32864
rect 16675 32823 16733 32824
rect 17163 32864 17205 32873
rect 17163 32824 17164 32864
rect 17204 32824 17205 32864
rect 17163 32815 17205 32824
rect 17259 32864 17301 32873
rect 17259 32824 17260 32864
rect 17300 32824 17301 32864
rect 17259 32815 17301 32824
rect 17643 32864 17685 32873
rect 17643 32824 17644 32864
rect 17684 32824 17685 32864
rect 17643 32815 17685 32824
rect 18211 32864 18269 32865
rect 18211 32824 18220 32864
rect 18260 32824 18269 32864
rect 18747 32833 18748 32873
rect 18788 32833 18789 32873
rect 18747 32824 18789 32833
rect 18211 32823 18269 32824
rect 6123 32780 6165 32789
rect 6123 32740 6124 32780
rect 6164 32740 6165 32780
rect 6123 32731 6165 32740
rect 7371 32780 7413 32789
rect 7371 32740 7372 32780
rect 7412 32740 7413 32780
rect 7371 32731 7413 32740
rect 16875 32780 16917 32789
rect 16875 32740 16876 32780
rect 16916 32740 16917 32780
rect 16875 32731 16917 32740
rect 18891 32780 18933 32789
rect 18891 32740 18892 32780
rect 18932 32740 18933 32780
rect 18891 32731 18933 32740
rect 9483 32696 9525 32705
rect 9483 32656 9484 32696
rect 9524 32656 9525 32696
rect 9483 32647 9525 32656
rect 11595 32696 11637 32705
rect 11595 32656 11596 32696
rect 11636 32656 11637 32696
rect 11595 32647 11637 32656
rect 14763 32696 14805 32705
rect 14763 32656 14764 32696
rect 14804 32656 14805 32696
rect 14763 32647 14805 32656
rect 1152 32528 20452 32552
rect 1152 32488 4928 32528
rect 4968 32488 5010 32528
rect 5050 32488 5092 32528
rect 5132 32488 5174 32528
rect 5214 32488 5256 32528
rect 5296 32488 20048 32528
rect 20088 32488 20130 32528
rect 20170 32488 20212 32528
rect 20252 32488 20294 32528
rect 20334 32488 20376 32528
rect 20416 32488 20452 32528
rect 1152 32464 20452 32488
rect 2763 32360 2805 32369
rect 2763 32320 2764 32360
rect 2804 32320 2805 32360
rect 2763 32311 2805 32320
rect 4779 32360 4821 32369
rect 4779 32320 4780 32360
rect 4820 32320 4821 32360
rect 4779 32311 4821 32320
rect 7851 32360 7893 32369
rect 7851 32320 7852 32360
rect 7892 32320 7893 32360
rect 7851 32311 7893 32320
rect 8323 32360 8381 32361
rect 8323 32320 8332 32360
rect 8372 32320 8381 32360
rect 8323 32319 8381 32320
rect 16491 32360 16533 32369
rect 16491 32320 16492 32360
rect 16532 32320 16533 32360
rect 16491 32311 16533 32320
rect 16875 32360 16917 32369
rect 16875 32320 16876 32360
rect 16916 32320 16917 32360
rect 16875 32311 16917 32320
rect 17259 32360 17301 32369
rect 17259 32320 17260 32360
rect 17300 32320 17301 32360
rect 17259 32311 17301 32320
rect 18891 32360 18933 32369
rect 18891 32320 18892 32360
rect 18932 32320 18933 32360
rect 18891 32311 18933 32320
rect 6891 32276 6933 32285
rect 6891 32236 6892 32276
rect 6932 32236 6933 32276
rect 6891 32227 6933 32236
rect 12171 32276 12213 32285
rect 12171 32236 12172 32276
rect 12212 32236 12213 32276
rect 12171 32227 12213 32236
rect 14187 32276 14229 32285
rect 14187 32236 14188 32276
rect 14228 32236 14229 32276
rect 14187 32227 14229 32236
rect 2955 32187 2997 32196
rect 2955 32147 2956 32187
rect 2996 32147 2997 32187
rect 3427 32192 3485 32193
rect 3427 32152 3436 32192
rect 3476 32152 3485 32192
rect 3427 32151 3485 32152
rect 4395 32192 4437 32201
rect 4395 32152 4396 32192
rect 4436 32152 4437 32192
rect 2955 32138 2997 32147
rect 4395 32143 4437 32152
rect 4491 32192 4533 32201
rect 4491 32152 4492 32192
rect 4532 32152 4533 32192
rect 4491 32143 4533 32152
rect 4963 32192 5021 32193
rect 4963 32152 4972 32192
rect 5012 32152 5021 32192
rect 4963 32151 5021 32152
rect 6211 32192 6269 32193
rect 6211 32152 6220 32192
rect 6260 32152 6269 32192
rect 6211 32151 6269 32152
rect 6499 32192 6557 32193
rect 6499 32152 6508 32192
rect 6548 32152 6557 32192
rect 6499 32151 6557 32152
rect 6795 32192 6837 32201
rect 6795 32152 6796 32192
rect 6836 32152 6837 32192
rect 6795 32143 6837 32152
rect 7659 32192 7701 32201
rect 7659 32152 7660 32192
rect 7700 32152 7701 32192
rect 8139 32192 8181 32201
rect 7659 32143 7701 32152
rect 8043 32147 8085 32156
rect 3915 32108 3957 32117
rect 3915 32068 3916 32108
rect 3956 32068 3957 32108
rect 3915 32059 3957 32068
rect 4011 32108 4053 32117
rect 4011 32068 4012 32108
rect 4052 32068 4053 32108
rect 8043 32107 8044 32147
rect 8084 32107 8085 32147
rect 8139 32152 8140 32192
rect 8180 32152 8181 32192
rect 8139 32143 8181 32152
rect 8235 32192 8277 32201
rect 8235 32152 8236 32192
rect 8276 32152 8277 32192
rect 8235 32143 8277 32152
rect 8611 32192 8669 32193
rect 8611 32152 8620 32192
rect 8660 32152 8669 32192
rect 8611 32151 8669 32152
rect 9859 32192 9917 32193
rect 9859 32152 9868 32192
rect 9908 32152 9917 32192
rect 9859 32151 9917 32152
rect 10723 32192 10781 32193
rect 10723 32152 10732 32192
rect 10772 32152 10781 32192
rect 10723 32151 10781 32152
rect 11971 32192 12029 32193
rect 11971 32152 11980 32192
rect 12020 32152 12029 32192
rect 11971 32151 12029 32152
rect 12459 32192 12501 32201
rect 12459 32152 12460 32192
rect 12500 32152 12501 32192
rect 12459 32143 12501 32152
rect 12555 32192 12597 32201
rect 12555 32152 12556 32192
rect 12596 32152 12597 32192
rect 12555 32143 12597 32152
rect 13507 32192 13565 32193
rect 13507 32152 13516 32192
rect 13556 32152 13565 32192
rect 14763 32192 14805 32201
rect 13507 32151 13565 32152
rect 13995 32178 14037 32187
rect 13995 32138 13996 32178
rect 14036 32138 14037 32178
rect 14763 32152 14764 32192
rect 14804 32152 14805 32192
rect 14763 32143 14805 32152
rect 14859 32192 14901 32201
rect 14859 32152 14860 32192
rect 14900 32152 14901 32192
rect 14859 32143 14901 32152
rect 15243 32192 15285 32201
rect 15243 32152 15244 32192
rect 15284 32152 15285 32192
rect 15243 32143 15285 32152
rect 15339 32192 15381 32201
rect 15339 32152 15340 32192
rect 15380 32152 15381 32192
rect 15339 32143 15381 32152
rect 15811 32192 15869 32193
rect 15811 32152 15820 32192
rect 15860 32152 15869 32192
rect 17443 32192 17501 32193
rect 15811 32151 15869 32152
rect 16299 32178 16341 32187
rect 13995 32129 14037 32138
rect 16299 32138 16300 32178
rect 16340 32138 16341 32178
rect 17443 32152 17452 32192
rect 17492 32152 17501 32192
rect 17443 32151 17501 32152
rect 18691 32192 18749 32193
rect 18691 32152 18700 32192
rect 18740 32152 18749 32192
rect 18691 32151 18749 32152
rect 16299 32129 16341 32138
rect 8043 32098 8085 32107
rect 12939 32108 12981 32117
rect 4011 32059 4053 32068
rect 12939 32068 12940 32108
rect 12980 32068 12981 32108
rect 12939 32059 12981 32068
rect 13035 32108 13077 32117
rect 13035 32068 13036 32108
rect 13076 32068 13077 32108
rect 13035 32059 13077 32068
rect 16675 32108 16733 32109
rect 16675 32068 16684 32108
rect 16724 32068 16733 32108
rect 16675 32067 16733 32068
rect 17059 32108 17117 32109
rect 17059 32068 17068 32108
rect 17108 32068 17117 32108
rect 17059 32067 17117 32068
rect 19363 32108 19421 32109
rect 19363 32068 19372 32108
rect 19412 32068 19421 32108
rect 19363 32067 19421 32068
rect 19747 32108 19805 32109
rect 19747 32068 19756 32108
rect 19796 32068 19805 32108
rect 19747 32067 19805 32068
rect 7171 32024 7229 32025
rect 7171 31984 7180 32024
rect 7220 31984 7229 32024
rect 7171 31983 7229 31984
rect 7659 32024 7701 32033
rect 7659 31984 7660 32024
rect 7700 31984 7701 32024
rect 7659 31975 7701 31984
rect 10059 31940 10101 31949
rect 10059 31900 10060 31940
rect 10100 31900 10101 31940
rect 10059 31891 10101 31900
rect 19563 31940 19605 31949
rect 19563 31900 19564 31940
rect 19604 31900 19605 31940
rect 19563 31891 19605 31900
rect 19947 31940 19989 31949
rect 19947 31900 19948 31940
rect 19988 31900 19989 31940
rect 19947 31891 19989 31900
rect 1152 31772 20352 31796
rect 1152 31732 3688 31772
rect 3728 31732 3770 31772
rect 3810 31732 3852 31772
rect 3892 31732 3934 31772
rect 3974 31732 4016 31772
rect 4056 31732 18808 31772
rect 18848 31732 18890 31772
rect 18930 31732 18972 31772
rect 19012 31732 19054 31772
rect 19094 31732 19136 31772
rect 19176 31732 20352 31772
rect 1152 31708 20352 31732
rect 13995 31604 14037 31613
rect 13995 31564 13996 31604
rect 14036 31564 14037 31604
rect 13995 31555 14037 31564
rect 16299 31604 16341 31613
rect 16299 31564 16300 31604
rect 16340 31564 16341 31604
rect 16299 31555 16341 31564
rect 8235 31436 8277 31445
rect 8235 31396 8236 31436
rect 8276 31396 8277 31436
rect 8235 31387 8277 31396
rect 10635 31436 10677 31445
rect 10635 31396 10636 31436
rect 10676 31396 10677 31436
rect 10635 31387 10677 31396
rect 20035 31436 20093 31437
rect 20035 31396 20044 31436
rect 20084 31396 20093 31436
rect 20035 31395 20093 31396
rect 9339 31361 9381 31370
rect 11595 31366 11637 31375
rect 1219 31352 1277 31353
rect 1219 31312 1228 31352
rect 1268 31312 1277 31352
rect 1219 31311 1277 31312
rect 2467 31352 2525 31353
rect 2467 31312 2476 31352
rect 2516 31312 2525 31352
rect 2467 31311 2525 31312
rect 3043 31352 3101 31353
rect 3043 31312 3052 31352
rect 3092 31312 3101 31352
rect 3043 31311 3101 31312
rect 4195 31352 4253 31353
rect 4195 31312 4204 31352
rect 4244 31312 4253 31352
rect 4195 31311 4253 31312
rect 4387 31352 4445 31353
rect 4387 31312 4396 31352
rect 4436 31312 4445 31352
rect 4387 31311 4445 31312
rect 5635 31352 5693 31353
rect 5635 31312 5644 31352
rect 5684 31312 5693 31352
rect 5635 31311 5693 31312
rect 6019 31352 6077 31353
rect 6019 31312 6028 31352
rect 6068 31312 6077 31352
rect 6019 31311 6077 31312
rect 7267 31352 7325 31353
rect 7267 31312 7276 31352
rect 7316 31312 7325 31352
rect 7267 31311 7325 31312
rect 7755 31352 7797 31361
rect 7755 31312 7756 31352
rect 7796 31312 7797 31352
rect 7755 31303 7797 31312
rect 7851 31352 7893 31361
rect 7851 31312 7852 31352
rect 7892 31312 7893 31352
rect 7851 31303 7893 31312
rect 8331 31352 8373 31361
rect 8331 31312 8332 31352
rect 8372 31312 8373 31352
rect 8331 31303 8373 31312
rect 8803 31352 8861 31353
rect 8803 31312 8812 31352
rect 8852 31312 8861 31352
rect 9339 31321 9340 31361
rect 9380 31321 9381 31361
rect 9339 31312 9381 31321
rect 10059 31352 10101 31361
rect 10059 31312 10060 31352
rect 10100 31312 10101 31352
rect 8803 31311 8861 31312
rect 10059 31303 10101 31312
rect 10155 31352 10197 31361
rect 10155 31312 10156 31352
rect 10196 31312 10197 31352
rect 10155 31303 10197 31312
rect 10539 31352 10581 31361
rect 10539 31312 10540 31352
rect 10580 31312 10581 31352
rect 10539 31303 10581 31312
rect 11107 31352 11165 31353
rect 11107 31312 11116 31352
rect 11156 31312 11165 31352
rect 11595 31326 11596 31366
rect 11636 31326 11637 31366
rect 11595 31317 11637 31326
rect 12547 31352 12605 31353
rect 11107 31311 11165 31312
rect 12547 31312 12556 31352
rect 12596 31312 12605 31352
rect 12547 31311 12605 31312
rect 13795 31352 13853 31353
rect 13795 31312 13804 31352
rect 13844 31312 13853 31352
rect 13795 31311 13853 31312
rect 14851 31352 14909 31353
rect 14851 31312 14860 31352
rect 14900 31312 14909 31352
rect 14851 31311 14909 31312
rect 16099 31352 16157 31353
rect 16099 31312 16108 31352
rect 16148 31312 16157 31352
rect 16099 31311 16157 31312
rect 16483 31352 16541 31353
rect 16483 31312 16492 31352
rect 16532 31312 16541 31352
rect 16483 31311 16541 31312
rect 17731 31352 17789 31353
rect 17731 31312 17740 31352
rect 17780 31312 17789 31352
rect 17731 31311 17789 31312
rect 18403 31352 18461 31353
rect 18403 31312 18412 31352
rect 18452 31312 18461 31352
rect 18403 31311 18461 31312
rect 19651 31352 19709 31353
rect 19651 31312 19660 31352
rect 19700 31312 19709 31352
rect 19651 31311 19709 31312
rect 7467 31268 7509 31277
rect 7467 31228 7468 31268
rect 7508 31228 7509 31268
rect 7467 31219 7509 31228
rect 2667 31184 2709 31193
rect 2667 31144 2668 31184
rect 2708 31144 2709 31184
rect 2667 31135 2709 31144
rect 3147 31184 3189 31193
rect 3147 31144 3148 31184
rect 3188 31144 3189 31184
rect 3147 31135 3189 31144
rect 4107 31184 4149 31193
rect 4107 31144 4108 31184
rect 4148 31144 4149 31184
rect 4107 31135 4149 31144
rect 5835 31184 5877 31193
rect 5835 31144 5836 31184
rect 5876 31144 5877 31184
rect 5835 31135 5877 31144
rect 9483 31184 9525 31193
rect 9483 31144 9484 31184
rect 9524 31144 9525 31184
rect 9483 31135 9525 31144
rect 11787 31184 11829 31193
rect 11787 31144 11788 31184
rect 11828 31144 11829 31184
rect 11787 31135 11829 31144
rect 17931 31184 17973 31193
rect 17931 31144 17932 31184
rect 17972 31144 17973 31184
rect 17931 31135 17973 31144
rect 19851 31184 19893 31193
rect 19851 31144 19852 31184
rect 19892 31144 19893 31184
rect 19851 31135 19893 31144
rect 20235 31184 20277 31193
rect 20235 31144 20236 31184
rect 20276 31144 20277 31184
rect 20235 31135 20277 31144
rect 1152 31016 20452 31040
rect 1152 30976 4928 31016
rect 4968 30976 5010 31016
rect 5050 30976 5092 31016
rect 5132 30976 5174 31016
rect 5214 30976 5256 31016
rect 5296 30976 20048 31016
rect 20088 30976 20130 31016
rect 20170 30976 20212 31016
rect 20252 30976 20294 31016
rect 20334 30976 20376 31016
rect 20416 30976 20452 31016
rect 1152 30952 20452 30976
rect 6595 30848 6653 30849
rect 6595 30808 6604 30848
rect 6644 30808 6653 30848
rect 6595 30807 6653 30808
rect 7083 30848 7125 30857
rect 7083 30808 7084 30848
rect 7124 30808 7125 30848
rect 7083 30799 7125 30808
rect 7467 30848 7509 30857
rect 7467 30808 7468 30848
rect 7508 30808 7509 30848
rect 7467 30799 7509 30808
rect 19467 30848 19509 30857
rect 19467 30808 19468 30848
rect 19508 30808 19509 30848
rect 19467 30799 19509 30808
rect 4107 30764 4149 30773
rect 4107 30724 4108 30764
rect 4148 30724 4149 30764
rect 4107 30715 4149 30724
rect 6123 30764 6165 30773
rect 6123 30724 6124 30764
rect 6164 30724 6165 30764
rect 6123 30715 6165 30724
rect 2187 30680 2229 30689
rect 2187 30640 2188 30680
rect 2228 30640 2229 30680
rect 2187 30631 2229 30640
rect 2379 30680 2421 30689
rect 2379 30640 2380 30680
rect 2420 30640 2421 30680
rect 2379 30631 2421 30640
rect 2475 30680 2517 30689
rect 2475 30640 2476 30680
rect 2516 30640 2517 30680
rect 2475 30631 2517 30640
rect 2659 30680 2717 30681
rect 2659 30640 2668 30680
rect 2708 30640 2717 30680
rect 2659 30639 2717 30640
rect 3907 30680 3965 30681
rect 3907 30640 3916 30680
rect 3956 30640 3965 30680
rect 3907 30639 3965 30640
rect 4395 30680 4437 30689
rect 4395 30640 4396 30680
rect 4436 30640 4437 30680
rect 4395 30631 4437 30640
rect 4491 30680 4533 30689
rect 4491 30640 4492 30680
rect 4532 30640 4533 30680
rect 4491 30631 4533 30640
rect 4875 30680 4917 30689
rect 4875 30640 4876 30680
rect 4916 30640 4917 30680
rect 4875 30631 4917 30640
rect 4971 30680 5013 30689
rect 4971 30640 4972 30680
rect 5012 30640 5013 30680
rect 4971 30631 5013 30640
rect 5443 30680 5501 30681
rect 5443 30640 5452 30680
rect 5492 30640 5501 30680
rect 5443 30639 5501 30640
rect 5931 30675 5973 30684
rect 5931 30635 5932 30675
rect 5972 30635 5973 30675
rect 5931 30626 5973 30635
rect 6315 30680 6357 30689
rect 6315 30640 6316 30680
rect 6356 30640 6357 30680
rect 6315 30631 6357 30640
rect 6411 30680 6453 30689
rect 6411 30640 6412 30680
rect 6452 30640 6453 30680
rect 6411 30631 6453 30640
rect 6507 30680 6549 30689
rect 6507 30640 6508 30680
rect 6548 30640 6549 30680
rect 6507 30631 6549 30640
rect 6987 30680 7029 30689
rect 6987 30640 6988 30680
rect 7028 30640 7029 30680
rect 6987 30631 7029 30640
rect 7179 30680 7221 30689
rect 7179 30640 7180 30680
rect 7220 30640 7221 30680
rect 7179 30631 7221 30640
rect 7363 30680 7421 30681
rect 7363 30640 7372 30680
rect 7412 30640 7421 30680
rect 7363 30639 7421 30640
rect 8899 30680 8957 30681
rect 8899 30640 8908 30680
rect 8948 30640 8957 30680
rect 8899 30639 8957 30640
rect 10147 30680 10205 30681
rect 10147 30640 10156 30680
rect 10196 30640 10205 30680
rect 10147 30639 10205 30640
rect 10819 30680 10877 30681
rect 10819 30640 10828 30680
rect 10868 30640 10877 30680
rect 10819 30639 10877 30640
rect 12067 30680 12125 30681
rect 12067 30640 12076 30680
rect 12116 30640 12125 30680
rect 12067 30639 12125 30640
rect 12451 30680 12509 30681
rect 12451 30640 12460 30680
rect 12500 30640 12509 30680
rect 12451 30639 12509 30640
rect 13699 30680 13757 30681
rect 13699 30640 13708 30680
rect 13748 30640 13757 30680
rect 13699 30639 13757 30640
rect 14083 30680 14141 30681
rect 14083 30640 14092 30680
rect 14132 30640 14141 30680
rect 14083 30639 14141 30640
rect 15331 30680 15389 30681
rect 15331 30640 15340 30680
rect 15380 30640 15389 30680
rect 15331 30639 15389 30640
rect 15715 30680 15773 30681
rect 15715 30640 15724 30680
rect 15764 30640 15773 30680
rect 15715 30639 15773 30640
rect 16963 30680 17021 30681
rect 16963 30640 16972 30680
rect 17012 30640 17021 30680
rect 16963 30639 17021 30640
rect 17739 30680 17781 30689
rect 17739 30640 17740 30680
rect 17780 30640 17781 30680
rect 17739 30631 17781 30640
rect 17835 30680 17877 30689
rect 17835 30640 17836 30680
rect 17876 30640 17877 30680
rect 17835 30631 17877 30640
rect 18219 30680 18261 30689
rect 18219 30640 18220 30680
rect 18260 30640 18261 30680
rect 18219 30631 18261 30640
rect 18315 30680 18357 30689
rect 18315 30640 18316 30680
rect 18356 30640 18357 30680
rect 18315 30631 18357 30640
rect 18787 30680 18845 30681
rect 18787 30640 18796 30680
rect 18836 30640 18845 30680
rect 18787 30639 18845 30640
rect 19275 30675 19317 30684
rect 19275 30635 19276 30675
rect 19316 30635 19317 30675
rect 19275 30626 19317 30635
rect 19651 30596 19709 30597
rect 19651 30556 19660 30596
rect 19700 30556 19709 30596
rect 19651 30555 19709 30556
rect 20035 30596 20093 30597
rect 20035 30556 20044 30596
rect 20084 30556 20093 30596
rect 20035 30555 20093 30556
rect 2283 30512 2325 30521
rect 2283 30472 2284 30512
rect 2324 30472 2325 30512
rect 2283 30463 2325 30472
rect 10347 30428 10389 30437
rect 10347 30388 10348 30428
rect 10388 30388 10389 30428
rect 10347 30379 10389 30388
rect 12267 30428 12309 30437
rect 12267 30388 12268 30428
rect 12308 30388 12309 30428
rect 12267 30379 12309 30388
rect 13899 30428 13941 30437
rect 13899 30388 13900 30428
rect 13940 30388 13941 30428
rect 13899 30379 13941 30388
rect 15531 30428 15573 30437
rect 15531 30388 15532 30428
rect 15572 30388 15573 30428
rect 15531 30379 15573 30388
rect 17163 30428 17205 30437
rect 17163 30388 17164 30428
rect 17204 30388 17205 30428
rect 17163 30379 17205 30388
rect 19851 30428 19893 30437
rect 19851 30388 19852 30428
rect 19892 30388 19893 30428
rect 19851 30379 19893 30388
rect 20235 30428 20277 30437
rect 20235 30388 20236 30428
rect 20276 30388 20277 30428
rect 20235 30379 20277 30388
rect 1152 30260 20352 30284
rect 1152 30220 3688 30260
rect 3728 30220 3770 30260
rect 3810 30220 3852 30260
rect 3892 30220 3934 30260
rect 3974 30220 4016 30260
rect 4056 30220 18808 30260
rect 18848 30220 18890 30260
rect 18930 30220 18972 30260
rect 19012 30220 19054 30260
rect 19094 30220 19136 30260
rect 19176 30220 20352 30260
rect 1152 30196 20352 30220
rect 16683 30092 16725 30101
rect 16683 30052 16684 30092
rect 16724 30052 16725 30092
rect 16683 30043 16725 30052
rect 2667 30008 2709 30017
rect 2667 29968 2668 30008
rect 2708 29968 2709 30008
rect 2667 29959 2709 29968
rect 16299 30008 16341 30017
rect 16299 29968 16300 30008
rect 16340 29968 16341 30008
rect 16299 29959 16341 29968
rect 7371 29924 7413 29933
rect 7371 29884 7372 29924
rect 7412 29884 7413 29924
rect 7371 29875 7413 29884
rect 7467 29924 7509 29933
rect 7467 29884 7468 29924
rect 7508 29884 7509 29924
rect 7467 29875 7509 29884
rect 11019 29924 11061 29933
rect 11019 29884 11020 29924
rect 11060 29884 11061 29924
rect 16099 29924 16157 29925
rect 11019 29875 11061 29884
rect 15483 29882 15525 29891
rect 16099 29884 16108 29924
rect 16148 29884 16157 29924
rect 16099 29883 16157 29884
rect 16483 29924 16541 29925
rect 16483 29884 16492 29924
rect 16532 29884 16541 29924
rect 16483 29883 16541 29884
rect 17643 29924 17685 29933
rect 17643 29884 17644 29924
rect 17684 29884 17685 29924
rect 11979 29854 12021 29863
rect 1219 29840 1277 29841
rect 1219 29800 1228 29840
rect 1268 29800 1277 29840
rect 1219 29799 1277 29800
rect 2467 29840 2525 29841
rect 2467 29800 2476 29840
rect 2516 29800 2525 29840
rect 2467 29799 2525 29800
rect 2851 29840 2909 29841
rect 2851 29800 2860 29840
rect 2900 29800 2909 29840
rect 2851 29799 2909 29800
rect 2947 29840 3005 29841
rect 2947 29800 2956 29840
rect 2996 29800 3005 29840
rect 2947 29799 3005 29800
rect 3147 29840 3189 29849
rect 3147 29800 3148 29840
rect 3188 29800 3189 29840
rect 3147 29791 3189 29800
rect 3243 29840 3285 29849
rect 3243 29800 3244 29840
rect 3284 29800 3285 29840
rect 3243 29791 3285 29800
rect 3336 29840 3394 29841
rect 3336 29800 3345 29840
rect 3385 29800 3394 29840
rect 3336 29799 3394 29800
rect 3627 29840 3669 29849
rect 3627 29800 3628 29840
rect 3668 29800 3669 29840
rect 3627 29791 3669 29800
rect 3723 29840 3765 29849
rect 3723 29800 3724 29840
rect 3764 29800 3765 29840
rect 3723 29791 3765 29800
rect 5155 29840 5213 29841
rect 5155 29800 5164 29840
rect 5204 29800 5213 29840
rect 5155 29799 5213 29800
rect 6403 29840 6461 29841
rect 6403 29800 6412 29840
rect 6452 29800 6461 29840
rect 6403 29799 6461 29800
rect 6891 29840 6933 29849
rect 6891 29800 6892 29840
rect 6932 29800 6933 29840
rect 6891 29791 6933 29800
rect 6987 29840 7029 29849
rect 8427 29845 8469 29854
rect 6987 29800 6988 29840
rect 7028 29800 7029 29840
rect 6987 29791 7029 29800
rect 7939 29840 7997 29841
rect 7939 29800 7948 29840
rect 7988 29800 7997 29840
rect 7939 29799 7997 29800
rect 8427 29805 8428 29845
rect 8468 29805 8469 29845
rect 8427 29796 8469 29805
rect 8803 29840 8861 29841
rect 8803 29800 8812 29840
rect 8852 29800 8861 29840
rect 8803 29799 8861 29800
rect 9763 29840 9821 29841
rect 9763 29800 9772 29840
rect 9812 29800 9821 29840
rect 9763 29799 9821 29800
rect 10443 29840 10485 29849
rect 10443 29800 10444 29840
rect 10484 29800 10485 29840
rect 10443 29791 10485 29800
rect 10539 29840 10581 29849
rect 10539 29800 10540 29840
rect 10580 29800 10581 29840
rect 10539 29791 10581 29800
rect 10923 29840 10965 29849
rect 10923 29800 10924 29840
rect 10964 29800 10965 29840
rect 10923 29791 10965 29800
rect 11491 29840 11549 29841
rect 11491 29800 11500 29840
rect 11540 29800 11549 29840
rect 11979 29814 11980 29854
rect 12020 29814 12021 29854
rect 11979 29805 12021 29814
rect 13899 29840 13941 29849
rect 11491 29799 11549 29800
rect 13899 29800 13900 29840
rect 13940 29800 13941 29840
rect 13899 29791 13941 29800
rect 13995 29840 14037 29849
rect 13995 29800 13996 29840
rect 14036 29800 14037 29840
rect 13995 29791 14037 29800
rect 14379 29840 14421 29849
rect 14379 29800 14380 29840
rect 14420 29800 14421 29840
rect 14379 29791 14421 29800
rect 14475 29840 14517 29849
rect 15483 29842 15484 29882
rect 15524 29842 15525 29882
rect 17643 29875 17685 29884
rect 19363 29924 19421 29925
rect 19363 29884 19372 29924
rect 19412 29884 19421 29924
rect 19363 29883 19421 29884
rect 19747 29924 19805 29925
rect 19747 29884 19756 29924
rect 19796 29884 19805 29924
rect 19747 29883 19805 29884
rect 18210 29882 18268 29883
rect 14475 29800 14476 29840
rect 14516 29800 14517 29840
rect 14475 29791 14517 29800
rect 14947 29840 15005 29841
rect 14947 29800 14956 29840
rect 14996 29800 15005 29840
rect 15483 29833 15525 29842
rect 17163 29840 17205 29849
rect 14947 29799 15005 29800
rect 17163 29800 17164 29840
rect 17204 29800 17205 29840
rect 17163 29791 17205 29800
rect 17259 29840 17301 29849
rect 17259 29800 17260 29840
rect 17300 29800 17301 29840
rect 17259 29791 17301 29800
rect 17739 29840 17781 29849
rect 18210 29842 18219 29882
rect 18259 29842 18268 29882
rect 18210 29841 18268 29842
rect 18699 29845 18741 29854
rect 17739 29800 17740 29840
rect 17780 29800 17781 29840
rect 17739 29791 17781 29800
rect 18699 29805 18700 29845
rect 18740 29805 18741 29845
rect 18699 29796 18741 29805
rect 6603 29756 6645 29765
rect 6603 29716 6604 29756
rect 6644 29716 6645 29756
rect 6603 29707 6645 29716
rect 8619 29756 8661 29765
rect 8619 29716 8620 29756
rect 8660 29716 8661 29756
rect 8619 29707 8661 29716
rect 12171 29756 12213 29765
rect 12171 29716 12172 29756
rect 12212 29716 12213 29756
rect 12171 29707 12213 29716
rect 15627 29756 15669 29765
rect 15627 29716 15628 29756
rect 15668 29716 15669 29756
rect 15627 29707 15669 29716
rect 18891 29756 18933 29765
rect 18891 29716 18892 29756
rect 18932 29716 18933 29756
rect 18891 29707 18933 29716
rect 3043 29672 3101 29673
rect 3043 29632 3052 29672
rect 3092 29632 3101 29672
rect 3043 29631 3101 29632
rect 3907 29672 3965 29673
rect 3907 29632 3916 29672
rect 3956 29632 3965 29672
rect 3907 29631 3965 29632
rect 19563 29672 19605 29681
rect 19563 29632 19564 29672
rect 19604 29632 19605 29672
rect 19563 29623 19605 29632
rect 19947 29672 19989 29681
rect 19947 29632 19948 29672
rect 19988 29632 19989 29672
rect 19947 29623 19989 29632
rect 1152 29504 20452 29528
rect 1152 29464 4928 29504
rect 4968 29464 5010 29504
rect 5050 29464 5092 29504
rect 5132 29464 5174 29504
rect 5214 29464 5256 29504
rect 5296 29464 20048 29504
rect 20088 29464 20130 29504
rect 20170 29464 20212 29504
rect 20252 29464 20294 29504
rect 20334 29464 20376 29504
rect 20416 29464 20452 29504
rect 1152 29440 20452 29464
rect 8427 29336 8469 29345
rect 8427 29296 8428 29336
rect 8468 29296 8469 29336
rect 8427 29287 8469 29296
rect 19947 29336 19989 29345
rect 19947 29296 19948 29336
rect 19988 29296 19989 29336
rect 19947 29287 19989 29296
rect 1507 29168 1565 29169
rect 1507 29128 1516 29168
rect 1556 29128 1565 29168
rect 1507 29127 1565 29128
rect 2755 29168 2813 29169
rect 2755 29128 2764 29168
rect 2804 29128 2813 29168
rect 2755 29127 2813 29128
rect 3811 29168 3869 29169
rect 3811 29128 3820 29168
rect 3860 29128 3869 29168
rect 3811 29127 3869 29128
rect 5059 29168 5117 29169
rect 5059 29128 5068 29168
rect 5108 29128 5117 29168
rect 5059 29127 5117 29128
rect 6979 29168 7037 29169
rect 6979 29128 6988 29168
rect 7028 29128 7037 29168
rect 6979 29127 7037 29128
rect 8227 29168 8285 29169
rect 8227 29128 8236 29168
rect 8276 29128 8285 29168
rect 8227 29127 8285 29128
rect 8707 29168 8765 29169
rect 8707 29128 8716 29168
rect 8756 29128 8765 29168
rect 8707 29127 8765 29128
rect 9955 29168 10013 29169
rect 9955 29128 9964 29168
rect 10004 29128 10013 29168
rect 9955 29127 10013 29128
rect 10339 29168 10397 29169
rect 10339 29128 10348 29168
rect 10388 29128 10397 29168
rect 10339 29127 10397 29128
rect 11587 29168 11645 29169
rect 11587 29128 11596 29168
rect 11636 29128 11645 29168
rect 11587 29127 11645 29128
rect 11971 29168 12029 29169
rect 11971 29128 11980 29168
rect 12020 29128 12029 29168
rect 11971 29127 12029 29128
rect 13219 29168 13277 29169
rect 13219 29128 13228 29168
rect 13268 29128 13277 29168
rect 13219 29127 13277 29128
rect 13603 29168 13661 29169
rect 13603 29128 13612 29168
rect 13652 29128 13661 29168
rect 13603 29127 13661 29128
rect 14851 29168 14909 29169
rect 14851 29128 14860 29168
rect 14900 29128 14909 29168
rect 14851 29127 14909 29128
rect 15235 29168 15293 29169
rect 15235 29128 15244 29168
rect 15284 29128 15293 29168
rect 15235 29127 15293 29128
rect 16483 29168 16541 29169
rect 16483 29128 16492 29168
rect 16532 29128 16541 29168
rect 16483 29127 16541 29128
rect 17059 29168 17117 29169
rect 17059 29128 17068 29168
rect 17108 29128 17117 29168
rect 17059 29127 17117 29128
rect 18307 29168 18365 29169
rect 18307 29128 18316 29168
rect 18356 29128 18365 29168
rect 18307 29127 18365 29128
rect 18499 29168 18557 29169
rect 18499 29128 18508 29168
rect 18548 29128 18557 29168
rect 18499 29127 18557 29128
rect 19747 29168 19805 29169
rect 19747 29128 19756 29168
rect 19796 29128 19805 29168
rect 19747 29127 19805 29128
rect 2955 28916 2997 28925
rect 2955 28876 2956 28916
rect 2996 28876 2997 28916
rect 2955 28867 2997 28876
rect 5259 28916 5301 28925
rect 5259 28876 5260 28916
rect 5300 28876 5301 28916
rect 5259 28867 5301 28876
rect 10155 28916 10197 28925
rect 10155 28876 10156 28916
rect 10196 28876 10197 28916
rect 10155 28867 10197 28876
rect 11787 28916 11829 28925
rect 11787 28876 11788 28916
rect 11828 28876 11829 28916
rect 11787 28867 11829 28876
rect 13419 28916 13461 28925
rect 13419 28876 13420 28916
rect 13460 28876 13461 28916
rect 13419 28867 13461 28876
rect 15051 28916 15093 28925
rect 15051 28876 15052 28916
rect 15092 28876 15093 28916
rect 15051 28867 15093 28876
rect 16683 28916 16725 28925
rect 16683 28876 16684 28916
rect 16724 28876 16725 28916
rect 16683 28867 16725 28876
rect 16875 28916 16917 28925
rect 16875 28876 16876 28916
rect 16916 28876 16917 28916
rect 16875 28867 16917 28876
rect 1152 28748 20352 28772
rect 1152 28708 3688 28748
rect 3728 28708 3770 28748
rect 3810 28708 3852 28748
rect 3892 28708 3934 28748
rect 3974 28708 4016 28748
rect 4056 28708 18808 28748
rect 18848 28708 18890 28748
rect 18930 28708 18972 28748
rect 19012 28708 19054 28748
rect 19094 28708 19136 28748
rect 19176 28708 20352 28748
rect 1152 28684 20352 28708
rect 10635 28412 10677 28421
rect 10635 28372 10636 28412
rect 10676 28372 10677 28412
rect 13899 28412 13941 28421
rect 10635 28363 10677 28372
rect 11739 28370 11781 28379
rect 5163 28342 5205 28351
rect 1891 28328 1949 28329
rect 1891 28288 1900 28328
rect 1940 28288 1949 28328
rect 1891 28287 1949 28288
rect 3139 28328 3197 28329
rect 3139 28288 3148 28328
rect 3188 28288 3197 28328
rect 3139 28287 3197 28288
rect 3627 28328 3669 28337
rect 3627 28288 3628 28328
rect 3668 28288 3669 28328
rect 3627 28279 3669 28288
rect 3723 28328 3765 28337
rect 3723 28288 3724 28328
rect 3764 28288 3765 28328
rect 3723 28279 3765 28288
rect 4107 28328 4149 28337
rect 4107 28288 4108 28328
rect 4148 28288 4149 28328
rect 4107 28279 4149 28288
rect 4203 28328 4245 28337
rect 4203 28288 4204 28328
rect 4244 28288 4245 28328
rect 4203 28279 4245 28288
rect 4675 28328 4733 28329
rect 4675 28288 4684 28328
rect 4724 28288 4733 28328
rect 5163 28302 5164 28342
rect 5204 28302 5205 28342
rect 10155 28347 10197 28356
rect 5163 28293 5205 28302
rect 5923 28328 5981 28329
rect 4675 28287 4733 28288
rect 5923 28288 5932 28328
rect 5972 28288 5981 28328
rect 5923 28287 5981 28288
rect 7171 28328 7229 28329
rect 7171 28288 7180 28328
rect 7220 28288 7229 28328
rect 7171 28287 7229 28288
rect 7747 28328 7805 28329
rect 7747 28288 7756 28328
rect 7796 28288 7805 28328
rect 7747 28287 7805 28288
rect 8995 28328 9053 28329
rect 8995 28288 9004 28328
rect 9044 28288 9053 28328
rect 10155 28307 10156 28347
rect 10196 28307 10197 28347
rect 10155 28298 10197 28307
rect 10251 28328 10293 28337
rect 8995 28287 9053 28288
rect 10251 28288 10252 28328
rect 10292 28288 10293 28328
rect 10251 28279 10293 28288
rect 10731 28328 10773 28337
rect 11739 28330 11740 28370
rect 11780 28330 11781 28370
rect 13899 28372 13900 28412
rect 13940 28372 13941 28412
rect 17059 28412 17117 28413
rect 13899 28363 13941 28372
rect 14907 28370 14949 28379
rect 17059 28372 17068 28412
rect 17108 28372 17117 28412
rect 17059 28371 17117 28372
rect 19459 28412 19517 28413
rect 19459 28372 19468 28412
rect 19508 28372 19517 28412
rect 19459 28371 19517 28372
rect 19843 28412 19901 28413
rect 19843 28372 19852 28412
rect 19892 28372 19901 28412
rect 19843 28371 19901 28372
rect 10731 28288 10732 28328
rect 10772 28288 10773 28328
rect 10731 28279 10773 28288
rect 11203 28328 11261 28329
rect 11203 28288 11212 28328
rect 11252 28288 11261 28328
rect 11739 28321 11781 28330
rect 13323 28328 13365 28337
rect 11203 28287 11261 28288
rect 13323 28288 13324 28328
rect 13364 28288 13365 28328
rect 13323 28279 13365 28288
rect 13419 28328 13461 28337
rect 13419 28288 13420 28328
rect 13460 28288 13461 28328
rect 13419 28279 13461 28288
rect 13803 28328 13845 28337
rect 14907 28330 14908 28370
rect 14948 28330 14949 28370
rect 19131 28337 19173 28346
rect 13803 28288 13804 28328
rect 13844 28288 13845 28328
rect 13803 28279 13845 28288
rect 14371 28328 14429 28329
rect 14371 28288 14380 28328
rect 14420 28288 14429 28328
rect 14907 28321 14949 28330
rect 15235 28328 15293 28329
rect 14371 28287 14429 28288
rect 15235 28288 15244 28328
rect 15284 28288 15293 28328
rect 15235 28287 15293 28288
rect 16483 28328 16541 28329
rect 16483 28288 16492 28328
rect 16532 28288 16541 28328
rect 16483 28287 16541 28288
rect 17547 28328 17589 28337
rect 17547 28288 17548 28328
rect 17588 28288 17589 28328
rect 17547 28279 17589 28288
rect 17643 28328 17685 28337
rect 17643 28288 17644 28328
rect 17684 28288 17685 28328
rect 17643 28279 17685 28288
rect 18027 28328 18069 28337
rect 18027 28288 18028 28328
rect 18068 28288 18069 28328
rect 18027 28279 18069 28288
rect 18123 28328 18165 28337
rect 18123 28288 18124 28328
rect 18164 28288 18165 28328
rect 18123 28279 18165 28288
rect 18595 28328 18653 28329
rect 18595 28288 18604 28328
rect 18644 28288 18653 28328
rect 19131 28297 19132 28337
rect 19172 28297 19173 28337
rect 19131 28288 19173 28297
rect 18595 28287 18653 28288
rect 5355 28244 5397 28253
rect 5355 28204 5356 28244
rect 5396 28204 5397 28244
rect 5355 28195 5397 28204
rect 11883 28244 11925 28253
rect 11883 28204 11884 28244
rect 11924 28204 11925 28244
rect 11883 28195 11925 28204
rect 15051 28244 15093 28253
rect 15051 28204 15052 28244
rect 15092 28204 15093 28244
rect 15051 28195 15093 28204
rect 3339 28160 3381 28169
rect 3339 28120 3340 28160
rect 3380 28120 3381 28160
rect 3339 28111 3381 28120
rect 7371 28160 7413 28169
rect 7371 28120 7372 28160
rect 7412 28120 7413 28160
rect 7371 28111 7413 28120
rect 9195 28160 9237 28169
rect 9195 28120 9196 28160
rect 9236 28120 9237 28160
rect 9195 28111 9237 28120
rect 16683 28160 16725 28169
rect 16683 28120 16684 28160
rect 16724 28120 16725 28160
rect 16683 28111 16725 28120
rect 17259 28160 17301 28169
rect 17259 28120 17260 28160
rect 17300 28120 17301 28160
rect 17259 28111 17301 28120
rect 19275 28160 19317 28169
rect 19275 28120 19276 28160
rect 19316 28120 19317 28160
rect 19275 28111 19317 28120
rect 19659 28160 19701 28169
rect 19659 28120 19660 28160
rect 19700 28120 19701 28160
rect 19659 28111 19701 28120
rect 20043 28160 20085 28169
rect 20043 28120 20044 28160
rect 20084 28120 20085 28160
rect 20043 28111 20085 28120
rect 1152 27992 20452 28016
rect 1152 27952 4928 27992
rect 4968 27952 5010 27992
rect 5050 27952 5092 27992
rect 5132 27952 5174 27992
rect 5214 27952 5256 27992
rect 5296 27952 20048 27992
rect 20088 27952 20130 27992
rect 20170 27952 20212 27992
rect 20252 27952 20294 27992
rect 20334 27952 20376 27992
rect 20416 27952 20452 27992
rect 1152 27928 20452 27952
rect 19755 27824 19797 27833
rect 19755 27784 19756 27824
rect 19796 27784 19797 27824
rect 19755 27775 19797 27784
rect 4203 27740 4245 27749
rect 4203 27700 4204 27740
rect 4244 27700 4245 27740
rect 4203 27691 4245 27700
rect 7275 27740 7317 27749
rect 7275 27700 7276 27740
rect 7316 27700 7317 27740
rect 7275 27691 7317 27700
rect 9291 27740 9333 27749
rect 9291 27700 9292 27740
rect 9332 27700 9333 27740
rect 9291 27691 9333 27700
rect 12171 27740 12213 27749
rect 12171 27700 12172 27740
rect 12212 27700 12213 27740
rect 12171 27691 12213 27700
rect 16491 27740 16533 27749
rect 16491 27700 16492 27740
rect 16532 27700 16533 27740
rect 16491 27691 16533 27700
rect 2475 27656 2517 27665
rect 2475 27616 2476 27656
rect 2516 27616 2517 27656
rect 2475 27607 2517 27616
rect 2571 27656 2613 27665
rect 2571 27616 2572 27656
rect 2612 27616 2613 27656
rect 2571 27607 2613 27616
rect 2955 27656 2997 27665
rect 2955 27616 2956 27656
rect 2996 27616 2997 27656
rect 2955 27607 2997 27616
rect 3523 27656 3581 27657
rect 3523 27616 3532 27656
rect 3572 27616 3581 27656
rect 3523 27615 3581 27616
rect 4011 27651 4053 27660
rect 4011 27611 4012 27651
rect 4052 27611 4053 27651
rect 4011 27602 4053 27611
rect 5547 27656 5589 27665
rect 5547 27616 5548 27656
rect 5588 27616 5589 27656
rect 5547 27607 5589 27616
rect 5643 27656 5685 27665
rect 5643 27616 5644 27656
rect 5684 27616 5685 27656
rect 5643 27607 5685 27616
rect 6595 27656 6653 27657
rect 6595 27616 6604 27656
rect 6644 27616 6653 27656
rect 7563 27656 7605 27665
rect 6595 27615 6653 27616
rect 7083 27642 7125 27651
rect 7083 27602 7084 27642
rect 7124 27602 7125 27642
rect 7563 27616 7564 27656
rect 7604 27616 7605 27656
rect 7563 27607 7605 27616
rect 7659 27656 7701 27665
rect 7659 27616 7660 27656
rect 7700 27616 7701 27656
rect 7659 27607 7701 27616
rect 8043 27656 8085 27665
rect 8043 27616 8044 27656
rect 8084 27616 8085 27656
rect 8043 27607 8085 27616
rect 8139 27656 8181 27665
rect 8139 27616 8140 27656
rect 8180 27616 8181 27656
rect 8139 27607 8181 27616
rect 8611 27656 8669 27657
rect 8611 27616 8620 27656
rect 8660 27616 8669 27656
rect 10443 27656 10485 27665
rect 8611 27615 8669 27616
rect 9147 27646 9189 27655
rect 7083 27593 7125 27602
rect 9147 27606 9148 27646
rect 9188 27606 9189 27646
rect 10443 27616 10444 27656
rect 10484 27616 10485 27656
rect 10443 27607 10485 27616
rect 10539 27656 10581 27665
rect 10539 27616 10540 27656
rect 10580 27616 10581 27656
rect 10539 27607 10581 27616
rect 11019 27656 11061 27665
rect 11019 27616 11020 27656
rect 11060 27616 11061 27656
rect 11019 27607 11061 27616
rect 11491 27656 11549 27657
rect 11491 27616 11500 27656
rect 11540 27616 11549 27656
rect 13027 27656 13085 27657
rect 11491 27615 11549 27616
rect 11979 27642 12021 27651
rect 9147 27597 9189 27606
rect 11979 27602 11980 27642
rect 12020 27602 12021 27642
rect 13027 27616 13036 27656
rect 13076 27616 13085 27656
rect 13027 27615 13085 27616
rect 14275 27656 14333 27657
rect 14275 27616 14284 27656
rect 14324 27616 14333 27656
rect 14275 27615 14333 27616
rect 14763 27656 14805 27665
rect 14763 27616 14764 27656
rect 14804 27616 14805 27656
rect 14763 27607 14805 27616
rect 14859 27656 14901 27665
rect 14859 27616 14860 27656
rect 14900 27616 14901 27656
rect 14859 27607 14901 27616
rect 15339 27656 15381 27665
rect 15339 27616 15340 27656
rect 15380 27616 15381 27656
rect 15339 27607 15381 27616
rect 15811 27656 15869 27657
rect 15811 27616 15820 27656
rect 15860 27616 15869 27656
rect 15811 27615 15869 27616
rect 16299 27651 16341 27660
rect 16299 27611 16300 27651
rect 16340 27611 16341 27651
rect 16675 27656 16733 27657
rect 16675 27616 16684 27656
rect 16724 27616 16733 27656
rect 16675 27615 16733 27616
rect 17923 27656 17981 27657
rect 17923 27616 17932 27656
rect 17972 27616 17981 27656
rect 17923 27615 17981 27616
rect 18307 27656 18365 27657
rect 18307 27616 18316 27656
rect 18356 27616 18365 27656
rect 18307 27615 18365 27616
rect 19555 27656 19613 27657
rect 19555 27616 19564 27656
rect 19604 27616 19613 27656
rect 19555 27615 19613 27616
rect 16299 27602 16341 27611
rect 11979 27593 12021 27602
rect 3051 27572 3093 27581
rect 3051 27532 3052 27572
rect 3092 27532 3093 27572
rect 3051 27523 3093 27532
rect 6027 27572 6069 27581
rect 6027 27532 6028 27572
rect 6068 27532 6069 27572
rect 6027 27523 6069 27532
rect 6123 27572 6165 27581
rect 6123 27532 6124 27572
rect 6164 27532 6165 27572
rect 6123 27523 6165 27532
rect 10923 27572 10965 27581
rect 10923 27532 10924 27572
rect 10964 27532 10965 27572
rect 10923 27523 10965 27532
rect 15243 27572 15285 27581
rect 15243 27532 15244 27572
rect 15284 27532 15285 27572
rect 15243 27523 15285 27532
rect 19939 27572 19997 27573
rect 19939 27532 19948 27572
rect 19988 27532 19997 27572
rect 19939 27531 19997 27532
rect 14475 27404 14517 27413
rect 14475 27364 14476 27404
rect 14516 27364 14517 27404
rect 14475 27355 14517 27364
rect 18123 27404 18165 27413
rect 18123 27364 18124 27404
rect 18164 27364 18165 27404
rect 18123 27355 18165 27364
rect 20139 27404 20181 27413
rect 20139 27364 20140 27404
rect 20180 27364 20181 27404
rect 20139 27355 20181 27364
rect 1152 27236 20352 27260
rect 1152 27196 3688 27236
rect 3728 27196 3770 27236
rect 3810 27196 3852 27236
rect 3892 27196 3934 27236
rect 3974 27196 4016 27236
rect 4056 27196 18808 27236
rect 18848 27196 18890 27236
rect 18930 27196 18972 27236
rect 19012 27196 19054 27236
rect 19094 27196 19136 27236
rect 19176 27196 20352 27236
rect 1152 27172 20352 27196
rect 2667 27068 2709 27077
rect 2667 27028 2668 27068
rect 2708 27028 2709 27068
rect 2667 27019 2709 27028
rect 5931 27068 5973 27077
rect 5931 27028 5932 27068
rect 5972 27028 5973 27068
rect 5931 27019 5973 27028
rect 7563 27068 7605 27077
rect 7563 27028 7564 27068
rect 7604 27028 7605 27068
rect 7563 27019 7605 27028
rect 10347 27068 10389 27077
rect 10347 27028 10348 27068
rect 10388 27028 10389 27068
rect 10347 27019 10389 27028
rect 18507 26984 18549 26993
rect 18507 26944 18508 26984
rect 18548 26944 18549 26984
rect 18507 26935 18549 26944
rect 17163 26900 17205 26909
rect 17163 26860 17164 26900
rect 17204 26860 17205 26900
rect 17163 26851 17205 26860
rect 18171 26825 18213 26834
rect 1219 26816 1277 26817
rect 1219 26776 1228 26816
rect 1268 26776 1277 26816
rect 1219 26775 1277 26776
rect 2467 26816 2525 26817
rect 2467 26776 2476 26816
rect 2516 26776 2525 26816
rect 2467 26775 2525 26776
rect 2851 26816 2909 26817
rect 2851 26776 2860 26816
rect 2900 26776 2909 26816
rect 2851 26775 2909 26776
rect 4099 26816 4157 26817
rect 4099 26776 4108 26816
rect 4148 26776 4157 26816
rect 4099 26775 4157 26776
rect 4483 26816 4541 26817
rect 4483 26776 4492 26816
rect 4532 26776 4541 26816
rect 4483 26775 4541 26776
rect 5731 26816 5789 26817
rect 5731 26776 5740 26816
rect 5780 26776 5789 26816
rect 5731 26775 5789 26776
rect 6115 26816 6173 26817
rect 6115 26776 6124 26816
rect 6164 26776 6173 26816
rect 6115 26775 6173 26776
rect 7363 26816 7421 26817
rect 7363 26776 7372 26816
rect 7412 26776 7421 26816
rect 7363 26775 7421 26776
rect 8899 26816 8957 26817
rect 8899 26776 8908 26816
rect 8948 26776 8957 26816
rect 8899 26775 8957 26776
rect 10147 26816 10205 26817
rect 10147 26776 10156 26816
rect 10196 26776 10205 26816
rect 10147 26775 10205 26776
rect 10819 26816 10877 26817
rect 10819 26776 10828 26816
rect 10868 26776 10877 26816
rect 10819 26775 10877 26776
rect 12067 26816 12125 26817
rect 12067 26776 12076 26816
rect 12116 26776 12125 26816
rect 12067 26775 12125 26776
rect 13603 26816 13661 26817
rect 13603 26776 13612 26816
rect 13652 26776 13661 26816
rect 13603 26775 13661 26776
rect 14851 26816 14909 26817
rect 14851 26776 14860 26816
rect 14900 26776 14909 26816
rect 14851 26775 14909 26776
rect 16587 26816 16629 26825
rect 16587 26776 16588 26816
rect 16628 26776 16629 26816
rect 16587 26767 16629 26776
rect 16683 26816 16725 26825
rect 16683 26776 16684 26816
rect 16724 26776 16725 26816
rect 16683 26767 16725 26776
rect 17067 26816 17109 26825
rect 17067 26776 17068 26816
rect 17108 26776 17109 26816
rect 17067 26767 17109 26776
rect 17635 26816 17693 26817
rect 17635 26776 17644 26816
rect 17684 26776 17693 26816
rect 18171 26785 18172 26825
rect 18212 26785 18213 26825
rect 18171 26776 18213 26785
rect 18691 26816 18749 26817
rect 18691 26776 18700 26816
rect 18740 26776 18749 26816
rect 17635 26775 17693 26776
rect 18691 26775 18749 26776
rect 19939 26816 19997 26817
rect 19939 26776 19948 26816
rect 19988 26776 19997 26816
rect 19939 26775 19997 26776
rect 4299 26648 4341 26657
rect 4299 26608 4300 26648
rect 4340 26608 4341 26648
rect 4299 26599 4341 26608
rect 12267 26648 12309 26657
rect 12267 26608 12268 26648
rect 12308 26608 12309 26648
rect 12267 26599 12309 26608
rect 15051 26648 15093 26657
rect 15051 26608 15052 26648
rect 15092 26608 15093 26648
rect 15051 26599 15093 26608
rect 18315 26648 18357 26657
rect 18315 26608 18316 26648
rect 18356 26608 18357 26648
rect 18315 26599 18357 26608
rect 1152 26480 20452 26504
rect 1152 26440 4928 26480
rect 4968 26440 5010 26480
rect 5050 26440 5092 26480
rect 5132 26440 5174 26480
rect 5214 26440 5256 26480
rect 5296 26440 20048 26480
rect 20088 26440 20130 26480
rect 20170 26440 20212 26480
rect 20252 26440 20294 26480
rect 20334 26440 20376 26480
rect 20416 26440 20452 26480
rect 1152 26416 20452 26440
rect 5067 26228 5109 26237
rect 5067 26188 5068 26228
rect 5108 26188 5109 26228
rect 5067 26179 5109 26188
rect 19179 26228 19221 26237
rect 19179 26188 19180 26228
rect 19220 26188 19221 26228
rect 19179 26179 19221 26188
rect 1603 26144 1661 26145
rect 1603 26104 1612 26144
rect 1652 26104 1661 26144
rect 1603 26103 1661 26104
rect 2851 26144 2909 26145
rect 2851 26104 2860 26144
rect 2900 26104 2909 26144
rect 3435 26144 3477 26153
rect 2851 26103 2909 26104
rect 3339 26125 3381 26134
rect 3339 26085 3340 26125
rect 3380 26085 3381 26125
rect 3435 26104 3436 26144
rect 3476 26104 3477 26144
rect 3435 26095 3477 26104
rect 4387 26144 4445 26145
rect 4387 26104 4396 26144
rect 4436 26104 4445 26144
rect 4387 26103 4445 26104
rect 4875 26139 4917 26148
rect 4875 26099 4876 26139
rect 4916 26099 4917 26139
rect 5443 26144 5501 26145
rect 5443 26104 5452 26144
rect 5492 26104 5501 26144
rect 5443 26103 5501 26104
rect 6691 26144 6749 26145
rect 6691 26104 6700 26144
rect 6740 26104 6749 26144
rect 6691 26103 6749 26104
rect 7075 26144 7133 26145
rect 7075 26104 7084 26144
rect 7124 26104 7133 26144
rect 7075 26103 7133 26104
rect 8323 26144 8381 26145
rect 8323 26104 8332 26144
rect 8372 26104 8381 26144
rect 8323 26103 8381 26104
rect 9187 26144 9245 26145
rect 9187 26104 9196 26144
rect 9236 26104 9245 26144
rect 9187 26103 9245 26104
rect 10435 26144 10493 26145
rect 10435 26104 10444 26144
rect 10484 26104 10493 26144
rect 10435 26103 10493 26104
rect 10819 26144 10877 26145
rect 10819 26104 10828 26144
rect 10868 26104 10877 26144
rect 10819 26103 10877 26104
rect 12067 26144 12125 26145
rect 12067 26104 12076 26144
rect 12116 26104 12125 26144
rect 12067 26103 12125 26104
rect 12451 26144 12509 26145
rect 12451 26104 12460 26144
rect 12500 26104 12509 26144
rect 12451 26103 12509 26104
rect 13699 26144 13757 26145
rect 13699 26104 13708 26144
rect 13748 26104 13757 26144
rect 13699 26103 13757 26104
rect 14851 26144 14909 26145
rect 14851 26104 14860 26144
rect 14900 26104 14909 26144
rect 14851 26103 14909 26104
rect 16099 26144 16157 26145
rect 16099 26104 16108 26144
rect 16148 26104 16157 26144
rect 16099 26103 16157 26104
rect 17451 26144 17493 26153
rect 17451 26104 17452 26144
rect 17492 26104 17493 26144
rect 4875 26090 4917 26099
rect 17451 26095 17493 26104
rect 17547 26144 17589 26153
rect 17547 26104 17548 26144
rect 17588 26104 17589 26144
rect 17547 26095 17589 26104
rect 18499 26144 18557 26145
rect 18499 26104 18508 26144
rect 18548 26104 18557 26144
rect 18499 26103 18557 26104
rect 19035 26102 19077 26111
rect 3339 26076 3381 26085
rect 3819 26060 3861 26069
rect 3819 26020 3820 26060
rect 3860 26020 3861 26060
rect 3819 26011 3861 26020
rect 3915 26060 3957 26069
rect 3915 26020 3916 26060
rect 3956 26020 3957 26060
rect 3915 26011 3957 26020
rect 17931 26060 17973 26069
rect 17931 26020 17932 26060
rect 17972 26020 17973 26060
rect 17931 26011 17973 26020
rect 18027 26060 18069 26069
rect 18027 26020 18028 26060
rect 18068 26020 18069 26060
rect 19035 26062 19036 26102
rect 19076 26062 19077 26102
rect 19035 26053 19077 26062
rect 19363 26060 19421 26061
rect 18027 26011 18069 26020
rect 19363 26020 19372 26060
rect 19412 26020 19421 26060
rect 19363 26019 19421 26020
rect 19747 26060 19805 26061
rect 19747 26020 19756 26060
rect 19796 26020 19805 26060
rect 19747 26019 19805 26020
rect 3051 25892 3093 25901
rect 3051 25852 3052 25892
rect 3092 25852 3093 25892
rect 3051 25843 3093 25852
rect 6891 25892 6933 25901
rect 6891 25852 6892 25892
rect 6932 25852 6933 25892
rect 6891 25843 6933 25852
rect 8523 25892 8565 25901
rect 8523 25852 8524 25892
rect 8564 25852 8565 25892
rect 8523 25843 8565 25852
rect 10635 25892 10677 25901
rect 10635 25852 10636 25892
rect 10676 25852 10677 25892
rect 10635 25843 10677 25852
rect 12267 25892 12309 25901
rect 12267 25852 12268 25892
rect 12308 25852 12309 25892
rect 12267 25843 12309 25852
rect 13899 25892 13941 25901
rect 13899 25852 13900 25892
rect 13940 25852 13941 25892
rect 13899 25843 13941 25852
rect 16299 25892 16341 25901
rect 16299 25852 16300 25892
rect 16340 25852 16341 25892
rect 16299 25843 16341 25852
rect 19563 25892 19605 25901
rect 19563 25852 19564 25892
rect 19604 25852 19605 25892
rect 19563 25843 19605 25852
rect 19947 25892 19989 25901
rect 19947 25852 19948 25892
rect 19988 25852 19989 25892
rect 19947 25843 19989 25852
rect 1152 25724 20352 25748
rect 1152 25684 3688 25724
rect 3728 25684 3770 25724
rect 3810 25684 3852 25724
rect 3892 25684 3934 25724
rect 3974 25684 4016 25724
rect 4056 25684 18808 25724
rect 18848 25684 18890 25724
rect 18930 25684 18972 25724
rect 19012 25684 19054 25724
rect 19094 25684 19136 25724
rect 19176 25684 20352 25724
rect 1152 25660 20352 25684
rect 3147 25556 3189 25565
rect 3147 25516 3148 25556
rect 3188 25516 3189 25556
rect 3147 25507 3189 25516
rect 19467 25556 19509 25565
rect 19467 25516 19468 25556
rect 19508 25516 19509 25556
rect 19467 25507 19509 25516
rect 19851 25472 19893 25481
rect 19851 25432 19852 25472
rect 19892 25432 19893 25472
rect 19851 25423 19893 25432
rect 4203 25388 4245 25397
rect 4203 25348 4204 25388
rect 4244 25348 4245 25388
rect 4203 25339 4245 25348
rect 4299 25388 4341 25397
rect 4299 25348 4300 25388
rect 4340 25348 4341 25388
rect 4299 25339 4341 25348
rect 11403 25388 11445 25397
rect 11403 25348 11404 25388
rect 11444 25348 11445 25388
rect 11403 25339 11445 25348
rect 19651 25388 19709 25389
rect 19651 25348 19660 25388
rect 19700 25348 19709 25388
rect 19651 25347 19709 25348
rect 20035 25388 20093 25389
rect 20035 25348 20044 25388
rect 20084 25348 20093 25388
rect 20035 25347 20093 25348
rect 5307 25313 5349 25322
rect 8619 25318 8661 25327
rect 1699 25304 1757 25305
rect 1699 25264 1708 25304
rect 1748 25264 1757 25304
rect 1699 25263 1757 25264
rect 2947 25304 3005 25305
rect 2947 25264 2956 25304
rect 2996 25264 3005 25304
rect 2947 25263 3005 25264
rect 3723 25304 3765 25313
rect 3723 25264 3724 25304
rect 3764 25264 3765 25304
rect 3723 25255 3765 25264
rect 3819 25304 3861 25313
rect 3819 25264 3820 25304
rect 3860 25264 3861 25304
rect 3819 25255 3861 25264
rect 4771 25304 4829 25305
rect 4771 25264 4780 25304
rect 4820 25264 4829 25304
rect 5307 25273 5308 25313
rect 5348 25273 5349 25313
rect 5307 25264 5349 25273
rect 7083 25303 7125 25312
rect 4771 25263 4829 25264
rect 7083 25263 7084 25303
rect 7124 25263 7125 25303
rect 7083 25254 7125 25263
rect 7179 25304 7221 25313
rect 7179 25264 7180 25304
rect 7220 25264 7221 25304
rect 7179 25255 7221 25264
rect 7563 25304 7605 25313
rect 7563 25264 7564 25304
rect 7604 25264 7605 25304
rect 7563 25255 7605 25264
rect 7659 25304 7701 25313
rect 7659 25264 7660 25304
rect 7700 25264 7701 25304
rect 7659 25255 7701 25264
rect 8131 25304 8189 25305
rect 8131 25264 8140 25304
rect 8180 25264 8189 25304
rect 8619 25278 8620 25318
rect 8660 25278 8661 25318
rect 12363 25318 12405 25327
rect 8619 25269 8661 25278
rect 9091 25304 9149 25305
rect 8131 25263 8189 25264
rect 9091 25264 9100 25304
rect 9140 25264 9149 25304
rect 9091 25263 9149 25264
rect 10339 25304 10397 25305
rect 10339 25264 10348 25304
rect 10388 25264 10397 25304
rect 10339 25263 10397 25264
rect 10827 25304 10869 25313
rect 10827 25264 10828 25304
rect 10868 25264 10869 25304
rect 10827 25255 10869 25264
rect 10923 25304 10965 25313
rect 10923 25264 10924 25304
rect 10964 25264 10965 25304
rect 10923 25255 10965 25264
rect 11307 25304 11349 25313
rect 11307 25264 11308 25304
rect 11348 25264 11349 25304
rect 11307 25255 11349 25264
rect 11875 25304 11933 25305
rect 11875 25264 11884 25304
rect 11924 25264 11933 25304
rect 12363 25278 12364 25318
rect 12404 25278 12405 25318
rect 15243 25318 15285 25327
rect 12363 25269 12405 25278
rect 13707 25304 13749 25313
rect 11875 25263 11933 25264
rect 13707 25264 13708 25304
rect 13748 25264 13749 25304
rect 13707 25255 13749 25264
rect 13803 25304 13845 25313
rect 13803 25264 13804 25304
rect 13844 25264 13845 25304
rect 13803 25255 13845 25264
rect 14187 25304 14229 25313
rect 14187 25264 14188 25304
rect 14228 25264 14229 25304
rect 14187 25255 14229 25264
rect 14283 25304 14325 25313
rect 14283 25264 14284 25304
rect 14324 25264 14325 25304
rect 14283 25255 14325 25264
rect 14755 25304 14813 25305
rect 14755 25264 14764 25304
rect 14804 25264 14813 25304
rect 15243 25278 15244 25318
rect 15284 25278 15285 25318
rect 15243 25269 15285 25278
rect 16387 25304 16445 25305
rect 14755 25263 14813 25264
rect 16387 25264 16396 25304
rect 16436 25264 16445 25304
rect 16387 25263 16445 25264
rect 17635 25304 17693 25305
rect 17635 25264 17644 25304
rect 17684 25264 17693 25304
rect 17635 25263 17693 25264
rect 18019 25304 18077 25305
rect 18019 25264 18028 25304
rect 18068 25264 18077 25304
rect 18019 25263 18077 25264
rect 19267 25304 19325 25305
rect 19267 25264 19276 25304
rect 19316 25264 19325 25304
rect 19267 25263 19325 25264
rect 5451 25220 5493 25229
rect 5451 25180 5452 25220
rect 5492 25180 5493 25220
rect 5451 25171 5493 25180
rect 8811 25220 8853 25229
rect 8811 25180 8812 25220
rect 8852 25180 8853 25220
rect 8811 25171 8853 25180
rect 10539 25220 10581 25229
rect 10539 25180 10540 25220
rect 10580 25180 10581 25220
rect 10539 25171 10581 25180
rect 12555 25136 12597 25145
rect 12555 25096 12556 25136
rect 12596 25096 12597 25136
rect 12555 25087 12597 25096
rect 15435 25136 15477 25145
rect 15435 25096 15436 25136
rect 15476 25096 15477 25136
rect 15435 25087 15477 25096
rect 17835 25136 17877 25145
rect 17835 25096 17836 25136
rect 17876 25096 17877 25136
rect 17835 25087 17877 25096
rect 20235 25136 20277 25145
rect 20235 25096 20236 25136
rect 20276 25096 20277 25136
rect 20235 25087 20277 25096
rect 1152 24968 20452 24992
rect 1152 24928 4928 24968
rect 4968 24928 5010 24968
rect 5050 24928 5092 24968
rect 5132 24928 5174 24968
rect 5214 24928 5256 24968
rect 5296 24928 20048 24968
rect 20088 24928 20130 24968
rect 20170 24928 20212 24968
rect 20252 24928 20294 24968
rect 20334 24928 20376 24968
rect 20416 24928 20452 24968
rect 1152 24904 20452 24928
rect 3139 24800 3197 24801
rect 3139 24760 3148 24800
rect 3188 24760 3197 24800
rect 3139 24759 3197 24760
rect 5067 24800 5109 24809
rect 5067 24760 5068 24800
rect 5108 24760 5109 24800
rect 5067 24751 5109 24760
rect 11691 24800 11733 24809
rect 11691 24760 11692 24800
rect 11732 24760 11733 24800
rect 11691 24751 11733 24760
rect 18795 24800 18837 24809
rect 18795 24760 18796 24800
rect 18836 24760 18837 24800
rect 18795 24751 18837 24760
rect 6699 24716 6741 24725
rect 6699 24676 6700 24716
rect 6740 24676 6741 24716
rect 6699 24667 6741 24676
rect 9675 24716 9717 24725
rect 9675 24676 9676 24716
rect 9716 24676 9717 24716
rect 9675 24667 9717 24676
rect 18219 24716 18261 24725
rect 18219 24676 18220 24716
rect 18260 24676 18261 24716
rect 18219 24667 18261 24676
rect 1219 24632 1277 24633
rect 1219 24592 1228 24632
rect 1268 24592 1277 24632
rect 1219 24591 1277 24592
rect 2467 24632 2525 24633
rect 2467 24592 2476 24632
rect 2516 24592 2525 24632
rect 2467 24591 2525 24592
rect 2859 24632 2901 24641
rect 2859 24592 2860 24632
rect 2900 24592 2901 24632
rect 2859 24583 2901 24592
rect 2955 24632 2997 24641
rect 2955 24592 2956 24632
rect 2996 24592 2997 24632
rect 2955 24583 2997 24592
rect 3619 24632 3677 24633
rect 3619 24592 3628 24632
rect 3668 24592 3677 24632
rect 3619 24591 3677 24592
rect 4867 24632 4925 24633
rect 4867 24592 4876 24632
rect 4916 24592 4925 24632
rect 4867 24591 4925 24592
rect 5251 24632 5309 24633
rect 5251 24592 5260 24632
rect 5300 24592 5309 24632
rect 5251 24591 5309 24592
rect 6499 24632 6557 24633
rect 6499 24592 6508 24632
rect 6548 24592 6557 24632
rect 6499 24591 6557 24592
rect 7171 24632 7229 24633
rect 7171 24592 7180 24632
rect 7220 24592 7229 24632
rect 7171 24591 7229 24592
rect 7467 24632 7509 24641
rect 7467 24592 7468 24632
rect 7508 24592 7509 24632
rect 7467 24583 7509 24592
rect 7563 24632 7605 24641
rect 7563 24592 7564 24632
rect 7604 24592 7605 24632
rect 7563 24583 7605 24592
rect 8227 24632 8285 24633
rect 8227 24592 8236 24632
rect 8276 24592 8285 24632
rect 8227 24591 8285 24592
rect 9475 24632 9533 24633
rect 9475 24592 9484 24632
rect 9524 24592 9533 24632
rect 9475 24591 9533 24592
rect 9963 24632 10005 24641
rect 9963 24592 9964 24632
rect 10004 24592 10005 24632
rect 9963 24583 10005 24592
rect 10059 24632 10101 24641
rect 10059 24592 10060 24632
rect 10100 24592 10101 24632
rect 10059 24583 10101 24592
rect 11011 24632 11069 24633
rect 11011 24592 11020 24632
rect 11060 24592 11069 24632
rect 11011 24591 11069 24592
rect 11499 24627 11541 24636
rect 11499 24587 11500 24627
rect 11540 24587 11541 24627
rect 13891 24632 13949 24633
rect 13891 24592 13900 24632
rect 13940 24592 13949 24632
rect 13891 24591 13949 24592
rect 15139 24632 15197 24633
rect 15139 24592 15148 24632
rect 15188 24592 15197 24632
rect 15139 24591 15197 24592
rect 16491 24632 16533 24641
rect 16491 24592 16492 24632
rect 16532 24592 16533 24632
rect 11499 24578 11541 24587
rect 16491 24583 16533 24592
rect 16587 24632 16629 24641
rect 16587 24592 16588 24632
rect 16628 24592 16629 24632
rect 16587 24583 16629 24592
rect 17539 24632 17597 24633
rect 17539 24592 17548 24632
rect 17588 24592 17597 24632
rect 17539 24591 17597 24592
rect 18027 24627 18069 24636
rect 18027 24587 18028 24627
rect 18068 24587 18069 24627
rect 18027 24578 18069 24587
rect 10443 24548 10485 24557
rect 10443 24508 10444 24548
rect 10484 24508 10485 24548
rect 10443 24499 10485 24508
rect 10539 24548 10581 24557
rect 10539 24508 10540 24548
rect 10580 24508 10581 24548
rect 10539 24499 10581 24508
rect 16971 24548 17013 24557
rect 16971 24508 16972 24548
rect 17012 24508 17013 24548
rect 16971 24499 17013 24508
rect 17067 24548 17109 24557
rect 17067 24508 17068 24548
rect 17108 24508 17109 24548
rect 17067 24499 17109 24508
rect 18595 24548 18653 24549
rect 18595 24508 18604 24548
rect 18644 24508 18653 24548
rect 18595 24507 18653 24508
rect 18979 24548 19037 24549
rect 18979 24508 18988 24548
rect 19028 24508 19037 24548
rect 18979 24507 19037 24508
rect 19363 24548 19421 24549
rect 19363 24508 19372 24548
rect 19412 24508 19421 24548
rect 19363 24507 19421 24508
rect 19747 24545 19805 24546
rect 19747 24505 19756 24545
rect 19796 24505 19805 24545
rect 19747 24504 19805 24505
rect 2667 24380 2709 24389
rect 2667 24340 2668 24380
rect 2708 24340 2709 24380
rect 2667 24331 2709 24340
rect 7843 24380 7901 24381
rect 7843 24340 7852 24380
rect 7892 24340 7901 24380
rect 7843 24339 7901 24340
rect 15339 24380 15381 24389
rect 15339 24340 15340 24380
rect 15380 24340 15381 24380
rect 15339 24331 15381 24340
rect 19179 24380 19221 24389
rect 19179 24340 19180 24380
rect 19220 24340 19221 24380
rect 19179 24331 19221 24340
rect 19563 24380 19605 24389
rect 19563 24340 19564 24380
rect 19604 24340 19605 24380
rect 19563 24331 19605 24340
rect 19947 24380 19989 24389
rect 19947 24340 19948 24380
rect 19988 24340 19989 24380
rect 19947 24331 19989 24340
rect 1152 24212 20352 24236
rect 1152 24172 3688 24212
rect 3728 24172 3770 24212
rect 3810 24172 3852 24212
rect 3892 24172 3934 24212
rect 3974 24172 4016 24212
rect 4056 24172 18808 24212
rect 18848 24172 18890 24212
rect 18930 24172 18972 24212
rect 19012 24172 19054 24212
rect 19094 24172 19136 24212
rect 19176 24172 20352 24212
rect 1152 24148 20352 24172
rect 2667 24044 2709 24053
rect 2667 24004 2668 24044
rect 2708 24004 2709 24044
rect 2667 23995 2709 24004
rect 15915 23960 15957 23969
rect 15915 23920 15916 23960
rect 15956 23920 15957 23960
rect 15915 23911 15957 23920
rect 4003 23876 4061 23877
rect 3339 23837 3381 23846
rect 1219 23792 1277 23793
rect 1219 23752 1228 23792
rect 1268 23752 1277 23792
rect 1219 23751 1277 23752
rect 2467 23792 2525 23793
rect 2467 23752 2476 23792
rect 2516 23752 2525 23792
rect 2955 23792 2997 23801
rect 2467 23751 2525 23752
rect 2859 23771 2901 23780
rect 2859 23731 2860 23771
rect 2900 23731 2901 23771
rect 2955 23752 2956 23792
rect 2996 23752 2997 23792
rect 2955 23743 2997 23752
rect 3051 23792 3093 23801
rect 3051 23752 3052 23792
rect 3092 23752 3093 23792
rect 3339 23797 3340 23837
rect 3380 23797 3381 23837
rect 4003 23836 4012 23876
rect 4052 23836 4061 23876
rect 4003 23835 4061 23836
rect 11307 23876 11349 23885
rect 11307 23836 11308 23876
rect 11348 23836 11349 23876
rect 3339 23788 3381 23797
rect 3427 23834 3485 23835
rect 3427 23794 3436 23834
rect 3476 23794 3485 23834
rect 11307 23827 11349 23836
rect 14379 23876 14421 23885
rect 14379 23836 14380 23876
rect 14420 23836 14421 23876
rect 14379 23827 14421 23836
rect 15715 23876 15773 23877
rect 15715 23836 15724 23876
rect 15764 23836 15773 23876
rect 15715 23835 15773 23836
rect 18411 23876 18453 23885
rect 18411 23836 18412 23876
rect 18452 23836 18453 23876
rect 18411 23827 18453 23836
rect 15339 23806 15381 23815
rect 3427 23793 3485 23794
rect 3531 23792 3573 23801
rect 3051 23743 3093 23752
rect 3531 23752 3532 23792
rect 3572 23752 3573 23792
rect 3531 23743 3573 23752
rect 4491 23792 4533 23801
rect 4491 23752 4492 23792
rect 4532 23752 4533 23792
rect 4491 23743 4533 23752
rect 4587 23792 4629 23801
rect 4587 23752 4588 23792
rect 4628 23752 4629 23792
rect 4587 23743 4629 23752
rect 4683 23792 4725 23801
rect 4683 23752 4684 23792
rect 4724 23752 4725 23792
rect 4683 23743 4725 23752
rect 5059 23792 5117 23793
rect 5059 23752 5068 23792
rect 5108 23752 5117 23792
rect 5059 23751 5117 23752
rect 5163 23792 5205 23801
rect 5163 23752 5164 23792
rect 5204 23752 5205 23792
rect 5163 23743 5205 23752
rect 5355 23792 5397 23801
rect 5355 23752 5356 23792
rect 5396 23752 5397 23792
rect 5355 23743 5397 23752
rect 5635 23792 5693 23793
rect 5635 23752 5644 23792
rect 5684 23752 5693 23792
rect 5635 23751 5693 23752
rect 6883 23792 6941 23793
rect 6883 23752 6892 23792
rect 6932 23752 6941 23792
rect 6883 23751 6941 23752
rect 7267 23792 7325 23793
rect 7267 23752 7276 23792
rect 7316 23752 7325 23792
rect 7267 23751 7325 23752
rect 8515 23792 8573 23793
rect 8515 23752 8524 23792
rect 8564 23752 8573 23792
rect 8515 23751 8573 23752
rect 8995 23792 9053 23793
rect 8995 23752 9004 23792
rect 9044 23752 9053 23792
rect 8995 23751 9053 23752
rect 10243 23792 10301 23793
rect 10243 23752 10252 23792
rect 10292 23752 10301 23792
rect 10243 23751 10301 23752
rect 10731 23791 10773 23800
rect 10731 23751 10732 23791
rect 10772 23751 10773 23791
rect 10731 23742 10773 23751
rect 10827 23792 10869 23801
rect 10827 23752 10828 23792
rect 10868 23752 10869 23792
rect 10827 23743 10869 23752
rect 11211 23792 11253 23801
rect 12267 23797 12309 23806
rect 11211 23752 11212 23792
rect 11252 23752 11253 23792
rect 11211 23743 11253 23752
rect 11779 23792 11837 23793
rect 11779 23752 11788 23792
rect 11828 23752 11837 23792
rect 11779 23751 11837 23752
rect 12267 23757 12268 23797
rect 12308 23757 12309 23797
rect 12267 23748 12309 23757
rect 13803 23792 13845 23801
rect 13803 23752 13804 23792
rect 13844 23752 13845 23792
rect 13803 23743 13845 23752
rect 13899 23792 13941 23801
rect 13899 23752 13900 23792
rect 13940 23752 13941 23792
rect 13899 23743 13941 23752
rect 14283 23792 14325 23801
rect 14283 23752 14284 23792
rect 14324 23752 14325 23792
rect 14283 23743 14325 23752
rect 14851 23792 14909 23793
rect 14851 23752 14860 23792
rect 14900 23752 14909 23792
rect 15339 23766 15340 23806
rect 15380 23766 15381 23806
rect 19419 23801 19461 23810
rect 15339 23757 15381 23766
rect 16099 23792 16157 23793
rect 14851 23751 14909 23752
rect 16099 23752 16108 23792
rect 16148 23752 16157 23792
rect 16099 23751 16157 23752
rect 17347 23792 17405 23793
rect 17347 23752 17356 23792
rect 17396 23752 17405 23792
rect 17347 23751 17405 23752
rect 17835 23792 17877 23801
rect 17835 23752 17836 23792
rect 17876 23752 17877 23792
rect 17835 23743 17877 23752
rect 17931 23792 17973 23801
rect 17931 23752 17932 23792
rect 17972 23752 17973 23792
rect 17931 23743 17973 23752
rect 18315 23792 18357 23801
rect 18315 23752 18316 23792
rect 18356 23752 18357 23792
rect 18315 23743 18357 23752
rect 18883 23792 18941 23793
rect 18883 23752 18892 23792
rect 18932 23752 18941 23792
rect 19419 23761 19420 23801
rect 19460 23761 19461 23801
rect 19419 23752 19461 23761
rect 18883 23751 18941 23752
rect 2859 23722 2901 23731
rect 10443 23708 10485 23717
rect 10443 23668 10444 23708
rect 10484 23668 10485 23708
rect 10443 23659 10485 23668
rect 17547 23708 17589 23717
rect 17547 23668 17548 23708
rect 17588 23668 17589 23708
rect 17547 23659 17589 23668
rect 3139 23624 3197 23625
rect 3139 23584 3148 23624
rect 3188 23584 3197 23624
rect 3139 23583 3197 23584
rect 3619 23624 3677 23625
rect 3619 23584 3628 23624
rect 3668 23584 3677 23624
rect 3619 23583 3677 23584
rect 3819 23624 3861 23633
rect 3819 23584 3820 23624
rect 3860 23584 3861 23624
rect 3819 23575 3861 23584
rect 4875 23624 4917 23633
rect 4875 23584 4876 23624
rect 4916 23584 4917 23624
rect 4875 23575 4917 23584
rect 5251 23624 5309 23625
rect 5251 23584 5260 23624
rect 5300 23584 5309 23624
rect 5251 23583 5309 23584
rect 7083 23624 7125 23633
rect 7083 23584 7084 23624
rect 7124 23584 7125 23624
rect 7083 23575 7125 23584
rect 8715 23624 8757 23633
rect 8715 23584 8716 23624
rect 8756 23584 8757 23624
rect 8715 23575 8757 23584
rect 12459 23624 12501 23633
rect 12459 23584 12460 23624
rect 12500 23584 12501 23624
rect 12459 23575 12501 23584
rect 15531 23624 15573 23633
rect 15531 23584 15532 23624
rect 15572 23584 15573 23624
rect 15531 23575 15573 23584
rect 19563 23624 19605 23633
rect 19563 23584 19564 23624
rect 19604 23584 19605 23624
rect 19563 23575 19605 23584
rect 1152 23456 20452 23480
rect 1152 23416 4928 23456
rect 4968 23416 5010 23456
rect 5050 23416 5092 23456
rect 5132 23416 5174 23456
rect 5214 23416 5256 23456
rect 5296 23416 20048 23456
rect 20088 23416 20130 23456
rect 20170 23416 20212 23456
rect 20252 23416 20294 23456
rect 20334 23416 20376 23456
rect 20416 23416 20452 23456
rect 1152 23392 20452 23416
rect 8995 23288 9053 23289
rect 8995 23248 9004 23288
rect 9044 23248 9053 23288
rect 8995 23247 9053 23248
rect 9763 23288 9821 23289
rect 9763 23248 9772 23288
rect 9812 23248 9821 23288
rect 9763 23247 9821 23248
rect 12171 23288 12213 23297
rect 12171 23248 12172 23288
rect 12212 23248 12213 23288
rect 12171 23239 12213 23248
rect 13803 23288 13845 23297
rect 13803 23248 13804 23288
rect 13844 23248 13845 23288
rect 13803 23239 13845 23248
rect 19755 23288 19797 23297
rect 19755 23248 19756 23288
rect 19796 23248 19797 23288
rect 19755 23239 19797 23248
rect 2859 23204 2901 23213
rect 2859 23164 2860 23204
rect 2900 23164 2901 23204
rect 2859 23155 2901 23164
rect 4971 23204 5013 23213
rect 4971 23164 4972 23204
rect 5012 23164 5013 23204
rect 4971 23155 5013 23164
rect 8331 23204 8373 23213
rect 8331 23164 8332 23204
rect 8372 23164 8373 23204
rect 8331 23155 8373 23164
rect 1411 23120 1469 23121
rect 1411 23080 1420 23120
rect 1460 23080 1469 23120
rect 1411 23079 1469 23080
rect 2659 23120 2717 23121
rect 2659 23080 2668 23120
rect 2708 23080 2717 23120
rect 2659 23079 2717 23080
rect 3243 23120 3285 23129
rect 3243 23080 3244 23120
rect 3284 23080 3285 23120
rect 3243 23071 3285 23080
rect 3339 23120 3381 23129
rect 3339 23080 3340 23120
rect 3380 23080 3381 23120
rect 3339 23071 3381 23080
rect 3819 23120 3861 23129
rect 3819 23080 3820 23120
rect 3860 23080 3861 23120
rect 3819 23071 3861 23080
rect 4291 23120 4349 23121
rect 4291 23080 4300 23120
rect 4340 23080 4349 23120
rect 5163 23120 5205 23129
rect 4291 23079 4349 23080
rect 4779 23106 4821 23115
rect 4779 23066 4780 23106
rect 4820 23066 4821 23106
rect 5163 23080 5164 23120
rect 5204 23080 5205 23120
rect 5163 23071 5205 23080
rect 5259 23120 5301 23129
rect 5259 23080 5260 23120
rect 5300 23080 5301 23120
rect 5259 23071 5301 23080
rect 5355 23120 5397 23129
rect 5355 23080 5356 23120
rect 5396 23080 5397 23120
rect 5355 23071 5397 23080
rect 5451 23120 5493 23129
rect 5451 23080 5452 23120
rect 5492 23080 5493 23120
rect 5451 23071 5493 23080
rect 5643 23120 5685 23129
rect 5643 23080 5644 23120
rect 5684 23080 5685 23120
rect 5643 23071 5685 23080
rect 5931 23120 5973 23129
rect 5931 23080 5932 23120
rect 5972 23080 5973 23120
rect 5931 23071 5973 23080
rect 6123 23120 6165 23129
rect 6123 23080 6124 23120
rect 6164 23080 6165 23120
rect 6123 23071 6165 23080
rect 6307 23120 6365 23121
rect 6307 23080 6316 23120
rect 6356 23080 6365 23120
rect 6307 23079 6365 23080
rect 6603 23120 6645 23129
rect 6603 23080 6604 23120
rect 6644 23080 6645 23120
rect 6603 23071 6645 23080
rect 6699 23120 6741 23129
rect 6699 23080 6700 23120
rect 6740 23080 6741 23120
rect 6699 23071 6741 23080
rect 7651 23120 7709 23121
rect 7651 23080 7660 23120
rect 7700 23080 7709 23120
rect 7651 23079 7709 23080
rect 8139 23115 8181 23124
rect 8139 23075 8140 23115
rect 8180 23075 8181 23115
rect 8139 23066 8181 23075
rect 8523 23120 8565 23129
rect 8523 23080 8524 23120
rect 8564 23080 8565 23120
rect 8523 23071 8565 23080
rect 8619 23120 8661 23129
rect 8619 23080 8620 23120
rect 8660 23080 8661 23120
rect 8619 23071 8661 23080
rect 8715 23120 8757 23129
rect 8715 23080 8716 23120
rect 8756 23080 8757 23120
rect 8715 23071 8757 23080
rect 8811 23120 8853 23129
rect 8811 23080 8812 23120
rect 8852 23080 8853 23120
rect 8811 23071 8853 23080
rect 9195 23120 9237 23129
rect 9195 23080 9196 23120
rect 9236 23080 9237 23120
rect 9195 23071 9237 23080
rect 9291 23120 9333 23129
rect 9291 23080 9292 23120
rect 9332 23080 9333 23120
rect 9291 23071 9333 23080
rect 9483 23120 9525 23129
rect 9483 23080 9484 23120
rect 9524 23080 9525 23120
rect 9483 23071 9525 23080
rect 9579 23120 9621 23129
rect 9579 23080 9580 23120
rect 9620 23080 9621 23120
rect 9579 23071 9621 23080
rect 9675 23120 9717 23129
rect 9675 23080 9676 23120
rect 9716 23080 9717 23120
rect 9675 23071 9717 23080
rect 10723 23120 10781 23121
rect 10723 23080 10732 23120
rect 10772 23080 10781 23120
rect 10723 23079 10781 23080
rect 11971 23120 12029 23121
rect 11971 23080 11980 23120
rect 12020 23080 12029 23120
rect 11971 23079 12029 23080
rect 12355 23120 12413 23121
rect 12355 23080 12364 23120
rect 12404 23080 12413 23120
rect 12355 23079 12413 23080
rect 13603 23120 13661 23121
rect 13603 23080 13612 23120
rect 13652 23080 13661 23120
rect 13603 23079 13661 23080
rect 18307 23120 18365 23121
rect 18307 23080 18316 23120
rect 18356 23080 18365 23120
rect 18307 23079 18365 23080
rect 19555 23120 19613 23121
rect 19555 23080 19564 23120
rect 19604 23080 19613 23120
rect 19555 23079 19613 23080
rect 4779 23057 4821 23066
rect 3723 23036 3765 23045
rect 3723 22996 3724 23036
rect 3764 22996 3765 23036
rect 3723 22987 3765 22996
rect 7083 23036 7125 23045
rect 7083 22996 7084 23036
rect 7124 22996 7125 23036
rect 7083 22987 7125 22996
rect 7179 23036 7221 23045
rect 7179 22996 7180 23036
rect 7220 22996 7221 23036
rect 7179 22987 7221 22996
rect 19939 23036 19997 23037
rect 19939 22996 19948 23036
rect 19988 22996 19997 23036
rect 19939 22995 19997 22996
rect 5643 22868 5685 22877
rect 5643 22828 5644 22868
rect 5684 22828 5685 22868
rect 5643 22819 5685 22828
rect 6219 22868 6261 22877
rect 6219 22828 6220 22868
rect 6260 22828 6261 22868
rect 6219 22819 6261 22828
rect 20139 22868 20181 22877
rect 20139 22828 20140 22868
rect 20180 22828 20181 22868
rect 20139 22819 20181 22828
rect 1152 22700 20352 22724
rect 1152 22660 3688 22700
rect 3728 22660 3770 22700
rect 3810 22660 3852 22700
rect 3892 22660 3934 22700
rect 3974 22660 4016 22700
rect 4056 22660 18808 22700
rect 18848 22660 18890 22700
rect 18930 22660 18972 22700
rect 19012 22660 19054 22700
rect 19094 22660 19136 22700
rect 19176 22660 20352 22700
rect 1152 22636 20352 22660
rect 4491 22532 4533 22541
rect 4491 22492 4492 22532
rect 4532 22492 4533 22532
rect 4491 22483 4533 22492
rect 7947 22532 7989 22541
rect 7947 22492 7948 22532
rect 7988 22492 7989 22532
rect 7947 22483 7989 22492
rect 19947 22532 19989 22541
rect 19947 22492 19948 22532
rect 19988 22492 19989 22532
rect 19947 22483 19989 22492
rect 4675 22448 4733 22449
rect 4675 22408 4684 22448
rect 4724 22408 4733 22448
rect 4675 22407 4733 22408
rect 10539 22364 10581 22373
rect 10539 22324 10540 22364
rect 10580 22324 10581 22364
rect 10539 22315 10581 22324
rect 18979 22364 19037 22365
rect 18979 22324 18988 22364
rect 19028 22324 19037 22364
rect 18979 22323 19037 22324
rect 19363 22364 19421 22365
rect 19363 22324 19372 22364
rect 19412 22324 19421 22364
rect 19363 22323 19421 22324
rect 19747 22364 19805 22365
rect 19747 22324 19756 22364
rect 19796 22324 19805 22364
rect 19747 22323 19805 22324
rect 14755 22301 14813 22302
rect 11011 22293 11069 22294
rect 1411 22280 1469 22281
rect 1411 22240 1420 22280
rect 1460 22240 1469 22280
rect 1411 22239 1469 22240
rect 2659 22280 2717 22281
rect 2659 22240 2668 22280
rect 2708 22240 2717 22280
rect 2659 22239 2717 22240
rect 3043 22280 3101 22281
rect 3043 22240 3052 22280
rect 3092 22240 3101 22280
rect 3043 22239 3101 22240
rect 4291 22280 4349 22281
rect 4291 22240 4300 22280
rect 4340 22240 4349 22280
rect 4291 22239 4349 22240
rect 4971 22280 5013 22289
rect 4971 22240 4972 22280
rect 5012 22240 5013 22280
rect 4971 22231 5013 22240
rect 5067 22280 5109 22289
rect 5067 22240 5068 22280
rect 5108 22240 5109 22280
rect 5067 22231 5109 22240
rect 5347 22280 5405 22281
rect 5347 22240 5356 22280
rect 5396 22240 5405 22280
rect 5347 22239 5405 22240
rect 6987 22280 7029 22289
rect 6987 22240 6988 22280
rect 7028 22240 7029 22280
rect 6987 22231 7029 22240
rect 7083 22280 7125 22289
rect 7083 22240 7084 22280
rect 7124 22240 7125 22280
rect 7083 22231 7125 22240
rect 7659 22280 7701 22289
rect 7659 22240 7660 22280
rect 7700 22240 7701 22280
rect 7659 22231 7701 22240
rect 7755 22280 7797 22289
rect 7755 22240 7756 22280
rect 7796 22240 7797 22280
rect 7755 22231 7797 22240
rect 8227 22280 8285 22281
rect 8227 22240 8236 22280
rect 8276 22240 8285 22280
rect 8227 22239 8285 22240
rect 9475 22280 9533 22281
rect 9475 22240 9484 22280
rect 9524 22240 9533 22280
rect 9475 22239 9533 22240
rect 9963 22280 10005 22289
rect 9963 22240 9964 22280
rect 10004 22240 10005 22280
rect 9963 22231 10005 22240
rect 10059 22280 10101 22289
rect 10059 22240 10060 22280
rect 10100 22240 10101 22280
rect 10059 22231 10101 22240
rect 10443 22280 10485 22289
rect 10443 22240 10444 22280
rect 10484 22240 10485 22280
rect 11011 22253 11020 22293
rect 11060 22253 11069 22293
rect 11011 22252 11069 22253
rect 11499 22285 11541 22294
rect 10443 22231 10485 22240
rect 11499 22245 11500 22285
rect 11540 22245 11541 22285
rect 11499 22236 11541 22245
rect 11875 22280 11933 22281
rect 11875 22240 11884 22280
rect 11924 22240 11933 22280
rect 11875 22239 11933 22240
rect 13123 22280 13181 22281
rect 13123 22240 13132 22280
rect 13172 22240 13181 22280
rect 13123 22239 13181 22240
rect 13507 22280 13565 22281
rect 13507 22240 13516 22280
rect 13556 22240 13565 22280
rect 14755 22261 14764 22301
rect 14804 22261 14813 22301
rect 14755 22260 14813 22261
rect 15235 22280 15293 22281
rect 13507 22239 13565 22240
rect 15235 22240 15244 22280
rect 15284 22240 15293 22280
rect 15235 22239 15293 22240
rect 16483 22280 16541 22281
rect 16483 22240 16492 22280
rect 16532 22240 16541 22280
rect 16483 22239 16541 22240
rect 17155 22280 17213 22281
rect 17155 22240 17164 22280
rect 17204 22240 17213 22280
rect 17155 22239 17213 22240
rect 18403 22280 18461 22281
rect 18403 22240 18412 22280
rect 18452 22240 18461 22280
rect 18403 22239 18461 22240
rect 2859 22196 2901 22205
rect 2859 22156 2860 22196
rect 2900 22156 2901 22196
rect 2859 22147 2901 22156
rect 9675 22196 9717 22205
rect 9675 22156 9676 22196
rect 9716 22156 9717 22196
rect 9675 22147 9717 22156
rect 11691 22196 11733 22205
rect 11691 22156 11692 22196
rect 11732 22156 11733 22196
rect 11691 22147 11733 22156
rect 7267 22112 7325 22113
rect 7267 22072 7276 22112
rect 7316 22072 7325 22112
rect 7267 22071 7325 22072
rect 7651 22112 7709 22113
rect 7651 22072 7660 22112
rect 7700 22072 7709 22112
rect 7651 22071 7709 22072
rect 13323 22112 13365 22121
rect 13323 22072 13324 22112
rect 13364 22072 13365 22112
rect 13323 22063 13365 22072
rect 14955 22112 14997 22121
rect 14955 22072 14956 22112
rect 14996 22072 14997 22112
rect 14955 22063 14997 22072
rect 16683 22112 16725 22121
rect 16683 22072 16684 22112
rect 16724 22072 16725 22112
rect 16683 22063 16725 22072
rect 18603 22112 18645 22121
rect 18603 22072 18604 22112
rect 18644 22072 18645 22112
rect 18603 22063 18645 22072
rect 19179 22112 19221 22121
rect 19179 22072 19180 22112
rect 19220 22072 19221 22112
rect 19179 22063 19221 22072
rect 19563 22112 19605 22121
rect 19563 22072 19564 22112
rect 19604 22072 19605 22112
rect 19563 22063 19605 22072
rect 1152 21944 20452 21968
rect 1152 21904 4928 21944
rect 4968 21904 5010 21944
rect 5050 21904 5092 21944
rect 5132 21904 5174 21944
rect 5214 21904 5256 21944
rect 5296 21904 20048 21944
rect 20088 21904 20130 21944
rect 20170 21904 20212 21944
rect 20252 21904 20294 21944
rect 20334 21904 20376 21944
rect 20416 21904 20452 21944
rect 1152 21880 20452 21904
rect 7083 21776 7125 21785
rect 7083 21736 7084 21776
rect 7124 21736 7125 21776
rect 7083 21727 7125 21736
rect 9195 21776 9237 21785
rect 9195 21736 9196 21776
rect 9236 21736 9237 21776
rect 9195 21727 9237 21736
rect 11307 21776 11349 21785
rect 11307 21736 11308 21776
rect 11348 21736 11349 21776
rect 11307 21727 11349 21736
rect 14571 21692 14613 21701
rect 14571 21652 14572 21692
rect 14612 21652 14613 21692
rect 14571 21643 14613 21652
rect 18699 21692 18741 21701
rect 18699 21652 18700 21692
rect 18740 21652 18741 21692
rect 18699 21643 18741 21652
rect 3243 21608 3285 21617
rect 3243 21568 3244 21608
rect 3284 21568 3285 21608
rect 3243 21559 3285 21568
rect 3339 21608 3381 21617
rect 3339 21568 3340 21608
rect 3380 21568 3381 21608
rect 3339 21559 3381 21568
rect 3619 21608 3677 21609
rect 3619 21568 3628 21608
rect 3668 21568 3677 21608
rect 3619 21567 3677 21568
rect 4003 21608 4061 21609
rect 4003 21568 4012 21608
rect 4052 21568 4061 21608
rect 4003 21567 4061 21568
rect 5251 21608 5309 21609
rect 5251 21568 5260 21608
rect 5300 21568 5309 21608
rect 5251 21567 5309 21568
rect 5635 21608 5693 21609
rect 5635 21568 5644 21608
rect 5684 21568 5693 21608
rect 5635 21567 5693 21568
rect 6883 21608 6941 21609
rect 6883 21568 6892 21608
rect 6932 21568 6941 21608
rect 6883 21567 6941 21568
rect 7467 21608 7509 21617
rect 7467 21568 7468 21608
rect 7508 21568 7509 21608
rect 7467 21559 7509 21568
rect 7563 21608 7605 21617
rect 7563 21568 7564 21608
rect 7604 21568 7605 21608
rect 7563 21559 7605 21568
rect 7947 21608 7989 21617
rect 7947 21568 7948 21608
rect 7988 21568 7989 21608
rect 7947 21559 7989 21568
rect 8043 21608 8085 21617
rect 8043 21568 8044 21608
rect 8084 21568 8085 21608
rect 8043 21559 8085 21568
rect 8515 21608 8573 21609
rect 8515 21568 8524 21608
rect 8564 21568 8573 21608
rect 9859 21608 9917 21609
rect 8515 21567 8573 21568
rect 9003 21594 9045 21603
rect 9003 21554 9004 21594
rect 9044 21554 9045 21594
rect 9859 21568 9868 21608
rect 9908 21568 9917 21608
rect 9859 21567 9917 21568
rect 11107 21608 11165 21609
rect 11107 21568 11116 21608
rect 11156 21568 11165 21608
rect 11107 21567 11165 21568
rect 12451 21608 12509 21609
rect 12451 21568 12460 21608
rect 12500 21568 12509 21608
rect 12451 21567 12509 21568
rect 12843 21608 12885 21617
rect 12843 21568 12844 21608
rect 12884 21568 12885 21608
rect 12843 21559 12885 21568
rect 12939 21608 12981 21617
rect 12939 21568 12940 21608
rect 12980 21568 12981 21608
rect 12939 21559 12981 21568
rect 13323 21608 13365 21617
rect 13323 21568 13324 21608
rect 13364 21568 13365 21608
rect 13323 21559 13365 21568
rect 13419 21608 13461 21617
rect 13419 21568 13420 21608
rect 13460 21568 13461 21608
rect 13419 21559 13461 21568
rect 13891 21608 13949 21609
rect 13891 21568 13900 21608
rect 13940 21568 13949 21608
rect 14851 21608 14909 21609
rect 13891 21567 13949 21568
rect 14379 21598 14421 21607
rect 9003 21545 9045 21554
rect 14379 21558 14380 21598
rect 14420 21558 14421 21598
rect 14851 21568 14860 21608
rect 14900 21568 14909 21608
rect 14851 21567 14909 21568
rect 16099 21608 16157 21609
rect 16099 21568 16108 21608
rect 16148 21568 16157 21608
rect 16099 21567 16157 21568
rect 16971 21608 17013 21617
rect 16971 21568 16972 21608
rect 17012 21568 17013 21608
rect 16971 21559 17013 21568
rect 17067 21608 17109 21617
rect 17067 21568 17068 21608
rect 17108 21568 17109 21608
rect 17067 21559 17109 21568
rect 17451 21608 17493 21617
rect 17451 21568 17452 21608
rect 17492 21568 17493 21608
rect 17451 21559 17493 21568
rect 18019 21608 18077 21609
rect 18019 21568 18028 21608
rect 18068 21568 18077 21608
rect 18019 21567 18077 21568
rect 18555 21598 18597 21607
rect 14379 21549 14421 21558
rect 18555 21558 18556 21598
rect 18596 21558 18597 21598
rect 18555 21549 18597 21558
rect 17547 21524 17589 21533
rect 17547 21484 17548 21524
rect 17588 21484 17589 21524
rect 17547 21475 17589 21484
rect 18979 21524 19037 21525
rect 18979 21484 18988 21524
rect 19028 21484 19037 21524
rect 18979 21483 19037 21484
rect 19363 21524 19421 21525
rect 19363 21484 19372 21524
rect 19412 21484 19421 21524
rect 19363 21483 19421 21484
rect 16299 21440 16341 21449
rect 16299 21400 16300 21440
rect 16340 21400 16341 21440
rect 16299 21391 16341 21400
rect 19563 21440 19605 21449
rect 19563 21400 19564 21440
rect 19604 21400 19605 21440
rect 19563 21391 19605 21400
rect 2947 21356 3005 21357
rect 2947 21316 2956 21356
rect 2996 21316 3005 21356
rect 2947 21315 3005 21316
rect 5451 21356 5493 21365
rect 5451 21316 5452 21356
rect 5492 21316 5493 21356
rect 5451 21307 5493 21316
rect 12555 21356 12597 21365
rect 12555 21316 12556 21356
rect 12596 21316 12597 21356
rect 12555 21307 12597 21316
rect 19179 21356 19221 21365
rect 19179 21316 19180 21356
rect 19220 21316 19221 21356
rect 19179 21307 19221 21316
rect 1152 21188 20352 21212
rect 1152 21148 3688 21188
rect 3728 21148 3770 21188
rect 3810 21148 3852 21188
rect 3892 21148 3934 21188
rect 3974 21148 4016 21188
rect 4056 21148 18808 21188
rect 18848 21148 18890 21188
rect 18930 21148 18972 21188
rect 19012 21148 19054 21188
rect 19094 21148 19136 21188
rect 19176 21148 20352 21188
rect 1152 21124 20352 21148
rect 9483 21020 9525 21029
rect 9483 20980 9484 21020
rect 9524 20980 9525 21020
rect 9483 20971 9525 20980
rect 4587 20852 4629 20861
rect 4587 20812 4588 20852
rect 4628 20812 4629 20852
rect 4587 20803 4629 20812
rect 4683 20852 4725 20861
rect 4683 20812 4684 20852
rect 4724 20812 4725 20852
rect 4683 20803 4725 20812
rect 15339 20852 15381 20861
rect 15339 20812 15340 20852
rect 15380 20812 15381 20852
rect 15339 20803 15381 20812
rect 18123 20852 18165 20861
rect 18123 20812 18124 20852
rect 18164 20812 18165 20852
rect 18123 20803 18165 20812
rect 19459 20852 19517 20853
rect 19459 20812 19468 20852
rect 19508 20812 19517 20852
rect 19459 20811 19517 20812
rect 19843 20852 19901 20853
rect 19843 20812 19852 20852
rect 19892 20812 19901 20852
rect 19843 20811 19901 20812
rect 16395 20782 16437 20791
rect 3627 20773 3669 20782
rect 1603 20768 1661 20769
rect 1603 20728 1612 20768
rect 1652 20728 1661 20768
rect 1603 20727 1661 20728
rect 2851 20768 2909 20769
rect 2851 20728 2860 20768
rect 2900 20728 2909 20768
rect 2851 20727 2909 20728
rect 3627 20733 3628 20773
rect 3668 20733 3669 20773
rect 3627 20724 3669 20733
rect 4099 20768 4157 20769
rect 4099 20728 4108 20768
rect 4148 20728 4157 20768
rect 4099 20727 4157 20728
rect 5067 20768 5109 20777
rect 5067 20728 5068 20768
rect 5108 20728 5109 20768
rect 5067 20719 5109 20728
rect 5163 20768 5205 20777
rect 5163 20728 5164 20768
rect 5204 20728 5205 20768
rect 5163 20719 5205 20728
rect 6123 20768 6165 20777
rect 6123 20728 6124 20768
rect 6164 20728 6165 20768
rect 6123 20719 6165 20728
rect 6219 20768 6261 20777
rect 6219 20728 6220 20768
rect 6260 20728 6261 20768
rect 6219 20719 6261 20728
rect 6603 20768 6645 20777
rect 6603 20728 6604 20768
rect 6644 20728 6645 20768
rect 6603 20719 6645 20728
rect 6699 20768 6741 20777
rect 7659 20773 7701 20782
rect 6699 20728 6700 20768
rect 6740 20728 6741 20768
rect 6699 20719 6741 20728
rect 7171 20768 7229 20769
rect 7171 20728 7180 20768
rect 7220 20728 7229 20768
rect 7171 20727 7229 20728
rect 7659 20733 7660 20773
rect 7700 20733 7701 20773
rect 7659 20724 7701 20733
rect 8035 20768 8093 20769
rect 8035 20728 8044 20768
rect 8084 20728 8093 20768
rect 8035 20727 8093 20728
rect 9283 20768 9341 20769
rect 9283 20728 9292 20768
rect 9332 20728 9341 20768
rect 9283 20727 9341 20728
rect 11011 20768 11069 20769
rect 11011 20728 11020 20768
rect 11060 20728 11069 20768
rect 11011 20727 11069 20728
rect 12259 20768 12317 20769
rect 12259 20728 12268 20768
rect 12308 20728 12317 20768
rect 12259 20727 12317 20728
rect 12651 20768 12693 20777
rect 12651 20728 12652 20768
rect 12692 20728 12693 20768
rect 12651 20719 12693 20728
rect 12843 20768 12885 20777
rect 12843 20728 12844 20768
rect 12884 20728 12885 20768
rect 12843 20719 12885 20728
rect 12939 20768 12981 20777
rect 12939 20728 12940 20768
rect 12980 20728 12981 20768
rect 12939 20719 12981 20728
rect 13123 20768 13181 20769
rect 13123 20728 13132 20768
rect 13172 20728 13181 20768
rect 13123 20727 13181 20728
rect 14371 20768 14429 20769
rect 14371 20728 14380 20768
rect 14420 20728 14429 20768
rect 14371 20727 14429 20728
rect 14859 20768 14901 20777
rect 14859 20728 14860 20768
rect 14900 20728 14901 20768
rect 14859 20719 14901 20728
rect 14955 20768 14997 20777
rect 14955 20728 14956 20768
rect 14996 20728 14997 20768
rect 14955 20719 14997 20728
rect 15435 20768 15477 20777
rect 15435 20728 15436 20768
rect 15476 20728 15477 20768
rect 15435 20719 15477 20728
rect 15907 20768 15965 20769
rect 15907 20728 15916 20768
rect 15956 20728 15965 20768
rect 16395 20742 16396 20782
rect 16436 20742 16437 20782
rect 19131 20777 19173 20786
rect 16395 20733 16437 20742
rect 17547 20768 17589 20777
rect 15907 20727 15965 20728
rect 17547 20728 17548 20768
rect 17588 20728 17589 20768
rect 17547 20719 17589 20728
rect 17643 20768 17685 20777
rect 17643 20728 17644 20768
rect 17684 20728 17685 20768
rect 17643 20719 17685 20728
rect 18027 20768 18069 20777
rect 18027 20728 18028 20768
rect 18068 20728 18069 20768
rect 18027 20719 18069 20728
rect 18595 20768 18653 20769
rect 18595 20728 18604 20768
rect 18644 20728 18653 20768
rect 19131 20737 19132 20777
rect 19172 20737 19173 20777
rect 19131 20728 19173 20737
rect 18595 20727 18653 20728
rect 3051 20684 3093 20693
rect 3051 20644 3052 20684
rect 3092 20644 3093 20684
rect 3051 20635 3093 20644
rect 3435 20684 3477 20693
rect 3435 20644 3436 20684
rect 3476 20644 3477 20684
rect 3435 20635 3477 20644
rect 14571 20684 14613 20693
rect 14571 20644 14572 20684
rect 14612 20644 14613 20684
rect 14571 20635 14613 20644
rect 16587 20684 16629 20693
rect 16587 20644 16588 20684
rect 16628 20644 16629 20684
rect 16587 20635 16629 20644
rect 7851 20600 7893 20609
rect 7851 20560 7852 20600
rect 7892 20560 7893 20600
rect 7851 20551 7893 20560
rect 12459 20600 12501 20609
rect 12459 20560 12460 20600
rect 12500 20560 12501 20600
rect 12459 20551 12501 20560
rect 12747 20600 12789 20609
rect 12747 20560 12748 20600
rect 12788 20560 12789 20600
rect 12747 20551 12789 20560
rect 19275 20600 19317 20609
rect 19275 20560 19276 20600
rect 19316 20560 19317 20600
rect 19275 20551 19317 20560
rect 19659 20600 19701 20609
rect 19659 20560 19660 20600
rect 19700 20560 19701 20600
rect 19659 20551 19701 20560
rect 20043 20600 20085 20609
rect 20043 20560 20044 20600
rect 20084 20560 20085 20600
rect 20043 20551 20085 20560
rect 1152 20432 20452 20456
rect 1152 20392 4928 20432
rect 4968 20392 5010 20432
rect 5050 20392 5092 20432
rect 5132 20392 5174 20432
rect 5214 20392 5256 20432
rect 5296 20392 20048 20432
rect 20088 20392 20130 20432
rect 20170 20392 20212 20432
rect 20252 20392 20294 20432
rect 20334 20392 20376 20432
rect 20416 20392 20452 20432
rect 1152 20368 20452 20392
rect 12171 20264 12213 20273
rect 12171 20224 12172 20264
rect 12212 20224 12213 20264
rect 12171 20215 12213 20224
rect 15427 20264 15485 20265
rect 15427 20224 15436 20264
rect 15476 20224 15485 20264
rect 15427 20223 15485 20224
rect 17259 20264 17301 20273
rect 17259 20224 17260 20264
rect 17300 20224 17301 20264
rect 17259 20215 17301 20224
rect 6795 20180 6837 20189
rect 6795 20140 6796 20180
rect 6836 20140 6837 20180
rect 6795 20131 6837 20140
rect 10443 20180 10485 20189
rect 10443 20140 10444 20180
rect 10484 20140 10485 20180
rect 10443 20131 10485 20140
rect 19659 20180 19701 20189
rect 19659 20140 19660 20180
rect 19700 20140 19701 20180
rect 19659 20131 19701 20140
rect 1507 20096 1565 20097
rect 1507 20056 1516 20096
rect 1556 20056 1565 20096
rect 1507 20055 1565 20056
rect 2755 20096 2813 20097
rect 2755 20056 2764 20096
rect 2804 20056 2813 20096
rect 2755 20055 2813 20056
rect 3243 20096 3285 20105
rect 3243 20056 3244 20096
rect 3284 20056 3285 20096
rect 3243 20047 3285 20056
rect 3339 20096 3381 20105
rect 3339 20056 3340 20096
rect 3380 20056 3381 20096
rect 3339 20047 3381 20056
rect 3531 20096 3573 20105
rect 3531 20056 3532 20096
rect 3572 20056 3573 20096
rect 3531 20047 3573 20056
rect 3915 20096 3957 20105
rect 3915 20056 3916 20096
rect 3956 20056 3957 20096
rect 3915 20047 3957 20056
rect 4011 20096 4053 20105
rect 4011 20056 4012 20096
rect 4052 20056 4053 20096
rect 4011 20047 4053 20056
rect 4107 20096 4149 20105
rect 4107 20056 4108 20096
rect 4148 20056 4149 20096
rect 4107 20047 4149 20056
rect 4395 20096 4437 20105
rect 4395 20056 4396 20096
rect 4436 20056 4437 20096
rect 4395 20047 4437 20056
rect 4587 20096 4629 20105
rect 4587 20056 4588 20096
rect 4628 20056 4629 20096
rect 4587 20047 4629 20056
rect 4675 20096 4733 20097
rect 4675 20056 4684 20096
rect 4724 20056 4733 20096
rect 4675 20055 4733 20056
rect 5347 20096 5405 20097
rect 5347 20056 5356 20096
rect 5396 20056 5405 20096
rect 5347 20055 5405 20056
rect 6595 20096 6653 20097
rect 6595 20056 6604 20096
rect 6644 20056 6653 20096
rect 6595 20055 6653 20056
rect 6979 20096 7037 20097
rect 6979 20056 6988 20096
rect 7028 20056 7037 20096
rect 6979 20055 7037 20056
rect 8227 20096 8285 20097
rect 8227 20056 8236 20096
rect 8276 20056 8285 20096
rect 8227 20055 8285 20056
rect 8715 20096 8757 20105
rect 8715 20056 8716 20096
rect 8756 20056 8757 20096
rect 8715 20047 8757 20056
rect 8811 20096 8853 20105
rect 8811 20056 8812 20096
rect 8852 20056 8853 20096
rect 8811 20047 8853 20056
rect 9195 20096 9237 20105
rect 9195 20056 9196 20096
rect 9236 20056 9237 20096
rect 9195 20047 9237 20056
rect 9763 20096 9821 20097
rect 9763 20056 9772 20096
rect 9812 20056 9821 20096
rect 10723 20096 10781 20097
rect 9763 20055 9821 20056
rect 10299 20054 10341 20063
rect 10723 20056 10732 20096
rect 10772 20056 10781 20096
rect 10723 20055 10781 20056
rect 11971 20096 12029 20097
rect 11971 20056 11980 20096
rect 12020 20056 12029 20096
rect 11971 20055 12029 20056
rect 12446 20096 12504 20097
rect 12446 20056 12455 20096
rect 12495 20056 12504 20096
rect 12446 20055 12504 20056
rect 12555 20096 12597 20105
rect 12555 20056 12556 20096
rect 12596 20056 12597 20096
rect 9291 20012 9333 20021
rect 9291 19972 9292 20012
rect 9332 19972 9333 20012
rect 10299 20014 10300 20054
rect 10340 20014 10341 20054
rect 12555 20047 12597 20056
rect 12651 20096 12693 20105
rect 12651 20056 12652 20096
rect 12692 20056 12693 20096
rect 12651 20047 12693 20056
rect 12835 20096 12893 20097
rect 12835 20056 12844 20096
rect 12884 20056 12893 20096
rect 12835 20055 12893 20056
rect 12931 20096 12989 20097
rect 12931 20056 12940 20096
rect 12980 20056 12989 20096
rect 12931 20055 12989 20056
rect 13699 20096 13757 20097
rect 13699 20056 13708 20096
rect 13748 20056 13757 20096
rect 13699 20055 13757 20056
rect 14947 20096 15005 20097
rect 14947 20056 14956 20096
rect 14996 20056 15005 20096
rect 14947 20055 15005 20056
rect 15147 20096 15189 20105
rect 15147 20056 15148 20096
rect 15188 20056 15189 20096
rect 15147 20047 15189 20056
rect 15243 20096 15285 20105
rect 15243 20056 15244 20096
rect 15284 20056 15285 20096
rect 15243 20047 15285 20056
rect 15811 20096 15869 20097
rect 15811 20056 15820 20096
rect 15860 20056 15869 20096
rect 15811 20055 15869 20056
rect 17059 20096 17117 20097
rect 17059 20056 17068 20096
rect 17108 20056 17117 20096
rect 17059 20055 17117 20056
rect 18211 20096 18269 20097
rect 18211 20056 18220 20096
rect 18260 20056 18269 20096
rect 18211 20055 18269 20056
rect 19459 20096 19517 20097
rect 19459 20056 19468 20096
rect 19508 20056 19517 20096
rect 19459 20055 19517 20056
rect 10299 20005 10341 20014
rect 19843 20012 19901 20013
rect 9291 19963 9333 19972
rect 19843 19972 19852 20012
rect 19892 19972 19901 20012
rect 19843 19971 19901 19972
rect 2955 19928 2997 19937
rect 2955 19888 2956 19928
rect 2996 19888 2997 19928
rect 2955 19879 2997 19888
rect 8427 19928 8469 19937
rect 8427 19888 8428 19928
rect 8468 19888 8469 19928
rect 8427 19879 8469 19888
rect 20043 19928 20085 19937
rect 20043 19888 20044 19928
rect 20084 19888 20085 19928
rect 20043 19879 20085 19888
rect 3715 19844 3773 19845
rect 3715 19804 3724 19844
rect 3764 19804 3773 19844
rect 3715 19803 3773 19804
rect 4395 19844 4437 19853
rect 4395 19804 4396 19844
rect 4436 19804 4437 19844
rect 4395 19795 4437 19804
rect 12939 19844 12981 19853
rect 12939 19804 12940 19844
rect 12980 19804 12981 19844
rect 12939 19795 12981 19804
rect 13515 19844 13557 19853
rect 13515 19804 13516 19844
rect 13556 19804 13557 19844
rect 13515 19795 13557 19804
rect 1152 19676 20352 19700
rect 1152 19636 3688 19676
rect 3728 19636 3770 19676
rect 3810 19636 3852 19676
rect 3892 19636 3934 19676
rect 3974 19636 4016 19676
rect 4056 19636 18808 19676
rect 18848 19636 18890 19676
rect 18930 19636 18972 19676
rect 19012 19636 19054 19676
rect 19094 19636 19136 19676
rect 19176 19636 20352 19676
rect 1152 19612 20352 19636
rect 2667 19508 2709 19517
rect 2667 19468 2668 19508
rect 2708 19468 2709 19508
rect 2667 19459 2709 19468
rect 10347 19508 10389 19517
rect 10347 19468 10348 19508
rect 10388 19468 10389 19508
rect 10347 19459 10389 19468
rect 15051 19508 15093 19517
rect 15051 19468 15052 19508
rect 15092 19468 15093 19508
rect 15051 19459 15093 19468
rect 19563 19508 19605 19517
rect 19563 19468 19564 19508
rect 19604 19468 19605 19508
rect 19563 19459 19605 19468
rect 17547 19340 17589 19349
rect 17547 19300 17548 19340
rect 17588 19300 17589 19340
rect 17547 19291 17589 19300
rect 18979 19340 19037 19341
rect 18979 19300 18988 19340
rect 19028 19300 19037 19340
rect 18979 19299 19037 19300
rect 19363 19340 19421 19341
rect 19363 19300 19372 19340
rect 19412 19300 19421 19340
rect 19363 19299 19421 19300
rect 19747 19340 19805 19341
rect 19747 19300 19756 19340
rect 19796 19300 19805 19340
rect 19747 19299 19805 19300
rect 13227 19266 13269 19275
rect 1219 19256 1277 19257
rect 1219 19216 1228 19256
rect 1268 19216 1277 19256
rect 1219 19215 1277 19216
rect 2467 19256 2525 19257
rect 2467 19216 2476 19256
rect 2516 19216 2525 19256
rect 2467 19215 2525 19216
rect 3723 19256 3765 19265
rect 3723 19216 3724 19256
rect 3764 19216 3765 19256
rect 3723 19207 3765 19216
rect 3819 19256 3861 19265
rect 3819 19216 3820 19256
rect 3860 19216 3861 19256
rect 3819 19207 3861 19216
rect 3915 19256 3957 19265
rect 3915 19216 3916 19256
rect 3956 19216 3957 19256
rect 3915 19207 3957 19216
rect 4099 19256 4157 19257
rect 4099 19216 4108 19256
rect 4148 19216 4157 19256
rect 4099 19215 4157 19216
rect 5347 19256 5405 19257
rect 5347 19216 5356 19256
rect 5396 19216 5405 19256
rect 5347 19215 5405 19216
rect 7267 19256 7325 19257
rect 7267 19216 7276 19256
rect 7316 19216 7325 19256
rect 7267 19215 7325 19216
rect 8515 19256 8573 19257
rect 8515 19216 8524 19256
rect 8564 19216 8573 19256
rect 8515 19215 8573 19216
rect 8899 19256 8957 19257
rect 8899 19216 8908 19256
rect 8948 19216 8957 19256
rect 8899 19215 8957 19216
rect 10147 19256 10205 19257
rect 10147 19216 10156 19256
rect 10196 19216 10205 19256
rect 10147 19215 10205 19216
rect 11587 19256 11645 19257
rect 11587 19216 11596 19256
rect 11636 19216 11645 19256
rect 11587 19215 11645 19216
rect 12835 19256 12893 19257
rect 12835 19216 12844 19256
rect 12884 19216 12893 19256
rect 13227 19226 13228 19266
rect 13268 19226 13269 19266
rect 18555 19265 18597 19274
rect 13227 19217 13269 19226
rect 13323 19256 13365 19265
rect 12835 19215 12893 19216
rect 13323 19216 13324 19256
rect 13364 19216 13365 19256
rect 13323 19207 13365 19216
rect 13891 19256 13949 19257
rect 13891 19216 13900 19256
rect 13940 19216 13949 19256
rect 13891 19215 13949 19216
rect 14283 19256 14325 19265
rect 14283 19216 14284 19256
rect 14324 19216 14325 19256
rect 14283 19207 14325 19216
rect 14379 19256 14421 19265
rect 14379 19216 14380 19256
rect 14420 19216 14421 19256
rect 14379 19207 14421 19216
rect 14659 19256 14717 19257
rect 14659 19216 14668 19256
rect 14708 19216 14717 19256
rect 14659 19215 14717 19216
rect 14763 19256 14805 19265
rect 14763 19216 14764 19256
rect 14804 19216 14805 19256
rect 14763 19207 14805 19216
rect 15235 19256 15293 19257
rect 15235 19216 15244 19256
rect 15284 19216 15293 19256
rect 15235 19215 15293 19216
rect 16483 19256 16541 19257
rect 16483 19216 16492 19256
rect 16532 19216 16541 19256
rect 16483 19215 16541 19216
rect 16971 19256 17013 19265
rect 16971 19216 16972 19256
rect 17012 19216 17013 19256
rect 16971 19207 17013 19216
rect 17067 19256 17109 19265
rect 17067 19216 17068 19256
rect 17108 19216 17109 19256
rect 17067 19207 17109 19216
rect 17451 19256 17493 19265
rect 17451 19216 17452 19256
rect 17492 19216 17493 19256
rect 17451 19207 17493 19216
rect 18019 19256 18077 19257
rect 18019 19216 18028 19256
rect 18068 19216 18077 19256
rect 18555 19225 18556 19265
rect 18596 19225 18597 19265
rect 18555 19216 18597 19225
rect 18019 19215 18077 19216
rect 13803 19172 13845 19181
rect 13803 19132 13804 19172
rect 13844 19132 13845 19172
rect 13803 19123 13845 19132
rect 16683 19172 16725 19181
rect 16683 19132 16684 19172
rect 16724 19132 16725 19172
rect 16683 19123 16725 19132
rect 18699 19172 18741 19181
rect 18699 19132 18700 19172
rect 18740 19132 18741 19172
rect 18699 19123 18741 19132
rect 3619 19088 3677 19089
rect 3619 19048 3628 19088
rect 3668 19048 3677 19088
rect 3619 19047 3677 19048
rect 5547 19088 5589 19097
rect 5547 19048 5548 19088
rect 5588 19048 5589 19088
rect 5547 19039 5589 19048
rect 8715 19088 8757 19097
rect 8715 19048 8716 19088
rect 8756 19048 8757 19088
rect 8715 19039 8757 19048
rect 13035 19088 13077 19097
rect 13035 19048 13036 19088
rect 13076 19048 13077 19088
rect 13035 19039 13077 19048
rect 13507 19088 13565 19089
rect 13507 19048 13516 19088
rect 13556 19048 13565 19088
rect 13507 19047 13565 19048
rect 14083 19088 14141 19089
rect 14083 19048 14092 19088
rect 14132 19048 14141 19088
rect 14083 19047 14141 19048
rect 19179 19088 19221 19097
rect 19179 19048 19180 19088
rect 19220 19048 19221 19088
rect 19179 19039 19221 19048
rect 19947 19088 19989 19097
rect 19947 19048 19948 19088
rect 19988 19048 19989 19088
rect 19947 19039 19989 19048
rect 14571 19030 14613 19039
rect 14571 18990 14572 19030
rect 14612 18990 14613 19030
rect 14571 18981 14613 18990
rect 1152 18920 20452 18944
rect 1152 18880 4928 18920
rect 4968 18880 5010 18920
rect 5050 18880 5092 18920
rect 5132 18880 5174 18920
rect 5214 18880 5256 18920
rect 5296 18880 20048 18920
rect 20088 18880 20130 18920
rect 20170 18880 20212 18920
rect 20252 18880 20294 18920
rect 20334 18880 20376 18920
rect 20416 18880 20452 18920
rect 1152 18856 20452 18880
rect 4203 18752 4245 18761
rect 4203 18712 4204 18752
rect 4244 18712 4245 18752
rect 4203 18703 4245 18712
rect 13323 18752 13365 18761
rect 13323 18712 13324 18752
rect 13364 18712 13365 18752
rect 13323 18703 13365 18712
rect 14955 18752 14997 18761
rect 14955 18712 14956 18752
rect 14996 18712 14997 18752
rect 14955 18703 14997 18712
rect 15619 18752 15677 18753
rect 15619 18712 15628 18752
rect 15668 18712 15677 18752
rect 15619 18711 15677 18712
rect 7179 18668 7221 18677
rect 7179 18628 7180 18668
rect 7220 18628 7221 18668
rect 7179 18619 7221 18628
rect 11307 18668 11349 18677
rect 11307 18628 11308 18668
rect 11348 18628 11349 18668
rect 11307 18619 11349 18628
rect 17451 18668 17493 18677
rect 17451 18628 17452 18668
rect 17492 18628 17493 18668
rect 17451 18619 17493 18628
rect 19467 18668 19509 18677
rect 19467 18628 19468 18668
rect 19508 18628 19509 18668
rect 19467 18619 19509 18628
rect 2475 18584 2517 18593
rect 2475 18544 2476 18584
rect 2516 18544 2517 18584
rect 2475 18535 2517 18544
rect 2571 18584 2613 18593
rect 2571 18544 2572 18584
rect 2612 18544 2613 18584
rect 2571 18535 2613 18544
rect 3523 18584 3581 18585
rect 3523 18544 3532 18584
rect 3572 18544 3581 18584
rect 5451 18584 5493 18593
rect 3523 18543 3581 18544
rect 4011 18570 4053 18579
rect 4011 18530 4012 18570
rect 4052 18530 4053 18570
rect 5451 18544 5452 18584
rect 5492 18544 5493 18584
rect 5451 18535 5493 18544
rect 5547 18584 5589 18593
rect 5547 18544 5548 18584
rect 5588 18544 5589 18584
rect 5547 18535 5589 18544
rect 6499 18584 6557 18585
rect 6499 18544 6508 18584
rect 6548 18544 6557 18584
rect 7459 18584 7517 18585
rect 6499 18543 6557 18544
rect 6987 18570 7029 18579
rect 4011 18521 4053 18530
rect 6987 18530 6988 18570
rect 7028 18530 7029 18570
rect 7459 18544 7468 18584
rect 7508 18544 7517 18584
rect 7459 18543 7517 18544
rect 8227 18584 8285 18585
rect 8227 18544 8236 18584
rect 8276 18544 8285 18584
rect 8227 18543 8285 18544
rect 9475 18584 9533 18585
rect 9475 18544 9484 18584
rect 9524 18544 9533 18584
rect 9475 18543 9533 18544
rect 9859 18584 9917 18585
rect 9859 18544 9868 18584
rect 9908 18544 9917 18584
rect 9859 18543 9917 18544
rect 11107 18584 11165 18585
rect 11107 18544 11116 18584
rect 11156 18544 11165 18584
rect 11107 18543 11165 18544
rect 11595 18584 11637 18593
rect 11595 18544 11596 18584
rect 11636 18544 11637 18584
rect 11595 18535 11637 18544
rect 11691 18584 11733 18593
rect 11691 18544 11692 18584
rect 11732 18544 11733 18584
rect 11691 18535 11733 18544
rect 12075 18584 12117 18593
rect 12075 18544 12076 18584
rect 12116 18544 12117 18584
rect 12075 18535 12117 18544
rect 12643 18584 12701 18585
rect 12643 18544 12652 18584
rect 12692 18544 12701 18584
rect 12643 18543 12701 18544
rect 13131 18579 13173 18588
rect 13131 18539 13132 18579
rect 13172 18539 13173 18579
rect 13507 18584 13565 18585
rect 13507 18544 13516 18584
rect 13556 18544 13565 18584
rect 13507 18543 13565 18544
rect 14755 18584 14813 18585
rect 14755 18544 14764 18584
rect 14804 18544 14813 18584
rect 14755 18543 14813 18544
rect 15139 18584 15197 18585
rect 15139 18544 15148 18584
rect 15188 18544 15197 18584
rect 15139 18543 15197 18544
rect 15235 18584 15293 18585
rect 15235 18544 15244 18584
rect 15284 18544 15293 18584
rect 15235 18543 15293 18544
rect 15435 18584 15477 18593
rect 15435 18544 15436 18584
rect 15476 18544 15477 18584
rect 13131 18530 13173 18539
rect 15435 18535 15477 18544
rect 15531 18584 15573 18593
rect 15531 18544 15532 18584
rect 15572 18544 15573 18584
rect 15531 18535 15573 18544
rect 15624 18584 15682 18585
rect 15624 18544 15633 18584
rect 15673 18544 15682 18584
rect 15624 18543 15682 18544
rect 16003 18584 16061 18585
rect 16003 18544 16012 18584
rect 16052 18544 16061 18584
rect 16003 18543 16061 18544
rect 17251 18584 17309 18585
rect 17251 18544 17260 18584
rect 17300 18544 17309 18584
rect 17251 18543 17309 18544
rect 17739 18584 17781 18593
rect 17739 18544 17740 18584
rect 17780 18544 17781 18584
rect 17739 18535 17781 18544
rect 17835 18584 17877 18593
rect 17835 18544 17836 18584
rect 17876 18544 17877 18584
rect 17835 18535 17877 18544
rect 18219 18584 18261 18593
rect 18219 18544 18220 18584
rect 18260 18544 18261 18584
rect 18219 18535 18261 18544
rect 18787 18584 18845 18585
rect 18787 18544 18796 18584
rect 18836 18544 18845 18584
rect 18787 18543 18845 18544
rect 19275 18570 19317 18579
rect 19275 18530 19276 18570
rect 19316 18530 19317 18570
rect 6987 18521 7029 18530
rect 19275 18521 19317 18530
rect 2955 18500 2997 18509
rect 2955 18460 2956 18500
rect 2996 18460 2997 18500
rect 2955 18451 2997 18460
rect 3051 18500 3093 18509
rect 3051 18460 3052 18500
rect 3092 18460 3093 18500
rect 3051 18451 3093 18460
rect 5931 18500 5973 18509
rect 5931 18460 5932 18500
rect 5972 18460 5973 18500
rect 5931 18451 5973 18460
rect 6027 18500 6069 18509
rect 6027 18460 6028 18500
rect 6068 18460 6069 18500
rect 6027 18451 6069 18460
rect 12171 18500 12213 18509
rect 12171 18460 12172 18500
rect 12212 18460 12213 18500
rect 12171 18451 12213 18460
rect 18315 18500 18357 18509
rect 18315 18460 18316 18500
rect 18356 18460 18357 18500
rect 18315 18451 18357 18460
rect 19651 18500 19709 18501
rect 19651 18460 19660 18500
rect 19700 18460 19709 18500
rect 19651 18459 19709 18460
rect 20035 18500 20093 18501
rect 20035 18460 20044 18500
rect 20084 18460 20093 18500
rect 20035 18459 20093 18460
rect 19851 18416 19893 18425
rect 19851 18376 19852 18416
rect 19892 18376 19893 18416
rect 19851 18367 19893 18376
rect 7371 18332 7413 18341
rect 7371 18292 7372 18332
rect 7412 18292 7413 18332
rect 7371 18283 7413 18292
rect 9675 18332 9717 18341
rect 9675 18292 9676 18332
rect 9716 18292 9717 18332
rect 9675 18283 9717 18292
rect 14955 18332 14997 18341
rect 14955 18292 14956 18332
rect 14996 18292 14997 18332
rect 14955 18283 14997 18292
rect 20235 18332 20277 18341
rect 20235 18292 20236 18332
rect 20276 18292 20277 18332
rect 20235 18283 20277 18292
rect 1152 18164 20352 18188
rect 1152 18124 3688 18164
rect 3728 18124 3770 18164
rect 3810 18124 3852 18164
rect 3892 18124 3934 18164
rect 3974 18124 4016 18164
rect 4056 18124 18808 18164
rect 18848 18124 18890 18164
rect 18930 18124 18972 18164
rect 19012 18124 19054 18164
rect 19094 18124 19136 18164
rect 19176 18124 20352 18164
rect 1152 18100 20352 18124
rect 4011 17996 4053 18005
rect 4011 17956 4012 17996
rect 4052 17956 4053 17996
rect 4011 17947 4053 17956
rect 6699 17996 6741 18005
rect 6699 17956 6700 17996
rect 6740 17956 6741 17996
rect 6699 17947 6741 17956
rect 16011 17996 16053 18005
rect 16011 17956 16012 17996
rect 16052 17956 16053 17996
rect 16011 17947 16053 17956
rect 18699 17996 18741 18005
rect 18699 17956 18700 17996
rect 18740 17956 18741 17996
rect 18699 17947 18741 17956
rect 19075 17912 19133 17913
rect 19075 17872 19084 17912
rect 19124 17872 19133 17912
rect 19075 17871 19133 17872
rect 7659 17828 7701 17837
rect 7659 17788 7660 17828
rect 7700 17788 7701 17828
rect 7659 17779 7701 17788
rect 9675 17828 9717 17837
rect 9675 17788 9676 17828
rect 9716 17788 9717 17828
rect 9675 17779 9717 17788
rect 15243 17828 15285 17837
rect 15243 17788 15244 17828
rect 15284 17788 15285 17828
rect 15243 17779 15285 17788
rect 8763 17753 8805 17762
rect 10731 17758 10773 17767
rect 16291 17763 16349 17764
rect 2563 17744 2621 17745
rect 2563 17704 2572 17744
rect 2612 17704 2621 17744
rect 2563 17703 2621 17704
rect 3811 17744 3869 17745
rect 3811 17704 3820 17744
rect 3860 17704 3869 17744
rect 3811 17703 3869 17704
rect 5251 17744 5309 17745
rect 5251 17704 5260 17744
rect 5300 17704 5309 17744
rect 5251 17703 5309 17704
rect 6499 17744 6557 17745
rect 6499 17704 6508 17744
rect 6548 17704 6557 17744
rect 6499 17703 6557 17704
rect 7179 17744 7221 17753
rect 7179 17704 7180 17744
rect 7220 17704 7221 17744
rect 7179 17695 7221 17704
rect 7275 17744 7317 17753
rect 7275 17704 7276 17744
rect 7316 17704 7317 17744
rect 7275 17695 7317 17704
rect 7755 17744 7797 17753
rect 7755 17704 7756 17744
rect 7796 17704 7797 17744
rect 7755 17695 7797 17704
rect 8227 17744 8285 17745
rect 8227 17704 8236 17744
rect 8276 17704 8285 17744
rect 8763 17713 8764 17753
rect 8804 17713 8805 17753
rect 8763 17704 8805 17713
rect 9195 17744 9237 17753
rect 9195 17704 9196 17744
rect 9236 17704 9237 17744
rect 8227 17703 8285 17704
rect 9195 17695 9237 17704
rect 9291 17744 9333 17753
rect 9291 17704 9292 17744
rect 9332 17704 9333 17744
rect 9291 17695 9333 17704
rect 9771 17744 9813 17753
rect 9771 17704 9772 17744
rect 9812 17704 9813 17744
rect 9771 17695 9813 17704
rect 10243 17744 10301 17745
rect 10243 17704 10252 17744
rect 10292 17704 10301 17744
rect 10731 17718 10732 17758
rect 10772 17718 10773 17758
rect 14187 17753 14229 17762
rect 10731 17709 10773 17718
rect 13699 17744 13757 17745
rect 10243 17703 10301 17704
rect 13699 17704 13708 17744
rect 13748 17704 13757 17744
rect 13699 17703 13757 17704
rect 13803 17744 13845 17753
rect 13803 17704 13804 17744
rect 13844 17704 13845 17744
rect 14187 17713 14188 17753
rect 14228 17713 14229 17753
rect 14187 17704 14229 17713
rect 14659 17744 14717 17745
rect 14659 17704 14668 17744
rect 14708 17704 14717 17744
rect 13803 17695 13845 17704
rect 14659 17703 14717 17704
rect 15147 17744 15189 17753
rect 15147 17704 15148 17744
rect 15188 17704 15189 17744
rect 15147 17695 15189 17704
rect 15627 17744 15669 17753
rect 15627 17704 15628 17744
rect 15668 17704 15669 17744
rect 15627 17695 15669 17704
rect 15723 17744 15765 17753
rect 15723 17704 15724 17744
rect 15764 17704 15765 17744
rect 15723 17695 15765 17704
rect 16011 17744 16053 17753
rect 16011 17704 16012 17744
rect 16052 17704 16053 17744
rect 16011 17695 16053 17704
rect 16203 17744 16245 17753
rect 16203 17704 16204 17744
rect 16244 17704 16245 17744
rect 16291 17723 16300 17763
rect 16340 17723 16349 17763
rect 16291 17722 16349 17723
rect 17251 17744 17309 17745
rect 16203 17695 16245 17704
rect 17251 17704 17260 17744
rect 17300 17704 17309 17744
rect 17251 17703 17309 17704
rect 18499 17744 18557 17745
rect 18499 17704 18508 17744
rect 18548 17704 18557 17744
rect 18499 17703 18557 17704
rect 19467 17744 19509 17753
rect 19467 17704 19468 17744
rect 19508 17704 19509 17744
rect 19467 17695 19509 17704
rect 19747 17744 19805 17745
rect 19747 17704 19756 17744
rect 19796 17704 19805 17744
rect 19747 17703 19805 17704
rect 13995 17660 14037 17669
rect 13995 17620 13996 17660
rect 14036 17620 14037 17660
rect 13995 17611 14037 17620
rect 19371 17660 19413 17669
rect 19371 17620 19372 17660
rect 19412 17620 19413 17660
rect 19371 17611 19413 17620
rect 8907 17576 8949 17585
rect 8907 17536 8908 17576
rect 8948 17536 8949 17576
rect 8907 17527 8949 17536
rect 10923 17576 10965 17585
rect 10923 17536 10924 17576
rect 10964 17536 10965 17576
rect 10923 17527 10965 17536
rect 1152 17408 20452 17432
rect 1152 17368 4928 17408
rect 4968 17368 5010 17408
rect 5050 17368 5092 17408
rect 5132 17368 5174 17408
rect 5214 17368 5256 17408
rect 5296 17368 20048 17408
rect 20088 17368 20130 17408
rect 20170 17368 20212 17408
rect 20252 17368 20294 17408
rect 20334 17368 20376 17408
rect 20416 17368 20452 17408
rect 1152 17344 20452 17368
rect 2667 17240 2709 17249
rect 2667 17200 2668 17240
rect 2708 17200 2709 17240
rect 2667 17191 2709 17200
rect 5539 17240 5597 17241
rect 5539 17200 5548 17240
rect 5588 17200 5597 17240
rect 5539 17199 5597 17200
rect 7179 17240 7221 17249
rect 7179 17200 7180 17240
rect 7220 17200 7221 17240
rect 7179 17191 7221 17200
rect 8907 17240 8949 17249
rect 8907 17200 8908 17240
rect 8948 17200 8949 17240
rect 8907 17191 8949 17200
rect 11403 17240 11445 17249
rect 11403 17200 11404 17240
rect 11444 17200 11445 17240
rect 11403 17191 11445 17200
rect 13419 17240 13461 17249
rect 13419 17200 13420 17240
rect 13460 17200 13461 17240
rect 13419 17191 13461 17200
rect 15427 17240 15485 17241
rect 15427 17200 15436 17240
rect 15476 17200 15485 17240
rect 15427 17199 15485 17200
rect 19851 17240 19893 17249
rect 19851 17200 19852 17240
rect 19892 17200 19893 17240
rect 19851 17191 19893 17200
rect 13707 17156 13749 17165
rect 13707 17116 13708 17156
rect 13748 17116 13749 17156
rect 13707 17107 13749 17116
rect 17547 17156 17589 17165
rect 17547 17116 17548 17156
rect 17588 17116 17589 17156
rect 17547 17107 17589 17116
rect 1219 17072 1277 17073
rect 1219 17032 1228 17072
rect 1268 17032 1277 17072
rect 1219 17031 1277 17032
rect 2467 17072 2525 17073
rect 2467 17032 2476 17072
rect 2516 17032 2525 17072
rect 2467 17031 2525 17032
rect 3051 17072 3093 17081
rect 3051 17032 3052 17072
rect 3092 17032 3093 17072
rect 3051 17023 3093 17032
rect 3339 17072 3381 17081
rect 3339 17032 3340 17072
rect 3380 17032 3381 17072
rect 3339 17023 3381 17032
rect 3523 17072 3581 17073
rect 3523 17032 3532 17072
rect 3572 17032 3581 17072
rect 3523 17031 3581 17032
rect 4771 17072 4829 17073
rect 4771 17032 4780 17072
rect 4820 17032 4829 17072
rect 4771 17031 4829 17032
rect 5259 17072 5301 17081
rect 5259 17032 5260 17072
rect 5300 17032 5301 17072
rect 5259 17023 5301 17032
rect 5355 17072 5397 17081
rect 5355 17032 5356 17072
rect 5396 17032 5397 17072
rect 5355 17023 5397 17032
rect 5731 17072 5789 17073
rect 5731 17032 5740 17072
rect 5780 17032 5789 17072
rect 5731 17031 5789 17032
rect 6979 17072 7037 17073
rect 6979 17032 6988 17072
rect 7028 17032 7037 17072
rect 6979 17031 7037 17032
rect 8707 17072 8765 17073
rect 8707 17032 8716 17072
rect 8756 17032 8765 17072
rect 8707 17031 8765 17032
rect 9955 17072 10013 17073
rect 9955 17032 9964 17072
rect 10004 17032 10013 17072
rect 9955 17031 10013 17032
rect 11203 17072 11261 17073
rect 11203 17032 11212 17072
rect 11252 17032 11261 17072
rect 11203 17031 11261 17032
rect 11691 17072 11733 17081
rect 11691 17032 11692 17072
rect 11732 17032 11733 17072
rect 7459 17030 7517 17031
rect 7459 16990 7468 17030
rect 7508 16990 7517 17030
rect 11691 17023 11733 17032
rect 11787 17072 11829 17081
rect 11787 17032 11788 17072
rect 11828 17032 11829 17072
rect 11787 17023 11829 17032
rect 12739 17072 12797 17073
rect 12739 17032 12748 17072
rect 12788 17032 12797 17072
rect 13891 17072 13949 17073
rect 12739 17031 12797 17032
rect 13227 17058 13269 17067
rect 13227 17018 13228 17058
rect 13268 17018 13269 17058
rect 13891 17032 13900 17072
rect 13940 17032 13949 17072
rect 13891 17031 13949 17032
rect 15139 17072 15197 17073
rect 15139 17032 15148 17072
rect 15188 17032 15197 17072
rect 15139 17031 15197 17032
rect 15339 17072 15381 17081
rect 15339 17032 15340 17072
rect 15380 17032 15381 17072
rect 15339 17023 15381 17032
rect 15531 17072 15573 17081
rect 15531 17032 15532 17072
rect 15572 17032 15573 17072
rect 15531 17023 15573 17032
rect 15619 17072 15677 17073
rect 15619 17032 15628 17072
rect 15668 17032 15677 17072
rect 15619 17031 15677 17032
rect 15907 17072 15965 17073
rect 15907 17032 15916 17072
rect 15956 17032 15965 17072
rect 15907 17031 15965 17032
rect 17155 17072 17213 17073
rect 17155 17032 17164 17072
rect 17204 17032 17213 17072
rect 17155 17031 17213 17032
rect 17739 17072 17781 17081
rect 17739 17032 17740 17072
rect 17780 17032 17781 17072
rect 17635 17030 17693 17031
rect 13227 17009 13269 17018
rect 7459 16989 7517 16990
rect 12171 16988 12213 16997
rect 12171 16948 12172 16988
rect 12212 16948 12213 16988
rect 12171 16939 12213 16948
rect 12267 16988 12309 16997
rect 17635 16990 17644 17030
rect 17684 16990 17693 17030
rect 17739 17023 17781 17032
rect 17835 17072 17877 17081
rect 17835 17032 17836 17072
rect 17876 17032 17877 17072
rect 17835 17023 17877 17032
rect 19651 17072 19709 17073
rect 19651 17032 19660 17072
rect 19700 17032 19709 17072
rect 19651 17031 19709 17032
rect 18403 17030 18461 17031
rect 17635 16989 17693 16990
rect 18403 16990 18412 17030
rect 18452 16990 18461 17030
rect 18403 16989 18461 16990
rect 12267 16948 12268 16988
rect 12308 16948 12309 16988
rect 12267 16939 12309 16948
rect 18019 16988 18077 16989
rect 18019 16948 18028 16988
rect 18068 16948 18077 16988
rect 18019 16947 18077 16948
rect 20035 16988 20093 16989
rect 20035 16948 20044 16988
rect 20084 16948 20093 16988
rect 20035 16947 20093 16948
rect 20235 16904 20277 16913
rect 20235 16864 20236 16904
rect 20276 16864 20277 16904
rect 20235 16855 20277 16864
rect 3339 16820 3381 16829
rect 3339 16780 3340 16820
rect 3380 16780 3381 16820
rect 3339 16771 3381 16780
rect 4971 16820 5013 16829
rect 4971 16780 4972 16820
rect 5012 16780 5013 16820
rect 4971 16771 5013 16780
rect 17355 16820 17397 16829
rect 17355 16780 17356 16820
rect 17396 16780 17397 16820
rect 17355 16771 17397 16780
rect 18219 16820 18261 16829
rect 18219 16780 18220 16820
rect 18260 16780 18261 16820
rect 18219 16771 18261 16780
rect 1152 16652 20352 16676
rect 1152 16612 3688 16652
rect 3728 16612 3770 16652
rect 3810 16612 3852 16652
rect 3892 16612 3934 16652
rect 3974 16612 4016 16652
rect 4056 16612 18808 16652
rect 18848 16612 18890 16652
rect 18930 16612 18972 16652
rect 19012 16612 19054 16652
rect 19094 16612 19136 16652
rect 19176 16612 20352 16652
rect 1152 16588 20352 16612
rect 2859 16484 2901 16493
rect 2859 16444 2860 16484
rect 2900 16444 2901 16484
rect 2859 16435 2901 16444
rect 13323 16484 13365 16493
rect 13323 16444 13324 16484
rect 13364 16444 13365 16484
rect 13323 16435 13365 16444
rect 16867 16484 16925 16485
rect 16867 16444 16876 16484
rect 16916 16444 16925 16484
rect 16867 16443 16925 16444
rect 6699 16400 6741 16409
rect 6699 16360 6700 16400
rect 6740 16360 6741 16400
rect 6699 16351 6741 16360
rect 15915 16400 15957 16409
rect 15915 16360 15916 16400
rect 15956 16360 15957 16400
rect 15915 16351 15957 16360
rect 17059 16400 17117 16401
rect 17059 16360 17068 16400
rect 17108 16360 17117 16400
rect 17059 16359 17117 16360
rect 19659 16400 19701 16409
rect 19659 16360 19660 16400
rect 19700 16360 19701 16400
rect 19659 16351 19701 16360
rect 3819 16316 3861 16325
rect 3819 16276 3820 16316
rect 3860 16276 3861 16316
rect 3819 16267 3861 16276
rect 3915 16316 3957 16325
rect 3915 16276 3916 16316
rect 3956 16276 3957 16316
rect 3915 16267 3957 16276
rect 4875 16246 4917 16255
rect 1411 16232 1469 16233
rect 1411 16192 1420 16232
rect 1460 16192 1469 16232
rect 1411 16191 1469 16192
rect 2659 16232 2717 16233
rect 2659 16192 2668 16232
rect 2708 16192 2717 16232
rect 2659 16191 2717 16192
rect 3339 16232 3381 16241
rect 3339 16192 3340 16232
rect 3380 16192 3381 16232
rect 3339 16183 3381 16192
rect 3435 16232 3477 16241
rect 3435 16192 3436 16232
rect 3476 16192 3477 16232
rect 3435 16183 3477 16192
rect 4387 16232 4445 16233
rect 4387 16192 4396 16232
rect 4436 16192 4445 16232
rect 4875 16206 4876 16246
rect 4916 16206 4917 16246
rect 4875 16197 4917 16206
rect 5251 16232 5309 16233
rect 4387 16191 4445 16192
rect 5251 16192 5260 16232
rect 5300 16192 5309 16232
rect 5251 16191 5309 16192
rect 6499 16232 6557 16233
rect 6499 16192 6508 16232
rect 6548 16192 6557 16232
rect 6499 16191 6557 16192
rect 6883 16232 6941 16233
rect 6883 16192 6892 16232
rect 6932 16192 6941 16232
rect 6883 16191 6941 16192
rect 6979 16232 7037 16233
rect 6979 16192 6988 16232
rect 7028 16192 7037 16232
rect 6979 16191 7037 16192
rect 7179 16232 7221 16241
rect 7179 16192 7180 16232
rect 7220 16192 7221 16232
rect 7179 16183 7221 16192
rect 7275 16232 7317 16241
rect 7275 16192 7276 16232
rect 7316 16192 7317 16232
rect 7275 16183 7317 16192
rect 7368 16232 7426 16233
rect 7368 16192 7377 16232
rect 7417 16192 7426 16232
rect 7368 16191 7426 16192
rect 7843 16232 7901 16233
rect 7843 16192 7852 16232
rect 7892 16192 7901 16232
rect 7843 16191 7901 16192
rect 9091 16232 9149 16233
rect 9091 16192 9100 16232
rect 9140 16192 9149 16232
rect 9091 16191 9149 16192
rect 9475 16232 9533 16233
rect 9475 16192 9484 16232
rect 9524 16192 9533 16232
rect 9475 16191 9533 16192
rect 10723 16232 10781 16233
rect 10723 16192 10732 16232
rect 10772 16192 10781 16232
rect 10723 16191 10781 16192
rect 11875 16232 11933 16233
rect 11875 16192 11884 16232
rect 11924 16192 11933 16232
rect 11875 16191 11933 16192
rect 13123 16232 13181 16233
rect 13123 16192 13132 16232
rect 13172 16192 13181 16232
rect 13123 16191 13181 16192
rect 15427 16232 15485 16233
rect 15427 16192 15436 16232
rect 15476 16192 15485 16232
rect 15427 16191 15485 16192
rect 15531 16232 15573 16241
rect 15531 16192 15532 16232
rect 15572 16192 15573 16232
rect 15531 16183 15573 16192
rect 15723 16232 15765 16241
rect 15723 16192 15724 16232
rect 15764 16192 15765 16232
rect 15723 16183 15765 16192
rect 15915 16232 15957 16241
rect 15915 16192 15916 16232
rect 15956 16192 15957 16232
rect 15915 16183 15957 16192
rect 16203 16232 16245 16241
rect 16203 16192 16204 16232
rect 16244 16192 16245 16232
rect 16203 16183 16245 16192
rect 16491 16232 16533 16241
rect 16491 16192 16492 16232
rect 16532 16192 16533 16232
rect 16491 16183 16533 16192
rect 16587 16232 16629 16241
rect 16587 16192 16588 16232
rect 16628 16192 16629 16232
rect 16587 16183 16629 16192
rect 16683 16232 16725 16241
rect 16683 16192 16684 16232
rect 16724 16192 16725 16232
rect 16683 16183 16725 16192
rect 17451 16232 17493 16241
rect 17451 16192 17452 16232
rect 17492 16192 17493 16232
rect 17451 16183 17493 16192
rect 17731 16232 17789 16233
rect 17731 16192 17740 16232
rect 17780 16192 17789 16232
rect 17731 16191 17789 16192
rect 18211 16232 18269 16233
rect 18211 16192 18220 16232
rect 18260 16192 18269 16232
rect 18211 16191 18269 16192
rect 19459 16232 19517 16233
rect 19459 16192 19468 16232
rect 19508 16192 19517 16232
rect 19459 16191 19517 16192
rect 19947 16232 19989 16241
rect 19947 16192 19948 16232
rect 19988 16192 19989 16232
rect 19947 16183 19989 16192
rect 20043 16232 20085 16241
rect 20043 16192 20044 16232
rect 20084 16192 20085 16232
rect 20043 16183 20085 16192
rect 20139 16211 20181 16220
rect 20139 16171 20140 16211
rect 20180 16171 20181 16211
rect 20139 16162 20181 16171
rect 5067 16148 5109 16157
rect 5067 16108 5068 16148
rect 5108 16108 5109 16148
rect 5067 16099 5109 16108
rect 15627 16148 15669 16157
rect 15627 16108 15628 16148
rect 15668 16108 15669 16148
rect 15627 16099 15669 16108
rect 17355 16148 17397 16157
rect 17355 16108 17356 16148
rect 17396 16108 17397 16148
rect 17355 16099 17397 16108
rect 2859 16064 2901 16073
rect 2859 16024 2860 16064
rect 2900 16024 2901 16064
rect 2859 16015 2901 16024
rect 7075 16064 7133 16065
rect 7075 16024 7084 16064
rect 7124 16024 7133 16064
rect 7075 16023 7133 16024
rect 9291 16064 9333 16073
rect 9291 16024 9292 16064
rect 9332 16024 9333 16064
rect 9291 16015 9333 16024
rect 10923 16064 10965 16073
rect 10923 16024 10924 16064
rect 10964 16024 10965 16064
rect 10923 16015 10965 16024
rect 19843 16064 19901 16065
rect 19843 16024 19852 16064
rect 19892 16024 19901 16064
rect 19843 16023 19901 16024
rect 1152 15896 20452 15920
rect 1152 15856 4928 15896
rect 4968 15856 5010 15896
rect 5050 15856 5092 15896
rect 5132 15856 5174 15896
rect 5214 15856 5256 15896
rect 5296 15856 20048 15896
rect 20088 15856 20130 15896
rect 20170 15856 20212 15896
rect 20252 15856 20294 15896
rect 20334 15856 20376 15896
rect 20416 15856 20452 15896
rect 1152 15832 20452 15856
rect 2667 15728 2709 15737
rect 2667 15688 2668 15728
rect 2708 15688 2709 15728
rect 2667 15679 2709 15688
rect 4203 15728 4245 15737
rect 4203 15688 4204 15728
rect 4244 15688 4245 15728
rect 4203 15679 4245 15688
rect 4587 15728 4629 15737
rect 4587 15688 4588 15728
rect 4628 15688 4629 15728
rect 4587 15679 4629 15688
rect 12555 15728 12597 15737
rect 12555 15688 12556 15728
rect 12596 15688 12597 15728
rect 12555 15679 12597 15688
rect 15915 15728 15957 15737
rect 15915 15688 15916 15728
rect 15956 15688 15957 15728
rect 15915 15679 15957 15688
rect 17931 15728 17973 15737
rect 17931 15688 17932 15728
rect 17972 15688 17973 15728
rect 17931 15679 17973 15688
rect 20235 15728 20277 15737
rect 20235 15688 20236 15728
rect 20276 15688 20277 15728
rect 20235 15679 20277 15688
rect 9675 15644 9717 15653
rect 9675 15604 9676 15644
rect 9716 15604 9717 15644
rect 9675 15595 9717 15604
rect 1219 15560 1277 15561
rect 1219 15520 1228 15560
rect 1268 15520 1277 15560
rect 1219 15519 1277 15520
rect 2467 15560 2525 15561
rect 2467 15520 2476 15560
rect 2516 15520 2525 15560
rect 2467 15519 2525 15520
rect 3051 15560 3093 15569
rect 3051 15520 3052 15560
rect 3092 15520 3093 15560
rect 3051 15511 3093 15520
rect 3147 15560 3189 15569
rect 3147 15520 3148 15560
rect 3188 15520 3189 15560
rect 3147 15511 3189 15520
rect 3243 15560 3285 15569
rect 3243 15520 3244 15560
rect 3284 15520 3285 15560
rect 3243 15511 3285 15520
rect 3627 15560 3669 15569
rect 3627 15520 3628 15560
rect 3668 15520 3669 15560
rect 3627 15511 3669 15520
rect 3819 15560 3861 15569
rect 3819 15520 3820 15560
rect 3860 15520 3861 15560
rect 3819 15511 3861 15520
rect 3907 15560 3965 15561
rect 3907 15520 3916 15560
rect 3956 15520 3965 15560
rect 3907 15519 3965 15520
rect 4107 15560 4149 15569
rect 4107 15520 4108 15560
rect 4148 15520 4149 15560
rect 4107 15511 4149 15520
rect 4299 15560 4341 15569
rect 4299 15520 4300 15560
rect 4340 15520 4341 15560
rect 4299 15511 4341 15520
rect 4395 15560 4437 15569
rect 4395 15520 4396 15560
rect 4436 15520 4437 15560
rect 4395 15511 4437 15520
rect 4771 15560 4829 15561
rect 4771 15520 4780 15560
rect 4820 15520 4829 15560
rect 4771 15519 4829 15520
rect 6019 15560 6077 15561
rect 6019 15520 6028 15560
rect 6068 15520 6077 15560
rect 6019 15519 6077 15520
rect 6211 15560 6269 15561
rect 6211 15520 6220 15560
rect 6260 15520 6269 15560
rect 6211 15519 6269 15520
rect 7459 15560 7517 15561
rect 7459 15520 7468 15560
rect 7508 15520 7517 15560
rect 7459 15519 7517 15520
rect 7947 15560 7989 15569
rect 7947 15520 7948 15560
rect 7988 15520 7989 15560
rect 7947 15511 7989 15520
rect 8043 15560 8085 15569
rect 8043 15520 8044 15560
rect 8084 15520 8085 15560
rect 8043 15511 8085 15520
rect 8427 15560 8469 15569
rect 8427 15520 8428 15560
rect 8468 15520 8469 15560
rect 8427 15511 8469 15520
rect 8523 15560 8565 15569
rect 8523 15520 8524 15560
rect 8564 15520 8565 15560
rect 8523 15511 8565 15520
rect 8995 15560 9053 15561
rect 8995 15520 9004 15560
rect 9044 15520 9053 15560
rect 8995 15519 9053 15520
rect 9483 15555 9525 15564
rect 9483 15515 9484 15555
rect 9524 15515 9525 15555
rect 9483 15506 9525 15515
rect 10827 15560 10869 15569
rect 10827 15520 10828 15560
rect 10868 15520 10869 15560
rect 10827 15511 10869 15520
rect 10923 15560 10965 15569
rect 10923 15520 10924 15560
rect 10964 15520 10965 15560
rect 10923 15511 10965 15520
rect 11403 15560 11445 15569
rect 11403 15520 11404 15560
rect 11444 15520 11445 15560
rect 11403 15511 11445 15520
rect 11875 15560 11933 15561
rect 11875 15520 11884 15560
rect 11924 15520 11933 15560
rect 12739 15560 12797 15561
rect 11875 15519 11933 15520
rect 12363 15546 12405 15555
rect 12363 15506 12364 15546
rect 12404 15506 12405 15546
rect 12739 15520 12748 15560
rect 12788 15520 12797 15560
rect 12739 15519 12797 15520
rect 13987 15560 14045 15561
rect 13987 15520 13996 15560
rect 14036 15520 14045 15560
rect 13987 15519 14045 15520
rect 14467 15560 14525 15561
rect 14467 15520 14476 15560
rect 14516 15520 14525 15560
rect 14467 15519 14525 15520
rect 15715 15560 15773 15561
rect 15715 15520 15724 15560
rect 15764 15520 15773 15560
rect 15715 15519 15773 15520
rect 16203 15560 16245 15569
rect 16203 15520 16204 15560
rect 16244 15520 16245 15560
rect 16203 15511 16245 15520
rect 16299 15560 16341 15569
rect 16299 15520 16300 15560
rect 16340 15520 16341 15560
rect 16299 15511 16341 15520
rect 16779 15560 16821 15569
rect 16779 15520 16780 15560
rect 16820 15520 16821 15560
rect 16779 15511 16821 15520
rect 17251 15560 17309 15561
rect 17251 15520 17260 15560
rect 17300 15520 17309 15560
rect 18507 15560 18549 15569
rect 17251 15519 17309 15520
rect 17787 15550 17829 15559
rect 12363 15497 12405 15506
rect 17787 15510 17788 15550
rect 17828 15510 17829 15550
rect 18507 15520 18508 15560
rect 18548 15520 18549 15560
rect 18507 15511 18549 15520
rect 18603 15560 18645 15569
rect 18603 15520 18604 15560
rect 18644 15520 18645 15560
rect 18603 15511 18645 15520
rect 18987 15560 19029 15569
rect 18987 15520 18988 15560
rect 19028 15520 19029 15560
rect 18987 15511 19029 15520
rect 19555 15560 19613 15561
rect 19555 15520 19564 15560
rect 19604 15520 19613 15560
rect 19555 15519 19613 15520
rect 20043 15546 20085 15555
rect 17787 15501 17829 15510
rect 20043 15506 20044 15546
rect 20084 15506 20085 15546
rect 20043 15497 20085 15506
rect 11307 15476 11349 15485
rect 11307 15436 11308 15476
rect 11348 15436 11349 15476
rect 11307 15427 11349 15436
rect 16683 15476 16725 15485
rect 16683 15436 16684 15476
rect 16724 15436 16725 15476
rect 16683 15427 16725 15436
rect 19083 15476 19125 15485
rect 19083 15436 19084 15476
rect 19124 15436 19125 15476
rect 19083 15427 19125 15436
rect 3427 15308 3485 15309
rect 3427 15268 3436 15308
rect 3476 15268 3485 15308
rect 3427 15267 3485 15268
rect 3627 15308 3669 15317
rect 3627 15268 3628 15308
rect 3668 15268 3669 15308
rect 3627 15259 3669 15268
rect 7659 15308 7701 15317
rect 7659 15268 7660 15308
rect 7700 15268 7701 15308
rect 7659 15259 7701 15268
rect 14187 15308 14229 15317
rect 14187 15268 14188 15308
rect 14228 15268 14229 15308
rect 14187 15259 14229 15268
rect 1152 15140 20352 15164
rect 1152 15100 3688 15140
rect 3728 15100 3770 15140
rect 3810 15100 3852 15140
rect 3892 15100 3934 15140
rect 3974 15100 4016 15140
rect 4056 15100 18808 15140
rect 18848 15100 18890 15140
rect 18930 15100 18972 15140
rect 19012 15100 19054 15140
rect 19094 15100 19136 15140
rect 19176 15100 20352 15140
rect 1152 15076 20352 15100
rect 2851 14972 2909 14973
rect 2851 14932 2860 14972
rect 2900 14932 2909 14972
rect 2851 14931 2909 14932
rect 7659 14972 7701 14981
rect 7659 14932 7660 14972
rect 7700 14932 7701 14972
rect 7659 14923 7701 14932
rect 12171 14972 12213 14981
rect 12171 14932 12172 14972
rect 12212 14932 12213 14972
rect 12171 14923 12213 14932
rect 13795 14972 13853 14973
rect 13795 14932 13804 14972
rect 13844 14932 13853 14972
rect 13795 14931 13853 14932
rect 16779 14972 16821 14981
rect 16779 14932 16780 14972
rect 16820 14932 16821 14972
rect 16779 14923 16821 14932
rect 19083 14972 19125 14981
rect 19083 14932 19084 14972
rect 19124 14932 19125 14972
rect 19083 14923 19125 14932
rect 19747 14972 19805 14973
rect 19747 14932 19756 14972
rect 19796 14932 19805 14972
rect 19747 14931 19805 14932
rect 19947 14972 19989 14981
rect 19947 14932 19948 14972
rect 19988 14932 19989 14972
rect 19947 14923 19989 14932
rect 12939 14888 12981 14897
rect 12939 14848 12940 14888
rect 12980 14848 12981 14888
rect 12939 14839 12981 14848
rect 8619 14804 8661 14813
rect 8619 14764 8620 14804
rect 8660 14764 8661 14804
rect 8619 14755 8661 14764
rect 9579 14734 9621 14743
rect 1219 14720 1277 14721
rect 1219 14680 1228 14720
rect 1268 14680 1277 14720
rect 1219 14679 1277 14680
rect 2467 14720 2525 14721
rect 2467 14680 2476 14720
rect 2516 14680 2525 14720
rect 2467 14679 2525 14680
rect 3243 14720 3285 14729
rect 3243 14680 3244 14720
rect 3284 14680 3285 14720
rect 3243 14671 3285 14680
rect 3523 14720 3581 14721
rect 3523 14680 3532 14720
rect 3572 14680 3581 14720
rect 3523 14679 3581 14680
rect 3915 14720 3957 14729
rect 3915 14680 3916 14720
rect 3956 14680 3957 14720
rect 3915 14671 3957 14680
rect 4011 14720 4053 14729
rect 4011 14680 4012 14720
rect 4052 14680 4053 14720
rect 4011 14671 4053 14680
rect 4107 14720 4149 14729
rect 4107 14680 4108 14720
rect 4148 14680 4149 14720
rect 4107 14671 4149 14680
rect 4387 14720 4445 14721
rect 4387 14680 4396 14720
rect 4436 14680 4445 14720
rect 4387 14679 4445 14680
rect 5635 14720 5693 14721
rect 5635 14680 5644 14720
rect 5684 14680 5693 14720
rect 5635 14679 5693 14680
rect 6211 14720 6269 14721
rect 6211 14680 6220 14720
rect 6260 14680 6269 14720
rect 6211 14679 6269 14680
rect 7459 14720 7517 14721
rect 7459 14680 7468 14720
rect 7508 14680 7517 14720
rect 7459 14679 7517 14680
rect 8043 14720 8085 14729
rect 8043 14680 8044 14720
rect 8084 14680 8085 14720
rect 8043 14671 8085 14680
rect 8139 14720 8181 14729
rect 8139 14680 8140 14720
rect 8180 14680 8181 14720
rect 8139 14671 8181 14680
rect 8523 14720 8565 14729
rect 8523 14680 8524 14720
rect 8564 14680 8565 14720
rect 8523 14671 8565 14680
rect 9091 14720 9149 14721
rect 9091 14680 9100 14720
rect 9140 14680 9149 14720
rect 9579 14694 9580 14734
rect 9620 14694 9621 14734
rect 20131 14734 20189 14735
rect 9579 14685 9621 14694
rect 10723 14720 10781 14721
rect 9091 14679 9149 14680
rect 10723 14680 10732 14720
rect 10772 14680 10781 14720
rect 10723 14679 10781 14680
rect 11971 14720 12029 14721
rect 11971 14680 11980 14720
rect 12020 14680 12029 14720
rect 11971 14679 12029 14680
rect 12643 14720 12701 14721
rect 12643 14680 12652 14720
rect 12692 14680 12701 14720
rect 12643 14679 12701 14680
rect 12747 14720 12789 14729
rect 12747 14680 12748 14720
rect 12788 14680 12789 14720
rect 12747 14671 12789 14680
rect 12939 14720 12981 14729
rect 12939 14680 12940 14720
rect 12980 14680 12981 14720
rect 12939 14671 12981 14680
rect 13227 14720 13269 14729
rect 13227 14680 13228 14720
rect 13268 14680 13269 14720
rect 13227 14671 13269 14680
rect 13323 14720 13365 14729
rect 13323 14680 13324 14720
rect 13364 14680 13365 14720
rect 13323 14671 13365 14680
rect 13419 14720 13461 14729
rect 13419 14680 13420 14720
rect 13460 14680 13461 14720
rect 13419 14671 13461 14680
rect 14187 14720 14229 14729
rect 14187 14680 14188 14720
rect 14228 14680 14229 14720
rect 14187 14671 14229 14680
rect 14467 14720 14525 14721
rect 14467 14680 14476 14720
rect 14516 14680 14525 14720
rect 14467 14679 14525 14680
rect 14763 14720 14805 14729
rect 14763 14680 14764 14720
rect 14804 14680 14805 14720
rect 14763 14671 14805 14680
rect 14859 14720 14901 14729
rect 14859 14680 14860 14720
rect 14900 14680 14901 14720
rect 14859 14671 14901 14680
rect 14955 14720 14997 14729
rect 14955 14680 14956 14720
rect 14996 14680 14997 14720
rect 14955 14671 14997 14680
rect 15051 14720 15093 14729
rect 15051 14680 15052 14720
rect 15092 14680 15093 14720
rect 15051 14671 15093 14680
rect 15331 14720 15389 14721
rect 15331 14680 15340 14720
rect 15380 14680 15389 14720
rect 15331 14679 15389 14680
rect 16579 14720 16637 14721
rect 16579 14680 16588 14720
rect 16628 14680 16637 14720
rect 16579 14679 16637 14680
rect 17635 14720 17693 14721
rect 17635 14680 17644 14720
rect 17684 14680 17693 14720
rect 17635 14679 17693 14680
rect 18883 14720 18941 14721
rect 18883 14680 18892 14720
rect 18932 14680 18941 14720
rect 18883 14679 18941 14680
rect 19371 14720 19413 14729
rect 19371 14680 19372 14720
rect 19412 14680 19413 14720
rect 19371 14671 19413 14680
rect 19467 14720 19509 14729
rect 19467 14680 19468 14720
rect 19508 14680 19509 14720
rect 19467 14671 19509 14680
rect 19563 14720 19605 14729
rect 19563 14680 19564 14720
rect 19604 14680 19605 14720
rect 19563 14671 19605 14680
rect 19947 14720 19989 14729
rect 19947 14680 19948 14720
rect 19988 14680 19989 14720
rect 20131 14694 20140 14734
rect 20180 14694 20189 14734
rect 20131 14693 20189 14694
rect 20227 14720 20285 14721
rect 19947 14671 19989 14680
rect 20227 14680 20236 14720
rect 20276 14680 20285 14720
rect 20227 14679 20285 14680
rect 3147 14636 3189 14645
rect 3147 14596 3148 14636
rect 3188 14596 3189 14636
rect 3147 14587 3189 14596
rect 3819 14636 3861 14645
rect 3819 14596 3820 14636
rect 3860 14596 3861 14636
rect 3819 14587 3861 14596
rect 14091 14636 14133 14645
rect 14091 14596 14092 14636
rect 14132 14596 14133 14636
rect 14091 14587 14133 14596
rect 2667 14552 2709 14561
rect 2667 14512 2668 14552
rect 2708 14512 2709 14552
rect 2667 14503 2709 14512
rect 5835 14552 5877 14561
rect 5835 14512 5836 14552
rect 5876 14512 5877 14552
rect 5835 14503 5877 14512
rect 9771 14552 9813 14561
rect 9771 14512 9772 14552
rect 9812 14512 9813 14552
rect 9771 14503 9813 14512
rect 13611 14552 13653 14561
rect 13611 14512 13612 14552
rect 13652 14512 13653 14552
rect 13611 14503 13653 14512
rect 1152 14384 20452 14408
rect 1152 14344 4928 14384
rect 4968 14344 5010 14384
rect 5050 14344 5092 14384
rect 5132 14344 5174 14384
rect 5214 14344 5256 14384
rect 5296 14344 20048 14384
rect 20088 14344 20130 14384
rect 20170 14344 20212 14384
rect 20252 14344 20294 14384
rect 20334 14344 20376 14384
rect 20416 14344 20452 14384
rect 1152 14320 20452 14344
rect 2667 14216 2709 14225
rect 2667 14176 2668 14216
rect 2708 14176 2709 14216
rect 2667 14167 2709 14176
rect 12459 14216 12501 14225
rect 12459 14176 12460 14216
rect 12500 14176 12501 14216
rect 12459 14167 12501 14176
rect 14283 14216 14325 14225
rect 14283 14176 14284 14216
rect 14324 14176 14325 14216
rect 14283 14167 14325 14176
rect 18411 14216 18453 14225
rect 18411 14176 18412 14216
rect 18452 14176 18453 14216
rect 18411 14167 18453 14176
rect 7659 14132 7701 14141
rect 7659 14092 7660 14132
rect 7700 14092 7701 14132
rect 7659 14083 7701 14092
rect 9195 14132 9237 14141
rect 9195 14092 9196 14132
rect 9236 14092 9237 14132
rect 9195 14083 9237 14092
rect 20139 14132 20181 14141
rect 20139 14092 20140 14132
rect 20180 14092 20181 14132
rect 20139 14083 20181 14092
rect 16683 14069 16725 14078
rect 2859 14043 2901 14052
rect 2859 14003 2860 14043
rect 2900 14003 2901 14043
rect 3331 14048 3389 14049
rect 3331 14008 3340 14048
rect 3380 14008 3389 14048
rect 3331 14007 3389 14008
rect 3915 14048 3957 14057
rect 3915 14008 3916 14048
rect 3956 14008 3957 14048
rect 2859 13994 2901 14003
rect 3915 13999 3957 14008
rect 4299 14048 4341 14057
rect 4299 14008 4300 14048
rect 4340 14008 4341 14048
rect 4299 13999 4341 14008
rect 4395 14048 4437 14057
rect 4395 14008 4396 14048
rect 4436 14008 4437 14048
rect 4395 13999 4437 14008
rect 5931 14048 5973 14057
rect 5931 14008 5932 14048
rect 5972 14008 5973 14048
rect 5931 13999 5973 14008
rect 6027 14048 6069 14057
rect 6027 14008 6028 14048
rect 6068 14008 6069 14048
rect 6027 13999 6069 14008
rect 6411 14048 6453 14057
rect 6411 14008 6412 14048
rect 6452 14008 6453 14048
rect 6411 13999 6453 14008
rect 6507 14048 6549 14057
rect 6507 14008 6508 14048
rect 6548 14008 6549 14048
rect 6507 13999 6549 14008
rect 6979 14048 7037 14049
rect 6979 14008 6988 14048
rect 7028 14008 7037 14048
rect 8419 14048 8477 14049
rect 6979 14007 7037 14008
rect 7467 14034 7509 14043
rect 7467 13994 7468 14034
rect 7508 13994 7509 14034
rect 8419 14008 8428 14048
rect 8468 14008 8477 14048
rect 8419 14007 8477 14008
rect 8523 14048 8565 14057
rect 8523 14008 8524 14048
rect 8564 14008 8565 14048
rect 8523 13999 8565 14008
rect 8715 14048 8757 14057
rect 8715 14008 8716 14048
rect 8756 14008 8757 14048
rect 8715 13999 8757 14008
rect 9291 14048 9333 14057
rect 9291 14008 9292 14048
rect 9332 14008 9333 14048
rect 9291 13999 9333 14008
rect 9571 14048 9629 14049
rect 9571 14008 9580 14048
rect 9620 14008 9629 14048
rect 9571 14007 9629 14008
rect 11011 14048 11069 14049
rect 11011 14008 11020 14048
rect 11060 14008 11069 14048
rect 11011 14007 11069 14008
rect 12259 14048 12317 14049
rect 12259 14008 12268 14048
rect 12308 14008 12317 14048
rect 12259 14007 12317 14008
rect 12835 14048 12893 14049
rect 12835 14008 12844 14048
rect 12884 14008 12893 14048
rect 12835 14007 12893 14008
rect 14083 14048 14141 14049
rect 14083 14008 14092 14048
rect 14132 14008 14141 14048
rect 14083 14007 14141 14008
rect 14475 14048 14517 14057
rect 14475 14008 14476 14048
rect 14516 14008 14517 14048
rect 14475 13999 14517 14008
rect 14763 14048 14805 14057
rect 14763 14008 14764 14048
rect 14804 14008 14805 14048
rect 14763 13999 14805 14008
rect 14947 14048 15005 14049
rect 14947 14008 14956 14048
rect 14996 14008 15005 14048
rect 14947 14007 15005 14008
rect 16195 14048 16253 14049
rect 16195 14008 16204 14048
rect 16244 14008 16253 14048
rect 16195 14007 16253 14008
rect 16587 14048 16629 14057
rect 16587 14008 16588 14048
rect 16628 14008 16629 14048
rect 16683 14029 16684 14069
rect 16724 14029 16725 14069
rect 16683 14020 16725 14029
rect 16779 14048 16821 14057
rect 16587 13999 16629 14008
rect 16779 14008 16780 14048
rect 16820 14008 16821 14048
rect 16779 13999 16821 14008
rect 16875 14048 16917 14057
rect 16875 14008 16876 14048
rect 16916 14008 16917 14048
rect 16875 13999 16917 14008
rect 17067 14048 17109 14057
rect 17067 14008 17068 14048
rect 17108 14008 17109 14048
rect 17067 13999 17109 14008
rect 17259 14048 17301 14057
rect 17259 14008 17260 14048
rect 17300 14008 17301 14048
rect 17259 13999 17301 14008
rect 17347 14048 17405 14049
rect 17347 14008 17356 14048
rect 17396 14008 17405 14048
rect 17347 14007 17405 14008
rect 18219 14048 18261 14057
rect 18219 14008 18220 14048
rect 18260 14008 18261 14048
rect 18219 13999 18261 14008
rect 18507 14048 18549 14057
rect 18507 14008 18508 14048
rect 18548 14008 18549 14048
rect 18507 13999 18549 14008
rect 18691 14048 18749 14049
rect 18691 14008 18700 14048
rect 18740 14008 18749 14048
rect 18691 14007 18749 14008
rect 19939 14048 19997 14049
rect 19939 14008 19948 14048
rect 19988 14008 19997 14048
rect 19939 14007 19997 14008
rect 7467 13985 7509 13994
rect 3819 13964 3861 13973
rect 3819 13924 3820 13964
rect 3860 13924 3861 13964
rect 3819 13915 3861 13924
rect 8899 13880 8957 13881
rect 8899 13840 8908 13880
rect 8948 13840 8957 13880
rect 8899 13839 8957 13840
rect 16395 13880 16437 13889
rect 16395 13840 16396 13880
rect 16436 13840 16437 13880
rect 16395 13831 16437 13840
rect 17067 13880 17109 13889
rect 17067 13840 17068 13880
rect 17108 13840 17109 13880
rect 17067 13831 17109 13840
rect 8715 13796 8757 13805
rect 8715 13756 8716 13796
rect 8756 13756 8757 13796
rect 8715 13747 8757 13756
rect 14283 13796 14325 13805
rect 14283 13756 14284 13796
rect 14324 13756 14325 13796
rect 14283 13747 14325 13756
rect 14475 13796 14517 13805
rect 14475 13756 14476 13796
rect 14516 13756 14517 13796
rect 14475 13747 14517 13756
rect 1152 13628 20352 13652
rect 1152 13588 3688 13628
rect 3728 13588 3770 13628
rect 3810 13588 3852 13628
rect 3892 13588 3934 13628
rect 3974 13588 4016 13628
rect 4056 13588 18808 13628
rect 18848 13588 18890 13628
rect 18930 13588 18972 13628
rect 19012 13588 19054 13628
rect 19094 13588 19136 13628
rect 19176 13588 20352 13628
rect 1152 13564 20352 13588
rect 7083 13460 7125 13469
rect 7083 13420 7084 13460
rect 7124 13420 7125 13460
rect 7083 13411 7125 13420
rect 8715 13460 8757 13469
rect 8715 13420 8716 13460
rect 8756 13420 8757 13460
rect 8715 13411 8757 13420
rect 14667 13460 14709 13469
rect 14667 13420 14668 13460
rect 14708 13420 14709 13460
rect 14667 13411 14709 13420
rect 16971 13376 17013 13385
rect 16971 13336 16972 13376
rect 17012 13336 17013 13376
rect 16971 13327 17013 13336
rect 11211 13292 11253 13301
rect 11211 13252 11212 13292
rect 11252 13252 11253 13292
rect 11211 13243 11253 13252
rect 15627 13292 15669 13301
rect 15627 13252 15628 13292
rect 15668 13252 15669 13292
rect 15627 13243 15669 13252
rect 17347 13251 17405 13252
rect 2763 13213 2805 13222
rect 12171 13217 12213 13226
rect 14187 13222 14229 13231
rect 2763 13173 2764 13213
rect 2804 13173 2805 13213
rect 2763 13164 2805 13173
rect 3235 13208 3293 13209
rect 3235 13168 3244 13208
rect 3284 13168 3293 13208
rect 3235 13167 3293 13168
rect 3723 13208 3765 13217
rect 3723 13168 3724 13208
rect 3764 13168 3765 13208
rect 3723 13159 3765 13168
rect 3819 13208 3861 13217
rect 3819 13168 3820 13208
rect 3860 13168 3861 13208
rect 3819 13159 3861 13168
rect 4203 13208 4245 13217
rect 4203 13168 4204 13208
rect 4244 13168 4245 13208
rect 4203 13159 4245 13168
rect 4299 13208 4341 13217
rect 4299 13168 4300 13208
rect 4340 13168 4341 13208
rect 4299 13159 4341 13168
rect 5635 13208 5693 13209
rect 5635 13168 5644 13208
rect 5684 13168 5693 13208
rect 5635 13167 5693 13168
rect 6883 13208 6941 13209
rect 6883 13168 6892 13208
rect 6932 13168 6941 13208
rect 6883 13167 6941 13168
rect 7267 13208 7325 13209
rect 7267 13168 7276 13208
rect 7316 13168 7325 13208
rect 7267 13167 7325 13168
rect 8515 13208 8573 13209
rect 8515 13168 8524 13208
rect 8564 13168 8573 13208
rect 8515 13167 8573 13168
rect 8899 13208 8957 13209
rect 8899 13168 8908 13208
rect 8948 13168 8957 13208
rect 8899 13167 8957 13168
rect 10147 13208 10205 13209
rect 10147 13168 10156 13208
rect 10196 13168 10205 13208
rect 10147 13167 10205 13168
rect 10635 13208 10677 13217
rect 10635 13168 10636 13208
rect 10676 13168 10677 13208
rect 10635 13159 10677 13168
rect 10731 13208 10773 13217
rect 10731 13168 10732 13208
rect 10772 13168 10773 13208
rect 10731 13159 10773 13168
rect 11115 13208 11157 13217
rect 11115 13168 11116 13208
rect 11156 13168 11157 13208
rect 11115 13159 11157 13168
rect 11683 13207 11741 13208
rect 11683 13167 11692 13207
rect 11732 13167 11741 13207
rect 12171 13177 12172 13217
rect 12212 13177 12213 13217
rect 12171 13168 12213 13177
rect 12651 13208 12693 13217
rect 12651 13168 12652 13208
rect 12692 13168 12693 13208
rect 11683 13166 11741 13167
rect 12651 13159 12693 13168
rect 12747 13208 12789 13217
rect 12747 13168 12748 13208
rect 12788 13168 12789 13208
rect 12747 13159 12789 13168
rect 13131 13208 13173 13217
rect 13131 13168 13132 13208
rect 13172 13168 13173 13208
rect 13131 13159 13173 13168
rect 13227 13208 13269 13217
rect 13227 13168 13228 13208
rect 13268 13168 13269 13208
rect 13227 13159 13269 13168
rect 13699 13208 13757 13209
rect 13699 13168 13708 13208
rect 13748 13168 13757 13208
rect 14187 13182 14188 13222
rect 14228 13182 14229 13222
rect 14187 13173 14229 13182
rect 14755 13208 14813 13209
rect 13699 13167 13757 13168
rect 14755 13168 14764 13208
rect 14804 13168 14813 13208
rect 14755 13167 14813 13168
rect 15051 13208 15093 13217
rect 15051 13168 15052 13208
rect 15092 13168 15093 13208
rect 15051 13159 15093 13168
rect 15147 13208 15189 13217
rect 15147 13168 15148 13208
rect 15188 13168 15189 13208
rect 15147 13159 15189 13168
rect 15531 13208 15573 13217
rect 16587 13213 16629 13222
rect 15531 13168 15532 13208
rect 15572 13168 15573 13208
rect 15531 13159 15573 13168
rect 16099 13208 16157 13209
rect 16099 13168 16108 13208
rect 16148 13168 16157 13208
rect 16099 13167 16157 13168
rect 16587 13173 16588 13213
rect 16628 13173 16629 13213
rect 16587 13164 16629 13173
rect 17259 13208 17301 13217
rect 17347 13211 17356 13251
rect 17396 13211 17405 13251
rect 17347 13210 17405 13211
rect 17259 13168 17260 13208
rect 17300 13168 17301 13208
rect 17259 13159 17301 13168
rect 17827 13208 17885 13209
rect 17827 13168 17836 13208
rect 17876 13168 17885 13208
rect 17827 13167 17885 13168
rect 19075 13208 19133 13209
rect 19075 13168 19084 13208
rect 19124 13168 19133 13208
rect 19075 13167 19133 13168
rect 19563 13208 19605 13217
rect 19563 13168 19564 13208
rect 19604 13168 19605 13208
rect 19563 13159 19605 13168
rect 19659 13208 19701 13217
rect 19659 13168 19660 13208
rect 19700 13168 19701 13208
rect 19659 13159 19701 13168
rect 19755 13208 19797 13217
rect 19755 13168 19756 13208
rect 19796 13168 19797 13208
rect 19755 13159 19797 13168
rect 2571 13124 2613 13133
rect 2571 13084 2572 13124
rect 2612 13084 2613 13124
rect 2571 13075 2613 13084
rect 10347 13124 10389 13133
rect 10347 13084 10348 13124
rect 10388 13084 10389 13124
rect 10347 13075 10389 13084
rect 12363 13124 12405 13133
rect 12363 13084 12364 13124
rect 12404 13084 12405 13124
rect 12363 13075 12405 13084
rect 14379 13124 14421 13133
rect 14379 13084 14380 13124
rect 14420 13084 14421 13124
rect 14379 13075 14421 13084
rect 16779 13082 16821 13091
rect 8715 13040 8757 13049
rect 8715 13000 8716 13040
rect 8756 13000 8757 13040
rect 16779 13042 16780 13082
rect 16820 13042 16821 13082
rect 16779 13033 16821 13042
rect 19275 13040 19317 13049
rect 8715 12991 8757 13000
rect 19275 13000 19276 13040
rect 19316 13000 19317 13040
rect 19275 12991 19317 13000
rect 19459 13040 19517 13041
rect 19459 13000 19468 13040
rect 19508 13000 19517 13040
rect 19459 12999 19517 13000
rect 17451 12982 17493 12991
rect 17451 12942 17452 12982
rect 17492 12942 17493 12982
rect 17451 12933 17493 12942
rect 1152 12872 20452 12896
rect 1152 12832 4928 12872
rect 4968 12832 5010 12872
rect 5050 12832 5092 12872
rect 5132 12832 5174 12872
rect 5214 12832 5256 12872
rect 5296 12832 20048 12872
rect 20088 12832 20130 12872
rect 20170 12832 20212 12872
rect 20252 12832 20294 12872
rect 20334 12832 20376 12872
rect 20416 12832 20452 12872
rect 1152 12808 20452 12832
rect 12267 12704 12309 12713
rect 12267 12664 12268 12704
rect 12308 12664 12309 12704
rect 12267 12655 12309 12664
rect 19851 12704 19893 12713
rect 19851 12664 19852 12704
rect 19892 12664 19893 12704
rect 19851 12655 19893 12664
rect 2283 12620 2325 12629
rect 2283 12580 2284 12620
rect 2324 12580 2325 12620
rect 2283 12571 2325 12580
rect 7371 12620 7413 12629
rect 7371 12580 7372 12620
rect 7412 12580 7413 12620
rect 7371 12571 7413 12580
rect 15243 12620 15285 12629
rect 15243 12580 15244 12620
rect 15284 12580 15285 12620
rect 15243 12571 15285 12580
rect 15531 12620 15573 12629
rect 15531 12580 15532 12620
rect 15572 12580 15573 12620
rect 15531 12571 15573 12580
rect 17643 12620 17685 12629
rect 17643 12580 17644 12620
rect 17684 12580 17685 12620
rect 17643 12571 17685 12580
rect 2467 12536 2525 12537
rect 2467 12496 2476 12536
rect 2516 12496 2525 12536
rect 2467 12495 2525 12496
rect 3715 12536 3773 12537
rect 3715 12496 3724 12536
rect 3764 12496 3773 12536
rect 3715 12495 3773 12496
rect 3907 12536 3965 12537
rect 3907 12496 3916 12536
rect 3956 12496 3965 12536
rect 3907 12495 3965 12496
rect 5155 12536 5213 12537
rect 5155 12496 5164 12536
rect 5204 12496 5213 12536
rect 5155 12495 5213 12496
rect 5643 12536 5685 12545
rect 5643 12496 5644 12536
rect 5684 12496 5685 12536
rect 5643 12487 5685 12496
rect 5739 12536 5781 12545
rect 5739 12496 5740 12536
rect 5780 12496 5781 12536
rect 5739 12487 5781 12496
rect 6123 12536 6165 12545
rect 6123 12496 6124 12536
rect 6164 12496 6165 12536
rect 6123 12487 6165 12496
rect 6219 12536 6261 12545
rect 6219 12496 6220 12536
rect 6260 12496 6261 12536
rect 6219 12487 6261 12496
rect 6691 12536 6749 12537
rect 6691 12496 6700 12536
rect 6740 12496 6749 12536
rect 7947 12536 7989 12545
rect 6691 12495 6749 12496
rect 7179 12522 7221 12531
rect 7179 12482 7180 12522
rect 7220 12482 7221 12522
rect 7947 12496 7948 12536
rect 7988 12496 7989 12536
rect 7947 12487 7989 12496
rect 8043 12536 8085 12545
rect 8043 12496 8044 12536
rect 8084 12496 8085 12536
rect 8043 12487 8085 12496
rect 8323 12536 8381 12537
rect 8323 12496 8332 12536
rect 8372 12496 8381 12536
rect 8323 12495 8381 12496
rect 8803 12536 8861 12537
rect 8803 12496 8812 12536
rect 8852 12496 8861 12536
rect 8803 12495 8861 12496
rect 10051 12536 10109 12537
rect 10051 12496 10060 12536
rect 10100 12496 10109 12536
rect 10051 12495 10109 12496
rect 10819 12536 10877 12537
rect 10819 12496 10828 12536
rect 10868 12496 10877 12536
rect 10819 12495 10877 12496
rect 12067 12536 12125 12537
rect 12067 12496 12076 12536
rect 12116 12496 12125 12536
rect 12067 12495 12125 12496
rect 12939 12536 12981 12545
rect 12939 12496 12940 12536
rect 12980 12496 12981 12536
rect 12939 12487 12981 12496
rect 13035 12536 13077 12545
rect 13035 12496 13036 12536
rect 13076 12496 13077 12536
rect 13035 12487 13077 12496
rect 13131 12536 13173 12545
rect 13131 12496 13132 12536
rect 13172 12496 13173 12536
rect 13131 12487 13173 12496
rect 13795 12536 13853 12537
rect 13795 12496 13804 12536
rect 13844 12496 13853 12536
rect 13795 12495 13853 12496
rect 15043 12536 15101 12537
rect 15043 12496 15052 12536
rect 15092 12496 15101 12536
rect 15043 12495 15101 12496
rect 15619 12536 15677 12537
rect 15619 12496 15628 12536
rect 15668 12496 15677 12536
rect 15619 12495 15677 12496
rect 15811 12536 15869 12537
rect 15811 12496 15820 12536
rect 15860 12496 15869 12536
rect 15811 12495 15869 12496
rect 15915 12536 15957 12545
rect 15915 12496 15916 12536
rect 15956 12496 15957 12536
rect 15915 12487 15957 12496
rect 16107 12536 16149 12545
rect 16107 12496 16108 12536
rect 16148 12496 16149 12536
rect 16107 12487 16149 12496
rect 16387 12536 16445 12537
rect 16387 12496 16396 12536
rect 16436 12496 16445 12536
rect 16387 12495 16445 12496
rect 16683 12536 16725 12545
rect 16683 12496 16684 12536
rect 16724 12496 16725 12536
rect 16683 12487 16725 12496
rect 16779 12536 16821 12545
rect 16779 12496 16780 12536
rect 16820 12496 16821 12536
rect 16779 12487 16821 12496
rect 17259 12536 17301 12545
rect 17259 12496 17260 12536
rect 17300 12496 17301 12536
rect 17259 12487 17301 12496
rect 17451 12536 17493 12545
rect 17451 12496 17452 12536
rect 17492 12496 17493 12536
rect 17451 12487 17493 12496
rect 17731 12536 17789 12537
rect 17731 12496 17740 12536
rect 17780 12496 17789 12536
rect 17731 12495 17789 12496
rect 17931 12536 17973 12545
rect 17931 12496 17932 12536
rect 17972 12496 17973 12536
rect 17931 12487 17973 12496
rect 18027 12536 18069 12545
rect 18027 12496 18028 12536
rect 18068 12496 18069 12536
rect 18027 12487 18069 12496
rect 18123 12536 18165 12545
rect 18123 12496 18124 12536
rect 18164 12496 18165 12536
rect 18123 12487 18165 12496
rect 18219 12536 18261 12545
rect 18219 12496 18220 12536
rect 18260 12496 18261 12536
rect 18219 12487 18261 12496
rect 18403 12536 18461 12537
rect 18403 12496 18412 12536
rect 18452 12496 18461 12536
rect 18403 12495 18461 12496
rect 19651 12536 19709 12537
rect 19651 12496 19660 12536
rect 19700 12496 19709 12536
rect 19651 12495 19709 12496
rect 7179 12473 7221 12482
rect 17355 12452 17397 12461
rect 17355 12412 17356 12452
rect 17396 12412 17397 12452
rect 17355 12403 17397 12412
rect 7651 12368 7709 12369
rect 7651 12328 7660 12368
rect 7700 12328 7709 12368
rect 7651 12327 7709 12328
rect 17059 12368 17117 12369
rect 17059 12328 17068 12368
rect 17108 12328 17117 12368
rect 17059 12327 17117 12328
rect 5355 12284 5397 12293
rect 5355 12244 5356 12284
rect 5396 12244 5397 12284
rect 5355 12235 5397 12244
rect 8619 12284 8661 12293
rect 8619 12244 8620 12284
rect 8660 12244 8661 12284
rect 8619 12235 8661 12244
rect 13315 12284 13373 12285
rect 13315 12244 13324 12284
rect 13364 12244 13373 12284
rect 13315 12243 13373 12244
rect 16107 12284 16149 12293
rect 16107 12244 16108 12284
rect 16148 12244 16149 12284
rect 16107 12235 16149 12244
rect 19851 12284 19893 12293
rect 19851 12244 19852 12284
rect 19892 12244 19893 12284
rect 19851 12235 19893 12244
rect 1152 12116 20352 12140
rect 1152 12076 3688 12116
rect 3728 12076 3770 12116
rect 3810 12076 3852 12116
rect 3892 12076 3934 12116
rect 3974 12076 4016 12116
rect 4056 12076 18808 12116
rect 18848 12076 18890 12116
rect 18930 12076 18972 12116
rect 19012 12076 19054 12116
rect 19094 12076 19136 12116
rect 19176 12076 20352 12116
rect 1152 12052 20352 12076
rect 2667 11948 2709 11957
rect 2667 11908 2668 11948
rect 2708 11908 2709 11948
rect 2667 11899 2709 11908
rect 6891 11948 6933 11957
rect 6891 11908 6892 11948
rect 6932 11908 6933 11948
rect 6891 11899 6933 11908
rect 8715 11948 8757 11957
rect 8715 11908 8716 11948
rect 8756 11908 8757 11948
rect 8715 11899 8757 11908
rect 9187 11948 9245 11949
rect 9187 11908 9196 11948
rect 9236 11908 9245 11948
rect 9187 11907 9245 11908
rect 16491 11948 16533 11957
rect 16491 11908 16492 11948
rect 16532 11908 16533 11948
rect 16491 11899 16533 11908
rect 18507 11948 18549 11957
rect 18507 11908 18508 11948
rect 18548 11908 18549 11948
rect 18507 11899 18549 11908
rect 18699 11864 18741 11873
rect 18699 11824 18700 11864
rect 18740 11824 18741 11864
rect 18699 11815 18741 11824
rect 19075 11864 19133 11865
rect 19075 11824 19084 11864
rect 19124 11824 19133 11864
rect 19075 11823 19133 11824
rect 20139 11864 20181 11873
rect 20139 11824 20140 11864
rect 20180 11824 20181 11864
rect 20139 11815 20181 11824
rect 12363 11780 12405 11789
rect 12363 11740 12364 11780
rect 12404 11740 12405 11780
rect 12363 11731 12405 11740
rect 12459 11780 12501 11789
rect 12459 11740 12460 11780
rect 12500 11740 12501 11780
rect 12459 11731 12501 11740
rect 13987 11710 14045 11711
rect 1219 11696 1277 11697
rect 1219 11656 1228 11696
rect 1268 11656 1277 11696
rect 1219 11655 1277 11656
rect 2467 11696 2525 11697
rect 2467 11656 2476 11696
rect 2516 11656 2525 11696
rect 2467 11655 2525 11656
rect 3627 11696 3669 11705
rect 3627 11656 3628 11696
rect 3668 11656 3669 11696
rect 3627 11647 3669 11656
rect 3723 11696 3765 11705
rect 3723 11656 3724 11696
rect 3764 11656 3765 11696
rect 3723 11647 3765 11656
rect 3819 11696 3861 11705
rect 3819 11656 3820 11696
rect 3860 11656 3861 11696
rect 3819 11647 3861 11656
rect 5443 11696 5501 11697
rect 5443 11656 5452 11696
rect 5492 11656 5501 11696
rect 5443 11655 5501 11656
rect 6691 11696 6749 11697
rect 6691 11656 6700 11696
rect 6740 11656 6749 11696
rect 6691 11655 6749 11656
rect 7075 11696 7133 11697
rect 7075 11656 7084 11696
rect 7124 11656 7133 11696
rect 7075 11655 7133 11656
rect 8323 11696 8381 11697
rect 8323 11656 8332 11696
rect 8372 11656 8381 11696
rect 8323 11655 8381 11656
rect 8715 11696 8757 11705
rect 8715 11656 8716 11696
rect 8756 11656 8757 11696
rect 8715 11647 8757 11656
rect 9003 11696 9045 11705
rect 9003 11656 9004 11696
rect 9044 11656 9045 11696
rect 9003 11647 9045 11656
rect 9579 11696 9621 11705
rect 9579 11656 9580 11696
rect 9620 11656 9621 11696
rect 9579 11647 9621 11656
rect 9859 11696 9917 11697
rect 9859 11656 9868 11696
rect 9908 11656 9917 11696
rect 9859 11655 9917 11656
rect 10147 11696 10205 11697
rect 10147 11656 10156 11696
rect 10196 11656 10205 11696
rect 10147 11655 10205 11656
rect 11395 11696 11453 11697
rect 11395 11656 11404 11696
rect 11444 11656 11453 11696
rect 11395 11655 11453 11656
rect 11883 11696 11925 11705
rect 11883 11656 11884 11696
rect 11924 11656 11925 11696
rect 11883 11647 11925 11656
rect 11979 11696 12021 11705
rect 13419 11701 13461 11710
rect 11979 11656 11980 11696
rect 12020 11656 12021 11696
rect 11979 11647 12021 11656
rect 12931 11696 12989 11697
rect 12931 11656 12940 11696
rect 12980 11656 12989 11696
rect 12931 11655 12989 11656
rect 13419 11661 13420 11701
rect 13460 11661 13461 11701
rect 13419 11652 13461 11661
rect 13803 11696 13845 11705
rect 13803 11656 13804 11696
rect 13844 11656 13845 11696
rect 13987 11670 13996 11710
rect 14036 11670 14045 11710
rect 13987 11669 14045 11670
rect 14083 11696 14141 11697
rect 13803 11647 13845 11656
rect 14083 11656 14092 11696
rect 14132 11656 14141 11696
rect 14083 11655 14141 11656
rect 14283 11696 14325 11705
rect 14283 11656 14284 11696
rect 14324 11656 14325 11696
rect 14283 11647 14325 11656
rect 14379 11696 14421 11705
rect 14379 11656 14380 11696
rect 14420 11656 14421 11696
rect 14379 11647 14421 11656
rect 14475 11696 14517 11705
rect 14475 11656 14476 11696
rect 14516 11656 14517 11696
rect 14475 11647 14517 11656
rect 15043 11696 15101 11697
rect 15043 11656 15052 11696
rect 15092 11656 15101 11696
rect 15043 11655 15101 11656
rect 16291 11696 16349 11697
rect 16291 11656 16300 11696
rect 16340 11656 16349 11696
rect 16291 11655 16349 11656
rect 16867 11696 16925 11697
rect 16867 11656 16876 11696
rect 16916 11656 16925 11696
rect 16867 11655 16925 11656
rect 18115 11696 18173 11697
rect 18115 11656 18124 11696
rect 18164 11656 18173 11696
rect 18115 11655 18173 11656
rect 18699 11696 18741 11705
rect 18699 11656 18700 11696
rect 18740 11656 18741 11696
rect 18699 11647 18741 11656
rect 19371 11696 19413 11705
rect 19371 11656 19372 11696
rect 19412 11656 19413 11696
rect 19371 11647 19413 11656
rect 19467 11696 19509 11705
rect 19467 11656 19468 11696
rect 19508 11656 19509 11696
rect 19467 11647 19509 11656
rect 19747 11696 19805 11697
rect 19747 11656 19756 11696
rect 19796 11656 19805 11696
rect 19747 11655 19805 11656
rect 20035 11696 20093 11697
rect 20035 11656 20044 11696
rect 20084 11656 20093 11696
rect 20035 11655 20093 11656
rect 9483 11612 9525 11621
rect 9483 11572 9484 11612
rect 9524 11572 9525 11612
rect 9483 11563 9525 11572
rect 18315 11612 18357 11621
rect 18315 11572 18316 11612
rect 18356 11572 18357 11612
rect 18315 11563 18357 11572
rect 3523 11528 3581 11529
rect 3523 11488 3532 11528
rect 3572 11488 3581 11528
rect 3523 11487 3581 11488
rect 8523 11528 8565 11537
rect 8523 11488 8524 11528
rect 8564 11488 8565 11528
rect 8523 11479 8565 11488
rect 11595 11528 11637 11537
rect 11595 11488 11596 11528
rect 11636 11488 11637 11528
rect 11595 11479 11637 11488
rect 13611 11528 13653 11537
rect 13611 11488 13612 11528
rect 13652 11488 13653 11528
rect 13611 11479 13653 11488
rect 13891 11528 13949 11529
rect 13891 11488 13900 11528
rect 13940 11488 13949 11528
rect 13891 11487 13949 11488
rect 14563 11528 14621 11529
rect 14563 11488 14572 11528
rect 14612 11488 14621 11528
rect 14563 11487 14621 11488
rect 1152 11360 20452 11384
rect 1152 11320 4928 11360
rect 4968 11320 5010 11360
rect 5050 11320 5092 11360
rect 5132 11320 5174 11360
rect 5214 11320 5256 11360
rect 5296 11320 20048 11360
rect 20088 11320 20130 11360
rect 20170 11320 20212 11360
rect 20252 11320 20294 11360
rect 20334 11320 20376 11360
rect 20416 11320 20452 11360
rect 1152 11296 20452 11320
rect 2667 11192 2709 11201
rect 2667 11152 2668 11192
rect 2708 11152 2709 11192
rect 2667 11143 2709 11152
rect 4963 11192 5021 11193
rect 4963 11152 4972 11192
rect 5012 11152 5021 11192
rect 4963 11151 5021 11152
rect 7275 11192 7317 11201
rect 7275 11152 7276 11192
rect 7316 11152 7317 11192
rect 7275 11143 7317 11152
rect 7755 11192 7797 11201
rect 7755 11152 7756 11192
rect 7796 11152 7797 11192
rect 7755 11143 7797 11152
rect 9763 11192 9821 11193
rect 9763 11152 9772 11192
rect 9812 11152 9821 11192
rect 9763 11151 9821 11152
rect 11979 11192 12021 11201
rect 11979 11152 11980 11192
rect 12020 11152 12021 11192
rect 11979 11143 12021 11152
rect 20043 11192 20085 11201
rect 20043 11152 20044 11192
rect 20084 11152 20085 11192
rect 20043 11143 20085 11152
rect 3339 11108 3381 11117
rect 3339 11068 3340 11108
rect 3380 11068 3381 11108
rect 3339 11059 3381 11068
rect 12747 11108 12789 11117
rect 12747 11068 12748 11108
rect 12788 11068 12789 11108
rect 12747 11059 12789 11068
rect 1219 11024 1277 11025
rect 1219 10984 1228 11024
rect 1268 10984 1277 11024
rect 1219 10983 1277 10984
rect 2467 11024 2525 11025
rect 2467 10984 2476 11024
rect 2516 10984 2525 11024
rect 3715 11024 3773 11025
rect 2467 10983 2525 10984
rect 3435 10982 3477 10991
rect 3715 10984 3724 11024
rect 3764 10984 3773 11024
rect 3715 10983 3773 10984
rect 4395 11024 4437 11033
rect 4395 10984 4396 11024
rect 4436 10984 4437 11024
rect 3435 10942 3436 10982
rect 3476 10942 3477 10982
rect 4395 10975 4437 10984
rect 4491 11024 4533 11033
rect 4491 10984 4492 11024
rect 4532 10984 4533 11024
rect 4491 10975 4533 10984
rect 4683 11024 4725 11033
rect 4683 10984 4684 11024
rect 4724 10984 4725 11024
rect 4683 10975 4725 10984
rect 4875 11024 4917 11033
rect 4875 10984 4876 11024
rect 4916 10984 4917 11024
rect 4875 10975 4917 10984
rect 5067 11024 5109 11033
rect 5067 10984 5068 11024
rect 5108 10984 5109 11024
rect 5067 10975 5109 10984
rect 5155 11024 5213 11025
rect 5155 10984 5164 11024
rect 5204 10984 5213 11024
rect 5155 10983 5213 10984
rect 5827 11024 5885 11025
rect 5827 10984 5836 11024
rect 5876 10984 5885 11024
rect 5827 10983 5885 10984
rect 7075 11024 7133 11025
rect 7075 10984 7084 11024
rect 7124 10984 7133 11024
rect 7075 10983 7133 10984
rect 7947 11019 7989 11028
rect 7947 10979 7948 11019
rect 7988 10979 7989 11019
rect 8419 11024 8477 11025
rect 8419 10984 8428 11024
rect 8468 10984 8477 11024
rect 8419 10983 8477 10984
rect 8907 11024 8949 11033
rect 8907 10984 8908 11024
rect 8948 10984 8949 11024
rect 7947 10970 7989 10979
rect 8907 10975 8949 10984
rect 9387 11024 9429 11033
rect 9387 10984 9388 11024
rect 9428 10984 9429 11024
rect 9387 10975 9429 10984
rect 9483 11024 9525 11033
rect 9483 10984 9484 11024
rect 9524 10984 9525 11024
rect 9483 10975 9525 10984
rect 9867 11024 9909 11033
rect 9867 10984 9868 11024
rect 9908 10984 9909 11024
rect 9867 10975 9909 10984
rect 9963 11024 10005 11033
rect 9963 10984 9964 11024
rect 10004 10984 10005 11024
rect 9963 10975 10005 10984
rect 10059 11024 10101 11033
rect 10059 10984 10060 11024
rect 10100 10984 10101 11024
rect 10059 10975 10101 10984
rect 10531 11024 10589 11025
rect 10531 10984 10540 11024
rect 10580 10984 10589 11024
rect 10531 10983 10589 10984
rect 11779 11024 11837 11025
rect 11779 10984 11788 11024
rect 11828 10984 11837 11024
rect 11779 10983 11837 10984
rect 12843 11024 12885 11033
rect 12843 10984 12844 11024
rect 12884 10984 12885 11024
rect 12843 10975 12885 10984
rect 13123 11024 13181 11025
rect 13123 10984 13132 11024
rect 13172 10984 13181 11024
rect 13123 10983 13181 10984
rect 13419 11024 13461 11033
rect 13419 10984 13420 11024
rect 13460 10984 13461 11024
rect 13419 10975 13461 10984
rect 13707 11024 13749 11033
rect 13707 10984 13708 11024
rect 13748 10984 13749 11024
rect 13707 10975 13749 10984
rect 17731 11024 17789 11025
rect 17731 10984 17740 11024
rect 17780 10984 17789 11024
rect 17731 10983 17789 10984
rect 17835 11024 17877 11033
rect 17835 10984 17836 11024
rect 17876 10984 17877 11024
rect 17835 10975 17877 10984
rect 18019 11024 18077 11025
rect 18019 10984 18028 11024
rect 18068 10984 18077 11024
rect 18019 10983 18077 10984
rect 18315 11024 18357 11033
rect 18315 10984 18316 11024
rect 18356 10984 18357 11024
rect 18315 10975 18357 10984
rect 18411 11024 18453 11033
rect 18411 10984 18412 11024
rect 18452 10984 18453 11024
rect 18411 10975 18453 10984
rect 19363 11024 19421 11025
rect 19363 10984 19372 11024
rect 19412 10984 19421 11024
rect 19363 10983 19421 10984
rect 19851 11019 19893 11028
rect 19851 10979 19852 11019
rect 19892 10979 19893 11019
rect 19851 10970 19893 10979
rect 3435 10933 3477 10942
rect 9003 10940 9045 10949
rect 9003 10900 9004 10940
rect 9044 10900 9045 10940
rect 9003 10891 9045 10900
rect 13515 10940 13557 10949
rect 13515 10900 13516 10940
rect 13556 10900 13557 10940
rect 13515 10891 13557 10900
rect 18795 10940 18837 10949
rect 18795 10900 18796 10940
rect 18836 10900 18837 10940
rect 18795 10891 18837 10900
rect 18891 10940 18933 10949
rect 18891 10900 18892 10940
rect 18932 10900 18933 10940
rect 18891 10891 18933 10900
rect 3043 10856 3101 10857
rect 3043 10816 3052 10856
rect 3092 10816 3101 10856
rect 3043 10815 3101 10816
rect 12451 10856 12509 10857
rect 12451 10816 12460 10856
rect 12500 10816 12509 10856
rect 12451 10815 12509 10816
rect 18027 10856 18069 10865
rect 18027 10816 18028 10856
rect 18068 10816 18069 10856
rect 18027 10807 18069 10816
rect 1152 10604 20352 10628
rect 1152 10564 3688 10604
rect 3728 10564 3770 10604
rect 3810 10564 3852 10604
rect 3892 10564 3934 10604
rect 3974 10564 4016 10604
rect 4056 10564 18808 10604
rect 18848 10564 18890 10604
rect 18930 10564 18972 10604
rect 19012 10564 19054 10604
rect 19094 10564 19136 10604
rect 19176 10564 20352 10604
rect 1152 10540 20352 10564
rect 2667 10436 2709 10445
rect 2667 10396 2668 10436
rect 2708 10396 2709 10436
rect 2667 10387 2709 10396
rect 10635 10436 10677 10445
rect 10635 10396 10636 10436
rect 10676 10396 10677 10436
rect 10635 10387 10677 10396
rect 12843 10436 12885 10445
rect 12843 10396 12844 10436
rect 12884 10396 12885 10436
rect 12843 10387 12885 10396
rect 7939 10352 7997 10353
rect 7939 10312 7948 10352
rect 7988 10312 7997 10352
rect 7939 10311 7997 10312
rect 19075 10352 19133 10353
rect 19075 10312 19084 10352
rect 19124 10312 19133 10352
rect 19075 10311 19133 10312
rect 9195 10268 9237 10277
rect 9195 10228 9196 10268
rect 9236 10228 9237 10268
rect 9195 10219 9237 10228
rect 9291 10268 9333 10277
rect 9291 10228 9292 10268
rect 9332 10228 9333 10268
rect 9291 10219 9333 10228
rect 15435 10268 15477 10277
rect 15435 10228 15436 10268
rect 15476 10228 15477 10268
rect 15435 10219 15477 10228
rect 3051 10198 3093 10207
rect 1219 10184 1277 10185
rect 1219 10144 1228 10184
rect 1268 10144 1277 10184
rect 1219 10143 1277 10144
rect 2467 10184 2525 10185
rect 2467 10144 2476 10184
rect 2516 10144 2525 10184
rect 3051 10158 3052 10198
rect 3092 10158 3093 10198
rect 3051 10149 3093 10158
rect 3523 10184 3581 10185
rect 2467 10143 2525 10144
rect 3523 10144 3532 10184
rect 3572 10144 3581 10184
rect 3523 10143 3581 10144
rect 4011 10184 4053 10193
rect 4011 10144 4012 10184
rect 4052 10144 4053 10184
rect 4011 10135 4053 10144
rect 4107 10184 4149 10193
rect 4107 10144 4108 10184
rect 4148 10144 4149 10184
rect 4107 10135 4149 10144
rect 4491 10184 4533 10193
rect 4491 10144 4492 10184
rect 4532 10144 4533 10184
rect 4491 10135 4533 10144
rect 4587 10184 4629 10193
rect 4587 10144 4588 10184
rect 4628 10144 4629 10184
rect 4587 10135 4629 10144
rect 7467 10184 7509 10193
rect 7467 10144 7468 10184
rect 7508 10144 7509 10184
rect 7467 10135 7509 10144
rect 7563 10184 7605 10193
rect 7563 10144 7564 10184
rect 7604 10144 7605 10184
rect 7563 10135 7605 10144
rect 7659 10184 7701 10193
rect 7659 10144 7660 10184
rect 7700 10144 7701 10184
rect 7659 10135 7701 10144
rect 7755 10184 7797 10193
rect 7755 10144 7756 10184
rect 7796 10144 7797 10184
rect 7755 10135 7797 10144
rect 8139 10184 8181 10193
rect 8139 10144 8140 10184
rect 8180 10144 8181 10184
rect 8139 10135 8181 10144
rect 8235 10184 8277 10193
rect 8235 10144 8236 10184
rect 8276 10144 8277 10184
rect 8235 10135 8277 10144
rect 8331 10184 8373 10193
rect 8331 10144 8332 10184
rect 8372 10144 8373 10184
rect 8331 10135 8373 10144
rect 8715 10184 8757 10193
rect 8715 10144 8716 10184
rect 8756 10144 8757 10184
rect 8715 10135 8757 10144
rect 8811 10184 8853 10193
rect 10251 10189 10293 10198
rect 16539 10193 16581 10202
rect 8811 10144 8812 10184
rect 8852 10144 8853 10184
rect 8811 10135 8853 10144
rect 9763 10184 9821 10185
rect 9763 10144 9772 10184
rect 9812 10144 9821 10184
rect 9763 10143 9821 10144
rect 10251 10149 10252 10189
rect 10292 10149 10293 10189
rect 10251 10140 10293 10149
rect 10635 10184 10677 10193
rect 10635 10144 10636 10184
rect 10676 10144 10677 10184
rect 10635 10135 10677 10144
rect 10827 10184 10869 10193
rect 10827 10144 10828 10184
rect 10868 10144 10869 10184
rect 10827 10135 10869 10144
rect 10915 10184 10973 10185
rect 10915 10144 10924 10184
rect 10964 10144 10973 10184
rect 10915 10143 10973 10144
rect 11395 10184 11453 10185
rect 11395 10144 11404 10184
rect 11444 10144 11453 10184
rect 11395 10143 11453 10144
rect 12643 10184 12701 10185
rect 12643 10144 12652 10184
rect 12692 10144 12701 10184
rect 12643 10143 12701 10144
rect 13219 10184 13277 10185
rect 13219 10144 13228 10184
rect 13268 10144 13277 10184
rect 13219 10143 13277 10144
rect 14467 10184 14525 10185
rect 14467 10144 14476 10184
rect 14516 10144 14525 10184
rect 14467 10143 14525 10144
rect 14955 10184 14997 10193
rect 14955 10144 14956 10184
rect 14996 10144 14997 10184
rect 14955 10135 14997 10144
rect 15051 10184 15093 10193
rect 15051 10144 15052 10184
rect 15092 10144 15093 10184
rect 15051 10135 15093 10144
rect 15531 10184 15573 10193
rect 15531 10144 15532 10184
rect 15572 10144 15573 10184
rect 15531 10135 15573 10144
rect 16003 10184 16061 10185
rect 16003 10144 16012 10184
rect 16052 10144 16061 10184
rect 16539 10153 16540 10193
rect 16580 10153 16581 10193
rect 16539 10144 16581 10153
rect 17443 10184 17501 10185
rect 17443 10144 17452 10184
rect 17492 10144 17501 10184
rect 16003 10143 16061 10144
rect 17443 10143 17501 10144
rect 18691 10184 18749 10185
rect 18691 10144 18700 10184
rect 18740 10144 18749 10184
rect 18691 10143 18749 10144
rect 19467 10184 19509 10193
rect 19467 10144 19468 10184
rect 19508 10144 19509 10184
rect 19467 10135 19509 10144
rect 19747 10184 19805 10185
rect 19747 10144 19756 10184
rect 19796 10144 19805 10184
rect 19747 10143 19805 10144
rect 2859 10100 2901 10109
rect 2859 10060 2860 10100
rect 2900 10060 2901 10100
rect 2859 10051 2901 10060
rect 10443 10100 10485 10109
rect 10443 10060 10444 10100
rect 10484 10060 10485 10100
rect 10443 10051 10485 10060
rect 14667 10100 14709 10109
rect 14667 10060 14668 10100
rect 14708 10060 14709 10100
rect 14667 10051 14709 10060
rect 16683 10100 16725 10109
rect 16683 10060 16684 10100
rect 16724 10060 16725 10100
rect 16683 10051 16725 10060
rect 18891 10100 18933 10109
rect 18891 10060 18892 10100
rect 18932 10060 18933 10100
rect 18891 10051 18933 10060
rect 19371 10100 19413 10109
rect 19371 10060 19372 10100
rect 19412 10060 19413 10100
rect 19371 10051 19413 10060
rect 1152 9848 20452 9872
rect 1152 9808 4928 9848
rect 4968 9808 5010 9848
rect 5050 9808 5092 9848
rect 5132 9808 5174 9848
rect 5214 9808 5256 9848
rect 5296 9808 20048 9848
rect 20088 9808 20130 9848
rect 20170 9808 20212 9848
rect 20252 9808 20294 9848
rect 20334 9808 20376 9848
rect 20416 9808 20452 9848
rect 1152 9784 20452 9808
rect 3723 9680 3765 9689
rect 3723 9640 3724 9680
rect 3764 9640 3765 9680
rect 3723 9631 3765 9640
rect 5739 9680 5781 9689
rect 5739 9640 5740 9680
rect 5780 9640 5781 9680
rect 5739 9631 5781 9640
rect 9675 9680 9717 9689
rect 9675 9640 9676 9680
rect 9716 9640 9717 9680
rect 9675 9631 9717 9640
rect 10539 9680 10581 9689
rect 10539 9640 10540 9680
rect 10580 9640 10581 9680
rect 10539 9631 10581 9640
rect 14667 9680 14709 9689
rect 14667 9640 14668 9680
rect 14708 9640 14709 9680
rect 14667 9631 14709 9640
rect 16587 9680 16629 9689
rect 16587 9640 16588 9680
rect 16628 9640 16629 9680
rect 16587 9631 16629 9640
rect 19755 9680 19797 9689
rect 19755 9640 19756 9680
rect 19796 9640 19797 9680
rect 19755 9631 19797 9640
rect 2955 9596 2997 9605
rect 2955 9556 2956 9596
rect 2996 9556 2997 9596
rect 2955 9547 2997 9556
rect 5547 9596 5589 9605
rect 5547 9556 5548 9596
rect 5588 9556 5589 9596
rect 5547 9547 5589 9556
rect 9195 9596 9237 9605
rect 9195 9556 9196 9596
rect 9236 9556 9237 9596
rect 9195 9547 9237 9556
rect 12651 9596 12693 9605
rect 12651 9556 12652 9596
rect 12692 9556 12693 9596
rect 12651 9547 12693 9556
rect 1507 9512 1565 9513
rect 1507 9472 1516 9512
rect 1556 9472 1565 9512
rect 1507 9471 1565 9472
rect 2755 9512 2813 9513
rect 2755 9472 2764 9512
rect 2804 9472 2813 9512
rect 2755 9471 2813 9472
rect 3339 9512 3381 9521
rect 3339 9472 3340 9512
rect 3380 9472 3381 9512
rect 3339 9463 3381 9472
rect 3435 9512 3477 9521
rect 3435 9472 3436 9512
rect 3476 9472 3477 9512
rect 3435 9463 3477 9472
rect 3531 9512 3573 9521
rect 3531 9472 3532 9512
rect 3572 9472 3573 9512
rect 3531 9463 3573 9472
rect 4099 9512 4157 9513
rect 4099 9472 4108 9512
rect 4148 9472 4157 9512
rect 4099 9471 4157 9472
rect 5347 9512 5405 9513
rect 5347 9472 5356 9512
rect 5396 9472 5405 9512
rect 6403 9512 6461 9513
rect 5347 9471 5405 9472
rect 5883 9470 5925 9479
rect 6403 9472 6412 9512
rect 6452 9472 6461 9512
rect 6403 9471 6461 9472
rect 6987 9512 7029 9521
rect 6987 9472 6988 9512
rect 7028 9472 7029 9512
rect 5883 9430 5884 9470
rect 5924 9430 5925 9470
rect 6987 9463 7029 9472
rect 7371 9512 7413 9521
rect 7371 9472 7372 9512
rect 7412 9472 7413 9512
rect 7371 9463 7413 9472
rect 7467 9512 7509 9521
rect 7467 9472 7468 9512
rect 7508 9472 7509 9512
rect 7467 9463 7509 9472
rect 7747 9512 7805 9513
rect 7747 9472 7756 9512
rect 7796 9472 7805 9512
rect 7747 9471 7805 9472
rect 8995 9512 9053 9513
rect 8995 9472 9004 9512
rect 9044 9472 9053 9512
rect 8995 9471 9053 9472
rect 9867 9512 9909 9521
rect 9867 9472 9868 9512
rect 9908 9472 9909 9512
rect 9867 9463 9909 9472
rect 10059 9512 10101 9521
rect 10059 9472 10060 9512
rect 10100 9472 10101 9512
rect 9955 9470 10013 9471
rect 5883 9421 5925 9430
rect 6891 9428 6933 9437
rect 9955 9430 9964 9470
rect 10004 9430 10013 9470
rect 10059 9463 10101 9472
rect 10347 9512 10389 9521
rect 10347 9472 10348 9512
rect 10388 9472 10389 9512
rect 10347 9463 10389 9472
rect 10635 9512 10677 9521
rect 10635 9472 10636 9512
rect 10676 9472 10677 9512
rect 10635 9463 10677 9472
rect 11203 9512 11261 9513
rect 11203 9472 11212 9512
rect 11252 9472 11261 9512
rect 11203 9471 11261 9472
rect 12451 9512 12509 9513
rect 12451 9472 12460 9512
rect 12500 9472 12509 9512
rect 12451 9471 12509 9472
rect 12939 9512 12981 9521
rect 12939 9472 12940 9512
rect 12980 9472 12981 9512
rect 12939 9463 12981 9472
rect 13035 9512 13077 9521
rect 13035 9472 13036 9512
rect 13076 9472 13077 9512
rect 13035 9463 13077 9472
rect 13515 9512 13557 9521
rect 13515 9472 13516 9512
rect 13556 9472 13557 9512
rect 13515 9463 13557 9472
rect 13987 9512 14045 9513
rect 13987 9472 13996 9512
rect 14036 9472 14045 9512
rect 14851 9512 14909 9513
rect 13987 9471 14045 9472
rect 14475 9498 14517 9507
rect 14475 9458 14476 9498
rect 14516 9458 14517 9498
rect 14851 9472 14860 9512
rect 14900 9472 14909 9512
rect 14851 9471 14909 9472
rect 15139 9512 15197 9513
rect 15139 9472 15148 9512
rect 15188 9472 15197 9512
rect 15139 9471 15197 9472
rect 16387 9512 16445 9513
rect 16387 9472 16396 9512
rect 16436 9472 16445 9512
rect 16387 9471 16445 9472
rect 16971 9512 17013 9521
rect 16971 9472 16972 9512
rect 17012 9472 17013 9512
rect 16971 9463 17013 9472
rect 17067 9512 17109 9521
rect 17067 9472 17068 9512
rect 17108 9472 17109 9512
rect 17067 9463 17109 9472
rect 17163 9512 17205 9521
rect 17163 9472 17164 9512
rect 17204 9472 17205 9512
rect 17163 9463 17205 9472
rect 17259 9512 17301 9521
rect 17259 9472 17260 9512
rect 17300 9472 17301 9512
rect 17259 9463 17301 9472
rect 17643 9512 17685 9521
rect 17643 9472 17644 9512
rect 17684 9472 17685 9512
rect 17643 9463 17685 9472
rect 18027 9512 18069 9521
rect 18027 9472 18028 9512
rect 18068 9472 18069 9512
rect 18027 9463 18069 9472
rect 18123 9512 18165 9521
rect 20139 9518 20181 9527
rect 18123 9472 18124 9512
rect 18164 9472 18165 9512
rect 18123 9463 18165 9472
rect 19075 9512 19133 9513
rect 19075 9472 19084 9512
rect 19124 9472 19133 9512
rect 19075 9471 19133 9472
rect 19563 9507 19605 9516
rect 19563 9467 19564 9507
rect 19604 9467 19605 9507
rect 19939 9512 19997 9513
rect 19939 9472 19948 9512
rect 19988 9472 19997 9512
rect 19939 9471 19997 9472
rect 20139 9478 20140 9518
rect 20180 9478 20181 9518
rect 20139 9469 20181 9478
rect 20227 9512 20285 9513
rect 20227 9472 20236 9512
rect 20276 9472 20285 9512
rect 20227 9471 20285 9472
rect 19563 9458 19605 9467
rect 14475 9449 14517 9458
rect 9955 9429 10013 9430
rect 6891 9388 6892 9428
rect 6932 9388 6933 9428
rect 6891 9379 6933 9388
rect 13419 9428 13461 9437
rect 13419 9388 13420 9428
rect 13460 9388 13461 9428
rect 13419 9379 13461 9388
rect 18507 9428 18549 9437
rect 18507 9388 18508 9428
rect 18548 9388 18549 9428
rect 18507 9379 18549 9388
rect 18603 9428 18645 9437
rect 18603 9388 18604 9428
rect 18644 9388 18645 9428
rect 18603 9379 18645 9388
rect 17451 9344 17493 9353
rect 17451 9304 17452 9344
rect 17492 9304 17493 9344
rect 17451 9295 17493 9304
rect 17643 9344 17685 9353
rect 17643 9304 17644 9344
rect 17684 9304 17685 9344
rect 17643 9295 17685 9304
rect 14955 9260 14997 9269
rect 14955 9220 14956 9260
rect 14996 9220 14997 9260
rect 14955 9211 14997 9220
rect 19947 9260 19989 9269
rect 19947 9220 19948 9260
rect 19988 9220 19989 9260
rect 19947 9211 19989 9220
rect 1152 9092 20352 9116
rect 1152 9052 3688 9092
rect 3728 9052 3770 9092
rect 3810 9052 3852 9092
rect 3892 9052 3934 9092
rect 3974 9052 4016 9092
rect 4056 9052 18808 9092
rect 18848 9052 18890 9092
rect 18930 9052 18972 9092
rect 19012 9052 19054 9092
rect 19094 9052 19136 9092
rect 19176 9052 20352 9092
rect 1152 9028 20352 9052
rect 2667 8924 2709 8933
rect 2667 8884 2668 8924
rect 2708 8884 2709 8924
rect 2667 8875 2709 8884
rect 5739 8924 5781 8933
rect 5739 8884 5740 8924
rect 5780 8884 5781 8924
rect 5739 8875 5781 8884
rect 14475 8924 14517 8933
rect 14475 8884 14476 8924
rect 14516 8884 14517 8924
rect 14475 8875 14517 8884
rect 3043 8840 3101 8841
rect 3043 8800 3052 8840
rect 3092 8800 3101 8840
rect 3043 8799 3101 8800
rect 4491 8840 4533 8849
rect 4491 8800 4492 8840
rect 4532 8800 4533 8840
rect 4491 8791 4533 8800
rect 9771 8840 9813 8849
rect 9771 8800 9772 8840
rect 9812 8800 9813 8840
rect 9771 8791 9813 8800
rect 14947 8840 15005 8841
rect 14947 8800 14956 8840
rect 14996 8800 15005 8840
rect 14947 8799 15005 8800
rect 19275 8840 19317 8849
rect 19275 8800 19276 8840
rect 19316 8800 19317 8840
rect 19275 8791 19317 8800
rect 20139 8840 20181 8849
rect 20139 8800 20140 8840
rect 20180 8800 20181 8840
rect 20139 8791 20181 8800
rect 10539 8756 10581 8765
rect 10539 8716 10540 8756
rect 10580 8716 10581 8756
rect 10539 8707 10581 8716
rect 10635 8756 10677 8765
rect 10635 8716 10636 8756
rect 10676 8716 10677 8756
rect 10635 8707 10677 8716
rect 19939 8756 19997 8757
rect 19939 8716 19948 8756
rect 19988 8716 19997 8756
rect 19939 8715 19997 8716
rect 4299 8683 4341 8692
rect 1219 8672 1277 8673
rect 1219 8632 1228 8672
rect 1268 8632 1277 8672
rect 1219 8631 1277 8632
rect 2467 8672 2525 8673
rect 2467 8632 2476 8672
rect 2516 8632 2525 8672
rect 2467 8631 2525 8632
rect 3435 8672 3477 8681
rect 3435 8632 3436 8672
rect 3476 8632 3477 8672
rect 3435 8623 3477 8632
rect 3715 8672 3773 8673
rect 3715 8632 3724 8672
rect 3764 8632 3773 8672
rect 3715 8631 3773 8632
rect 4003 8672 4061 8673
rect 4003 8632 4012 8672
rect 4052 8632 4061 8672
rect 4003 8631 4061 8632
rect 4107 8672 4149 8681
rect 4107 8632 4108 8672
rect 4148 8632 4149 8672
rect 4299 8643 4300 8683
rect 4340 8643 4341 8683
rect 4299 8634 4341 8643
rect 4491 8672 4533 8681
rect 4107 8623 4149 8632
rect 4491 8632 4492 8672
rect 4532 8632 4533 8672
rect 4491 8623 4533 8632
rect 4779 8672 4821 8681
rect 4779 8632 4780 8672
rect 4820 8632 4821 8672
rect 4779 8623 4821 8632
rect 5923 8672 5981 8673
rect 5923 8632 5932 8672
rect 5972 8632 5981 8672
rect 5923 8631 5981 8632
rect 7171 8672 7229 8673
rect 7171 8632 7180 8672
rect 7220 8632 7229 8672
rect 7171 8631 7229 8632
rect 8323 8672 8381 8673
rect 8323 8632 8332 8672
rect 8372 8632 8381 8672
rect 8323 8631 8381 8632
rect 9571 8672 9629 8673
rect 9571 8632 9580 8672
rect 9620 8632 9629 8672
rect 9571 8631 9629 8632
rect 10059 8672 10101 8681
rect 10059 8632 10060 8672
rect 10100 8632 10101 8672
rect 10059 8623 10101 8632
rect 10155 8672 10197 8681
rect 11595 8677 11637 8686
rect 10155 8632 10156 8672
rect 10196 8632 10197 8672
rect 10155 8623 10197 8632
rect 11107 8672 11165 8673
rect 11107 8632 11116 8672
rect 11156 8632 11165 8672
rect 11107 8631 11165 8632
rect 11595 8637 11596 8677
rect 11636 8637 11637 8677
rect 11595 8628 11637 8637
rect 13027 8672 13085 8673
rect 13027 8632 13036 8672
rect 13076 8632 13085 8672
rect 13027 8631 13085 8632
rect 14275 8672 14333 8673
rect 14275 8632 14284 8672
rect 14324 8632 14333 8672
rect 14275 8631 14333 8632
rect 14763 8672 14805 8681
rect 14763 8632 14764 8672
rect 14804 8632 14805 8672
rect 14763 8623 14805 8632
rect 14955 8672 14997 8681
rect 14955 8632 14956 8672
rect 14996 8632 14997 8672
rect 14955 8623 14997 8632
rect 15051 8672 15093 8681
rect 15051 8632 15052 8672
rect 15092 8632 15093 8672
rect 15051 8623 15093 8632
rect 15235 8672 15293 8673
rect 15235 8632 15244 8672
rect 15284 8632 15293 8672
rect 15235 8631 15293 8632
rect 15331 8672 15389 8673
rect 15331 8632 15340 8672
rect 15380 8632 15389 8672
rect 15331 8631 15389 8632
rect 15531 8672 15573 8681
rect 15531 8632 15532 8672
rect 15572 8632 15573 8672
rect 15531 8623 15573 8632
rect 15627 8672 15669 8681
rect 15627 8632 15628 8672
rect 15668 8632 15669 8672
rect 15627 8623 15669 8632
rect 15720 8672 15778 8673
rect 15720 8632 15729 8672
rect 15769 8632 15778 8672
rect 15720 8631 15778 8632
rect 16195 8672 16253 8673
rect 16195 8632 16204 8672
rect 16244 8632 16253 8672
rect 16195 8631 16253 8632
rect 17443 8672 17501 8673
rect 17443 8632 17452 8672
rect 17492 8632 17501 8672
rect 17443 8631 17501 8632
rect 17827 8672 17885 8673
rect 17827 8632 17836 8672
rect 17876 8632 17885 8672
rect 17827 8631 17885 8632
rect 19075 8672 19133 8673
rect 19075 8632 19084 8672
rect 19124 8632 19133 8672
rect 19075 8631 19133 8632
rect 19467 8672 19509 8681
rect 19467 8632 19468 8672
rect 19508 8632 19509 8672
rect 19467 8623 19509 8632
rect 19563 8672 19605 8681
rect 19563 8632 19564 8672
rect 19604 8632 19605 8672
rect 19563 8623 19605 8632
rect 19659 8672 19701 8681
rect 19659 8632 19660 8672
rect 19700 8632 19701 8672
rect 19659 8623 19701 8632
rect 3339 8588 3381 8597
rect 3339 8548 3340 8588
rect 3380 8548 3381 8588
rect 3339 8539 3381 8548
rect 11787 8588 11829 8597
rect 11787 8548 11788 8588
rect 11828 8548 11829 8588
rect 11787 8539 11829 8548
rect 4195 8504 4253 8505
rect 4195 8464 4204 8504
rect 4244 8464 4253 8504
rect 4195 8463 4253 8464
rect 15427 8504 15485 8505
rect 15427 8464 15436 8504
rect 15476 8464 15485 8504
rect 15427 8463 15485 8464
rect 17643 8504 17685 8513
rect 17643 8464 17644 8504
rect 17684 8464 17685 8504
rect 17643 8455 17685 8464
rect 19747 8504 19805 8505
rect 19747 8464 19756 8504
rect 19796 8464 19805 8504
rect 19747 8463 19805 8464
rect 1152 8336 20452 8360
rect 1152 8296 4928 8336
rect 4968 8296 5010 8336
rect 5050 8296 5092 8336
rect 5132 8296 5174 8336
rect 5214 8296 5256 8336
rect 5296 8296 20048 8336
rect 20088 8296 20130 8336
rect 20170 8296 20212 8336
rect 20252 8296 20294 8336
rect 20334 8296 20376 8336
rect 20416 8296 20452 8336
rect 1152 8272 20452 8296
rect 4395 8168 4437 8177
rect 4395 8128 4396 8168
rect 4436 8128 4437 8168
rect 4395 8119 4437 8128
rect 9867 8168 9909 8177
rect 9867 8128 9868 8168
rect 9908 8128 9909 8168
rect 9867 8119 9909 8128
rect 11499 8168 11541 8177
rect 11499 8128 11500 8168
rect 11540 8128 11541 8168
rect 11499 8119 11541 8128
rect 15339 8168 15381 8177
rect 15339 8128 15340 8168
rect 15380 8128 15381 8168
rect 15339 8119 15381 8128
rect 18603 8168 18645 8177
rect 18603 8128 18604 8168
rect 18644 8128 18645 8168
rect 18603 8119 18645 8128
rect 8139 8084 8181 8093
rect 8139 8044 8140 8084
rect 8180 8044 8181 8084
rect 8139 8035 8181 8044
rect 1995 8000 2037 8009
rect 1995 7960 1996 8000
rect 2036 7960 2037 8000
rect 1995 7951 2037 7960
rect 2091 8000 2133 8009
rect 2091 7960 2092 8000
rect 2132 7960 2133 8000
rect 2091 7951 2133 7960
rect 2187 8000 2229 8009
rect 2187 7960 2188 8000
rect 2228 7960 2229 8000
rect 2187 7951 2229 7960
rect 2667 8000 2709 8009
rect 2667 7960 2668 8000
rect 2708 7960 2709 8000
rect 2667 7951 2709 7960
rect 2763 8000 2805 8009
rect 2763 7960 2764 8000
rect 2804 7960 2805 8000
rect 2763 7951 2805 7960
rect 3715 8000 3773 8001
rect 3715 7960 3724 8000
rect 3764 7960 3773 8000
rect 4675 8000 4733 8001
rect 3715 7959 3773 7960
rect 4203 7986 4245 7995
rect 4203 7946 4204 7986
rect 4244 7946 4245 7986
rect 4675 7960 4684 8000
rect 4724 7960 4733 8000
rect 4675 7959 4733 7960
rect 5923 8000 5981 8001
rect 5923 7960 5932 8000
rect 5972 7960 5981 8000
rect 5923 7959 5981 7960
rect 6411 8000 6453 8009
rect 6411 7960 6412 8000
rect 6452 7960 6453 8000
rect 6411 7951 6453 7960
rect 6507 8000 6549 8009
rect 6507 7960 6508 8000
rect 6548 7960 6549 8000
rect 6507 7951 6549 7960
rect 6987 8000 7029 8009
rect 6987 7960 6988 8000
rect 7028 7960 7029 8000
rect 6987 7951 7029 7960
rect 7459 8000 7517 8001
rect 7459 7960 7468 8000
rect 7508 7960 7517 8000
rect 8419 8000 8477 8001
rect 7459 7959 7517 7960
rect 7947 7986 7989 7995
rect 4203 7937 4245 7946
rect 7947 7946 7948 7986
rect 7988 7946 7989 7986
rect 8419 7960 8428 8000
rect 8468 7960 8477 8000
rect 8419 7959 8477 7960
rect 9667 8000 9725 8001
rect 9667 7960 9676 8000
rect 9716 7960 9725 8000
rect 9667 7959 9725 7960
rect 10051 8000 10109 8001
rect 10051 7960 10060 8000
rect 10100 7960 10109 8000
rect 10051 7959 10109 7960
rect 11299 8000 11357 8001
rect 11299 7960 11308 8000
rect 11348 7960 11357 8000
rect 11299 7959 11357 7960
rect 11683 8000 11741 8001
rect 11683 7960 11692 8000
rect 11732 7960 11741 8000
rect 11683 7959 11741 7960
rect 12931 8000 12989 8001
rect 12931 7960 12940 8000
rect 12980 7960 12989 8000
rect 12931 7959 12989 7960
rect 13891 8000 13949 8001
rect 13891 7960 13900 8000
rect 13940 7960 13949 8000
rect 13891 7959 13949 7960
rect 15139 8000 15197 8001
rect 15139 7960 15148 8000
rect 15188 7960 15197 8000
rect 15139 7959 15197 7960
rect 15523 8000 15581 8001
rect 15523 7960 15532 8000
rect 15572 7960 15581 8000
rect 15523 7959 15581 7960
rect 16771 8000 16829 8001
rect 16771 7960 16780 8000
rect 16820 7960 16829 8000
rect 16771 7959 16829 7960
rect 18027 8000 18069 8009
rect 18027 7960 18028 8000
rect 18068 7960 18069 8000
rect 18027 7951 18069 7960
rect 18315 8000 18357 8009
rect 18315 7960 18316 8000
rect 18356 7960 18357 8000
rect 18315 7951 18357 7960
rect 18499 8000 18557 8001
rect 18499 7960 18508 8000
rect 18548 7960 18557 8000
rect 18499 7959 18557 7960
rect 19371 8000 19413 8009
rect 19371 7960 19372 8000
rect 19412 7960 19413 8000
rect 19371 7951 19413 7960
rect 19467 8000 19509 8009
rect 19467 7960 19468 8000
rect 19508 7960 19509 8000
rect 19467 7951 19509 7960
rect 19747 8000 19805 8001
rect 19747 7960 19756 8000
rect 19796 7960 19805 8000
rect 19747 7959 19805 7960
rect 7947 7937 7989 7946
rect 3147 7916 3189 7925
rect 3147 7876 3148 7916
rect 3188 7876 3189 7916
rect 3147 7867 3189 7876
rect 3243 7916 3285 7925
rect 3243 7876 3244 7916
rect 3284 7876 3285 7916
rect 3243 7867 3285 7876
rect 6891 7916 6933 7925
rect 6891 7876 6892 7916
rect 6932 7876 6933 7916
rect 6891 7867 6933 7876
rect 6123 7832 6165 7841
rect 6123 7792 6124 7832
rect 6164 7792 6165 7832
rect 6123 7783 6165 7792
rect 2371 7748 2429 7749
rect 2371 7708 2380 7748
rect 2420 7708 2429 7748
rect 2371 7707 2429 7708
rect 13131 7748 13173 7757
rect 13131 7708 13132 7748
rect 13172 7708 13173 7748
rect 13131 7699 13173 7708
rect 16971 7748 17013 7757
rect 16971 7708 16972 7748
rect 17012 7708 17013 7748
rect 16971 7699 17013 7708
rect 18315 7748 18357 7757
rect 18315 7708 18316 7748
rect 18356 7708 18357 7748
rect 18315 7699 18357 7708
rect 19075 7748 19133 7749
rect 19075 7708 19084 7748
rect 19124 7708 19133 7748
rect 19075 7707 19133 7708
rect 1152 7580 20352 7604
rect 1152 7540 3688 7580
rect 3728 7540 3770 7580
rect 3810 7540 3852 7580
rect 3892 7540 3934 7580
rect 3974 7540 4016 7580
rect 4056 7540 18808 7580
rect 18848 7540 18890 7580
rect 18930 7540 18972 7580
rect 19012 7540 19054 7580
rect 19094 7540 19136 7580
rect 19176 7540 20352 7580
rect 1152 7516 20352 7540
rect 2667 7412 2709 7421
rect 2667 7372 2668 7412
rect 2708 7372 2709 7412
rect 2667 7363 2709 7372
rect 2859 7412 2901 7421
rect 2859 7372 2860 7412
rect 2900 7372 2901 7412
rect 2859 7363 2901 7372
rect 7851 7412 7893 7421
rect 7851 7372 7852 7412
rect 7892 7372 7893 7412
rect 7851 7363 7893 7372
rect 15723 7412 15765 7421
rect 15723 7372 15724 7412
rect 15764 7372 15765 7412
rect 15723 7363 15765 7372
rect 19755 7412 19797 7421
rect 19755 7372 19756 7412
rect 19796 7372 19797 7412
rect 19755 7363 19797 7372
rect 13227 7174 13269 7183
rect 1219 7160 1277 7161
rect 1219 7120 1228 7160
rect 1268 7120 1277 7160
rect 1219 7119 1277 7120
rect 2467 7160 2525 7161
rect 2467 7120 2476 7160
rect 2516 7120 2525 7160
rect 2467 7119 2525 7120
rect 3043 7160 3101 7161
rect 3043 7120 3052 7160
rect 3092 7120 3101 7160
rect 3043 7119 3101 7120
rect 4291 7160 4349 7161
rect 4291 7120 4300 7160
rect 4340 7120 4349 7160
rect 4291 7119 4349 7120
rect 4491 7160 4533 7169
rect 4491 7120 4492 7160
rect 4532 7120 4533 7160
rect 4491 7111 4533 7120
rect 4587 7160 4629 7169
rect 4587 7120 4588 7160
rect 4628 7120 4629 7160
rect 4587 7111 4629 7120
rect 4683 7160 4725 7169
rect 4683 7120 4684 7160
rect 4724 7120 4725 7160
rect 4683 7111 4725 7120
rect 6403 7160 6461 7161
rect 6403 7120 6412 7160
rect 6452 7120 6461 7160
rect 6403 7119 6461 7120
rect 7651 7160 7709 7161
rect 7651 7120 7660 7160
rect 7700 7120 7709 7160
rect 7651 7119 7709 7120
rect 8323 7160 8381 7161
rect 8323 7120 8332 7160
rect 8372 7120 8381 7160
rect 8323 7119 8381 7120
rect 9571 7160 9629 7161
rect 9571 7120 9580 7160
rect 9620 7120 9629 7160
rect 9571 7119 9629 7120
rect 9955 7160 10013 7161
rect 9955 7120 9964 7160
rect 10004 7120 10013 7160
rect 9955 7119 10013 7120
rect 11203 7160 11261 7161
rect 11203 7120 11212 7160
rect 11252 7120 11261 7160
rect 11203 7119 11261 7120
rect 11691 7160 11733 7169
rect 11691 7120 11692 7160
rect 11732 7120 11733 7160
rect 11691 7111 11733 7120
rect 11787 7160 11829 7169
rect 11787 7120 11788 7160
rect 11828 7120 11829 7160
rect 11787 7111 11829 7120
rect 12171 7160 12213 7169
rect 12171 7120 12172 7160
rect 12212 7120 12213 7160
rect 12171 7111 12213 7120
rect 12267 7160 12309 7169
rect 12267 7120 12268 7160
rect 12308 7120 12309 7160
rect 12267 7111 12309 7120
rect 12739 7160 12797 7161
rect 12739 7120 12748 7160
rect 12788 7120 12797 7160
rect 13227 7134 13228 7174
rect 13268 7134 13269 7174
rect 13227 7125 13269 7134
rect 14275 7160 14333 7161
rect 12739 7119 12797 7120
rect 14275 7120 14284 7160
rect 14324 7120 14333 7160
rect 14275 7119 14333 7120
rect 15523 7160 15581 7161
rect 15523 7120 15532 7160
rect 15572 7120 15581 7160
rect 15523 7119 15581 7120
rect 15915 7160 15957 7169
rect 15915 7120 15916 7160
rect 15956 7120 15957 7160
rect 15915 7111 15957 7120
rect 16011 7160 16053 7169
rect 16011 7120 16012 7160
rect 16052 7120 16053 7160
rect 16011 7111 16053 7120
rect 16387 7160 16445 7161
rect 16387 7120 16396 7160
rect 16436 7120 16445 7160
rect 16387 7119 16445 7120
rect 16675 7160 16733 7161
rect 16675 7120 16684 7160
rect 16724 7120 16733 7160
rect 16675 7119 16733 7120
rect 17923 7160 17981 7161
rect 17923 7120 17932 7160
rect 17972 7120 17981 7160
rect 17923 7119 17981 7120
rect 18307 7160 18365 7161
rect 18307 7120 18316 7160
rect 18356 7120 18365 7160
rect 18307 7119 18365 7120
rect 19555 7160 19613 7161
rect 19555 7120 19564 7160
rect 19604 7120 19613 7160
rect 19555 7119 19613 7120
rect 11403 7076 11445 7085
rect 11403 7036 11404 7076
rect 11444 7036 11445 7076
rect 11403 7027 11445 7036
rect 18123 7076 18165 7085
rect 18123 7036 18124 7076
rect 18164 7036 18165 7076
rect 18123 7027 18165 7036
rect 2667 6992 2709 7001
rect 2667 6952 2668 6992
rect 2708 6952 2709 6992
rect 2667 6943 2709 6952
rect 4771 6992 4829 6993
rect 4771 6952 4780 6992
rect 4820 6952 4829 6992
rect 4771 6951 4829 6952
rect 9771 6992 9813 7001
rect 9771 6952 9772 6992
rect 9812 6952 9813 6992
rect 9771 6943 9813 6952
rect 13419 6992 13461 7001
rect 13419 6952 13420 6992
rect 13460 6952 13461 6992
rect 13419 6943 13461 6952
rect 16195 6992 16253 6993
rect 16195 6952 16204 6992
rect 16244 6952 16253 6992
rect 16195 6951 16253 6952
rect 16491 6992 16533 7001
rect 16491 6952 16492 6992
rect 16532 6952 16533 6992
rect 16491 6943 16533 6952
rect 1152 6824 20452 6848
rect 1152 6784 4928 6824
rect 4968 6784 5010 6824
rect 5050 6784 5092 6824
rect 5132 6784 5174 6824
rect 5214 6784 5256 6824
rect 5296 6784 20048 6824
rect 20088 6784 20130 6824
rect 20170 6784 20212 6824
rect 20252 6784 20294 6824
rect 20334 6784 20376 6824
rect 20416 6784 20452 6824
rect 1152 6760 20452 6784
rect 16683 6714 16725 6723
rect 16683 6674 16684 6714
rect 16724 6674 16725 6714
rect 16683 6665 16725 6674
rect 2667 6656 2709 6665
rect 2667 6616 2668 6656
rect 2708 6616 2709 6656
rect 2667 6607 2709 6616
rect 3235 6656 3293 6657
rect 3235 6616 3244 6656
rect 3284 6616 3293 6656
rect 3235 6615 3293 6616
rect 6891 6656 6933 6665
rect 6891 6616 6892 6656
rect 6932 6616 6933 6656
rect 6891 6607 6933 6616
rect 20043 6656 20085 6665
rect 20043 6616 20044 6656
rect 20084 6616 20085 6656
rect 20043 6607 20085 6616
rect 10443 6572 10485 6581
rect 10443 6532 10444 6572
rect 10484 6532 10485 6572
rect 10443 6523 10485 6532
rect 12651 6572 12693 6581
rect 12651 6532 12652 6572
rect 12692 6532 12693 6572
rect 12651 6523 12693 6532
rect 14667 6572 14709 6581
rect 14667 6532 14668 6572
rect 14708 6532 14709 6572
rect 14667 6523 14709 6532
rect 1219 6488 1277 6489
rect 1219 6448 1228 6488
rect 1268 6448 1277 6488
rect 1219 6447 1277 6448
rect 2467 6488 2525 6489
rect 2467 6448 2476 6488
rect 2516 6448 2525 6488
rect 2467 6447 2525 6448
rect 2955 6488 2997 6497
rect 2955 6448 2956 6488
rect 2996 6448 2997 6488
rect 2955 6439 2997 6448
rect 3051 6488 3093 6497
rect 3051 6448 3052 6488
rect 3092 6448 3093 6488
rect 3051 6439 3093 6448
rect 3147 6488 3189 6497
rect 3147 6448 3148 6488
rect 3188 6448 3189 6488
rect 3147 6439 3189 6448
rect 3427 6488 3485 6489
rect 3427 6448 3436 6488
rect 3476 6448 3485 6488
rect 3427 6447 3485 6448
rect 5163 6488 5205 6497
rect 5163 6448 5164 6488
rect 5204 6448 5205 6488
rect 4675 6446 4733 6447
rect 4675 6406 4684 6446
rect 4724 6406 4733 6446
rect 5163 6439 5205 6448
rect 5259 6488 5301 6497
rect 5259 6448 5260 6488
rect 5300 6448 5301 6488
rect 5259 6439 5301 6448
rect 5643 6488 5685 6497
rect 5643 6448 5644 6488
rect 5684 6448 5685 6488
rect 5643 6439 5685 6448
rect 6211 6488 6269 6489
rect 6211 6448 6220 6488
rect 6260 6448 6269 6488
rect 7075 6488 7133 6489
rect 6211 6447 6269 6448
rect 6699 6474 6741 6483
rect 6699 6434 6700 6474
rect 6740 6434 6741 6474
rect 7075 6448 7084 6488
rect 7124 6448 7133 6488
rect 7075 6447 7133 6448
rect 8715 6488 8757 6497
rect 8715 6448 8716 6488
rect 8756 6448 8757 6488
rect 8715 6439 8757 6448
rect 8811 6488 8853 6497
rect 8811 6448 8812 6488
rect 8852 6448 8853 6488
rect 8811 6439 8853 6448
rect 9195 6488 9237 6497
rect 9195 6448 9196 6488
rect 9236 6448 9237 6488
rect 9195 6439 9237 6448
rect 9291 6488 9333 6497
rect 9291 6448 9292 6488
rect 9332 6448 9333 6488
rect 9291 6439 9333 6448
rect 9763 6488 9821 6489
rect 9763 6448 9772 6488
rect 9812 6448 9821 6488
rect 9763 6447 9821 6448
rect 10251 6483 10293 6492
rect 10251 6443 10252 6483
rect 10292 6443 10293 6483
rect 11203 6488 11261 6489
rect 11203 6448 11212 6488
rect 11252 6448 11261 6488
rect 11203 6447 11261 6448
rect 12451 6488 12509 6489
rect 12451 6448 12460 6488
rect 12500 6448 12509 6488
rect 12451 6447 12509 6448
rect 12939 6488 12981 6497
rect 12939 6448 12940 6488
rect 12980 6448 12981 6488
rect 10251 6434 10293 6443
rect 12939 6439 12981 6448
rect 13035 6488 13077 6497
rect 13035 6448 13036 6488
rect 13076 6448 13077 6488
rect 13035 6439 13077 6448
rect 13419 6488 13461 6497
rect 13419 6448 13420 6488
rect 13460 6448 13461 6488
rect 13419 6439 13461 6448
rect 13987 6488 14045 6489
rect 13987 6448 13996 6488
rect 14036 6448 14045 6488
rect 15723 6488 15765 6497
rect 13987 6447 14045 6448
rect 14523 6446 14565 6455
rect 6699 6425 6741 6434
rect 4675 6405 4733 6406
rect 5739 6404 5781 6413
rect 5739 6364 5740 6404
rect 5780 6364 5781 6404
rect 5739 6355 5781 6364
rect 13515 6404 13557 6413
rect 13515 6364 13516 6404
rect 13556 6364 13557 6404
rect 14523 6406 14524 6446
rect 14564 6406 14565 6446
rect 15723 6448 15724 6488
rect 15764 6448 15765 6488
rect 15723 6439 15765 6448
rect 15915 6488 15957 6497
rect 15915 6448 15916 6488
rect 15956 6448 15957 6488
rect 15915 6439 15957 6448
rect 16003 6488 16061 6489
rect 16003 6448 16012 6488
rect 16052 6448 16061 6488
rect 16003 6447 16061 6448
rect 16491 6488 16533 6497
rect 16491 6448 16492 6488
rect 16532 6448 16533 6488
rect 16491 6439 16533 6448
rect 16579 6488 16637 6489
rect 16579 6448 16588 6488
rect 16628 6448 16637 6488
rect 16579 6447 16637 6448
rect 16875 6488 16917 6497
rect 16875 6448 16876 6488
rect 16916 6448 16917 6488
rect 16875 6439 16917 6448
rect 17067 6488 17109 6497
rect 17067 6448 17068 6488
rect 17108 6448 17109 6488
rect 17067 6439 17109 6448
rect 17155 6488 17213 6489
rect 17155 6448 17164 6488
rect 17204 6448 17213 6488
rect 17155 6447 17213 6448
rect 17643 6488 17685 6497
rect 17643 6448 17644 6488
rect 17684 6448 17685 6488
rect 17643 6439 17685 6448
rect 17739 6488 17781 6497
rect 17739 6448 17740 6488
rect 17780 6448 17781 6488
rect 17739 6439 17781 6448
rect 17835 6488 17877 6497
rect 17835 6448 17836 6488
rect 17876 6448 17877 6488
rect 17835 6439 17877 6448
rect 18315 6488 18357 6497
rect 18315 6448 18316 6488
rect 18356 6448 18357 6488
rect 18315 6439 18357 6448
rect 18411 6488 18453 6497
rect 18411 6448 18412 6488
rect 18452 6448 18453 6488
rect 18411 6439 18453 6448
rect 18891 6488 18933 6497
rect 18891 6448 18892 6488
rect 18932 6448 18933 6488
rect 18891 6439 18933 6448
rect 19363 6488 19421 6489
rect 19363 6448 19372 6488
rect 19412 6448 19421 6488
rect 19363 6447 19421 6448
rect 19851 6483 19893 6492
rect 19851 6443 19852 6483
rect 19892 6443 19893 6483
rect 19851 6434 19893 6443
rect 14523 6397 14565 6406
rect 18795 6404 18837 6413
rect 13515 6355 13557 6364
rect 18795 6364 18796 6404
rect 18836 6364 18837 6404
rect 18795 6355 18837 6364
rect 4875 6320 4917 6329
rect 4875 6280 4876 6320
rect 4916 6280 4917 6320
rect 4875 6271 4917 6280
rect 16875 6320 16917 6329
rect 16875 6280 16876 6320
rect 16916 6280 16917 6320
rect 16875 6271 16917 6280
rect 18019 6320 18077 6321
rect 18019 6280 18028 6320
rect 18068 6280 18077 6320
rect 18019 6279 18077 6280
rect 7179 6236 7221 6245
rect 7179 6196 7180 6236
rect 7220 6196 7221 6236
rect 7179 6187 7221 6196
rect 15723 6236 15765 6245
rect 15723 6196 15724 6236
rect 15764 6196 15765 6236
rect 15723 6187 15765 6196
rect 16203 6236 16245 6245
rect 16203 6196 16204 6236
rect 16244 6196 16245 6236
rect 16203 6187 16245 6196
rect 1152 6068 20352 6092
rect 1152 6028 3688 6068
rect 3728 6028 3770 6068
rect 3810 6028 3852 6068
rect 3892 6028 3934 6068
rect 3974 6028 4016 6068
rect 4056 6028 18808 6068
rect 18848 6028 18890 6068
rect 18930 6028 18972 6068
rect 19012 6028 19054 6068
rect 19094 6028 19136 6068
rect 19176 6028 20352 6068
rect 1152 6004 20352 6028
rect 1507 5900 1565 5901
rect 1507 5860 1516 5900
rect 1556 5860 1565 5900
rect 1507 5859 1565 5860
rect 4963 5900 5021 5901
rect 4963 5860 4972 5900
rect 5012 5860 5021 5900
rect 4963 5859 5021 5860
rect 6603 5900 6645 5909
rect 6603 5860 6604 5900
rect 6644 5860 6645 5900
rect 6603 5851 6645 5860
rect 8427 5900 8469 5909
rect 8427 5860 8428 5900
rect 8468 5860 8469 5900
rect 8427 5851 8469 5860
rect 14667 5900 14709 5909
rect 14667 5860 14668 5900
rect 14708 5860 14709 5900
rect 14667 5851 14709 5860
rect 19755 5900 19797 5909
rect 19755 5860 19756 5900
rect 19796 5860 19797 5900
rect 19755 5851 19797 5860
rect 15627 5816 15669 5825
rect 15627 5776 15628 5816
rect 15668 5776 15669 5816
rect 15627 5767 15669 5776
rect 16003 5816 16061 5817
rect 16003 5776 16012 5816
rect 16052 5776 16061 5816
rect 16003 5775 16061 5776
rect 16971 5816 17013 5825
rect 16971 5776 16972 5816
rect 17012 5776 17013 5816
rect 16971 5767 17013 5776
rect 3627 5732 3669 5741
rect 3627 5692 3628 5732
rect 3668 5692 3669 5732
rect 3627 5683 3669 5692
rect 3723 5732 3765 5741
rect 3723 5692 3724 5732
rect 3764 5692 3765 5732
rect 3723 5683 3765 5692
rect 9195 5732 9237 5741
rect 9195 5692 9196 5732
rect 9236 5692 9237 5732
rect 9195 5683 9237 5692
rect 9291 5732 9333 5741
rect 9291 5692 9292 5732
rect 9332 5692 9333 5732
rect 9291 5683 9333 5692
rect 15531 5732 15573 5741
rect 15531 5692 15532 5732
rect 15572 5692 15573 5732
rect 15531 5683 15573 5692
rect 15723 5732 15765 5741
rect 15723 5692 15724 5732
rect 15764 5692 15765 5732
rect 17931 5693 17973 5702
rect 15723 5683 15765 5692
rect 17347 5691 17405 5692
rect 10251 5662 10293 5671
rect 1803 5648 1845 5657
rect 1803 5608 1804 5648
rect 1844 5608 1845 5648
rect 1803 5599 1845 5608
rect 1899 5648 1941 5657
rect 2667 5653 2709 5662
rect 1899 5608 1900 5648
rect 1940 5608 1941 5648
rect 1899 5599 1941 5608
rect 2179 5648 2237 5649
rect 2179 5608 2188 5648
rect 2228 5608 2237 5648
rect 2179 5607 2237 5608
rect 2667 5613 2668 5653
rect 2708 5613 2709 5653
rect 2667 5604 2709 5613
rect 3139 5648 3197 5649
rect 3139 5608 3148 5648
rect 3188 5608 3197 5648
rect 3139 5607 3197 5608
rect 4107 5648 4149 5657
rect 4107 5608 4108 5648
rect 4148 5608 4149 5648
rect 4107 5599 4149 5608
rect 4203 5648 4245 5657
rect 4203 5608 4204 5648
rect 4244 5608 4245 5648
rect 4203 5599 4245 5608
rect 4587 5648 4629 5657
rect 4587 5608 4588 5648
rect 4628 5608 4629 5648
rect 4587 5599 4629 5608
rect 4683 5648 4725 5657
rect 4683 5608 4684 5648
rect 4724 5608 4725 5648
rect 4683 5599 4725 5608
rect 4779 5648 4821 5657
rect 4779 5608 4780 5648
rect 4820 5608 4821 5648
rect 4779 5599 4821 5608
rect 5155 5648 5213 5649
rect 5155 5608 5164 5648
rect 5204 5608 5213 5648
rect 5155 5607 5213 5608
rect 6403 5648 6461 5649
rect 6403 5608 6412 5648
rect 6452 5608 6461 5648
rect 6403 5607 6461 5608
rect 6979 5648 7037 5649
rect 6979 5608 6988 5648
rect 7028 5608 7037 5648
rect 6979 5607 7037 5608
rect 8227 5648 8285 5649
rect 8227 5608 8236 5648
rect 8276 5608 8285 5648
rect 8227 5607 8285 5608
rect 8715 5648 8757 5657
rect 8715 5608 8716 5648
rect 8756 5608 8757 5648
rect 8715 5599 8757 5608
rect 8811 5648 8853 5657
rect 8811 5608 8812 5648
rect 8852 5608 8853 5648
rect 8811 5599 8853 5608
rect 9763 5648 9821 5649
rect 9763 5608 9772 5648
rect 9812 5608 9821 5648
rect 10251 5622 10252 5662
rect 10292 5622 10293 5662
rect 10251 5613 10293 5622
rect 11395 5648 11453 5649
rect 9763 5607 9821 5608
rect 11395 5608 11404 5648
rect 11444 5608 11453 5648
rect 11395 5607 11453 5608
rect 12643 5648 12701 5649
rect 12643 5608 12652 5648
rect 12692 5608 12701 5648
rect 12643 5607 12701 5608
rect 13219 5648 13277 5649
rect 13219 5608 13228 5648
rect 13268 5608 13277 5648
rect 13219 5607 13277 5608
rect 14467 5648 14525 5649
rect 14467 5608 14476 5648
rect 14516 5608 14525 5648
rect 14467 5607 14525 5608
rect 14955 5648 14997 5657
rect 14955 5608 14956 5648
rect 14996 5608 14997 5648
rect 14955 5599 14997 5608
rect 15051 5648 15093 5657
rect 15051 5608 15052 5648
rect 15092 5608 15093 5648
rect 15051 5599 15093 5608
rect 15147 5648 15189 5657
rect 15147 5608 15148 5648
rect 15188 5608 15189 5648
rect 15147 5599 15189 5608
rect 15243 5648 15285 5657
rect 15243 5608 15244 5648
rect 15284 5608 15285 5648
rect 15243 5599 15285 5608
rect 15427 5648 15485 5649
rect 15427 5608 15436 5648
rect 15476 5608 15485 5648
rect 15427 5607 15485 5608
rect 15819 5648 15861 5657
rect 15819 5608 15820 5648
rect 15860 5608 15861 5648
rect 15819 5599 15861 5608
rect 16395 5648 16437 5657
rect 16395 5608 16396 5648
rect 16436 5608 16437 5648
rect 16395 5599 16437 5608
rect 16675 5648 16733 5649
rect 16675 5608 16684 5648
rect 16724 5608 16733 5648
rect 16675 5607 16733 5608
rect 17259 5648 17301 5657
rect 17347 5651 17356 5691
rect 17396 5651 17405 5691
rect 17347 5650 17405 5651
rect 17259 5608 17260 5648
rect 17300 5608 17301 5648
rect 17259 5599 17301 5608
rect 17643 5648 17685 5657
rect 17643 5608 17644 5648
rect 17684 5608 17685 5648
rect 17643 5599 17685 5608
rect 17739 5656 17781 5665
rect 17739 5616 17740 5656
rect 17780 5616 17781 5656
rect 17739 5607 17781 5616
rect 17835 5648 17877 5657
rect 17835 5608 17836 5648
rect 17876 5608 17877 5648
rect 17931 5653 17932 5693
rect 17972 5653 17973 5693
rect 20131 5690 20189 5691
rect 17931 5644 17973 5653
rect 18307 5648 18365 5649
rect 17835 5599 17877 5608
rect 18307 5608 18316 5648
rect 18356 5608 18365 5648
rect 18307 5607 18365 5608
rect 19555 5648 19613 5649
rect 19555 5608 19564 5648
rect 19604 5608 19613 5648
rect 19555 5607 19613 5608
rect 19947 5648 19989 5657
rect 19947 5608 19948 5648
rect 19988 5608 19989 5648
rect 19947 5599 19989 5608
rect 20043 5648 20085 5657
rect 20131 5650 20140 5690
rect 20180 5650 20189 5690
rect 20131 5649 20189 5650
rect 20043 5608 20044 5648
rect 20084 5608 20085 5648
rect 20043 5599 20085 5608
rect 20235 5648 20277 5657
rect 20235 5608 20236 5648
rect 20276 5608 20277 5648
rect 20235 5599 20277 5608
rect 16299 5564 16341 5573
rect 16299 5524 16300 5564
rect 16340 5524 16341 5564
rect 16299 5515 16341 5524
rect 2475 5480 2517 5489
rect 2475 5440 2476 5480
rect 2516 5440 2517 5480
rect 2475 5431 2517 5440
rect 10443 5480 10485 5489
rect 10443 5440 10444 5480
rect 10484 5440 10485 5480
rect 10443 5431 10485 5440
rect 12843 5480 12885 5489
rect 12843 5440 12844 5480
rect 12884 5440 12885 5480
rect 12843 5431 12885 5440
rect 17451 5422 17493 5431
rect 17451 5382 17452 5422
rect 17492 5382 17493 5422
rect 17451 5373 17493 5382
rect 1152 5312 20452 5336
rect 1152 5272 4928 5312
rect 4968 5272 5010 5312
rect 5050 5272 5092 5312
rect 5132 5272 5174 5312
rect 5214 5272 5256 5312
rect 5296 5272 20048 5312
rect 20088 5272 20130 5312
rect 20170 5272 20212 5312
rect 20252 5272 20294 5312
rect 20334 5272 20376 5312
rect 20416 5272 20452 5312
rect 1152 5248 20452 5272
rect 8811 5060 8853 5069
rect 8811 5020 8812 5060
rect 8852 5020 8853 5060
rect 8811 5011 8853 5020
rect 12843 5060 12885 5069
rect 12843 5020 12844 5060
rect 12884 5020 12885 5060
rect 12843 5011 12885 5020
rect 14859 5060 14901 5069
rect 14859 5020 14860 5060
rect 14900 5020 14901 5060
rect 14859 5011 14901 5020
rect 16491 5060 16533 5069
rect 16491 5020 16492 5060
rect 16532 5020 16533 5060
rect 16491 5011 16533 5020
rect 18411 5018 18453 5027
rect 13131 4996 13173 5005
rect 1219 4976 1277 4977
rect 1219 4936 1228 4976
rect 1268 4936 1277 4976
rect 1219 4935 1277 4936
rect 2467 4976 2525 4977
rect 2467 4936 2476 4976
rect 2516 4936 2525 4976
rect 2467 4935 2525 4936
rect 2851 4976 2909 4977
rect 2851 4936 2860 4976
rect 2900 4936 2909 4976
rect 2851 4935 2909 4936
rect 4099 4976 4157 4977
rect 4099 4936 4108 4976
rect 4148 4936 4157 4976
rect 4099 4935 4157 4936
rect 4491 4976 4533 4985
rect 4491 4936 4492 4976
rect 4532 4936 4533 4976
rect 4491 4927 4533 4936
rect 4779 4976 4821 4985
rect 4779 4936 4780 4976
rect 4820 4936 4821 4976
rect 4779 4927 4821 4936
rect 5251 4976 5309 4977
rect 5251 4936 5260 4976
rect 5300 4936 5309 4976
rect 5251 4935 5309 4936
rect 6499 4976 6557 4977
rect 6499 4936 6508 4976
rect 6548 4936 6557 4976
rect 6499 4935 6557 4936
rect 7083 4976 7125 4985
rect 7083 4936 7084 4976
rect 7124 4936 7125 4976
rect 7083 4927 7125 4936
rect 7179 4976 7221 4985
rect 7179 4936 7180 4976
rect 7220 4936 7221 4976
rect 7179 4927 7221 4936
rect 8131 4976 8189 4977
rect 8131 4936 8140 4976
rect 8180 4936 8189 4976
rect 9763 4976 9821 4977
rect 8131 4935 8189 4936
rect 8619 4962 8661 4971
rect 8619 4922 8620 4962
rect 8660 4922 8661 4962
rect 9763 4936 9772 4976
rect 9812 4936 9821 4976
rect 9763 4935 9821 4936
rect 11011 4976 11069 4977
rect 11011 4936 11020 4976
rect 11060 4936 11069 4976
rect 11011 4935 11069 4936
rect 11395 4976 11453 4977
rect 11395 4936 11404 4976
rect 11444 4936 11453 4976
rect 11395 4935 11453 4936
rect 12643 4976 12701 4977
rect 12643 4936 12652 4976
rect 12692 4936 12701 4976
rect 13131 4956 13132 4996
rect 13172 4956 13173 4996
rect 13131 4947 13173 4956
rect 13227 4976 13269 4985
rect 12643 4935 12701 4936
rect 13227 4936 13228 4976
rect 13268 4936 13269 4976
rect 13227 4927 13269 4936
rect 13611 4976 13653 4985
rect 13611 4936 13612 4976
rect 13652 4936 13653 4976
rect 13611 4927 13653 4936
rect 13707 4976 13749 4985
rect 13707 4936 13708 4976
rect 13748 4936 13749 4976
rect 13707 4927 13749 4936
rect 14179 4976 14237 4977
rect 14179 4936 14188 4976
rect 14228 4936 14237 4976
rect 15043 4976 15101 4977
rect 14179 4935 14237 4936
rect 14667 4962 14709 4971
rect 8619 4913 8661 4922
rect 14667 4922 14668 4962
rect 14708 4922 14709 4962
rect 15043 4936 15052 4976
rect 15092 4936 15101 4976
rect 15043 4935 15101 4936
rect 16291 4976 16349 4977
rect 16291 4936 16300 4976
rect 16340 4936 16349 4976
rect 16291 4935 16349 4936
rect 16771 4976 16829 4977
rect 16771 4936 16780 4976
rect 16820 4936 16829 4976
rect 16771 4935 16829 4936
rect 17067 4976 17109 4985
rect 18411 4978 18412 5018
rect 18452 4978 18453 5018
rect 17067 4936 17068 4976
rect 17108 4936 17109 4976
rect 17067 4927 17109 4936
rect 17731 4976 17789 4977
rect 17731 4936 17740 4976
rect 17780 4936 17789 4976
rect 17731 4935 17789 4936
rect 18307 4976 18365 4977
rect 18307 4936 18316 4976
rect 18356 4936 18365 4976
rect 18411 4969 18453 4978
rect 18603 4976 18645 4985
rect 18307 4935 18365 4936
rect 18603 4936 18604 4976
rect 18644 4936 18645 4976
rect 17155 4934 17213 4935
rect 14667 4913 14709 4922
rect 7563 4892 7605 4901
rect 7563 4852 7564 4892
rect 7604 4852 7605 4892
rect 7563 4843 7605 4852
rect 7659 4892 7701 4901
rect 17155 4894 17164 4934
rect 17204 4894 17213 4934
rect 18603 4927 18645 4936
rect 19371 4976 19413 4985
rect 19371 4936 19372 4976
rect 19412 4936 19413 4976
rect 19371 4927 19413 4936
rect 19467 4976 19509 4985
rect 19467 4936 19468 4976
rect 19508 4936 19509 4976
rect 19467 4927 19509 4936
rect 19747 4976 19805 4977
rect 19747 4936 19756 4976
rect 19796 4936 19805 4976
rect 19747 4935 19805 4936
rect 17155 4893 17213 4894
rect 7659 4852 7660 4892
rect 7700 4852 7701 4892
rect 7659 4843 7701 4852
rect 2667 4808 2709 4817
rect 2667 4768 2668 4808
rect 2708 4768 2709 4808
rect 2667 4759 2709 4768
rect 17443 4808 17501 4809
rect 17443 4768 17452 4808
rect 17492 4768 17501 4808
rect 17443 4767 17501 4768
rect 19075 4808 19133 4809
rect 19075 4768 19084 4808
rect 19124 4768 19133 4808
rect 19075 4767 19133 4768
rect 4299 4724 4341 4733
rect 4299 4684 4300 4724
rect 4340 4684 4341 4724
rect 4299 4675 4341 4684
rect 4491 4724 4533 4733
rect 4491 4684 4492 4724
rect 4532 4684 4533 4724
rect 4491 4675 4533 4684
rect 6699 4724 6741 4733
rect 6699 4684 6700 4724
rect 6740 4684 6741 4724
rect 6699 4675 6741 4684
rect 11211 4724 11253 4733
rect 11211 4684 11212 4724
rect 11252 4684 11253 4724
rect 11211 4675 11253 4684
rect 17643 4724 17685 4733
rect 17643 4684 17644 4724
rect 17684 4684 17685 4724
rect 17643 4675 17685 4684
rect 18603 4724 18645 4733
rect 18603 4684 18604 4724
rect 18644 4684 18645 4724
rect 18603 4675 18645 4684
rect 1152 4556 20352 4580
rect 1152 4516 3688 4556
rect 3728 4516 3770 4556
rect 3810 4516 3852 4556
rect 3892 4516 3934 4556
rect 3974 4516 4016 4556
rect 4056 4516 18808 4556
rect 18848 4516 18890 4556
rect 18930 4516 18972 4556
rect 19012 4516 19054 4556
rect 19094 4516 19136 4556
rect 19176 4516 20352 4556
rect 1152 4492 20352 4516
rect 3147 4388 3189 4397
rect 3147 4348 3148 4388
rect 3188 4348 3189 4388
rect 3147 4339 3189 4348
rect 8715 4388 8757 4397
rect 8715 4348 8716 4388
rect 8756 4348 8757 4388
rect 8715 4339 8757 4348
rect 14763 4388 14805 4397
rect 14763 4348 14764 4388
rect 14804 4348 14805 4388
rect 14763 4339 14805 4348
rect 16299 4388 16341 4397
rect 16299 4348 16300 4388
rect 16340 4348 16341 4388
rect 16299 4339 16341 4348
rect 16587 4388 16629 4397
rect 16587 4348 16588 4388
rect 16628 4348 16629 4388
rect 16587 4339 16629 4348
rect 4971 4304 5013 4313
rect 4971 4264 4972 4304
rect 5012 4264 5013 4304
rect 4971 4255 5013 4264
rect 17635 4304 17693 4305
rect 17635 4264 17644 4304
rect 17684 4264 17693 4304
rect 17635 4263 17693 4264
rect 5835 4220 5877 4229
rect 5835 4180 5836 4220
rect 5876 4180 5877 4220
rect 5835 4171 5877 4180
rect 11883 4220 11925 4229
rect 11883 4180 11884 4220
rect 11924 4180 11925 4220
rect 11883 4171 11925 4180
rect 18987 4220 19029 4229
rect 18987 4180 18988 4220
rect 19028 4180 19029 4220
rect 18987 4171 19029 4180
rect 19083 4220 19125 4229
rect 19083 4180 19084 4220
rect 19124 4180 19125 4220
rect 19083 4171 19125 4180
rect 12939 4150 12981 4159
rect 1219 4136 1277 4137
rect 1219 4096 1228 4136
rect 1268 4096 1277 4136
rect 1219 4095 1277 4096
rect 2467 4136 2525 4137
rect 2467 4096 2476 4136
rect 2516 4096 2525 4136
rect 2467 4095 2525 4096
rect 2851 4136 2909 4137
rect 2851 4096 2860 4136
rect 2900 4096 2909 4136
rect 2851 4095 2909 4096
rect 2955 4136 2997 4145
rect 2955 4096 2956 4136
rect 2996 4096 2997 4136
rect 2955 4087 2997 4096
rect 3147 4136 3189 4145
rect 3147 4096 3148 4136
rect 3188 4096 3189 4136
rect 3147 4087 3189 4096
rect 3331 4136 3389 4137
rect 3331 4096 3340 4136
rect 3380 4096 3389 4136
rect 3331 4095 3389 4096
rect 4579 4136 4637 4137
rect 4579 4096 4588 4136
rect 4628 4096 4637 4136
rect 4579 4095 4637 4096
rect 5355 4136 5397 4145
rect 5355 4096 5356 4136
rect 5396 4096 5397 4136
rect 5355 4087 5397 4096
rect 5451 4136 5493 4145
rect 5451 4096 5452 4136
rect 5492 4096 5493 4136
rect 5451 4087 5493 4096
rect 5931 4136 5973 4145
rect 6891 4141 6933 4150
rect 5931 4096 5932 4136
rect 5972 4096 5973 4136
rect 5931 4087 5973 4096
rect 6403 4136 6461 4137
rect 6403 4096 6412 4136
rect 6452 4096 6461 4136
rect 6403 4095 6461 4096
rect 6891 4101 6892 4141
rect 6932 4101 6933 4141
rect 6891 4092 6933 4101
rect 7267 4136 7325 4137
rect 7267 4096 7276 4136
rect 7316 4096 7325 4136
rect 7267 4095 7325 4096
rect 8515 4136 8573 4137
rect 8515 4096 8524 4136
rect 8564 4096 8573 4136
rect 8515 4095 8573 4096
rect 8995 4136 9053 4137
rect 8995 4096 9004 4136
rect 9044 4096 9053 4136
rect 8995 4095 9053 4096
rect 10243 4136 10301 4137
rect 10243 4096 10252 4136
rect 10292 4096 10301 4136
rect 10243 4095 10301 4096
rect 11403 4136 11445 4145
rect 11403 4096 11404 4136
rect 11444 4096 11445 4136
rect 11403 4087 11445 4096
rect 11499 4136 11541 4145
rect 11499 4096 11500 4136
rect 11540 4096 11541 4136
rect 11499 4087 11541 4096
rect 11979 4136 12021 4145
rect 11979 4096 11980 4136
rect 12020 4096 12021 4136
rect 11979 4087 12021 4096
rect 12450 4127 12508 4128
rect 12450 4087 12459 4127
rect 12499 4087 12508 4127
rect 12939 4110 12940 4150
rect 12980 4110 12981 4150
rect 12939 4101 12981 4110
rect 13315 4136 13373 4137
rect 13315 4096 13324 4136
rect 13364 4096 13373 4136
rect 13315 4095 13373 4096
rect 14563 4136 14621 4137
rect 14563 4096 14572 4136
rect 14612 4096 14621 4136
rect 14563 4095 14621 4096
rect 16387 4136 16445 4137
rect 16387 4096 16396 4136
rect 16436 4096 16445 4136
rect 16387 4095 16445 4096
rect 16675 4136 16733 4137
rect 16675 4096 16684 4136
rect 16724 4096 16733 4136
rect 16675 4095 16733 4096
rect 16963 4136 17021 4137
rect 16963 4096 16972 4136
rect 17012 4096 17021 4136
rect 16963 4095 17021 4096
rect 17259 4136 17301 4145
rect 17259 4096 17260 4136
rect 17300 4096 17301 4136
rect 17259 4087 17301 4096
rect 17355 4136 17397 4145
rect 17355 4096 17356 4136
rect 17396 4096 17397 4136
rect 17355 4087 17397 4096
rect 18507 4136 18549 4145
rect 18507 4096 18508 4136
rect 18548 4096 18549 4136
rect 18507 4087 18549 4096
rect 18603 4136 18645 4145
rect 20043 4141 20085 4150
rect 18603 4096 18604 4136
rect 18644 4096 18645 4136
rect 18603 4087 18645 4096
rect 19555 4136 19613 4137
rect 19555 4096 19564 4136
rect 19604 4096 19613 4136
rect 19555 4095 19613 4096
rect 20043 4101 20044 4141
rect 20084 4101 20085 4141
rect 20043 4092 20085 4101
rect 12450 4086 12508 4087
rect 4779 4052 4821 4061
rect 4779 4012 4780 4052
rect 4820 4012 4821 4052
rect 4779 4003 4821 4012
rect 7083 4052 7125 4061
rect 7083 4012 7084 4052
rect 7124 4012 7125 4052
rect 7083 4003 7125 4012
rect 20235 4052 20277 4061
rect 20235 4012 20236 4052
rect 20276 4012 20277 4052
rect 20235 4003 20277 4012
rect 2667 3968 2709 3977
rect 2667 3928 2668 3968
rect 2708 3928 2709 3968
rect 2667 3919 2709 3928
rect 10443 3968 10485 3977
rect 10443 3928 10444 3968
rect 10484 3928 10485 3968
rect 10443 3919 10485 3928
rect 13131 3968 13173 3977
rect 13131 3928 13132 3968
rect 13172 3928 13173 3968
rect 13131 3919 13173 3928
rect 1152 3800 20452 3824
rect 1152 3760 4928 3800
rect 4968 3760 5010 3800
rect 5050 3760 5092 3800
rect 5132 3760 5174 3800
rect 5214 3760 5256 3800
rect 5296 3760 20048 3800
rect 20088 3760 20130 3800
rect 20170 3760 20212 3800
rect 20252 3760 20294 3800
rect 20334 3760 20376 3800
rect 20416 3760 20452 3800
rect 1152 3736 20452 3760
rect 17259 3690 17301 3699
rect 17259 3650 17260 3690
rect 17300 3650 17301 3690
rect 5067 3636 5109 3645
rect 17259 3641 17301 3650
rect 5067 3596 5068 3636
rect 5108 3596 5109 3636
rect 5067 3587 5109 3596
rect 6699 3632 6741 3641
rect 6699 3592 6700 3632
rect 6740 3592 6741 3632
rect 6699 3583 6741 3592
rect 7075 3632 7133 3633
rect 7075 3592 7084 3632
rect 7124 3592 7133 3632
rect 15627 3632 15669 3641
rect 7075 3591 7133 3592
rect 8235 3590 8277 3599
rect 2475 3548 2517 3557
rect 2475 3508 2476 3548
rect 2516 3508 2517 3548
rect 8235 3550 8236 3590
rect 8276 3550 8277 3590
rect 15627 3592 15628 3632
rect 15668 3592 15669 3632
rect 15627 3583 15669 3592
rect 17443 3632 17501 3633
rect 17443 3592 17452 3632
rect 17492 3592 17501 3632
rect 17443 3591 17501 3592
rect 19563 3632 19605 3641
rect 19563 3592 19564 3632
rect 19604 3592 19605 3632
rect 19563 3583 19605 3592
rect 8235 3541 8277 3550
rect 2475 3499 2517 3508
rect 16195 3506 16253 3507
rect 3139 3464 3197 3465
rect 2667 3450 2709 3459
rect 2667 3410 2668 3450
rect 2708 3410 2709 3450
rect 3139 3424 3148 3464
rect 3188 3424 3197 3464
rect 3139 3423 3197 3424
rect 3627 3464 3669 3473
rect 3627 3424 3628 3464
rect 3668 3424 3669 3464
rect 3627 3415 3669 3424
rect 4107 3464 4149 3473
rect 4107 3424 4108 3464
rect 4148 3424 4149 3464
rect 4107 3415 4149 3424
rect 4203 3464 4245 3473
rect 4203 3424 4204 3464
rect 4244 3424 4245 3464
rect 4203 3415 4245 3424
rect 4875 3464 4917 3473
rect 4875 3424 4876 3464
rect 4916 3424 4917 3464
rect 4875 3415 4917 3424
rect 4963 3464 5021 3465
rect 4963 3424 4972 3464
rect 5012 3424 5021 3464
rect 4963 3423 5021 3424
rect 5251 3464 5309 3465
rect 5251 3424 5260 3464
rect 5300 3424 5309 3464
rect 5251 3423 5309 3424
rect 6499 3464 6557 3465
rect 6499 3424 6508 3464
rect 6548 3424 6557 3464
rect 6499 3423 6557 3424
rect 6987 3464 7029 3473
rect 6987 3424 6988 3464
rect 7028 3424 7029 3464
rect 6987 3415 7029 3424
rect 7179 3464 7221 3473
rect 7179 3424 7180 3464
rect 7220 3424 7221 3464
rect 7467 3464 7509 3473
rect 7179 3415 7221 3424
rect 7267 3445 7325 3446
rect 2667 3401 2709 3410
rect 7267 3405 7276 3445
rect 7316 3405 7325 3445
rect 7467 3424 7468 3464
rect 7508 3424 7509 3464
rect 7467 3415 7509 3424
rect 7843 3464 7901 3465
rect 7843 3424 7852 3464
rect 7892 3424 7901 3464
rect 7843 3423 7901 3424
rect 8035 3464 8093 3465
rect 8035 3424 8044 3464
rect 8084 3424 8093 3464
rect 8035 3423 8093 3424
rect 8427 3464 8469 3473
rect 8427 3424 8428 3464
rect 8468 3424 8469 3464
rect 8427 3415 8469 3424
rect 8611 3464 8669 3465
rect 8611 3424 8620 3464
rect 8660 3424 8669 3464
rect 8611 3423 8669 3424
rect 9003 3464 9045 3473
rect 16195 3466 16204 3506
rect 16244 3466 16253 3506
rect 16195 3465 16253 3466
rect 9003 3424 9004 3464
rect 9044 3424 9045 3464
rect 9003 3415 9045 3424
rect 9187 3464 9245 3465
rect 9187 3424 9196 3464
rect 9236 3424 9245 3464
rect 9187 3423 9245 3424
rect 10435 3464 10493 3465
rect 10435 3424 10444 3464
rect 10484 3424 10493 3464
rect 10435 3423 10493 3424
rect 11203 3464 11261 3465
rect 11203 3424 11212 3464
rect 11252 3424 11261 3464
rect 11203 3423 11261 3424
rect 12451 3464 12509 3465
rect 12451 3424 12460 3464
rect 12500 3424 12509 3464
rect 12451 3423 12509 3424
rect 14179 3464 14237 3465
rect 14179 3424 14188 3464
rect 14228 3424 14237 3464
rect 14179 3423 14237 3424
rect 15427 3464 15485 3465
rect 15427 3424 15436 3464
rect 15476 3424 15485 3464
rect 15427 3423 15485 3424
rect 16587 3464 16629 3473
rect 16587 3424 16588 3464
rect 16628 3424 16629 3464
rect 16587 3415 16629 3424
rect 17067 3464 17109 3473
rect 17067 3424 17068 3464
rect 17108 3424 17109 3464
rect 17067 3415 17109 3424
rect 17547 3464 17589 3473
rect 17547 3424 17548 3464
rect 17588 3424 17589 3464
rect 17155 3422 17213 3423
rect 7267 3404 7325 3405
rect 3723 3380 3765 3389
rect 3723 3340 3724 3380
rect 3764 3340 3765 3380
rect 3723 3331 3765 3340
rect 7563 3380 7605 3389
rect 7563 3340 7564 3380
rect 7604 3340 7605 3380
rect 7563 3331 7605 3340
rect 7755 3380 7797 3389
rect 7755 3340 7756 3380
rect 7796 3340 7797 3380
rect 7755 3331 7797 3340
rect 8139 3380 8181 3389
rect 8139 3340 8140 3380
rect 8180 3340 8181 3380
rect 8139 3331 8181 3340
rect 8331 3380 8373 3389
rect 8331 3340 8332 3380
rect 8372 3340 8373 3380
rect 8331 3331 8373 3340
rect 8715 3380 8757 3389
rect 8715 3340 8716 3380
rect 8756 3340 8757 3380
rect 8715 3331 8757 3340
rect 8907 3380 8949 3389
rect 8907 3340 8908 3380
rect 8948 3340 8949 3380
rect 8907 3331 8949 3340
rect 16003 3380 16061 3381
rect 16003 3340 16012 3380
rect 16052 3340 16061 3380
rect 16003 3339 16061 3340
rect 16299 3380 16341 3389
rect 16299 3340 16300 3380
rect 16340 3340 16341 3380
rect 16299 3331 16341 3340
rect 16491 3380 16533 3389
rect 17155 3382 17164 3422
rect 17204 3382 17213 3422
rect 17547 3415 17589 3424
rect 17643 3464 17685 3473
rect 17643 3424 17644 3464
rect 17684 3424 17685 3464
rect 17643 3415 17685 3424
rect 17739 3464 17781 3473
rect 17739 3424 17740 3464
rect 17780 3424 17781 3464
rect 17739 3415 17781 3424
rect 18115 3464 18173 3465
rect 18115 3424 18124 3464
rect 18164 3424 18173 3464
rect 18115 3423 18173 3424
rect 19363 3464 19421 3465
rect 19363 3424 19372 3464
rect 19412 3424 19421 3464
rect 19363 3423 19421 3424
rect 19755 3464 19797 3473
rect 19755 3424 19756 3464
rect 19796 3424 19797 3464
rect 19755 3415 19797 3424
rect 20043 3464 20085 3473
rect 20043 3424 20044 3464
rect 20084 3424 20085 3464
rect 20043 3415 20085 3424
rect 17155 3381 17213 3382
rect 16491 3340 16492 3380
rect 16532 3340 16533 3380
rect 16491 3331 16533 3340
rect 19947 3380 19989 3389
rect 19947 3340 19948 3380
rect 19988 3340 19989 3380
rect 19947 3331 19989 3340
rect 4587 3296 4629 3305
rect 4587 3256 4588 3296
rect 4628 3256 4629 3296
rect 4587 3247 4629 3256
rect 7659 3296 7701 3305
rect 7659 3256 7660 3296
rect 7700 3256 7701 3296
rect 7659 3247 7701 3256
rect 8811 3296 8853 3305
rect 8811 3256 8812 3296
rect 8852 3256 8853 3296
rect 8811 3247 8853 3256
rect 16395 3296 16437 3305
rect 16395 3256 16396 3296
rect 16436 3256 16437 3296
rect 16395 3247 16437 3256
rect 16779 3296 16821 3305
rect 16779 3256 16780 3296
rect 16820 3256 16821 3296
rect 16779 3247 16821 3256
rect 10635 3212 10677 3221
rect 10635 3172 10636 3212
rect 10676 3172 10677 3212
rect 10635 3163 10677 3172
rect 12651 3212 12693 3221
rect 12651 3172 12652 3212
rect 12692 3172 12693 3212
rect 12651 3163 12693 3172
rect 15819 3212 15861 3221
rect 15819 3172 15820 3212
rect 15860 3172 15861 3212
rect 15819 3163 15861 3172
rect 1152 3044 20352 3068
rect 1152 3004 3688 3044
rect 3728 3004 3770 3044
rect 3810 3004 3852 3044
rect 3892 3004 3934 3044
rect 3974 3004 4016 3044
rect 4056 3004 18808 3044
rect 18848 3004 18890 3044
rect 18930 3004 18972 3044
rect 19012 3004 19054 3044
rect 19094 3004 19136 3044
rect 19176 3004 20352 3044
rect 1152 2980 20352 3004
rect 3435 2876 3477 2885
rect 3435 2836 3436 2876
rect 3476 2836 3477 2876
rect 3435 2827 3477 2836
rect 5259 2876 5301 2885
rect 5259 2836 5260 2876
rect 5300 2836 5301 2876
rect 5259 2827 5301 2836
rect 8715 2876 8757 2885
rect 8715 2836 8716 2876
rect 8756 2836 8757 2876
rect 8715 2827 8757 2836
rect 9483 2876 9525 2885
rect 9483 2836 9484 2876
rect 9524 2836 9525 2876
rect 9483 2827 9525 2836
rect 16203 2876 16245 2885
rect 16203 2836 16204 2876
rect 16244 2836 16245 2876
rect 16203 2827 16245 2836
rect 18123 2876 18165 2885
rect 18123 2836 18124 2876
rect 18164 2836 18165 2876
rect 18123 2827 18165 2836
rect 5827 2792 5885 2793
rect 5827 2752 5836 2792
rect 5876 2752 5885 2792
rect 5827 2751 5885 2752
rect 7651 2792 7709 2793
rect 7651 2752 7660 2792
rect 7700 2752 7709 2792
rect 7651 2751 7709 2752
rect 9291 2792 9333 2801
rect 9291 2752 9292 2792
rect 9332 2752 9333 2792
rect 9291 2743 9333 2752
rect 10627 2792 10685 2793
rect 10627 2752 10636 2792
rect 10676 2752 10685 2792
rect 10627 2751 10685 2752
rect 17635 2792 17693 2793
rect 17635 2752 17644 2792
rect 17684 2752 17693 2792
rect 17635 2751 17693 2752
rect 18979 2792 19037 2793
rect 18979 2752 18988 2792
rect 19028 2752 19037 2792
rect 18979 2751 19037 2752
rect 5443 2708 5501 2709
rect 5443 2668 5452 2708
rect 5492 2668 5501 2708
rect 5443 2667 5501 2668
rect 11403 2708 11445 2717
rect 11403 2668 11404 2708
rect 11444 2668 11445 2708
rect 11403 2659 11445 2668
rect 11499 2708 11541 2717
rect 11499 2668 11500 2708
rect 11540 2668 11541 2708
rect 13987 2708 14045 2709
rect 11499 2659 11541 2668
rect 12507 2666 12549 2675
rect 13987 2668 13996 2708
rect 14036 2668 14045 2708
rect 13987 2667 14045 2668
rect 14179 2708 14237 2709
rect 14179 2668 14188 2708
rect 14228 2668 14237 2708
rect 14179 2667 14237 2668
rect 1611 2624 1653 2633
rect 1611 2584 1612 2624
rect 1652 2584 1653 2624
rect 1611 2575 1653 2584
rect 1795 2624 1853 2625
rect 1795 2584 1804 2624
rect 1844 2584 1853 2624
rect 1795 2583 1853 2584
rect 1987 2624 2045 2625
rect 1987 2584 1996 2624
rect 2036 2584 2045 2624
rect 1987 2583 2045 2584
rect 3235 2624 3293 2625
rect 3235 2584 3244 2624
rect 3284 2584 3293 2624
rect 3235 2583 3293 2584
rect 3811 2624 3869 2625
rect 3811 2584 3820 2624
rect 3860 2584 3869 2624
rect 3811 2583 3869 2584
rect 5059 2624 5117 2625
rect 5059 2584 5068 2624
rect 5108 2584 5117 2624
rect 5059 2583 5117 2584
rect 6123 2624 6165 2633
rect 6123 2584 6124 2624
rect 6164 2584 6165 2624
rect 6123 2575 6165 2584
rect 6219 2624 6261 2633
rect 6219 2584 6220 2624
rect 6260 2584 6261 2624
rect 6219 2575 6261 2584
rect 6499 2624 6557 2625
rect 6499 2584 6508 2624
rect 6548 2584 6557 2624
rect 6499 2583 6557 2584
rect 6787 2624 6845 2625
rect 6787 2584 6796 2624
rect 6836 2584 6845 2624
rect 6787 2583 6845 2584
rect 6883 2624 6941 2625
rect 6883 2584 6892 2624
rect 6932 2584 6941 2624
rect 6883 2583 6941 2584
rect 7083 2624 7125 2633
rect 7083 2584 7084 2624
rect 7124 2584 7125 2624
rect 7083 2575 7125 2584
rect 7179 2624 7221 2633
rect 7179 2584 7180 2624
rect 7220 2584 7221 2624
rect 7179 2575 7221 2584
rect 7272 2624 7330 2625
rect 7272 2584 7281 2624
rect 7321 2584 7330 2624
rect 7272 2583 7330 2584
rect 7947 2624 7989 2633
rect 7947 2584 7948 2624
rect 7988 2584 7989 2624
rect 7947 2575 7989 2584
rect 8043 2624 8085 2633
rect 8043 2584 8044 2624
rect 8084 2584 8085 2624
rect 8043 2575 8085 2584
rect 8323 2624 8381 2625
rect 8323 2584 8332 2624
rect 8372 2584 8381 2624
rect 8323 2583 8381 2584
rect 8715 2624 8757 2633
rect 8715 2584 8716 2624
rect 8756 2584 8757 2624
rect 8715 2575 8757 2584
rect 9003 2624 9045 2633
rect 9003 2584 9004 2624
rect 9044 2584 9045 2624
rect 9003 2575 9045 2584
rect 9483 2624 9525 2633
rect 9483 2584 9484 2624
rect 9524 2584 9525 2624
rect 9483 2575 9525 2584
rect 9675 2624 9717 2633
rect 9675 2584 9676 2624
rect 9716 2584 9717 2624
rect 9675 2575 9717 2584
rect 9955 2624 10013 2625
rect 9955 2584 9964 2624
rect 10004 2584 10013 2624
rect 9955 2583 10013 2584
rect 10251 2624 10293 2633
rect 10251 2584 10252 2624
rect 10292 2584 10293 2624
rect 10251 2575 10293 2584
rect 10347 2624 10389 2633
rect 10347 2584 10348 2624
rect 10388 2584 10389 2624
rect 10347 2575 10389 2584
rect 10923 2624 10965 2633
rect 10923 2584 10924 2624
rect 10964 2584 10965 2624
rect 10923 2575 10965 2584
rect 11019 2624 11061 2633
rect 12507 2626 12508 2666
rect 12548 2626 12549 2666
rect 11019 2584 11020 2624
rect 11060 2584 11061 2624
rect 11019 2575 11061 2584
rect 11971 2624 12029 2625
rect 11971 2584 11980 2624
rect 12020 2584 12029 2624
rect 12507 2617 12549 2626
rect 14755 2624 14813 2625
rect 11971 2583 12029 2584
rect 14755 2584 14764 2624
rect 14804 2584 14813 2624
rect 14755 2583 14813 2584
rect 16003 2624 16061 2625
rect 16003 2584 16012 2624
rect 16052 2584 16061 2624
rect 16003 2583 16061 2584
rect 16491 2624 16533 2633
rect 16491 2584 16492 2624
rect 16532 2584 16533 2624
rect 16491 2575 16533 2584
rect 16587 2624 16629 2633
rect 16587 2584 16588 2624
rect 16628 2584 16629 2624
rect 16587 2575 16629 2584
rect 16683 2624 16725 2633
rect 16683 2584 16684 2624
rect 16724 2584 16725 2624
rect 16683 2575 16725 2584
rect 16963 2624 17021 2625
rect 16963 2584 16972 2624
rect 17012 2584 17021 2624
rect 16963 2583 17021 2584
rect 17259 2624 17301 2633
rect 17259 2584 17260 2624
rect 17300 2584 17301 2624
rect 17259 2575 17301 2584
rect 17355 2624 17397 2633
rect 17355 2584 17356 2624
rect 17396 2584 17397 2624
rect 17355 2575 17397 2584
rect 17827 2624 17885 2625
rect 17827 2584 17836 2624
rect 17876 2584 17885 2624
rect 17827 2583 17885 2584
rect 17931 2624 17973 2633
rect 17931 2584 17932 2624
rect 17972 2584 17973 2624
rect 17931 2575 17973 2584
rect 18123 2624 18165 2633
rect 18123 2584 18124 2624
rect 18164 2584 18165 2624
rect 18123 2575 18165 2584
rect 18507 2624 18549 2633
rect 18507 2584 18508 2624
rect 18548 2584 18549 2624
rect 18507 2575 18549 2584
rect 18603 2624 18645 2633
rect 18603 2584 18604 2624
rect 18644 2584 18645 2624
rect 18603 2575 18645 2584
rect 18699 2624 18741 2633
rect 18699 2584 18700 2624
rect 18740 2584 18741 2624
rect 18699 2575 18741 2584
rect 18795 2624 18837 2633
rect 18795 2584 18796 2624
rect 18836 2584 18837 2624
rect 18795 2575 18837 2584
rect 19179 2624 19221 2633
rect 19179 2584 19180 2624
rect 19220 2584 19221 2624
rect 19179 2575 19221 2584
rect 19275 2624 19317 2633
rect 19275 2584 19276 2624
rect 19316 2584 19317 2624
rect 19275 2575 19317 2584
rect 19371 2624 19413 2633
rect 19371 2584 19372 2624
rect 19412 2584 19413 2624
rect 19371 2575 19413 2584
rect 19651 2624 19709 2625
rect 19651 2584 19660 2624
rect 19700 2584 19709 2624
rect 19651 2583 19709 2584
rect 19755 2624 19797 2633
rect 19755 2584 19756 2624
rect 19796 2584 19797 2624
rect 19755 2575 19797 2584
rect 19947 2624 19989 2633
rect 19947 2584 19948 2624
rect 19988 2584 19989 2624
rect 19947 2575 19989 2584
rect 1707 2540 1749 2549
rect 1707 2500 1708 2540
rect 1748 2500 1749 2540
rect 1707 2491 1749 2500
rect 12651 2540 12693 2549
rect 12651 2500 12652 2540
rect 12692 2500 12693 2540
rect 12651 2491 12693 2500
rect 19851 2540 19893 2549
rect 19851 2500 19852 2540
rect 19892 2500 19893 2540
rect 19851 2491 19893 2500
rect 5643 2456 5685 2465
rect 5643 2416 5644 2456
rect 5684 2416 5685 2456
rect 5643 2407 5685 2416
rect 6979 2456 7037 2457
rect 6979 2416 6988 2456
rect 7028 2416 7037 2456
rect 6979 2415 7037 2416
rect 9187 2456 9245 2457
rect 9187 2416 9196 2456
rect 9236 2416 9245 2456
rect 9187 2415 9245 2416
rect 13803 2456 13845 2465
rect 13803 2416 13804 2456
rect 13844 2416 13845 2456
rect 13803 2407 13845 2416
rect 14379 2456 14421 2465
rect 14379 2416 14380 2456
rect 14420 2416 14421 2456
rect 14379 2407 14421 2416
rect 16387 2456 16445 2457
rect 16387 2416 16396 2456
rect 16436 2416 16445 2456
rect 16387 2415 16445 2416
rect 1152 2288 20452 2312
rect 1152 2248 4928 2288
rect 4968 2248 5010 2288
rect 5050 2248 5092 2288
rect 5132 2248 5174 2288
rect 5214 2248 5256 2288
rect 5296 2248 20048 2288
rect 20088 2248 20130 2288
rect 20170 2248 20212 2288
rect 20252 2248 20294 2288
rect 20334 2248 20376 2288
rect 20416 2248 20452 2288
rect 1152 2224 20452 2248
rect 2763 2120 2805 2129
rect 2763 2080 2764 2120
rect 2804 2080 2805 2120
rect 2763 2071 2805 2080
rect 8323 2120 8381 2121
rect 8323 2080 8332 2120
rect 8372 2080 8381 2120
rect 8323 2079 8381 2080
rect 8611 2120 8669 2121
rect 8611 2080 8620 2120
rect 8660 2080 8669 2120
rect 8611 2079 8669 2080
rect 8899 2120 8957 2121
rect 8899 2080 8908 2120
rect 8948 2080 8957 2120
rect 8899 2079 8957 2080
rect 9867 2120 9909 2129
rect 9867 2080 9868 2120
rect 9908 2080 9909 2120
rect 9867 2071 9909 2080
rect 14955 2120 14997 2129
rect 14955 2080 14956 2120
rect 14996 2080 14997 2120
rect 14955 2071 14997 2080
rect 17355 2124 17397 2133
rect 17355 2084 17356 2124
rect 17396 2084 17397 2124
rect 17355 2075 17397 2084
rect 19851 2120 19893 2129
rect 19851 2080 19852 2120
rect 19892 2080 19893 2120
rect 19851 2071 19893 2080
rect 12939 2036 12981 2045
rect 12939 1996 12940 2036
rect 12980 1996 12981 2036
rect 12939 1987 12981 1996
rect 1315 1952 1373 1953
rect 1315 1912 1324 1952
rect 1364 1912 1373 1952
rect 1315 1911 1373 1912
rect 2563 1952 2621 1953
rect 2563 1912 2572 1952
rect 2612 1912 2621 1952
rect 2563 1911 2621 1912
rect 3523 1952 3581 1953
rect 3523 1912 3532 1952
rect 3572 1912 3581 1952
rect 3523 1911 3581 1912
rect 4771 1952 4829 1953
rect 4771 1912 4780 1952
rect 4820 1912 4829 1952
rect 4771 1911 4829 1912
rect 4963 1952 5021 1953
rect 4963 1912 4972 1952
rect 5012 1912 5021 1952
rect 4963 1911 5021 1912
rect 6211 1952 6269 1953
rect 6211 1912 6220 1952
rect 6260 1912 6269 1952
rect 6211 1911 6269 1912
rect 6987 1952 7029 1961
rect 6987 1912 6988 1952
rect 7028 1912 7029 1952
rect 6987 1903 7029 1912
rect 7179 1952 7221 1961
rect 7179 1912 7180 1952
rect 7220 1912 7221 1952
rect 7179 1903 7221 1912
rect 7267 1952 7325 1953
rect 7267 1912 7276 1952
rect 7316 1912 7325 1952
rect 7267 1911 7325 1912
rect 7659 1952 7701 1961
rect 7659 1912 7660 1952
rect 7700 1912 7701 1952
rect 7659 1903 7701 1912
rect 7755 1952 7797 1961
rect 7755 1912 7756 1952
rect 7796 1912 7797 1952
rect 7755 1903 7797 1912
rect 7851 1952 7893 1961
rect 7851 1912 7852 1952
rect 7892 1912 7893 1952
rect 7851 1903 7893 1912
rect 7947 1952 7989 1961
rect 7947 1912 7948 1952
rect 7988 1912 7989 1952
rect 7947 1903 7989 1912
rect 8131 1952 8189 1953
rect 8131 1912 8140 1952
rect 8180 1912 8189 1952
rect 8131 1911 8189 1912
rect 8235 1952 8277 1961
rect 8235 1912 8236 1952
rect 8276 1912 8277 1952
rect 8707 1952 8765 1953
rect 8235 1903 8277 1912
rect 8427 1941 8469 1950
rect 8427 1901 8428 1941
rect 8468 1901 8469 1941
rect 8707 1912 8716 1952
rect 8756 1912 8765 1952
rect 8707 1911 8765 1912
rect 9771 1952 9813 1961
rect 9771 1912 9772 1952
rect 9812 1912 9813 1952
rect 9771 1903 9813 1912
rect 10059 1952 10101 1961
rect 10059 1912 10060 1952
rect 10100 1912 10101 1952
rect 10059 1903 10101 1912
rect 11491 1952 11549 1953
rect 11491 1912 11500 1952
rect 11540 1912 11549 1952
rect 11491 1911 11549 1912
rect 12739 1952 12797 1953
rect 12739 1912 12748 1952
rect 12788 1912 12797 1952
rect 12739 1911 12797 1912
rect 13227 1952 13269 1961
rect 13227 1912 13228 1952
rect 13268 1912 13269 1952
rect 13227 1903 13269 1912
rect 13323 1952 13365 1961
rect 13323 1912 13324 1952
rect 13364 1912 13365 1952
rect 13323 1903 13365 1912
rect 13707 1952 13749 1961
rect 13707 1912 13708 1952
rect 13748 1912 13749 1952
rect 13707 1903 13749 1912
rect 14275 1952 14333 1953
rect 14275 1912 14284 1952
rect 14324 1912 14333 1952
rect 15235 1952 15293 1953
rect 14275 1911 14333 1912
rect 14763 1938 14805 1947
rect 8427 1892 8469 1901
rect 14763 1898 14764 1938
rect 14804 1898 14805 1938
rect 15235 1912 15244 1952
rect 15284 1912 15293 1952
rect 15235 1911 15293 1912
rect 16483 1952 16541 1953
rect 16483 1912 16492 1952
rect 16532 1912 16541 1952
rect 16483 1911 16541 1912
rect 17163 1952 17205 1961
rect 17163 1912 17164 1952
rect 17204 1912 17205 1952
rect 17163 1903 17205 1912
rect 17251 1952 17309 1953
rect 17251 1912 17260 1952
rect 17300 1912 17309 1952
rect 17251 1911 17309 1912
rect 17539 1952 17597 1953
rect 17539 1912 17548 1952
rect 17588 1912 17597 1952
rect 17539 1911 17597 1912
rect 17643 1952 17685 1961
rect 17643 1912 17644 1952
rect 17684 1912 17685 1952
rect 17643 1903 17685 1912
rect 17835 1952 17877 1961
rect 17835 1912 17836 1952
rect 17876 1912 17877 1952
rect 17835 1903 17877 1912
rect 18027 1952 18069 1961
rect 18027 1912 18028 1952
rect 18068 1912 18069 1952
rect 18027 1903 18069 1912
rect 18115 1952 18173 1953
rect 18115 1912 18124 1952
rect 18164 1912 18173 1952
rect 18115 1911 18173 1912
rect 18403 1952 18461 1953
rect 18403 1912 18412 1952
rect 18452 1912 18461 1952
rect 18403 1911 18461 1912
rect 19651 1952 19709 1953
rect 19651 1912 19660 1952
rect 19700 1912 19709 1952
rect 19651 1911 19709 1912
rect 14763 1889 14805 1898
rect 2947 1868 3005 1869
rect 2947 1828 2956 1868
rect 2996 1828 3005 1868
rect 2947 1827 3005 1828
rect 6595 1868 6653 1869
rect 6595 1828 6604 1868
rect 6644 1828 6653 1868
rect 6595 1827 6653 1828
rect 9187 1868 9245 1869
rect 9187 1828 9196 1868
rect 9236 1828 9245 1868
rect 9187 1827 9245 1828
rect 10339 1868 10397 1869
rect 10339 1828 10348 1868
rect 10388 1828 10397 1868
rect 10339 1827 10397 1828
rect 10723 1868 10781 1869
rect 10723 1828 10732 1868
rect 10772 1828 10781 1868
rect 10723 1827 10781 1828
rect 11107 1868 11165 1869
rect 11107 1828 11116 1868
rect 11156 1828 11165 1868
rect 11107 1827 11165 1828
rect 13803 1868 13845 1877
rect 13803 1828 13804 1868
rect 13844 1828 13845 1868
rect 13803 1819 13845 1828
rect 6987 1784 7029 1793
rect 6987 1744 6988 1784
rect 7028 1744 7029 1784
rect 6987 1735 7029 1744
rect 16875 1784 16917 1793
rect 16875 1744 16876 1784
rect 16916 1744 16917 1784
rect 16875 1735 16917 1744
rect 17835 1784 17877 1793
rect 17835 1744 17836 1784
rect 17876 1744 17877 1784
rect 17835 1735 17877 1744
rect 3147 1700 3189 1709
rect 3147 1660 3148 1700
rect 3188 1660 3189 1700
rect 3147 1651 3189 1660
rect 3339 1700 3381 1709
rect 3339 1660 3340 1700
rect 3380 1660 3381 1700
rect 3339 1651 3381 1660
rect 6411 1700 6453 1709
rect 6411 1660 6412 1700
rect 6452 1660 6453 1700
rect 6411 1651 6453 1660
rect 6795 1700 6837 1709
rect 6795 1660 6796 1700
rect 6836 1660 6837 1700
rect 6795 1651 6837 1660
rect 9387 1700 9429 1709
rect 9387 1660 9388 1700
rect 9428 1660 9429 1700
rect 9387 1651 9429 1660
rect 10539 1700 10581 1709
rect 10539 1660 10540 1700
rect 10580 1660 10581 1700
rect 10539 1651 10581 1660
rect 10923 1700 10965 1709
rect 10923 1660 10924 1700
rect 10964 1660 10965 1700
rect 10923 1651 10965 1660
rect 11307 1700 11349 1709
rect 11307 1660 11308 1700
rect 11348 1660 11349 1700
rect 11307 1651 11349 1660
rect 16683 1700 16725 1709
rect 16683 1660 16684 1700
rect 16724 1660 16725 1700
rect 16683 1651 16725 1660
rect 1152 1532 20352 1556
rect 1152 1492 3688 1532
rect 3728 1492 3770 1532
rect 3810 1492 3852 1532
rect 3892 1492 3934 1532
rect 3974 1492 4016 1532
rect 4056 1492 18808 1532
rect 18848 1492 18890 1532
rect 18930 1492 18972 1532
rect 19012 1492 19054 1532
rect 19094 1492 19136 1532
rect 19176 1492 20352 1532
rect 1152 1468 20352 1492
rect 6019 1364 6077 1365
rect 6019 1324 6028 1364
rect 6068 1324 6077 1364
rect 6019 1323 6077 1324
rect 14667 1364 14709 1373
rect 14667 1324 14668 1364
rect 14708 1324 14709 1364
rect 14667 1315 14709 1324
rect 17355 1364 17397 1373
rect 17355 1324 17356 1364
rect 17396 1324 17397 1364
rect 17355 1315 17397 1324
rect 17739 1364 17781 1373
rect 17739 1324 17740 1364
rect 17780 1324 17781 1364
rect 17739 1315 17781 1324
rect 6219 1280 6261 1289
rect 6219 1240 6220 1280
rect 6260 1240 6261 1280
rect 6219 1231 6261 1240
rect 9195 1280 9237 1289
rect 9195 1240 9196 1280
rect 9236 1240 9237 1280
rect 9195 1231 9237 1240
rect 17163 1280 17205 1289
rect 17163 1240 17164 1280
rect 17204 1240 17205 1280
rect 17163 1231 17205 1240
rect 19563 1280 19605 1289
rect 19563 1240 19564 1280
rect 19604 1240 19605 1280
rect 19563 1231 19605 1240
rect 2371 1196 2429 1197
rect 2371 1156 2380 1196
rect 2420 1156 2429 1196
rect 2371 1155 2429 1156
rect 4387 1196 4445 1197
rect 4387 1156 4396 1196
rect 4436 1156 4445 1196
rect 4387 1155 4445 1156
rect 7651 1196 7709 1197
rect 7651 1156 7660 1196
rect 7700 1156 7709 1196
rect 7651 1155 7709 1156
rect 8035 1196 8093 1197
rect 8035 1156 8044 1196
rect 8084 1156 8093 1196
rect 8035 1155 8093 1156
rect 8419 1196 8477 1197
rect 8419 1156 8428 1196
rect 8468 1156 8477 1196
rect 8419 1155 8477 1156
rect 8803 1196 8861 1197
rect 8803 1156 8812 1196
rect 8852 1156 8861 1196
rect 8803 1155 8861 1156
rect 9571 1196 9629 1197
rect 9571 1156 9580 1196
rect 9620 1156 9629 1196
rect 9571 1155 9629 1156
rect 9955 1196 10013 1197
rect 9955 1156 9964 1196
rect 10004 1156 10013 1196
rect 9955 1155 10013 1156
rect 10339 1196 10397 1197
rect 10339 1156 10348 1196
rect 10388 1156 10397 1196
rect 10339 1155 10397 1156
rect 10915 1196 10973 1197
rect 10915 1156 10924 1196
rect 10964 1156 10973 1196
rect 10915 1155 10973 1156
rect 11203 1196 11261 1197
rect 11203 1156 11212 1196
rect 11252 1156 11261 1196
rect 11203 1155 11261 1156
rect 11779 1196 11837 1197
rect 11779 1156 11788 1196
rect 11828 1156 11837 1196
rect 11779 1155 11837 1156
rect 14851 1196 14909 1197
rect 14851 1156 14860 1196
rect 14900 1156 14909 1196
rect 14851 1155 14909 1156
rect 15523 1196 15581 1197
rect 15523 1156 15532 1196
rect 15572 1156 15581 1196
rect 15523 1155 15581 1156
rect 2755 1112 2813 1113
rect 2755 1072 2764 1112
rect 2804 1072 2813 1112
rect 2755 1071 2813 1072
rect 4003 1112 4061 1113
rect 4003 1072 4012 1112
rect 4052 1072 4061 1112
rect 4003 1071 4061 1072
rect 4779 1112 4821 1121
rect 4779 1072 4780 1112
rect 4820 1072 4821 1112
rect 4779 1063 4821 1072
rect 4875 1112 4917 1121
rect 4875 1072 4876 1112
rect 4916 1072 4917 1112
rect 4875 1063 4917 1072
rect 4971 1112 5013 1121
rect 4971 1072 4972 1112
rect 5012 1072 5013 1112
rect 4971 1063 5013 1072
rect 5067 1112 5109 1121
rect 5067 1072 5068 1112
rect 5108 1072 5109 1112
rect 5067 1063 5109 1072
rect 5347 1112 5405 1113
rect 5347 1072 5356 1112
rect 5396 1072 5405 1112
rect 5347 1071 5405 1072
rect 5643 1112 5685 1121
rect 5643 1072 5644 1112
rect 5684 1072 5685 1112
rect 5643 1063 5685 1072
rect 6307 1112 6365 1113
rect 6307 1072 6316 1112
rect 6356 1072 6365 1112
rect 6307 1071 6365 1072
rect 6507 1112 6549 1121
rect 6507 1072 6508 1112
rect 6548 1072 6549 1112
rect 6507 1063 6549 1072
rect 6603 1112 6645 1121
rect 6603 1072 6604 1112
rect 6644 1072 6645 1112
rect 6603 1063 6645 1072
rect 7371 1112 7413 1121
rect 7371 1072 7372 1112
rect 7412 1072 7413 1112
rect 13219 1112 13277 1113
rect 7371 1063 7413 1072
rect 7464 1103 7522 1104
rect 7464 1063 7473 1103
rect 7513 1063 7522 1103
rect 13219 1072 13228 1112
rect 13268 1072 13277 1112
rect 13219 1071 13277 1072
rect 14467 1112 14525 1113
rect 14467 1072 14476 1112
rect 14516 1072 14525 1112
rect 14467 1071 14525 1072
rect 15715 1112 15773 1113
rect 15715 1072 15724 1112
rect 15764 1072 15773 1112
rect 15715 1071 15773 1072
rect 16963 1112 17021 1113
rect 16963 1072 16972 1112
rect 17012 1072 17021 1112
rect 16963 1071 17021 1072
rect 17443 1112 17501 1113
rect 17443 1072 17452 1112
rect 17492 1072 17501 1112
rect 17443 1071 17501 1072
rect 17635 1112 17693 1113
rect 17635 1072 17644 1112
rect 17684 1072 17693 1112
rect 17635 1071 17693 1072
rect 18115 1112 18173 1113
rect 18115 1072 18124 1112
rect 18164 1072 18173 1112
rect 18115 1071 18173 1072
rect 19363 1112 19421 1113
rect 19363 1072 19372 1112
rect 19412 1072 19421 1112
rect 19363 1071 19421 1072
rect 7464 1062 7522 1063
rect 4203 1028 4245 1037
rect 4203 988 4204 1028
rect 4244 988 4245 1028
rect 4203 979 4245 988
rect 5739 1028 5781 1037
rect 5739 988 5740 1028
rect 5780 988 5781 1028
rect 5739 979 5781 988
rect 2571 944 2613 953
rect 2571 904 2572 944
rect 2612 904 2613 944
rect 2571 895 2613 904
rect 4587 944 4629 953
rect 4587 904 4588 944
rect 4628 904 4629 944
rect 4587 895 4629 904
rect 6787 944 6845 945
rect 6787 904 6796 944
rect 6836 904 6845 944
rect 6787 903 6845 904
rect 7171 944 7229 945
rect 7171 904 7180 944
rect 7220 904 7229 944
rect 7171 903 7229 904
rect 7851 944 7893 953
rect 7851 904 7852 944
rect 7892 904 7893 944
rect 7851 895 7893 904
rect 8235 944 8277 953
rect 8235 904 8236 944
rect 8276 904 8277 944
rect 8235 895 8277 904
rect 8619 944 8661 953
rect 8619 904 8620 944
rect 8660 904 8661 944
rect 8619 895 8661 904
rect 9003 944 9045 953
rect 9003 904 9004 944
rect 9044 904 9045 944
rect 9003 895 9045 904
rect 9771 944 9813 953
rect 9771 904 9772 944
rect 9812 904 9813 944
rect 9771 895 9813 904
rect 10155 944 10197 953
rect 10155 904 10156 944
rect 10196 904 10197 944
rect 10155 895 10197 904
rect 10539 944 10581 953
rect 10539 904 10540 944
rect 10580 904 10581 944
rect 10539 895 10581 904
rect 10731 944 10773 953
rect 10731 904 10732 944
rect 10772 904 10773 944
rect 10731 895 10773 904
rect 11403 944 11445 953
rect 11403 904 11404 944
rect 11444 904 11445 944
rect 11403 895 11445 904
rect 11595 944 11637 953
rect 11595 904 11596 944
rect 11636 904 11637 944
rect 11595 895 11637 904
rect 15051 944 15093 953
rect 15051 904 15052 944
rect 15092 904 15093 944
rect 15051 895 15093 904
rect 15339 944 15381 953
rect 15339 904 15340 944
rect 15380 904 15381 944
rect 15339 895 15381 904
rect 1152 776 20452 800
rect 1152 736 4928 776
rect 4968 736 5010 776
rect 5050 736 5092 776
rect 5132 736 5174 776
rect 5214 736 5256 776
rect 5296 736 20048 776
rect 20088 736 20130 776
rect 20170 736 20212 776
rect 20252 736 20294 776
rect 20334 736 20376 776
rect 20416 736 20452 776
rect 1152 712 20452 736
<< via1 >>
rect 4928 41560 4968 41600
rect 5010 41560 5050 41600
rect 5092 41560 5132 41600
rect 5174 41560 5214 41600
rect 5256 41560 5296 41600
rect 20048 41560 20088 41600
rect 20130 41560 20170 41600
rect 20212 41560 20252 41600
rect 20294 41560 20334 41600
rect 20376 41560 20416 41600
rect 8236 41392 8276 41432
rect 18604 41392 18644 41432
rect 18988 41392 19028 41432
rect 19372 41392 19412 41432
rect 1804 41224 1844 41264
rect 3052 41224 3092 41264
rect 3436 41224 3476 41264
rect 4684 41224 4724 41264
rect 6316 41224 6356 41264
rect 7564 41224 7604 41264
rect 8716 41224 8756 41264
rect 9964 41224 10004 41264
rect 10348 41224 10388 41264
rect 11596 41224 11636 41264
rect 12172 41224 12212 41264
rect 13420 41224 13460 41264
rect 13804 41224 13844 41264
rect 15052 41224 15092 41264
rect 16684 41224 16724 41264
rect 17932 41224 17972 41264
rect 8044 41140 8084 41180
rect 15436 41140 15476 41180
rect 15820 41140 15860 41180
rect 16204 41140 16244 41180
rect 18796 41140 18836 41180
rect 19180 41140 19220 41180
rect 19564 41140 19604 41180
rect 19756 41140 19796 41180
rect 1324 41056 1364 41096
rect 18316 41056 18356 41096
rect 3244 40972 3284 41012
rect 4876 40972 4916 41012
rect 6124 40972 6164 41012
rect 10156 40972 10196 41012
rect 11788 40972 11828 41012
rect 11980 40972 12020 41012
rect 13612 40972 13652 41012
rect 15244 40972 15284 41012
rect 15628 40972 15668 41012
rect 16012 40972 16052 41012
rect 18124 40972 18164 41012
rect 19948 40972 19988 41012
rect 3688 40804 3728 40844
rect 3770 40804 3810 40844
rect 3852 40804 3892 40844
rect 3934 40804 3974 40844
rect 4016 40804 4056 40844
rect 18808 40804 18848 40844
rect 18890 40804 18930 40844
rect 18972 40804 19012 40844
rect 19054 40804 19094 40844
rect 19136 40804 19176 40844
rect 1708 40636 1748 40676
rect 3916 40636 3956 40676
rect 6220 40636 6260 40676
rect 13708 40636 13748 40676
rect 17452 40636 17492 40676
rect 18316 40636 18356 40676
rect 19084 40636 19124 40676
rect 19468 40636 19508 40676
rect 19852 40636 19892 40676
rect 1324 40552 1364 40592
rect 3532 40552 3572 40592
rect 14092 40552 14132 40592
rect 14476 40552 14516 40592
rect 14860 40552 14900 40592
rect 15244 40552 15284 40592
rect 15628 40552 15668 40592
rect 16012 40552 16052 40592
rect 16396 40552 16436 40592
rect 17644 40552 17684 40592
rect 18700 40552 18740 40592
rect 1516 40468 1556 40508
rect 3724 40468 3764 40508
rect 6028 40468 6068 40508
rect 13900 40468 13940 40508
rect 14284 40468 14324 40508
rect 14668 40468 14708 40508
rect 15052 40468 15092 40508
rect 15436 40468 15476 40508
rect 15820 40468 15860 40508
rect 16204 40468 16244 40508
rect 16588 40479 16628 40519
rect 16972 40468 17012 40508
rect 17260 40468 17300 40508
rect 17836 40468 17876 40508
rect 18028 40468 18068 40508
rect 2092 40384 2132 40424
rect 3340 40384 3380 40424
rect 4108 40384 4148 40424
rect 5356 40384 5396 40424
rect 6412 40384 6452 40424
rect 7660 40384 7700 40424
rect 8140 40384 8180 40424
rect 9388 40384 9428 40424
rect 10156 40384 10196 40424
rect 10252 40384 10292 40424
rect 10636 40384 10676 40424
rect 11740 40426 11780 40466
rect 18508 40468 18548 40508
rect 18892 40468 18932 40508
rect 19276 40468 19316 40508
rect 19660 40468 19700 40508
rect 20044 40468 20084 40508
rect 10732 40384 10772 40424
rect 11212 40384 11252 40424
rect 12268 40384 12308 40424
rect 13516 40384 13556 40424
rect 5548 40300 5588 40340
rect 9772 40300 9812 40340
rect 7852 40216 7892 40256
rect 9580 40216 9620 40256
rect 11884 40174 11924 40214
rect 12076 40216 12116 40256
rect 16780 40216 16820 40256
rect 4928 40048 4968 40088
rect 5010 40048 5050 40088
rect 5092 40048 5132 40088
rect 5174 40048 5214 40088
rect 5256 40048 5296 40088
rect 20048 40048 20088 40088
rect 20130 40048 20170 40088
rect 20212 40048 20252 40088
rect 20294 40048 20334 40088
rect 20376 40048 20416 40088
rect 1420 39880 1460 39920
rect 3532 39880 3572 39920
rect 10252 39880 10292 39920
rect 13132 39880 13172 39920
rect 17548 39880 17588 39920
rect 18412 39880 18452 39920
rect 18604 39880 18644 39920
rect 18988 39880 19028 39920
rect 12748 39796 12788 39836
rect 1708 39712 1748 39752
rect 2956 39712 2996 39752
rect 4396 39712 4436 39752
rect 5644 39712 5684 39752
rect 6988 39712 7028 39752
rect 8236 39712 8276 39752
rect 8620 39712 8660 39752
rect 9868 39712 9908 39752
rect 11020 39712 11060 39752
rect 11116 39712 11156 39752
rect 12076 39712 12116 39752
rect 12556 39707 12596 39747
rect 13324 39712 13364 39752
rect 14572 39712 14612 39752
rect 15244 39712 15284 39752
rect 16492 39712 16532 39752
rect 1228 39628 1268 39668
rect 3340 39628 3380 39668
rect 10444 39628 10484 39668
rect 11500 39628 11540 39668
rect 11596 39628 11636 39668
rect 12940 39628 12980 39668
rect 17068 39628 17108 39668
rect 17740 39628 17780 39668
rect 18220 39628 18260 39668
rect 18796 39628 18836 39668
rect 19180 39628 19220 39668
rect 19372 39628 19412 39668
rect 19756 39628 19796 39668
rect 3820 39544 3860 39584
rect 6028 39544 6068 39584
rect 10636 39544 10676 39584
rect 17260 39544 17300 39584
rect 18028 39544 18068 39584
rect 20140 39544 20180 39584
rect 3148 39460 3188 39500
rect 5836 39460 5876 39500
rect 8428 39460 8468 39500
rect 10060 39460 10100 39500
rect 14764 39460 14804 39500
rect 16684 39460 16724 39500
rect 16876 39460 16916 39500
rect 19564 39460 19604 39500
rect 19948 39460 19988 39500
rect 3688 39292 3728 39332
rect 3770 39292 3810 39332
rect 3852 39292 3892 39332
rect 3934 39292 3974 39332
rect 4016 39292 4056 39332
rect 18808 39292 18848 39332
rect 18890 39292 18930 39332
rect 18972 39292 19012 39332
rect 19054 39292 19094 39332
rect 19136 39292 19176 39332
rect 17452 39124 17492 39164
rect 1516 39040 1556 39080
rect 4396 39040 4436 39080
rect 14668 39040 14708 39080
rect 17644 39040 17684 39080
rect 18508 39040 18548 39080
rect 1324 38956 1364 38996
rect 4204 38956 4244 38996
rect 6316 38956 6356 38996
rect 8332 38956 8372 38996
rect 12076 38956 12116 38996
rect 14476 38956 14516 38996
rect 15532 38956 15572 38996
rect 16876 38956 16916 38996
rect 17260 38956 17300 38996
rect 17836 38956 17876 38996
rect 18700 38956 18740 38996
rect 19276 38956 19316 38996
rect 19660 38956 19700 38996
rect 20044 38956 20084 38996
rect 1708 38872 1748 38912
rect 2956 38872 2996 38912
rect 5836 38872 5876 38912
rect 5932 38872 5972 38912
rect 6412 38872 6452 38912
rect 6892 38872 6932 38912
rect 7372 38886 7412 38926
rect 7852 38872 7892 38912
rect 7948 38872 7988 38912
rect 8428 38872 8468 38912
rect 8908 38872 8948 38912
rect 9388 38886 9428 38926
rect 10252 38872 10292 38912
rect 11500 38872 11540 38912
rect 12556 38872 12596 38912
rect 13804 38872 13844 38912
rect 14956 38872 14996 38912
rect 15052 38872 15092 38912
rect 15436 38872 15476 38912
rect 16012 38872 16052 38912
rect 16540 38881 16580 38921
rect 3148 38704 3188 38744
rect 3340 38704 3380 38744
rect 7564 38704 7604 38744
rect 9580 38704 9620 38744
rect 11692 38704 11732 38744
rect 12268 38704 12308 38744
rect 13996 38704 14036 38744
rect 16684 38704 16724 38744
rect 17068 38704 17108 38744
rect 18220 38704 18260 38744
rect 18988 38704 19028 38744
rect 19468 38704 19508 38744
rect 19852 38704 19892 38744
rect 20236 38704 20276 38744
rect 4928 38536 4968 38576
rect 5010 38536 5050 38576
rect 5092 38536 5132 38576
rect 5174 38536 5214 38576
rect 5256 38536 5296 38576
rect 20048 38536 20088 38576
rect 20130 38536 20170 38576
rect 20212 38536 20252 38576
rect 20294 38536 20334 38576
rect 20376 38536 20416 38576
rect 1420 38368 1460 38408
rect 1804 38368 1844 38408
rect 6892 38368 6932 38408
rect 7276 38368 7316 38408
rect 12268 38368 12308 38408
rect 12652 38368 12692 38408
rect 13036 38368 13076 38408
rect 13420 38368 13460 38408
rect 17068 38368 17108 38408
rect 19180 38368 19220 38408
rect 4204 38284 4244 38324
rect 6508 38284 6548 38324
rect 11692 38284 11732 38324
rect 20140 38284 20180 38324
rect 2476 38200 2516 38240
rect 2572 38200 2612 38240
rect 3532 38200 3572 38240
rect 4012 38195 4052 38235
rect 4780 38200 4820 38240
rect 4876 38200 4916 38240
rect 5836 38200 5876 38240
rect 7852 38200 7892 38240
rect 9100 38200 9140 38240
rect 9580 38200 9620 38240
rect 1228 38116 1268 38156
rect 1612 38116 1652 38156
rect 1996 38116 2036 38156
rect 2956 38116 2996 38156
rect 3052 38116 3092 38156
rect 5260 38116 5300 38156
rect 5356 38116 5396 38156
rect 6364 38158 6404 38198
rect 9964 38200 10004 38240
rect 10060 38200 10100 38240
rect 10540 38200 10580 38240
rect 11020 38200 11060 38240
rect 11548 38190 11588 38230
rect 13612 38200 13652 38240
rect 14860 38200 14900 38240
rect 15340 38200 15380 38240
rect 15436 38200 15476 38240
rect 15820 38200 15860 38240
rect 15916 38200 15956 38240
rect 16396 38200 16436 38240
rect 16876 38186 16916 38226
rect 17452 38200 17492 38240
rect 18700 38200 18740 38240
rect 7084 38116 7124 38156
rect 7468 38116 7508 38156
rect 10444 38116 10484 38156
rect 12076 38116 12116 38156
rect 12460 38116 12500 38156
rect 12844 38116 12884 38156
rect 13228 38116 13268 38156
rect 18988 38116 19028 38156
rect 19372 38116 19412 38156
rect 19756 38116 19796 38156
rect 15052 38032 15092 38072
rect 2188 37948 2228 37988
rect 9292 37948 9332 37988
rect 17260 37948 17300 37988
rect 19564 37948 19604 37988
rect 19948 37948 19988 37988
rect 3688 37780 3728 37820
rect 3770 37780 3810 37820
rect 3852 37780 3892 37820
rect 3934 37780 3974 37820
rect 4016 37780 4056 37820
rect 18808 37780 18848 37820
rect 18890 37780 18930 37820
rect 18972 37780 19012 37820
rect 19054 37780 19094 37820
rect 19136 37780 19176 37820
rect 1804 37612 1844 37652
rect 4684 37612 4724 37652
rect 5068 37612 5108 37652
rect 5452 37612 5492 37652
rect 15436 37612 15476 37652
rect 17068 37612 17108 37652
rect 1420 37528 1460 37568
rect 7372 37528 7412 37568
rect 17452 37528 17492 37568
rect 1228 37444 1268 37484
rect 1612 37444 1652 37484
rect 4492 37444 4532 37484
rect 4876 37444 4916 37484
rect 5260 37444 5300 37484
rect 2476 37360 2516 37400
rect 2572 37360 2612 37400
rect 2956 37360 2996 37400
rect 4060 37402 4100 37442
rect 15244 37444 15284 37484
rect 17260 37444 17300 37484
rect 18220 37444 18260 37484
rect 3052 37360 3092 37400
rect 3532 37360 3572 37400
rect 5644 37360 5684 37400
rect 6892 37360 6932 37400
rect 7660 37360 7700 37400
rect 7756 37360 7796 37400
rect 8140 37360 8180 37400
rect 9244 37402 9284 37442
rect 19660 37444 19700 37484
rect 20044 37444 20084 37484
rect 8236 37360 8276 37400
rect 8716 37360 8756 37400
rect 9772 37360 9812 37400
rect 11020 37360 11060 37400
rect 11500 37360 11540 37400
rect 12748 37360 12788 37400
rect 13324 37360 13364 37400
rect 14572 37360 14612 37400
rect 15628 37360 15668 37400
rect 16876 37360 16916 37400
rect 17740 37360 17780 37400
rect 17836 37360 17876 37400
rect 18316 37360 18356 37400
rect 18796 37360 18836 37400
rect 19276 37374 19316 37414
rect 7084 37276 7124 37316
rect 19468 37276 19508 37316
rect 1996 37192 2036 37232
rect 4204 37192 4244 37232
rect 7276 37192 7316 37232
rect 9388 37150 9428 37190
rect 9580 37192 9620 37232
rect 12940 37192 12980 37232
rect 14764 37192 14804 37232
rect 19852 37192 19892 37232
rect 20236 37192 20276 37232
rect 4928 37024 4968 37064
rect 5010 37024 5050 37064
rect 5092 37024 5132 37064
rect 5174 37024 5214 37064
rect 5256 37024 5296 37064
rect 20048 37024 20088 37064
rect 20130 37024 20170 37064
rect 20212 37024 20252 37064
rect 20294 37024 20334 37064
rect 20376 37024 20416 37064
rect 1516 36856 1556 36896
rect 1900 36856 1940 36896
rect 3820 36856 3860 36896
rect 4684 36856 4724 36896
rect 7084 36856 7124 36896
rect 14668 36856 14708 36896
rect 15052 36856 15092 36896
rect 17068 36856 17108 36896
rect 19180 36856 19220 36896
rect 19564 36856 19604 36896
rect 12172 36772 12212 36812
rect 14188 36772 14228 36812
rect 4972 36688 5012 36728
rect 6220 36688 6260 36728
rect 7468 36688 7508 36728
rect 8716 36688 8756 36728
rect 9100 36688 9140 36728
rect 10348 36688 10388 36728
rect 10732 36688 10772 36728
rect 12460 36688 12500 36728
rect 1324 36604 1364 36644
rect 1708 36604 1748 36644
rect 2188 36604 2228 36644
rect 11980 36646 12020 36686
rect 12556 36688 12596 36728
rect 13516 36688 13556 36728
rect 13996 36683 14036 36723
rect 15340 36688 15380 36728
rect 15436 36688 15476 36728
rect 16396 36688 16436 36728
rect 16876 36674 16916 36714
rect 17452 36688 17492 36728
rect 18700 36688 18740 36728
rect 4300 36604 4340 36644
rect 4492 36604 4532 36644
rect 6892 36604 6932 36644
rect 12940 36604 12980 36644
rect 13036 36604 13076 36644
rect 14476 36604 14516 36644
rect 14860 36604 14900 36644
rect 15820 36604 15860 36644
rect 15916 36604 15956 36644
rect 18988 36604 19028 36644
rect 19372 36604 19412 36644
rect 19756 36604 19796 36644
rect 2380 36520 2420 36560
rect 6700 36520 6740 36560
rect 19948 36520 19988 36560
rect 6412 36436 6452 36476
rect 8908 36436 8948 36476
rect 10540 36436 10580 36476
rect 17260 36436 17300 36476
rect 3688 36268 3728 36308
rect 3770 36268 3810 36308
rect 3852 36268 3892 36308
rect 3934 36268 3974 36308
rect 4016 36268 4056 36308
rect 18808 36268 18848 36308
rect 18890 36268 18930 36308
rect 18972 36268 19012 36308
rect 19054 36268 19094 36308
rect 19136 36268 19176 36308
rect 1516 36100 1556 36140
rect 3436 36100 3476 36140
rect 4012 36100 4052 36140
rect 11596 36100 11636 36140
rect 12364 36100 12404 36140
rect 15052 36100 15092 36140
rect 16684 36100 16724 36140
rect 1324 35932 1364 35972
rect 3628 35932 3668 35972
rect 3820 35932 3860 35972
rect 6988 35932 7028 35972
rect 7084 35932 7124 35972
rect 11404 35932 11444 35972
rect 19948 35932 19988 35972
rect 4972 35848 5012 35888
rect 6220 35848 6260 35888
rect 6508 35848 6548 35888
rect 6604 35848 6644 35888
rect 7564 35848 7604 35888
rect 8044 35853 8084 35893
rect 9484 35848 9524 35888
rect 9580 35848 9620 35888
rect 9964 35848 10004 35888
rect 10060 35848 10100 35888
rect 10540 35848 10580 35888
rect 11020 35862 11060 35902
rect 11884 35848 11924 35888
rect 13132 35848 13172 35888
rect 13228 35848 13268 35888
rect 13612 35848 13652 35888
rect 14716 35890 14756 35930
rect 13708 35848 13748 35888
rect 14188 35848 14228 35888
rect 15244 35848 15284 35888
rect 16492 35848 16532 35888
rect 16876 35848 16916 35888
rect 18124 35848 18164 35888
rect 18316 35848 18356 35888
rect 19564 35848 19604 35888
rect 8236 35764 8276 35804
rect 2188 35680 2228 35720
rect 4492 35680 4532 35720
rect 4780 35680 4820 35720
rect 11212 35680 11252 35720
rect 14860 35680 14900 35720
rect 19756 35680 19796 35720
rect 20140 35680 20180 35720
rect 4928 35512 4968 35552
rect 5010 35512 5050 35552
rect 5092 35512 5132 35552
rect 5174 35512 5214 35552
rect 5256 35512 5296 35552
rect 20048 35512 20088 35552
rect 20130 35512 20170 35552
rect 20212 35512 20252 35552
rect 20294 35512 20334 35552
rect 20376 35512 20416 35552
rect 7564 35344 7604 35384
rect 3628 35260 3668 35300
rect 5644 35260 5684 35300
rect 19276 35260 19316 35300
rect 1900 35176 1940 35216
rect 1996 35176 2036 35216
rect 2476 35176 2516 35216
rect 2956 35176 2996 35216
rect 3436 35162 3476 35202
rect 3916 35176 3956 35216
rect 4012 35176 4052 35216
rect 4972 35176 5012 35216
rect 5452 35171 5492 35211
rect 6124 35176 6164 35216
rect 7372 35176 7412 35216
rect 7756 35176 7796 35216
rect 9004 35176 9044 35216
rect 9388 35176 9428 35216
rect 10636 35176 10676 35216
rect 11020 35176 11060 35216
rect 12268 35176 12308 35216
rect 12652 35176 12692 35216
rect 13900 35176 13940 35216
rect 15724 35176 15764 35216
rect 17548 35176 17588 35216
rect 1420 35092 1460 35132
rect 2380 35092 2420 35132
rect 4396 35092 4436 35132
rect 14476 35134 14516 35174
rect 17644 35176 17684 35216
rect 18028 35176 18068 35216
rect 18124 35176 18164 35216
rect 18604 35176 18644 35216
rect 19084 35171 19124 35211
rect 4492 35092 4532 35132
rect 15916 35092 15956 35132
rect 16300 35092 16340 35132
rect 16684 35092 16724 35132
rect 17068 35092 17108 35132
rect 19468 35092 19508 35132
rect 19852 35092 19892 35132
rect 1612 35008 1652 35048
rect 16108 35008 16148 35048
rect 16492 35008 16532 35048
rect 16876 35008 16916 35048
rect 17260 35008 17300 35048
rect 9196 34924 9236 34964
rect 10828 34924 10868 34964
rect 12460 34924 12500 34964
rect 14092 34924 14132 34964
rect 14284 34924 14324 34964
rect 19660 34924 19700 34964
rect 20044 34924 20084 34964
rect 3688 34756 3728 34796
rect 3770 34756 3810 34796
rect 3852 34756 3892 34796
rect 3934 34756 3974 34796
rect 4016 34756 4056 34796
rect 18808 34756 18848 34796
rect 18890 34756 18930 34796
rect 18972 34756 19012 34796
rect 19054 34756 19094 34796
rect 19136 34756 19176 34796
rect 2956 34588 2996 34628
rect 3148 34420 3188 34460
rect 3916 34420 3956 34460
rect 8428 34420 8468 34460
rect 13804 34420 13844 34460
rect 18604 34420 18644 34460
rect 18988 34420 19028 34460
rect 19372 34420 19412 34460
rect 19756 34420 19796 34460
rect 1228 34336 1268 34376
rect 2476 34336 2516 34376
rect 3340 34336 3380 34376
rect 3436 34336 3476 34376
rect 3628 34336 3668 34376
rect 4204 34336 4244 34376
rect 5452 34336 5492 34376
rect 6028 34336 6068 34376
rect 6220 34336 6260 34376
rect 7468 34336 7508 34376
rect 7948 34336 7988 34376
rect 8044 34336 8084 34376
rect 8524 34336 8564 34376
rect 9004 34336 9044 34376
rect 9484 34350 9524 34390
rect 11020 34336 11060 34376
rect 12268 34336 12308 34376
rect 13324 34336 13364 34376
rect 13420 34336 13460 34376
rect 13900 34336 13940 34376
rect 14380 34336 14420 34376
rect 14860 34350 14900 34390
rect 15244 34336 15284 34376
rect 16492 34336 16532 34376
rect 16876 34336 16916 34376
rect 18124 34336 18164 34376
rect 5644 34252 5684 34292
rect 7660 34252 7700 34292
rect 2668 34168 2708 34208
rect 3532 34168 3572 34208
rect 5932 34168 5972 34208
rect 9676 34168 9716 34208
rect 12460 34168 12500 34208
rect 15052 34168 15092 34208
rect 16684 34168 16724 34208
rect 18316 34168 18356 34208
rect 18796 34168 18836 34208
rect 19180 34168 19220 34208
rect 19564 34168 19604 34208
rect 19948 34168 19988 34208
rect 4928 34000 4968 34040
rect 5010 34000 5050 34040
rect 5092 34000 5132 34040
rect 5174 34000 5214 34040
rect 5256 34000 5296 34040
rect 20048 34000 20088 34040
rect 20130 34000 20170 34040
rect 20212 34000 20252 34040
rect 20294 34000 20334 34040
rect 20376 34000 20416 34040
rect 1612 33832 1652 33872
rect 3916 33832 3956 33872
rect 5644 33832 5684 33872
rect 5836 33832 5876 33872
rect 15724 33832 15764 33872
rect 17740 33832 17780 33872
rect 3628 33748 3668 33788
rect 9676 33748 9716 33788
rect 11692 33748 11732 33788
rect 14188 33748 14228 33788
rect 1900 33664 1940 33704
rect 1996 33664 2036 33704
rect 2476 33664 2516 33704
rect 2967 33651 3007 33691
rect 3436 33659 3476 33699
rect 4204 33664 4244 33704
rect 5452 33664 5492 33704
rect 6028 33664 6068 33704
rect 7276 33664 7316 33704
rect 7468 33664 7508 33704
rect 7852 33664 7892 33704
rect 8236 33664 8276 33704
rect 9484 33664 9524 33704
rect 9964 33664 10004 33704
rect 10060 33664 10100 33704
rect 10444 33664 10484 33704
rect 10540 33664 10580 33704
rect 11020 33664 11060 33704
rect 11500 33659 11540 33699
rect 12460 33664 12500 33704
rect 12556 33664 12596 33704
rect 13516 33664 13556 33704
rect 14044 33654 14084 33694
rect 16012 33664 16052 33704
rect 16108 33664 16148 33704
rect 17068 33664 17108 33704
rect 17548 33659 17588 33699
rect 1420 33580 1460 33620
rect 2380 33580 2420 33620
rect 7564 33580 7604 33620
rect 7756 33580 7796 33620
rect 12940 33580 12980 33620
rect 13036 33580 13076 33620
rect 15532 33580 15572 33620
rect 16492 33580 16532 33620
rect 16588 33580 16628 33620
rect 18220 33580 18260 33620
rect 18604 33580 18644 33620
rect 18988 33580 19028 33620
rect 19372 33580 19412 33620
rect 19756 33580 19796 33620
rect 7660 33496 7700 33536
rect 15340 33496 15380 33536
rect 19180 33496 19220 33536
rect 5644 33412 5684 33452
rect 18412 33412 18452 33452
rect 18796 33412 18836 33452
rect 19564 33412 19604 33452
rect 19948 33412 19988 33452
rect 3688 33244 3728 33284
rect 3770 33244 3810 33284
rect 3852 33244 3892 33284
rect 3934 33244 3974 33284
rect 4016 33244 4056 33284
rect 18808 33244 18848 33284
rect 18890 33244 18930 33284
rect 18972 33244 19012 33284
rect 19054 33244 19094 33284
rect 19136 33244 19176 33284
rect 1516 33076 1556 33116
rect 1900 33076 1940 33116
rect 5452 33076 5492 33116
rect 5836 33076 5876 33116
rect 7084 33076 7124 33116
rect 19564 33076 19604 33116
rect 2284 32992 2324 33032
rect 19948 32992 19988 33032
rect 1324 32908 1364 32948
rect 1708 32908 1748 32948
rect 11884 32908 11924 32948
rect 17740 32908 17780 32948
rect 19372 32908 19412 32948
rect 19756 32908 19796 32948
rect 2476 32824 2516 32864
rect 3724 32824 3764 32864
rect 4012 32824 4052 32864
rect 5260 32824 5300 32864
rect 6220 32824 6260 32864
rect 6508 32824 6548 32864
rect 6796 32824 6836 32864
rect 6892 32824 6932 32864
rect 7084 32824 7124 32864
rect 7276 32824 7316 32864
rect 7468 32824 7508 32864
rect 7564 32824 7604 32864
rect 7756 32824 7796 32864
rect 7852 32824 7892 32864
rect 8044 32824 8084 32864
rect 9292 32824 9332 32864
rect 10156 32824 10196 32864
rect 11404 32824 11444 32864
rect 12652 32824 12692 32864
rect 13324 32824 13364 32864
rect 14572 32824 14612 32864
rect 15436 32824 15476 32864
rect 16684 32824 16724 32864
rect 17164 32824 17204 32864
rect 17260 32824 17300 32864
rect 17644 32824 17684 32864
rect 18220 32824 18260 32864
rect 18748 32833 18788 32873
rect 6124 32740 6164 32780
rect 7372 32740 7412 32780
rect 16876 32740 16916 32780
rect 18892 32740 18932 32780
rect 9484 32656 9524 32696
rect 11596 32656 11636 32696
rect 14764 32656 14804 32696
rect 4928 32488 4968 32528
rect 5010 32488 5050 32528
rect 5092 32488 5132 32528
rect 5174 32488 5214 32528
rect 5256 32488 5296 32528
rect 20048 32488 20088 32528
rect 20130 32488 20170 32528
rect 20212 32488 20252 32528
rect 20294 32488 20334 32528
rect 20376 32488 20416 32528
rect 2764 32320 2804 32360
rect 4780 32320 4820 32360
rect 7852 32320 7892 32360
rect 8332 32320 8372 32360
rect 16492 32320 16532 32360
rect 16876 32320 16916 32360
rect 17260 32320 17300 32360
rect 18892 32320 18932 32360
rect 6892 32236 6932 32276
rect 12172 32236 12212 32276
rect 14188 32236 14228 32276
rect 2956 32147 2996 32187
rect 3436 32152 3476 32192
rect 4396 32152 4436 32192
rect 4492 32152 4532 32192
rect 4972 32152 5012 32192
rect 6220 32152 6260 32192
rect 6508 32152 6548 32192
rect 6796 32152 6836 32192
rect 7660 32152 7700 32192
rect 3916 32068 3956 32108
rect 4012 32068 4052 32108
rect 8044 32107 8084 32147
rect 8140 32152 8180 32192
rect 8236 32152 8276 32192
rect 8620 32152 8660 32192
rect 9868 32152 9908 32192
rect 10732 32152 10772 32192
rect 11980 32152 12020 32192
rect 12460 32152 12500 32192
rect 12556 32152 12596 32192
rect 13516 32152 13556 32192
rect 13996 32138 14036 32178
rect 14764 32152 14804 32192
rect 14860 32152 14900 32192
rect 15244 32152 15284 32192
rect 15340 32152 15380 32192
rect 15820 32152 15860 32192
rect 16300 32138 16340 32178
rect 17452 32152 17492 32192
rect 18700 32152 18740 32192
rect 12940 32068 12980 32108
rect 13036 32068 13076 32108
rect 16684 32068 16724 32108
rect 17068 32068 17108 32108
rect 19372 32068 19412 32108
rect 19756 32068 19796 32108
rect 7180 31984 7220 32024
rect 7660 31984 7700 32024
rect 10060 31900 10100 31940
rect 19564 31900 19604 31940
rect 19948 31900 19988 31940
rect 3688 31732 3728 31772
rect 3770 31732 3810 31772
rect 3852 31732 3892 31772
rect 3934 31732 3974 31772
rect 4016 31732 4056 31772
rect 18808 31732 18848 31772
rect 18890 31732 18930 31772
rect 18972 31732 19012 31772
rect 19054 31732 19094 31772
rect 19136 31732 19176 31772
rect 13996 31564 14036 31604
rect 16300 31564 16340 31604
rect 8236 31396 8276 31436
rect 10636 31396 10676 31436
rect 20044 31396 20084 31436
rect 1228 31312 1268 31352
rect 2476 31312 2516 31352
rect 3052 31312 3092 31352
rect 4204 31312 4244 31352
rect 4396 31312 4436 31352
rect 5644 31312 5684 31352
rect 6028 31312 6068 31352
rect 7276 31312 7316 31352
rect 7756 31312 7796 31352
rect 7852 31312 7892 31352
rect 8332 31312 8372 31352
rect 8812 31312 8852 31352
rect 9340 31321 9380 31361
rect 10060 31312 10100 31352
rect 10156 31312 10196 31352
rect 10540 31312 10580 31352
rect 11116 31312 11156 31352
rect 11596 31326 11636 31366
rect 12556 31312 12596 31352
rect 13804 31312 13844 31352
rect 14860 31312 14900 31352
rect 16108 31312 16148 31352
rect 16492 31312 16532 31352
rect 17740 31312 17780 31352
rect 18412 31312 18452 31352
rect 19660 31312 19700 31352
rect 7468 31228 7508 31268
rect 2668 31144 2708 31184
rect 3148 31144 3188 31184
rect 4108 31144 4148 31184
rect 5836 31144 5876 31184
rect 9484 31144 9524 31184
rect 11788 31144 11828 31184
rect 17932 31144 17972 31184
rect 19852 31144 19892 31184
rect 20236 31144 20276 31184
rect 4928 30976 4968 31016
rect 5010 30976 5050 31016
rect 5092 30976 5132 31016
rect 5174 30976 5214 31016
rect 5256 30976 5296 31016
rect 20048 30976 20088 31016
rect 20130 30976 20170 31016
rect 20212 30976 20252 31016
rect 20294 30976 20334 31016
rect 20376 30976 20416 31016
rect 6604 30808 6644 30848
rect 7084 30808 7124 30848
rect 7468 30808 7508 30848
rect 19468 30808 19508 30848
rect 4108 30724 4148 30764
rect 6124 30724 6164 30764
rect 2188 30640 2228 30680
rect 2380 30640 2420 30680
rect 2476 30640 2516 30680
rect 2668 30640 2708 30680
rect 3916 30640 3956 30680
rect 4396 30640 4436 30680
rect 4492 30640 4532 30680
rect 4876 30640 4916 30680
rect 4972 30640 5012 30680
rect 5452 30640 5492 30680
rect 5932 30635 5972 30675
rect 6316 30640 6356 30680
rect 6412 30640 6452 30680
rect 6508 30640 6548 30680
rect 6988 30640 7028 30680
rect 7180 30640 7220 30680
rect 7372 30640 7412 30680
rect 8908 30640 8948 30680
rect 10156 30640 10196 30680
rect 10828 30640 10868 30680
rect 12076 30640 12116 30680
rect 12460 30640 12500 30680
rect 13708 30640 13748 30680
rect 14092 30640 14132 30680
rect 15340 30640 15380 30680
rect 15724 30640 15764 30680
rect 16972 30640 17012 30680
rect 17740 30640 17780 30680
rect 17836 30640 17876 30680
rect 18220 30640 18260 30680
rect 18316 30640 18356 30680
rect 18796 30640 18836 30680
rect 19276 30635 19316 30675
rect 19660 30556 19700 30596
rect 20044 30556 20084 30596
rect 2284 30472 2324 30512
rect 10348 30388 10388 30428
rect 12268 30388 12308 30428
rect 13900 30388 13940 30428
rect 15532 30388 15572 30428
rect 17164 30388 17204 30428
rect 19852 30388 19892 30428
rect 20236 30388 20276 30428
rect 3688 30220 3728 30260
rect 3770 30220 3810 30260
rect 3852 30220 3892 30260
rect 3934 30220 3974 30260
rect 4016 30220 4056 30260
rect 18808 30220 18848 30260
rect 18890 30220 18930 30260
rect 18972 30220 19012 30260
rect 19054 30220 19094 30260
rect 19136 30220 19176 30260
rect 16684 30052 16724 30092
rect 2668 29968 2708 30008
rect 16300 29968 16340 30008
rect 7372 29884 7412 29924
rect 7468 29884 7508 29924
rect 11020 29884 11060 29924
rect 16108 29884 16148 29924
rect 16492 29884 16532 29924
rect 17644 29884 17684 29924
rect 1228 29800 1268 29840
rect 2476 29800 2516 29840
rect 2860 29800 2900 29840
rect 2956 29800 2996 29840
rect 3148 29800 3188 29840
rect 3244 29800 3284 29840
rect 3345 29800 3385 29840
rect 3628 29800 3668 29840
rect 3724 29800 3764 29840
rect 5164 29800 5204 29840
rect 6412 29800 6452 29840
rect 6892 29800 6932 29840
rect 6988 29800 7028 29840
rect 7948 29800 7988 29840
rect 8428 29805 8468 29845
rect 8812 29800 8852 29840
rect 9772 29800 9812 29840
rect 10444 29800 10484 29840
rect 10540 29800 10580 29840
rect 10924 29800 10964 29840
rect 11500 29800 11540 29840
rect 11980 29814 12020 29854
rect 13900 29800 13940 29840
rect 13996 29800 14036 29840
rect 14380 29800 14420 29840
rect 15484 29842 15524 29882
rect 19372 29884 19412 29924
rect 19756 29884 19796 29924
rect 14476 29800 14516 29840
rect 14956 29800 14996 29840
rect 17164 29800 17204 29840
rect 17260 29800 17300 29840
rect 18219 29842 18259 29882
rect 17740 29800 17780 29840
rect 18700 29805 18740 29845
rect 6604 29716 6644 29756
rect 8620 29716 8660 29756
rect 12172 29716 12212 29756
rect 15628 29716 15668 29756
rect 18892 29716 18932 29756
rect 3052 29632 3092 29672
rect 3916 29632 3956 29672
rect 19564 29632 19604 29672
rect 19948 29632 19988 29672
rect 4928 29464 4968 29504
rect 5010 29464 5050 29504
rect 5092 29464 5132 29504
rect 5174 29464 5214 29504
rect 5256 29464 5296 29504
rect 20048 29464 20088 29504
rect 20130 29464 20170 29504
rect 20212 29464 20252 29504
rect 20294 29464 20334 29504
rect 20376 29464 20416 29504
rect 8428 29296 8468 29336
rect 19948 29296 19988 29336
rect 1516 29128 1556 29168
rect 2764 29128 2804 29168
rect 3820 29128 3860 29168
rect 5068 29128 5108 29168
rect 6988 29128 7028 29168
rect 8236 29128 8276 29168
rect 8716 29128 8756 29168
rect 9964 29128 10004 29168
rect 10348 29128 10388 29168
rect 11596 29128 11636 29168
rect 11980 29128 12020 29168
rect 13228 29128 13268 29168
rect 13612 29128 13652 29168
rect 14860 29128 14900 29168
rect 15244 29128 15284 29168
rect 16492 29128 16532 29168
rect 17068 29128 17108 29168
rect 18316 29128 18356 29168
rect 18508 29128 18548 29168
rect 19756 29128 19796 29168
rect 2956 28876 2996 28916
rect 5260 28876 5300 28916
rect 10156 28876 10196 28916
rect 11788 28876 11828 28916
rect 13420 28876 13460 28916
rect 15052 28876 15092 28916
rect 16684 28876 16724 28916
rect 16876 28876 16916 28916
rect 3688 28708 3728 28748
rect 3770 28708 3810 28748
rect 3852 28708 3892 28748
rect 3934 28708 3974 28748
rect 4016 28708 4056 28748
rect 18808 28708 18848 28748
rect 18890 28708 18930 28748
rect 18972 28708 19012 28748
rect 19054 28708 19094 28748
rect 19136 28708 19176 28748
rect 10636 28372 10676 28412
rect 1900 28288 1940 28328
rect 3148 28288 3188 28328
rect 3628 28288 3668 28328
rect 3724 28288 3764 28328
rect 4108 28288 4148 28328
rect 4204 28288 4244 28328
rect 4684 28288 4724 28328
rect 5164 28302 5204 28342
rect 5932 28288 5972 28328
rect 7180 28288 7220 28328
rect 7756 28288 7796 28328
rect 9004 28288 9044 28328
rect 10156 28307 10196 28347
rect 10252 28288 10292 28328
rect 11740 28330 11780 28370
rect 13900 28372 13940 28412
rect 17068 28372 17108 28412
rect 19468 28372 19508 28412
rect 19852 28372 19892 28412
rect 10732 28288 10772 28328
rect 11212 28288 11252 28328
rect 13324 28288 13364 28328
rect 13420 28288 13460 28328
rect 14908 28330 14948 28370
rect 13804 28288 13844 28328
rect 14380 28288 14420 28328
rect 15244 28288 15284 28328
rect 16492 28288 16532 28328
rect 17548 28288 17588 28328
rect 17644 28288 17684 28328
rect 18028 28288 18068 28328
rect 18124 28288 18164 28328
rect 18604 28288 18644 28328
rect 19132 28297 19172 28337
rect 5356 28204 5396 28244
rect 11884 28204 11924 28244
rect 15052 28204 15092 28244
rect 3340 28120 3380 28160
rect 7372 28120 7412 28160
rect 9196 28120 9236 28160
rect 16684 28120 16724 28160
rect 17260 28120 17300 28160
rect 19276 28120 19316 28160
rect 19660 28120 19700 28160
rect 20044 28120 20084 28160
rect 4928 27952 4968 27992
rect 5010 27952 5050 27992
rect 5092 27952 5132 27992
rect 5174 27952 5214 27992
rect 5256 27952 5296 27992
rect 20048 27952 20088 27992
rect 20130 27952 20170 27992
rect 20212 27952 20252 27992
rect 20294 27952 20334 27992
rect 20376 27952 20416 27992
rect 19756 27784 19796 27824
rect 4204 27700 4244 27740
rect 7276 27700 7316 27740
rect 9292 27700 9332 27740
rect 12172 27700 12212 27740
rect 16492 27700 16532 27740
rect 2476 27616 2516 27656
rect 2572 27616 2612 27656
rect 2956 27616 2996 27656
rect 3532 27616 3572 27656
rect 4012 27611 4052 27651
rect 5548 27616 5588 27656
rect 5644 27616 5684 27656
rect 6604 27616 6644 27656
rect 7084 27602 7124 27642
rect 7564 27616 7604 27656
rect 7660 27616 7700 27656
rect 8044 27616 8084 27656
rect 8140 27616 8180 27656
rect 8620 27616 8660 27656
rect 9148 27606 9188 27646
rect 10444 27616 10484 27656
rect 10540 27616 10580 27656
rect 11020 27616 11060 27656
rect 11500 27616 11540 27656
rect 11980 27602 12020 27642
rect 13036 27616 13076 27656
rect 14284 27616 14324 27656
rect 14764 27616 14804 27656
rect 14860 27616 14900 27656
rect 15340 27616 15380 27656
rect 15820 27616 15860 27656
rect 16300 27611 16340 27651
rect 16684 27616 16724 27656
rect 17932 27616 17972 27656
rect 18316 27616 18356 27656
rect 19564 27616 19604 27656
rect 3052 27532 3092 27572
rect 6028 27532 6068 27572
rect 6124 27532 6164 27572
rect 10924 27532 10964 27572
rect 15244 27532 15284 27572
rect 19948 27532 19988 27572
rect 14476 27364 14516 27404
rect 18124 27364 18164 27404
rect 20140 27364 20180 27404
rect 3688 27196 3728 27236
rect 3770 27196 3810 27236
rect 3852 27196 3892 27236
rect 3934 27196 3974 27236
rect 4016 27196 4056 27236
rect 18808 27196 18848 27236
rect 18890 27196 18930 27236
rect 18972 27196 19012 27236
rect 19054 27196 19094 27236
rect 19136 27196 19176 27236
rect 2668 27028 2708 27068
rect 5932 27028 5972 27068
rect 7564 27028 7604 27068
rect 10348 27028 10388 27068
rect 18508 26944 18548 26984
rect 17164 26860 17204 26900
rect 1228 26776 1268 26816
rect 2476 26776 2516 26816
rect 2860 26776 2900 26816
rect 4108 26776 4148 26816
rect 4492 26776 4532 26816
rect 5740 26776 5780 26816
rect 6124 26776 6164 26816
rect 7372 26776 7412 26816
rect 8908 26776 8948 26816
rect 10156 26776 10196 26816
rect 10828 26776 10868 26816
rect 12076 26776 12116 26816
rect 13612 26776 13652 26816
rect 14860 26776 14900 26816
rect 16588 26776 16628 26816
rect 16684 26776 16724 26816
rect 17068 26776 17108 26816
rect 17644 26776 17684 26816
rect 18172 26785 18212 26825
rect 18700 26776 18740 26816
rect 19948 26776 19988 26816
rect 4300 26608 4340 26648
rect 12268 26608 12308 26648
rect 15052 26608 15092 26648
rect 18316 26608 18356 26648
rect 4928 26440 4968 26480
rect 5010 26440 5050 26480
rect 5092 26440 5132 26480
rect 5174 26440 5214 26480
rect 5256 26440 5296 26480
rect 20048 26440 20088 26480
rect 20130 26440 20170 26480
rect 20212 26440 20252 26480
rect 20294 26440 20334 26480
rect 20376 26440 20416 26480
rect 5068 26188 5108 26228
rect 19180 26188 19220 26228
rect 1612 26104 1652 26144
rect 2860 26104 2900 26144
rect 3340 26085 3380 26125
rect 3436 26104 3476 26144
rect 4396 26104 4436 26144
rect 4876 26099 4916 26139
rect 5452 26104 5492 26144
rect 6700 26104 6740 26144
rect 7084 26104 7124 26144
rect 8332 26104 8372 26144
rect 9196 26104 9236 26144
rect 10444 26104 10484 26144
rect 10828 26104 10868 26144
rect 12076 26104 12116 26144
rect 12460 26104 12500 26144
rect 13708 26104 13748 26144
rect 14860 26104 14900 26144
rect 16108 26104 16148 26144
rect 17452 26104 17492 26144
rect 17548 26104 17588 26144
rect 18508 26104 18548 26144
rect 3820 26020 3860 26060
rect 3916 26020 3956 26060
rect 17932 26020 17972 26060
rect 18028 26020 18068 26060
rect 19036 26062 19076 26102
rect 19372 26020 19412 26060
rect 19756 26020 19796 26060
rect 3052 25852 3092 25892
rect 6892 25852 6932 25892
rect 8524 25852 8564 25892
rect 10636 25852 10676 25892
rect 12268 25852 12308 25892
rect 13900 25852 13940 25892
rect 16300 25852 16340 25892
rect 19564 25852 19604 25892
rect 19948 25852 19988 25892
rect 3688 25684 3728 25724
rect 3770 25684 3810 25724
rect 3852 25684 3892 25724
rect 3934 25684 3974 25724
rect 4016 25684 4056 25724
rect 18808 25684 18848 25724
rect 18890 25684 18930 25724
rect 18972 25684 19012 25724
rect 19054 25684 19094 25724
rect 19136 25684 19176 25724
rect 3148 25516 3188 25556
rect 19468 25516 19508 25556
rect 19852 25432 19892 25472
rect 4204 25348 4244 25388
rect 4300 25348 4340 25388
rect 11404 25348 11444 25388
rect 19660 25348 19700 25388
rect 20044 25348 20084 25388
rect 1708 25264 1748 25304
rect 2956 25264 2996 25304
rect 3724 25264 3764 25304
rect 3820 25264 3860 25304
rect 4780 25264 4820 25304
rect 5308 25273 5348 25313
rect 7084 25263 7124 25303
rect 7180 25264 7220 25304
rect 7564 25264 7604 25304
rect 7660 25264 7700 25304
rect 8140 25264 8180 25304
rect 8620 25278 8660 25318
rect 9100 25264 9140 25304
rect 10348 25264 10388 25304
rect 10828 25264 10868 25304
rect 10924 25264 10964 25304
rect 11308 25264 11348 25304
rect 11884 25264 11924 25304
rect 12364 25278 12404 25318
rect 13708 25264 13748 25304
rect 13804 25264 13844 25304
rect 14188 25264 14228 25304
rect 14284 25264 14324 25304
rect 14764 25264 14804 25304
rect 15244 25278 15284 25318
rect 16396 25264 16436 25304
rect 17644 25264 17684 25304
rect 18028 25264 18068 25304
rect 19276 25264 19316 25304
rect 5452 25180 5492 25220
rect 8812 25180 8852 25220
rect 10540 25180 10580 25220
rect 12556 25096 12596 25136
rect 15436 25096 15476 25136
rect 17836 25096 17876 25136
rect 20236 25096 20276 25136
rect 4928 24928 4968 24968
rect 5010 24928 5050 24968
rect 5092 24928 5132 24968
rect 5174 24928 5214 24968
rect 5256 24928 5296 24968
rect 20048 24928 20088 24968
rect 20130 24928 20170 24968
rect 20212 24928 20252 24968
rect 20294 24928 20334 24968
rect 20376 24928 20416 24968
rect 3148 24760 3188 24800
rect 5068 24760 5108 24800
rect 11692 24760 11732 24800
rect 18796 24760 18836 24800
rect 6700 24676 6740 24716
rect 9676 24676 9716 24716
rect 18220 24676 18260 24716
rect 1228 24592 1268 24632
rect 2476 24592 2516 24632
rect 2860 24592 2900 24632
rect 2956 24592 2996 24632
rect 3628 24592 3668 24632
rect 4876 24592 4916 24632
rect 5260 24592 5300 24632
rect 6508 24592 6548 24632
rect 7180 24592 7220 24632
rect 7468 24592 7508 24632
rect 7564 24592 7604 24632
rect 8236 24592 8276 24632
rect 9484 24592 9524 24632
rect 9964 24592 10004 24632
rect 10060 24592 10100 24632
rect 11020 24592 11060 24632
rect 11500 24587 11540 24627
rect 13900 24592 13940 24632
rect 15148 24592 15188 24632
rect 16492 24592 16532 24632
rect 16588 24592 16628 24632
rect 17548 24592 17588 24632
rect 18028 24587 18068 24627
rect 10444 24508 10484 24548
rect 10540 24508 10580 24548
rect 16972 24508 17012 24548
rect 17068 24508 17108 24548
rect 18604 24508 18644 24548
rect 18988 24508 19028 24548
rect 19372 24508 19412 24548
rect 19756 24505 19796 24545
rect 2668 24340 2708 24380
rect 7852 24340 7892 24380
rect 15340 24340 15380 24380
rect 19180 24340 19220 24380
rect 19564 24340 19604 24380
rect 19948 24340 19988 24380
rect 3688 24172 3728 24212
rect 3770 24172 3810 24212
rect 3852 24172 3892 24212
rect 3934 24172 3974 24212
rect 4016 24172 4056 24212
rect 18808 24172 18848 24212
rect 18890 24172 18930 24212
rect 18972 24172 19012 24212
rect 19054 24172 19094 24212
rect 19136 24172 19176 24212
rect 2668 24004 2708 24044
rect 15916 23920 15956 23960
rect 1228 23752 1268 23792
rect 2476 23752 2516 23792
rect 2860 23731 2900 23771
rect 2956 23752 2996 23792
rect 3052 23752 3092 23792
rect 3340 23797 3380 23837
rect 4012 23836 4052 23876
rect 11308 23836 11348 23876
rect 3436 23794 3476 23834
rect 14380 23836 14420 23876
rect 15724 23836 15764 23876
rect 18412 23836 18452 23876
rect 3532 23752 3572 23792
rect 4492 23752 4532 23792
rect 4588 23752 4628 23792
rect 4684 23752 4724 23792
rect 5068 23752 5108 23792
rect 5164 23752 5204 23792
rect 5356 23752 5396 23792
rect 5644 23752 5684 23792
rect 6892 23752 6932 23792
rect 7276 23752 7316 23792
rect 8524 23752 8564 23792
rect 9004 23752 9044 23792
rect 10252 23752 10292 23792
rect 10732 23751 10772 23791
rect 10828 23752 10868 23792
rect 11212 23752 11252 23792
rect 11788 23752 11828 23792
rect 12268 23757 12308 23797
rect 13804 23752 13844 23792
rect 13900 23752 13940 23792
rect 14284 23752 14324 23792
rect 14860 23752 14900 23792
rect 15340 23766 15380 23806
rect 16108 23752 16148 23792
rect 17356 23752 17396 23792
rect 17836 23752 17876 23792
rect 17932 23752 17972 23792
rect 18316 23752 18356 23792
rect 18892 23752 18932 23792
rect 19420 23761 19460 23801
rect 10444 23668 10484 23708
rect 17548 23668 17588 23708
rect 3148 23584 3188 23624
rect 3628 23584 3668 23624
rect 3820 23584 3860 23624
rect 4876 23584 4916 23624
rect 5260 23584 5300 23624
rect 7084 23584 7124 23624
rect 8716 23584 8756 23624
rect 12460 23584 12500 23624
rect 15532 23584 15572 23624
rect 19564 23584 19604 23624
rect 4928 23416 4968 23456
rect 5010 23416 5050 23456
rect 5092 23416 5132 23456
rect 5174 23416 5214 23456
rect 5256 23416 5296 23456
rect 20048 23416 20088 23456
rect 20130 23416 20170 23456
rect 20212 23416 20252 23456
rect 20294 23416 20334 23456
rect 20376 23416 20416 23456
rect 9004 23248 9044 23288
rect 9772 23248 9812 23288
rect 12172 23248 12212 23288
rect 13804 23248 13844 23288
rect 19756 23248 19796 23288
rect 2860 23164 2900 23204
rect 4972 23164 5012 23204
rect 8332 23164 8372 23204
rect 1420 23080 1460 23120
rect 2668 23080 2708 23120
rect 3244 23080 3284 23120
rect 3340 23080 3380 23120
rect 3820 23080 3860 23120
rect 4300 23080 4340 23120
rect 4780 23066 4820 23106
rect 5164 23080 5204 23120
rect 5260 23080 5300 23120
rect 5356 23080 5396 23120
rect 5452 23080 5492 23120
rect 5644 23080 5684 23120
rect 5932 23080 5972 23120
rect 6124 23080 6164 23120
rect 6316 23080 6356 23120
rect 6604 23080 6644 23120
rect 6700 23080 6740 23120
rect 7660 23080 7700 23120
rect 8140 23075 8180 23115
rect 8524 23080 8564 23120
rect 8620 23080 8660 23120
rect 8716 23080 8756 23120
rect 8812 23080 8852 23120
rect 9196 23080 9236 23120
rect 9292 23080 9332 23120
rect 9484 23080 9524 23120
rect 9580 23080 9620 23120
rect 9676 23080 9716 23120
rect 10732 23080 10772 23120
rect 11980 23080 12020 23120
rect 12364 23080 12404 23120
rect 13612 23080 13652 23120
rect 18316 23080 18356 23120
rect 19564 23080 19604 23120
rect 3724 22996 3764 23036
rect 7084 22996 7124 23036
rect 7180 22996 7220 23036
rect 19948 22996 19988 23036
rect 5644 22828 5684 22868
rect 6220 22828 6260 22868
rect 20140 22828 20180 22868
rect 3688 22660 3728 22700
rect 3770 22660 3810 22700
rect 3852 22660 3892 22700
rect 3934 22660 3974 22700
rect 4016 22660 4056 22700
rect 18808 22660 18848 22700
rect 18890 22660 18930 22700
rect 18972 22660 19012 22700
rect 19054 22660 19094 22700
rect 19136 22660 19176 22700
rect 4492 22492 4532 22532
rect 7948 22492 7988 22532
rect 19948 22492 19988 22532
rect 4684 22408 4724 22448
rect 10540 22324 10580 22364
rect 18988 22324 19028 22364
rect 19372 22324 19412 22364
rect 19756 22324 19796 22364
rect 1420 22240 1460 22280
rect 2668 22240 2708 22280
rect 3052 22240 3092 22280
rect 4300 22240 4340 22280
rect 4972 22240 5012 22280
rect 5068 22240 5108 22280
rect 5356 22240 5396 22280
rect 6988 22240 7028 22280
rect 7084 22240 7124 22280
rect 7660 22240 7700 22280
rect 7756 22240 7796 22280
rect 8236 22240 8276 22280
rect 9484 22240 9524 22280
rect 9964 22240 10004 22280
rect 10060 22240 10100 22280
rect 10444 22240 10484 22280
rect 11020 22253 11060 22293
rect 11500 22245 11540 22285
rect 11884 22240 11924 22280
rect 13132 22240 13172 22280
rect 13516 22240 13556 22280
rect 14764 22261 14804 22301
rect 15244 22240 15284 22280
rect 16492 22240 16532 22280
rect 17164 22240 17204 22280
rect 18412 22240 18452 22280
rect 2860 22156 2900 22196
rect 9676 22156 9716 22196
rect 11692 22156 11732 22196
rect 7276 22072 7316 22112
rect 7660 22072 7700 22112
rect 13324 22072 13364 22112
rect 14956 22072 14996 22112
rect 16684 22072 16724 22112
rect 18604 22072 18644 22112
rect 19180 22072 19220 22112
rect 19564 22072 19604 22112
rect 4928 21904 4968 21944
rect 5010 21904 5050 21944
rect 5092 21904 5132 21944
rect 5174 21904 5214 21944
rect 5256 21904 5296 21944
rect 20048 21904 20088 21944
rect 20130 21904 20170 21944
rect 20212 21904 20252 21944
rect 20294 21904 20334 21944
rect 20376 21904 20416 21944
rect 7084 21736 7124 21776
rect 9196 21736 9236 21776
rect 11308 21736 11348 21776
rect 14572 21652 14612 21692
rect 18700 21652 18740 21692
rect 3244 21568 3284 21608
rect 3340 21568 3380 21608
rect 3628 21568 3668 21608
rect 4012 21568 4052 21608
rect 5260 21568 5300 21608
rect 5644 21568 5684 21608
rect 6892 21568 6932 21608
rect 7468 21568 7508 21608
rect 7564 21568 7604 21608
rect 7948 21568 7988 21608
rect 8044 21568 8084 21608
rect 8524 21568 8564 21608
rect 9004 21554 9044 21594
rect 9868 21568 9908 21608
rect 11116 21568 11156 21608
rect 12460 21568 12500 21608
rect 12844 21568 12884 21608
rect 12940 21568 12980 21608
rect 13324 21568 13364 21608
rect 13420 21568 13460 21608
rect 13900 21568 13940 21608
rect 14380 21558 14420 21598
rect 14860 21568 14900 21608
rect 16108 21568 16148 21608
rect 16972 21568 17012 21608
rect 17068 21568 17108 21608
rect 17452 21568 17492 21608
rect 18028 21568 18068 21608
rect 18556 21558 18596 21598
rect 17548 21484 17588 21524
rect 18988 21484 19028 21524
rect 19372 21484 19412 21524
rect 16300 21400 16340 21440
rect 19564 21400 19604 21440
rect 2956 21316 2996 21356
rect 5452 21316 5492 21356
rect 12556 21316 12596 21356
rect 19180 21316 19220 21356
rect 3688 21148 3728 21188
rect 3770 21148 3810 21188
rect 3852 21148 3892 21188
rect 3934 21148 3974 21188
rect 4016 21148 4056 21188
rect 18808 21148 18848 21188
rect 18890 21148 18930 21188
rect 18972 21148 19012 21188
rect 19054 21148 19094 21188
rect 19136 21148 19176 21188
rect 9484 20980 9524 21020
rect 4588 20812 4628 20852
rect 4684 20812 4724 20852
rect 15340 20812 15380 20852
rect 18124 20812 18164 20852
rect 19468 20812 19508 20852
rect 19852 20812 19892 20852
rect 1612 20728 1652 20768
rect 2860 20728 2900 20768
rect 3628 20733 3668 20773
rect 4108 20728 4148 20768
rect 5068 20728 5108 20768
rect 5164 20728 5204 20768
rect 6124 20728 6164 20768
rect 6220 20728 6260 20768
rect 6604 20728 6644 20768
rect 6700 20728 6740 20768
rect 7180 20728 7220 20768
rect 7660 20733 7700 20773
rect 8044 20728 8084 20768
rect 9292 20728 9332 20768
rect 11020 20728 11060 20768
rect 12268 20728 12308 20768
rect 12652 20728 12692 20768
rect 12844 20728 12884 20768
rect 12940 20728 12980 20768
rect 13132 20728 13172 20768
rect 14380 20728 14420 20768
rect 14860 20728 14900 20768
rect 14956 20728 14996 20768
rect 15436 20728 15476 20768
rect 15916 20728 15956 20768
rect 16396 20742 16436 20782
rect 17548 20728 17588 20768
rect 17644 20728 17684 20768
rect 18028 20728 18068 20768
rect 18604 20728 18644 20768
rect 19132 20737 19172 20777
rect 3052 20644 3092 20684
rect 3436 20644 3476 20684
rect 14572 20644 14612 20684
rect 16588 20644 16628 20684
rect 7852 20560 7892 20600
rect 12460 20560 12500 20600
rect 12748 20560 12788 20600
rect 19276 20560 19316 20600
rect 19660 20560 19700 20600
rect 20044 20560 20084 20600
rect 4928 20392 4968 20432
rect 5010 20392 5050 20432
rect 5092 20392 5132 20432
rect 5174 20392 5214 20432
rect 5256 20392 5296 20432
rect 20048 20392 20088 20432
rect 20130 20392 20170 20432
rect 20212 20392 20252 20432
rect 20294 20392 20334 20432
rect 20376 20392 20416 20432
rect 12172 20224 12212 20264
rect 15436 20224 15476 20264
rect 17260 20224 17300 20264
rect 6796 20140 6836 20180
rect 10444 20140 10484 20180
rect 19660 20140 19700 20180
rect 1516 20056 1556 20096
rect 2764 20056 2804 20096
rect 3244 20056 3284 20096
rect 3340 20056 3380 20096
rect 3532 20056 3572 20096
rect 3916 20056 3956 20096
rect 4012 20056 4052 20096
rect 4108 20056 4148 20096
rect 4396 20056 4436 20096
rect 4588 20056 4628 20096
rect 4684 20056 4724 20096
rect 5356 20056 5396 20096
rect 6604 20056 6644 20096
rect 6988 20056 7028 20096
rect 8236 20056 8276 20096
rect 8716 20056 8756 20096
rect 8812 20056 8852 20096
rect 9196 20056 9236 20096
rect 9772 20056 9812 20096
rect 10732 20056 10772 20096
rect 11980 20056 12020 20096
rect 12455 20056 12495 20096
rect 12556 20056 12596 20096
rect 9292 19972 9332 20012
rect 10300 20014 10340 20054
rect 12652 20056 12692 20096
rect 12844 20056 12884 20096
rect 12940 20056 12980 20096
rect 13708 20056 13748 20096
rect 14956 20056 14996 20096
rect 15148 20056 15188 20096
rect 15244 20056 15284 20096
rect 15820 20056 15860 20096
rect 17068 20056 17108 20096
rect 18220 20056 18260 20096
rect 19468 20056 19508 20096
rect 19852 19972 19892 20012
rect 2956 19888 2996 19928
rect 8428 19888 8468 19928
rect 20044 19888 20084 19928
rect 3724 19804 3764 19844
rect 4396 19804 4436 19844
rect 12940 19804 12980 19844
rect 13516 19804 13556 19844
rect 3688 19636 3728 19676
rect 3770 19636 3810 19676
rect 3852 19636 3892 19676
rect 3934 19636 3974 19676
rect 4016 19636 4056 19676
rect 18808 19636 18848 19676
rect 18890 19636 18930 19676
rect 18972 19636 19012 19676
rect 19054 19636 19094 19676
rect 19136 19636 19176 19676
rect 2668 19468 2708 19508
rect 10348 19468 10388 19508
rect 15052 19468 15092 19508
rect 19564 19468 19604 19508
rect 17548 19300 17588 19340
rect 18988 19300 19028 19340
rect 19372 19300 19412 19340
rect 19756 19300 19796 19340
rect 1228 19216 1268 19256
rect 2476 19216 2516 19256
rect 3724 19216 3764 19256
rect 3820 19216 3860 19256
rect 3916 19216 3956 19256
rect 4108 19216 4148 19256
rect 5356 19216 5396 19256
rect 7276 19216 7316 19256
rect 8524 19216 8564 19256
rect 8908 19216 8948 19256
rect 10156 19216 10196 19256
rect 11596 19216 11636 19256
rect 12844 19216 12884 19256
rect 13228 19226 13268 19266
rect 13324 19216 13364 19256
rect 13900 19216 13940 19256
rect 14284 19216 14324 19256
rect 14380 19216 14420 19256
rect 14668 19216 14708 19256
rect 14764 19216 14804 19256
rect 15244 19216 15284 19256
rect 16492 19216 16532 19256
rect 16972 19216 17012 19256
rect 17068 19216 17108 19256
rect 17452 19216 17492 19256
rect 18028 19216 18068 19256
rect 18556 19225 18596 19265
rect 13804 19132 13844 19172
rect 16684 19132 16724 19172
rect 18700 19132 18740 19172
rect 3628 19048 3668 19088
rect 5548 19048 5588 19088
rect 8716 19048 8756 19088
rect 13036 19048 13076 19088
rect 13516 19048 13556 19088
rect 14092 19048 14132 19088
rect 19180 19048 19220 19088
rect 19948 19048 19988 19088
rect 14572 18990 14612 19030
rect 4928 18880 4968 18920
rect 5010 18880 5050 18920
rect 5092 18880 5132 18920
rect 5174 18880 5214 18920
rect 5256 18880 5296 18920
rect 20048 18880 20088 18920
rect 20130 18880 20170 18920
rect 20212 18880 20252 18920
rect 20294 18880 20334 18920
rect 20376 18880 20416 18920
rect 4204 18712 4244 18752
rect 13324 18712 13364 18752
rect 14956 18712 14996 18752
rect 15628 18712 15668 18752
rect 7180 18628 7220 18668
rect 11308 18628 11348 18668
rect 17452 18628 17492 18668
rect 19468 18628 19508 18668
rect 2476 18544 2516 18584
rect 2572 18544 2612 18584
rect 3532 18544 3572 18584
rect 4012 18530 4052 18570
rect 5452 18544 5492 18584
rect 5548 18544 5588 18584
rect 6508 18544 6548 18584
rect 6988 18530 7028 18570
rect 7468 18544 7508 18584
rect 8236 18544 8276 18584
rect 9484 18544 9524 18584
rect 9868 18544 9908 18584
rect 11116 18544 11156 18584
rect 11596 18544 11636 18584
rect 11692 18544 11732 18584
rect 12076 18544 12116 18584
rect 12652 18544 12692 18584
rect 13132 18539 13172 18579
rect 13516 18544 13556 18584
rect 14764 18544 14804 18584
rect 15148 18544 15188 18584
rect 15244 18544 15284 18584
rect 15436 18544 15476 18584
rect 15532 18544 15572 18584
rect 15633 18544 15673 18584
rect 16012 18544 16052 18584
rect 17260 18544 17300 18584
rect 17740 18544 17780 18584
rect 17836 18544 17876 18584
rect 18220 18544 18260 18584
rect 18796 18544 18836 18584
rect 19276 18530 19316 18570
rect 2956 18460 2996 18500
rect 3052 18460 3092 18500
rect 5932 18460 5972 18500
rect 6028 18460 6068 18500
rect 12172 18460 12212 18500
rect 18316 18460 18356 18500
rect 19660 18460 19700 18500
rect 20044 18460 20084 18500
rect 19852 18376 19892 18416
rect 7372 18292 7412 18332
rect 9676 18292 9716 18332
rect 14956 18292 14996 18332
rect 20236 18292 20276 18332
rect 3688 18124 3728 18164
rect 3770 18124 3810 18164
rect 3852 18124 3892 18164
rect 3934 18124 3974 18164
rect 4016 18124 4056 18164
rect 18808 18124 18848 18164
rect 18890 18124 18930 18164
rect 18972 18124 19012 18164
rect 19054 18124 19094 18164
rect 19136 18124 19176 18164
rect 4012 17956 4052 17996
rect 6700 17956 6740 17996
rect 16012 17956 16052 17996
rect 18700 17956 18740 17996
rect 19084 17872 19124 17912
rect 7660 17788 7700 17828
rect 9676 17788 9716 17828
rect 15244 17788 15284 17828
rect 2572 17704 2612 17744
rect 3820 17704 3860 17744
rect 5260 17704 5300 17744
rect 6508 17704 6548 17744
rect 7180 17704 7220 17744
rect 7276 17704 7316 17744
rect 7756 17704 7796 17744
rect 8236 17704 8276 17744
rect 8764 17713 8804 17753
rect 9196 17704 9236 17744
rect 9292 17704 9332 17744
rect 9772 17704 9812 17744
rect 10252 17704 10292 17744
rect 10732 17718 10772 17758
rect 13708 17704 13748 17744
rect 13804 17704 13844 17744
rect 14188 17713 14228 17753
rect 14668 17704 14708 17744
rect 15148 17704 15188 17744
rect 15628 17704 15668 17744
rect 15724 17704 15764 17744
rect 16012 17704 16052 17744
rect 16204 17704 16244 17744
rect 16300 17723 16340 17763
rect 17260 17704 17300 17744
rect 18508 17704 18548 17744
rect 19468 17704 19508 17744
rect 19756 17704 19796 17744
rect 13996 17620 14036 17660
rect 19372 17620 19412 17660
rect 8908 17536 8948 17576
rect 10924 17536 10964 17576
rect 4928 17368 4968 17408
rect 5010 17368 5050 17408
rect 5092 17368 5132 17408
rect 5174 17368 5214 17408
rect 5256 17368 5296 17408
rect 20048 17368 20088 17408
rect 20130 17368 20170 17408
rect 20212 17368 20252 17408
rect 20294 17368 20334 17408
rect 20376 17368 20416 17408
rect 2668 17200 2708 17240
rect 5548 17200 5588 17240
rect 7180 17200 7220 17240
rect 8908 17200 8948 17240
rect 11404 17200 11444 17240
rect 13420 17200 13460 17240
rect 15436 17200 15476 17240
rect 19852 17200 19892 17240
rect 13708 17116 13748 17156
rect 17548 17116 17588 17156
rect 1228 17032 1268 17072
rect 2476 17032 2516 17072
rect 3052 17032 3092 17072
rect 3340 17032 3380 17072
rect 3532 17032 3572 17072
rect 4780 17032 4820 17072
rect 5260 17032 5300 17072
rect 5356 17032 5396 17072
rect 5740 17032 5780 17072
rect 6988 17032 7028 17072
rect 8716 17032 8756 17072
rect 9964 17032 10004 17072
rect 11212 17032 11252 17072
rect 11692 17032 11732 17072
rect 7468 16990 7508 17030
rect 11788 17032 11828 17072
rect 12748 17032 12788 17072
rect 13228 17018 13268 17058
rect 13900 17032 13940 17072
rect 15148 17032 15188 17072
rect 15340 17032 15380 17072
rect 15532 17032 15572 17072
rect 15628 17032 15668 17072
rect 15916 17032 15956 17072
rect 17164 17032 17204 17072
rect 17740 17032 17780 17072
rect 12172 16948 12212 16988
rect 17644 16990 17684 17030
rect 17836 17032 17876 17072
rect 19660 17032 19700 17072
rect 18412 16990 18452 17030
rect 12268 16948 12308 16988
rect 18028 16948 18068 16988
rect 20044 16948 20084 16988
rect 20236 16864 20276 16904
rect 3340 16780 3380 16820
rect 4972 16780 5012 16820
rect 17356 16780 17396 16820
rect 18220 16780 18260 16820
rect 3688 16612 3728 16652
rect 3770 16612 3810 16652
rect 3852 16612 3892 16652
rect 3934 16612 3974 16652
rect 4016 16612 4056 16652
rect 18808 16612 18848 16652
rect 18890 16612 18930 16652
rect 18972 16612 19012 16652
rect 19054 16612 19094 16652
rect 19136 16612 19176 16652
rect 2860 16444 2900 16484
rect 13324 16444 13364 16484
rect 16876 16444 16916 16484
rect 6700 16360 6740 16400
rect 15916 16360 15956 16400
rect 17068 16360 17108 16400
rect 19660 16360 19700 16400
rect 3820 16276 3860 16316
rect 3916 16276 3956 16316
rect 1420 16192 1460 16232
rect 2668 16192 2708 16232
rect 3340 16192 3380 16232
rect 3436 16192 3476 16232
rect 4396 16192 4436 16232
rect 4876 16206 4916 16246
rect 5260 16192 5300 16232
rect 6508 16192 6548 16232
rect 6892 16192 6932 16232
rect 6988 16192 7028 16232
rect 7180 16192 7220 16232
rect 7276 16192 7316 16232
rect 7377 16192 7417 16232
rect 7852 16192 7892 16232
rect 9100 16192 9140 16232
rect 9484 16192 9524 16232
rect 10732 16192 10772 16232
rect 11884 16192 11924 16232
rect 13132 16192 13172 16232
rect 15436 16192 15476 16232
rect 15532 16192 15572 16232
rect 15724 16192 15764 16232
rect 15916 16192 15956 16232
rect 16204 16192 16244 16232
rect 16492 16192 16532 16232
rect 16588 16192 16628 16232
rect 16684 16192 16724 16232
rect 17452 16192 17492 16232
rect 17740 16192 17780 16232
rect 18220 16192 18260 16232
rect 19468 16192 19508 16232
rect 19948 16192 19988 16232
rect 20044 16192 20084 16232
rect 20140 16171 20180 16211
rect 5068 16108 5108 16148
rect 15628 16108 15668 16148
rect 17356 16108 17396 16148
rect 2860 16024 2900 16064
rect 7084 16024 7124 16064
rect 9292 16024 9332 16064
rect 10924 16024 10964 16064
rect 19852 16024 19892 16064
rect 4928 15856 4968 15896
rect 5010 15856 5050 15896
rect 5092 15856 5132 15896
rect 5174 15856 5214 15896
rect 5256 15856 5296 15896
rect 20048 15856 20088 15896
rect 20130 15856 20170 15896
rect 20212 15856 20252 15896
rect 20294 15856 20334 15896
rect 20376 15856 20416 15896
rect 2668 15688 2708 15728
rect 4204 15688 4244 15728
rect 4588 15688 4628 15728
rect 12556 15688 12596 15728
rect 15916 15688 15956 15728
rect 17932 15688 17972 15728
rect 20236 15688 20276 15728
rect 9676 15604 9716 15644
rect 1228 15520 1268 15560
rect 2476 15520 2516 15560
rect 3052 15520 3092 15560
rect 3148 15520 3188 15560
rect 3244 15520 3284 15560
rect 3628 15520 3668 15560
rect 3820 15520 3860 15560
rect 3916 15520 3956 15560
rect 4108 15520 4148 15560
rect 4300 15520 4340 15560
rect 4396 15520 4436 15560
rect 4780 15520 4820 15560
rect 6028 15520 6068 15560
rect 6220 15520 6260 15560
rect 7468 15520 7508 15560
rect 7948 15520 7988 15560
rect 8044 15520 8084 15560
rect 8428 15520 8468 15560
rect 8524 15520 8564 15560
rect 9004 15520 9044 15560
rect 9484 15515 9524 15555
rect 10828 15520 10868 15560
rect 10924 15520 10964 15560
rect 11404 15520 11444 15560
rect 11884 15520 11924 15560
rect 12364 15506 12404 15546
rect 12748 15520 12788 15560
rect 13996 15520 14036 15560
rect 14476 15520 14516 15560
rect 15724 15520 15764 15560
rect 16204 15520 16244 15560
rect 16300 15520 16340 15560
rect 16780 15520 16820 15560
rect 17260 15520 17300 15560
rect 17788 15510 17828 15550
rect 18508 15520 18548 15560
rect 18604 15520 18644 15560
rect 18988 15520 19028 15560
rect 19564 15520 19604 15560
rect 20044 15506 20084 15546
rect 11308 15436 11348 15476
rect 16684 15436 16724 15476
rect 19084 15436 19124 15476
rect 3436 15268 3476 15308
rect 3628 15268 3668 15308
rect 7660 15268 7700 15308
rect 14188 15268 14228 15308
rect 3688 15100 3728 15140
rect 3770 15100 3810 15140
rect 3852 15100 3892 15140
rect 3934 15100 3974 15140
rect 4016 15100 4056 15140
rect 18808 15100 18848 15140
rect 18890 15100 18930 15140
rect 18972 15100 19012 15140
rect 19054 15100 19094 15140
rect 19136 15100 19176 15140
rect 2860 14932 2900 14972
rect 7660 14932 7700 14972
rect 12172 14932 12212 14972
rect 13804 14932 13844 14972
rect 16780 14932 16820 14972
rect 19084 14932 19124 14972
rect 19756 14932 19796 14972
rect 19948 14932 19988 14972
rect 12940 14848 12980 14888
rect 8620 14764 8660 14804
rect 1228 14680 1268 14720
rect 2476 14680 2516 14720
rect 3244 14680 3284 14720
rect 3532 14680 3572 14720
rect 3916 14680 3956 14720
rect 4012 14680 4052 14720
rect 4108 14680 4148 14720
rect 4396 14680 4436 14720
rect 5644 14680 5684 14720
rect 6220 14680 6260 14720
rect 7468 14680 7508 14720
rect 8044 14680 8084 14720
rect 8140 14680 8180 14720
rect 8524 14680 8564 14720
rect 9100 14680 9140 14720
rect 9580 14694 9620 14734
rect 10732 14680 10772 14720
rect 11980 14680 12020 14720
rect 12652 14680 12692 14720
rect 12748 14680 12788 14720
rect 12940 14680 12980 14720
rect 13228 14680 13268 14720
rect 13324 14680 13364 14720
rect 13420 14680 13460 14720
rect 14188 14680 14228 14720
rect 14476 14680 14516 14720
rect 14764 14680 14804 14720
rect 14860 14680 14900 14720
rect 14956 14680 14996 14720
rect 15052 14680 15092 14720
rect 15340 14680 15380 14720
rect 16588 14680 16628 14720
rect 17644 14680 17684 14720
rect 18892 14680 18932 14720
rect 19372 14680 19412 14720
rect 19468 14680 19508 14720
rect 19564 14680 19604 14720
rect 19948 14680 19988 14720
rect 20140 14694 20180 14734
rect 20236 14680 20276 14720
rect 3148 14596 3188 14636
rect 3820 14596 3860 14636
rect 14092 14596 14132 14636
rect 2668 14512 2708 14552
rect 5836 14512 5876 14552
rect 9772 14512 9812 14552
rect 13612 14512 13652 14552
rect 4928 14344 4968 14384
rect 5010 14344 5050 14384
rect 5092 14344 5132 14384
rect 5174 14344 5214 14384
rect 5256 14344 5296 14384
rect 20048 14344 20088 14384
rect 20130 14344 20170 14384
rect 20212 14344 20252 14384
rect 20294 14344 20334 14384
rect 20376 14344 20416 14384
rect 2668 14176 2708 14216
rect 12460 14176 12500 14216
rect 14284 14176 14324 14216
rect 18412 14176 18452 14216
rect 7660 14092 7700 14132
rect 9196 14092 9236 14132
rect 20140 14092 20180 14132
rect 2860 14003 2900 14043
rect 3340 14008 3380 14048
rect 3916 14008 3956 14048
rect 4300 14008 4340 14048
rect 4396 14008 4436 14048
rect 5932 14008 5972 14048
rect 6028 14008 6068 14048
rect 6412 14008 6452 14048
rect 6508 14008 6548 14048
rect 6988 14008 7028 14048
rect 7468 13994 7508 14034
rect 8428 14008 8468 14048
rect 8524 14008 8564 14048
rect 8716 14008 8756 14048
rect 9292 14008 9332 14048
rect 9580 14008 9620 14048
rect 11020 14008 11060 14048
rect 12268 14008 12308 14048
rect 12844 14008 12884 14048
rect 14092 14008 14132 14048
rect 14476 14008 14516 14048
rect 14764 14008 14804 14048
rect 14956 14008 14996 14048
rect 16204 14008 16244 14048
rect 16588 14008 16628 14048
rect 16684 14029 16724 14069
rect 16780 14008 16820 14048
rect 16876 14008 16916 14048
rect 17068 14008 17108 14048
rect 17260 14008 17300 14048
rect 17356 14008 17396 14048
rect 18220 14008 18260 14048
rect 18508 14008 18548 14048
rect 18700 14008 18740 14048
rect 19948 14008 19988 14048
rect 3820 13924 3860 13964
rect 8908 13840 8948 13880
rect 16396 13840 16436 13880
rect 17068 13840 17108 13880
rect 8716 13756 8756 13796
rect 14284 13756 14324 13796
rect 14476 13756 14516 13796
rect 3688 13588 3728 13628
rect 3770 13588 3810 13628
rect 3852 13588 3892 13628
rect 3934 13588 3974 13628
rect 4016 13588 4056 13628
rect 18808 13588 18848 13628
rect 18890 13588 18930 13628
rect 18972 13588 19012 13628
rect 19054 13588 19094 13628
rect 19136 13588 19176 13628
rect 7084 13420 7124 13460
rect 8716 13420 8756 13460
rect 14668 13420 14708 13460
rect 16972 13336 17012 13376
rect 11212 13252 11252 13292
rect 15628 13252 15668 13292
rect 2764 13173 2804 13213
rect 3244 13168 3284 13208
rect 3724 13168 3764 13208
rect 3820 13168 3860 13208
rect 4204 13168 4244 13208
rect 4300 13168 4340 13208
rect 5644 13168 5684 13208
rect 6892 13168 6932 13208
rect 7276 13168 7316 13208
rect 8524 13168 8564 13208
rect 8908 13168 8948 13208
rect 10156 13168 10196 13208
rect 10636 13168 10676 13208
rect 10732 13168 10772 13208
rect 11116 13168 11156 13208
rect 11692 13167 11732 13207
rect 12172 13177 12212 13217
rect 12652 13168 12692 13208
rect 12748 13168 12788 13208
rect 13132 13168 13172 13208
rect 13228 13168 13268 13208
rect 13708 13168 13748 13208
rect 14188 13182 14228 13222
rect 14764 13168 14804 13208
rect 15052 13168 15092 13208
rect 15148 13168 15188 13208
rect 15532 13168 15572 13208
rect 16108 13168 16148 13208
rect 16588 13173 16628 13213
rect 17356 13211 17396 13251
rect 17260 13168 17300 13208
rect 17836 13168 17876 13208
rect 19084 13168 19124 13208
rect 19564 13168 19604 13208
rect 19660 13168 19700 13208
rect 19756 13168 19796 13208
rect 2572 13084 2612 13124
rect 10348 13084 10388 13124
rect 12364 13084 12404 13124
rect 14380 13084 14420 13124
rect 8716 13000 8756 13040
rect 16780 13042 16820 13082
rect 19276 13000 19316 13040
rect 19468 13000 19508 13040
rect 17452 12942 17492 12982
rect 4928 12832 4968 12872
rect 5010 12832 5050 12872
rect 5092 12832 5132 12872
rect 5174 12832 5214 12872
rect 5256 12832 5296 12872
rect 20048 12832 20088 12872
rect 20130 12832 20170 12872
rect 20212 12832 20252 12872
rect 20294 12832 20334 12872
rect 20376 12832 20416 12872
rect 12268 12664 12308 12704
rect 19852 12664 19892 12704
rect 2284 12580 2324 12620
rect 7372 12580 7412 12620
rect 15244 12580 15284 12620
rect 15532 12580 15572 12620
rect 17644 12580 17684 12620
rect 2476 12496 2516 12536
rect 3724 12496 3764 12536
rect 3916 12496 3956 12536
rect 5164 12496 5204 12536
rect 5644 12496 5684 12536
rect 5740 12496 5780 12536
rect 6124 12496 6164 12536
rect 6220 12496 6260 12536
rect 6700 12496 6740 12536
rect 7180 12482 7220 12522
rect 7948 12496 7988 12536
rect 8044 12496 8084 12536
rect 8332 12496 8372 12536
rect 8812 12496 8852 12536
rect 10060 12496 10100 12536
rect 10828 12496 10868 12536
rect 12076 12496 12116 12536
rect 12940 12496 12980 12536
rect 13036 12496 13076 12536
rect 13132 12496 13172 12536
rect 13804 12496 13844 12536
rect 15052 12496 15092 12536
rect 15628 12496 15668 12536
rect 15820 12496 15860 12536
rect 15916 12496 15956 12536
rect 16108 12496 16148 12536
rect 16396 12496 16436 12536
rect 16684 12496 16724 12536
rect 16780 12496 16820 12536
rect 17260 12496 17300 12536
rect 17452 12496 17492 12536
rect 17740 12496 17780 12536
rect 17932 12496 17972 12536
rect 18028 12496 18068 12536
rect 18124 12496 18164 12536
rect 18220 12496 18260 12536
rect 18412 12496 18452 12536
rect 19660 12496 19700 12536
rect 17356 12412 17396 12452
rect 7660 12328 7700 12368
rect 17068 12328 17108 12368
rect 5356 12244 5396 12284
rect 8620 12244 8660 12284
rect 13324 12244 13364 12284
rect 16108 12244 16148 12284
rect 19852 12244 19892 12284
rect 3688 12076 3728 12116
rect 3770 12076 3810 12116
rect 3852 12076 3892 12116
rect 3934 12076 3974 12116
rect 4016 12076 4056 12116
rect 18808 12076 18848 12116
rect 18890 12076 18930 12116
rect 18972 12076 19012 12116
rect 19054 12076 19094 12116
rect 19136 12076 19176 12116
rect 2668 11908 2708 11948
rect 6892 11908 6932 11948
rect 8716 11908 8756 11948
rect 9196 11908 9236 11948
rect 16492 11908 16532 11948
rect 18508 11908 18548 11948
rect 18700 11824 18740 11864
rect 19084 11824 19124 11864
rect 20140 11824 20180 11864
rect 12364 11740 12404 11780
rect 12460 11740 12500 11780
rect 1228 11656 1268 11696
rect 2476 11656 2516 11696
rect 3628 11656 3668 11696
rect 3724 11656 3764 11696
rect 3820 11656 3860 11696
rect 5452 11656 5492 11696
rect 6700 11656 6740 11696
rect 7084 11656 7124 11696
rect 8332 11656 8372 11696
rect 8716 11656 8756 11696
rect 9004 11656 9044 11696
rect 9580 11656 9620 11696
rect 9868 11656 9908 11696
rect 10156 11656 10196 11696
rect 11404 11656 11444 11696
rect 11884 11656 11924 11696
rect 11980 11656 12020 11696
rect 12940 11656 12980 11696
rect 13420 11661 13460 11701
rect 13804 11656 13844 11696
rect 13996 11670 14036 11710
rect 14092 11656 14132 11696
rect 14284 11656 14324 11696
rect 14380 11656 14420 11696
rect 14476 11656 14516 11696
rect 15052 11656 15092 11696
rect 16300 11656 16340 11696
rect 16876 11656 16916 11696
rect 18124 11656 18164 11696
rect 18700 11656 18740 11696
rect 19372 11656 19412 11696
rect 19468 11656 19508 11696
rect 19756 11656 19796 11696
rect 20044 11656 20084 11696
rect 9484 11572 9524 11612
rect 18316 11572 18356 11612
rect 3532 11488 3572 11528
rect 8524 11488 8564 11528
rect 11596 11488 11636 11528
rect 13612 11488 13652 11528
rect 13900 11488 13940 11528
rect 14572 11488 14612 11528
rect 4928 11320 4968 11360
rect 5010 11320 5050 11360
rect 5092 11320 5132 11360
rect 5174 11320 5214 11360
rect 5256 11320 5296 11360
rect 20048 11320 20088 11360
rect 20130 11320 20170 11360
rect 20212 11320 20252 11360
rect 20294 11320 20334 11360
rect 20376 11320 20416 11360
rect 2668 11152 2708 11192
rect 4972 11152 5012 11192
rect 7276 11152 7316 11192
rect 7756 11152 7796 11192
rect 9772 11152 9812 11192
rect 11980 11152 12020 11192
rect 20044 11152 20084 11192
rect 3340 11068 3380 11108
rect 12748 11068 12788 11108
rect 1228 10984 1268 11024
rect 2476 10984 2516 11024
rect 3724 10984 3764 11024
rect 4396 10984 4436 11024
rect 3436 10942 3476 10982
rect 4492 10984 4532 11024
rect 4684 10984 4724 11024
rect 4876 10984 4916 11024
rect 5068 10984 5108 11024
rect 5164 10984 5204 11024
rect 5836 10984 5876 11024
rect 7084 10984 7124 11024
rect 7948 10979 7988 11019
rect 8428 10984 8468 11024
rect 8908 10984 8948 11024
rect 9388 10984 9428 11024
rect 9484 10984 9524 11024
rect 9868 10984 9908 11024
rect 9964 10984 10004 11024
rect 10060 10984 10100 11024
rect 10540 10984 10580 11024
rect 11788 10984 11828 11024
rect 12844 10984 12884 11024
rect 13132 10984 13172 11024
rect 13420 10984 13460 11024
rect 13708 10984 13748 11024
rect 17740 10984 17780 11024
rect 17836 10984 17876 11024
rect 18028 10984 18068 11024
rect 18316 10984 18356 11024
rect 18412 10984 18452 11024
rect 19372 10984 19412 11024
rect 19852 10979 19892 11019
rect 9004 10900 9044 10940
rect 13516 10900 13556 10940
rect 18796 10900 18836 10940
rect 18892 10900 18932 10940
rect 3052 10816 3092 10856
rect 12460 10816 12500 10856
rect 18028 10816 18068 10856
rect 3688 10564 3728 10604
rect 3770 10564 3810 10604
rect 3852 10564 3892 10604
rect 3934 10564 3974 10604
rect 4016 10564 4056 10604
rect 18808 10564 18848 10604
rect 18890 10564 18930 10604
rect 18972 10564 19012 10604
rect 19054 10564 19094 10604
rect 19136 10564 19176 10604
rect 2668 10396 2708 10436
rect 10636 10396 10676 10436
rect 12844 10396 12884 10436
rect 7948 10312 7988 10352
rect 19084 10312 19124 10352
rect 9196 10228 9236 10268
rect 9292 10228 9332 10268
rect 15436 10228 15476 10268
rect 1228 10144 1268 10184
rect 2476 10144 2516 10184
rect 3052 10158 3092 10198
rect 3532 10144 3572 10184
rect 4012 10144 4052 10184
rect 4108 10144 4148 10184
rect 4492 10144 4532 10184
rect 4588 10144 4628 10184
rect 7468 10144 7508 10184
rect 7564 10144 7604 10184
rect 7660 10144 7700 10184
rect 7756 10144 7796 10184
rect 8140 10144 8180 10184
rect 8236 10144 8276 10184
rect 8332 10144 8372 10184
rect 8716 10144 8756 10184
rect 8812 10144 8852 10184
rect 9772 10144 9812 10184
rect 10252 10149 10292 10189
rect 10636 10144 10676 10184
rect 10828 10144 10868 10184
rect 10924 10144 10964 10184
rect 11404 10144 11444 10184
rect 12652 10144 12692 10184
rect 13228 10144 13268 10184
rect 14476 10144 14516 10184
rect 14956 10144 14996 10184
rect 15052 10144 15092 10184
rect 15532 10144 15572 10184
rect 16012 10144 16052 10184
rect 16540 10153 16580 10193
rect 17452 10144 17492 10184
rect 18700 10144 18740 10184
rect 19468 10144 19508 10184
rect 19756 10144 19796 10184
rect 2860 10060 2900 10100
rect 10444 10060 10484 10100
rect 14668 10060 14708 10100
rect 16684 10060 16724 10100
rect 18892 10060 18932 10100
rect 19372 10060 19412 10100
rect 4928 9808 4968 9848
rect 5010 9808 5050 9848
rect 5092 9808 5132 9848
rect 5174 9808 5214 9848
rect 5256 9808 5296 9848
rect 20048 9808 20088 9848
rect 20130 9808 20170 9848
rect 20212 9808 20252 9848
rect 20294 9808 20334 9848
rect 20376 9808 20416 9848
rect 3724 9640 3764 9680
rect 5740 9640 5780 9680
rect 9676 9640 9716 9680
rect 10540 9640 10580 9680
rect 14668 9640 14708 9680
rect 16588 9640 16628 9680
rect 19756 9640 19796 9680
rect 2956 9556 2996 9596
rect 5548 9556 5588 9596
rect 9196 9556 9236 9596
rect 12652 9556 12692 9596
rect 1516 9472 1556 9512
rect 2764 9472 2804 9512
rect 3340 9472 3380 9512
rect 3436 9472 3476 9512
rect 3532 9472 3572 9512
rect 4108 9472 4148 9512
rect 5356 9472 5396 9512
rect 6412 9472 6452 9512
rect 6988 9472 7028 9512
rect 5884 9430 5924 9470
rect 7372 9472 7412 9512
rect 7468 9472 7508 9512
rect 7756 9472 7796 9512
rect 9004 9472 9044 9512
rect 9868 9472 9908 9512
rect 10060 9472 10100 9512
rect 9964 9430 10004 9470
rect 10348 9472 10388 9512
rect 10636 9472 10676 9512
rect 11212 9472 11252 9512
rect 12460 9472 12500 9512
rect 12940 9472 12980 9512
rect 13036 9472 13076 9512
rect 13516 9472 13556 9512
rect 13996 9472 14036 9512
rect 14476 9458 14516 9498
rect 14860 9472 14900 9512
rect 15148 9472 15188 9512
rect 16396 9472 16436 9512
rect 16972 9472 17012 9512
rect 17068 9472 17108 9512
rect 17164 9472 17204 9512
rect 17260 9472 17300 9512
rect 17644 9472 17684 9512
rect 18028 9472 18068 9512
rect 18124 9472 18164 9512
rect 19084 9472 19124 9512
rect 19564 9467 19604 9507
rect 19948 9472 19988 9512
rect 20140 9478 20180 9518
rect 20236 9472 20276 9512
rect 6892 9388 6932 9428
rect 13420 9388 13460 9428
rect 18508 9388 18548 9428
rect 18604 9388 18644 9428
rect 17452 9304 17492 9344
rect 17644 9304 17684 9344
rect 14956 9220 14996 9260
rect 19948 9220 19988 9260
rect 3688 9052 3728 9092
rect 3770 9052 3810 9092
rect 3852 9052 3892 9092
rect 3934 9052 3974 9092
rect 4016 9052 4056 9092
rect 18808 9052 18848 9092
rect 18890 9052 18930 9092
rect 18972 9052 19012 9092
rect 19054 9052 19094 9092
rect 19136 9052 19176 9092
rect 2668 8884 2708 8924
rect 5740 8884 5780 8924
rect 14476 8884 14516 8924
rect 3052 8800 3092 8840
rect 4492 8800 4532 8840
rect 9772 8800 9812 8840
rect 14956 8800 14996 8840
rect 19276 8800 19316 8840
rect 20140 8800 20180 8840
rect 10540 8716 10580 8756
rect 10636 8716 10676 8756
rect 19948 8716 19988 8756
rect 1228 8632 1268 8672
rect 2476 8632 2516 8672
rect 3436 8632 3476 8672
rect 3724 8632 3764 8672
rect 4012 8632 4052 8672
rect 4108 8632 4148 8672
rect 4300 8643 4340 8683
rect 4492 8632 4532 8672
rect 4780 8632 4820 8672
rect 5932 8632 5972 8672
rect 7180 8632 7220 8672
rect 8332 8632 8372 8672
rect 9580 8632 9620 8672
rect 10060 8632 10100 8672
rect 10156 8632 10196 8672
rect 11116 8632 11156 8672
rect 11596 8637 11636 8677
rect 13036 8632 13076 8672
rect 14284 8632 14324 8672
rect 14764 8632 14804 8672
rect 14956 8632 14996 8672
rect 15052 8632 15092 8672
rect 15244 8632 15284 8672
rect 15340 8632 15380 8672
rect 15532 8632 15572 8672
rect 15628 8632 15668 8672
rect 15729 8632 15769 8672
rect 16204 8632 16244 8672
rect 17452 8632 17492 8672
rect 17836 8632 17876 8672
rect 19084 8632 19124 8672
rect 19468 8632 19508 8672
rect 19564 8632 19604 8672
rect 19660 8632 19700 8672
rect 3340 8548 3380 8588
rect 11788 8548 11828 8588
rect 4204 8464 4244 8504
rect 15436 8464 15476 8504
rect 17644 8464 17684 8504
rect 19756 8464 19796 8504
rect 4928 8296 4968 8336
rect 5010 8296 5050 8336
rect 5092 8296 5132 8336
rect 5174 8296 5214 8336
rect 5256 8296 5296 8336
rect 20048 8296 20088 8336
rect 20130 8296 20170 8336
rect 20212 8296 20252 8336
rect 20294 8296 20334 8336
rect 20376 8296 20416 8336
rect 4396 8128 4436 8168
rect 9868 8128 9908 8168
rect 11500 8128 11540 8168
rect 15340 8128 15380 8168
rect 18604 8128 18644 8168
rect 8140 8044 8180 8084
rect 1996 7960 2036 8000
rect 2092 7960 2132 8000
rect 2188 7960 2228 8000
rect 2668 7960 2708 8000
rect 2764 7960 2804 8000
rect 3724 7960 3764 8000
rect 4204 7946 4244 7986
rect 4684 7960 4724 8000
rect 5932 7960 5972 8000
rect 6412 7960 6452 8000
rect 6508 7960 6548 8000
rect 6988 7960 7028 8000
rect 7468 7960 7508 8000
rect 7948 7946 7988 7986
rect 8428 7960 8468 8000
rect 9676 7960 9716 8000
rect 10060 7960 10100 8000
rect 11308 7960 11348 8000
rect 11692 7960 11732 8000
rect 12940 7960 12980 8000
rect 13900 7960 13940 8000
rect 15148 7960 15188 8000
rect 15532 7960 15572 8000
rect 16780 7960 16820 8000
rect 18028 7960 18068 8000
rect 18316 7960 18356 8000
rect 18508 7960 18548 8000
rect 19372 7960 19412 8000
rect 19468 7960 19508 8000
rect 19756 7960 19796 8000
rect 3148 7876 3188 7916
rect 3244 7876 3284 7916
rect 6892 7876 6932 7916
rect 6124 7792 6164 7832
rect 2380 7708 2420 7748
rect 13132 7708 13172 7748
rect 16972 7708 17012 7748
rect 18316 7708 18356 7748
rect 19084 7708 19124 7748
rect 3688 7540 3728 7580
rect 3770 7540 3810 7580
rect 3852 7540 3892 7580
rect 3934 7540 3974 7580
rect 4016 7540 4056 7580
rect 18808 7540 18848 7580
rect 18890 7540 18930 7580
rect 18972 7540 19012 7580
rect 19054 7540 19094 7580
rect 19136 7540 19176 7580
rect 2668 7372 2708 7412
rect 2860 7372 2900 7412
rect 7852 7372 7892 7412
rect 15724 7372 15764 7412
rect 19756 7372 19796 7412
rect 1228 7120 1268 7160
rect 2476 7120 2516 7160
rect 3052 7120 3092 7160
rect 4300 7120 4340 7160
rect 4492 7120 4532 7160
rect 4588 7120 4628 7160
rect 4684 7120 4724 7160
rect 6412 7120 6452 7160
rect 7660 7120 7700 7160
rect 8332 7120 8372 7160
rect 9580 7120 9620 7160
rect 9964 7120 10004 7160
rect 11212 7120 11252 7160
rect 11692 7120 11732 7160
rect 11788 7120 11828 7160
rect 12172 7120 12212 7160
rect 12268 7120 12308 7160
rect 12748 7120 12788 7160
rect 13228 7134 13268 7174
rect 14284 7120 14324 7160
rect 15532 7120 15572 7160
rect 15916 7120 15956 7160
rect 16012 7120 16052 7160
rect 16396 7120 16436 7160
rect 16684 7120 16724 7160
rect 17932 7120 17972 7160
rect 18316 7120 18356 7160
rect 19564 7120 19604 7160
rect 11404 7036 11444 7076
rect 18124 7036 18164 7076
rect 2668 6952 2708 6992
rect 4780 6952 4820 6992
rect 9772 6952 9812 6992
rect 13420 6952 13460 6992
rect 16204 6952 16244 6992
rect 16492 6952 16532 6992
rect 4928 6784 4968 6824
rect 5010 6784 5050 6824
rect 5092 6784 5132 6824
rect 5174 6784 5214 6824
rect 5256 6784 5296 6824
rect 20048 6784 20088 6824
rect 20130 6784 20170 6824
rect 20212 6784 20252 6824
rect 20294 6784 20334 6824
rect 20376 6784 20416 6824
rect 16684 6674 16724 6714
rect 2668 6616 2708 6656
rect 3244 6616 3284 6656
rect 6892 6616 6932 6656
rect 20044 6616 20084 6656
rect 10444 6532 10484 6572
rect 12652 6532 12692 6572
rect 14668 6532 14708 6572
rect 1228 6448 1268 6488
rect 2476 6448 2516 6488
rect 2956 6448 2996 6488
rect 3052 6448 3092 6488
rect 3148 6448 3188 6488
rect 3436 6448 3476 6488
rect 5164 6448 5204 6488
rect 4684 6406 4724 6446
rect 5260 6448 5300 6488
rect 5644 6448 5684 6488
rect 6220 6448 6260 6488
rect 6700 6434 6740 6474
rect 7084 6448 7124 6488
rect 8716 6448 8756 6488
rect 8812 6448 8852 6488
rect 9196 6448 9236 6488
rect 9292 6448 9332 6488
rect 9772 6448 9812 6488
rect 10252 6443 10292 6483
rect 11212 6448 11252 6488
rect 12460 6448 12500 6488
rect 12940 6448 12980 6488
rect 13036 6448 13076 6488
rect 13420 6448 13460 6488
rect 13996 6448 14036 6488
rect 5740 6364 5780 6404
rect 13516 6364 13556 6404
rect 14524 6406 14564 6446
rect 15724 6448 15764 6488
rect 15916 6448 15956 6488
rect 16012 6448 16052 6488
rect 16492 6448 16532 6488
rect 16588 6448 16628 6488
rect 16876 6448 16916 6488
rect 17068 6448 17108 6488
rect 17164 6448 17204 6488
rect 17644 6448 17684 6488
rect 17740 6448 17780 6488
rect 17836 6448 17876 6488
rect 18316 6448 18356 6488
rect 18412 6448 18452 6488
rect 18892 6448 18932 6488
rect 19372 6448 19412 6488
rect 19852 6443 19892 6483
rect 18796 6364 18836 6404
rect 4876 6280 4916 6320
rect 16876 6280 16916 6320
rect 18028 6280 18068 6320
rect 7180 6196 7220 6236
rect 15724 6196 15764 6236
rect 16204 6196 16244 6236
rect 3688 6028 3728 6068
rect 3770 6028 3810 6068
rect 3852 6028 3892 6068
rect 3934 6028 3974 6068
rect 4016 6028 4056 6068
rect 18808 6028 18848 6068
rect 18890 6028 18930 6068
rect 18972 6028 19012 6068
rect 19054 6028 19094 6068
rect 19136 6028 19176 6068
rect 1516 5860 1556 5900
rect 4972 5860 5012 5900
rect 6604 5860 6644 5900
rect 8428 5860 8468 5900
rect 14668 5860 14708 5900
rect 19756 5860 19796 5900
rect 15628 5776 15668 5816
rect 16012 5776 16052 5816
rect 16972 5776 17012 5816
rect 3628 5692 3668 5732
rect 3724 5692 3764 5732
rect 9196 5692 9236 5732
rect 9292 5692 9332 5732
rect 15532 5692 15572 5732
rect 15724 5692 15764 5732
rect 1804 5608 1844 5648
rect 1900 5608 1940 5648
rect 2188 5608 2228 5648
rect 2668 5613 2708 5653
rect 3148 5608 3188 5648
rect 4108 5608 4148 5648
rect 4204 5608 4244 5648
rect 4588 5608 4628 5648
rect 4684 5608 4724 5648
rect 4780 5608 4820 5648
rect 5164 5608 5204 5648
rect 6412 5608 6452 5648
rect 6988 5608 7028 5648
rect 8236 5608 8276 5648
rect 8716 5608 8756 5648
rect 8812 5608 8852 5648
rect 9772 5608 9812 5648
rect 10252 5622 10292 5662
rect 11404 5608 11444 5648
rect 12652 5608 12692 5648
rect 13228 5608 13268 5648
rect 14476 5608 14516 5648
rect 14956 5608 14996 5648
rect 15052 5608 15092 5648
rect 15148 5608 15188 5648
rect 15244 5608 15284 5648
rect 15436 5608 15476 5648
rect 15820 5608 15860 5648
rect 16396 5608 16436 5648
rect 16684 5608 16724 5648
rect 17356 5651 17396 5691
rect 17260 5608 17300 5648
rect 17644 5608 17684 5648
rect 17740 5616 17780 5656
rect 17836 5608 17876 5648
rect 17932 5653 17972 5693
rect 18316 5608 18356 5648
rect 19564 5608 19604 5648
rect 19948 5608 19988 5648
rect 20140 5650 20180 5690
rect 20044 5608 20084 5648
rect 20236 5608 20276 5648
rect 16300 5524 16340 5564
rect 2476 5440 2516 5480
rect 10444 5440 10484 5480
rect 12844 5440 12884 5480
rect 17452 5382 17492 5422
rect 4928 5272 4968 5312
rect 5010 5272 5050 5312
rect 5092 5272 5132 5312
rect 5174 5272 5214 5312
rect 5256 5272 5296 5312
rect 20048 5272 20088 5312
rect 20130 5272 20170 5312
rect 20212 5272 20252 5312
rect 20294 5272 20334 5312
rect 20376 5272 20416 5312
rect 8812 5020 8852 5060
rect 12844 5020 12884 5060
rect 14860 5020 14900 5060
rect 16492 5020 16532 5060
rect 1228 4936 1268 4976
rect 2476 4936 2516 4976
rect 2860 4936 2900 4976
rect 4108 4936 4148 4976
rect 4492 4936 4532 4976
rect 4780 4936 4820 4976
rect 5260 4936 5300 4976
rect 6508 4936 6548 4976
rect 7084 4936 7124 4976
rect 7180 4936 7220 4976
rect 8140 4936 8180 4976
rect 8620 4922 8660 4962
rect 9772 4936 9812 4976
rect 11020 4936 11060 4976
rect 11404 4936 11444 4976
rect 12652 4936 12692 4976
rect 13132 4956 13172 4996
rect 13228 4936 13268 4976
rect 13612 4936 13652 4976
rect 13708 4936 13748 4976
rect 14188 4936 14228 4976
rect 14668 4922 14708 4962
rect 15052 4936 15092 4976
rect 16300 4936 16340 4976
rect 16780 4936 16820 4976
rect 18412 4978 18452 5018
rect 17068 4936 17108 4976
rect 17740 4936 17780 4976
rect 18316 4936 18356 4976
rect 18604 4936 18644 4976
rect 7564 4852 7604 4892
rect 17164 4894 17204 4934
rect 19372 4936 19412 4976
rect 19468 4936 19508 4976
rect 19756 4936 19796 4976
rect 7660 4852 7700 4892
rect 2668 4768 2708 4808
rect 17452 4768 17492 4808
rect 19084 4768 19124 4808
rect 4300 4684 4340 4724
rect 4492 4684 4532 4724
rect 6700 4684 6740 4724
rect 11212 4684 11252 4724
rect 17644 4684 17684 4724
rect 18604 4684 18644 4724
rect 3688 4516 3728 4556
rect 3770 4516 3810 4556
rect 3852 4516 3892 4556
rect 3934 4516 3974 4556
rect 4016 4516 4056 4556
rect 18808 4516 18848 4556
rect 18890 4516 18930 4556
rect 18972 4516 19012 4556
rect 19054 4516 19094 4556
rect 19136 4516 19176 4556
rect 3148 4348 3188 4388
rect 8716 4348 8756 4388
rect 14764 4348 14804 4388
rect 16300 4348 16340 4388
rect 16588 4348 16628 4388
rect 4972 4264 5012 4304
rect 17644 4264 17684 4304
rect 5836 4180 5876 4220
rect 11884 4180 11924 4220
rect 18988 4180 19028 4220
rect 19084 4180 19124 4220
rect 1228 4096 1268 4136
rect 2476 4096 2516 4136
rect 2860 4096 2900 4136
rect 2956 4096 2996 4136
rect 3148 4096 3188 4136
rect 3340 4096 3380 4136
rect 4588 4096 4628 4136
rect 5356 4096 5396 4136
rect 5452 4096 5492 4136
rect 5932 4096 5972 4136
rect 6412 4096 6452 4136
rect 6892 4101 6932 4141
rect 7276 4096 7316 4136
rect 8524 4096 8564 4136
rect 9004 4096 9044 4136
rect 10252 4096 10292 4136
rect 11404 4096 11444 4136
rect 11500 4096 11540 4136
rect 11980 4096 12020 4136
rect 12459 4087 12499 4127
rect 12940 4110 12980 4150
rect 13324 4096 13364 4136
rect 14572 4096 14612 4136
rect 16396 4096 16436 4136
rect 16684 4096 16724 4136
rect 16972 4096 17012 4136
rect 17260 4096 17300 4136
rect 17356 4096 17396 4136
rect 18508 4096 18548 4136
rect 18604 4096 18644 4136
rect 19564 4096 19604 4136
rect 20044 4101 20084 4141
rect 4780 4012 4820 4052
rect 7084 4012 7124 4052
rect 20236 4012 20276 4052
rect 2668 3928 2708 3968
rect 10444 3928 10484 3968
rect 13132 3928 13172 3968
rect 4928 3760 4968 3800
rect 5010 3760 5050 3800
rect 5092 3760 5132 3800
rect 5174 3760 5214 3800
rect 5256 3760 5296 3800
rect 20048 3760 20088 3800
rect 20130 3760 20170 3800
rect 20212 3760 20252 3800
rect 20294 3760 20334 3800
rect 20376 3760 20416 3800
rect 17260 3650 17300 3690
rect 5068 3596 5108 3636
rect 6700 3592 6740 3632
rect 7084 3592 7124 3632
rect 2476 3508 2516 3548
rect 8236 3550 8276 3590
rect 15628 3592 15668 3632
rect 17452 3592 17492 3632
rect 19564 3592 19604 3632
rect 2668 3410 2708 3450
rect 3148 3424 3188 3464
rect 3628 3424 3668 3464
rect 4108 3424 4148 3464
rect 4204 3424 4244 3464
rect 4876 3424 4916 3464
rect 4972 3424 5012 3464
rect 5260 3424 5300 3464
rect 6508 3424 6548 3464
rect 6988 3424 7028 3464
rect 7180 3424 7220 3464
rect 7276 3405 7316 3445
rect 7468 3424 7508 3464
rect 7852 3424 7892 3464
rect 8044 3424 8084 3464
rect 8428 3424 8468 3464
rect 8620 3424 8660 3464
rect 16204 3466 16244 3506
rect 9004 3424 9044 3464
rect 9196 3424 9236 3464
rect 10444 3424 10484 3464
rect 11212 3424 11252 3464
rect 12460 3424 12500 3464
rect 14188 3424 14228 3464
rect 15436 3424 15476 3464
rect 16588 3424 16628 3464
rect 17068 3424 17108 3464
rect 17548 3424 17588 3464
rect 3724 3340 3764 3380
rect 7564 3340 7604 3380
rect 7756 3340 7796 3380
rect 8140 3340 8180 3380
rect 8332 3340 8372 3380
rect 8716 3340 8756 3380
rect 8908 3340 8948 3380
rect 16012 3340 16052 3380
rect 16300 3340 16340 3380
rect 17164 3382 17204 3422
rect 17644 3424 17684 3464
rect 17740 3424 17780 3464
rect 18124 3424 18164 3464
rect 19372 3424 19412 3464
rect 19756 3424 19796 3464
rect 20044 3424 20084 3464
rect 16492 3340 16532 3380
rect 19948 3340 19988 3380
rect 4588 3256 4628 3296
rect 7660 3256 7700 3296
rect 8812 3256 8852 3296
rect 16396 3256 16436 3296
rect 16780 3256 16820 3296
rect 10636 3172 10676 3212
rect 12652 3172 12692 3212
rect 15820 3172 15860 3212
rect 3688 3004 3728 3044
rect 3770 3004 3810 3044
rect 3852 3004 3892 3044
rect 3934 3004 3974 3044
rect 4016 3004 4056 3044
rect 18808 3004 18848 3044
rect 18890 3004 18930 3044
rect 18972 3004 19012 3044
rect 19054 3004 19094 3044
rect 19136 3004 19176 3044
rect 3436 2836 3476 2876
rect 5260 2836 5300 2876
rect 8716 2836 8756 2876
rect 9484 2836 9524 2876
rect 16204 2836 16244 2876
rect 18124 2836 18164 2876
rect 5836 2752 5876 2792
rect 7660 2752 7700 2792
rect 9292 2752 9332 2792
rect 10636 2752 10676 2792
rect 17644 2752 17684 2792
rect 18988 2752 19028 2792
rect 5452 2668 5492 2708
rect 11404 2668 11444 2708
rect 11500 2668 11540 2708
rect 13996 2668 14036 2708
rect 14188 2668 14228 2708
rect 1612 2584 1652 2624
rect 1804 2584 1844 2624
rect 1996 2584 2036 2624
rect 3244 2584 3284 2624
rect 3820 2584 3860 2624
rect 5068 2584 5108 2624
rect 6124 2584 6164 2624
rect 6220 2584 6260 2624
rect 6508 2584 6548 2624
rect 6796 2584 6836 2624
rect 6892 2584 6932 2624
rect 7084 2584 7124 2624
rect 7180 2584 7220 2624
rect 7281 2584 7321 2624
rect 7948 2584 7988 2624
rect 8044 2584 8084 2624
rect 8332 2584 8372 2624
rect 8716 2584 8756 2624
rect 9004 2584 9044 2624
rect 9484 2584 9524 2624
rect 9676 2584 9716 2624
rect 9964 2584 10004 2624
rect 10252 2584 10292 2624
rect 10348 2584 10388 2624
rect 10924 2584 10964 2624
rect 12508 2626 12548 2666
rect 11020 2584 11060 2624
rect 11980 2584 12020 2624
rect 14764 2584 14804 2624
rect 16012 2584 16052 2624
rect 16492 2584 16532 2624
rect 16588 2584 16628 2624
rect 16684 2584 16724 2624
rect 16972 2584 17012 2624
rect 17260 2584 17300 2624
rect 17356 2584 17396 2624
rect 17836 2584 17876 2624
rect 17932 2584 17972 2624
rect 18124 2584 18164 2624
rect 18508 2584 18548 2624
rect 18604 2584 18644 2624
rect 18700 2584 18740 2624
rect 18796 2584 18836 2624
rect 19180 2584 19220 2624
rect 19276 2584 19316 2624
rect 19372 2584 19412 2624
rect 19660 2584 19700 2624
rect 19756 2584 19796 2624
rect 19948 2584 19988 2624
rect 1708 2500 1748 2540
rect 12652 2500 12692 2540
rect 19852 2500 19892 2540
rect 5644 2416 5684 2456
rect 6988 2416 7028 2456
rect 9196 2416 9236 2456
rect 13804 2416 13844 2456
rect 14380 2416 14420 2456
rect 16396 2416 16436 2456
rect 4928 2248 4968 2288
rect 5010 2248 5050 2288
rect 5092 2248 5132 2288
rect 5174 2248 5214 2288
rect 5256 2248 5296 2288
rect 20048 2248 20088 2288
rect 20130 2248 20170 2288
rect 20212 2248 20252 2288
rect 20294 2248 20334 2288
rect 20376 2248 20416 2288
rect 2764 2080 2804 2120
rect 8332 2080 8372 2120
rect 8620 2080 8660 2120
rect 8908 2080 8948 2120
rect 9868 2080 9908 2120
rect 14956 2080 14996 2120
rect 17356 2084 17396 2124
rect 19852 2080 19892 2120
rect 12940 1996 12980 2036
rect 1324 1912 1364 1952
rect 2572 1912 2612 1952
rect 3532 1912 3572 1952
rect 4780 1912 4820 1952
rect 4972 1912 5012 1952
rect 6220 1912 6260 1952
rect 6988 1912 7028 1952
rect 7180 1912 7220 1952
rect 7276 1912 7316 1952
rect 7660 1912 7700 1952
rect 7756 1912 7796 1952
rect 7852 1912 7892 1952
rect 7948 1912 7988 1952
rect 8140 1912 8180 1952
rect 8236 1912 8276 1952
rect 8428 1901 8468 1941
rect 8716 1912 8756 1952
rect 9772 1912 9812 1952
rect 10060 1912 10100 1952
rect 11500 1912 11540 1952
rect 12748 1912 12788 1952
rect 13228 1912 13268 1952
rect 13324 1912 13364 1952
rect 13708 1912 13748 1952
rect 14284 1912 14324 1952
rect 14764 1898 14804 1938
rect 15244 1912 15284 1952
rect 16492 1912 16532 1952
rect 17164 1912 17204 1952
rect 17260 1912 17300 1952
rect 17548 1912 17588 1952
rect 17644 1912 17684 1952
rect 17836 1912 17876 1952
rect 18028 1912 18068 1952
rect 18124 1912 18164 1952
rect 18412 1912 18452 1952
rect 19660 1912 19700 1952
rect 2956 1828 2996 1868
rect 6604 1828 6644 1868
rect 9196 1828 9236 1868
rect 10348 1828 10388 1868
rect 10732 1828 10772 1868
rect 11116 1828 11156 1868
rect 13804 1828 13844 1868
rect 6988 1744 7028 1784
rect 16876 1744 16916 1784
rect 17836 1744 17876 1784
rect 3148 1660 3188 1700
rect 3340 1660 3380 1700
rect 6412 1660 6452 1700
rect 6796 1660 6836 1700
rect 9388 1660 9428 1700
rect 10540 1660 10580 1700
rect 10924 1660 10964 1700
rect 11308 1660 11348 1700
rect 16684 1660 16724 1700
rect 3688 1492 3728 1532
rect 3770 1492 3810 1532
rect 3852 1492 3892 1532
rect 3934 1492 3974 1532
rect 4016 1492 4056 1532
rect 18808 1492 18848 1532
rect 18890 1492 18930 1532
rect 18972 1492 19012 1532
rect 19054 1492 19094 1532
rect 19136 1492 19176 1532
rect 6028 1324 6068 1364
rect 14668 1324 14708 1364
rect 17356 1324 17396 1364
rect 17740 1324 17780 1364
rect 6220 1240 6260 1280
rect 9196 1240 9236 1280
rect 17164 1240 17204 1280
rect 19564 1240 19604 1280
rect 2380 1156 2420 1196
rect 4396 1156 4436 1196
rect 7660 1156 7700 1196
rect 8044 1156 8084 1196
rect 8428 1156 8468 1196
rect 8812 1156 8852 1196
rect 9580 1156 9620 1196
rect 9964 1156 10004 1196
rect 10348 1156 10388 1196
rect 10924 1156 10964 1196
rect 11212 1156 11252 1196
rect 11788 1156 11828 1196
rect 14860 1156 14900 1196
rect 15532 1156 15572 1196
rect 2764 1072 2804 1112
rect 4012 1072 4052 1112
rect 4780 1072 4820 1112
rect 4876 1072 4916 1112
rect 4972 1072 5012 1112
rect 5068 1072 5108 1112
rect 5356 1072 5396 1112
rect 5644 1072 5684 1112
rect 6316 1072 6356 1112
rect 6508 1072 6548 1112
rect 6604 1072 6644 1112
rect 7372 1072 7412 1112
rect 7473 1063 7513 1103
rect 13228 1072 13268 1112
rect 14476 1072 14516 1112
rect 15724 1072 15764 1112
rect 16972 1072 17012 1112
rect 17452 1072 17492 1112
rect 17644 1072 17684 1112
rect 18124 1072 18164 1112
rect 19372 1072 19412 1112
rect 4204 988 4244 1028
rect 5740 988 5780 1028
rect 2572 904 2612 944
rect 4588 904 4628 944
rect 6796 904 6836 944
rect 7180 904 7220 944
rect 7852 904 7892 944
rect 8236 904 8276 944
rect 8620 904 8660 944
rect 9004 904 9044 944
rect 9772 904 9812 944
rect 10156 904 10196 944
rect 10540 904 10580 944
rect 10732 904 10772 944
rect 11404 904 11444 944
rect 11596 904 11636 944
rect 15052 904 15092 944
rect 15340 904 15380 944
rect 4928 736 4968 776
rect 5010 736 5050 776
rect 5092 736 5132 776
rect 5174 736 5214 776
rect 5256 736 5296 776
rect 20048 736 20088 776
rect 20130 736 20170 776
rect 20212 736 20252 776
rect 20294 736 20334 776
rect 20376 736 20416 776
<< metal2 >>
rect 1784 42928 1864 43008
rect 1976 42928 2056 43008
rect 2168 42928 2248 43008
rect 2360 42928 2440 43008
rect 2552 42928 2632 43008
rect 2744 42928 2824 43008
rect 2936 42928 3016 43008
rect 3128 42928 3208 43008
rect 3320 42928 3400 43008
rect 3512 42928 3592 43008
rect 3704 42928 3784 43008
rect 3896 42928 3976 43008
rect 4088 42928 4168 43008
rect 4280 42928 4360 43008
rect 4472 42928 4552 43008
rect 4664 42928 4744 43008
rect 4856 42928 4936 43008
rect 5048 42928 5128 43008
rect 5240 42928 5320 43008
rect 5432 42928 5512 43008
rect 5624 42928 5704 43008
rect 5816 42928 5896 43008
rect 6008 42928 6088 43008
rect 6200 42928 6280 43008
rect 6392 42928 6472 43008
rect 6584 42928 6664 43008
rect 6776 42928 6856 43008
rect 6968 42928 7048 43008
rect 7160 42928 7240 43008
rect 7352 42928 7432 43008
rect 7544 42928 7624 43008
rect 7736 42928 7816 43008
rect 7928 42928 8008 43008
rect 8120 42928 8200 43008
rect 8312 42928 8392 43008
rect 8504 42928 8584 43008
rect 8696 42928 8776 43008
rect 8888 42928 8968 43008
rect 9080 42928 9160 43008
rect 9272 42928 9352 43008
rect 9464 42928 9544 43008
rect 9656 42928 9736 43008
rect 9848 42928 9928 43008
rect 10040 42928 10120 43008
rect 10232 42928 10312 43008
rect 10424 42928 10504 43008
rect 10616 42928 10696 43008
rect 10808 42928 10888 43008
rect 11000 42928 11080 43008
rect 11192 42928 11272 43008
rect 11384 42928 11464 43008
rect 11576 42928 11656 43008
rect 11768 42928 11848 43008
rect 11960 42928 12040 43008
rect 12152 42928 12232 43008
rect 12344 42928 12424 43008
rect 12536 42928 12616 43008
rect 12728 42928 12808 43008
rect 12920 42928 13000 43008
rect 13112 42928 13192 43008
rect 13304 42928 13384 43008
rect 13496 42928 13576 43008
rect 13688 42928 13768 43008
rect 13880 42928 13960 43008
rect 14072 42928 14152 43008
rect 14264 42928 14344 43008
rect 14456 42928 14536 43008
rect 14648 42928 14728 43008
rect 14840 42928 14920 43008
rect 15032 42928 15112 43008
rect 15224 42928 15304 43008
rect 15416 42928 15496 43008
rect 15608 42928 15688 43008
rect 15800 42928 15880 43008
rect 15992 42928 16072 43008
rect 16184 42928 16264 43008
rect 16376 42928 16456 43008
rect 16568 42928 16648 43008
rect 16760 42928 16840 43008
rect 16952 42928 17032 43008
rect 17144 42928 17224 43008
rect 17336 42928 17416 43008
rect 17528 42928 17608 43008
rect 17720 42928 17800 43008
rect 17912 42928 17992 43008
rect 18104 42928 18184 43008
rect 18296 42928 18376 43008
rect 18488 42928 18568 43008
rect 18680 42928 18760 43008
rect 18872 42928 18952 43008
rect 19064 42928 19144 43008
rect 19256 42928 19336 43008
rect 19448 42928 19528 43008
rect 1804 42860 1844 42928
rect 1612 42820 1844 42860
rect 1324 41096 1364 41105
rect 1324 40601 1364 41056
rect 1419 41012 1461 41021
rect 1419 40972 1420 41012
rect 1460 40972 1461 41012
rect 1419 40963 1461 40972
rect 1323 40592 1365 40601
rect 1323 40552 1324 40592
rect 1364 40552 1365 40592
rect 1323 40543 1365 40552
rect 1324 40458 1364 40543
rect 1420 39920 1460 40963
rect 1515 40592 1557 40601
rect 1515 40552 1516 40592
rect 1556 40552 1557 40592
rect 1515 40543 1557 40552
rect 1516 40508 1556 40543
rect 1516 40457 1556 40468
rect 1420 39871 1460 39880
rect 1228 39668 1268 39677
rect 940 39628 1228 39668
rect 843 38156 885 38165
rect 843 38116 844 38156
rect 884 38116 885 38156
rect 843 38107 885 38116
rect 844 28253 884 38107
rect 843 28244 885 28253
rect 843 28204 844 28244
rect 884 28204 885 28244
rect 843 28195 885 28204
rect 75 26732 117 26741
rect 75 26692 76 26732
rect 116 26692 117 26732
rect 75 26683 117 26692
rect 76 26489 116 26683
rect 75 26480 117 26489
rect 75 26440 76 26480
rect 116 26440 117 26480
rect 75 26431 117 26440
rect 171 25808 213 25817
rect 171 25768 172 25808
rect 212 25768 213 25808
rect 171 25759 213 25768
rect 75 17912 117 17921
rect 75 17872 76 17912
rect 116 17872 117 17912
rect 75 17863 117 17872
rect 76 6077 116 17863
rect 172 13889 212 25759
rect 555 19424 597 19433
rect 555 19384 556 19424
rect 596 19384 597 19424
rect 555 19375 597 19384
rect 267 18500 309 18509
rect 267 18460 268 18500
rect 308 18460 309 18500
rect 267 18451 309 18460
rect 171 13880 213 13889
rect 171 13840 172 13880
rect 212 13840 213 13880
rect 171 13831 213 13840
rect 75 6068 117 6077
rect 75 6028 76 6068
rect 116 6028 117 6068
rect 75 6019 117 6028
rect 268 3305 308 18451
rect 459 17660 501 17669
rect 459 17620 460 17660
rect 500 17620 501 17660
rect 459 17611 501 17620
rect 363 14048 405 14057
rect 363 14008 364 14048
rect 404 14008 405 14048
rect 363 13999 405 14008
rect 364 4313 404 13999
rect 363 4304 405 4313
rect 363 4264 364 4304
rect 404 4264 405 4304
rect 363 4255 405 4264
rect 267 3296 309 3305
rect 267 3256 268 3296
rect 308 3256 309 3296
rect 267 3247 309 3256
rect 460 2801 500 17611
rect 556 11285 596 19375
rect 651 18332 693 18341
rect 651 18292 652 18332
rect 692 18292 693 18332
rect 651 18283 693 18292
rect 555 11276 597 11285
rect 555 11236 556 11276
rect 596 11236 597 11276
rect 555 11227 597 11236
rect 652 7337 692 18283
rect 940 13133 980 39628
rect 1228 39619 1268 39628
rect 1419 39584 1461 39593
rect 1419 39544 1420 39584
rect 1460 39544 1461 39584
rect 1419 39535 1461 39544
rect 1323 38996 1365 39005
rect 1323 38956 1324 38996
rect 1364 38956 1365 38996
rect 1323 38947 1365 38956
rect 1324 38862 1364 38947
rect 1420 38576 1460 39535
rect 1516 39080 1556 39089
rect 1516 38921 1556 39040
rect 1515 38912 1557 38921
rect 1515 38872 1516 38912
rect 1556 38872 1557 38912
rect 1515 38863 1557 38872
rect 1324 38536 1460 38576
rect 1035 38492 1077 38501
rect 1035 38452 1036 38492
rect 1076 38452 1077 38492
rect 1035 38443 1077 38452
rect 1036 21113 1076 38443
rect 1227 38156 1269 38165
rect 1227 38116 1228 38156
rect 1268 38116 1269 38156
rect 1227 38107 1269 38116
rect 1228 38022 1268 38107
rect 1228 37484 1268 37493
rect 1132 37444 1228 37484
rect 1035 21104 1077 21113
rect 1035 21064 1036 21104
rect 1076 21064 1077 21104
rect 1035 21055 1077 21064
rect 1132 16409 1172 37444
rect 1228 37435 1268 37444
rect 1324 36821 1364 38536
rect 1419 38408 1461 38417
rect 1419 38368 1420 38408
rect 1460 38368 1461 38408
rect 1419 38359 1461 38368
rect 1420 38274 1460 38359
rect 1612 38324 1652 42820
rect 1707 42524 1749 42533
rect 1707 42484 1708 42524
rect 1748 42484 1749 42524
rect 1707 42475 1749 42484
rect 1708 40676 1748 42475
rect 1996 41600 2036 42928
rect 1900 41560 2036 41600
rect 1803 41264 1845 41273
rect 1803 41224 1804 41264
rect 1844 41224 1845 41264
rect 1803 41215 1845 41224
rect 1804 41130 1844 41215
rect 1708 40627 1748 40636
rect 1707 39752 1749 39761
rect 1707 39712 1708 39752
rect 1748 39712 1749 39752
rect 1707 39703 1749 39712
rect 1708 39618 1748 39703
rect 1707 38912 1749 38921
rect 1707 38872 1708 38912
rect 1748 38872 1749 38912
rect 1707 38863 1749 38872
rect 1708 38778 1748 38863
rect 1803 38744 1845 38753
rect 1803 38704 1804 38744
rect 1844 38704 1845 38744
rect 1803 38695 1845 38704
rect 1804 38408 1844 38695
rect 1804 38359 1844 38368
rect 1612 38284 1748 38324
rect 1612 38156 1652 38165
rect 1612 37913 1652 38116
rect 1611 37904 1653 37913
rect 1611 37864 1612 37904
rect 1652 37864 1653 37904
rect 1611 37855 1653 37864
rect 1515 37736 1557 37745
rect 1515 37696 1516 37736
rect 1556 37696 1557 37736
rect 1515 37687 1557 37696
rect 1419 37568 1461 37577
rect 1419 37528 1420 37568
rect 1460 37528 1461 37568
rect 1419 37519 1461 37528
rect 1420 37434 1460 37519
rect 1516 37316 1556 37687
rect 1611 37484 1653 37493
rect 1611 37444 1612 37484
rect 1652 37444 1653 37484
rect 1611 37435 1653 37444
rect 1612 37350 1652 37435
rect 1420 37276 1556 37316
rect 1323 36812 1365 36821
rect 1228 36772 1324 36812
rect 1364 36772 1365 36812
rect 1228 35720 1268 36772
rect 1323 36763 1365 36772
rect 1323 36644 1365 36653
rect 1323 36604 1324 36644
rect 1364 36604 1365 36644
rect 1323 36595 1365 36604
rect 1324 36510 1364 36595
rect 1323 35972 1365 35981
rect 1323 35932 1324 35972
rect 1364 35932 1365 35972
rect 1420 35972 1460 37276
rect 1611 37064 1653 37073
rect 1611 37024 1612 37064
rect 1652 37024 1653 37064
rect 1611 37015 1653 37024
rect 1515 36980 1557 36989
rect 1515 36940 1516 36980
rect 1556 36940 1557 36980
rect 1515 36931 1557 36940
rect 1516 36896 1556 36931
rect 1516 36845 1556 36856
rect 1516 36140 1556 36149
rect 1612 36140 1652 37015
rect 1708 36812 1748 38284
rect 1803 37652 1845 37661
rect 1803 37612 1804 37652
rect 1844 37612 1845 37652
rect 1803 37603 1845 37612
rect 1804 37518 1844 37603
rect 1900 37073 1940 41560
rect 2091 40676 2133 40685
rect 2091 40636 2092 40676
rect 2132 40636 2133 40676
rect 2091 40627 2133 40636
rect 2092 40424 2132 40627
rect 1996 40384 2092 40424
rect 1996 38669 2036 40384
rect 2092 40375 2132 40384
rect 2091 40004 2133 40013
rect 2091 39964 2092 40004
rect 2132 39964 2133 40004
rect 2091 39955 2133 39964
rect 1995 38660 2037 38669
rect 1995 38620 1996 38660
rect 2036 38620 2037 38660
rect 1995 38611 2037 38620
rect 2092 38333 2132 39955
rect 2091 38324 2133 38333
rect 2091 38284 2092 38324
rect 2132 38284 2133 38324
rect 2091 38275 2133 38284
rect 1996 38156 2036 38165
rect 2188 38156 2228 42928
rect 2283 40928 2325 40937
rect 2283 40888 2284 40928
rect 2324 40888 2325 40928
rect 2283 40879 2325 40888
rect 1996 37241 2036 38116
rect 2092 38116 2228 38156
rect 1995 37232 2037 37241
rect 1995 37192 1996 37232
rect 2036 37192 2037 37232
rect 1995 37183 2037 37192
rect 1996 37098 2036 37183
rect 1899 37064 1941 37073
rect 1899 37024 1900 37064
rect 1940 37024 1941 37064
rect 1899 37015 1941 37024
rect 1899 36896 1941 36905
rect 1899 36856 1900 36896
rect 1940 36856 1941 36896
rect 1899 36847 1941 36856
rect 1708 36772 1844 36812
rect 1708 36644 1748 36653
rect 1708 36485 1748 36604
rect 1707 36476 1749 36485
rect 1707 36436 1708 36476
rect 1748 36436 1749 36476
rect 1707 36427 1749 36436
rect 1556 36100 1652 36140
rect 1516 36091 1556 36100
rect 1707 36056 1749 36065
rect 1707 36016 1708 36056
rect 1748 36016 1749 36056
rect 1707 36007 1749 36016
rect 1420 35932 1556 35972
rect 1323 35923 1365 35932
rect 1324 35838 1364 35923
rect 1228 35680 1364 35720
rect 1227 34376 1269 34385
rect 1227 34336 1228 34376
rect 1268 34336 1269 34376
rect 1227 34327 1269 34336
rect 1228 34242 1268 34327
rect 1324 33368 1364 35680
rect 1419 35132 1461 35141
rect 1419 35092 1420 35132
rect 1460 35092 1461 35132
rect 1419 35083 1461 35092
rect 1420 34998 1460 35083
rect 1516 34973 1556 35932
rect 1611 35048 1653 35057
rect 1611 35008 1612 35048
rect 1652 35008 1653 35048
rect 1611 34999 1653 35008
rect 1515 34964 1557 34973
rect 1515 34924 1516 34964
rect 1556 34924 1557 34964
rect 1515 34915 1557 34924
rect 1516 33704 1556 34915
rect 1612 34914 1652 34999
rect 1611 33956 1653 33965
rect 1611 33916 1612 33956
rect 1652 33916 1653 33956
rect 1611 33907 1653 33916
rect 1612 33872 1652 33907
rect 1612 33821 1652 33832
rect 1516 33664 1652 33704
rect 1419 33620 1461 33629
rect 1419 33580 1420 33620
rect 1460 33580 1461 33620
rect 1419 33571 1461 33580
rect 1420 33486 1460 33571
rect 1324 33328 1460 33368
rect 1323 32948 1365 32957
rect 1323 32908 1324 32948
rect 1364 32908 1365 32948
rect 1323 32899 1365 32908
rect 1324 32814 1364 32899
rect 1228 31352 1268 31361
rect 1323 31352 1365 31361
rect 1268 31312 1324 31352
rect 1364 31312 1365 31352
rect 1228 31303 1268 31312
rect 1323 31303 1365 31312
rect 1228 29840 1268 29849
rect 1323 29840 1365 29849
rect 1268 29800 1324 29840
rect 1364 29800 1365 29840
rect 1228 29791 1268 29800
rect 1323 29791 1365 29800
rect 1227 26816 1269 26825
rect 1227 26776 1228 26816
rect 1268 26776 1269 26816
rect 1227 26767 1269 26776
rect 1228 26682 1268 26767
rect 1227 24632 1269 24641
rect 1227 24592 1228 24632
rect 1268 24592 1269 24632
rect 1227 24583 1269 24592
rect 1228 24498 1268 24583
rect 1227 23792 1269 23801
rect 1227 23752 1228 23792
rect 1268 23752 1269 23792
rect 1227 23743 1269 23752
rect 1228 22196 1268 23743
rect 1324 22280 1364 29791
rect 1420 29000 1460 33328
rect 1515 33200 1557 33209
rect 1515 33160 1516 33200
rect 1556 33160 1557 33200
rect 1515 33151 1557 33160
rect 1516 33116 1556 33151
rect 1516 33065 1556 33076
rect 1515 32864 1557 32873
rect 1515 32824 1516 32864
rect 1556 32824 1557 32864
rect 1515 32815 1557 32824
rect 1516 29849 1556 32815
rect 1612 32789 1652 33664
rect 1708 33116 1748 36007
rect 1804 33965 1844 36772
rect 1900 36762 1940 36847
rect 1899 35384 1941 35393
rect 1899 35344 1900 35384
rect 1940 35344 1941 35384
rect 1899 35335 1941 35344
rect 1900 35216 1940 35335
rect 1900 35167 1940 35176
rect 1995 35216 2037 35225
rect 1995 35176 1996 35216
rect 2036 35176 2037 35216
rect 1995 35167 2037 35176
rect 1803 33956 1845 33965
rect 1803 33916 1804 33956
rect 1844 33916 1845 33956
rect 1803 33907 1845 33916
rect 1899 33872 1941 33881
rect 1899 33832 1900 33872
rect 1940 33832 1941 33872
rect 1899 33823 1941 33832
rect 1900 33704 1940 33823
rect 1900 33655 1940 33664
rect 1996 33704 2036 35167
rect 2092 35057 2132 38116
rect 2187 37988 2229 37997
rect 2187 37948 2188 37988
rect 2228 37948 2229 37988
rect 2187 37939 2229 37948
rect 2188 37854 2228 37939
rect 2284 37661 2324 40879
rect 2283 37652 2325 37661
rect 2283 37612 2284 37652
rect 2324 37612 2325 37652
rect 2283 37603 2325 37612
rect 2283 37064 2325 37073
rect 2283 37024 2284 37064
rect 2324 37024 2325 37064
rect 2283 37015 2325 37024
rect 2188 36644 2228 36653
rect 2188 35729 2228 36604
rect 2187 35720 2229 35729
rect 2187 35680 2188 35720
rect 2228 35680 2229 35720
rect 2187 35671 2229 35680
rect 2188 35586 2228 35671
rect 2091 35048 2133 35057
rect 2091 35008 2092 35048
rect 2132 35008 2133 35048
rect 2091 34999 2133 35008
rect 2091 34544 2133 34553
rect 2091 34504 2092 34544
rect 2132 34504 2133 34544
rect 2091 34495 2133 34504
rect 1899 33200 1941 33209
rect 1899 33160 1900 33200
rect 1940 33160 1941 33200
rect 1899 33151 1941 33160
rect 1900 33116 1940 33151
rect 1708 33076 1844 33116
rect 1707 32948 1749 32957
rect 1707 32908 1708 32948
rect 1748 32908 1749 32948
rect 1707 32899 1749 32908
rect 1708 32814 1748 32899
rect 1611 32780 1653 32789
rect 1611 32740 1612 32780
rect 1652 32740 1653 32780
rect 1611 32731 1653 32740
rect 1804 32528 1844 33076
rect 1900 33065 1940 33076
rect 1899 32780 1941 32789
rect 1899 32740 1900 32780
rect 1940 32740 1941 32780
rect 1899 32731 1941 32740
rect 1708 32488 1844 32528
rect 1515 29840 1557 29849
rect 1515 29800 1516 29840
rect 1556 29800 1557 29840
rect 1515 29791 1557 29800
rect 1516 29168 1556 29177
rect 1708 29168 1748 32488
rect 1803 31100 1845 31109
rect 1803 31060 1804 31100
rect 1844 31060 1845 31100
rect 1803 31051 1845 31060
rect 1804 29345 1844 31051
rect 1803 29336 1845 29345
rect 1803 29296 1804 29336
rect 1844 29296 1845 29336
rect 1803 29287 1845 29296
rect 1556 29128 1748 29168
rect 1516 29119 1556 29128
rect 1420 28960 1652 29000
rect 1612 26144 1652 28960
rect 1708 27245 1748 29128
rect 1707 27236 1749 27245
rect 1707 27196 1708 27236
rect 1748 27196 1749 27236
rect 1707 27187 1749 27196
rect 1707 27068 1749 27077
rect 1707 27028 1708 27068
rect 1748 27028 1749 27068
rect 1707 27019 1749 27028
rect 1515 25976 1557 25985
rect 1515 25936 1516 25976
rect 1556 25936 1557 25976
rect 1515 25927 1557 25936
rect 1419 25472 1461 25481
rect 1419 25432 1420 25472
rect 1460 25432 1461 25472
rect 1419 25423 1461 25432
rect 1420 23885 1460 25423
rect 1516 24641 1556 25927
rect 1612 25061 1652 26104
rect 1708 25304 1748 27019
rect 1804 26825 1844 29287
rect 1900 28925 1940 32731
rect 1996 30596 2036 33664
rect 2092 31109 2132 34495
rect 2284 33200 2324 37015
rect 2380 36989 2420 42928
rect 2572 42869 2612 42928
rect 2571 42860 2613 42869
rect 2571 42820 2572 42860
rect 2612 42820 2613 42860
rect 2571 42811 2613 42820
rect 2764 41768 2804 42928
rect 2764 41728 2900 41768
rect 2763 40760 2805 40769
rect 2763 40720 2764 40760
rect 2804 40720 2805 40760
rect 2763 40711 2805 40720
rect 2667 40424 2709 40433
rect 2667 40384 2668 40424
rect 2708 40384 2709 40424
rect 2667 40375 2709 40384
rect 2475 38660 2517 38669
rect 2475 38620 2476 38660
rect 2516 38620 2517 38660
rect 2475 38611 2517 38620
rect 2476 38240 2516 38611
rect 2476 38191 2516 38200
rect 2572 38240 2612 38249
rect 2475 38072 2517 38081
rect 2475 38032 2476 38072
rect 2516 38032 2517 38072
rect 2475 38023 2517 38032
rect 2476 37400 2516 38023
rect 2572 37409 2612 38200
rect 2668 37661 2708 40375
rect 2667 37652 2709 37661
rect 2667 37612 2668 37652
rect 2708 37612 2709 37652
rect 2667 37603 2709 37612
rect 2476 37351 2516 37360
rect 2571 37400 2613 37409
rect 2571 37360 2572 37400
rect 2612 37360 2613 37400
rect 2571 37351 2613 37360
rect 2572 37266 2612 37351
rect 2667 37316 2709 37325
rect 2667 37276 2668 37316
rect 2708 37276 2709 37316
rect 2667 37267 2709 37276
rect 2379 36980 2421 36989
rect 2379 36940 2380 36980
rect 2420 36940 2421 36980
rect 2379 36931 2421 36940
rect 2379 36728 2421 36737
rect 2379 36688 2380 36728
rect 2420 36688 2421 36728
rect 2379 36679 2421 36688
rect 2380 36560 2420 36679
rect 2380 36511 2420 36520
rect 2668 35468 2708 37267
rect 2764 36821 2804 40711
rect 2763 36812 2805 36821
rect 2763 36772 2764 36812
rect 2804 36772 2805 36812
rect 2763 36763 2805 36772
rect 2763 35972 2805 35981
rect 2763 35932 2764 35972
rect 2804 35932 2805 35972
rect 2763 35923 2805 35932
rect 2380 35428 2708 35468
rect 2380 35132 2420 35428
rect 2469 35309 2509 35333
rect 2468 35300 2510 35309
rect 2468 35260 2469 35300
rect 2509 35260 2516 35300
rect 2468 35251 2516 35260
rect 2476 35216 2516 35251
rect 2516 35176 2612 35216
rect 2476 35148 2516 35176
rect 2380 33620 2420 35092
rect 2476 34376 2516 34385
rect 2476 33965 2516 34336
rect 2475 33956 2517 33965
rect 2475 33916 2476 33956
rect 2516 33916 2517 33956
rect 2475 33907 2517 33916
rect 2476 33704 2516 33713
rect 2572 33704 2612 35176
rect 2516 33664 2612 33704
rect 2476 33655 2516 33664
rect 2380 33209 2420 33580
rect 2475 33452 2517 33461
rect 2475 33412 2476 33452
rect 2516 33412 2517 33452
rect 2475 33403 2517 33412
rect 2188 33160 2324 33200
rect 2379 33200 2421 33209
rect 2379 33160 2380 33200
rect 2420 33160 2421 33200
rect 2188 31361 2228 33160
rect 2379 33151 2421 33160
rect 2283 33032 2325 33041
rect 2283 32992 2284 33032
rect 2324 32992 2325 33032
rect 2283 32983 2325 32992
rect 2284 32898 2324 32983
rect 2476 32864 2516 33403
rect 2476 31697 2516 32824
rect 2572 31865 2612 33664
rect 2668 34208 2708 34217
rect 2668 32201 2708 34168
rect 2764 32360 2804 35923
rect 2860 34628 2900 41728
rect 2956 40676 2996 42928
rect 3052 41264 3092 41273
rect 3052 40853 3092 41224
rect 3051 40844 3093 40853
rect 3051 40804 3052 40844
rect 3092 40804 3093 40844
rect 3051 40795 3093 40804
rect 2956 40636 3092 40676
rect 2955 40508 2997 40517
rect 2955 40468 2956 40508
rect 2996 40468 2997 40508
rect 2955 40459 2997 40468
rect 2956 39752 2996 40459
rect 2956 38912 2996 39712
rect 2956 38333 2996 38872
rect 3052 38417 3092 40636
rect 3148 40433 3188 42928
rect 3244 41012 3284 41021
rect 3147 40424 3189 40433
rect 3147 40384 3148 40424
rect 3188 40384 3189 40424
rect 3147 40375 3189 40384
rect 3244 40349 3284 40972
rect 3340 40592 3380 42928
rect 3435 41264 3477 41273
rect 3435 41224 3436 41264
rect 3476 41224 3477 41264
rect 3435 41215 3477 41224
rect 3436 41130 3476 41215
rect 3532 40769 3572 42928
rect 3724 41021 3764 42928
rect 3916 42197 3956 42928
rect 4108 42281 4148 42928
rect 4107 42272 4149 42281
rect 4107 42232 4108 42272
rect 4148 42232 4149 42272
rect 4107 42223 4149 42232
rect 3915 42188 3957 42197
rect 3915 42148 3916 42188
rect 3956 42148 3957 42188
rect 3915 42139 3957 42148
rect 4107 41768 4149 41777
rect 4107 41728 4108 41768
rect 4148 41728 4149 41768
rect 4107 41719 4149 41728
rect 3723 41012 3765 41021
rect 3723 40972 3724 41012
rect 3764 40972 3765 41012
rect 3723 40963 3765 40972
rect 3688 40844 4056 40853
rect 3728 40804 3770 40844
rect 3810 40804 3852 40844
rect 3892 40804 3934 40844
rect 3974 40804 4016 40844
rect 3688 40795 4056 40804
rect 3531 40760 3573 40769
rect 3531 40720 3532 40760
rect 3572 40720 3573 40760
rect 3531 40711 3573 40720
rect 3916 40676 3956 40685
rect 4108 40676 4148 41719
rect 4300 40937 4340 42928
rect 4492 42113 4532 42928
rect 4491 42104 4533 42113
rect 4491 42064 4492 42104
rect 4532 42064 4533 42104
rect 4491 42055 4533 42064
rect 4684 41432 4724 42928
rect 4876 42533 4916 42928
rect 4875 42524 4917 42533
rect 4875 42484 4876 42524
rect 4916 42484 4917 42524
rect 4875 42475 4917 42484
rect 5068 41768 5108 42928
rect 5260 41945 5300 42928
rect 5259 41936 5301 41945
rect 5259 41896 5260 41936
rect 5300 41896 5301 41936
rect 5259 41887 5301 41896
rect 5068 41728 5396 41768
rect 4928 41600 5296 41609
rect 4968 41560 5010 41600
rect 5050 41560 5092 41600
rect 5132 41560 5174 41600
rect 5214 41560 5256 41600
rect 4928 41551 5296 41560
rect 4588 41392 4724 41432
rect 4299 40928 4341 40937
rect 4299 40888 4300 40928
rect 4340 40888 4341 40928
rect 4299 40879 4341 40888
rect 3956 40636 4148 40676
rect 3916 40627 3956 40636
rect 3531 40592 3573 40601
rect 3340 40552 3476 40592
rect 3340 40424 3380 40433
rect 3243 40340 3285 40349
rect 3243 40300 3244 40340
rect 3284 40300 3285 40340
rect 3243 40291 3285 40300
rect 3340 40265 3380 40384
rect 3339 40256 3381 40265
rect 3339 40216 3340 40256
rect 3380 40216 3381 40256
rect 3339 40207 3381 40216
rect 3340 39845 3380 40207
rect 3339 39836 3381 39845
rect 3339 39796 3340 39836
rect 3380 39796 3381 39836
rect 3339 39787 3381 39796
rect 3340 39668 3380 39677
rect 3148 39500 3188 39509
rect 3188 39460 3284 39500
rect 3148 39451 3188 39460
rect 3148 38744 3188 38753
rect 3051 38408 3093 38417
rect 3051 38368 3052 38408
rect 3092 38368 3093 38408
rect 3051 38359 3093 38368
rect 2955 38324 2997 38333
rect 2955 38284 2956 38324
rect 2996 38284 2997 38324
rect 2955 38275 2997 38284
rect 2956 38156 2996 38165
rect 2956 37400 2996 38116
rect 3052 38156 3092 38167
rect 3052 38081 3092 38116
rect 3051 38072 3093 38081
rect 3051 38032 3052 38072
rect 3092 38032 3093 38072
rect 3051 38023 3093 38032
rect 2956 37325 2996 37360
rect 3052 37400 3092 38023
rect 3148 37829 3188 38704
rect 3147 37820 3189 37829
rect 3147 37780 3148 37820
rect 3188 37780 3189 37820
rect 3147 37771 3189 37780
rect 2955 37316 2997 37325
rect 2955 37276 2956 37316
rect 2996 37276 2997 37316
rect 2955 37267 2997 37276
rect 3052 35309 3092 37360
rect 3051 35300 3093 35309
rect 3051 35260 3052 35300
rect 3092 35260 3093 35300
rect 3051 35251 3093 35260
rect 2956 35216 2996 35225
rect 2956 35141 2996 35176
rect 2955 35132 2997 35141
rect 2955 35092 2956 35132
rect 2996 35092 2997 35132
rect 2955 35083 2997 35092
rect 2956 34796 2996 35083
rect 2956 34756 3092 34796
rect 2956 34628 2996 34637
rect 2860 34588 2956 34628
rect 2956 34579 2996 34588
rect 2967 33699 3007 33700
rect 3052 33699 3092 34756
rect 2967 33691 3092 33699
rect 3007 33659 3092 33691
rect 2967 33642 3007 33651
rect 3052 33545 3092 33659
rect 3148 34460 3188 34469
rect 3051 33536 3093 33545
rect 3051 33496 3052 33536
rect 3092 33496 3093 33536
rect 3051 33487 3093 33496
rect 2955 33032 2997 33041
rect 2955 32992 2956 33032
rect 2996 32992 2997 33032
rect 2955 32983 2997 32992
rect 2859 32444 2901 32453
rect 2859 32404 2860 32444
rect 2900 32404 2901 32444
rect 2859 32395 2901 32404
rect 2764 32311 2804 32320
rect 2667 32192 2709 32201
rect 2667 32152 2668 32192
rect 2708 32152 2709 32192
rect 2667 32143 2709 32152
rect 2860 32024 2900 32395
rect 2956 32187 2996 32983
rect 3148 32873 3188 34420
rect 3244 33699 3284 39460
rect 3340 38744 3380 39628
rect 3340 38501 3380 38704
rect 3339 38492 3381 38501
rect 3339 38452 3340 38492
rect 3380 38452 3381 38492
rect 3339 38443 3381 38452
rect 3339 38324 3381 38333
rect 3339 38284 3340 38324
rect 3380 38284 3381 38324
rect 3339 38275 3381 38284
rect 3340 35897 3380 38275
rect 3436 36140 3476 40552
rect 3531 40552 3532 40592
rect 3572 40552 3573 40592
rect 3531 40543 3573 40552
rect 3532 40458 3572 40543
rect 3627 40508 3669 40517
rect 3627 40468 3628 40508
rect 3668 40468 3669 40508
rect 3627 40459 3669 40468
rect 3724 40508 3764 40517
rect 3764 40468 3860 40508
rect 3724 40459 3764 40468
rect 3532 39920 3572 39929
rect 3628 39920 3668 40459
rect 3572 39880 3668 39920
rect 3532 39871 3572 39880
rect 3820 39584 3860 40468
rect 4108 40424 4148 40433
rect 4011 40340 4053 40349
rect 4011 40300 4012 40340
rect 4052 40300 4053 40340
rect 4011 40291 4053 40300
rect 3820 39509 3860 39544
rect 3819 39500 3861 39509
rect 3819 39460 3820 39500
rect 3860 39460 3861 39500
rect 4012 39500 4052 40291
rect 4108 39677 4148 40384
rect 4396 39752 4436 39761
rect 4107 39668 4149 39677
rect 4107 39628 4108 39668
rect 4148 39628 4149 39668
rect 4107 39619 4149 39628
rect 4396 39593 4436 39712
rect 4491 39668 4533 39677
rect 4491 39628 4492 39668
rect 4532 39628 4533 39668
rect 4491 39619 4533 39628
rect 4395 39584 4437 39593
rect 4395 39544 4396 39584
rect 4436 39544 4437 39584
rect 4395 39535 4437 39544
rect 4012 39460 4148 39500
rect 3819 39451 3861 39460
rect 3688 39332 4056 39341
rect 3728 39292 3770 39332
rect 3810 39292 3852 39332
rect 3892 39292 3934 39332
rect 3974 39292 4016 39332
rect 3688 39283 4056 39292
rect 4011 39164 4053 39173
rect 4011 39124 4012 39164
rect 4052 39124 4053 39164
rect 4011 39115 4053 39124
rect 3436 36091 3476 36100
rect 3532 38240 3572 38249
rect 3532 37400 3572 38200
rect 4012 38235 4052 39115
rect 4012 38186 4052 38195
rect 3688 37820 4056 37829
rect 3728 37780 3770 37820
rect 3810 37780 3852 37820
rect 3892 37780 3934 37820
rect 3974 37780 4016 37820
rect 3688 37771 4056 37780
rect 3915 37652 3957 37661
rect 3915 37612 3916 37652
rect 3956 37612 3957 37652
rect 3915 37603 3957 37612
rect 3339 35888 3381 35897
rect 3339 35848 3340 35888
rect 3380 35848 3381 35888
rect 3339 35839 3381 35848
rect 3340 34637 3380 35839
rect 3436 35202 3476 35211
rect 3339 34628 3381 34637
rect 3339 34588 3340 34628
rect 3380 34588 3381 34628
rect 3339 34579 3381 34588
rect 3436 34553 3476 35162
rect 3532 35141 3572 37360
rect 3916 37316 3956 37603
rect 4108 37484 4148 39460
rect 4395 39416 4437 39425
rect 4395 39376 4396 39416
rect 4436 39376 4437 39416
rect 4395 39367 4437 39376
rect 4396 39080 4436 39367
rect 4396 39031 4436 39040
rect 4204 38996 4244 39005
rect 4204 38501 4244 38956
rect 4492 38828 4532 39619
rect 4396 38788 4532 38828
rect 4203 38492 4245 38501
rect 4203 38452 4204 38492
rect 4244 38452 4245 38492
rect 4203 38443 4245 38452
rect 4060 37444 4148 37484
rect 4204 38324 4244 38333
rect 4060 37442 4100 37444
rect 4204 37409 4244 38284
rect 4060 37393 4100 37402
rect 4203 37400 4245 37409
rect 4203 37360 4204 37400
rect 4244 37360 4245 37400
rect 4203 37351 4245 37360
rect 3916 37276 4148 37316
rect 3819 36896 3861 36905
rect 3819 36856 3820 36896
rect 3860 36856 3861 36896
rect 3819 36847 3861 36856
rect 3820 36762 3860 36847
rect 3688 36308 4056 36317
rect 3728 36268 3770 36308
rect 3810 36268 3852 36308
rect 3892 36268 3934 36308
rect 3974 36268 4016 36308
rect 3688 36259 4056 36268
rect 4011 36140 4053 36149
rect 4011 36100 4012 36140
rect 4052 36100 4053 36140
rect 4011 36091 4053 36100
rect 3819 36056 3861 36065
rect 3819 36016 3820 36056
rect 3860 36016 3861 36056
rect 3819 36007 3861 36016
rect 3627 35972 3669 35981
rect 3627 35932 3628 35972
rect 3668 35932 3669 35972
rect 3627 35923 3669 35932
rect 3820 35972 3860 36007
rect 4012 36006 4052 36091
rect 3628 35838 3668 35923
rect 3820 35921 3860 35932
rect 4108 35888 4148 37276
rect 4204 37232 4244 37241
rect 4204 36821 4244 37192
rect 4203 36812 4245 36821
rect 4203 36772 4204 36812
rect 4244 36772 4245 36812
rect 4396 36812 4436 38788
rect 4491 37736 4533 37745
rect 4491 37696 4492 37736
rect 4532 37696 4533 37736
rect 4491 37687 4533 37696
rect 4492 37484 4532 37687
rect 4492 37241 4532 37444
rect 4491 37232 4533 37241
rect 4491 37192 4492 37232
rect 4532 37192 4533 37232
rect 4491 37183 4533 37192
rect 4588 36896 4628 41392
rect 4684 41264 4724 41273
rect 4684 40433 4724 41224
rect 4876 41012 4916 41021
rect 4780 40972 4876 41012
rect 4683 40424 4725 40433
rect 4683 40384 4684 40424
rect 4724 40384 4725 40424
rect 4683 40375 4725 40384
rect 4780 38240 4820 40972
rect 4876 40963 4916 40972
rect 5259 41012 5301 41021
rect 5259 40972 5260 41012
rect 5300 40972 5301 41012
rect 5259 40963 5301 40972
rect 5260 40256 5300 40963
rect 5356 40769 5396 41728
rect 5355 40760 5397 40769
rect 5355 40720 5356 40760
rect 5396 40720 5397 40760
rect 5355 40711 5397 40720
rect 5356 40433 5396 40518
rect 5355 40424 5397 40433
rect 5355 40384 5356 40424
rect 5396 40384 5397 40424
rect 5355 40375 5397 40384
rect 5260 40216 5396 40256
rect 4928 40088 5296 40097
rect 4968 40048 5010 40088
rect 5050 40048 5092 40088
rect 5132 40048 5174 40088
rect 5214 40048 5256 40088
rect 4928 40039 5296 40048
rect 5259 39920 5301 39929
rect 5259 39880 5260 39920
rect 5300 39880 5301 39920
rect 5259 39871 5301 39880
rect 4971 39836 5013 39845
rect 4971 39796 4972 39836
rect 5012 39796 5013 39836
rect 4971 39787 5013 39796
rect 4972 39173 5012 39787
rect 4971 39164 5013 39173
rect 4971 39124 4972 39164
rect 5012 39124 5013 39164
rect 4971 39115 5013 39124
rect 5260 38753 5300 39871
rect 5259 38744 5301 38753
rect 5259 38704 5260 38744
rect 5300 38704 5301 38744
rect 5259 38695 5301 38704
rect 5356 38669 5396 40216
rect 5355 38660 5397 38669
rect 5355 38620 5356 38660
rect 5396 38620 5397 38660
rect 5355 38611 5397 38620
rect 4928 38576 5296 38585
rect 4968 38536 5010 38576
rect 5050 38536 5092 38576
rect 5132 38536 5174 38576
rect 5214 38536 5256 38576
rect 4928 38527 5296 38536
rect 5452 38408 5492 42928
rect 5644 42104 5684 42928
rect 5548 42064 5684 42104
rect 5548 40853 5588 42064
rect 5643 41936 5685 41945
rect 5643 41896 5644 41936
rect 5684 41896 5685 41936
rect 5643 41887 5685 41896
rect 5547 40844 5589 40853
rect 5547 40804 5548 40844
rect 5588 40804 5589 40844
rect 5547 40795 5589 40804
rect 5547 40340 5589 40349
rect 5547 40300 5548 40340
rect 5588 40300 5589 40340
rect 5547 40291 5589 40300
rect 5548 40206 5588 40291
rect 5547 40088 5589 40097
rect 5547 40048 5548 40088
rect 5588 40048 5589 40088
rect 5547 40039 5589 40048
rect 5164 38368 5492 38408
rect 4780 38191 4820 38200
rect 4876 38240 4916 38249
rect 4876 37745 4916 38200
rect 5164 37820 5204 38368
rect 5068 37780 5204 37820
rect 5260 38156 5300 38165
rect 4875 37736 4917 37745
rect 4875 37696 4876 37736
rect 4916 37696 4917 37736
rect 4875 37687 4917 37696
rect 4683 37652 4725 37661
rect 4683 37612 4684 37652
rect 4724 37612 4725 37652
rect 4683 37603 4725 37612
rect 5068 37652 5108 37780
rect 5260 37652 5300 38116
rect 5356 38156 5396 38165
rect 5356 37829 5396 38116
rect 5355 37820 5397 37829
rect 5355 37780 5356 37820
rect 5396 37780 5397 37820
rect 5355 37771 5397 37780
rect 5452 37652 5492 37661
rect 5548 37652 5588 40039
rect 5644 39929 5684 41887
rect 5739 40592 5781 40601
rect 5739 40552 5740 40592
rect 5780 40552 5781 40592
rect 5739 40543 5781 40552
rect 5643 39920 5685 39929
rect 5643 39880 5644 39920
rect 5684 39880 5685 39920
rect 5643 39871 5685 39880
rect 5643 39752 5685 39761
rect 5643 39712 5644 39752
rect 5684 39712 5685 39752
rect 5643 39703 5685 39712
rect 5644 39618 5684 39703
rect 5740 38912 5780 40543
rect 5836 40433 5876 42928
rect 6028 40676 6068 42928
rect 6220 42617 6260 42928
rect 6219 42608 6261 42617
rect 6219 42568 6220 42608
rect 6260 42568 6261 42608
rect 6219 42559 6261 42568
rect 6219 41684 6261 41693
rect 6219 41644 6220 41684
rect 6260 41644 6261 41684
rect 6219 41635 6261 41644
rect 6124 41021 6164 41106
rect 6123 41012 6165 41021
rect 6123 40972 6124 41012
rect 6164 40972 6165 41012
rect 6123 40963 6165 40972
rect 6123 40760 6165 40769
rect 6123 40720 6124 40760
rect 6164 40720 6165 40760
rect 6123 40711 6165 40720
rect 5932 40636 6068 40676
rect 5835 40424 5877 40433
rect 5835 40384 5836 40424
rect 5876 40384 5877 40424
rect 5835 40375 5877 40384
rect 5932 40097 5972 40636
rect 6028 40508 6068 40517
rect 5931 40088 5973 40097
rect 5931 40048 5932 40088
rect 5972 40048 5973 40088
rect 5931 40039 5973 40048
rect 6028 39584 6068 40468
rect 5835 39500 5877 39509
rect 5835 39460 5836 39500
rect 5876 39460 5877 39500
rect 5835 39451 5877 39460
rect 5836 39366 5876 39451
rect 5836 38912 5876 38921
rect 5740 38872 5836 38912
rect 5836 38863 5876 38872
rect 5931 38912 5973 38921
rect 5931 38872 5932 38912
rect 5972 38872 5973 38912
rect 5931 38863 5973 38872
rect 5932 38778 5972 38863
rect 5835 38660 5877 38669
rect 5835 38620 5836 38660
rect 5876 38620 5877 38660
rect 5835 38611 5877 38620
rect 5836 38240 5876 38611
rect 5836 38191 5876 38200
rect 5260 37612 5396 37652
rect 5068 37603 5108 37612
rect 4684 37518 4724 37603
rect 4875 37568 4917 37577
rect 4875 37528 4876 37568
rect 4916 37528 4917 37568
rect 4875 37519 4917 37528
rect 4876 37484 4916 37519
rect 4876 37433 4916 37444
rect 5259 37484 5301 37493
rect 5259 37444 5260 37484
rect 5300 37444 5301 37484
rect 5259 37435 5301 37444
rect 5260 37350 5300 37435
rect 4928 37064 5296 37073
rect 4968 37024 5010 37064
rect 5050 37024 5092 37064
rect 5132 37024 5174 37064
rect 5214 37024 5256 37064
rect 4928 37015 5296 37024
rect 4684 36896 4724 36905
rect 4588 36856 4684 36896
rect 4684 36847 4724 36856
rect 4971 36896 5013 36905
rect 4971 36856 4972 36896
rect 5012 36856 5013 36896
rect 4971 36847 5013 36856
rect 4396 36772 4628 36812
rect 4203 36763 4245 36772
rect 4300 36644 4340 36653
rect 4300 36560 4340 36604
rect 4492 36644 4532 36653
rect 4492 36560 4532 36604
rect 4300 36520 4532 36560
rect 4299 36056 4341 36065
rect 4299 36016 4300 36056
rect 4340 36016 4341 36056
rect 4299 36007 4341 36016
rect 3916 35848 4148 35888
rect 3628 35300 3668 35309
rect 3531 35132 3573 35141
rect 3531 35092 3532 35132
rect 3572 35092 3573 35132
rect 3531 35083 3573 35092
rect 3628 34973 3668 35260
rect 3916 35216 3956 35848
rect 3916 35167 3956 35176
rect 4011 35216 4053 35225
rect 4011 35176 4012 35216
rect 4052 35176 4053 35216
rect 4011 35167 4053 35176
rect 4012 35082 4052 35167
rect 4107 35048 4149 35057
rect 4107 35008 4108 35048
rect 4148 35008 4149 35048
rect 4107 34999 4149 35008
rect 3627 34964 3669 34973
rect 3627 34924 3628 34964
rect 3668 34924 3669 34964
rect 3627 34915 3669 34924
rect 3688 34796 4056 34805
rect 3728 34756 3770 34796
rect 3810 34756 3852 34796
rect 3892 34756 3934 34796
rect 3974 34756 4016 34796
rect 3688 34747 4056 34756
rect 3435 34544 3477 34553
rect 3435 34504 3436 34544
rect 3476 34504 3477 34544
rect 3435 34495 3477 34504
rect 3915 34460 3957 34469
rect 3915 34420 3916 34460
rect 3956 34420 3957 34460
rect 3915 34411 3957 34420
rect 3339 34376 3381 34385
rect 3339 34336 3340 34376
rect 3380 34336 3381 34376
rect 3339 34327 3381 34336
rect 3436 34376 3476 34385
rect 3340 34242 3380 34327
rect 3436 34133 3476 34336
rect 3628 34376 3668 34385
rect 3531 34208 3573 34217
rect 3531 34168 3532 34208
rect 3572 34168 3573 34208
rect 3531 34159 3573 34168
rect 3435 34124 3477 34133
rect 3435 34084 3436 34124
rect 3476 34084 3477 34124
rect 3435 34075 3477 34084
rect 3532 34074 3572 34159
rect 3628 33965 3668 34336
rect 3627 33956 3669 33965
rect 3627 33916 3628 33956
rect 3668 33916 3669 33956
rect 3627 33907 3669 33916
rect 3916 33872 3956 34411
rect 4108 34376 4148 34999
rect 4204 34376 4244 34385
rect 4108 34336 4204 34376
rect 4204 34327 4244 34336
rect 3916 33823 3956 33832
rect 3628 33788 3668 33797
rect 3532 33748 3628 33788
rect 3436 33699 3476 33708
rect 3244 33659 3436 33699
rect 3436 33650 3476 33659
rect 3147 32864 3189 32873
rect 3147 32824 3148 32864
rect 3188 32824 3189 32864
rect 3147 32815 3189 32824
rect 3339 32612 3381 32621
rect 3339 32572 3340 32612
rect 3380 32572 3381 32612
rect 3339 32563 3381 32572
rect 2956 32138 2996 32147
rect 2764 31984 2900 32024
rect 2571 31856 2613 31865
rect 2571 31816 2572 31856
rect 2612 31816 2613 31856
rect 2571 31807 2613 31816
rect 2475 31688 2517 31697
rect 2475 31648 2476 31688
rect 2516 31648 2517 31688
rect 2475 31639 2517 31648
rect 2187 31352 2229 31361
rect 2187 31312 2188 31352
rect 2228 31312 2229 31352
rect 2187 31303 2229 31312
rect 2475 31352 2517 31361
rect 2475 31312 2476 31352
rect 2516 31312 2517 31352
rect 2475 31303 2517 31312
rect 2091 31100 2133 31109
rect 2091 31060 2092 31100
rect 2132 31060 2133 31100
rect 2091 31051 2133 31060
rect 2188 30941 2228 31303
rect 2476 31218 2516 31303
rect 2668 31184 2708 31193
rect 2572 31144 2668 31184
rect 2187 30932 2229 30941
rect 2187 30892 2188 30932
rect 2228 30892 2229 30932
rect 2187 30883 2229 30892
rect 2572 30689 2612 31144
rect 2668 31135 2708 31144
rect 2188 30680 2228 30689
rect 2188 30596 2228 30640
rect 2379 30680 2421 30689
rect 2379 30640 2380 30680
rect 2420 30640 2421 30680
rect 2379 30631 2421 30640
rect 2476 30680 2516 30689
rect 1996 30556 2228 30596
rect 1899 28916 1941 28925
rect 1899 28876 1900 28916
rect 1940 28876 1941 28916
rect 1899 28867 1941 28876
rect 1900 28328 1940 28867
rect 1900 28279 1940 28288
rect 2188 27665 2228 30556
rect 2380 30546 2420 30631
rect 2284 30512 2324 30521
rect 2284 30101 2324 30472
rect 2476 30185 2516 30640
rect 2571 30680 2613 30689
rect 2571 30640 2572 30680
rect 2612 30640 2613 30680
rect 2571 30631 2613 30640
rect 2668 30680 2708 30689
rect 2764 30680 2804 31984
rect 2859 31856 2901 31865
rect 2859 31816 2860 31856
rect 2900 31816 2901 31856
rect 2859 31807 2901 31816
rect 2708 30640 2804 30680
rect 2860 31352 2900 31807
rect 3052 31352 3092 31361
rect 2860 31312 3052 31352
rect 2668 30631 2708 30640
rect 2860 30596 2900 31312
rect 3052 31303 3092 31312
rect 3051 31184 3093 31193
rect 3051 31144 3052 31184
rect 3092 31144 3093 31184
rect 3051 31135 3093 31144
rect 3148 31184 3188 31193
rect 3188 31144 3284 31184
rect 3148 31135 3188 31144
rect 2955 30680 2997 30689
rect 2955 30640 2956 30680
rect 2996 30640 2997 30680
rect 2955 30631 2997 30640
rect 2764 30556 2900 30596
rect 2475 30176 2517 30185
rect 2475 30136 2476 30176
rect 2516 30136 2517 30176
rect 2475 30127 2517 30136
rect 2667 30176 2709 30185
rect 2667 30136 2668 30176
rect 2708 30136 2709 30176
rect 2667 30127 2709 30136
rect 2283 30092 2325 30101
rect 2283 30052 2284 30092
rect 2324 30052 2325 30092
rect 2283 30043 2325 30052
rect 2668 30008 2708 30127
rect 2668 29959 2708 29968
rect 2475 29840 2517 29849
rect 2475 29800 2476 29840
rect 2516 29800 2517 29840
rect 2475 29791 2517 29800
rect 2476 29706 2516 29791
rect 2764 29672 2804 30556
rect 2859 30092 2901 30101
rect 2859 30052 2860 30092
rect 2900 30052 2901 30092
rect 2859 30043 2901 30052
rect 2860 29840 2900 30043
rect 2860 29791 2900 29800
rect 2956 29840 2996 30631
rect 2956 29791 2996 29800
rect 3052 29672 3092 31135
rect 3148 29840 3188 29849
rect 3148 29681 3188 29800
rect 3244 29840 3284 31144
rect 3340 31025 3380 32563
rect 3436 32192 3476 32201
rect 3436 31193 3476 32152
rect 3532 32117 3572 33748
rect 3628 33739 3668 33748
rect 4203 33704 4245 33713
rect 4203 33664 4204 33704
rect 4244 33664 4245 33704
rect 4203 33655 4245 33664
rect 4204 33570 4244 33655
rect 4203 33368 4245 33377
rect 4203 33328 4204 33368
rect 4244 33328 4245 33368
rect 4203 33319 4245 33328
rect 3688 33284 4056 33293
rect 3728 33244 3770 33284
rect 3810 33244 3852 33284
rect 3892 33244 3934 33284
rect 3974 33244 4016 33284
rect 3688 33235 4056 33244
rect 4011 33116 4053 33125
rect 4011 33076 4012 33116
rect 4052 33076 4053 33116
rect 4011 33067 4053 33076
rect 3724 32864 3764 32873
rect 3724 32621 3764 32824
rect 4012 32864 4052 33067
rect 4012 32815 4052 32824
rect 3723 32612 3765 32621
rect 3723 32572 3724 32612
rect 3764 32572 3765 32612
rect 3723 32563 3765 32572
rect 3531 32108 3573 32117
rect 3531 32068 3532 32108
rect 3572 32068 3573 32108
rect 3531 32059 3573 32068
rect 3915 32108 3957 32117
rect 3915 32068 3916 32108
rect 3956 32068 3957 32108
rect 3915 32059 3957 32068
rect 4012 32108 4052 32117
rect 4052 32068 4148 32108
rect 4012 32059 4052 32068
rect 3916 31974 3956 32059
rect 3688 31772 4056 31781
rect 3728 31732 3770 31772
rect 3810 31732 3852 31772
rect 3892 31732 3934 31772
rect 3974 31732 4016 31772
rect 3688 31723 4056 31732
rect 3531 31688 3573 31697
rect 3531 31648 3532 31688
rect 3572 31648 3573 31688
rect 3531 31639 3573 31648
rect 3435 31184 3477 31193
rect 3435 31144 3436 31184
rect 3476 31144 3477 31184
rect 3435 31135 3477 31144
rect 3339 31016 3381 31025
rect 3339 30976 3340 31016
rect 3380 30976 3381 31016
rect 3339 30967 3381 30976
rect 3435 30932 3477 30941
rect 3435 30892 3436 30932
rect 3476 30892 3477 30932
rect 3435 30883 3477 30892
rect 3339 30176 3381 30185
rect 3339 30136 3340 30176
rect 3380 30136 3381 30176
rect 3339 30127 3381 30136
rect 3340 29849 3380 30127
rect 3340 29840 3386 29849
rect 3340 29800 3345 29840
rect 3385 29800 3386 29840
rect 3244 29791 3284 29800
rect 3344 29791 3386 29800
rect 3345 29706 3385 29791
rect 2764 29632 2900 29672
rect 2763 29252 2805 29261
rect 2763 29212 2764 29252
rect 2804 29212 2805 29252
rect 2763 29203 2805 29212
rect 2764 29168 2804 29203
rect 2764 29117 2804 29128
rect 2763 28412 2805 28421
rect 2763 28372 2764 28412
rect 2804 28372 2805 28412
rect 2763 28363 2805 28372
rect 1995 27656 2037 27665
rect 1995 27616 1996 27656
rect 2036 27616 2037 27656
rect 1995 27607 2037 27616
rect 2187 27656 2229 27665
rect 2187 27616 2188 27656
rect 2228 27616 2229 27656
rect 2187 27607 2229 27616
rect 2476 27656 2516 27665
rect 1803 26816 1845 26825
rect 1803 26776 1804 26816
rect 1844 26776 1845 26816
rect 1803 26767 1845 26776
rect 1708 25255 1748 25264
rect 1611 25052 1653 25061
rect 1611 25012 1612 25052
rect 1652 25012 1653 25052
rect 1611 25003 1653 25012
rect 1515 24632 1557 24641
rect 1515 24592 1516 24632
rect 1556 24592 1557 24632
rect 1515 24583 1557 24592
rect 1611 23960 1653 23969
rect 1611 23920 1612 23960
rect 1652 23920 1653 23960
rect 1611 23911 1653 23920
rect 1419 23876 1461 23885
rect 1419 23836 1420 23876
rect 1460 23836 1461 23876
rect 1419 23827 1461 23836
rect 1419 23120 1461 23129
rect 1419 23080 1420 23120
rect 1460 23080 1556 23120
rect 1419 23071 1461 23080
rect 1420 22986 1460 23071
rect 1420 22280 1460 22289
rect 1324 22240 1420 22280
rect 1420 22231 1460 22240
rect 1228 22156 1364 22196
rect 1324 20096 1364 22156
rect 1516 22037 1556 23080
rect 1515 22028 1557 22037
rect 1515 21988 1516 22028
rect 1556 21988 1557 22028
rect 1515 21979 1557 21988
rect 1612 20768 1652 23911
rect 1804 23633 1844 26767
rect 1899 24632 1941 24641
rect 1899 24592 1900 24632
rect 1940 24592 1941 24632
rect 1899 24583 1941 24592
rect 1803 23624 1845 23633
rect 1803 23584 1804 23624
rect 1844 23584 1845 23624
rect 1803 23575 1845 23584
rect 1803 21944 1845 21953
rect 1803 21904 1804 21944
rect 1844 21904 1845 21944
rect 1803 21895 1845 21904
rect 1612 20719 1652 20728
rect 1516 20096 1556 20105
rect 1324 20056 1516 20096
rect 1323 19424 1365 19433
rect 1323 19384 1324 19424
rect 1364 19384 1365 19424
rect 1323 19375 1365 19384
rect 1228 19256 1268 19265
rect 1324 19256 1364 19375
rect 1268 19216 1364 19256
rect 1228 19207 1268 19216
rect 1419 17492 1461 17501
rect 1419 17452 1420 17492
rect 1460 17452 1461 17492
rect 1419 17443 1461 17452
rect 1323 17156 1365 17165
rect 1228 17116 1324 17156
rect 1364 17116 1365 17156
rect 1228 17072 1268 17116
rect 1323 17107 1365 17116
rect 1228 17023 1268 17032
rect 1131 16400 1173 16409
rect 1131 16360 1132 16400
rect 1172 16360 1173 16400
rect 1131 16351 1173 16360
rect 1420 16232 1460 17443
rect 1420 16183 1460 16192
rect 1228 15560 1268 15569
rect 1323 15560 1365 15569
rect 1268 15520 1324 15560
rect 1364 15520 1365 15560
rect 1228 15511 1268 15520
rect 1323 15511 1365 15520
rect 1323 15056 1365 15065
rect 1323 15016 1324 15056
rect 1364 15016 1365 15056
rect 1323 15007 1365 15016
rect 1228 14720 1268 14729
rect 1324 14720 1364 15007
rect 1268 14680 1364 14720
rect 1228 14671 1268 14680
rect 1516 13973 1556 20056
rect 1707 16652 1749 16661
rect 1707 16612 1708 16652
rect 1748 16612 1749 16652
rect 1707 16603 1749 16612
rect 1611 14132 1653 14141
rect 1611 14092 1612 14132
rect 1652 14092 1653 14132
rect 1611 14083 1653 14092
rect 1515 13964 1557 13973
rect 1515 13924 1516 13964
rect 1556 13924 1557 13964
rect 1515 13915 1557 13924
rect 939 13124 981 13133
rect 939 13084 940 13124
rect 980 13084 981 13124
rect 939 13075 981 13084
rect 1323 11864 1365 11873
rect 1323 11824 1324 11864
rect 1364 11824 1365 11864
rect 1323 11815 1365 11824
rect 1228 11696 1268 11705
rect 1324 11696 1364 11815
rect 1268 11656 1364 11696
rect 1228 11647 1268 11656
rect 1419 11528 1461 11537
rect 1419 11488 1420 11528
rect 1460 11488 1461 11528
rect 1419 11479 1461 11488
rect 1227 11024 1269 11033
rect 1227 10984 1228 11024
rect 1268 10984 1269 11024
rect 1227 10975 1269 10984
rect 1228 10890 1268 10975
rect 1323 10940 1365 10949
rect 1323 10900 1324 10940
rect 1364 10900 1365 10940
rect 1323 10891 1365 10900
rect 1227 10184 1269 10193
rect 1227 10144 1228 10184
rect 1268 10144 1269 10184
rect 1227 10135 1269 10144
rect 1228 10050 1268 10135
rect 1228 8672 1268 8681
rect 1324 8672 1364 10891
rect 1268 8632 1364 8672
rect 1228 8623 1268 8632
rect 1324 7841 1364 8632
rect 1323 7832 1365 7841
rect 1323 7792 1324 7832
rect 1364 7792 1365 7832
rect 1323 7783 1365 7792
rect 651 7328 693 7337
rect 651 7288 652 7328
rect 692 7288 693 7328
rect 651 7279 693 7288
rect 1323 7244 1365 7253
rect 1228 7204 1324 7244
rect 1364 7204 1365 7244
rect 1228 7160 1268 7204
rect 1323 7195 1365 7204
rect 1228 7111 1268 7120
rect 1323 7076 1365 7085
rect 1323 7036 1324 7076
rect 1364 7036 1365 7076
rect 1323 7027 1365 7036
rect 1228 6488 1268 6497
rect 1324 6488 1364 7027
rect 1268 6448 1364 6488
rect 1228 6439 1268 6448
rect 1228 4976 1268 4985
rect 1268 4936 1364 4976
rect 1228 4927 1268 4936
rect 1324 4733 1364 4936
rect 1323 4724 1365 4733
rect 1323 4684 1324 4724
rect 1364 4684 1365 4724
rect 1323 4675 1365 4684
rect 1323 4304 1365 4313
rect 1323 4264 1324 4304
rect 1364 4264 1365 4304
rect 1323 4255 1365 4264
rect 1228 4136 1268 4145
rect 1324 4136 1364 4255
rect 1268 4096 1364 4136
rect 1228 4087 1268 4096
rect 1420 3221 1460 11479
rect 1612 11117 1652 14083
rect 1708 13889 1748 16603
rect 1707 13880 1749 13889
rect 1707 13840 1708 13880
rect 1748 13840 1749 13880
rect 1707 13831 1749 13840
rect 1611 11108 1653 11117
rect 1611 11068 1612 11108
rect 1652 11068 1653 11108
rect 1611 11059 1653 11068
rect 1612 10277 1652 11059
rect 1611 10268 1653 10277
rect 1611 10228 1612 10268
rect 1652 10228 1653 10268
rect 1611 10219 1653 10228
rect 1611 9764 1653 9773
rect 1611 9724 1612 9764
rect 1652 9724 1653 9764
rect 1611 9715 1653 9724
rect 1516 9512 1556 9521
rect 1516 6581 1556 9472
rect 1515 6572 1557 6581
rect 1515 6532 1516 6572
rect 1556 6532 1557 6572
rect 1515 6523 1557 6532
rect 1515 6068 1557 6077
rect 1515 6028 1516 6068
rect 1556 6028 1557 6068
rect 1515 6019 1557 6028
rect 1516 5900 1556 6019
rect 1516 5851 1556 5860
rect 1419 3212 1461 3221
rect 1419 3172 1420 3212
rect 1460 3172 1461 3212
rect 1419 3163 1461 3172
rect 1612 3137 1652 9715
rect 1804 8849 1844 21895
rect 1900 19433 1940 24583
rect 1899 19424 1941 19433
rect 1899 19384 1900 19424
rect 1940 19384 1941 19424
rect 1899 19375 1941 19384
rect 1899 18752 1941 18761
rect 1899 18712 1900 18752
rect 1940 18712 1941 18752
rect 1899 18703 1941 18712
rect 1900 15569 1940 18703
rect 1899 15560 1941 15569
rect 1899 15520 1900 15560
rect 1940 15520 1941 15560
rect 1899 15511 1941 15520
rect 1900 10949 1940 15511
rect 1899 10940 1941 10949
rect 1899 10900 1900 10940
rect 1940 10900 1941 10940
rect 1899 10891 1941 10900
rect 1803 8840 1845 8849
rect 1803 8800 1804 8840
rect 1844 8800 1845 8840
rect 1803 8791 1845 8800
rect 1996 8672 2036 27607
rect 2187 27236 2229 27245
rect 2187 27196 2188 27236
rect 2228 27196 2229 27236
rect 2187 27187 2229 27196
rect 2091 25052 2133 25061
rect 2091 25012 2092 25052
rect 2132 25012 2133 25052
rect 2091 25003 2133 25012
rect 2092 19601 2132 25003
rect 2188 23792 2228 27187
rect 2476 27161 2516 27616
rect 2571 27656 2613 27665
rect 2571 27616 2572 27656
rect 2612 27616 2613 27656
rect 2571 27607 2613 27616
rect 2572 27522 2612 27607
rect 2475 27152 2517 27161
rect 2475 27112 2476 27152
rect 2516 27112 2517 27152
rect 2475 27103 2517 27112
rect 2667 27152 2709 27161
rect 2667 27112 2668 27152
rect 2708 27112 2709 27152
rect 2667 27103 2709 27112
rect 2668 27068 2708 27103
rect 2668 27017 2708 27028
rect 2475 26816 2517 26825
rect 2475 26776 2476 26816
rect 2516 26776 2517 26816
rect 2475 26767 2517 26776
rect 2476 26682 2516 26767
rect 2379 24968 2421 24977
rect 2379 24928 2380 24968
rect 2420 24928 2421 24968
rect 2379 24919 2421 24928
rect 2380 23969 2420 24919
rect 2764 24809 2804 28363
rect 2860 27656 2900 29632
rect 3052 29623 3092 29632
rect 3147 29672 3189 29681
rect 3147 29632 3148 29672
rect 3188 29632 3189 29672
rect 3147 29623 3189 29632
rect 3436 29588 3476 30883
rect 3340 29548 3476 29588
rect 2956 28916 2996 28925
rect 2956 28337 2996 28876
rect 3340 28421 3380 29548
rect 3532 29261 3572 31639
rect 4108 31352 4148 32068
rect 4012 31312 4148 31352
rect 4204 31352 4244 33319
rect 4300 31529 4340 36007
rect 4492 35729 4532 36520
rect 4491 35720 4533 35729
rect 4491 35680 4492 35720
rect 4532 35680 4533 35720
rect 4491 35671 4533 35680
rect 4492 35586 4532 35671
rect 4396 35132 4436 35141
rect 4396 34049 4436 35092
rect 4491 35132 4533 35141
rect 4491 35092 4492 35132
rect 4532 35092 4533 35132
rect 4491 35083 4533 35092
rect 4492 34469 4532 35083
rect 4491 34460 4533 34469
rect 4491 34420 4492 34460
rect 4532 34420 4533 34460
rect 4491 34411 4533 34420
rect 4588 34301 4628 36772
rect 4972 36728 5012 36847
rect 4972 36679 5012 36688
rect 4971 35888 5013 35897
rect 4971 35848 4972 35888
rect 5012 35848 5013 35888
rect 4971 35839 5013 35848
rect 4972 35754 5012 35839
rect 4779 35720 4821 35729
rect 4779 35680 4780 35720
rect 4820 35680 4821 35720
rect 4779 35671 4821 35680
rect 4780 35586 4820 35671
rect 4683 35552 4725 35561
rect 4683 35512 4684 35552
rect 4724 35512 4725 35552
rect 4683 35503 4725 35512
rect 4928 35552 5296 35561
rect 4968 35512 5010 35552
rect 5050 35512 5092 35552
rect 5132 35512 5174 35552
rect 5214 35512 5256 35552
rect 4928 35503 5296 35512
rect 4587 34292 4629 34301
rect 4587 34252 4588 34292
rect 4628 34252 4629 34292
rect 4587 34243 4629 34252
rect 4684 34124 4724 35503
rect 4779 35384 4821 35393
rect 4779 35344 4780 35384
rect 4820 35344 4821 35384
rect 4779 35335 4821 35344
rect 4971 35384 5013 35393
rect 4971 35344 4972 35384
rect 5012 35344 5013 35384
rect 4971 35335 5013 35344
rect 4588 34084 4724 34124
rect 4395 34040 4437 34049
rect 4395 34000 4396 34040
rect 4436 34000 4437 34040
rect 4395 33991 4437 34000
rect 4395 32360 4437 32369
rect 4395 32320 4396 32360
rect 4436 32320 4437 32360
rect 4395 32311 4437 32320
rect 4396 32192 4436 32311
rect 4299 31520 4341 31529
rect 4299 31480 4300 31520
rect 4340 31480 4341 31520
rect 4396 31520 4436 32152
rect 4491 32192 4533 32201
rect 4491 32152 4492 32192
rect 4532 32152 4533 32192
rect 4491 32143 4533 32152
rect 4492 32058 4532 32143
rect 4396 31480 4532 31520
rect 4299 31471 4341 31480
rect 3916 30680 3956 30689
rect 3916 30521 3956 30640
rect 3915 30512 3957 30521
rect 3915 30472 3916 30512
rect 3956 30472 3957 30512
rect 4012 30512 4052 31312
rect 4204 31303 4244 31312
rect 4396 31352 4436 31361
rect 4108 31184 4148 31193
rect 4108 30941 4148 31144
rect 4396 31109 4436 31312
rect 4395 31100 4437 31109
rect 4395 31060 4396 31100
rect 4436 31060 4437 31100
rect 4395 31051 4437 31060
rect 4107 30932 4149 30941
rect 4107 30892 4108 30932
rect 4148 30892 4149 30932
rect 4107 30883 4149 30892
rect 4108 30764 4148 30773
rect 4148 30724 4436 30764
rect 4108 30715 4148 30724
rect 4396 30680 4436 30724
rect 4396 30631 4436 30640
rect 4492 30680 4532 31480
rect 4588 30932 4628 34084
rect 4683 33032 4725 33041
rect 4683 32992 4684 33032
rect 4724 32992 4725 33032
rect 4683 32983 4725 32992
rect 4684 31109 4724 32983
rect 4780 32360 4820 35335
rect 4972 35216 5012 35335
rect 4972 35167 5012 35176
rect 4928 34040 5296 34049
rect 4968 34000 5010 34040
rect 5050 34000 5092 34040
rect 5132 34000 5174 34040
rect 5214 34000 5256 34040
rect 4928 33991 5296 34000
rect 5259 32864 5301 32873
rect 5259 32824 5260 32864
rect 5300 32824 5301 32864
rect 5259 32815 5301 32824
rect 5260 32730 5300 32815
rect 4928 32528 5296 32537
rect 4968 32488 5010 32528
rect 5050 32488 5092 32528
rect 5132 32488 5174 32528
rect 5214 32488 5256 32528
rect 4928 32479 5296 32488
rect 4780 32311 4820 32320
rect 5356 32285 5396 37612
rect 5492 37612 5588 37652
rect 5452 37603 5492 37612
rect 5644 37400 5684 37409
rect 5684 37360 5780 37400
rect 5644 37351 5684 37360
rect 5451 35720 5493 35729
rect 5451 35680 5452 35720
rect 5492 35680 5493 35720
rect 5451 35671 5493 35680
rect 5452 35211 5492 35671
rect 5643 35300 5685 35309
rect 5643 35260 5644 35300
rect 5684 35260 5685 35300
rect 5643 35251 5685 35260
rect 5452 35162 5492 35171
rect 5644 35166 5684 35251
rect 5547 34964 5589 34973
rect 5547 34924 5548 34964
rect 5588 34924 5589 34964
rect 5547 34915 5589 34924
rect 5452 34376 5492 34385
rect 5452 33704 5492 34336
rect 5548 34049 5588 34915
rect 5740 34889 5780 37360
rect 5739 34880 5781 34889
rect 5739 34840 5740 34880
rect 5780 34840 5781 34880
rect 5739 34831 5781 34840
rect 5740 34721 5780 34831
rect 5739 34712 5781 34721
rect 5739 34672 5740 34712
rect 5780 34672 5781 34712
rect 5739 34663 5781 34672
rect 5835 34544 5877 34553
rect 5835 34504 5836 34544
rect 5876 34504 5877 34544
rect 6028 34544 6068 39544
rect 6124 37661 6164 40711
rect 6220 40676 6260 41635
rect 6220 40627 6260 40636
rect 6316 41264 6356 41273
rect 6316 40433 6356 41224
rect 6412 40601 6452 42928
rect 6411 40592 6453 40601
rect 6411 40552 6412 40592
rect 6452 40552 6453 40592
rect 6411 40543 6453 40552
rect 6315 40424 6357 40433
rect 6315 40384 6316 40424
rect 6356 40384 6357 40424
rect 6315 40375 6357 40384
rect 6412 40424 6452 40433
rect 6316 39761 6356 40375
rect 6315 39752 6357 39761
rect 6315 39712 6316 39752
rect 6356 39712 6357 39752
rect 6315 39703 6357 39712
rect 6412 39248 6452 40384
rect 6507 40340 6549 40349
rect 6507 40300 6508 40340
rect 6548 40300 6549 40340
rect 6507 40291 6549 40300
rect 6220 39208 6452 39248
rect 6220 38828 6260 39208
rect 6411 39080 6453 39089
rect 6316 39040 6412 39080
rect 6452 39040 6453 39080
rect 6316 38996 6356 39040
rect 6411 39031 6453 39040
rect 6316 38947 6356 38956
rect 6412 38912 6452 38923
rect 6412 38837 6452 38872
rect 6411 38828 6453 38837
rect 6220 38788 6356 38828
rect 6316 38333 6356 38788
rect 6411 38788 6412 38828
rect 6452 38788 6453 38828
rect 6411 38779 6453 38788
rect 6508 38492 6548 40291
rect 6412 38452 6548 38492
rect 6315 38324 6357 38333
rect 6315 38284 6316 38324
rect 6356 38284 6357 38324
rect 6315 38275 6357 38284
rect 6412 38230 6452 38452
rect 6604 38417 6644 42928
rect 6699 40424 6741 40433
rect 6699 40384 6700 40424
rect 6740 40384 6741 40424
rect 6699 40375 6741 40384
rect 6603 38408 6645 38417
rect 6603 38368 6604 38408
rect 6644 38368 6645 38408
rect 6603 38359 6645 38368
rect 6364 38198 6452 38230
rect 6404 38190 6452 38198
rect 6508 38324 6548 38333
rect 6364 38149 6404 38158
rect 6508 37820 6548 38284
rect 6508 37780 6644 37820
rect 6123 37652 6165 37661
rect 6123 37612 6124 37652
rect 6164 37612 6165 37652
rect 6123 37603 6165 37612
rect 6507 37484 6549 37493
rect 6507 37444 6508 37484
rect 6548 37444 6549 37484
rect 6507 37435 6549 37444
rect 6220 36728 6260 36737
rect 6124 36688 6220 36728
rect 6124 35384 6164 36688
rect 6220 36679 6260 36688
rect 6508 36569 6548 37435
rect 6507 36560 6549 36569
rect 6507 36520 6508 36560
rect 6548 36520 6549 36560
rect 6507 36511 6549 36520
rect 6412 36476 6452 36485
rect 6220 35888 6260 35897
rect 6412 35888 6452 36436
rect 6604 36056 6644 37780
rect 6700 37400 6740 40375
rect 6796 39173 6836 42928
rect 6988 40517 7028 42928
rect 6987 40508 7029 40517
rect 6987 40468 6988 40508
rect 7028 40468 7029 40508
rect 6987 40459 7029 40468
rect 6988 39752 7028 39761
rect 6988 39257 7028 39712
rect 6987 39248 7029 39257
rect 6987 39208 6988 39248
rect 7028 39208 7124 39248
rect 6987 39199 7029 39208
rect 6795 39164 6837 39173
rect 6795 39124 6796 39164
rect 6836 39124 6837 39164
rect 6795 39115 6837 39124
rect 6892 38912 6932 38921
rect 6932 38872 7028 38912
rect 6892 38863 6932 38872
rect 6891 38408 6933 38417
rect 6891 38368 6892 38408
rect 6932 38368 6933 38408
rect 6891 38359 6933 38368
rect 6892 38274 6932 38359
rect 6892 37400 6932 37409
rect 6700 37360 6892 37400
rect 6796 37073 6836 37360
rect 6892 37351 6932 37360
rect 6795 37064 6837 37073
rect 6795 37024 6796 37064
rect 6836 37024 6837 37064
rect 6795 37015 6837 37024
rect 6699 36560 6741 36569
rect 6699 36520 6700 36560
rect 6740 36520 6741 36560
rect 6699 36511 6741 36520
rect 6700 36426 6740 36511
rect 6604 36016 6740 36056
rect 6508 35888 6548 35897
rect 6412 35848 6508 35888
rect 6220 35468 6260 35848
rect 6508 35839 6548 35848
rect 6603 35888 6645 35897
rect 6603 35848 6604 35888
rect 6644 35848 6645 35888
rect 6603 35839 6645 35848
rect 6604 35754 6644 35839
rect 6220 35428 6452 35468
rect 6124 35344 6260 35384
rect 6220 35225 6260 35344
rect 6315 35300 6357 35309
rect 6315 35260 6316 35300
rect 6356 35260 6357 35300
rect 6315 35251 6357 35260
rect 6124 35216 6164 35225
rect 6124 34805 6164 35176
rect 6219 35216 6261 35225
rect 6219 35176 6220 35216
rect 6260 35176 6261 35216
rect 6219 35167 6261 35176
rect 6123 34796 6165 34805
rect 6123 34756 6124 34796
rect 6164 34756 6165 34796
rect 6123 34747 6165 34756
rect 6028 34504 6164 34544
rect 5835 34495 5877 34504
rect 5739 34376 5781 34385
rect 5739 34336 5740 34376
rect 5780 34336 5781 34376
rect 5739 34327 5781 34336
rect 5643 34292 5685 34301
rect 5643 34252 5644 34292
rect 5684 34252 5685 34292
rect 5643 34243 5685 34252
rect 5644 34158 5684 34243
rect 5547 34040 5589 34049
rect 5547 34000 5548 34040
rect 5588 34000 5589 34040
rect 5547 33991 5589 34000
rect 5643 33956 5685 33965
rect 5643 33916 5644 33956
rect 5684 33916 5685 33956
rect 5643 33907 5685 33916
rect 5644 33872 5684 33907
rect 5644 33821 5684 33832
rect 5492 33664 5588 33704
rect 5452 33655 5492 33664
rect 5451 33368 5493 33377
rect 5451 33328 5452 33368
rect 5492 33328 5493 33368
rect 5451 33319 5493 33328
rect 5452 33116 5492 33319
rect 5452 33067 5492 33076
rect 5451 32948 5493 32957
rect 5451 32908 5452 32948
rect 5492 32908 5493 32948
rect 5451 32899 5493 32908
rect 5355 32276 5397 32285
rect 5355 32236 5356 32276
rect 5396 32236 5397 32276
rect 5355 32227 5397 32236
rect 4971 32192 5013 32201
rect 4971 32152 4972 32192
rect 5012 32152 5013 32192
rect 4971 32143 5013 32152
rect 4779 32108 4821 32117
rect 4779 32068 4780 32108
rect 4820 32068 4821 32108
rect 4779 32059 4821 32068
rect 4683 31100 4725 31109
rect 4683 31060 4684 31100
rect 4724 31060 4725 31100
rect 4683 31051 4725 31060
rect 4588 30892 4724 30932
rect 4532 30640 4628 30680
rect 4492 30631 4532 30640
rect 4012 30472 4148 30512
rect 3915 30463 3957 30472
rect 3688 30260 4056 30269
rect 3728 30220 3770 30260
rect 3810 30220 3852 30260
rect 3892 30220 3934 30260
rect 3974 30220 4016 30260
rect 3688 30211 4056 30220
rect 3627 29840 3669 29849
rect 3627 29800 3628 29840
rect 3668 29800 3669 29840
rect 3627 29791 3669 29800
rect 3724 29840 3764 29849
rect 3628 29706 3668 29791
rect 3531 29252 3573 29261
rect 3531 29212 3532 29252
rect 3572 29212 3573 29252
rect 3531 29203 3573 29212
rect 3724 29000 3764 29800
rect 3915 29672 3957 29681
rect 3915 29632 3916 29672
rect 3956 29632 3957 29672
rect 3915 29623 3957 29632
rect 3916 29538 3956 29623
rect 3819 29420 3861 29429
rect 3819 29380 3820 29420
rect 3860 29380 3861 29420
rect 3819 29371 3861 29380
rect 3820 29168 3860 29371
rect 3820 29119 3860 29128
rect 3436 28960 3764 29000
rect 3339 28412 3381 28421
rect 3339 28372 3340 28412
rect 3380 28372 3381 28412
rect 3339 28363 3381 28372
rect 2955 28328 2997 28337
rect 2955 28288 2956 28328
rect 2996 28288 2997 28328
rect 2955 28279 2997 28288
rect 3148 28328 3188 28337
rect 2956 27656 2996 27665
rect 2860 27616 2956 27656
rect 2956 27607 2996 27616
rect 3051 27572 3093 27581
rect 3051 27532 3052 27572
rect 3092 27532 3093 27572
rect 3051 27523 3093 27532
rect 3052 27438 3092 27523
rect 2859 27236 2901 27245
rect 2859 27196 2860 27236
rect 2900 27196 2901 27236
rect 2859 27187 2901 27196
rect 2860 26825 2900 27187
rect 3148 26909 3188 28288
rect 3339 28160 3381 28169
rect 3339 28120 3340 28160
rect 3380 28120 3381 28160
rect 3339 28111 3381 28120
rect 3340 28026 3380 28111
rect 3436 27908 3476 28960
rect 3688 28748 4056 28757
rect 3728 28708 3770 28748
rect 3810 28708 3852 28748
rect 3892 28708 3934 28748
rect 3974 28708 4016 28748
rect 3688 28699 4056 28708
rect 3627 28328 3669 28337
rect 3627 28288 3628 28328
rect 3668 28288 3669 28328
rect 3627 28279 3669 28288
rect 3724 28328 3764 28337
rect 4108 28328 4148 30472
rect 4395 30428 4437 30437
rect 4395 30388 4396 30428
rect 4436 30388 4437 30428
rect 4395 30379 4437 30388
rect 4203 29588 4245 29597
rect 4203 29548 4204 29588
rect 4244 29548 4245 29588
rect 4203 29539 4245 29548
rect 4204 29000 4244 29539
rect 4204 28960 4340 29000
rect 3628 28194 3668 28279
rect 3340 27868 3476 27908
rect 3147 26900 3189 26909
rect 3147 26860 3148 26900
rect 3188 26860 3189 26900
rect 3147 26851 3189 26860
rect 2859 26816 2901 26825
rect 2859 26776 2860 26816
rect 2900 26776 2901 26816
rect 2859 26767 2901 26776
rect 2860 26682 2900 26767
rect 2859 26480 2901 26489
rect 2859 26440 2860 26480
rect 2900 26440 2901 26480
rect 2859 26431 2901 26440
rect 2860 26144 2900 26431
rect 3340 26237 3380 27868
rect 3435 27740 3477 27749
rect 3435 27700 3436 27740
rect 3476 27700 3477 27740
rect 3435 27691 3477 27700
rect 3436 26312 3476 27691
rect 3531 27656 3573 27665
rect 3531 27616 3532 27656
rect 3572 27616 3573 27656
rect 3531 27607 3573 27616
rect 3532 27522 3572 27607
rect 3724 27404 3764 28288
rect 3916 28288 4108 28328
rect 3916 27749 3956 28288
rect 4108 28279 4148 28288
rect 4204 28328 4244 28337
rect 4011 28160 4053 28169
rect 4011 28120 4012 28160
rect 4052 28120 4053 28160
rect 4011 28111 4053 28120
rect 3915 27740 3957 27749
rect 3915 27700 3916 27740
rect 3956 27700 3957 27740
rect 3915 27691 3957 27700
rect 4012 27651 4052 28111
rect 4204 27908 4244 28288
rect 4012 27602 4052 27611
rect 4108 27868 4244 27908
rect 3532 27364 3764 27404
rect 3532 26480 3572 27364
rect 3688 27236 4056 27245
rect 3728 27196 3770 27236
rect 3810 27196 3852 27236
rect 3892 27196 3934 27236
rect 3974 27196 4016 27236
rect 3688 27187 4056 27196
rect 4108 26984 4148 27868
rect 4204 27740 4244 27749
rect 4300 27740 4340 28960
rect 4244 27700 4340 27740
rect 4204 27691 4244 27700
rect 4012 26944 4148 26984
rect 3532 26440 3668 26480
rect 3436 26272 3572 26312
rect 3339 26228 3381 26237
rect 3339 26188 3340 26228
rect 3380 26188 3381 26228
rect 3339 26179 3381 26188
rect 3435 26144 3477 26153
rect 2860 25304 2900 26104
rect 3340 26125 3380 26134
rect 3435 26104 3436 26144
rect 3476 26104 3477 26144
rect 3435 26095 3477 26104
rect 3052 25892 3092 25901
rect 3052 25397 3092 25852
rect 3340 25565 3380 26085
rect 3436 26010 3476 26095
rect 3147 25556 3189 25565
rect 3147 25516 3148 25556
rect 3188 25516 3189 25556
rect 3147 25507 3189 25516
rect 3339 25556 3381 25565
rect 3339 25516 3340 25556
rect 3380 25516 3381 25556
rect 3339 25507 3381 25516
rect 3148 25422 3188 25507
rect 3051 25388 3093 25397
rect 3051 25348 3052 25388
rect 3092 25348 3093 25388
rect 3051 25339 3093 25348
rect 2956 25304 2996 25313
rect 2860 25264 2956 25304
rect 2956 25255 2996 25264
rect 2763 24800 2805 24809
rect 2763 24760 2764 24800
rect 2804 24760 2805 24800
rect 2763 24751 2805 24760
rect 3147 24800 3189 24809
rect 3147 24760 3148 24800
rect 3188 24760 3189 24800
rect 3147 24751 3189 24760
rect 3435 24800 3477 24809
rect 3435 24760 3436 24800
rect 3476 24760 3477 24800
rect 3435 24751 3477 24760
rect 3148 24666 3188 24751
rect 2476 24632 2516 24641
rect 2860 24632 2900 24641
rect 2379 23960 2421 23969
rect 2379 23920 2380 23960
rect 2420 23920 2421 23960
rect 2379 23911 2421 23920
rect 2476 23792 2516 24592
rect 2764 24592 2860 24632
rect 2667 24380 2709 24389
rect 2667 24340 2668 24380
rect 2708 24340 2709 24380
rect 2667 24331 2709 24340
rect 2668 24246 2708 24331
rect 2668 24044 2708 24053
rect 2764 24044 2804 24592
rect 2860 24583 2900 24592
rect 2955 24632 2997 24641
rect 2955 24592 2956 24632
rect 2996 24592 2997 24632
rect 2955 24583 2997 24592
rect 2956 24498 2996 24583
rect 2955 24380 2997 24389
rect 2955 24340 2956 24380
rect 2996 24340 2997 24380
rect 2955 24331 2997 24340
rect 2708 24004 2804 24044
rect 2668 23995 2708 24004
rect 2764 23801 2804 24004
rect 2956 23885 2996 24331
rect 3340 23885 3380 23932
rect 2955 23876 2997 23885
rect 2955 23836 2956 23876
rect 2996 23836 2997 23876
rect 2955 23827 2997 23836
rect 3339 23876 3381 23885
rect 3339 23827 3340 23876
rect 2188 23752 2420 23792
rect 2283 23624 2325 23633
rect 2283 23584 2284 23624
rect 2324 23584 2325 23624
rect 2283 23575 2325 23584
rect 2187 21692 2229 21701
rect 2187 21652 2188 21692
rect 2228 21652 2229 21692
rect 2187 21643 2229 21652
rect 2091 19592 2133 19601
rect 2091 19552 2092 19592
rect 2132 19552 2133 19592
rect 2091 19543 2133 19552
rect 2091 19256 2133 19265
rect 2091 19216 2092 19256
rect 2132 19216 2133 19256
rect 2091 19207 2133 19216
rect 2092 14141 2132 19207
rect 2188 18761 2228 21643
rect 2187 18752 2229 18761
rect 2187 18712 2188 18752
rect 2228 18712 2229 18752
rect 2187 18703 2229 18712
rect 2187 18584 2229 18593
rect 2187 18544 2188 18584
rect 2228 18544 2229 18584
rect 2187 18535 2229 18544
rect 2091 14132 2133 14141
rect 2091 14092 2092 14132
rect 2132 14092 2133 14132
rect 2091 14083 2133 14092
rect 2091 13880 2133 13889
rect 2091 13840 2092 13880
rect 2132 13840 2133 13880
rect 2091 13831 2133 13840
rect 2092 10193 2132 13831
rect 2188 11033 2228 18535
rect 2284 17585 2324 23575
rect 2283 17576 2325 17585
rect 2283 17536 2284 17576
rect 2324 17536 2325 17576
rect 2283 17527 2325 17536
rect 2284 17165 2324 17527
rect 2283 17156 2325 17165
rect 2283 17116 2284 17156
rect 2324 17116 2325 17156
rect 2283 17107 2325 17116
rect 2283 15392 2325 15401
rect 2283 15352 2284 15392
rect 2324 15352 2325 15392
rect 2283 15343 2325 15352
rect 2284 12788 2324 15343
rect 2380 15065 2420 23752
rect 2476 23549 2516 23752
rect 2763 23792 2805 23801
rect 2763 23752 2764 23792
rect 2804 23752 2805 23792
rect 2956 23792 2996 23827
rect 2763 23743 2805 23752
rect 2860 23771 2900 23780
rect 2956 23742 2996 23752
rect 3051 23792 3093 23801
rect 3051 23752 3052 23792
rect 3092 23752 3093 23792
rect 3380 23827 3381 23876
rect 3436 23834 3476 24751
rect 3532 24632 3572 26272
rect 3628 26237 3668 26440
rect 3627 26228 3669 26237
rect 3627 26188 3628 26228
rect 3668 26188 3669 26228
rect 3627 26179 3669 26188
rect 3820 26060 3860 26069
rect 3820 25901 3860 26020
rect 3915 26060 3957 26069
rect 3915 26020 3916 26060
rect 3956 26020 3957 26060
rect 3915 26011 3957 26020
rect 3916 25926 3956 26011
rect 3819 25892 3861 25901
rect 3819 25852 3820 25892
rect 3860 25852 3861 25892
rect 4012 25892 4052 26944
rect 4108 26816 4148 26825
rect 4108 26489 4148 26776
rect 4300 26648 4340 26657
rect 4107 26480 4149 26489
rect 4107 26440 4108 26480
rect 4148 26440 4149 26480
rect 4107 26431 4149 26440
rect 4300 26237 4340 26608
rect 4396 26312 4436 30379
rect 4492 26825 4532 26910
rect 4491 26816 4533 26825
rect 4491 26776 4492 26816
rect 4532 26776 4533 26816
rect 4491 26767 4533 26776
rect 4396 26272 4532 26312
rect 4299 26228 4341 26237
rect 4299 26188 4300 26228
rect 4340 26188 4341 26228
rect 4299 26179 4341 26188
rect 4396 26144 4436 26153
rect 4396 25901 4436 26104
rect 4395 25892 4437 25901
rect 4012 25852 4148 25892
rect 3819 25843 3861 25852
rect 3688 25724 4056 25733
rect 3728 25684 3770 25724
rect 3810 25684 3852 25724
rect 3892 25684 3934 25724
rect 3974 25684 4016 25724
rect 3688 25675 4056 25684
rect 3723 25388 3765 25397
rect 3723 25348 3724 25388
rect 3764 25348 3765 25388
rect 3723 25339 3765 25348
rect 3724 25304 3764 25339
rect 3724 25253 3764 25264
rect 3819 25304 3861 25313
rect 3819 25264 3820 25304
rect 3860 25264 3861 25304
rect 3819 25255 3861 25264
rect 3820 25170 3860 25255
rect 3628 24632 3668 24641
rect 3532 24592 3628 24632
rect 3532 23960 3572 24592
rect 3628 24583 3668 24592
rect 3688 24212 4056 24221
rect 3728 24172 3770 24212
rect 3810 24172 3852 24212
rect 3892 24172 3934 24212
rect 3974 24172 4016 24212
rect 3688 24163 4056 24172
rect 4108 24044 4148 25852
rect 4395 25852 4396 25892
rect 4436 25852 4437 25892
rect 4395 25843 4437 25852
rect 4203 25808 4245 25817
rect 4203 25768 4204 25808
rect 4244 25768 4245 25808
rect 4203 25759 4245 25768
rect 4204 25388 4244 25759
rect 4204 25339 4244 25348
rect 4300 25388 4340 25397
rect 4492 25388 4532 26272
rect 4340 25348 4532 25388
rect 3916 24004 4244 24044
rect 3532 23920 3764 23960
rect 3340 23788 3380 23797
rect 3436 23785 3476 23794
rect 3532 23792 3572 23801
rect 3051 23743 3093 23752
rect 2475 23540 2517 23549
rect 2475 23500 2476 23540
rect 2516 23500 2517 23540
rect 2475 23491 2517 23500
rect 2860 23372 2900 23731
rect 3052 23658 3092 23743
rect 3532 23633 3572 23752
rect 3147 23624 3189 23633
rect 3147 23584 3148 23624
rect 3188 23584 3189 23624
rect 3147 23575 3189 23584
rect 3531 23624 3573 23633
rect 3531 23584 3532 23624
rect 3572 23584 3573 23624
rect 3531 23575 3573 23584
rect 3628 23624 3668 23633
rect 3148 23490 3188 23575
rect 2572 23332 2900 23372
rect 3339 23372 3381 23381
rect 3339 23332 3340 23372
rect 3380 23332 3381 23372
rect 2475 19256 2517 19265
rect 2475 19216 2476 19256
rect 2516 19216 2517 19256
rect 2475 19207 2517 19216
rect 2476 19122 2516 19207
rect 2572 18593 2612 23332
rect 3339 23323 3381 23332
rect 2859 23204 2901 23213
rect 2859 23164 2860 23204
rect 2900 23164 2901 23204
rect 2859 23155 2901 23164
rect 3243 23204 3285 23213
rect 3243 23164 3244 23204
rect 3284 23164 3285 23204
rect 3243 23155 3285 23164
rect 2668 23120 2708 23129
rect 2668 22280 2708 23080
rect 2860 23070 2900 23155
rect 3244 23120 3284 23155
rect 3244 23069 3284 23080
rect 3340 23120 3380 23323
rect 3531 23204 3573 23213
rect 3531 23164 3532 23204
rect 3572 23164 3573 23204
rect 3531 23155 3573 23164
rect 3340 23071 3380 23080
rect 2763 22280 2805 22289
rect 3052 22280 3092 22289
rect 2708 22240 2764 22280
rect 2804 22240 2805 22280
rect 2668 22231 2708 22240
rect 2763 22231 2805 22240
rect 2956 22240 3052 22280
rect 2764 20768 2804 22231
rect 2859 22196 2901 22205
rect 2859 22156 2860 22196
rect 2900 22156 2901 22196
rect 2859 22147 2901 22156
rect 2860 22062 2900 22147
rect 2956 22121 2996 22240
rect 3052 22231 3092 22240
rect 2955 22112 2997 22121
rect 2955 22072 2956 22112
rect 2996 22072 2997 22112
rect 2955 22063 2997 22072
rect 3244 21608 3284 21617
rect 2956 21356 2996 21365
rect 2860 20768 2900 20777
rect 2764 20728 2860 20768
rect 2764 20096 2804 20728
rect 2860 20719 2900 20728
rect 2956 20180 2996 21316
rect 3052 20693 3092 20778
rect 3051 20684 3093 20693
rect 3051 20644 3052 20684
rect 3092 20644 3093 20684
rect 3051 20635 3093 20644
rect 3147 20684 3189 20693
rect 3147 20644 3148 20684
rect 3188 20644 3189 20684
rect 3147 20635 3189 20644
rect 2667 19508 2709 19517
rect 2667 19468 2668 19508
rect 2708 19468 2709 19508
rect 2667 19459 2709 19468
rect 2668 19374 2708 19459
rect 2764 19265 2804 20056
rect 2860 20140 2996 20180
rect 2763 19256 2805 19265
rect 2763 19216 2764 19256
rect 2804 19216 2805 19256
rect 2763 19207 2805 19216
rect 2476 18584 2516 18593
rect 2476 17240 2516 18544
rect 2571 18584 2613 18593
rect 2571 18544 2572 18584
rect 2612 18544 2613 18584
rect 2571 18535 2613 18544
rect 2572 18450 2612 18535
rect 2572 17744 2612 17753
rect 2572 17501 2612 17704
rect 2571 17492 2613 17501
rect 2571 17452 2572 17492
rect 2612 17452 2613 17492
rect 2571 17443 2613 17452
rect 2860 17417 2900 20140
rect 3148 20012 3188 20635
rect 3244 20348 3284 21568
rect 3340 21608 3380 21617
rect 3380 21568 3476 21608
rect 3340 21559 3380 21568
rect 3436 20684 3476 21568
rect 3436 20635 3476 20644
rect 3244 20308 3476 20348
rect 3244 20096 3284 20106
rect 3244 20021 3284 20056
rect 3339 20096 3381 20105
rect 3339 20056 3340 20096
rect 3380 20056 3381 20096
rect 3339 20047 3381 20056
rect 3243 20012 3285 20021
rect 3148 19972 3244 20012
rect 3284 19972 3285 20012
rect 3243 19963 3285 19972
rect 3340 19962 3380 20047
rect 2955 19928 2997 19937
rect 2955 19888 2956 19928
rect 2996 19888 2997 19928
rect 2955 19879 2997 19888
rect 2956 19794 2996 19879
rect 3243 19760 3285 19769
rect 3243 19720 3244 19760
rect 3284 19720 3285 19760
rect 3243 19711 3285 19720
rect 3244 18929 3284 19711
rect 3339 19592 3381 19601
rect 3339 19552 3340 19592
rect 3380 19552 3381 19592
rect 3339 19543 3381 19552
rect 3243 18920 3285 18929
rect 3243 18880 3244 18920
rect 3284 18880 3285 18920
rect 3243 18871 3285 18880
rect 3340 18836 3380 19543
rect 3436 19088 3476 20308
rect 3532 20273 3572 23155
rect 3628 22961 3668 23584
rect 3724 23213 3764 23920
rect 3820 23624 3860 23633
rect 3820 23465 3860 23584
rect 3819 23456 3861 23465
rect 3819 23416 3820 23456
rect 3860 23416 3861 23456
rect 3819 23407 3861 23416
rect 3723 23204 3765 23213
rect 3723 23164 3724 23204
rect 3764 23164 3765 23204
rect 3723 23155 3765 23164
rect 3820 23120 3860 23129
rect 3916 23120 3956 24004
rect 4011 23876 4053 23885
rect 4011 23836 4012 23876
rect 4052 23836 4053 23876
rect 4011 23827 4053 23836
rect 4012 23742 4052 23827
rect 4107 23624 4149 23633
rect 4107 23584 4108 23624
rect 4148 23584 4149 23624
rect 4107 23575 4149 23584
rect 3860 23080 3956 23120
rect 3820 23071 3860 23080
rect 3723 23036 3765 23045
rect 3723 22996 3724 23036
rect 3764 22996 3765 23036
rect 3723 22987 3765 22996
rect 3627 22952 3669 22961
rect 3627 22912 3628 22952
rect 3668 22912 3669 22952
rect 3627 22903 3669 22912
rect 3724 22902 3764 22987
rect 4108 22877 4148 23575
rect 4107 22868 4149 22877
rect 4107 22828 4108 22868
rect 4148 22828 4149 22868
rect 4107 22819 4149 22828
rect 3688 22700 4056 22709
rect 3728 22660 3770 22700
rect 3810 22660 3852 22700
rect 3892 22660 3934 22700
rect 3974 22660 4016 22700
rect 3688 22651 4056 22660
rect 3627 21608 3669 21617
rect 3627 21568 3628 21608
rect 3668 21568 3669 21608
rect 3627 21559 3669 21568
rect 4011 21608 4053 21617
rect 4011 21568 4012 21608
rect 4052 21568 4053 21608
rect 4011 21559 4053 21568
rect 3628 21474 3668 21559
rect 4012 21474 4052 21559
rect 3688 21188 4056 21197
rect 3728 21148 3770 21188
rect 3810 21148 3852 21188
rect 3892 21148 3934 21188
rect 3974 21148 4016 21188
rect 4108 21188 4148 22819
rect 4204 21272 4244 24004
rect 4300 23717 4340 25348
rect 4588 23960 4628 30640
rect 4684 29420 4724 30892
rect 4780 30689 4820 32059
rect 4972 32058 5012 32143
rect 5452 31352 5492 32899
rect 5548 32864 5588 33664
rect 5644 33452 5684 33461
rect 5644 33041 5684 33412
rect 5740 33116 5780 34327
rect 5836 33872 5876 34495
rect 6027 34376 6069 34385
rect 6027 34336 6028 34376
rect 6068 34336 6069 34376
rect 6027 34327 6069 34336
rect 6028 34242 6068 34327
rect 5932 34208 5972 34219
rect 5932 34133 5972 34168
rect 5931 34124 5973 34133
rect 5931 34084 5932 34124
rect 5972 34084 5973 34124
rect 5931 34075 5973 34084
rect 5931 33956 5973 33965
rect 5931 33916 5932 33956
rect 5972 33916 5973 33956
rect 5931 33907 5973 33916
rect 5836 33823 5876 33832
rect 5836 33116 5876 33125
rect 5740 33076 5836 33116
rect 5836 33067 5876 33076
rect 5643 33032 5685 33041
rect 5643 32992 5644 33032
rect 5684 32992 5685 33032
rect 5643 32983 5685 32992
rect 5643 32864 5685 32873
rect 5548 32824 5644 32864
rect 5684 32824 5685 32864
rect 5643 32815 5685 32824
rect 5547 31520 5589 31529
rect 5547 31480 5548 31520
rect 5588 31480 5589 31520
rect 5547 31471 5589 31480
rect 5356 31312 5492 31352
rect 4928 31016 5296 31025
rect 4968 30976 5010 31016
rect 5050 30976 5092 31016
rect 5132 30976 5174 31016
rect 5214 30976 5256 31016
rect 4928 30967 5296 30976
rect 4875 30848 4917 30857
rect 4875 30808 4876 30848
rect 4916 30808 4917 30848
rect 4875 30799 4917 30808
rect 4779 30680 4821 30689
rect 4779 30640 4780 30680
rect 4820 30640 4821 30680
rect 4779 30631 4821 30640
rect 4876 30680 4916 30799
rect 4876 30631 4916 30640
rect 4971 30680 5013 30689
rect 4971 30640 4972 30680
rect 5012 30640 5013 30680
rect 4971 30631 5013 30640
rect 4972 30437 5012 30631
rect 4971 30428 5013 30437
rect 4971 30388 4972 30428
rect 5012 30388 5013 30428
rect 4971 30379 5013 30388
rect 5164 29840 5204 29849
rect 5356 29840 5396 31312
rect 5451 31184 5493 31193
rect 5451 31144 5452 31184
rect 5492 31144 5493 31184
rect 5451 31135 5493 31144
rect 5452 30680 5492 31135
rect 5452 30631 5492 30640
rect 5204 29800 5492 29840
rect 5164 29791 5204 29800
rect 4928 29504 5296 29513
rect 4968 29464 5010 29504
rect 5050 29464 5092 29504
rect 5132 29464 5174 29504
rect 5214 29464 5256 29504
rect 4928 29455 5296 29464
rect 4779 29420 4821 29429
rect 4684 29380 4780 29420
rect 4820 29380 4821 29420
rect 4779 29371 4821 29380
rect 5355 29420 5397 29429
rect 5355 29380 5356 29420
rect 5396 29380 5397 29420
rect 5355 29371 5397 29380
rect 4683 28580 4725 28589
rect 4683 28540 4684 28580
rect 4724 28540 4725 28580
rect 4683 28531 4725 28540
rect 4684 28328 4724 28531
rect 4684 28279 4724 28288
rect 4780 27077 4820 29371
rect 5067 29252 5109 29261
rect 5356 29252 5396 29371
rect 5452 29252 5492 29800
rect 5067 29212 5068 29252
rect 5108 29212 5396 29252
rect 5439 29212 5492 29252
rect 5067 29203 5109 29212
rect 5068 29168 5108 29203
rect 5439 29168 5479 29212
rect 5068 29118 5108 29128
rect 5356 29128 5479 29168
rect 5260 28916 5300 28925
rect 5164 28876 5260 28916
rect 5164 28342 5204 28876
rect 5260 28867 5300 28876
rect 5356 28421 5396 29128
rect 5548 29093 5588 31471
rect 5644 31352 5684 32815
rect 5739 32696 5781 32705
rect 5739 32656 5740 32696
rect 5780 32656 5781 32696
rect 5739 32647 5781 32656
rect 5644 30521 5684 31312
rect 5643 30512 5685 30521
rect 5643 30472 5644 30512
rect 5684 30472 5685 30512
rect 5643 30463 5685 30472
rect 5643 30260 5685 30269
rect 5643 30220 5644 30260
rect 5684 30220 5685 30260
rect 5643 30211 5685 30220
rect 5547 29084 5589 29093
rect 5547 29044 5548 29084
rect 5588 29044 5589 29084
rect 5547 29035 5589 29044
rect 5451 29000 5493 29009
rect 5451 28960 5452 29000
rect 5492 28960 5493 29000
rect 5644 29000 5684 30211
rect 5740 30101 5780 32647
rect 5932 31361 5972 33907
rect 6028 33713 6068 33798
rect 6027 33704 6069 33713
rect 6027 33664 6028 33704
rect 6068 33664 6069 33704
rect 6027 33655 6069 33664
rect 6124 33536 6164 34504
rect 6028 33496 6164 33536
rect 6220 34376 6260 34385
rect 6028 32612 6068 33496
rect 6220 33293 6260 34336
rect 6219 33284 6261 33293
rect 6219 33244 6220 33284
rect 6260 33244 6261 33284
rect 6219 33235 6261 33244
rect 6124 32789 6164 32874
rect 6220 32864 6260 32873
rect 6123 32780 6165 32789
rect 6123 32740 6124 32780
rect 6164 32740 6165 32780
rect 6123 32731 6165 32740
rect 6028 32572 6164 32612
rect 6027 32024 6069 32033
rect 6027 31984 6028 32024
rect 6068 31984 6069 32024
rect 6027 31975 6069 31984
rect 6028 31529 6068 31975
rect 6027 31520 6069 31529
rect 6027 31480 6028 31520
rect 6068 31480 6069 31520
rect 6027 31471 6069 31480
rect 5931 31352 5973 31361
rect 5931 31312 5932 31352
rect 5972 31312 5973 31352
rect 5931 31303 5973 31312
rect 6028 31352 6068 31471
rect 6124 31361 6164 32572
rect 6220 32369 6260 32824
rect 6219 32360 6261 32369
rect 6219 32320 6220 32360
rect 6260 32320 6261 32360
rect 6219 32311 6261 32320
rect 6220 32192 6260 32201
rect 6028 31303 6068 31312
rect 6123 31352 6165 31361
rect 6123 31312 6124 31352
rect 6164 31312 6165 31352
rect 6123 31303 6165 31312
rect 5836 31184 5876 31193
rect 6027 31184 6069 31193
rect 5876 31144 5972 31184
rect 5836 31135 5876 31144
rect 5932 30675 5972 31144
rect 6027 31144 6028 31184
rect 6068 31144 6069 31184
rect 6027 31135 6069 31144
rect 5932 30626 5972 30635
rect 5739 30092 5781 30101
rect 5739 30052 5740 30092
rect 5780 30052 5781 30092
rect 5739 30043 5781 30052
rect 5644 28960 5876 29000
rect 5451 28951 5493 28960
rect 5355 28412 5397 28421
rect 5355 28372 5356 28412
rect 5396 28372 5397 28412
rect 5355 28363 5397 28372
rect 5164 28293 5204 28302
rect 5355 28244 5397 28253
rect 5355 28204 5356 28244
rect 5396 28204 5397 28244
rect 5355 28195 5397 28204
rect 5356 28110 5396 28195
rect 4928 27992 5296 28001
rect 4968 27952 5010 27992
rect 5050 27952 5092 27992
rect 5132 27952 5174 27992
rect 5214 27952 5256 27992
rect 4928 27943 5296 27952
rect 4779 27068 4821 27077
rect 4779 27028 4780 27068
rect 4820 27028 4821 27068
rect 4779 27019 4821 27028
rect 4780 26825 4820 27019
rect 4779 26816 4821 26825
rect 4779 26776 4780 26816
rect 4820 26776 4821 26816
rect 4779 26767 4821 26776
rect 4683 26480 4725 26489
rect 4683 26440 4684 26480
rect 4724 26440 4725 26480
rect 4683 26431 4725 26440
rect 4928 26480 5296 26489
rect 4968 26440 5010 26480
rect 5050 26440 5092 26480
rect 5132 26440 5174 26480
rect 5214 26440 5256 26480
rect 4928 26431 5296 26440
rect 4684 24627 4724 26431
rect 5452 26312 5492 28951
rect 5548 27656 5588 27665
rect 5548 27077 5588 27616
rect 5644 27656 5684 27665
rect 5547 27068 5589 27077
rect 5547 27028 5548 27068
rect 5588 27028 5589 27068
rect 5547 27019 5589 27028
rect 5452 26272 5588 26312
rect 4875 26228 4917 26237
rect 4875 26188 4876 26228
rect 4916 26188 4917 26228
rect 4875 26179 4917 26188
rect 5067 26228 5109 26237
rect 5067 26188 5068 26228
rect 5108 26188 5109 26228
rect 5067 26179 5109 26188
rect 4876 26139 4916 26179
rect 4876 26090 4916 26099
rect 5068 26094 5108 26179
rect 5452 26144 5492 26155
rect 5452 26069 5492 26104
rect 5451 26060 5493 26069
rect 5451 26020 5452 26060
rect 5492 26020 5493 26060
rect 5451 26011 5493 26020
rect 5451 25388 5493 25397
rect 5451 25348 5452 25388
rect 5492 25348 5493 25388
rect 5451 25339 5493 25348
rect 5308 25313 5348 25322
rect 4780 25304 4820 25313
rect 5348 25273 5396 25304
rect 5308 25264 5396 25273
rect 4780 24800 4820 25264
rect 4928 24968 5296 24977
rect 4968 24928 5010 24968
rect 5050 24928 5092 24968
rect 5132 24928 5174 24968
rect 5214 24928 5256 24968
rect 4928 24919 5296 24928
rect 5068 24800 5108 24809
rect 5356 24800 5396 25264
rect 5452 25220 5492 25339
rect 5452 25171 5492 25180
rect 5451 24884 5493 24893
rect 5548 24884 5588 26272
rect 5644 25313 5684 27616
rect 5739 26816 5781 26825
rect 5739 26776 5740 26816
rect 5780 26776 5781 26816
rect 5739 26767 5781 26776
rect 5740 26682 5780 26767
rect 5836 26657 5876 28960
rect 5931 28916 5973 28925
rect 5931 28876 5932 28916
rect 5972 28876 5973 28916
rect 5931 28867 5973 28876
rect 5932 28337 5972 28867
rect 5931 28328 5973 28337
rect 5931 28288 5932 28328
rect 5972 28288 5973 28328
rect 5931 28279 5973 28288
rect 5932 28194 5972 28279
rect 6028 27572 6068 31135
rect 6124 30764 6164 30773
rect 6124 29177 6164 30724
rect 6220 30269 6260 32152
rect 6316 31688 6356 35251
rect 6412 34805 6452 35428
rect 6411 34796 6453 34805
rect 6411 34756 6412 34796
rect 6452 34756 6453 34796
rect 6411 34747 6453 34756
rect 6411 34376 6453 34385
rect 6411 34336 6412 34376
rect 6452 34336 6453 34376
rect 6411 34327 6453 34336
rect 6412 32024 6452 34327
rect 6507 33368 6549 33377
rect 6507 33328 6508 33368
rect 6548 33328 6549 33368
rect 6507 33319 6549 33328
rect 6508 32864 6548 33319
rect 6508 32201 6548 32824
rect 6700 32360 6740 36016
rect 6796 33713 6836 37015
rect 6988 36737 7028 38872
rect 7084 38753 7124 39208
rect 7083 38744 7125 38753
rect 7083 38704 7084 38744
rect 7124 38704 7125 38744
rect 7083 38695 7125 38704
rect 7083 38156 7125 38165
rect 7083 38116 7084 38156
rect 7124 38116 7125 38156
rect 7083 38107 7125 38116
rect 7084 38022 7124 38107
rect 7083 37316 7125 37325
rect 7083 37276 7084 37316
rect 7124 37276 7125 37316
rect 7083 37267 7125 37276
rect 7084 37182 7124 37267
rect 7084 36896 7124 36905
rect 7180 36896 7220 42928
rect 7372 41777 7412 42928
rect 7371 41768 7413 41777
rect 7371 41728 7372 41768
rect 7412 41728 7413 41768
rect 7371 41719 7413 41728
rect 7564 41432 7604 42928
rect 7756 41693 7796 42928
rect 7755 41684 7797 41693
rect 7755 41644 7756 41684
rect 7796 41644 7797 41684
rect 7755 41635 7797 41644
rect 7564 41392 7796 41432
rect 7563 41264 7605 41273
rect 7563 41224 7564 41264
rect 7604 41224 7605 41264
rect 7563 41215 7605 41224
rect 7564 41130 7604 41215
rect 7275 40592 7317 40601
rect 7275 40552 7276 40592
rect 7316 40552 7317 40592
rect 7275 40543 7317 40552
rect 7276 38408 7316 40543
rect 7659 40424 7701 40433
rect 7659 40384 7660 40424
rect 7700 40384 7701 40424
rect 7659 40375 7701 40384
rect 7660 40097 7700 40375
rect 7756 40181 7796 41392
rect 7948 40769 7988 42928
rect 8043 41180 8085 41189
rect 8043 41140 8044 41180
rect 8084 41140 8085 41180
rect 8043 41131 8085 41140
rect 8044 41046 8084 41131
rect 8140 40844 8180 42928
rect 8236 41432 8276 41441
rect 8332 41432 8372 42928
rect 8276 41392 8372 41432
rect 8236 41383 8276 41392
rect 8044 40804 8180 40844
rect 7947 40760 7989 40769
rect 7947 40720 7948 40760
rect 7988 40720 7989 40760
rect 7947 40711 7989 40720
rect 7852 40256 7892 40265
rect 7755 40172 7797 40181
rect 7755 40132 7756 40172
rect 7796 40132 7797 40172
rect 7755 40123 7797 40132
rect 7659 40088 7701 40097
rect 7659 40048 7660 40088
rect 7700 40048 7701 40088
rect 7659 40039 7701 40048
rect 7371 39500 7413 39509
rect 7371 39460 7372 39500
rect 7412 39460 7413 39500
rect 7371 39451 7413 39460
rect 7372 38926 7412 39451
rect 7372 38877 7412 38886
rect 7755 38912 7797 38921
rect 7755 38872 7756 38912
rect 7796 38872 7797 38912
rect 7755 38863 7797 38872
rect 7852 38912 7892 40216
rect 8044 39425 8084 40804
rect 8524 40601 8564 42928
rect 8716 41516 8756 42928
rect 8620 41476 8756 41516
rect 8523 40592 8565 40601
rect 8523 40552 8524 40592
rect 8564 40552 8565 40592
rect 8523 40543 8565 40552
rect 8140 40424 8180 40433
rect 8180 40384 8564 40424
rect 8140 40375 8180 40384
rect 8235 40088 8277 40097
rect 8235 40048 8236 40088
rect 8276 40048 8277 40088
rect 8235 40039 8277 40048
rect 8236 39752 8276 40039
rect 8236 39703 8276 39712
rect 8427 39500 8469 39509
rect 8427 39460 8428 39500
rect 8468 39460 8469 39500
rect 8427 39451 8469 39460
rect 8043 39416 8085 39425
rect 8043 39376 8044 39416
rect 8084 39376 8085 39416
rect 8043 39367 8085 39376
rect 8428 39366 8468 39451
rect 8139 39080 8181 39089
rect 8139 39040 8140 39080
rect 8180 39040 8181 39080
rect 8139 39031 8181 39040
rect 8331 39080 8373 39089
rect 8331 39040 8332 39080
rect 8372 39040 8373 39080
rect 8331 39031 8373 39040
rect 7852 38863 7892 38872
rect 7947 38912 7989 38921
rect 7947 38872 7948 38912
rect 7988 38872 7989 38912
rect 7947 38863 7989 38872
rect 7276 38359 7316 38368
rect 7564 38744 7604 38753
rect 7275 38240 7317 38249
rect 7275 38200 7276 38240
rect 7316 38200 7317 38240
rect 7275 38191 7317 38200
rect 7276 37400 7316 38191
rect 7468 38156 7508 38165
rect 7468 37820 7508 38116
rect 7372 37780 7508 37820
rect 7372 37568 7412 37780
rect 7372 37519 7412 37528
rect 7276 37360 7412 37400
rect 7275 37232 7317 37241
rect 7275 37192 7276 37232
rect 7316 37192 7317 37232
rect 7275 37183 7317 37192
rect 7276 37098 7316 37183
rect 7372 36905 7412 37360
rect 7124 36856 7220 36896
rect 7371 36896 7413 36905
rect 7371 36856 7372 36896
rect 7412 36856 7413 36896
rect 7084 36847 7124 36856
rect 7371 36847 7413 36856
rect 7275 36812 7317 36821
rect 7180 36772 7276 36812
rect 7316 36772 7317 36812
rect 6987 36728 7029 36737
rect 6987 36688 6988 36728
rect 7028 36688 7029 36728
rect 6987 36679 7029 36688
rect 6892 36644 6932 36655
rect 6892 36569 6932 36604
rect 6891 36560 6933 36569
rect 6891 36520 6892 36560
rect 6932 36520 6933 36560
rect 6891 36511 6933 36520
rect 6988 35972 7028 36679
rect 6988 35923 7028 35932
rect 7084 35972 7124 35981
rect 7180 35972 7220 36772
rect 7275 36763 7317 36772
rect 7468 36728 7508 36737
rect 7275 36560 7317 36569
rect 7275 36520 7276 36560
rect 7316 36520 7317 36560
rect 7275 36511 7317 36520
rect 7124 35932 7220 35972
rect 6891 34124 6933 34133
rect 6891 34084 6892 34124
rect 6932 34084 6933 34124
rect 6891 34075 6933 34084
rect 6795 33704 6837 33713
rect 6795 33664 6796 33704
rect 6836 33664 6837 33704
rect 6795 33655 6837 33664
rect 6892 32957 6932 34075
rect 7084 33284 7124 35932
rect 7276 35813 7316 36511
rect 7275 35804 7317 35813
rect 7275 35764 7276 35804
rect 7316 35764 7317 35804
rect 7275 35755 7317 35764
rect 7276 35057 7316 35755
rect 7468 35477 7508 36688
rect 7564 36065 7604 38704
rect 7660 37400 7700 37411
rect 7660 37325 7700 37360
rect 7756 37400 7796 38863
rect 7948 38778 7988 38863
rect 7851 38576 7893 38585
rect 7851 38536 7852 38576
rect 7892 38536 7893 38576
rect 7851 38527 7893 38536
rect 7852 38240 7892 38527
rect 7852 38191 7892 38200
rect 8043 37652 8085 37661
rect 8043 37612 8044 37652
rect 8084 37612 8085 37652
rect 8043 37603 8085 37612
rect 7659 37316 7701 37325
rect 7659 37276 7660 37316
rect 7700 37276 7701 37316
rect 7659 37267 7701 37276
rect 7563 36056 7605 36065
rect 7563 36016 7564 36056
rect 7604 36016 7605 36056
rect 7563 36007 7605 36016
rect 7564 35888 7604 35897
rect 7564 35561 7604 35848
rect 7659 35720 7701 35729
rect 7659 35680 7660 35720
rect 7700 35680 7701 35720
rect 7659 35671 7701 35680
rect 7563 35552 7605 35561
rect 7563 35512 7564 35552
rect 7604 35512 7605 35552
rect 7563 35503 7605 35512
rect 7467 35468 7509 35477
rect 7467 35428 7468 35468
rect 7508 35428 7509 35468
rect 7467 35419 7509 35428
rect 7564 35384 7604 35393
rect 7660 35384 7700 35671
rect 7604 35344 7700 35384
rect 7756 35384 7796 37360
rect 7947 37400 7989 37409
rect 7947 37360 7948 37400
rect 7988 37360 7989 37400
rect 7947 37351 7989 37360
rect 7851 37316 7893 37325
rect 7851 37276 7852 37316
rect 7892 37276 7893 37316
rect 7851 37267 7893 37276
rect 7852 35645 7892 37267
rect 7948 35897 7988 37351
rect 8044 37232 8084 37603
rect 8140 37409 8180 39031
rect 8332 38996 8372 39031
rect 8332 38945 8372 38956
rect 8427 38912 8469 38921
rect 8427 38872 8428 38912
rect 8468 38872 8469 38912
rect 8427 38863 8469 38872
rect 8331 38492 8373 38501
rect 8331 38452 8332 38492
rect 8372 38452 8373 38492
rect 8331 38443 8373 38452
rect 8332 37661 8372 38443
rect 8331 37652 8373 37661
rect 8331 37612 8332 37652
rect 8372 37612 8373 37652
rect 8331 37603 8373 37612
rect 8428 37484 8468 38863
rect 8524 37829 8564 40384
rect 8620 40097 8660 41476
rect 8716 41264 8756 41273
rect 8716 40685 8756 41224
rect 8715 40676 8757 40685
rect 8715 40636 8716 40676
rect 8756 40636 8757 40676
rect 8715 40627 8757 40636
rect 8619 40088 8661 40097
rect 8619 40048 8620 40088
rect 8660 40048 8661 40088
rect 8619 40039 8661 40048
rect 8620 39752 8660 39761
rect 8620 38417 8660 39712
rect 8908 39668 8948 42928
rect 8812 39628 8948 39668
rect 8619 38408 8661 38417
rect 8619 38368 8620 38408
rect 8660 38368 8661 38408
rect 8619 38359 8661 38368
rect 8523 37820 8565 37829
rect 8523 37780 8524 37820
rect 8564 37780 8565 37820
rect 8620 37820 8660 38359
rect 8812 38081 8852 39628
rect 8907 38996 8949 39005
rect 8907 38956 8908 38996
rect 8948 38956 8949 38996
rect 8907 38947 8949 38956
rect 8908 38912 8948 38947
rect 9100 38921 9140 42928
rect 9195 40256 9237 40265
rect 9195 40216 9196 40256
rect 9236 40216 9237 40256
rect 9195 40207 9237 40216
rect 8811 38072 8853 38081
rect 8811 38032 8812 38072
rect 8852 38032 8853 38072
rect 8811 38023 8853 38032
rect 8908 37820 8948 38872
rect 9099 38912 9141 38921
rect 9099 38872 9100 38912
rect 9140 38872 9141 38912
rect 9099 38863 9141 38872
rect 8620 37780 8755 37820
rect 8523 37771 8565 37780
rect 8715 37652 8755 37780
rect 8236 37444 8468 37484
rect 8524 37612 8755 37652
rect 8812 37780 8948 37820
rect 9100 38240 9140 38249
rect 8139 37400 8181 37409
rect 8139 37360 8140 37400
rect 8180 37360 8181 37400
rect 8139 37351 8181 37360
rect 8236 37400 8276 37444
rect 8044 37192 8180 37232
rect 7947 35888 7989 35897
rect 7947 35848 7948 35888
rect 7988 35848 7989 35888
rect 7947 35839 7989 35848
rect 8044 35893 8084 35902
rect 8044 35729 8084 35853
rect 8043 35720 8085 35729
rect 8043 35680 8044 35720
rect 8084 35680 8085 35720
rect 8043 35671 8085 35680
rect 7851 35636 7893 35645
rect 7851 35596 7852 35636
rect 7892 35596 7893 35636
rect 7851 35587 7893 35596
rect 7756 35344 8084 35384
rect 7564 35335 7604 35344
rect 7371 35216 7413 35225
rect 7371 35176 7372 35216
rect 7412 35176 7413 35216
rect 7371 35167 7413 35176
rect 7756 35216 7796 35225
rect 7372 35082 7412 35167
rect 7275 35048 7317 35057
rect 7275 35008 7276 35048
rect 7316 35008 7317 35048
rect 7275 34999 7317 35008
rect 7467 35048 7509 35057
rect 7467 35008 7468 35048
rect 7508 35008 7509 35048
rect 7467 34999 7509 35008
rect 7275 34796 7317 34805
rect 7275 34756 7276 34796
rect 7316 34756 7317 34796
rect 7275 34747 7317 34756
rect 7276 33704 7316 34747
rect 7468 34376 7508 34999
rect 7756 34973 7796 35176
rect 7755 34964 7797 34973
rect 7755 34924 7756 34964
rect 7796 34924 7797 34964
rect 7755 34915 7797 34924
rect 7756 34637 7796 34915
rect 7755 34628 7797 34637
rect 7755 34588 7756 34628
rect 7796 34588 7797 34628
rect 7755 34579 7797 34588
rect 8044 34385 8084 35344
rect 7468 34327 7508 34336
rect 7948 34376 7988 34385
rect 7660 34292 7700 34301
rect 7948 34292 7988 34336
rect 8043 34376 8085 34385
rect 8043 34336 8044 34376
rect 8084 34336 8085 34376
rect 8043 34327 8085 34336
rect 7700 34252 7988 34292
rect 7660 34243 7700 34252
rect 8044 34242 8084 34327
rect 7563 34208 7605 34217
rect 7563 34168 7564 34208
rect 7604 34168 7605 34208
rect 7563 34159 7605 34168
rect 7276 33293 7316 33664
rect 7468 33704 7508 33713
rect 6988 33244 7124 33284
rect 7275 33284 7317 33293
rect 7275 33244 7276 33284
rect 7316 33244 7317 33284
rect 6891 32948 6933 32957
rect 6891 32908 6892 32948
rect 6932 32908 6933 32948
rect 6891 32899 6933 32908
rect 6796 32864 6836 32873
rect 6796 32537 6836 32824
rect 6892 32864 6932 32899
rect 6892 32814 6932 32824
rect 6988 32612 7028 33244
rect 7275 33235 7317 33244
rect 7084 33116 7124 33125
rect 7468 33116 7508 33664
rect 7564 33620 7604 34159
rect 8140 34124 8180 37192
rect 8236 36821 8276 37360
rect 8524 36980 8564 37612
rect 8716 37400 8756 37409
rect 8812 37400 8852 37780
rect 9100 37736 9140 38200
rect 8756 37360 8852 37400
rect 8908 37696 9140 37736
rect 8619 37316 8661 37325
rect 8619 37276 8620 37316
rect 8660 37276 8661 37316
rect 8619 37267 8661 37276
rect 8428 36940 8564 36980
rect 8235 36812 8277 36821
rect 8235 36772 8236 36812
rect 8276 36772 8277 36812
rect 8235 36763 8277 36772
rect 8235 35804 8277 35813
rect 8235 35764 8236 35804
rect 8276 35764 8277 35804
rect 8235 35755 8277 35764
rect 8236 35670 8276 35755
rect 8235 35552 8277 35561
rect 8235 35512 8236 35552
rect 8276 35512 8277 35552
rect 8235 35503 8277 35512
rect 7564 33571 7604 33580
rect 7660 34084 8180 34124
rect 7660 33536 7700 34084
rect 8236 33872 8276 35503
rect 8428 34628 8468 36940
rect 8620 36905 8660 37267
rect 8619 36896 8661 36905
rect 8619 36856 8620 36896
rect 8660 36856 8661 36896
rect 8716 36896 8756 37360
rect 8908 37073 8948 37696
rect 9196 37568 9236 40207
rect 9292 38333 9332 42928
rect 9387 41264 9429 41273
rect 9387 41224 9388 41264
rect 9428 41224 9429 41264
rect 9387 41215 9429 41224
rect 9388 40424 9428 41215
rect 9388 40375 9428 40384
rect 9387 39500 9429 39509
rect 9387 39460 9388 39500
rect 9428 39460 9429 39500
rect 9387 39451 9429 39460
rect 9388 38926 9428 39451
rect 9388 38877 9428 38886
rect 9387 38744 9429 38753
rect 9387 38704 9388 38744
rect 9428 38704 9429 38744
rect 9387 38695 9429 38704
rect 9291 38324 9333 38333
rect 9291 38284 9292 38324
rect 9332 38284 9333 38324
rect 9291 38275 9333 38284
rect 9388 38081 9428 38695
rect 9387 38072 9429 38081
rect 9387 38032 9388 38072
rect 9428 38032 9429 38072
rect 9387 38023 9429 38032
rect 9004 37528 9236 37568
rect 9292 37988 9332 37997
rect 8907 37064 8949 37073
rect 8907 37024 8908 37064
rect 8948 37024 8949 37064
rect 8907 37015 8949 37024
rect 8716 36856 8852 36896
rect 8619 36847 8661 36856
rect 8523 36812 8565 36821
rect 8523 36772 8524 36812
rect 8564 36772 8565 36812
rect 8523 36763 8565 36772
rect 8140 33832 8276 33872
rect 8332 34588 8468 34628
rect 7852 33704 7892 33713
rect 7892 33664 7988 33704
rect 7852 33655 7892 33664
rect 7755 33620 7797 33629
rect 7755 33580 7756 33620
rect 7796 33580 7797 33620
rect 7755 33571 7797 33580
rect 7660 33487 7700 33496
rect 7756 33486 7796 33571
rect 7124 33076 7508 33116
rect 7084 33067 7124 33076
rect 7755 33032 7797 33041
rect 7755 32992 7756 33032
rect 7796 32992 7797 33032
rect 7755 32983 7797 32992
rect 7275 32948 7317 32957
rect 7275 32908 7276 32948
rect 7316 32908 7317 32948
rect 7275 32899 7317 32908
rect 7083 32864 7125 32873
rect 7083 32824 7084 32864
rect 7124 32824 7125 32864
rect 7083 32815 7125 32824
rect 7276 32864 7316 32899
rect 7084 32730 7124 32815
rect 7276 32813 7316 32824
rect 7468 32864 7508 32873
rect 7371 32780 7413 32789
rect 7371 32740 7372 32780
rect 7412 32740 7413 32780
rect 7371 32731 7413 32740
rect 7372 32646 7412 32731
rect 6988 32572 7124 32612
rect 6795 32528 6837 32537
rect 6795 32488 6796 32528
rect 6836 32488 6837 32528
rect 6795 32479 6837 32488
rect 6604 32320 6740 32360
rect 6507 32192 6549 32201
rect 6507 32152 6508 32192
rect 6548 32152 6549 32192
rect 6507 32143 6549 32152
rect 6412 31984 6548 32024
rect 6316 31648 6452 31688
rect 6315 31268 6357 31277
rect 6315 31228 6316 31268
rect 6356 31228 6357 31268
rect 6315 31219 6357 31228
rect 6316 30941 6356 31219
rect 6315 30932 6357 30941
rect 6315 30892 6316 30932
rect 6356 30892 6357 30932
rect 6315 30883 6357 30892
rect 6316 30680 6356 30883
rect 6316 30631 6356 30640
rect 6412 30680 6452 31648
rect 6412 30512 6452 30640
rect 6508 30680 6548 31984
rect 6604 31613 6644 32320
rect 6891 32276 6933 32285
rect 6891 32236 6892 32276
rect 6932 32236 6933 32276
rect 6891 32227 6933 32236
rect 6699 32192 6741 32201
rect 6699 32152 6700 32192
rect 6740 32152 6741 32192
rect 6699 32143 6741 32152
rect 6796 32192 6836 32201
rect 6603 31604 6645 31613
rect 6603 31564 6604 31604
rect 6644 31564 6645 31604
rect 6603 31555 6645 31564
rect 6603 31436 6645 31445
rect 6603 31396 6604 31436
rect 6644 31396 6645 31436
rect 6603 31387 6645 31396
rect 6604 30848 6644 31387
rect 6604 30799 6644 30808
rect 6700 30680 6740 32143
rect 6796 30857 6836 32152
rect 6892 32142 6932 32227
rect 7084 32201 7124 32572
rect 7179 32528 7221 32537
rect 7179 32488 7180 32528
rect 7220 32488 7221 32528
rect 7179 32479 7221 32488
rect 7083 32192 7125 32201
rect 7083 32152 7084 32192
rect 7124 32152 7125 32192
rect 7083 32143 7125 32152
rect 7180 32024 7220 32479
rect 7180 31975 7220 31984
rect 6891 31520 6933 31529
rect 6891 31480 6892 31520
rect 6932 31480 6933 31520
rect 6891 31471 6933 31480
rect 7083 31520 7125 31529
rect 7083 31480 7084 31520
rect 7124 31480 7125 31520
rect 7083 31471 7125 31480
rect 6892 31109 6932 31471
rect 6891 31100 6933 31109
rect 6891 31060 6892 31100
rect 6932 31060 6933 31100
rect 6891 31051 6933 31060
rect 6795 30848 6837 30857
rect 6795 30808 6796 30848
rect 6836 30808 6837 30848
rect 6795 30799 6837 30808
rect 7084 30848 7124 31471
rect 7468 31366 7508 32824
rect 7564 32864 7604 32873
rect 7564 32360 7604 32824
rect 7756 32864 7796 32983
rect 7756 32815 7796 32824
rect 7851 32864 7893 32873
rect 7851 32824 7852 32864
rect 7892 32824 7893 32864
rect 7851 32815 7893 32824
rect 7852 32730 7892 32815
rect 7852 32360 7892 32369
rect 7948 32360 7988 33664
rect 8043 33032 8085 33041
rect 8043 32992 8044 33032
rect 8084 32992 8085 33032
rect 8043 32983 8085 32992
rect 7564 32320 7796 32360
rect 7660 32192 7700 32201
rect 7564 32152 7660 32192
rect 7564 31529 7604 32152
rect 7660 32143 7700 32152
rect 7660 32024 7700 32033
rect 7563 31520 7605 31529
rect 7563 31480 7564 31520
rect 7604 31480 7605 31520
rect 7563 31471 7605 31480
rect 7660 31445 7700 31984
rect 7756 31529 7796 32320
rect 7892 32320 7988 32360
rect 8044 32864 8084 32983
rect 7852 32311 7892 32320
rect 8044 32276 8084 32824
rect 8140 32369 8180 33832
rect 8332 33788 8372 34588
rect 8427 34460 8469 34469
rect 8427 34420 8428 34460
rect 8468 34420 8469 34460
rect 8427 34411 8469 34420
rect 8428 34326 8468 34411
rect 8524 34376 8564 36763
rect 8332 33748 8468 33788
rect 8235 33704 8277 33713
rect 8235 33664 8236 33704
rect 8276 33664 8277 33704
rect 8235 33655 8277 33664
rect 8236 33570 8276 33655
rect 8331 33620 8373 33629
rect 8331 33580 8332 33620
rect 8372 33580 8373 33620
rect 8331 33571 8373 33580
rect 8235 32780 8277 32789
rect 8235 32740 8236 32780
rect 8276 32740 8277 32780
rect 8235 32731 8277 32740
rect 8139 32360 8181 32369
rect 8139 32320 8140 32360
rect 8180 32320 8181 32360
rect 8139 32311 8181 32320
rect 7948 32236 8084 32276
rect 7948 31697 7988 32236
rect 8139 32192 8181 32201
rect 8044 32147 8084 32156
rect 8139 32152 8140 32192
rect 8180 32152 8181 32192
rect 8139 32143 8181 32152
rect 8236 32192 8276 32731
rect 8332 32360 8372 33571
rect 8428 32369 8468 33748
rect 8332 32311 8372 32320
rect 8427 32360 8469 32369
rect 8427 32320 8428 32360
rect 8468 32320 8469 32360
rect 8427 32311 8469 32320
rect 8236 32143 8276 32152
rect 7947 31688 7989 31697
rect 7947 31648 7948 31688
rect 7988 31648 7989 31688
rect 7947 31639 7989 31648
rect 8044 31529 8084 32107
rect 8140 31604 8180 32143
rect 8140 31564 8468 31604
rect 7755 31520 7797 31529
rect 7755 31480 7756 31520
rect 7796 31480 7797 31520
rect 7755 31471 7797 31480
rect 8043 31520 8085 31529
rect 8043 31480 8044 31520
rect 8084 31480 8085 31520
rect 8043 31471 8085 31480
rect 7659 31436 7701 31445
rect 7659 31396 7660 31436
rect 7700 31396 7701 31436
rect 7659 31387 7701 31396
rect 8235 31436 8277 31445
rect 8235 31396 8236 31436
rect 8276 31396 8277 31436
rect 8235 31387 8277 31396
rect 7276 31352 7316 31361
rect 7179 31184 7221 31193
rect 7179 31144 7180 31184
rect 7220 31144 7221 31184
rect 7179 31135 7221 31144
rect 7084 30799 7124 30808
rect 6988 30680 7028 30689
rect 6700 30640 6988 30680
rect 6508 30631 6548 30640
rect 6988 30631 7028 30640
rect 7180 30680 7220 31135
rect 7180 30631 7220 30640
rect 6412 30472 6548 30512
rect 6219 30260 6261 30269
rect 6219 30220 6220 30260
rect 6260 30220 6261 30260
rect 6219 30211 6261 30220
rect 6219 30092 6261 30101
rect 6219 30052 6220 30092
rect 6260 30052 6261 30092
rect 6219 30043 6261 30052
rect 6123 29168 6165 29177
rect 6123 29128 6124 29168
rect 6164 29128 6165 29168
rect 6123 29119 6165 29128
rect 6220 27833 6260 30043
rect 6315 30008 6357 30017
rect 6315 29968 6316 30008
rect 6356 29968 6357 30008
rect 6315 29959 6357 29968
rect 6316 29765 6356 29959
rect 6411 29840 6453 29849
rect 6411 29800 6412 29840
rect 6452 29800 6453 29840
rect 6411 29791 6453 29800
rect 6315 29756 6357 29765
rect 6315 29716 6316 29756
rect 6356 29716 6357 29756
rect 6315 29707 6357 29716
rect 6219 27824 6261 27833
rect 6219 27784 6220 27824
rect 6260 27784 6261 27824
rect 6219 27775 6261 27784
rect 5931 27068 5973 27077
rect 5931 27028 5932 27068
rect 5972 27028 5973 27068
rect 5931 27019 5973 27028
rect 5932 26934 5972 27019
rect 5931 26732 5973 26741
rect 5931 26692 5932 26732
rect 5972 26692 5973 26732
rect 5931 26683 5973 26692
rect 5835 26648 5877 26657
rect 5835 26608 5836 26648
rect 5876 26608 5877 26648
rect 5835 26599 5877 26608
rect 5643 25304 5685 25313
rect 5643 25264 5644 25304
rect 5684 25264 5685 25304
rect 5643 25255 5685 25264
rect 5451 24844 5452 24884
rect 5492 24844 5588 24884
rect 5451 24835 5493 24844
rect 4780 24760 5012 24800
rect 4876 24632 4916 24641
rect 4684 24592 4876 24627
rect 4684 24587 4916 24592
rect 4876 24053 4916 24587
rect 4875 24044 4917 24053
rect 4875 24004 4876 24044
rect 4916 24004 4917 24044
rect 4875 23995 4917 24004
rect 4396 23920 4628 23960
rect 4299 23708 4341 23717
rect 4299 23668 4300 23708
rect 4340 23668 4341 23708
rect 4299 23659 4341 23668
rect 4396 23381 4436 23920
rect 4491 23792 4533 23801
rect 4491 23752 4492 23792
rect 4532 23752 4533 23792
rect 4491 23743 4533 23752
rect 4588 23792 4628 23801
rect 4395 23372 4437 23381
rect 4395 23332 4396 23372
rect 4436 23332 4437 23372
rect 4395 23323 4437 23332
rect 4492 23297 4532 23743
rect 4588 23633 4628 23752
rect 4684 23792 4724 23801
rect 4587 23624 4629 23633
rect 4587 23584 4588 23624
rect 4628 23584 4629 23624
rect 4587 23575 4629 23584
rect 4491 23288 4533 23297
rect 4491 23248 4492 23288
rect 4532 23248 4533 23288
rect 4491 23239 4533 23248
rect 4300 23120 4340 23129
rect 4684 23120 4724 23752
rect 4972 23633 5012 24760
rect 5108 24760 5396 24800
rect 5068 24751 5108 24760
rect 5260 24632 5300 24641
rect 5452 24632 5492 24835
rect 5300 24592 5492 24632
rect 5260 24583 5300 24592
rect 5739 24044 5781 24053
rect 5739 24004 5740 24044
rect 5780 24004 5781 24044
rect 5739 23995 5781 24004
rect 5068 23792 5108 23803
rect 5068 23717 5108 23752
rect 5163 23792 5205 23801
rect 5163 23752 5164 23792
rect 5204 23752 5205 23792
rect 5163 23743 5205 23752
rect 5356 23792 5396 23801
rect 5643 23792 5685 23801
rect 5396 23752 5492 23792
rect 5356 23743 5396 23752
rect 5067 23708 5109 23717
rect 5067 23668 5068 23708
rect 5108 23668 5109 23708
rect 5067 23659 5109 23668
rect 5164 23658 5204 23743
rect 5452 23633 5492 23752
rect 5643 23752 5644 23792
rect 5684 23752 5685 23792
rect 5643 23743 5685 23752
rect 5644 23658 5684 23743
rect 4876 23624 4916 23633
rect 4780 23584 4876 23624
rect 4780 23297 4820 23584
rect 4876 23575 4916 23584
rect 4971 23624 5013 23633
rect 4971 23584 4972 23624
rect 5012 23584 5013 23624
rect 4971 23575 5013 23584
rect 5260 23624 5300 23633
rect 5451 23624 5493 23633
rect 5300 23584 5396 23624
rect 5260 23575 5300 23584
rect 4928 23456 5296 23465
rect 4968 23416 5010 23456
rect 5050 23416 5092 23456
rect 5132 23416 5174 23456
rect 5214 23416 5256 23456
rect 4928 23407 5296 23416
rect 4779 23288 4821 23297
rect 5356 23288 5396 23584
rect 5451 23584 5452 23624
rect 5492 23584 5493 23624
rect 5451 23575 5493 23584
rect 5643 23456 5685 23465
rect 5643 23416 5644 23456
rect 5684 23416 5685 23456
rect 5643 23407 5685 23416
rect 4779 23248 4780 23288
rect 4820 23248 4821 23288
rect 4779 23239 4821 23248
rect 5260 23248 5396 23288
rect 5644 23288 5684 23407
rect 5644 23248 5689 23288
rect 4972 23204 5012 23213
rect 5012 23164 5108 23204
rect 4972 23155 5012 23164
rect 4340 23080 4628 23120
rect 4684 23106 4820 23120
rect 4684 23080 4780 23106
rect 4300 23071 4340 23080
rect 4491 22952 4533 22961
rect 4491 22912 4492 22952
rect 4532 22912 4533 22952
rect 4491 22903 4533 22912
rect 4492 22532 4532 22903
rect 4492 22483 4532 22492
rect 4299 22280 4341 22289
rect 4299 22240 4300 22280
rect 4340 22240 4341 22280
rect 4299 22231 4341 22240
rect 4300 22146 4340 22231
rect 4588 21356 4628 23080
rect 4780 22961 4820 23066
rect 4779 22952 4821 22961
rect 4779 22912 4780 22952
rect 4820 22912 4821 22952
rect 4779 22903 4821 22912
rect 4684 22448 4724 22457
rect 4684 21533 4724 22408
rect 4971 22280 5013 22289
rect 4971 22240 4972 22280
rect 5012 22240 5013 22280
rect 4971 22231 5013 22240
rect 5068 22280 5108 23164
rect 5164 23120 5204 23129
rect 5164 22961 5204 23080
rect 5260 23120 5300 23248
rect 5649 23204 5689 23248
rect 5644 23164 5689 23204
rect 5260 23071 5300 23080
rect 5355 23120 5397 23129
rect 5355 23080 5356 23120
rect 5396 23080 5397 23120
rect 5355 23071 5397 23080
rect 5452 23120 5492 23129
rect 5356 22986 5396 23071
rect 5163 22952 5205 22961
rect 5163 22912 5164 22952
rect 5204 22912 5205 22952
rect 5163 22903 5205 22912
rect 5068 22231 5108 22240
rect 5356 22280 5396 22291
rect 5452 22289 5492 23080
rect 5644 23120 5684 23164
rect 5644 23071 5684 23080
rect 5547 22952 5589 22961
rect 5547 22912 5548 22952
rect 5588 22912 5589 22952
rect 5547 22903 5589 22912
rect 4972 22146 5012 22231
rect 5356 22205 5396 22240
rect 5451 22280 5493 22289
rect 5451 22240 5452 22280
rect 5492 22240 5493 22280
rect 5451 22231 5493 22240
rect 5355 22196 5397 22205
rect 5355 22156 5356 22196
rect 5396 22156 5397 22196
rect 5355 22147 5397 22156
rect 4928 21944 5296 21953
rect 4968 21904 5010 21944
rect 5050 21904 5092 21944
rect 5132 21904 5174 21944
rect 5214 21904 5256 21944
rect 4928 21895 5296 21904
rect 5259 21776 5301 21785
rect 5259 21736 5260 21776
rect 5300 21736 5301 21776
rect 5259 21727 5301 21736
rect 5260 21608 5300 21727
rect 5260 21559 5300 21568
rect 4683 21524 4725 21533
rect 4683 21484 4684 21524
rect 4724 21484 4725 21524
rect 4683 21475 4725 21484
rect 5451 21356 5493 21365
rect 4588 21316 4724 21356
rect 4204 21232 4628 21272
rect 4108 21148 4244 21188
rect 3688 21139 4056 21148
rect 4107 20936 4149 20945
rect 4107 20896 4108 20936
rect 4148 20896 4149 20936
rect 4107 20887 4149 20896
rect 3628 20773 3668 20782
rect 3628 20693 3668 20733
rect 4108 20768 4148 20887
rect 4108 20719 4148 20728
rect 3627 20684 3669 20693
rect 3627 20644 3628 20684
rect 3668 20644 3669 20684
rect 3627 20635 3669 20644
rect 4204 20600 4244 21148
rect 4299 21020 4341 21029
rect 4299 20980 4300 21020
rect 4340 20980 4341 21020
rect 4299 20971 4341 20980
rect 4012 20560 4244 20600
rect 3531 20264 3573 20273
rect 3531 20224 3532 20264
rect 3572 20224 3573 20264
rect 3531 20215 3573 20224
rect 3532 20096 3572 20105
rect 3532 20012 3572 20056
rect 3916 20096 3956 20105
rect 3532 19972 3860 20012
rect 3820 19853 3860 19972
rect 3916 19937 3956 20056
rect 4012 20096 4052 20560
rect 4012 20047 4052 20056
rect 4108 20096 4148 20107
rect 4108 20021 4148 20056
rect 4107 20012 4149 20021
rect 4107 19972 4108 20012
rect 4148 19972 4149 20012
rect 4107 19963 4149 19972
rect 3915 19928 3957 19937
rect 3915 19888 3916 19928
rect 3956 19888 3957 19928
rect 3915 19879 3957 19888
rect 3724 19844 3764 19853
rect 3532 19804 3724 19844
rect 3532 19256 3572 19804
rect 3724 19795 3764 19804
rect 3819 19844 3861 19853
rect 3819 19804 3820 19844
rect 3860 19804 3861 19844
rect 3819 19795 3861 19804
rect 3688 19676 4056 19685
rect 3728 19636 3770 19676
rect 3810 19636 3852 19676
rect 3892 19636 3934 19676
rect 3974 19636 4016 19676
rect 3688 19627 4056 19636
rect 3819 19340 3861 19349
rect 3819 19300 3820 19340
rect 3860 19300 3861 19340
rect 3819 19291 3861 19300
rect 3724 19256 3764 19265
rect 3532 19216 3724 19256
rect 3724 19207 3764 19216
rect 3820 19256 3860 19291
rect 3820 19205 3860 19216
rect 3915 19256 3957 19265
rect 3915 19216 3916 19256
rect 3956 19216 3957 19256
rect 3915 19207 3957 19216
rect 4108 19256 4148 19265
rect 3916 19122 3956 19207
rect 3628 19088 3668 19097
rect 3436 19048 3628 19088
rect 3628 19039 3668 19048
rect 4108 18845 4148 19216
rect 4107 18836 4149 18845
rect 3340 18796 3476 18836
rect 3339 18668 3381 18677
rect 3339 18628 3340 18668
rect 3380 18628 3381 18668
rect 3339 18619 3381 18628
rect 3243 18584 3285 18593
rect 3243 18544 3244 18584
rect 3284 18544 3285 18584
rect 3243 18535 3285 18544
rect 2956 18500 2996 18509
rect 2859 17408 2901 17417
rect 2859 17368 2860 17408
rect 2900 17368 2901 17408
rect 2859 17359 2901 17368
rect 2668 17240 2708 17249
rect 2476 17200 2668 17240
rect 2668 17191 2708 17200
rect 2475 17072 2517 17081
rect 2475 17032 2476 17072
rect 2516 17032 2517 17072
rect 2475 17023 2517 17032
rect 2476 15560 2516 17023
rect 2859 16988 2901 16997
rect 2859 16948 2860 16988
rect 2900 16948 2901 16988
rect 2859 16939 2901 16948
rect 2860 16484 2900 16939
rect 2860 16435 2900 16444
rect 2668 16232 2708 16241
rect 2476 15485 2516 15520
rect 2572 16192 2668 16232
rect 2475 15476 2517 15485
rect 2475 15436 2476 15476
rect 2516 15436 2517 15476
rect 2475 15427 2517 15436
rect 2572 15140 2612 16192
rect 2668 16183 2708 16192
rect 2763 16232 2805 16241
rect 2763 16192 2764 16232
rect 2804 16192 2805 16232
rect 2763 16183 2805 16192
rect 2668 15728 2708 15737
rect 2764 15728 2804 16183
rect 2859 16064 2901 16073
rect 2859 16024 2860 16064
rect 2900 16024 2901 16064
rect 2859 16015 2901 16024
rect 2860 15930 2900 16015
rect 2708 15688 2804 15728
rect 2668 15679 2708 15688
rect 2859 15308 2901 15317
rect 2859 15268 2860 15308
rect 2900 15268 2901 15308
rect 2859 15259 2901 15268
rect 2476 15100 2612 15140
rect 2379 15056 2421 15065
rect 2379 15016 2380 15056
rect 2420 15016 2421 15056
rect 2379 15007 2421 15016
rect 2476 14720 2516 15100
rect 2860 14972 2900 15259
rect 2956 15149 2996 18460
rect 3052 18500 3092 18509
rect 3052 17417 3092 18460
rect 3147 18248 3189 18257
rect 3147 18208 3148 18248
rect 3188 18208 3189 18248
rect 3147 18199 3189 18208
rect 3051 17408 3093 17417
rect 3051 17368 3052 17408
rect 3092 17368 3093 17408
rect 3051 17359 3093 17368
rect 3051 17240 3093 17249
rect 3051 17200 3052 17240
rect 3092 17200 3093 17240
rect 3051 17191 3093 17200
rect 3052 17072 3092 17191
rect 3052 16829 3092 17032
rect 3051 16820 3093 16829
rect 3051 16780 3052 16820
rect 3092 16780 3093 16820
rect 3051 16771 3093 16780
rect 3051 16064 3093 16073
rect 3051 16024 3052 16064
rect 3092 16024 3093 16064
rect 3051 16015 3093 16024
rect 3052 15569 3092 16015
rect 3051 15560 3093 15569
rect 3051 15520 3052 15560
rect 3092 15520 3093 15560
rect 3051 15511 3093 15520
rect 3148 15560 3188 18199
rect 3244 15728 3284 18535
rect 3340 17249 3380 18619
rect 3339 17240 3381 17249
rect 3339 17200 3340 17240
rect 3380 17200 3381 17240
rect 3339 17191 3381 17200
rect 3340 17072 3380 17083
rect 3340 16997 3380 17032
rect 3339 16988 3381 16997
rect 3339 16948 3340 16988
rect 3380 16948 3381 16988
rect 3339 16939 3381 16948
rect 3340 16820 3380 16829
rect 3340 16493 3380 16780
rect 3339 16484 3381 16493
rect 3339 16444 3340 16484
rect 3380 16444 3381 16484
rect 3339 16435 3381 16444
rect 3436 16409 3476 18796
rect 4107 18796 4108 18836
rect 4148 18796 4149 18836
rect 4107 18787 4149 18796
rect 4203 18752 4245 18761
rect 4203 18712 4204 18752
rect 4244 18712 4245 18752
rect 4203 18703 4245 18712
rect 4204 18618 4244 18703
rect 3532 18584 3572 18593
rect 3532 18257 3572 18544
rect 4012 18570 4052 18579
rect 4012 18332 4052 18530
rect 4012 18292 4148 18332
rect 3531 18248 3573 18257
rect 3531 18208 3532 18248
rect 3572 18208 3573 18248
rect 3531 18199 3573 18208
rect 3688 18164 4056 18173
rect 3728 18124 3770 18164
rect 3810 18124 3852 18164
rect 3892 18124 3934 18164
rect 3974 18124 4016 18164
rect 3688 18115 4056 18124
rect 4012 17996 4052 18005
rect 4108 17996 4148 18292
rect 4052 17956 4148 17996
rect 4012 17947 4052 17956
rect 3820 17744 3860 17753
rect 3531 17156 3573 17165
rect 3531 17116 3532 17156
rect 3572 17116 3573 17156
rect 3531 17107 3573 17116
rect 3532 17072 3572 17107
rect 3820 17081 3860 17704
rect 3532 16661 3572 17032
rect 3819 17072 3861 17081
rect 3819 17032 3820 17072
rect 3860 17032 3861 17072
rect 3819 17023 3861 17032
rect 3531 16652 3573 16661
rect 3531 16612 3532 16652
rect 3572 16612 3573 16652
rect 3531 16603 3573 16612
rect 3688 16652 4056 16661
rect 3728 16612 3770 16652
rect 3810 16612 3852 16652
rect 3892 16612 3934 16652
rect 3974 16612 4016 16652
rect 3688 16603 4056 16612
rect 3627 16484 3669 16493
rect 3627 16444 3628 16484
rect 3668 16444 3669 16484
rect 3627 16435 3669 16444
rect 3819 16484 3861 16493
rect 4300 16484 4340 20971
rect 4588 20852 4628 21232
rect 4684 20861 4724 21316
rect 5451 21316 5452 21356
rect 5492 21316 5493 21356
rect 5451 21307 5493 21316
rect 5452 21222 5492 21307
rect 5548 21029 5588 22903
rect 5644 22868 5684 22879
rect 5644 22793 5684 22828
rect 5643 22784 5685 22793
rect 5643 22744 5644 22784
rect 5684 22744 5685 22784
rect 5643 22735 5685 22744
rect 5643 22616 5685 22625
rect 5643 22576 5644 22616
rect 5684 22576 5685 22616
rect 5643 22567 5685 22576
rect 5644 21701 5684 22567
rect 5740 21785 5780 23995
rect 5836 23801 5876 26599
rect 5835 23792 5877 23801
rect 5835 23752 5836 23792
rect 5876 23752 5877 23792
rect 5835 23743 5877 23752
rect 5932 23288 5972 26683
rect 6028 24968 6068 27532
rect 6124 27572 6164 27581
rect 6219 27572 6261 27581
rect 6164 27532 6220 27572
rect 6260 27532 6261 27572
rect 6124 27523 6164 27532
rect 6219 27523 6261 27532
rect 6124 26816 6164 26827
rect 6124 26741 6164 26776
rect 6123 26732 6165 26741
rect 6123 26692 6124 26732
rect 6164 26692 6165 26732
rect 6123 26683 6165 26692
rect 6123 26564 6165 26573
rect 6123 26524 6124 26564
rect 6164 26524 6165 26564
rect 6123 26515 6165 26524
rect 6124 25145 6164 26515
rect 6220 26153 6260 27523
rect 6316 26489 6356 29707
rect 6412 29706 6452 29791
rect 6508 27656 6548 30472
rect 7276 29849 7316 31312
rect 7372 31326 7508 31366
rect 7756 31352 7796 31361
rect 7372 30848 7412 31326
rect 7468 31268 7508 31277
rect 7756 31268 7796 31312
rect 7852 31352 7892 31361
rect 7892 31312 7988 31352
rect 7852 31303 7892 31312
rect 7508 31228 7796 31268
rect 7468 31219 7508 31228
rect 7468 30848 7508 30857
rect 7372 30808 7468 30848
rect 7468 30799 7508 30808
rect 7371 30680 7413 30689
rect 7371 30640 7372 30680
rect 7412 30640 7413 30680
rect 7371 30631 7413 30640
rect 7372 30546 7412 30631
rect 7948 30260 7988 31312
rect 8236 31302 8276 31387
rect 8332 31352 8372 31361
rect 8332 31193 8372 31312
rect 8331 31184 8373 31193
rect 8331 31144 8332 31184
rect 8372 31144 8373 31184
rect 8331 31135 8373 31144
rect 7948 30220 8180 30260
rect 7371 30008 7413 30017
rect 7371 29968 7372 30008
rect 7412 29968 7413 30008
rect 7371 29959 7413 29968
rect 7851 30008 7893 30017
rect 7851 29968 7852 30008
rect 7892 29968 7893 30008
rect 7851 29959 7893 29968
rect 7372 29924 7412 29959
rect 7372 29873 7412 29884
rect 7467 29924 7509 29933
rect 7467 29884 7468 29924
rect 7508 29884 7509 29924
rect 7467 29875 7509 29884
rect 6892 29840 6932 29849
rect 6604 29756 6644 29765
rect 6892 29756 6932 29800
rect 6644 29716 6932 29756
rect 6988 29840 7028 29849
rect 6604 29707 6644 29716
rect 6988 29420 7028 29800
rect 7275 29840 7317 29849
rect 7275 29800 7276 29840
rect 7316 29800 7317 29840
rect 7275 29791 7317 29800
rect 7468 29790 7508 29875
rect 6796 29380 7028 29420
rect 6699 28412 6741 28421
rect 6699 28372 6700 28412
rect 6740 28372 6741 28412
rect 6699 28363 6741 28372
rect 6604 27656 6644 27665
rect 6508 27616 6604 27656
rect 6507 26900 6549 26909
rect 6507 26860 6508 26900
rect 6548 26860 6549 26900
rect 6507 26851 6549 26860
rect 6315 26480 6357 26489
rect 6315 26440 6316 26480
rect 6356 26440 6357 26480
rect 6315 26431 6357 26440
rect 6219 26144 6261 26153
rect 6219 26104 6220 26144
rect 6260 26104 6261 26144
rect 6219 26095 6261 26104
rect 6123 25136 6165 25145
rect 6123 25096 6124 25136
rect 6164 25096 6165 25136
rect 6123 25087 6165 25096
rect 6220 24977 6260 26095
rect 6219 24968 6261 24977
rect 6028 24928 6164 24968
rect 6027 23708 6069 23717
rect 6027 23668 6028 23708
rect 6068 23668 6069 23708
rect 6027 23659 6069 23668
rect 6028 23465 6068 23659
rect 6027 23456 6069 23465
rect 6027 23416 6028 23456
rect 6068 23416 6069 23456
rect 6027 23407 6069 23416
rect 6124 23297 6164 24928
rect 6219 24928 6220 24968
rect 6260 24928 6261 24968
rect 6219 24919 6261 24928
rect 6508 24632 6548 26851
rect 6604 25985 6644 27616
rect 6700 27404 6740 28363
rect 6796 27581 6836 29380
rect 6891 29252 6933 29261
rect 6891 29212 6892 29252
rect 6932 29212 6933 29252
rect 6891 29203 6933 29212
rect 6795 27572 6837 27581
rect 6795 27532 6796 27572
rect 6836 27532 6837 27572
rect 6795 27523 6837 27532
rect 6892 27497 6932 29203
rect 6987 29168 7029 29177
rect 6987 29128 6988 29168
rect 7028 29128 7029 29168
rect 6987 29119 7029 29128
rect 6988 29034 7028 29119
rect 7755 28412 7797 28421
rect 7755 28372 7756 28412
rect 7796 28372 7797 28412
rect 7755 28363 7797 28372
rect 7180 28328 7220 28337
rect 6987 27656 7029 27665
rect 6987 27616 6988 27656
rect 7028 27616 7029 27656
rect 6987 27607 7029 27616
rect 7084 27642 7124 27651
rect 6891 27488 6933 27497
rect 6891 27448 6892 27488
rect 6932 27448 6933 27488
rect 6891 27439 6933 27448
rect 6700 27364 6836 27404
rect 6699 26816 6741 26825
rect 6699 26776 6700 26816
rect 6740 26776 6741 26816
rect 6699 26767 6741 26776
rect 6700 26573 6740 26767
rect 6699 26564 6741 26573
rect 6699 26524 6700 26564
rect 6740 26524 6741 26564
rect 6699 26515 6741 26524
rect 6700 26144 6740 26515
rect 6796 26153 6836 27364
rect 6988 26480 7028 27607
rect 7084 27077 7124 27602
rect 7083 27068 7125 27077
rect 7083 27028 7084 27068
rect 7124 27028 7125 27068
rect 7083 27019 7125 27028
rect 7180 26816 7220 28288
rect 7756 28328 7796 28363
rect 7372 28160 7412 28169
rect 7412 28120 7508 28160
rect 7372 28111 7412 28120
rect 7276 27740 7316 27749
rect 7276 27497 7316 27700
rect 7468 27656 7508 28120
rect 7564 27656 7604 27665
rect 7468 27616 7564 27656
rect 7564 27607 7604 27616
rect 7659 27656 7701 27665
rect 7659 27616 7660 27656
rect 7700 27616 7701 27656
rect 7659 27607 7701 27616
rect 7660 27522 7700 27607
rect 7275 27488 7317 27497
rect 7275 27448 7276 27488
rect 7316 27448 7317 27488
rect 7275 27439 7317 27448
rect 7467 27404 7509 27413
rect 7467 27364 7468 27404
rect 7508 27364 7509 27404
rect 7467 27355 7509 27364
rect 7372 26816 7412 26825
rect 7180 26776 7372 26816
rect 7372 26573 7412 26776
rect 7371 26564 7413 26573
rect 7371 26524 7372 26564
rect 7412 26524 7413 26564
rect 7371 26515 7413 26524
rect 7275 26480 7317 26489
rect 6988 26440 7220 26480
rect 6700 26095 6740 26104
rect 6795 26144 6837 26153
rect 6795 26104 6796 26144
rect 6836 26104 6837 26144
rect 6795 26095 6837 26104
rect 7083 26144 7125 26153
rect 7083 26104 7084 26144
rect 7124 26104 7125 26144
rect 7083 26095 7125 26104
rect 7084 26010 7124 26095
rect 6603 25976 6645 25985
rect 6603 25936 6604 25976
rect 6644 25936 6645 25976
rect 6603 25927 6645 25936
rect 6795 25892 6837 25901
rect 6795 25852 6796 25892
rect 6836 25852 6837 25892
rect 6795 25843 6837 25852
rect 6892 25892 6932 25901
rect 6932 25852 7028 25892
rect 6892 25843 6932 25852
rect 6700 24716 6740 24727
rect 6700 24641 6740 24676
rect 6699 24632 6741 24641
rect 6508 23801 6548 24592
rect 6604 24592 6700 24632
rect 6740 24592 6741 24632
rect 6507 23792 6549 23801
rect 6507 23752 6508 23792
rect 6548 23752 6549 23792
rect 6507 23743 6549 23752
rect 5836 23248 5972 23288
rect 6123 23288 6165 23297
rect 6123 23248 6124 23288
rect 6164 23248 6165 23288
rect 5739 21776 5781 21785
rect 5739 21736 5740 21776
rect 5780 21736 5781 21776
rect 5739 21727 5781 21736
rect 5643 21692 5685 21701
rect 5643 21652 5644 21692
rect 5684 21652 5685 21692
rect 5643 21643 5685 21652
rect 5644 21608 5684 21643
rect 5644 21557 5684 21568
rect 5739 21608 5781 21617
rect 5739 21568 5740 21608
rect 5780 21568 5781 21608
rect 5739 21559 5781 21568
rect 5547 21020 5589 21029
rect 5547 20980 5548 21020
rect 5588 20980 5589 21020
rect 5547 20971 5589 20980
rect 4588 20600 4628 20812
rect 4683 20852 4725 20861
rect 4683 20812 4684 20852
rect 4724 20812 4725 20852
rect 4683 20803 4725 20812
rect 4684 20718 4724 20803
rect 5067 20768 5109 20777
rect 5067 20728 5068 20768
rect 5108 20728 5109 20768
rect 5067 20719 5109 20728
rect 5164 20768 5204 20777
rect 5204 20728 5396 20768
rect 5164 20719 5204 20728
rect 5068 20634 5108 20719
rect 4588 20560 4820 20600
rect 4683 20348 4725 20357
rect 4683 20308 4684 20348
rect 4724 20308 4725 20348
rect 4683 20299 4725 20308
rect 4395 20096 4437 20105
rect 4395 20056 4396 20096
rect 4436 20056 4437 20096
rect 4395 20047 4437 20056
rect 4588 20096 4628 20107
rect 4396 19962 4436 20047
rect 4588 20021 4628 20056
rect 4684 20096 4724 20299
rect 4684 20047 4724 20056
rect 4587 20012 4629 20021
rect 4587 19972 4588 20012
rect 4628 19972 4629 20012
rect 4587 19963 4629 19972
rect 4491 19928 4533 19937
rect 4491 19888 4492 19928
rect 4532 19888 4533 19928
rect 4491 19879 4533 19888
rect 4396 19844 4436 19853
rect 4396 19349 4436 19804
rect 4395 19340 4437 19349
rect 4395 19300 4396 19340
rect 4436 19300 4437 19340
rect 4395 19291 4437 19300
rect 4492 19265 4532 19879
rect 4491 19256 4533 19265
rect 4491 19216 4492 19256
rect 4532 19216 4533 19256
rect 4491 19207 4533 19216
rect 4780 17240 4820 20560
rect 4928 20432 5296 20441
rect 4968 20392 5010 20432
rect 5050 20392 5092 20432
rect 5132 20392 5174 20432
rect 5214 20392 5256 20432
rect 4928 20383 5296 20392
rect 5356 20264 5396 20728
rect 5260 20224 5396 20264
rect 5260 19937 5300 20224
rect 5355 20096 5397 20105
rect 5355 20056 5356 20096
rect 5396 20056 5397 20096
rect 5355 20047 5397 20056
rect 5356 19962 5396 20047
rect 5259 19928 5301 19937
rect 5259 19888 5260 19928
rect 5300 19888 5301 19928
rect 5259 19879 5301 19888
rect 5355 19256 5397 19265
rect 5355 19216 5356 19256
rect 5396 19216 5397 19256
rect 5355 19207 5397 19216
rect 5356 19122 5396 19207
rect 5548 19088 5588 19097
rect 5452 19048 5548 19088
rect 4928 18920 5296 18929
rect 4968 18880 5010 18920
rect 5050 18880 5092 18920
rect 5132 18880 5174 18920
rect 5214 18880 5256 18920
rect 4928 18871 5296 18880
rect 5163 18752 5205 18761
rect 5163 18712 5164 18752
rect 5204 18712 5205 18752
rect 5163 18703 5205 18712
rect 5164 17576 5204 18703
rect 5452 18584 5492 19048
rect 5548 19039 5588 19048
rect 5740 18920 5780 21559
rect 5452 18535 5492 18544
rect 5548 18880 5780 18920
rect 5548 18584 5588 18880
rect 5548 18509 5588 18544
rect 5547 18500 5589 18509
rect 5547 18460 5548 18500
rect 5588 18460 5589 18500
rect 5547 18451 5589 18460
rect 5548 18420 5588 18451
rect 5259 17912 5301 17921
rect 5259 17872 5260 17912
rect 5300 17872 5301 17912
rect 5259 17863 5301 17872
rect 5260 17744 5300 17863
rect 5260 17695 5300 17704
rect 5164 17536 5396 17576
rect 4928 17408 5296 17417
rect 4968 17368 5010 17408
rect 5050 17368 5092 17408
rect 5132 17368 5174 17408
rect 5214 17368 5256 17408
rect 4928 17359 5296 17368
rect 5356 17240 5396 17536
rect 3819 16444 3820 16484
rect 3860 16444 3861 16484
rect 3819 16435 3861 16444
rect 4012 16444 4340 16484
rect 4684 17200 4820 17240
rect 5164 17200 5396 17240
rect 5548 17240 5588 17249
rect 3435 16400 3477 16409
rect 3435 16360 3436 16400
rect 3476 16360 3477 16400
rect 3435 16351 3477 16360
rect 3340 16241 3380 16326
rect 3339 16232 3381 16241
rect 3339 16192 3340 16232
rect 3380 16192 3381 16232
rect 3339 16183 3381 16192
rect 3436 16232 3476 16241
rect 3244 15688 3380 15728
rect 2955 15140 2997 15149
rect 2955 15100 2956 15140
rect 2996 15100 2997 15140
rect 2955 15091 2997 15100
rect 2860 14923 2900 14932
rect 3052 14720 3092 15511
rect 3148 15401 3188 15520
rect 3244 15560 3284 15569
rect 3147 15392 3189 15401
rect 3147 15352 3148 15392
rect 3188 15352 3189 15392
rect 3147 15343 3189 15352
rect 3244 14897 3284 15520
rect 3243 14888 3285 14897
rect 3243 14848 3244 14888
rect 3284 14848 3285 14888
rect 3243 14839 3285 14848
rect 2476 12872 2516 14680
rect 2860 14680 3092 14720
rect 3244 14720 3284 14729
rect 2667 14552 2709 14561
rect 2667 14512 2668 14552
rect 2708 14512 2709 14552
rect 2667 14503 2709 14512
rect 2668 14418 2708 14503
rect 2763 14384 2805 14393
rect 2763 14344 2764 14384
rect 2804 14344 2805 14384
rect 2763 14335 2805 14344
rect 2668 14216 2708 14225
rect 2764 14216 2804 14335
rect 2708 14176 2804 14216
rect 2668 14167 2708 14176
rect 2860 14043 2900 14680
rect 3147 14636 3189 14645
rect 3147 14596 3148 14636
rect 3188 14596 3189 14636
rect 3147 14587 3189 14596
rect 3148 14502 3188 14587
rect 3244 14393 3284 14680
rect 3243 14384 3285 14393
rect 3243 14344 3244 14384
rect 3284 14344 3285 14384
rect 3243 14335 3285 14344
rect 3340 14225 3380 15688
rect 3436 15485 3476 16192
rect 3628 15560 3668 16435
rect 3820 16316 3860 16435
rect 3820 16267 3860 16276
rect 3915 16316 3957 16325
rect 3915 16276 3916 16316
rect 3956 16276 3957 16316
rect 3915 16267 3957 16276
rect 3916 16182 3956 16267
rect 3628 15511 3668 15520
rect 3819 15560 3861 15569
rect 3819 15520 3820 15560
rect 3860 15520 3861 15560
rect 3819 15511 3861 15520
rect 3916 15560 3956 15569
rect 4012 15560 4052 16444
rect 4491 16400 4533 16409
rect 4491 16360 4492 16400
rect 4532 16360 4533 16400
rect 4491 16351 4533 16360
rect 4396 16232 4436 16241
rect 4396 16073 4436 16192
rect 4395 16064 4437 16073
rect 4395 16024 4396 16064
rect 4436 16024 4437 16064
rect 4395 16015 4437 16024
rect 4299 15812 4341 15821
rect 4299 15772 4300 15812
rect 4340 15772 4341 15812
rect 4299 15763 4341 15772
rect 4203 15728 4245 15737
rect 4203 15688 4204 15728
rect 4244 15688 4245 15728
rect 4203 15679 4245 15688
rect 4108 15569 4148 15654
rect 4204 15594 4244 15679
rect 3956 15520 4052 15560
rect 4107 15560 4149 15569
rect 4107 15520 4108 15560
rect 4148 15520 4149 15560
rect 3916 15511 3956 15520
rect 4107 15511 4149 15520
rect 4300 15560 4340 15763
rect 4300 15511 4340 15520
rect 4396 15560 4436 15569
rect 4492 15560 4532 16351
rect 4587 15812 4629 15821
rect 4587 15772 4588 15812
rect 4628 15772 4629 15812
rect 4587 15763 4629 15772
rect 4588 15728 4628 15763
rect 4588 15677 4628 15688
rect 4436 15520 4532 15560
rect 4396 15511 4436 15520
rect 3435 15476 3477 15485
rect 3435 15436 3436 15476
rect 3476 15436 3477 15476
rect 3435 15427 3477 15436
rect 3820 15426 3860 15511
rect 3628 15317 3668 15402
rect 4491 15392 4533 15401
rect 4491 15352 4492 15392
rect 4532 15352 4533 15392
rect 4491 15343 4533 15352
rect 3436 15308 3476 15317
rect 3436 15140 3476 15268
rect 3627 15308 3669 15317
rect 3627 15268 3628 15308
rect 3668 15268 3669 15308
rect 3627 15259 3669 15268
rect 4107 15308 4149 15317
rect 4107 15268 4108 15308
rect 4148 15268 4149 15308
rect 4107 15259 4149 15268
rect 3688 15140 4056 15149
rect 3436 15100 3572 15140
rect 3532 14972 3572 15100
rect 3728 15100 3770 15140
rect 3810 15100 3852 15140
rect 3892 15100 3934 15140
rect 3974 15100 4016 15140
rect 3688 15091 4056 15100
rect 4108 14972 4148 15259
rect 3532 14932 3956 14972
rect 3532 14720 3572 14729
rect 3532 14561 3572 14680
rect 3916 14720 3956 14932
rect 3916 14671 3956 14680
rect 4012 14932 4148 14972
rect 4012 14720 4052 14932
rect 4108 14813 4148 14844
rect 4107 14804 4149 14813
rect 4107 14764 4108 14804
rect 4148 14764 4149 14804
rect 4107 14755 4149 14764
rect 4012 14671 4052 14680
rect 4108 14720 4148 14755
rect 3819 14636 3861 14645
rect 3819 14596 3820 14636
rect 3860 14596 3861 14636
rect 3819 14587 3861 14596
rect 3531 14552 3573 14561
rect 3531 14512 3532 14552
rect 3572 14512 3573 14552
rect 3531 14503 3573 14512
rect 3820 14502 3860 14587
rect 3531 14384 3573 14393
rect 3531 14344 3532 14384
rect 3572 14344 3573 14384
rect 3531 14335 3573 14344
rect 2955 14216 2997 14225
rect 2955 14176 2956 14216
rect 2996 14176 2997 14216
rect 2955 14167 2997 14176
rect 3339 14216 3381 14225
rect 3339 14176 3340 14216
rect 3380 14176 3381 14216
rect 3339 14167 3381 14176
rect 2860 13994 2900 14003
rect 2859 13880 2901 13889
rect 2859 13840 2860 13880
rect 2900 13840 2901 13880
rect 2859 13831 2901 13840
rect 2764 13213 2804 13222
rect 2571 13124 2613 13133
rect 2571 13084 2572 13124
rect 2612 13084 2613 13124
rect 2571 13075 2613 13084
rect 2572 12990 2612 13075
rect 2476 12832 2612 12872
rect 2284 12748 2516 12788
rect 2283 12620 2325 12629
rect 2283 12580 2284 12620
rect 2324 12580 2325 12620
rect 2283 12571 2325 12580
rect 2284 12486 2324 12571
rect 2476 12545 2516 12748
rect 2475 12536 2517 12545
rect 2475 12496 2476 12536
rect 2516 12496 2517 12536
rect 2475 12487 2517 12496
rect 2283 12368 2325 12377
rect 2572 12368 2612 12832
rect 2764 12629 2804 13173
rect 2763 12620 2805 12629
rect 2763 12580 2764 12620
rect 2804 12580 2805 12620
rect 2763 12571 2805 12580
rect 2283 12328 2284 12368
rect 2324 12328 2325 12368
rect 2283 12319 2325 12328
rect 2476 12328 2612 12368
rect 2187 11024 2229 11033
rect 2187 10984 2188 11024
rect 2228 10984 2229 11024
rect 2187 10975 2229 10984
rect 2284 11024 2324 12319
rect 2476 11705 2516 12328
rect 2668 11948 2708 11957
rect 2860 11948 2900 13831
rect 2708 11908 2900 11948
rect 2668 11899 2708 11908
rect 2475 11696 2517 11705
rect 2475 11656 2476 11696
rect 2516 11656 2517 11696
rect 2475 11647 2517 11656
rect 2476 11562 2516 11647
rect 2667 11276 2709 11285
rect 2667 11236 2668 11276
rect 2708 11236 2709 11276
rect 2667 11227 2709 11236
rect 2668 11192 2708 11227
rect 2668 11141 2708 11152
rect 2476 11024 2516 11033
rect 2284 10984 2476 11024
rect 2284 10352 2324 10984
rect 2476 10975 2516 10984
rect 2571 10772 2613 10781
rect 2571 10732 2572 10772
rect 2612 10732 2613 10772
rect 2571 10723 2613 10732
rect 2188 10312 2324 10352
rect 2091 10184 2133 10193
rect 2091 10144 2092 10184
rect 2132 10144 2133 10184
rect 2091 10135 2133 10144
rect 2188 9605 2228 10312
rect 2475 10268 2517 10277
rect 2475 10228 2476 10268
rect 2516 10228 2517 10268
rect 2475 10219 2517 10228
rect 2283 10184 2325 10193
rect 2283 10144 2284 10184
rect 2324 10144 2325 10184
rect 2283 10135 2325 10144
rect 2476 10184 2516 10219
rect 2187 9596 2229 9605
rect 2187 9556 2188 9596
rect 2228 9556 2229 9596
rect 2187 9547 2229 9556
rect 1708 8632 2036 8672
rect 1708 3212 1748 8632
rect 1996 8009 2036 8094
rect 1995 8000 2037 8009
rect 1995 7960 1996 8000
rect 2036 7960 2037 8000
rect 1995 7951 2037 7960
rect 2092 8000 2132 8009
rect 1995 7832 2037 7841
rect 1995 7792 1996 7832
rect 2036 7792 2037 7832
rect 1995 7783 2037 7792
rect 1803 6992 1845 7001
rect 1803 6952 1804 6992
rect 1844 6952 1845 6992
rect 1803 6943 1845 6952
rect 1804 5648 1844 6943
rect 1804 5599 1844 5608
rect 1900 5648 1940 5657
rect 1900 5489 1940 5608
rect 1899 5480 1941 5489
rect 1899 5440 1900 5480
rect 1940 5440 1941 5480
rect 1899 5431 1941 5440
rect 1996 4649 2036 7783
rect 2092 7505 2132 7960
rect 2187 8000 2229 8009
rect 2187 7960 2188 8000
rect 2228 7960 2229 8000
rect 2187 7951 2229 7960
rect 2188 7866 2228 7951
rect 2091 7496 2133 7505
rect 2091 7456 2092 7496
rect 2132 7456 2133 7496
rect 2091 7447 2133 7456
rect 2091 5984 2133 5993
rect 2091 5944 2092 5984
rect 2132 5944 2133 5984
rect 2091 5935 2133 5944
rect 1995 4640 2037 4649
rect 1995 4600 1996 4640
rect 2036 4600 2037 4640
rect 1995 4591 2037 4600
rect 1995 3716 2037 3725
rect 1995 3676 1996 3716
rect 2036 3676 2037 3716
rect 1995 3667 2037 3676
rect 1708 3172 1940 3212
rect 1611 3128 1653 3137
rect 1611 3088 1612 3128
rect 1652 3088 1653 3128
rect 1611 3079 1653 3088
rect 459 2792 501 2801
rect 459 2752 460 2792
rect 500 2752 501 2792
rect 459 2743 501 2752
rect 1611 2624 1653 2633
rect 1611 2584 1612 2624
rect 1652 2584 1653 2624
rect 1611 2575 1653 2584
rect 1804 2624 1844 2633
rect 1612 2490 1652 2575
rect 1707 2540 1749 2549
rect 1707 2500 1708 2540
rect 1748 2500 1749 2540
rect 1707 2491 1749 2500
rect 1708 2406 1748 2491
rect 1323 1952 1365 1961
rect 1323 1912 1324 1952
rect 1364 1912 1365 1952
rect 1323 1903 1365 1912
rect 1324 1818 1364 1903
rect 1804 1709 1844 2584
rect 1803 1700 1845 1709
rect 1803 1660 1804 1700
rect 1844 1660 1845 1700
rect 1803 1651 1845 1660
rect 1803 1532 1845 1541
rect 1803 1492 1804 1532
rect 1844 1492 1845 1532
rect 1803 1483 1845 1492
rect 1804 188 1844 1483
rect 1900 281 1940 3172
rect 1996 2624 2036 3667
rect 1996 2575 2036 2584
rect 2092 1541 2132 5935
rect 2188 5648 2228 5657
rect 2188 4817 2228 5608
rect 2284 5069 2324 10135
rect 2476 9437 2516 10144
rect 2475 9428 2517 9437
rect 2475 9388 2476 9428
rect 2516 9388 2517 9428
rect 2475 9379 2517 9388
rect 2476 8672 2516 9379
rect 2380 7748 2420 7757
rect 2380 6497 2420 7708
rect 2476 7169 2516 8632
rect 2572 7589 2612 10723
rect 2667 10604 2709 10613
rect 2667 10564 2668 10604
rect 2708 10564 2709 10604
rect 2667 10555 2709 10564
rect 2668 10436 2708 10555
rect 2668 10387 2708 10396
rect 2859 10100 2901 10109
rect 2859 10060 2860 10100
rect 2900 10060 2901 10100
rect 2859 10051 2901 10060
rect 2860 9966 2900 10051
rect 2956 9764 2996 14167
rect 3340 14048 3380 14057
rect 3243 13796 3285 13805
rect 3243 13756 3244 13796
rect 3284 13756 3285 13796
rect 3243 13747 3285 13756
rect 3244 13208 3284 13747
rect 3340 13721 3380 14008
rect 3339 13712 3381 13721
rect 3339 13672 3340 13712
rect 3380 13672 3381 13712
rect 3339 13663 3381 13672
rect 3244 12125 3284 13168
rect 3532 12545 3572 14335
rect 3915 14216 3957 14225
rect 3915 14176 3916 14216
rect 3956 14176 3957 14216
rect 3915 14167 3957 14176
rect 3916 14048 3956 14167
rect 3916 13999 3956 14008
rect 4108 13973 4148 14680
rect 4396 14720 4436 14729
rect 4396 14561 4436 14680
rect 4395 14552 4437 14561
rect 4395 14512 4396 14552
rect 4436 14512 4437 14552
rect 4395 14503 4437 14512
rect 4300 14048 4340 14057
rect 4204 14008 4300 14048
rect 3820 13964 3860 13973
rect 3820 13796 3860 13924
rect 4107 13964 4149 13973
rect 4107 13924 4108 13964
rect 4148 13924 4149 13964
rect 4107 13915 4149 13924
rect 3820 13756 4148 13796
rect 3688 13628 4056 13637
rect 3728 13588 3770 13628
rect 3810 13588 3852 13628
rect 3892 13588 3934 13628
rect 3974 13588 4016 13628
rect 3688 13579 4056 13588
rect 4108 13217 4148 13756
rect 3723 13208 3765 13217
rect 3723 13168 3724 13208
rect 3764 13168 3765 13208
rect 3723 13159 3765 13168
rect 3820 13208 3860 13217
rect 3724 13074 3764 13159
rect 3531 12536 3573 12545
rect 3724 12536 3764 12545
rect 3531 12496 3532 12536
rect 3572 12496 3724 12536
rect 3531 12487 3573 12496
rect 3724 12487 3764 12496
rect 3532 12402 3572 12487
rect 3820 12293 3860 13168
rect 4107 13208 4149 13217
rect 4107 13168 4108 13208
rect 4148 13168 4149 13208
rect 4107 13159 4149 13168
rect 4204 13208 4244 14008
rect 4300 13999 4340 14008
rect 4396 14048 4436 14057
rect 4396 13889 4436 14008
rect 4395 13880 4437 13889
rect 4395 13840 4396 13880
rect 4436 13840 4437 13880
rect 4395 13831 4437 13840
rect 3915 12536 3957 12545
rect 3915 12496 3916 12536
rect 3956 12496 3957 12536
rect 3915 12487 3957 12496
rect 3916 12402 3956 12487
rect 3819 12284 3861 12293
rect 3819 12244 3820 12284
rect 3860 12244 3861 12284
rect 3819 12235 3861 12244
rect 3243 12116 3285 12125
rect 3243 12076 3244 12116
rect 3284 12076 3285 12116
rect 3243 12067 3285 12076
rect 3688 12116 4056 12125
rect 3728 12076 3770 12116
rect 3810 12076 3852 12116
rect 3892 12076 3934 12116
rect 3974 12076 4016 12116
rect 3688 12067 4056 12076
rect 3628 11696 3668 11705
rect 3532 11528 3572 11537
rect 3051 11192 3093 11201
rect 3051 11152 3052 11192
rect 3092 11152 3093 11192
rect 3051 11143 3093 11152
rect 3052 10856 3092 11143
rect 3340 11108 3380 11117
rect 3532 11108 3572 11488
rect 3380 11068 3572 11108
rect 3340 11059 3380 11068
rect 3052 10807 3092 10816
rect 3436 10982 3476 10991
rect 3051 10436 3093 10445
rect 3051 10396 3052 10436
rect 3092 10396 3093 10436
rect 3051 10387 3093 10396
rect 3052 10198 3092 10387
rect 3092 10158 3188 10198
rect 3052 10149 3092 10158
rect 2956 9724 3092 9764
rect 3052 9680 3092 9724
rect 3051 9640 3092 9680
rect 2956 9596 2996 9607
rect 3051 9596 3091 9640
rect 3051 9556 3092 9596
rect 2764 9512 2804 9523
rect 2956 9521 2996 9556
rect 2764 9437 2804 9472
rect 2955 9512 2997 9521
rect 2955 9472 2956 9512
rect 2996 9472 2997 9512
rect 2955 9463 2997 9472
rect 2763 9428 2805 9437
rect 2763 9388 2764 9428
rect 2804 9388 2805 9428
rect 3052 9428 3092 9556
rect 3148 9512 3188 10158
rect 3436 10109 3476 10942
rect 3628 10772 3668 11656
rect 3724 11696 3764 11705
rect 3724 11201 3764 11656
rect 3820 11696 3860 11705
rect 3723 11192 3765 11201
rect 3723 11152 3724 11192
rect 3764 11152 3765 11192
rect 3723 11143 3765 11152
rect 3724 11024 3764 11033
rect 3724 10865 3764 10984
rect 3723 10856 3765 10865
rect 3723 10816 3724 10856
rect 3764 10816 3765 10856
rect 3723 10807 3765 10816
rect 3820 10781 3860 11656
rect 3532 10732 3668 10772
rect 3819 10772 3861 10781
rect 3819 10732 3820 10772
rect 3860 10732 3861 10772
rect 3532 10352 3572 10732
rect 3819 10723 3861 10732
rect 3688 10604 4056 10613
rect 3728 10564 3770 10604
rect 3810 10564 3852 10604
rect 3892 10564 3934 10604
rect 3974 10564 4016 10604
rect 3688 10555 4056 10564
rect 4108 10352 4148 13159
rect 4204 10856 4244 13168
rect 4300 13208 4340 13217
rect 4300 11285 4340 13168
rect 4492 12209 4532 15343
rect 4587 14216 4629 14225
rect 4587 14176 4588 14216
rect 4628 14176 4629 14216
rect 4587 14167 4629 14176
rect 4491 12200 4533 12209
rect 4491 12160 4492 12200
rect 4532 12160 4533 12200
rect 4491 12151 4533 12160
rect 4588 11369 4628 14167
rect 4684 14141 4724 17200
rect 4779 17072 4821 17081
rect 4779 17032 4780 17072
rect 4820 17032 4821 17072
rect 4779 17023 4821 17032
rect 4780 16938 4820 17023
rect 4779 16820 4821 16829
rect 4972 16820 5012 16829
rect 4779 16780 4780 16820
rect 4820 16780 4821 16820
rect 4779 16771 4821 16780
rect 4876 16780 4972 16820
rect 4780 15728 4820 16771
rect 4876 16246 4916 16780
rect 4972 16771 5012 16780
rect 5164 16241 5204 17200
rect 5260 17072 5300 17081
rect 5260 16409 5300 17032
rect 5356 17072 5396 17081
rect 5259 16400 5301 16409
rect 5259 16360 5260 16400
rect 5300 16360 5301 16400
rect 5259 16351 5301 16360
rect 4876 16197 4916 16206
rect 5163 16232 5205 16241
rect 5260 16232 5300 16241
rect 5163 16192 5164 16232
rect 5204 16192 5260 16232
rect 5163 16183 5205 16192
rect 5260 16183 5300 16192
rect 5067 16148 5109 16157
rect 5067 16108 5068 16148
rect 5108 16108 5109 16148
rect 5067 16099 5109 16108
rect 5068 16014 5108 16099
rect 5164 16098 5204 16183
rect 4928 15896 5296 15905
rect 4968 15856 5010 15896
rect 5050 15856 5092 15896
rect 5132 15856 5174 15896
rect 5214 15856 5256 15896
rect 4928 15847 5296 15856
rect 4780 15688 4916 15728
rect 4779 15560 4821 15569
rect 4779 15520 4780 15560
rect 4820 15520 4821 15560
rect 4779 15511 4821 15520
rect 4683 14132 4725 14141
rect 4683 14092 4684 14132
rect 4724 14092 4725 14132
rect 4683 14083 4725 14092
rect 4587 11360 4629 11369
rect 4587 11320 4588 11360
rect 4628 11320 4629 11360
rect 4587 11311 4629 11320
rect 4299 11276 4341 11285
rect 4299 11236 4300 11276
rect 4340 11236 4341 11276
rect 4299 11227 4341 11236
rect 4396 11024 4436 11033
rect 4396 10865 4436 10984
rect 4491 11024 4533 11033
rect 4491 10984 4492 11024
rect 4532 10984 4533 11024
rect 4491 10975 4533 10984
rect 4684 11024 4724 11033
rect 4492 10890 4532 10975
rect 4395 10856 4437 10865
rect 4204 10816 4340 10856
rect 3532 10312 3764 10352
rect 3532 10184 3572 10193
rect 3435 10100 3477 10109
rect 3435 10060 3436 10100
rect 3476 10060 3477 10100
rect 3435 10051 3477 10060
rect 3532 10025 3572 10144
rect 3531 10016 3573 10025
rect 3531 9976 3532 10016
rect 3572 9976 3573 10016
rect 3531 9967 3573 9976
rect 3724 9680 3764 10312
rect 4012 10312 4148 10352
rect 4012 10184 4052 10312
rect 4012 9680 4052 10144
rect 4107 10184 4149 10193
rect 4107 10144 4108 10184
rect 4148 10144 4149 10184
rect 4300 10184 4340 10816
rect 4395 10816 4396 10856
rect 4436 10816 4437 10856
rect 4395 10807 4437 10816
rect 4396 10445 4436 10807
rect 4684 10781 4724 10984
rect 4491 10772 4533 10781
rect 4683 10772 4725 10781
rect 4491 10732 4492 10772
rect 4532 10732 4628 10772
rect 4491 10723 4533 10732
rect 4395 10436 4437 10445
rect 4395 10396 4396 10436
rect 4436 10396 4437 10436
rect 4395 10387 4437 10396
rect 4492 10184 4532 10193
rect 4300 10144 4492 10184
rect 4107 10135 4149 10144
rect 4108 10050 4148 10135
rect 4012 9640 4244 9680
rect 3724 9631 3764 9640
rect 3339 9512 3381 9521
rect 3148 9472 3340 9512
rect 3380 9472 3381 9512
rect 3339 9463 3381 9472
rect 3436 9512 3476 9523
rect 3052 9388 3284 9428
rect 2763 9379 2805 9388
rect 3147 9260 3189 9269
rect 3147 9220 3148 9260
rect 3188 9220 3189 9260
rect 3147 9211 3189 9220
rect 2667 8924 2709 8933
rect 2667 8884 2668 8924
rect 2708 8884 2709 8924
rect 2667 8875 2709 8884
rect 2668 8790 2708 8875
rect 3051 8840 3093 8849
rect 3051 8800 3052 8840
rect 3092 8800 3093 8840
rect 3051 8791 3093 8800
rect 3052 8706 3092 8791
rect 3051 8588 3093 8597
rect 3051 8548 3052 8588
rect 3092 8548 3093 8588
rect 3051 8539 3093 8548
rect 2955 8504 2997 8513
rect 2955 8464 2956 8504
rect 2996 8464 2997 8504
rect 2955 8455 2997 8464
rect 2667 8000 2709 8009
rect 2667 7960 2668 8000
rect 2708 7960 2709 8000
rect 2667 7951 2709 7960
rect 2764 8000 2804 8009
rect 2571 7580 2613 7589
rect 2571 7540 2572 7580
rect 2612 7540 2613 7580
rect 2571 7531 2613 7540
rect 2571 7412 2613 7421
rect 2571 7372 2572 7412
rect 2612 7372 2613 7412
rect 2571 7363 2613 7372
rect 2668 7412 2708 7951
rect 2764 7757 2804 7960
rect 2859 7916 2901 7925
rect 2859 7876 2860 7916
rect 2900 7876 2901 7916
rect 2859 7867 2901 7876
rect 2763 7748 2805 7757
rect 2763 7708 2764 7748
rect 2804 7708 2805 7748
rect 2763 7699 2805 7708
rect 2668 7363 2708 7372
rect 2860 7412 2900 7867
rect 2860 7363 2900 7372
rect 2475 7160 2517 7169
rect 2475 7120 2476 7160
rect 2516 7120 2517 7160
rect 2475 7111 2517 7120
rect 2379 6488 2421 6497
rect 2379 6448 2380 6488
rect 2420 6448 2421 6488
rect 2379 6439 2421 6448
rect 2476 6488 2516 7111
rect 2476 6320 2516 6448
rect 2572 6329 2612 7363
rect 2668 6992 2708 7001
rect 2708 6952 2804 6992
rect 2668 6943 2708 6952
rect 2667 6656 2709 6665
rect 2667 6616 2668 6656
rect 2708 6616 2709 6656
rect 2667 6607 2709 6616
rect 2668 6522 2708 6607
rect 2764 6488 2804 6952
rect 2956 6908 2996 8455
rect 3052 7328 3092 8539
rect 3148 7916 3188 9211
rect 3148 7748 3188 7876
rect 3244 7916 3284 9388
rect 3340 9378 3380 9463
rect 3436 9437 3476 9472
rect 3531 9512 3573 9521
rect 3531 9472 3532 9512
rect 3572 9472 3573 9512
rect 3531 9463 3573 9472
rect 4108 9512 4148 9523
rect 3435 9428 3477 9437
rect 3435 9388 3436 9428
rect 3476 9388 3477 9428
rect 3435 9379 3477 9388
rect 3532 8933 3572 9463
rect 4108 9437 4148 9472
rect 4107 9428 4149 9437
rect 4107 9388 4108 9428
rect 4148 9388 4149 9428
rect 4107 9379 4149 9388
rect 3688 9092 4056 9101
rect 3728 9052 3770 9092
rect 3810 9052 3852 9092
rect 3892 9052 3934 9092
rect 3974 9052 4016 9092
rect 3688 9043 4056 9052
rect 3531 8924 3573 8933
rect 3531 8884 3532 8924
rect 3572 8884 3573 8924
rect 3531 8875 3573 8884
rect 3819 8924 3861 8933
rect 3819 8884 3820 8924
rect 3860 8884 3861 8924
rect 3819 8875 3861 8884
rect 3436 8672 3476 8681
rect 3724 8672 3764 8681
rect 3339 8588 3381 8597
rect 3339 8548 3340 8588
rect 3380 8548 3381 8588
rect 3339 8539 3381 8548
rect 3340 8454 3380 8539
rect 3436 8177 3476 8632
rect 3532 8632 3724 8672
rect 3435 8168 3477 8177
rect 3435 8128 3436 8168
rect 3476 8128 3477 8168
rect 3435 8119 3477 8128
rect 3244 7832 3284 7876
rect 3244 7792 3476 7832
rect 3148 7708 3380 7748
rect 3052 7288 3188 7328
rect 3148 7244 3188 7288
rect 3148 7204 3284 7244
rect 3051 7160 3093 7169
rect 3051 7120 3052 7160
rect 3092 7120 3093 7160
rect 3051 7111 3093 7120
rect 3052 7026 3092 7111
rect 2956 6868 3092 6908
rect 2956 6488 2996 6497
rect 2764 6448 2956 6488
rect 2956 6439 2996 6448
rect 3052 6488 3092 6868
rect 3244 6656 3284 7204
rect 3244 6607 3284 6616
rect 3052 6439 3092 6448
rect 3147 6488 3189 6497
rect 3147 6448 3148 6488
rect 3188 6448 3189 6488
rect 3147 6439 3189 6448
rect 3148 6354 3188 6439
rect 2380 6280 2516 6320
rect 2571 6320 2613 6329
rect 2571 6280 2572 6320
rect 2612 6280 2613 6320
rect 2283 5060 2325 5069
rect 2283 5020 2284 5060
rect 2324 5020 2325 5060
rect 2283 5011 2325 5020
rect 2380 4976 2420 6280
rect 2571 6271 2613 6280
rect 3051 6320 3093 6329
rect 3051 6280 3052 6320
rect 3092 6280 3093 6320
rect 3051 6271 3093 6280
rect 3243 6320 3285 6329
rect 3243 6280 3244 6320
rect 3284 6280 3285 6320
rect 3243 6271 3285 6280
rect 2668 5653 2708 5662
rect 2764 5657 2804 5676
rect 2763 5648 2805 5657
rect 2708 5613 2764 5648
rect 2668 5608 2764 5613
rect 2804 5608 2805 5648
rect 2475 5480 2517 5489
rect 2475 5440 2476 5480
rect 2516 5440 2517 5480
rect 2475 5431 2517 5440
rect 2476 5346 2516 5431
rect 2668 5144 2708 5608
rect 2763 5599 2805 5608
rect 2668 5104 2804 5144
rect 2476 4976 2516 4985
rect 2380 4936 2476 4976
rect 2187 4808 2229 4817
rect 2187 4768 2188 4808
rect 2228 4768 2229 4808
rect 2187 4759 2229 4768
rect 2476 4136 2516 4936
rect 2667 4808 2709 4817
rect 2667 4768 2668 4808
rect 2708 4768 2709 4808
rect 2667 4759 2709 4768
rect 2668 4674 2708 4759
rect 2516 4096 2612 4136
rect 2476 4087 2516 4096
rect 2476 3548 2516 3557
rect 2187 3212 2229 3221
rect 2187 3172 2188 3212
rect 2228 3172 2229 3212
rect 2187 3163 2229 3172
rect 2091 1532 2133 1541
rect 2091 1492 2092 1532
rect 2132 1492 2133 1532
rect 2091 1483 2133 1492
rect 1899 272 1941 281
rect 1899 232 1900 272
rect 1940 232 1941 272
rect 1899 223 1941 232
rect 1804 148 1847 188
rect 1807 104 1847 148
rect 1804 80 1847 104
rect 1995 104 2037 113
rect 1995 80 1996 104
rect 1784 0 1864 80
rect 1976 64 1996 80
rect 2036 80 2037 104
rect 2188 80 2228 3163
rect 2283 3128 2325 3137
rect 2283 3088 2284 3128
rect 2324 3088 2325 3128
rect 2283 3079 2325 3088
rect 2284 1028 2324 3079
rect 2380 1196 2420 1205
rect 2476 1196 2516 3508
rect 2572 1952 2612 4096
rect 2667 3968 2709 3977
rect 2667 3928 2668 3968
rect 2708 3928 2709 3968
rect 2667 3919 2709 3928
rect 2668 3834 2708 3919
rect 2668 3450 2708 3459
rect 2668 2885 2708 3410
rect 2667 2876 2709 2885
rect 2667 2836 2668 2876
rect 2708 2836 2709 2876
rect 2667 2827 2709 2836
rect 2764 2120 2804 5104
rect 2860 4985 2900 5066
rect 2854 4976 2900 4985
rect 2854 4936 2855 4976
rect 2854 4927 2900 4936
rect 2955 4976 2997 4985
rect 2955 4936 2956 4976
rect 2996 4936 2997 4976
rect 2955 4927 2997 4936
rect 2859 4808 2901 4817
rect 2859 4768 2860 4808
rect 2900 4768 2901 4808
rect 2859 4759 2901 4768
rect 2860 4136 2900 4759
rect 2860 4087 2900 4096
rect 2956 4136 2996 4927
rect 2859 3968 2901 3977
rect 2859 3928 2860 3968
rect 2900 3928 2901 3968
rect 2859 3919 2901 3928
rect 2764 2071 2804 2080
rect 2572 1903 2612 1912
rect 2420 1156 2516 1196
rect 2380 1147 2420 1156
rect 2764 1112 2804 1121
rect 2860 1112 2900 3919
rect 2956 3893 2996 4096
rect 2955 3884 2997 3893
rect 2955 3844 2956 3884
rect 2996 3844 2997 3884
rect 2955 3835 2997 3844
rect 2955 1868 2997 1877
rect 2955 1828 2956 1868
rect 2996 1828 2997 1868
rect 2955 1819 2997 1828
rect 2956 1734 2996 1819
rect 3052 1280 3092 6271
rect 3147 5816 3189 5825
rect 3147 5776 3148 5816
rect 3188 5776 3189 5816
rect 3147 5767 3189 5776
rect 3148 5648 3188 5767
rect 3148 5599 3188 5608
rect 3147 5480 3189 5489
rect 3147 5440 3148 5480
rect 3188 5440 3189 5480
rect 3147 5431 3189 5440
rect 3148 4817 3188 5431
rect 3147 4808 3189 4817
rect 3147 4768 3148 4808
rect 3188 4768 3189 4808
rect 3147 4759 3189 4768
rect 3148 4388 3188 4397
rect 3244 4388 3284 6271
rect 3340 5909 3380 7708
rect 3436 7673 3476 7792
rect 3435 7664 3477 7673
rect 3435 7624 3436 7664
rect 3476 7624 3477 7664
rect 3435 7615 3477 7624
rect 3435 7160 3477 7169
rect 3435 7120 3436 7160
rect 3476 7120 3477 7160
rect 3435 7111 3477 7120
rect 3436 6581 3476 7111
rect 3532 6665 3572 8632
rect 3724 8623 3764 8632
rect 3820 8504 3860 8875
rect 4204 8765 4244 9640
rect 4492 9185 4532 10144
rect 4588 10184 4628 10732
rect 4683 10732 4684 10772
rect 4724 10732 4725 10772
rect 4683 10723 4725 10732
rect 4588 9521 4628 10144
rect 4587 9512 4629 9521
rect 4587 9472 4588 9512
rect 4628 9472 4629 9512
rect 4587 9463 4629 9472
rect 4683 9428 4725 9437
rect 4683 9388 4684 9428
rect 4724 9388 4725 9428
rect 4683 9379 4725 9388
rect 4491 9176 4533 9185
rect 4491 9136 4492 9176
rect 4532 9136 4533 9176
rect 4491 9127 4533 9136
rect 4492 8840 4532 8849
rect 4684 8840 4724 9379
rect 4300 8800 4492 8840
rect 4203 8756 4245 8765
rect 4203 8716 4204 8756
rect 4244 8716 4245 8756
rect 4203 8707 4245 8716
rect 4300 8683 4340 8800
rect 4492 8791 4532 8800
rect 4588 8800 4724 8840
rect 4780 8840 4820 15511
rect 4876 15401 4916 15688
rect 4875 15392 4917 15401
rect 4875 15352 4876 15392
rect 4916 15352 4917 15392
rect 4875 15343 4917 15352
rect 4928 14384 5296 14393
rect 4968 14344 5010 14384
rect 5050 14344 5092 14384
rect 5132 14344 5174 14384
rect 5214 14344 5256 14384
rect 4928 14335 5296 14344
rect 4928 12872 5296 12881
rect 4968 12832 5010 12872
rect 5050 12832 5092 12872
rect 5132 12832 5174 12872
rect 5214 12832 5256 12872
rect 4928 12823 5296 12832
rect 5356 12620 5396 17032
rect 5451 16316 5493 16325
rect 5451 16276 5452 16316
rect 5492 16276 5493 16316
rect 5451 16267 5493 16276
rect 5452 12881 5492 16267
rect 5548 16241 5588 17200
rect 5740 17072 5780 17081
rect 5836 17072 5876 23248
rect 6123 23239 6165 23248
rect 6604 23213 6644 24592
rect 6699 24583 6741 24592
rect 6699 23372 6741 23381
rect 6699 23332 6700 23372
rect 6740 23332 6741 23372
rect 6699 23323 6741 23332
rect 6315 23204 6357 23213
rect 6315 23164 6316 23204
rect 6356 23164 6357 23204
rect 6315 23155 6357 23164
rect 6603 23204 6645 23213
rect 6603 23164 6604 23204
rect 6644 23164 6645 23204
rect 6603 23155 6645 23164
rect 5932 23120 5972 23131
rect 6124 23120 6164 23129
rect 5932 23045 5972 23080
rect 6028 23080 6124 23120
rect 5931 23036 5973 23045
rect 5931 22996 5932 23036
rect 5972 22996 5973 23036
rect 5931 22987 5973 22996
rect 6028 22877 6068 23080
rect 6124 23071 6164 23080
rect 6316 23120 6356 23155
rect 6316 23069 6356 23080
rect 6604 23120 6644 23155
rect 6604 23070 6644 23080
rect 6700 23120 6740 23323
rect 6700 23071 6740 23080
rect 6315 22952 6357 22961
rect 6315 22912 6316 22952
rect 6356 22912 6357 22952
rect 6315 22903 6357 22912
rect 6027 22868 6069 22877
rect 6027 22828 6028 22868
rect 6068 22828 6069 22868
rect 6027 22819 6069 22828
rect 6220 22868 6260 22877
rect 6220 22373 6260 22828
rect 6219 22364 6261 22373
rect 6219 22324 6220 22364
rect 6260 22324 6261 22364
rect 6219 22315 6261 22324
rect 6219 22196 6261 22205
rect 6219 22156 6220 22196
rect 6260 22156 6261 22196
rect 6219 22147 6261 22156
rect 6123 21356 6165 21365
rect 6123 21316 6124 21356
rect 6164 21316 6165 21356
rect 6123 21307 6165 21316
rect 6124 20768 6164 21307
rect 6124 20719 6164 20728
rect 6220 20768 6260 22147
rect 5931 20684 5973 20693
rect 5931 20644 5932 20684
rect 5972 20644 5973 20684
rect 5931 20635 5973 20644
rect 5932 18500 5972 20635
rect 5932 18257 5972 18460
rect 6028 18500 6068 18509
rect 6028 18341 6068 18460
rect 6027 18332 6069 18341
rect 6027 18292 6028 18332
rect 6068 18292 6069 18332
rect 6027 18283 6069 18292
rect 5931 18248 5973 18257
rect 5931 18208 5932 18248
rect 5972 18208 5973 18248
rect 5931 18199 5973 18208
rect 6027 17912 6069 17921
rect 6027 17872 6028 17912
rect 6068 17872 6069 17912
rect 6027 17863 6069 17872
rect 5780 17032 5876 17072
rect 5547 16232 5589 16241
rect 5547 16192 5548 16232
rect 5588 16192 5589 16232
rect 5547 16183 5589 16192
rect 5740 15644 5780 17032
rect 5548 15604 5780 15644
rect 5548 13889 5588 15604
rect 6028 15560 6068 17863
rect 6220 17660 6260 20728
rect 5739 15476 5781 15485
rect 5739 15436 5740 15476
rect 5780 15436 5781 15476
rect 5739 15427 5781 15436
rect 5643 14888 5685 14897
rect 5643 14848 5644 14888
rect 5684 14848 5685 14888
rect 5643 14839 5685 14848
rect 5644 14720 5684 14839
rect 5644 14671 5684 14680
rect 5740 14645 5780 15427
rect 5739 14636 5781 14645
rect 5739 14596 5740 14636
rect 5780 14596 5781 14636
rect 5739 14587 5781 14596
rect 5547 13880 5589 13889
rect 5547 13840 5548 13880
rect 5588 13840 5589 13880
rect 5547 13831 5589 13840
rect 5643 13208 5685 13217
rect 5643 13168 5644 13208
rect 5684 13168 5685 13208
rect 5643 13159 5685 13168
rect 5644 13074 5684 13159
rect 5451 12872 5493 12881
rect 5451 12832 5452 12872
rect 5492 12832 5493 12872
rect 5451 12823 5493 12832
rect 5260 12580 5396 12620
rect 5164 12536 5204 12545
rect 5164 12293 5204 12496
rect 5163 12284 5205 12293
rect 5163 12244 5164 12284
rect 5204 12244 5205 12284
rect 5163 12235 5205 12244
rect 5260 11528 5300 12580
rect 5644 12536 5684 12545
rect 5356 12496 5644 12536
rect 5356 12284 5396 12496
rect 5644 12487 5684 12496
rect 5740 12536 5780 14587
rect 5836 14552 5876 14561
rect 5836 14048 5876 14512
rect 6028 14309 6068 15520
rect 6124 17620 6260 17660
rect 6027 14300 6069 14309
rect 6027 14260 6028 14300
rect 6068 14260 6069 14300
rect 6027 14251 6069 14260
rect 5932 14048 5972 14057
rect 5836 14008 5932 14048
rect 5932 13999 5972 14008
rect 6027 14048 6069 14057
rect 6027 14008 6028 14048
rect 6068 14008 6069 14048
rect 6027 13999 6069 14008
rect 6028 13914 6068 13999
rect 5835 13880 5877 13889
rect 5835 13840 5836 13880
rect 5876 13840 5877 13880
rect 5835 13831 5877 13840
rect 5356 12235 5396 12244
rect 5451 12032 5493 12041
rect 5451 11992 5452 12032
rect 5492 11992 5493 12032
rect 5451 11983 5493 11992
rect 5452 11696 5492 11983
rect 5452 11647 5492 11656
rect 5260 11488 5396 11528
rect 4928 11360 5296 11369
rect 4968 11320 5010 11360
rect 5050 11320 5092 11360
rect 5132 11320 5174 11360
rect 5214 11320 5256 11360
rect 4928 11311 5296 11320
rect 4971 11192 5013 11201
rect 4971 11152 4972 11192
rect 5012 11152 5013 11192
rect 4971 11143 5013 11152
rect 4972 11058 5012 11143
rect 4875 11024 4917 11033
rect 4875 10984 4876 11024
rect 4916 10984 4917 11024
rect 4875 10975 4917 10984
rect 5068 11024 5108 11033
rect 4876 10890 4916 10975
rect 5068 10865 5108 10984
rect 5163 11024 5205 11033
rect 5163 10984 5164 11024
rect 5204 10984 5205 11024
rect 5163 10975 5205 10984
rect 5164 10890 5204 10975
rect 5067 10856 5109 10865
rect 5067 10816 5068 10856
rect 5108 10816 5109 10856
rect 5067 10807 5109 10816
rect 5356 9857 5396 11488
rect 5740 11360 5780 12496
rect 5836 11873 5876 13831
rect 6124 13796 6164 17620
rect 6219 16148 6261 16157
rect 6219 16108 6220 16148
rect 6260 16108 6261 16148
rect 6219 16099 6261 16108
rect 6220 15653 6260 16099
rect 6219 15644 6261 15653
rect 6219 15604 6220 15644
rect 6260 15604 6261 15644
rect 6219 15595 6261 15604
rect 6220 15560 6260 15595
rect 6220 15509 6260 15520
rect 6220 14720 6260 14729
rect 6220 13889 6260 14680
rect 6219 13880 6261 13889
rect 6219 13840 6220 13880
rect 6260 13840 6261 13880
rect 6219 13831 6261 13840
rect 6028 13756 6164 13796
rect 5931 12536 5973 12545
rect 5931 12496 5932 12536
rect 5972 12496 5973 12536
rect 5931 12487 5973 12496
rect 5835 11864 5877 11873
rect 5835 11824 5836 11864
rect 5876 11824 5877 11864
rect 5835 11815 5877 11824
rect 5932 11789 5972 12487
rect 5931 11780 5973 11789
rect 5931 11740 5932 11780
rect 5972 11740 5973 11780
rect 5931 11731 5973 11740
rect 5932 11360 5972 11731
rect 5644 11320 5780 11360
rect 5836 11320 5972 11360
rect 4928 9848 5296 9857
rect 4968 9808 5010 9848
rect 5050 9808 5092 9848
rect 5132 9808 5174 9848
rect 5214 9808 5256 9848
rect 4928 9799 5296 9808
rect 5355 9848 5397 9857
rect 5355 9808 5356 9848
rect 5396 9808 5397 9848
rect 5355 9799 5397 9808
rect 5356 9605 5396 9636
rect 5355 9596 5397 9605
rect 5355 9556 5356 9596
rect 5396 9556 5397 9596
rect 5355 9547 5397 9556
rect 5547 9596 5589 9605
rect 5547 9556 5548 9596
rect 5588 9556 5589 9596
rect 5547 9547 5589 9556
rect 5356 9512 5396 9547
rect 5356 9185 5396 9472
rect 5548 9462 5588 9547
rect 5355 9176 5397 9185
rect 5355 9136 5356 9176
rect 5396 9136 5397 9176
rect 5355 9127 5397 9136
rect 4780 8800 4916 8840
rect 4012 8672 4052 8683
rect 4012 8597 4052 8632
rect 4107 8672 4149 8681
rect 4107 8632 4108 8672
rect 4148 8632 4149 8672
rect 4300 8634 4340 8643
rect 4491 8672 4533 8681
rect 4107 8623 4149 8632
rect 4491 8632 4492 8672
rect 4532 8632 4533 8672
rect 4491 8623 4533 8632
rect 4011 8588 4053 8597
rect 4011 8548 4012 8588
rect 4052 8548 4053 8588
rect 4011 8539 4053 8548
rect 3724 8464 3860 8504
rect 3724 8000 3764 8464
rect 4108 8084 4148 8623
rect 4492 8538 4532 8623
rect 4203 8504 4245 8513
rect 4203 8464 4204 8504
rect 4244 8464 4245 8504
rect 4203 8455 4245 8464
rect 4204 8370 4244 8455
rect 4395 8168 4437 8177
rect 4395 8128 4396 8168
rect 4436 8128 4437 8168
rect 4395 8119 4437 8128
rect 4108 8044 4244 8084
rect 3724 7841 3764 7960
rect 4204 7986 4244 8044
rect 4396 8034 4436 8119
rect 4204 7925 4244 7946
rect 4203 7916 4245 7925
rect 4203 7876 4204 7916
rect 4244 7876 4245 7916
rect 4203 7867 4245 7876
rect 3723 7832 3765 7841
rect 3723 7792 3724 7832
rect 3764 7792 3765 7832
rect 3723 7783 3765 7792
rect 4107 7748 4149 7757
rect 4107 7708 4108 7748
rect 4148 7708 4149 7748
rect 4107 7699 4149 7708
rect 3688 7580 4056 7589
rect 3728 7540 3770 7580
rect 3810 7540 3852 7580
rect 3892 7540 3934 7580
rect 3974 7540 4016 7580
rect 3688 7531 4056 7540
rect 3531 6656 3573 6665
rect 3531 6616 3532 6656
rect 3572 6616 3573 6656
rect 3531 6607 3573 6616
rect 3435 6572 3477 6581
rect 3435 6532 3436 6572
rect 3476 6532 3477 6572
rect 3435 6523 3477 6532
rect 3436 6488 3476 6523
rect 3436 6438 3476 6448
rect 4108 6245 4148 7699
rect 4395 7496 4437 7505
rect 4395 7456 4396 7496
rect 4436 7456 4437 7496
rect 4395 7447 4437 7456
rect 4299 7244 4341 7253
rect 4299 7204 4300 7244
rect 4340 7204 4341 7244
rect 4299 7195 4341 7204
rect 4300 7160 4340 7195
rect 4300 7109 4340 7120
rect 4107 6236 4149 6245
rect 4107 6196 4108 6236
rect 4148 6196 4149 6236
rect 4107 6187 4149 6196
rect 4299 6236 4341 6245
rect 4299 6196 4300 6236
rect 4340 6196 4341 6236
rect 4299 6187 4341 6196
rect 3688 6068 4056 6077
rect 3728 6028 3770 6068
rect 3810 6028 3852 6068
rect 3892 6028 3934 6068
rect 3974 6028 4016 6068
rect 3688 6019 4056 6028
rect 3339 5900 3381 5909
rect 3339 5860 3340 5900
rect 3380 5860 3381 5900
rect 3339 5851 3381 5860
rect 3723 5900 3765 5909
rect 3723 5860 3724 5900
rect 3764 5860 3765 5900
rect 3723 5851 3765 5860
rect 3627 5732 3669 5741
rect 3627 5692 3628 5732
rect 3668 5692 3669 5732
rect 3627 5683 3669 5692
rect 3724 5732 3764 5851
rect 3724 5683 3764 5692
rect 3628 5598 3668 5683
rect 4108 5648 4148 5659
rect 4108 5573 4148 5608
rect 4204 5648 4244 5657
rect 4107 5564 4149 5573
rect 4107 5524 4108 5564
rect 4148 5524 4149 5564
rect 4107 5515 4149 5524
rect 4204 5069 4244 5608
rect 4300 5153 4340 6187
rect 4396 5405 4436 7447
rect 4588 7421 4628 8800
rect 4780 8672 4820 8681
rect 4683 8000 4725 8009
rect 4683 7960 4684 8000
rect 4724 7960 4725 8000
rect 4683 7951 4725 7960
rect 4684 7866 4724 7951
rect 4780 7589 4820 8632
rect 4876 8513 4916 8800
rect 5355 8672 5397 8681
rect 5355 8632 5356 8672
rect 5396 8632 5397 8672
rect 5355 8623 5397 8632
rect 4875 8504 4917 8513
rect 4875 8464 4876 8504
rect 4916 8464 4917 8504
rect 4875 8455 4917 8464
rect 4928 8336 5296 8345
rect 4968 8296 5010 8336
rect 5050 8296 5092 8336
rect 5132 8296 5174 8336
rect 5214 8296 5256 8336
rect 4928 8287 5296 8296
rect 4779 7580 4821 7589
rect 4779 7540 4780 7580
rect 4820 7540 4821 7580
rect 4779 7531 4821 7540
rect 4587 7412 4629 7421
rect 4587 7372 4588 7412
rect 4628 7372 4629 7412
rect 4587 7363 4629 7372
rect 4492 7160 4532 7169
rect 4492 5816 4532 7120
rect 4588 7160 4628 7169
rect 4588 6329 4628 7120
rect 4684 7160 4724 7169
rect 4684 6740 4724 7120
rect 4779 6992 4821 7001
rect 4779 6952 4780 6992
rect 4820 6952 4821 6992
rect 4779 6943 4821 6952
rect 4780 6858 4820 6943
rect 4928 6824 5296 6833
rect 4968 6784 5010 6824
rect 5050 6784 5092 6824
rect 5132 6784 5174 6824
rect 5214 6784 5256 6824
rect 4928 6775 5296 6784
rect 4684 6700 4826 6740
rect 4786 6572 4826 6700
rect 4780 6532 4826 6572
rect 4684 6446 4724 6455
rect 4587 6320 4629 6329
rect 4587 6280 4588 6320
rect 4628 6280 4629 6320
rect 4587 6271 4629 6280
rect 4684 6245 4724 6406
rect 4683 6236 4725 6245
rect 4683 6196 4684 6236
rect 4724 6196 4725 6236
rect 4683 6187 4725 6196
rect 4780 6152 4820 6532
rect 5164 6488 5204 6497
rect 4876 6448 5164 6488
rect 4876 6320 4916 6448
rect 5164 6439 5204 6448
rect 5260 6488 5300 6499
rect 5260 6413 5300 6448
rect 5259 6404 5301 6413
rect 5259 6364 5260 6404
rect 5300 6364 5301 6404
rect 5259 6355 5301 6364
rect 4876 6271 4916 6280
rect 4780 6112 5012 6152
rect 4972 5900 5012 6112
rect 4972 5851 5012 5860
rect 4492 5776 4820 5816
rect 4780 5657 4820 5776
rect 4588 5653 4628 5657
rect 4492 5648 4628 5653
rect 4492 5613 4588 5648
rect 4395 5396 4437 5405
rect 4395 5356 4396 5396
rect 4436 5356 4437 5396
rect 4395 5347 4437 5356
rect 4299 5144 4341 5153
rect 4299 5104 4300 5144
rect 4340 5104 4341 5144
rect 4299 5095 4341 5104
rect 3339 5060 3381 5069
rect 3339 5020 3340 5060
rect 3380 5020 3381 5060
rect 3339 5011 3381 5020
rect 4203 5060 4245 5069
rect 4203 5020 4204 5060
rect 4244 5020 4245 5060
rect 4203 5011 4245 5020
rect 3188 4348 3284 4388
rect 3148 4339 3188 4348
rect 3243 4220 3285 4229
rect 3243 4180 3244 4220
rect 3284 4180 3285 4220
rect 3243 4171 3285 4180
rect 3147 4136 3189 4145
rect 3147 4096 3148 4136
rect 3188 4096 3189 4136
rect 3147 4087 3189 4096
rect 3148 4002 3188 4087
rect 3147 3632 3189 3641
rect 3147 3592 3148 3632
rect 3188 3592 3189 3632
rect 3147 3583 3189 3592
rect 3148 3464 3188 3583
rect 3148 3415 3188 3424
rect 3244 2624 3284 4171
rect 3340 4136 3380 5011
rect 4108 4976 4148 4985
rect 4108 4817 4148 4936
rect 4300 4892 4340 5095
rect 4492 4985 4532 5613
rect 4588 5599 4628 5608
rect 4684 5648 4724 5657
rect 4684 5405 4724 5608
rect 4779 5648 4821 5657
rect 4779 5608 4780 5648
rect 4820 5608 4821 5648
rect 4779 5599 4821 5608
rect 5163 5648 5205 5657
rect 5163 5608 5164 5648
rect 5204 5608 5205 5648
rect 5163 5599 5205 5608
rect 5164 5514 5204 5599
rect 4683 5396 4725 5405
rect 4683 5356 4684 5396
rect 4724 5356 4725 5396
rect 4683 5347 4725 5356
rect 4491 4976 4533 4985
rect 4491 4936 4492 4976
rect 4532 4936 4533 4976
rect 4491 4927 4533 4936
rect 4204 4852 4340 4892
rect 4395 4892 4437 4901
rect 4395 4852 4396 4892
rect 4436 4852 4437 4892
rect 4107 4808 4149 4817
rect 4107 4768 4108 4808
rect 4148 4768 4149 4808
rect 4107 4759 4149 4768
rect 3688 4556 4056 4565
rect 3728 4516 3770 4556
rect 3810 4516 3852 4556
rect 3892 4516 3934 4556
rect 3974 4516 4016 4556
rect 3688 4507 4056 4516
rect 3531 4304 3573 4313
rect 3531 4264 3532 4304
rect 3572 4264 3573 4304
rect 3531 4255 3573 4264
rect 3340 4087 3380 4096
rect 3435 2876 3477 2885
rect 3435 2836 3436 2876
rect 3476 2836 3477 2876
rect 3435 2827 3477 2836
rect 3436 2742 3476 2827
rect 3244 2575 3284 2584
rect 3532 2540 3572 4255
rect 4108 4229 4148 4759
rect 4107 4220 4149 4229
rect 4107 4180 4108 4220
rect 4148 4180 4149 4220
rect 4107 4171 4149 4180
rect 4204 4052 4244 4852
rect 4395 4843 4437 4852
rect 4108 4012 4244 4052
rect 4300 4724 4340 4733
rect 3627 3464 3669 3473
rect 3627 3424 3628 3464
rect 3668 3424 3669 3464
rect 3627 3415 3669 3424
rect 4108 3464 4148 4012
rect 4108 3415 4148 3424
rect 4204 3464 4244 3473
rect 4300 3464 4340 4684
rect 4244 3424 4340 3464
rect 4204 3415 4244 3424
rect 3628 3330 3668 3415
rect 3723 3380 3765 3389
rect 3723 3340 3724 3380
rect 3764 3340 3765 3380
rect 3723 3331 3765 3340
rect 3724 3246 3764 3331
rect 3688 3044 4056 3053
rect 3728 3004 3770 3044
rect 3810 3004 3852 3044
rect 3892 3004 3934 3044
rect 3974 3004 4016 3044
rect 3688 2995 4056 3004
rect 3915 2708 3957 2717
rect 3820 2668 3916 2708
rect 3956 2668 3957 2708
rect 3820 2624 3860 2668
rect 3915 2659 3957 2668
rect 3820 2575 3860 2584
rect 3436 2500 3572 2540
rect 3147 1700 3189 1709
rect 3147 1660 3148 1700
rect 3188 1660 3189 1700
rect 3147 1651 3189 1660
rect 3340 1700 3380 1711
rect 3148 1566 3188 1651
rect 3340 1625 3380 1660
rect 3339 1616 3381 1625
rect 3339 1576 3340 1616
rect 3380 1576 3381 1616
rect 3339 1567 3381 1576
rect 3436 1448 3476 2500
rect 3532 1952 3572 1961
rect 3532 1793 3572 1912
rect 3531 1784 3573 1793
rect 3531 1744 3532 1784
rect 3572 1744 3573 1784
rect 3531 1735 3573 1744
rect 4107 1784 4149 1793
rect 4107 1744 4108 1784
rect 4148 1744 4149 1784
rect 4107 1735 4149 1744
rect 3688 1532 4056 1541
rect 3728 1492 3770 1532
rect 3810 1492 3852 1532
rect 3892 1492 3934 1532
rect 3974 1492 4016 1532
rect 3688 1483 4056 1492
rect 2804 1072 2900 1112
rect 2956 1240 3092 1280
rect 3148 1408 3476 1448
rect 2764 1063 2804 1072
rect 2284 988 2420 1028
rect 2380 80 2420 988
rect 2572 944 2612 953
rect 2763 944 2805 953
rect 2612 904 2708 944
rect 2572 895 2612 904
rect 2571 776 2613 785
rect 2571 736 2572 776
rect 2612 736 2613 776
rect 2571 727 2613 736
rect 2572 80 2612 727
rect 2668 701 2708 904
rect 2763 904 2764 944
rect 2804 904 2805 944
rect 2763 895 2805 904
rect 2667 692 2709 701
rect 2667 652 2668 692
rect 2708 652 2709 692
rect 2667 643 2709 652
rect 2764 80 2804 895
rect 2956 80 2996 1240
rect 3148 80 3188 1408
rect 3339 1280 3381 1289
rect 3339 1240 3340 1280
rect 3380 1240 3381 1280
rect 3339 1231 3381 1240
rect 3723 1280 3765 1289
rect 3723 1240 3724 1280
rect 3764 1240 3765 1280
rect 3723 1231 3765 1240
rect 3340 80 3380 1231
rect 3531 1028 3573 1037
rect 3531 988 3532 1028
rect 3572 988 3573 1028
rect 3531 979 3573 988
rect 3532 80 3572 979
rect 3724 80 3764 1231
rect 3915 1196 3957 1205
rect 3915 1156 3916 1196
rect 3956 1156 3957 1196
rect 3915 1147 3957 1156
rect 3916 80 3956 1147
rect 4012 1112 4052 1121
rect 4108 1112 4148 1735
rect 4396 1196 4436 4843
rect 4492 4724 4532 4733
rect 4492 4145 4532 4684
rect 4587 4220 4629 4229
rect 4587 4180 4588 4220
rect 4628 4180 4629 4220
rect 4587 4171 4629 4180
rect 4491 4136 4533 4145
rect 4491 4096 4492 4136
rect 4532 4096 4533 4136
rect 4491 4087 4533 4096
rect 4588 4136 4628 4171
rect 4588 4085 4628 4096
rect 4684 3641 4724 5347
rect 4928 5312 5296 5321
rect 4968 5272 5010 5312
rect 5050 5272 5092 5312
rect 5132 5272 5174 5312
rect 5214 5272 5256 5312
rect 4928 5263 5296 5272
rect 4779 5060 4821 5069
rect 4779 5020 4780 5060
rect 4820 5020 4821 5060
rect 4779 5011 4821 5020
rect 4780 4976 4820 5011
rect 4780 4925 4820 4936
rect 5260 4976 5300 4985
rect 5356 4976 5396 8623
rect 5451 8504 5493 8513
rect 5451 8464 5452 8504
rect 5492 8464 5493 8504
rect 5451 8455 5493 8464
rect 5452 6245 5492 8455
rect 5547 8084 5589 8093
rect 5547 8044 5548 8084
rect 5588 8044 5589 8084
rect 5547 8035 5589 8044
rect 5451 6236 5493 6245
rect 5451 6196 5452 6236
rect 5492 6196 5493 6236
rect 5451 6187 5493 6196
rect 5300 4936 5396 4976
rect 5260 4927 5300 4936
rect 5259 4640 5301 4649
rect 5259 4600 5260 4640
rect 5300 4600 5301 4640
rect 5259 4591 5301 4600
rect 4971 4304 5013 4313
rect 4971 4264 4972 4304
rect 5012 4264 5013 4304
rect 4971 4255 5013 4264
rect 4972 4170 5012 4255
rect 4779 4052 4821 4061
rect 4779 4012 4780 4052
rect 4820 4012 4821 4052
rect 4779 4003 4821 4012
rect 4780 3918 4820 4003
rect 5260 3977 5300 4591
rect 5451 4304 5493 4313
rect 5451 4264 5452 4304
rect 5492 4264 5493 4304
rect 5451 4255 5493 4264
rect 5356 4136 5396 4147
rect 5356 4061 5396 4096
rect 5452 4136 5492 4255
rect 5452 4087 5492 4096
rect 5355 4052 5397 4061
rect 5355 4012 5356 4052
rect 5396 4012 5397 4052
rect 5355 4003 5397 4012
rect 5259 3968 5301 3977
rect 5259 3928 5260 3968
rect 5300 3928 5301 3968
rect 5259 3919 5301 3928
rect 5355 3884 5397 3893
rect 5355 3844 5356 3884
rect 5396 3844 5397 3884
rect 5355 3835 5397 3844
rect 4928 3800 5296 3809
rect 4968 3760 5010 3800
rect 5050 3760 5092 3800
rect 5132 3760 5174 3800
rect 5214 3760 5256 3800
rect 4928 3751 5296 3760
rect 5068 3641 5108 3645
rect 4683 3632 4725 3641
rect 4683 3592 4684 3632
rect 4724 3592 4725 3632
rect 4683 3583 4725 3592
rect 5067 3636 5109 3641
rect 5067 3592 5068 3636
rect 5108 3592 5109 3636
rect 5067 3583 5109 3592
rect 4587 3548 4629 3557
rect 4587 3508 4588 3548
rect 4628 3508 4629 3548
rect 4587 3499 4629 3508
rect 5068 3501 5108 3583
rect 4588 3296 4628 3499
rect 4876 3464 4916 3473
rect 4876 3305 4916 3424
rect 4972 3464 5012 3473
rect 4588 3247 4628 3256
rect 4875 3296 4917 3305
rect 4875 3256 4876 3296
rect 4916 3256 4917 3296
rect 4875 3247 4917 3256
rect 4972 2885 5012 3424
rect 5260 3464 5300 3473
rect 5356 3464 5396 3835
rect 5300 3424 5396 3464
rect 5260 3415 5300 3424
rect 5260 2885 5300 2970
rect 4971 2876 5013 2885
rect 4971 2836 4972 2876
rect 5012 2836 5013 2876
rect 4971 2827 5013 2836
rect 5259 2876 5301 2885
rect 5259 2836 5260 2876
rect 5300 2836 5301 2876
rect 5259 2827 5301 2836
rect 5452 2708 5492 2717
rect 5548 2708 5588 8035
rect 5644 7757 5684 11320
rect 5836 11024 5876 11320
rect 5836 10975 5876 10984
rect 5739 9680 5781 9689
rect 5739 9640 5740 9680
rect 5780 9640 5781 9680
rect 5739 9631 5781 9640
rect 5740 9546 5780 9631
rect 5884 9470 5924 9479
rect 5884 9428 5924 9430
rect 5740 9388 5924 9428
rect 5740 8924 5780 9388
rect 5931 9176 5973 9185
rect 5931 9136 5932 9176
rect 5972 9136 5973 9176
rect 5931 9127 5973 9136
rect 5740 8875 5780 8884
rect 5932 8672 5972 9127
rect 5932 8623 5972 8632
rect 6028 8504 6068 13756
rect 6219 12872 6261 12881
rect 6219 12832 6220 12872
rect 6260 12832 6261 12872
rect 6219 12823 6261 12832
rect 6123 12536 6165 12545
rect 6123 12496 6124 12536
rect 6164 12496 6165 12536
rect 6123 12487 6165 12496
rect 6220 12536 6260 12823
rect 6124 12402 6164 12487
rect 6123 12284 6165 12293
rect 6123 12244 6124 12284
rect 6164 12244 6165 12284
rect 6123 12235 6165 12244
rect 5836 8464 6068 8504
rect 5643 7748 5685 7757
rect 5643 7708 5644 7748
rect 5684 7708 5685 7748
rect 5643 7699 5685 7708
rect 5643 6488 5685 6497
rect 5643 6448 5644 6488
rect 5684 6448 5685 6488
rect 5643 6439 5685 6448
rect 5644 6354 5684 6439
rect 5740 6404 5780 6413
rect 5164 2668 5396 2708
rect 5068 2624 5108 2633
rect 5164 2624 5204 2668
rect 5108 2584 5204 2624
rect 5068 2575 5108 2584
rect 4928 2288 5296 2297
rect 4968 2248 5010 2288
rect 5050 2248 5092 2288
rect 5132 2248 5174 2288
rect 5214 2248 5256 2288
rect 4928 2239 5296 2248
rect 4779 2120 4821 2129
rect 4779 2080 4780 2120
rect 4820 2080 4821 2120
rect 4779 2071 4821 2080
rect 4780 1961 4820 2071
rect 4779 1952 4821 1961
rect 4779 1912 4780 1952
rect 4820 1912 4821 1952
rect 4779 1903 4821 1912
rect 4971 1952 5013 1961
rect 4971 1912 4972 1952
rect 5012 1912 5013 1952
rect 4971 1903 5013 1912
rect 4780 1818 4820 1903
rect 4972 1818 5012 1903
rect 5356 1793 5396 2668
rect 5492 2668 5588 2708
rect 5452 2659 5492 2668
rect 5644 2456 5684 2465
rect 5644 2045 5684 2416
rect 5643 2036 5685 2045
rect 5643 1996 5644 2036
rect 5684 1996 5685 2036
rect 5643 1987 5685 1996
rect 5355 1784 5397 1793
rect 5355 1744 5356 1784
rect 5396 1744 5397 1784
rect 5355 1735 5397 1744
rect 4971 1532 5013 1541
rect 4971 1492 4972 1532
rect 5012 1492 5013 1532
rect 4971 1483 5013 1492
rect 4875 1448 4917 1457
rect 4875 1408 4876 1448
rect 4916 1408 4917 1448
rect 4875 1399 4917 1408
rect 4396 1147 4436 1156
rect 4780 1121 4820 1206
rect 4052 1072 4148 1112
rect 4203 1112 4245 1121
rect 4203 1072 4204 1112
rect 4244 1072 4245 1112
rect 4012 1063 4052 1072
rect 4203 1063 4245 1072
rect 4779 1112 4821 1121
rect 4779 1072 4780 1112
rect 4820 1072 4821 1112
rect 4779 1063 4821 1072
rect 4876 1112 4916 1399
rect 4204 1028 4244 1063
rect 4204 977 4244 988
rect 4491 1028 4533 1037
rect 4491 988 4492 1028
rect 4532 988 4533 1028
rect 4491 979 4533 988
rect 4107 944 4149 953
rect 4107 904 4108 944
rect 4148 904 4149 944
rect 4107 895 4149 904
rect 4108 80 4148 895
rect 4299 608 4341 617
rect 4299 568 4300 608
rect 4340 568 4341 608
rect 4299 559 4341 568
rect 4300 80 4340 559
rect 4492 80 4532 979
rect 4587 944 4629 953
rect 4876 944 4916 1072
rect 4972 1112 5012 1483
rect 5451 1280 5493 1289
rect 5451 1240 5452 1280
rect 5492 1240 5493 1280
rect 5451 1231 5493 1240
rect 4972 1063 5012 1072
rect 5067 1112 5109 1121
rect 5067 1072 5068 1112
rect 5108 1072 5109 1112
rect 5067 1063 5109 1072
rect 5356 1112 5396 1121
rect 5068 978 5108 1063
rect 5356 953 5396 1072
rect 4587 904 4588 944
rect 4628 904 4629 944
rect 4587 895 4629 904
rect 4684 904 4916 944
rect 5355 944 5397 953
rect 5355 904 5356 944
rect 5396 904 5397 944
rect 4588 810 4628 895
rect 4684 80 4724 904
rect 5355 895 5397 904
rect 4928 776 5296 785
rect 4968 736 5010 776
rect 5050 736 5092 776
rect 5132 736 5174 776
rect 5214 736 5256 776
rect 4928 727 5296 736
rect 4875 608 4917 617
rect 4875 568 4876 608
rect 4916 568 4917 608
rect 4875 559 4917 568
rect 5259 608 5301 617
rect 5259 568 5260 608
rect 5300 568 5301 608
rect 5259 559 5301 568
rect 4876 80 4916 559
rect 5067 524 5109 533
rect 5067 484 5068 524
rect 5108 484 5109 524
rect 5067 475 5109 484
rect 5068 80 5108 475
rect 5260 80 5300 559
rect 5452 80 5492 1231
rect 5643 1196 5685 1205
rect 5643 1156 5644 1196
rect 5684 1156 5685 1196
rect 5643 1147 5685 1156
rect 5644 1112 5684 1147
rect 5644 1061 5684 1072
rect 5740 1037 5780 6364
rect 5836 6161 5876 8464
rect 6124 8420 6164 12235
rect 6220 8597 6260 12496
rect 6316 11033 6356 22903
rect 6796 20861 6836 25843
rect 6988 25304 7028 25852
rect 7180 25313 7220 26440
rect 7275 26440 7276 26480
rect 7316 26440 7317 26480
rect 7275 26431 7317 26440
rect 7084 25304 7124 25312
rect 6988 25303 7124 25304
rect 6988 25264 7084 25303
rect 7084 25254 7124 25263
rect 7179 25304 7221 25313
rect 7179 25264 7180 25304
rect 7220 25264 7221 25304
rect 7179 25255 7221 25264
rect 7180 25170 7220 25255
rect 7179 24632 7221 24641
rect 7179 24592 7180 24632
rect 7220 24592 7221 24632
rect 7179 24583 7221 24592
rect 7180 24498 7220 24583
rect 6891 23792 6933 23801
rect 6891 23752 6892 23792
rect 6932 23752 6933 23792
rect 6891 23743 6933 23752
rect 7276 23792 7316 26431
rect 7468 24632 7508 27355
rect 7563 27068 7605 27077
rect 7563 27028 7564 27068
rect 7604 27028 7605 27068
rect 7563 27019 7605 27028
rect 7564 26934 7604 27019
rect 7659 26480 7701 26489
rect 7659 26440 7660 26480
rect 7700 26440 7701 26480
rect 7659 26431 7701 26440
rect 7563 25304 7605 25313
rect 7563 25264 7564 25304
rect 7604 25264 7605 25304
rect 7563 25255 7605 25264
rect 7660 25304 7700 26431
rect 7564 25170 7604 25255
rect 7660 25052 7700 25264
rect 7276 23743 7316 23752
rect 7372 24592 7468 24632
rect 6892 23658 6932 23743
rect 7083 23624 7125 23633
rect 7083 23584 7084 23624
rect 7124 23584 7125 23624
rect 7083 23575 7125 23584
rect 7084 23490 7124 23575
rect 6891 23456 6933 23465
rect 6891 23416 6892 23456
rect 6932 23416 6933 23456
rect 6891 23407 6933 23416
rect 6892 22709 6932 23407
rect 6987 23204 7029 23213
rect 6987 23164 6988 23204
rect 7028 23164 7029 23204
rect 6987 23155 7029 23164
rect 6891 22700 6933 22709
rect 6891 22660 6892 22700
rect 6932 22660 6933 22700
rect 6891 22651 6933 22660
rect 6988 22280 7028 23155
rect 7083 23036 7125 23045
rect 7083 22996 7084 23036
rect 7124 22996 7125 23036
rect 7083 22987 7125 22996
rect 7180 23036 7220 23045
rect 7084 22902 7124 22987
rect 7180 22877 7220 22996
rect 7179 22868 7221 22877
rect 7179 22828 7180 22868
rect 7220 22828 7221 22868
rect 7179 22819 7221 22828
rect 7083 22700 7125 22709
rect 7083 22660 7084 22700
rect 7124 22660 7125 22700
rect 7083 22651 7125 22660
rect 6988 22231 7028 22240
rect 7084 22280 7124 22651
rect 7084 22231 7124 22240
rect 7275 22280 7317 22289
rect 7275 22240 7276 22280
rect 7316 22240 7317 22280
rect 7275 22231 7317 22240
rect 7276 22112 7316 22231
rect 7276 22063 7316 22072
rect 6891 21776 6933 21785
rect 6891 21736 6892 21776
rect 6932 21736 6933 21776
rect 6891 21727 6933 21736
rect 7083 21776 7125 21785
rect 7083 21736 7084 21776
rect 7124 21736 7125 21776
rect 7083 21727 7125 21736
rect 6892 21608 6932 21727
rect 7084 21642 7124 21727
rect 6795 20852 6837 20861
rect 6795 20812 6796 20852
rect 6836 20812 6837 20852
rect 6892 20852 6932 21568
rect 7179 20852 7221 20861
rect 6892 20812 7028 20852
rect 6795 20803 6837 20812
rect 6604 20768 6644 20779
rect 6604 20693 6644 20728
rect 6699 20768 6741 20777
rect 6699 20728 6700 20768
rect 6740 20728 6741 20768
rect 6699 20719 6741 20728
rect 6603 20684 6645 20693
rect 6603 20644 6604 20684
rect 6644 20644 6645 20684
rect 6603 20635 6645 20644
rect 6700 20634 6740 20719
rect 6988 20516 7028 20812
rect 7179 20812 7180 20852
rect 7220 20812 7221 20852
rect 7179 20803 7221 20812
rect 6604 20476 7028 20516
rect 7180 20768 7220 20803
rect 6604 20096 6644 20476
rect 6796 20180 6836 20220
rect 6796 20105 6836 20140
rect 6604 20047 6644 20056
rect 6795 20096 6837 20105
rect 6795 20056 6796 20096
rect 6836 20056 6837 20096
rect 6795 20047 6837 20056
rect 6988 20096 7028 20105
rect 6796 20045 6836 20047
rect 6988 19769 7028 20056
rect 6987 19760 7029 19769
rect 6987 19720 6988 19760
rect 7028 19720 7029 19760
rect 6987 19711 7029 19720
rect 6988 19517 7028 19711
rect 6987 19508 7029 19517
rect 6987 19468 6988 19508
rect 7028 19468 7029 19508
rect 6987 19459 7029 19468
rect 6411 19256 6453 19265
rect 6411 19216 6412 19256
rect 6452 19216 6453 19256
rect 6411 19207 6453 19216
rect 6412 17744 6452 19207
rect 7180 18836 7220 20728
rect 7372 20357 7412 24592
rect 7468 24583 7508 24592
rect 7564 25012 7700 25052
rect 7564 24632 7604 25012
rect 7564 24464 7604 24592
rect 7468 24424 7604 24464
rect 7468 22961 7508 24424
rect 7563 23624 7605 23633
rect 7563 23584 7564 23624
rect 7604 23584 7605 23624
rect 7563 23575 7605 23584
rect 7467 22952 7509 22961
rect 7467 22912 7468 22952
rect 7508 22912 7509 22952
rect 7467 22903 7509 22912
rect 7564 22112 7604 23575
rect 7659 23120 7701 23129
rect 7659 23080 7660 23120
rect 7700 23080 7701 23120
rect 7659 23071 7701 23080
rect 7660 22986 7700 23071
rect 7756 22625 7796 28288
rect 7852 26489 7892 29959
rect 8043 29924 8085 29933
rect 8043 29884 8044 29924
rect 8084 29884 8085 29924
rect 8043 29875 8085 29884
rect 7948 29840 7988 29849
rect 7948 28589 7988 29800
rect 7947 28580 7989 28589
rect 7947 28540 7948 28580
rect 7988 28540 7989 28580
rect 7947 28531 7989 28540
rect 8044 27656 8084 29875
rect 8044 27413 8084 27616
rect 8140 27656 8180 30220
rect 8428 30017 8468 31564
rect 8427 30008 8469 30017
rect 8427 29968 8428 30008
rect 8468 29968 8469 30008
rect 8427 29959 8469 29968
rect 8235 29840 8277 29849
rect 8235 29800 8236 29840
rect 8276 29800 8277 29840
rect 8235 29791 8277 29800
rect 8428 29845 8468 29854
rect 8236 29168 8276 29791
rect 8428 29336 8468 29805
rect 8428 29287 8468 29296
rect 8236 29119 8276 29128
rect 8524 29000 8564 34336
rect 8620 33713 8660 36847
rect 8812 36737 8852 36856
rect 8716 36728 8756 36737
rect 8716 36569 8756 36688
rect 8811 36728 8853 36737
rect 8811 36688 8812 36728
rect 8852 36688 8853 36728
rect 8811 36679 8853 36688
rect 8715 36560 8757 36569
rect 8715 36520 8716 36560
rect 8756 36520 8757 36560
rect 8715 36511 8757 36520
rect 8715 36056 8757 36065
rect 8715 36016 8716 36056
rect 8756 36016 8757 36056
rect 8715 36007 8757 36016
rect 8619 33704 8661 33713
rect 8619 33664 8620 33704
rect 8660 33664 8661 33704
rect 8619 33655 8661 33664
rect 8619 32192 8661 32201
rect 8619 32152 8620 32192
rect 8660 32152 8661 32192
rect 8619 32143 8661 32152
rect 8620 32058 8660 32143
rect 8716 31361 8756 36007
rect 8812 34376 8852 36679
rect 8908 36485 8948 36570
rect 8907 36476 8949 36485
rect 8907 36436 8908 36476
rect 8948 36436 8949 36476
rect 8907 36427 8949 36436
rect 9004 36308 9044 37528
rect 9292 37484 9332 37948
rect 9244 37444 9332 37484
rect 9388 37484 9428 38023
rect 9484 37568 9524 42928
rect 9676 40265 9716 42928
rect 9868 41609 9908 42928
rect 10060 41609 10100 42928
rect 9867 41600 9909 41609
rect 9867 41560 9868 41600
rect 9908 41560 9909 41600
rect 9867 41551 9909 41560
rect 10059 41600 10101 41609
rect 10059 41560 10060 41600
rect 10100 41560 10101 41600
rect 10059 41551 10101 41560
rect 9963 41264 10005 41273
rect 9963 41224 9964 41264
rect 10004 41224 10005 41264
rect 9963 41215 10005 41224
rect 9771 40508 9813 40517
rect 9771 40468 9772 40508
rect 9812 40468 9813 40508
rect 9771 40459 9813 40468
rect 9772 40349 9812 40459
rect 9771 40340 9813 40349
rect 9771 40300 9772 40340
rect 9812 40300 9813 40340
rect 9771 40291 9813 40300
rect 9580 40256 9620 40265
rect 9580 39929 9620 40216
rect 9675 40256 9717 40265
rect 9675 40216 9676 40256
rect 9716 40216 9717 40256
rect 9675 40207 9717 40216
rect 9772 40206 9812 40291
rect 9579 39920 9621 39929
rect 9579 39880 9580 39920
rect 9620 39880 9621 39920
rect 9579 39871 9621 39880
rect 9868 39752 9908 39761
rect 9964 39752 10004 41215
rect 10156 41012 10196 41021
rect 10059 40844 10101 40853
rect 10059 40804 10060 40844
rect 10100 40804 10101 40844
rect 10059 40795 10101 40804
rect 9908 39712 10004 39752
rect 9580 38744 9620 38753
rect 9620 38704 9716 38744
rect 9580 38695 9620 38704
rect 9579 38240 9621 38249
rect 9579 38200 9580 38240
rect 9620 38200 9621 38240
rect 9579 38191 9621 38200
rect 9580 38106 9620 38191
rect 9676 37652 9716 38704
rect 9868 37820 9908 39712
rect 10060 39668 10100 40795
rect 10156 40424 10196 40972
rect 10252 40685 10292 42928
rect 10348 41264 10388 41273
rect 10251 40676 10293 40685
rect 10251 40636 10252 40676
rect 10292 40636 10293 40676
rect 10251 40627 10293 40636
rect 10156 40375 10196 40384
rect 10252 40424 10292 40433
rect 10252 40265 10292 40384
rect 10251 40256 10293 40265
rect 10251 40216 10252 40256
rect 10292 40216 10293 40256
rect 10251 40207 10293 40216
rect 10155 40172 10197 40181
rect 10155 40132 10156 40172
rect 10196 40132 10197 40172
rect 10155 40123 10197 40132
rect 10156 39920 10196 40123
rect 10252 39920 10292 39929
rect 10156 39880 10252 39920
rect 10252 39871 10292 39880
rect 10348 39752 10388 41224
rect 10444 40853 10484 42928
rect 10443 40844 10485 40853
rect 10443 40804 10444 40844
rect 10484 40804 10485 40844
rect 10443 40795 10485 40804
rect 10443 40676 10485 40685
rect 10443 40636 10444 40676
rect 10484 40636 10485 40676
rect 10443 40627 10485 40636
rect 10444 40466 10484 40627
rect 10636 40592 10676 42928
rect 10828 42440 10868 42928
rect 10828 42400 10964 42440
rect 10924 40685 10964 42400
rect 10923 40676 10965 40685
rect 10923 40636 10924 40676
rect 10964 40636 10965 40676
rect 10923 40627 10965 40636
rect 10636 40552 10772 40592
rect 10443 40426 10484 40466
rect 10539 40508 10581 40517
rect 10539 40468 10540 40508
rect 10580 40468 10676 40508
rect 10539 40459 10581 40468
rect 10443 40340 10483 40426
rect 10636 40424 10676 40468
rect 10732 40433 10772 40552
rect 10636 40375 10676 40384
rect 10731 40424 10773 40433
rect 10731 40384 10732 40424
rect 10772 40384 10773 40424
rect 10731 40375 10773 40384
rect 10443 40300 10484 40340
rect 10444 39836 10484 40300
rect 10732 40290 10772 40375
rect 11020 40181 11060 42928
rect 11212 40592 11252 42928
rect 11404 41609 11444 42928
rect 11596 41609 11636 42928
rect 11788 42617 11828 42928
rect 11787 42608 11829 42617
rect 11787 42568 11788 42608
rect 11828 42568 11829 42608
rect 11787 42559 11829 42568
rect 11403 41600 11445 41609
rect 11403 41560 11404 41600
rect 11444 41560 11445 41600
rect 11403 41551 11445 41560
rect 11595 41600 11637 41609
rect 11595 41560 11596 41600
rect 11636 41560 11637 41600
rect 11595 41551 11637 41560
rect 11307 41432 11349 41441
rect 11307 41392 11308 41432
rect 11348 41392 11349 41432
rect 11307 41383 11349 41392
rect 11116 40552 11252 40592
rect 11116 40256 11156 40552
rect 11212 40424 11252 40433
rect 11308 40424 11348 41383
rect 11596 41273 11636 41358
rect 11595 41264 11637 41273
rect 11500 41224 11596 41264
rect 11636 41224 11637 41264
rect 11403 41180 11445 41189
rect 11403 41140 11404 41180
rect 11444 41140 11445 41180
rect 11403 41131 11445 41140
rect 11252 40384 11348 40424
rect 11212 40375 11252 40384
rect 11116 40216 11252 40256
rect 10731 40172 10773 40181
rect 10731 40132 10732 40172
rect 10772 40132 10773 40172
rect 10731 40123 10773 40132
rect 11019 40172 11061 40181
rect 11019 40132 11020 40172
rect 11060 40132 11061 40172
rect 11019 40123 11061 40132
rect 10444 39796 10580 39836
rect 10252 39712 10388 39752
rect 10060 39628 10196 39668
rect 10060 39500 10100 39509
rect 9964 39460 10060 39500
rect 9964 38240 10004 39460
rect 10060 39451 10100 39460
rect 10156 38996 10196 39628
rect 10252 39593 10292 39712
rect 10444 39668 10484 39677
rect 10348 39628 10444 39668
rect 10251 39584 10293 39593
rect 10251 39544 10252 39584
rect 10292 39544 10293 39584
rect 10251 39535 10293 39544
rect 10060 38956 10196 38996
rect 10060 38837 10100 38956
rect 10252 38912 10292 38921
rect 10156 38872 10252 38912
rect 10059 38828 10101 38837
rect 10059 38788 10060 38828
rect 10100 38788 10101 38828
rect 10059 38779 10101 38788
rect 9964 38191 10004 38200
rect 10059 38240 10101 38249
rect 10059 38200 10060 38240
rect 10100 38200 10101 38240
rect 10059 38191 10101 38200
rect 10060 38106 10100 38191
rect 9868 37780 10100 37820
rect 9676 37612 10004 37652
rect 9484 37528 9908 37568
rect 9388 37444 9524 37484
rect 9244 37442 9284 37444
rect 9244 37393 9284 37402
rect 9388 37190 9428 37199
rect 9388 37148 9428 37150
rect 9292 37108 9428 37148
rect 8908 36268 9044 36308
rect 9100 36728 9140 36737
rect 8908 35141 8948 36268
rect 9100 35561 9140 36688
rect 9099 35552 9141 35561
rect 9099 35512 9100 35552
rect 9140 35512 9141 35552
rect 9099 35503 9141 35512
rect 9292 35309 9332 37108
rect 9484 37064 9524 37444
rect 9771 37400 9813 37409
rect 9771 37360 9772 37400
rect 9812 37360 9813 37400
rect 9771 37351 9813 37360
rect 9580 37232 9620 37241
rect 9620 37192 9716 37232
rect 9580 37183 9620 37192
rect 9388 37024 9524 37064
rect 9003 35300 9045 35309
rect 9003 35260 9004 35300
rect 9044 35260 9045 35300
rect 9003 35251 9045 35260
rect 9291 35300 9333 35309
rect 9291 35260 9292 35300
rect 9332 35260 9333 35300
rect 9291 35251 9333 35260
rect 9004 35216 9044 35251
rect 8907 35132 8949 35141
rect 8907 35092 8908 35132
rect 8948 35092 8949 35132
rect 8907 35083 8949 35092
rect 8908 34721 8948 35083
rect 9004 35057 9044 35176
rect 9388 35216 9428 37024
rect 9483 36476 9525 36485
rect 9483 36436 9484 36476
rect 9524 36436 9525 36476
rect 9483 36427 9525 36436
rect 9484 35888 9524 36427
rect 9484 35839 9524 35848
rect 9580 35888 9620 35897
rect 9580 35477 9620 35848
rect 9579 35468 9621 35477
rect 9579 35428 9580 35468
rect 9620 35428 9621 35468
rect 9579 35419 9621 35428
rect 9388 35132 9428 35176
rect 9100 35092 9428 35132
rect 9003 35048 9045 35057
rect 9003 35008 9004 35048
rect 9044 35008 9045 35048
rect 9003 34999 9045 35008
rect 8907 34712 8949 34721
rect 8907 34672 8908 34712
rect 8948 34672 8949 34712
rect 8907 34663 8949 34672
rect 9004 34376 9044 34385
rect 8812 34336 9004 34376
rect 9004 34327 9044 34336
rect 8907 34208 8949 34217
rect 8907 34168 8908 34208
rect 8948 34168 8949 34208
rect 8907 34159 8949 34168
rect 8715 31352 8757 31361
rect 8715 31312 8716 31352
rect 8756 31312 8757 31352
rect 8715 31303 8757 31312
rect 8812 31352 8852 31361
rect 8619 31268 8661 31277
rect 8619 31228 8620 31268
rect 8660 31228 8661 31268
rect 8619 31219 8661 31228
rect 8620 29756 8660 31219
rect 8715 31100 8757 31109
rect 8715 31060 8716 31100
rect 8756 31060 8757 31100
rect 8715 31051 8757 31060
rect 8620 29707 8660 29716
rect 8716 29588 8756 31051
rect 8812 30941 8852 31312
rect 8811 30932 8853 30941
rect 8811 30892 8812 30932
rect 8852 30892 8853 30932
rect 8811 30883 8853 30892
rect 8908 30680 8948 34159
rect 8428 28960 8564 29000
rect 8620 29548 8756 29588
rect 8812 29840 8852 29849
rect 8235 28328 8277 28337
rect 8235 28288 8236 28328
rect 8276 28288 8277 28328
rect 8235 28279 8277 28288
rect 8043 27404 8085 27413
rect 8043 27364 8044 27404
rect 8084 27364 8085 27404
rect 8043 27355 8085 27364
rect 7851 26480 7893 26489
rect 8140 26480 8180 27616
rect 7851 26440 7852 26480
rect 7892 26440 7893 26480
rect 7851 26431 7893 26440
rect 7948 26440 8180 26480
rect 7851 25136 7893 25145
rect 7851 25096 7852 25136
rect 7892 25096 7893 25136
rect 7851 25087 7893 25096
rect 7852 24641 7892 25087
rect 7851 24632 7893 24641
rect 7851 24592 7852 24632
rect 7892 24592 7893 24632
rect 7851 24583 7893 24592
rect 7851 24380 7893 24389
rect 7851 24340 7852 24380
rect 7892 24340 7893 24380
rect 7851 24331 7893 24340
rect 7852 24246 7892 24331
rect 7948 24128 7988 26440
rect 8139 25976 8181 25985
rect 8139 25936 8140 25976
rect 8180 25936 8181 25976
rect 8139 25927 8181 25936
rect 8140 25313 8180 25927
rect 8139 25304 8181 25313
rect 8139 25264 8140 25304
rect 8180 25264 8181 25304
rect 8139 25255 8181 25264
rect 8140 25170 8180 25255
rect 8236 24809 8276 28279
rect 8331 26480 8373 26489
rect 8331 26440 8332 26480
rect 8372 26440 8373 26480
rect 8331 26431 8373 26440
rect 8332 26144 8372 26431
rect 8332 26095 8372 26104
rect 8331 25976 8373 25985
rect 8331 25936 8332 25976
rect 8372 25936 8373 25976
rect 8331 25927 8373 25936
rect 8235 24800 8277 24809
rect 8235 24760 8236 24800
rect 8276 24760 8277 24800
rect 8235 24751 8277 24760
rect 8235 24632 8277 24641
rect 8235 24592 8236 24632
rect 8276 24592 8277 24632
rect 8235 24583 8277 24592
rect 8236 24498 8276 24583
rect 7852 24088 7988 24128
rect 7755 22616 7797 22625
rect 7755 22576 7756 22616
rect 7796 22576 7797 22616
rect 7755 22567 7797 22576
rect 7660 22289 7700 22374
rect 7755 22364 7797 22373
rect 7755 22324 7756 22364
rect 7796 22324 7797 22364
rect 7755 22315 7797 22324
rect 7659 22280 7701 22289
rect 7659 22240 7660 22280
rect 7700 22240 7701 22280
rect 7659 22231 7701 22240
rect 7756 22280 7796 22315
rect 7756 22229 7796 22240
rect 7660 22112 7700 22121
rect 7852 22112 7892 24088
rect 8332 23633 8372 25927
rect 8139 23624 8181 23633
rect 8139 23584 8140 23624
rect 8180 23584 8181 23624
rect 8139 23575 8181 23584
rect 8331 23624 8373 23633
rect 8331 23584 8332 23624
rect 8372 23584 8373 23624
rect 8331 23575 8373 23584
rect 8140 23115 8180 23575
rect 8428 23372 8468 28960
rect 8620 27656 8660 29548
rect 8716 29168 8756 29177
rect 8716 28841 8756 29128
rect 8715 28832 8757 28841
rect 8715 28792 8716 28832
rect 8756 28792 8757 28832
rect 8715 28783 8757 28792
rect 8716 27749 8756 28783
rect 8715 27740 8757 27749
rect 8715 27700 8716 27740
rect 8756 27700 8757 27740
rect 8715 27691 8757 27700
rect 8620 26069 8660 27616
rect 8812 26480 8852 29800
rect 8908 28673 8948 30640
rect 9003 29168 9045 29177
rect 9003 29128 9004 29168
rect 9044 29128 9045 29168
rect 9003 29119 9045 29128
rect 8907 28664 8949 28673
rect 8907 28624 8908 28664
rect 8948 28624 8949 28664
rect 8907 28615 8949 28624
rect 8907 28496 8949 28505
rect 8907 28456 8908 28496
rect 8948 28456 8949 28496
rect 8907 28447 8949 28456
rect 8908 26816 8948 28447
rect 9004 28328 9044 29119
rect 9100 28589 9140 35092
rect 9196 34964 9236 34973
rect 9236 34924 9524 34964
rect 9196 34915 9236 34924
rect 9484 34390 9524 34924
rect 9676 34376 9716 37192
rect 9772 36737 9812 37351
rect 9771 36728 9813 36737
rect 9771 36688 9772 36728
rect 9812 36688 9813 36728
rect 9771 36679 9813 36688
rect 9772 36569 9812 36679
rect 9771 36560 9813 36569
rect 9771 36520 9772 36560
rect 9812 36520 9813 36560
rect 9771 36511 9813 36520
rect 9868 35729 9908 37528
rect 9964 36569 10004 37612
rect 10060 37409 10100 37780
rect 10059 37400 10101 37409
rect 10059 37360 10060 37400
rect 10100 37360 10101 37400
rect 10059 37351 10101 37360
rect 10059 37064 10101 37073
rect 10059 37024 10060 37064
rect 10100 37024 10101 37064
rect 10059 37015 10101 37024
rect 9963 36560 10005 36569
rect 9963 36520 9964 36560
rect 10004 36520 10005 36560
rect 9963 36511 10005 36520
rect 10060 36401 10100 37015
rect 10156 36905 10196 38872
rect 10252 38863 10292 38872
rect 10348 37820 10388 39628
rect 10444 39619 10484 39628
rect 10540 38249 10580 39796
rect 10636 39584 10676 39593
rect 10636 39257 10676 39544
rect 10635 39248 10677 39257
rect 10635 39208 10636 39248
rect 10676 39208 10677 39248
rect 10635 39199 10677 39208
rect 10732 39080 10772 40123
rect 10923 39920 10965 39929
rect 10923 39880 10924 39920
rect 10964 39880 10965 39920
rect 10923 39871 10965 39880
rect 10924 39747 10964 39871
rect 11020 39752 11060 39761
rect 10924 39712 11020 39747
rect 10924 39707 11060 39712
rect 11020 39703 11060 39707
rect 11116 39752 11156 39761
rect 11019 39164 11061 39173
rect 11019 39124 11020 39164
rect 11060 39124 11061 39164
rect 11019 39115 11061 39124
rect 10636 39040 10772 39080
rect 10827 39080 10869 39089
rect 10827 39040 10828 39080
rect 10868 39040 10869 39080
rect 10539 38240 10581 38249
rect 10539 38200 10540 38240
rect 10580 38200 10581 38240
rect 10539 38191 10581 38200
rect 10443 38156 10485 38165
rect 10443 38116 10444 38156
rect 10484 38116 10485 38156
rect 10443 38107 10485 38116
rect 10444 38022 10484 38107
rect 10540 38106 10580 38191
rect 10252 37780 10388 37820
rect 10155 36896 10197 36905
rect 10155 36856 10156 36896
rect 10196 36856 10197 36896
rect 10155 36847 10197 36856
rect 10059 36392 10101 36401
rect 10059 36352 10060 36392
rect 10100 36352 10101 36392
rect 10059 36343 10101 36352
rect 9963 35888 10005 35897
rect 9963 35848 9964 35888
rect 10004 35848 10005 35888
rect 9963 35839 10005 35848
rect 10060 35888 10100 35897
rect 9964 35754 10004 35839
rect 10060 35729 10100 35848
rect 9867 35720 9909 35729
rect 9867 35680 9868 35720
rect 9908 35680 9909 35720
rect 9867 35671 9909 35680
rect 10059 35720 10101 35729
rect 10059 35680 10060 35720
rect 10100 35680 10101 35720
rect 10059 35671 10101 35680
rect 9484 34341 9524 34350
rect 9580 34336 9716 34376
rect 9483 34124 9525 34133
rect 9483 34084 9484 34124
rect 9524 34084 9525 34124
rect 9483 34075 9525 34084
rect 9484 33704 9524 34075
rect 9580 33881 9620 34336
rect 9675 34208 9717 34217
rect 9675 34168 9676 34208
rect 9716 34168 9717 34208
rect 9675 34159 9717 34168
rect 9676 34074 9716 34159
rect 9579 33872 9621 33881
rect 9579 33832 9580 33872
rect 9620 33832 9621 33872
rect 9579 33823 9621 33832
rect 9676 33788 9716 33797
rect 9716 33748 10004 33788
rect 9676 33739 9716 33748
rect 9964 33704 10004 33748
rect 9524 33664 9620 33704
rect 9484 33655 9524 33664
rect 9291 32864 9333 32873
rect 9291 32824 9292 32864
rect 9332 32824 9333 32864
rect 9291 32815 9333 32824
rect 9292 32730 9332 32815
rect 9484 32696 9524 32705
rect 9195 32192 9237 32201
rect 9195 32152 9196 32192
rect 9236 32152 9237 32192
rect 9195 32143 9237 32152
rect 9099 28580 9141 28589
rect 9099 28540 9100 28580
rect 9140 28540 9141 28580
rect 9099 28531 9141 28540
rect 9196 28505 9236 32143
rect 9340 31361 9380 31370
rect 9484 31361 9524 32656
rect 9380 31321 9524 31361
rect 9340 31312 9380 31321
rect 9483 31184 9525 31193
rect 9483 31144 9484 31184
rect 9524 31144 9525 31184
rect 9483 31135 9525 31144
rect 9484 31050 9524 31135
rect 9580 29177 9620 33664
rect 9964 33655 10004 33664
rect 10060 33704 10100 33713
rect 10060 33209 10100 33664
rect 10156 33461 10196 36847
rect 10155 33452 10197 33461
rect 10155 33412 10156 33452
rect 10196 33412 10197 33452
rect 10155 33403 10197 33412
rect 10252 33293 10292 37780
rect 10443 36812 10485 36821
rect 10443 36772 10444 36812
rect 10484 36772 10485 36812
rect 10443 36763 10485 36772
rect 10347 36728 10389 36737
rect 10347 36688 10348 36728
rect 10388 36688 10389 36728
rect 10347 36679 10389 36688
rect 10348 36594 10388 36679
rect 10444 36476 10484 36763
rect 10348 36436 10484 36476
rect 10539 36476 10581 36485
rect 10539 36436 10540 36476
rect 10580 36436 10581 36476
rect 10348 34805 10388 36436
rect 10539 36427 10581 36436
rect 10540 36342 10580 36427
rect 10540 35888 10580 35897
rect 10636 35888 10676 39040
rect 10827 39031 10869 39040
rect 10731 38240 10773 38249
rect 10731 38200 10732 38240
rect 10772 38200 10773 38240
rect 10731 38191 10773 38200
rect 10732 37997 10772 38191
rect 10731 37988 10773 37997
rect 10731 37948 10732 37988
rect 10772 37948 10773 37988
rect 10731 37939 10773 37948
rect 10731 37736 10773 37745
rect 10731 37696 10732 37736
rect 10772 37696 10773 37736
rect 10731 37687 10773 37696
rect 10732 36728 10772 37687
rect 10828 37073 10868 39031
rect 11020 38240 11060 39115
rect 11020 38191 11060 38200
rect 11116 37577 11156 39712
rect 11115 37568 11157 37577
rect 11115 37528 11116 37568
rect 11156 37528 11157 37568
rect 11115 37519 11157 37528
rect 11020 37400 11060 37409
rect 11060 37360 11156 37400
rect 11020 37351 11060 37360
rect 10827 37064 10869 37073
rect 10827 37024 10828 37064
rect 10868 37024 10869 37064
rect 10827 37015 10869 37024
rect 11019 36980 11061 36989
rect 11019 36940 11020 36980
rect 11060 36940 11061 36980
rect 11019 36931 11061 36940
rect 10732 36679 10772 36688
rect 11020 36644 11060 36931
rect 10924 36604 11060 36644
rect 10731 36560 10773 36569
rect 10731 36520 10732 36560
rect 10772 36520 10773 36560
rect 10731 36511 10773 36520
rect 10580 35848 10676 35888
rect 10540 35839 10580 35848
rect 10635 35216 10677 35225
rect 10635 35176 10636 35216
rect 10676 35176 10677 35216
rect 10635 35167 10677 35176
rect 10347 34796 10389 34805
rect 10347 34756 10348 34796
rect 10388 34756 10389 34796
rect 10347 34747 10389 34756
rect 10251 33284 10293 33293
rect 10251 33244 10252 33284
rect 10292 33244 10293 33284
rect 10251 33235 10293 33244
rect 10059 33200 10101 33209
rect 10059 33160 10060 33200
rect 10100 33160 10101 33200
rect 10059 33151 10101 33160
rect 9771 32948 9813 32957
rect 9771 32908 9772 32948
rect 9812 32908 9813 32948
rect 9771 32899 9813 32908
rect 9772 29840 9812 32899
rect 9867 32864 9909 32873
rect 9867 32824 9868 32864
rect 9908 32824 9909 32864
rect 9867 32815 9909 32824
rect 10155 32864 10197 32873
rect 10348 32864 10388 34747
rect 10636 34133 10676 35167
rect 10732 35132 10772 36511
rect 10924 35216 10964 36604
rect 11019 36476 11061 36485
rect 11019 36436 11020 36476
rect 11060 36436 11061 36476
rect 11019 36427 11061 36436
rect 11020 35902 11060 36427
rect 11020 35853 11060 35862
rect 11020 35216 11060 35225
rect 10924 35176 11020 35216
rect 11020 35167 11060 35176
rect 10732 35092 10964 35132
rect 10827 34964 10869 34973
rect 10827 34924 10828 34964
rect 10868 34924 10869 34964
rect 10827 34915 10869 34924
rect 10828 34830 10868 34915
rect 10635 34124 10677 34133
rect 10635 34084 10636 34124
rect 10676 34084 10677 34124
rect 10635 34075 10677 34084
rect 10443 33704 10485 33713
rect 10443 33664 10444 33704
rect 10484 33664 10485 33704
rect 10443 33655 10485 33664
rect 10540 33704 10580 33713
rect 10924 33704 10964 35092
rect 11116 34553 11156 37360
rect 11212 36560 11252 40216
rect 11404 38669 11444 41131
rect 11500 39836 11540 41224
rect 11595 41215 11637 41224
rect 11980 41189 12020 42928
rect 12172 41441 12212 42928
rect 12171 41432 12213 41441
rect 12171 41392 12172 41432
rect 12212 41392 12213 41432
rect 12171 41383 12213 41392
rect 12171 41264 12213 41273
rect 12171 41224 12172 41264
rect 12212 41224 12213 41264
rect 12171 41215 12213 41224
rect 11979 41180 12021 41189
rect 11979 41140 11980 41180
rect 12020 41140 12021 41180
rect 11979 41131 12021 41140
rect 12172 41130 12212 41215
rect 11595 41096 11637 41105
rect 11595 41056 11596 41096
rect 11636 41056 11637 41096
rect 11595 41047 11637 41056
rect 11596 40349 11636 41047
rect 11788 41012 11828 41021
rect 11980 41012 12020 41021
rect 11788 40508 11828 40972
rect 11740 40468 11828 40508
rect 11884 40972 11980 41012
rect 11740 40466 11780 40468
rect 11740 40417 11780 40426
rect 11595 40340 11637 40349
rect 11884 40340 11924 40972
rect 11980 40963 12020 40972
rect 12364 40844 12404 42928
rect 12459 41348 12501 41357
rect 12459 41308 12460 41348
rect 12500 41308 12501 41348
rect 12459 41299 12501 41308
rect 11595 40300 11596 40340
rect 11636 40300 11637 40340
rect 11595 40291 11637 40300
rect 11788 40300 11924 40340
rect 11980 40804 12404 40844
rect 11788 40013 11828 40300
rect 11884 40214 11924 40223
rect 11787 40004 11829 40013
rect 11787 39964 11788 40004
rect 11828 39964 11829 40004
rect 11787 39955 11829 39964
rect 11500 39796 11732 39836
rect 11500 39668 11540 39677
rect 11500 39257 11540 39628
rect 11595 39668 11637 39677
rect 11595 39628 11596 39668
rect 11636 39628 11637 39668
rect 11595 39619 11637 39628
rect 11596 39534 11636 39619
rect 11499 39248 11541 39257
rect 11499 39208 11500 39248
rect 11540 39208 11541 39248
rect 11499 39199 11541 39208
rect 11500 38912 11540 38921
rect 11692 38912 11732 39796
rect 11540 38872 11732 38912
rect 11500 38863 11540 38872
rect 11692 38744 11732 38753
rect 11596 38704 11692 38744
rect 11403 38660 11445 38669
rect 11403 38620 11404 38660
rect 11444 38620 11445 38660
rect 11403 38611 11445 38620
rect 11596 38240 11636 38704
rect 11692 38695 11732 38704
rect 11548 38230 11636 38240
rect 11588 38200 11636 38230
rect 11692 38324 11732 38333
rect 11548 38181 11588 38190
rect 11403 38156 11445 38165
rect 11308 38116 11404 38156
rect 11444 38116 11445 38156
rect 11308 36821 11348 38116
rect 11403 38107 11445 38116
rect 11500 37400 11540 37409
rect 11404 37360 11500 37400
rect 11307 36812 11349 36821
rect 11307 36772 11308 36812
rect 11348 36772 11349 36812
rect 11307 36763 11349 36772
rect 11212 36520 11348 36560
rect 11212 35720 11252 35729
rect 11115 34544 11157 34553
rect 11115 34504 11116 34544
rect 11156 34504 11157 34544
rect 11115 34495 11157 34504
rect 11020 34376 11060 34385
rect 11060 34336 11156 34376
rect 11020 34327 11060 34336
rect 11019 34208 11061 34217
rect 11019 34168 11020 34208
rect 11060 34168 11061 34208
rect 11019 34159 11061 34168
rect 11020 33713 11060 34159
rect 11116 33797 11156 34336
rect 11115 33788 11157 33797
rect 11115 33748 11116 33788
rect 11156 33748 11157 33788
rect 11115 33739 11157 33748
rect 10580 33664 10964 33704
rect 10540 33655 10580 33664
rect 10444 33570 10484 33655
rect 10443 33452 10485 33461
rect 10443 33412 10444 33452
rect 10484 33412 10485 33452
rect 10443 33403 10485 33412
rect 10155 32824 10156 32864
rect 10196 32824 10388 32864
rect 10155 32815 10197 32824
rect 9868 32192 9908 32815
rect 10156 32730 10196 32815
rect 9868 31445 9908 32152
rect 10060 31940 10100 31949
rect 9867 31436 9909 31445
rect 9867 31396 9868 31436
rect 9908 31396 9909 31436
rect 9867 31387 9909 31396
rect 9868 30680 9908 31387
rect 10060 31352 10100 31900
rect 10060 31303 10100 31312
rect 10156 31352 10196 31361
rect 10196 31312 10292 31352
rect 10156 31303 10196 31312
rect 10156 30680 10196 30689
rect 9868 30640 10156 30680
rect 10060 29849 10100 30640
rect 10156 30631 10196 30640
rect 9772 29791 9812 29800
rect 10059 29840 10101 29849
rect 10059 29800 10060 29840
rect 10100 29800 10101 29840
rect 10059 29791 10101 29800
rect 9579 29168 9621 29177
rect 9579 29128 9580 29168
rect 9620 29128 9621 29168
rect 9579 29119 9621 29128
rect 9963 29168 10005 29177
rect 9963 29128 9964 29168
rect 10004 29128 10005 29168
rect 9963 29119 10005 29128
rect 9964 29034 10004 29119
rect 10156 28916 10196 28925
rect 9483 28664 9525 28673
rect 9483 28624 9484 28664
rect 9524 28624 9525 28664
rect 9483 28615 9525 28624
rect 9387 28580 9429 28589
rect 9387 28540 9388 28580
rect 9428 28540 9429 28580
rect 9387 28531 9429 28540
rect 9195 28496 9237 28505
rect 9195 28456 9196 28496
rect 9236 28456 9237 28496
rect 9195 28447 9237 28456
rect 9004 28279 9044 28288
rect 9196 28160 9236 28169
rect 9196 27656 9236 28120
rect 9291 28076 9333 28085
rect 9291 28036 9292 28076
rect 9332 28036 9333 28076
rect 9291 28027 9333 28036
rect 9292 27740 9332 28027
rect 9292 27691 9332 27700
rect 9148 27646 9236 27656
rect 9188 27616 9236 27646
rect 9148 27597 9188 27606
rect 9291 27572 9333 27581
rect 9291 27532 9292 27572
rect 9332 27532 9333 27572
rect 9291 27523 9333 27532
rect 9195 27404 9237 27413
rect 9195 27364 9196 27404
rect 9236 27364 9237 27404
rect 9195 27355 9237 27364
rect 9099 26984 9141 26993
rect 9099 26944 9100 26984
rect 9140 26944 9141 26984
rect 9099 26935 9141 26944
rect 8948 26776 9044 26816
rect 8908 26767 8948 26776
rect 8812 26440 8948 26480
rect 8619 26060 8661 26069
rect 8619 26020 8620 26060
rect 8660 26020 8661 26060
rect 8619 26011 8661 26020
rect 8524 25892 8564 25901
rect 8715 25892 8757 25901
rect 8564 25852 8660 25892
rect 8524 25843 8564 25852
rect 8620 25318 8660 25852
rect 8715 25852 8716 25892
rect 8756 25852 8757 25892
rect 8715 25843 8757 25852
rect 8716 25649 8756 25843
rect 8715 25640 8757 25649
rect 8715 25600 8716 25640
rect 8756 25600 8757 25640
rect 8715 25591 8757 25600
rect 8811 25556 8853 25565
rect 8811 25516 8812 25556
rect 8852 25516 8853 25556
rect 8811 25507 8853 25516
rect 8620 25269 8660 25278
rect 8812 25220 8852 25507
rect 8812 25171 8852 25180
rect 8908 23885 8948 26440
rect 9004 26321 9044 26776
rect 9003 26312 9045 26321
rect 9003 26272 9004 26312
rect 9044 26272 9045 26312
rect 9003 26263 9045 26272
rect 9100 25304 9140 26935
rect 9196 26144 9236 27355
rect 9196 26095 9236 26104
rect 8907 23876 8949 23885
rect 8907 23836 8908 23876
rect 8948 23836 8949 23876
rect 8907 23827 8949 23836
rect 8524 23792 8564 23803
rect 8524 23717 8564 23752
rect 9003 23792 9045 23801
rect 9003 23752 9004 23792
rect 9044 23752 9045 23792
rect 9003 23743 9045 23752
rect 8523 23708 8565 23717
rect 8523 23668 8524 23708
rect 8564 23668 8565 23708
rect 8523 23659 8565 23668
rect 9004 23658 9044 23743
rect 8715 23624 8757 23633
rect 8715 23584 8716 23624
rect 8756 23584 8757 23624
rect 8715 23575 8757 23584
rect 8716 23490 8756 23575
rect 8140 23045 8180 23075
rect 8236 23332 8468 23372
rect 8139 23036 8181 23045
rect 8139 22996 8140 23036
rect 8180 22996 8181 23036
rect 8139 22987 8181 22996
rect 8140 22951 8180 22987
rect 7947 22616 7989 22625
rect 7947 22576 7948 22616
rect 7988 22576 7989 22616
rect 7947 22567 7989 22576
rect 7948 22532 7988 22567
rect 7948 22481 7988 22492
rect 8139 22448 8181 22457
rect 8139 22408 8140 22448
rect 8180 22408 8181 22448
rect 8236 22448 8276 23332
rect 8619 23288 8661 23297
rect 9004 23288 9044 23297
rect 8619 23248 8620 23288
rect 8660 23248 8661 23288
rect 8619 23239 8661 23248
rect 8716 23248 9004 23288
rect 8331 23204 8373 23213
rect 8331 23164 8332 23204
rect 8372 23164 8373 23204
rect 8331 23155 8373 23164
rect 8332 23070 8372 23155
rect 8524 23120 8564 23129
rect 8428 23080 8524 23120
rect 8428 22709 8468 23080
rect 8524 23071 8564 23080
rect 8620 23120 8660 23239
rect 8620 23071 8660 23080
rect 8716 23120 8756 23248
rect 9004 23239 9044 23248
rect 8716 23071 8756 23080
rect 8811 23120 8853 23129
rect 9100 23120 9140 25264
rect 9292 23792 9332 27523
rect 9388 23876 9428 28531
rect 9484 26993 9524 28615
rect 10156 28347 10196 28876
rect 10252 28505 10292 31312
rect 10444 31025 10484 33403
rect 10635 33368 10677 33377
rect 10635 33328 10636 33368
rect 10676 33328 10677 33368
rect 10635 33319 10677 33328
rect 10636 31436 10676 33319
rect 10827 32696 10869 32705
rect 10827 32656 10828 32696
rect 10868 32656 10869 32696
rect 10827 32647 10869 32656
rect 10732 32192 10772 32201
rect 10732 31613 10772 32152
rect 10731 31604 10773 31613
rect 10731 31564 10732 31604
rect 10772 31564 10773 31604
rect 10731 31555 10773 31564
rect 10539 31352 10581 31361
rect 10539 31312 10540 31352
rect 10580 31312 10581 31352
rect 10539 31303 10581 31312
rect 10540 31218 10580 31303
rect 10443 31016 10485 31025
rect 10443 30976 10444 31016
rect 10484 30976 10485 31016
rect 10443 30967 10485 30976
rect 10348 30428 10388 30437
rect 10348 29840 10388 30388
rect 10444 30017 10484 30967
rect 10443 30008 10485 30017
rect 10443 29968 10444 30008
rect 10484 29968 10485 30008
rect 10443 29959 10485 29968
rect 10444 29840 10484 29849
rect 10348 29800 10444 29840
rect 10444 29791 10484 29800
rect 10540 29840 10580 29849
rect 10347 29336 10389 29345
rect 10347 29296 10348 29336
rect 10388 29296 10389 29336
rect 10347 29287 10389 29296
rect 10348 29168 10388 29287
rect 10348 29093 10388 29128
rect 10347 29084 10389 29093
rect 10347 29044 10348 29084
rect 10388 29044 10389 29084
rect 10347 29035 10389 29044
rect 10348 29004 10388 29035
rect 10251 28496 10293 28505
rect 10251 28456 10252 28496
rect 10292 28456 10293 28496
rect 10251 28447 10293 28456
rect 10156 28298 10196 28307
rect 10252 28328 10292 28337
rect 9867 27740 9909 27749
rect 9867 27700 9868 27740
rect 9908 27700 9909 27740
rect 9867 27691 9909 27700
rect 9483 26984 9525 26993
rect 9483 26944 9484 26984
rect 9524 26944 9525 26984
rect 9483 26935 9525 26944
rect 9483 26732 9525 26741
rect 9483 26692 9484 26732
rect 9524 26692 9525 26732
rect 9483 26683 9525 26692
rect 9484 26573 9524 26683
rect 9483 26564 9525 26573
rect 9483 26524 9484 26564
rect 9524 26524 9525 26564
rect 9483 26515 9525 26524
rect 9484 24632 9524 26515
rect 9675 24716 9717 24725
rect 9675 24676 9676 24716
rect 9716 24676 9717 24716
rect 9675 24667 9717 24676
rect 9484 24583 9524 24592
rect 9676 24582 9716 24667
rect 9579 24380 9621 24389
rect 9579 24340 9580 24380
rect 9620 24340 9621 24380
rect 9579 24331 9621 24340
rect 9388 23836 9524 23876
rect 9292 23752 9428 23792
rect 9291 23624 9333 23633
rect 9291 23584 9292 23624
rect 9332 23584 9333 23624
rect 9291 23575 9333 23584
rect 9195 23204 9237 23213
rect 9195 23164 9196 23204
rect 9236 23164 9237 23204
rect 9195 23155 9237 23164
rect 8811 23080 8812 23120
rect 8852 23080 8853 23120
rect 8811 23071 8853 23080
rect 8908 23080 9140 23120
rect 9196 23120 9236 23155
rect 9292 23129 9332 23575
rect 8812 22986 8852 23071
rect 8908 22868 8948 23080
rect 9196 23069 9236 23080
rect 9291 23120 9333 23129
rect 9291 23080 9292 23120
rect 9332 23080 9333 23120
rect 9291 23071 9333 23080
rect 9292 22986 9332 23071
rect 8716 22828 8948 22868
rect 8523 22784 8565 22793
rect 8523 22744 8524 22784
rect 8564 22744 8565 22784
rect 8523 22735 8565 22744
rect 8427 22700 8469 22709
rect 8427 22660 8428 22700
rect 8468 22660 8469 22700
rect 8427 22651 8469 22660
rect 8427 22532 8469 22541
rect 8427 22492 8428 22532
rect 8468 22492 8469 22532
rect 8427 22483 8469 22492
rect 8236 22408 8372 22448
rect 8139 22399 8181 22408
rect 7564 22072 7660 22112
rect 7660 22063 7700 22072
rect 7756 22072 7892 22112
rect 7467 21776 7509 21785
rect 7467 21736 7468 21776
rect 7508 21736 7509 21776
rect 7467 21727 7509 21736
rect 7468 21608 7508 21727
rect 7468 21559 7508 21568
rect 7564 21608 7604 21617
rect 7756 21608 7796 22072
rect 7948 21617 7988 21702
rect 7604 21568 7796 21608
rect 7564 21559 7604 21568
rect 7563 21440 7605 21449
rect 7563 21400 7564 21440
rect 7604 21400 7605 21440
rect 7563 21391 7605 21400
rect 7371 20348 7413 20357
rect 7371 20308 7372 20348
rect 7412 20308 7413 20348
rect 7371 20299 7413 20308
rect 7275 19760 7317 19769
rect 7275 19720 7276 19760
rect 7316 19720 7317 19760
rect 7275 19711 7317 19720
rect 7276 19256 7316 19711
rect 7276 19207 7316 19216
rect 6892 18796 7220 18836
rect 6508 18584 6548 18593
rect 6892 18584 6932 18796
rect 6548 18544 6932 18584
rect 7180 18668 7220 18677
rect 6988 18570 7028 18579
rect 6508 18535 6548 18544
rect 6508 17753 6548 17838
rect 6507 17744 6549 17753
rect 6412 17704 6508 17744
rect 6548 17704 6549 17744
rect 6507 17695 6549 17704
rect 6508 16232 6548 16241
rect 6508 15989 6548 16192
rect 6507 15980 6549 15989
rect 6507 15940 6508 15980
rect 6548 15940 6549 15980
rect 6507 15931 6549 15940
rect 6508 15569 6548 15931
rect 6507 15560 6549 15569
rect 6507 15520 6508 15560
rect 6548 15520 6549 15560
rect 6507 15511 6549 15520
rect 6411 14804 6453 14813
rect 6411 14764 6412 14804
rect 6452 14764 6453 14804
rect 6411 14755 6453 14764
rect 6412 14048 6452 14755
rect 6507 14132 6549 14141
rect 6507 14092 6508 14132
rect 6548 14092 6549 14132
rect 6507 14083 6549 14092
rect 6412 12545 6452 14008
rect 6508 14048 6548 14083
rect 6508 13997 6548 14008
rect 6604 13805 6644 18544
rect 6988 18080 7028 18530
rect 7180 18089 7220 18628
rect 7468 18584 7508 18593
rect 7564 18584 7604 21391
rect 7660 20773 7700 20782
rect 7660 20189 7700 20733
rect 7659 20180 7701 20189
rect 7659 20140 7660 20180
rect 7700 20140 7701 20180
rect 7659 20131 7701 20140
rect 7756 20021 7796 21568
rect 7947 21608 7989 21617
rect 7947 21568 7948 21608
rect 7988 21568 7989 21608
rect 7947 21559 7989 21568
rect 8044 21608 8084 21617
rect 8044 21365 8084 21568
rect 8043 21356 8085 21365
rect 8043 21316 8044 21356
rect 8084 21316 8085 21356
rect 8043 21307 8085 21316
rect 8140 20861 8180 22399
rect 8236 22280 8276 22289
rect 8139 20852 8181 20861
rect 8139 20812 8140 20852
rect 8180 20812 8181 20852
rect 8139 20803 8181 20812
rect 8043 20768 8085 20777
rect 8043 20728 8044 20768
rect 8084 20728 8085 20768
rect 8043 20719 8085 20728
rect 8044 20634 8084 20719
rect 8139 20684 8181 20693
rect 8139 20644 8140 20684
rect 8180 20644 8181 20684
rect 8139 20635 8181 20644
rect 7852 20600 7892 20609
rect 7755 20012 7797 20021
rect 7755 19972 7756 20012
rect 7796 19972 7797 20012
rect 7755 19963 7797 19972
rect 7852 19349 7892 20560
rect 8043 20516 8085 20525
rect 8043 20476 8044 20516
rect 8084 20476 8085 20516
rect 8043 20467 8085 20476
rect 7851 19340 7893 19349
rect 7851 19300 7852 19340
rect 7892 19300 7893 19340
rect 7851 19291 7893 19300
rect 7508 18544 7700 18584
rect 7468 18535 7508 18544
rect 7372 18332 7412 18341
rect 6700 18040 7028 18080
rect 7179 18080 7221 18089
rect 7179 18040 7180 18080
rect 7220 18040 7221 18080
rect 6700 17996 6740 18040
rect 7179 18031 7221 18040
rect 6700 17947 6740 17956
rect 7275 17828 7317 17837
rect 7275 17788 7276 17828
rect 7316 17788 7317 17828
rect 7275 17779 7317 17788
rect 6987 17744 7029 17753
rect 6987 17704 6988 17744
rect 7028 17704 7029 17744
rect 6987 17695 7029 17704
rect 7180 17744 7220 17753
rect 6988 17072 7028 17695
rect 7180 17240 7220 17704
rect 7276 17744 7316 17779
rect 7276 17693 7316 17704
rect 7372 17240 7412 18292
rect 7467 18248 7509 18257
rect 7467 18208 7468 18248
rect 7508 18208 7509 18248
rect 7467 18199 7509 18208
rect 7468 17324 7508 18199
rect 7660 17828 7700 18544
rect 7755 18500 7797 18509
rect 7755 18460 7756 18500
rect 7796 18460 7797 18500
rect 7755 18451 7797 18460
rect 7660 17779 7700 17788
rect 7756 17744 7796 18451
rect 7756 17669 7796 17704
rect 7755 17660 7797 17669
rect 7755 17620 7756 17660
rect 7796 17620 7797 17660
rect 7755 17611 7797 17620
rect 7947 17660 7989 17669
rect 7947 17620 7948 17660
rect 7988 17620 7989 17660
rect 7947 17611 7989 17620
rect 7468 17284 7604 17324
rect 7180 17191 7220 17200
rect 7276 17200 7412 17240
rect 6988 17023 7028 17032
rect 6795 16988 6837 16997
rect 6795 16948 6796 16988
rect 6836 16948 6837 16988
rect 6795 16939 6837 16948
rect 6699 16400 6741 16409
rect 6699 16360 6700 16400
rect 6740 16360 6741 16400
rect 6699 16351 6741 16360
rect 6700 16266 6740 16351
rect 6699 16064 6741 16073
rect 6699 16024 6700 16064
rect 6740 16024 6741 16064
rect 6699 16015 6741 16024
rect 6603 13796 6645 13805
rect 6603 13756 6604 13796
rect 6644 13756 6645 13796
rect 6603 13747 6645 13756
rect 6603 13628 6645 13637
rect 6603 13588 6604 13628
rect 6644 13588 6645 13628
rect 6603 13579 6645 13588
rect 6507 13292 6549 13301
rect 6507 13252 6508 13292
rect 6548 13252 6549 13292
rect 6507 13243 6549 13252
rect 6411 12536 6453 12545
rect 6411 12496 6412 12536
rect 6452 12496 6453 12536
rect 6411 12487 6453 12496
rect 6315 11024 6357 11033
rect 6315 10984 6316 11024
rect 6356 10984 6357 11024
rect 6315 10975 6357 10984
rect 6412 9512 6452 9521
rect 6412 8765 6452 9472
rect 6411 8756 6453 8765
rect 6411 8716 6412 8756
rect 6452 8716 6453 8756
rect 6411 8707 6453 8716
rect 6219 8588 6261 8597
rect 6219 8548 6220 8588
rect 6260 8548 6261 8588
rect 6219 8539 6261 8548
rect 5932 8380 6164 8420
rect 5932 8000 5972 8380
rect 6508 8177 6548 13243
rect 6604 9101 6644 13579
rect 6700 12536 6740 16015
rect 6796 15065 6836 16939
rect 6892 16232 6932 16241
rect 6892 15737 6932 16192
rect 6988 16232 7028 16241
rect 6988 15821 7028 16192
rect 7179 16232 7221 16241
rect 7179 16192 7180 16232
rect 7220 16192 7221 16232
rect 7179 16183 7221 16192
rect 7276 16232 7316 17200
rect 7468 17030 7508 17039
rect 7371 16988 7413 16997
rect 7468 16988 7508 16990
rect 7371 16948 7372 16988
rect 7412 16948 7508 16988
rect 7371 16939 7413 16948
rect 7564 16904 7604 17284
rect 7468 16864 7604 16904
rect 7376 16400 7418 16409
rect 7376 16360 7377 16400
rect 7417 16360 7418 16400
rect 7376 16351 7418 16360
rect 7276 16183 7316 16192
rect 7377 16232 7417 16351
rect 7377 16183 7417 16192
rect 7180 16098 7220 16183
rect 7083 16064 7125 16073
rect 7468 16064 7508 16864
rect 7851 16232 7893 16241
rect 7851 16192 7852 16232
rect 7892 16192 7893 16232
rect 7851 16183 7893 16192
rect 7852 16098 7892 16183
rect 7083 16024 7084 16064
rect 7124 16024 7125 16064
rect 7083 16015 7125 16024
rect 7372 16024 7508 16064
rect 7084 15930 7124 16015
rect 6987 15812 7029 15821
rect 6987 15772 6988 15812
rect 7028 15772 7029 15812
rect 6987 15763 7029 15772
rect 6891 15728 6933 15737
rect 6891 15688 6892 15728
rect 6932 15688 6933 15728
rect 6891 15679 6933 15688
rect 6795 15056 6837 15065
rect 6795 15016 6796 15056
rect 6836 15016 6837 15056
rect 6795 15007 6837 15016
rect 6700 12487 6740 12496
rect 6699 12284 6741 12293
rect 6699 12244 6700 12284
rect 6740 12244 6741 12284
rect 6699 12235 6741 12244
rect 6700 11696 6740 12235
rect 6700 11647 6740 11656
rect 6796 11360 6836 15007
rect 6891 14888 6933 14897
rect 6891 14848 6892 14888
rect 6932 14848 6933 14888
rect 6891 14839 6933 14848
rect 6892 13208 6932 14839
rect 6987 14048 7029 14057
rect 6987 14008 6988 14048
rect 7028 14008 7029 14048
rect 6987 13999 7029 14008
rect 6988 13914 7028 13999
rect 7083 13460 7125 13469
rect 7083 13420 7084 13460
rect 7124 13420 7125 13460
rect 7083 13411 7125 13420
rect 7084 13326 7124 13411
rect 6892 12293 6932 13168
rect 7276 13208 7316 13217
rect 7372 13208 7412 16024
rect 7948 15737 7988 17611
rect 8044 17585 8084 20467
rect 8043 17576 8085 17585
rect 8043 17536 8044 17576
rect 8084 17536 8085 17576
rect 8043 17527 8085 17536
rect 8044 17081 8084 17527
rect 8043 17072 8085 17081
rect 8043 17032 8044 17072
rect 8084 17032 8085 17072
rect 8043 17023 8085 17032
rect 8043 16400 8085 16409
rect 8043 16360 8044 16400
rect 8084 16360 8085 16400
rect 8043 16351 8085 16360
rect 7947 15728 7989 15737
rect 7947 15688 7948 15728
rect 7988 15688 7989 15728
rect 7947 15679 7989 15688
rect 7467 15560 7509 15569
rect 7948 15560 7988 15569
rect 7467 15520 7468 15560
rect 7508 15520 7509 15560
rect 7467 15511 7509 15520
rect 7756 15520 7948 15560
rect 7468 14897 7508 15511
rect 7660 15308 7700 15317
rect 7564 15268 7660 15308
rect 7467 14888 7509 14897
rect 7467 14848 7468 14888
rect 7508 14848 7509 14888
rect 7467 14839 7509 14848
rect 7468 14720 7508 14839
rect 7468 14671 7508 14680
rect 7564 14057 7604 15268
rect 7660 15259 7700 15268
rect 7660 14972 7700 14981
rect 7756 14972 7796 15520
rect 7948 15511 7988 15520
rect 8044 15560 8084 16351
rect 8044 15511 8084 15520
rect 7700 14932 8084 14972
rect 7660 14923 7700 14932
rect 8044 14720 8084 14932
rect 8140 14888 8180 20635
rect 8236 20525 8276 22240
rect 8332 21449 8372 22408
rect 8331 21440 8373 21449
rect 8331 21400 8332 21440
rect 8372 21400 8373 21440
rect 8331 21391 8373 21400
rect 8235 20516 8277 20525
rect 8235 20476 8236 20516
rect 8276 20476 8277 20516
rect 8235 20467 8277 20476
rect 8428 20180 8468 22483
rect 8524 21617 8564 22735
rect 8619 21944 8661 21953
rect 8619 21904 8620 21944
rect 8660 21904 8661 21944
rect 8619 21895 8661 21904
rect 8523 21608 8565 21617
rect 8523 21568 8524 21608
rect 8564 21568 8565 21608
rect 8523 21559 8565 21568
rect 8620 21365 8660 21895
rect 8619 21356 8661 21365
rect 8619 21316 8620 21356
rect 8660 21316 8661 21356
rect 8619 21307 8661 21316
rect 8716 20693 8756 22828
rect 9195 22364 9237 22373
rect 9195 22324 9196 22364
rect 9236 22324 9237 22364
rect 9195 22315 9237 22324
rect 9196 21953 9236 22315
rect 9291 22280 9333 22289
rect 9291 22240 9292 22280
rect 9332 22240 9333 22280
rect 9291 22231 9333 22240
rect 9195 21944 9237 21953
rect 9100 21904 9196 21944
rect 9236 21904 9237 21944
rect 9004 21594 9044 21603
rect 9004 21029 9044 21554
rect 9003 21020 9045 21029
rect 9003 20980 9004 21020
rect 9044 20980 9045 21020
rect 9003 20971 9045 20980
rect 8715 20684 8757 20693
rect 8715 20644 8716 20684
rect 8756 20644 8757 20684
rect 8715 20635 8757 20644
rect 8332 20140 8468 20180
rect 8235 20096 8277 20105
rect 8332 20096 8372 20140
rect 8235 20056 8236 20096
rect 8276 20056 8277 20096
rect 8235 20047 8277 20056
rect 8324 20056 8372 20096
rect 8619 20096 8661 20105
rect 8619 20056 8620 20096
rect 8660 20056 8661 20096
rect 8236 19962 8276 20047
rect 8324 20012 8364 20056
rect 8619 20047 8661 20056
rect 8716 20096 8756 20105
rect 8324 19972 8372 20012
rect 8235 18584 8277 18593
rect 8235 18544 8236 18584
rect 8276 18544 8277 18584
rect 8235 18535 8277 18544
rect 8236 18450 8276 18535
rect 8235 17996 8277 18005
rect 8235 17956 8236 17996
rect 8276 17956 8277 17996
rect 8235 17947 8277 17956
rect 8236 17744 8276 17947
rect 8236 15476 8276 17704
rect 8332 15560 8372 19972
rect 8427 19928 8469 19937
rect 8427 19888 8428 19928
rect 8468 19888 8469 19928
rect 8427 19879 8469 19888
rect 8428 19794 8468 19879
rect 8620 19265 8660 20047
rect 8716 19937 8756 20056
rect 8812 20096 8852 20105
rect 8715 19928 8757 19937
rect 8715 19888 8716 19928
rect 8756 19888 8757 19928
rect 8715 19879 8757 19888
rect 8524 19256 8564 19265
rect 8619 19256 8661 19265
rect 8564 19216 8620 19256
rect 8660 19216 8661 19256
rect 8524 19207 8564 19216
rect 8619 19207 8661 19216
rect 8523 19088 8565 19097
rect 8523 19048 8524 19088
rect 8564 19048 8565 19088
rect 8523 19039 8565 19048
rect 8427 18584 8469 18593
rect 8427 18544 8428 18584
rect 8468 18544 8469 18584
rect 8427 18535 8469 18544
rect 8428 15737 8468 18535
rect 8524 17165 8564 19039
rect 8523 17156 8565 17165
rect 8523 17116 8524 17156
rect 8564 17116 8565 17156
rect 8523 17107 8565 17116
rect 8524 16829 8564 17107
rect 8620 17072 8660 19207
rect 8716 19088 8756 19097
rect 8716 17921 8756 19048
rect 8812 18929 8852 20056
rect 8907 20096 8949 20105
rect 9100 20096 9140 21904
rect 9195 21895 9237 21904
rect 9292 21869 9332 22231
rect 9388 21953 9428 23752
rect 9484 23465 9524 23836
rect 9483 23456 9525 23465
rect 9483 23416 9484 23456
rect 9524 23416 9525 23456
rect 9483 23407 9525 23416
rect 9484 23120 9524 23131
rect 9484 23045 9524 23080
rect 9580 23120 9620 24331
rect 9771 23288 9813 23297
rect 9771 23248 9772 23288
rect 9812 23248 9813 23288
rect 9771 23239 9813 23248
rect 9772 23154 9812 23239
rect 9580 23071 9620 23080
rect 9675 23120 9717 23129
rect 9675 23080 9676 23120
rect 9716 23080 9717 23120
rect 9675 23071 9717 23080
rect 9483 23036 9525 23045
rect 9483 22996 9484 23036
rect 9524 22996 9525 23036
rect 9483 22987 9525 22996
rect 9676 22986 9716 23071
rect 9579 22952 9621 22961
rect 9579 22912 9580 22952
rect 9620 22912 9621 22952
rect 9579 22903 9621 22912
rect 9483 22280 9525 22289
rect 9483 22240 9484 22280
rect 9524 22240 9525 22280
rect 9483 22231 9525 22240
rect 9484 22146 9524 22231
rect 9387 21944 9429 21953
rect 9387 21904 9388 21944
rect 9428 21904 9429 21944
rect 9387 21895 9429 21904
rect 9291 21860 9333 21869
rect 9291 21820 9292 21860
rect 9332 21820 9333 21860
rect 9291 21811 9333 21820
rect 9195 21776 9237 21785
rect 9195 21736 9196 21776
rect 9236 21736 9237 21776
rect 9195 21727 9237 21736
rect 9196 21642 9236 21727
rect 9292 20768 9332 21811
rect 9292 20719 9332 20728
rect 9196 20096 9236 20105
rect 8907 20056 8908 20096
rect 8948 20056 8949 20096
rect 8907 20047 8949 20056
rect 9004 20056 9196 20096
rect 8908 19685 8948 20047
rect 8907 19676 8949 19685
rect 8907 19636 8908 19676
rect 8948 19636 8949 19676
rect 8907 19627 8949 19636
rect 8908 19256 8948 19627
rect 8908 19207 8948 19216
rect 8811 18920 8853 18929
rect 8811 18880 8812 18920
rect 8852 18880 8853 18920
rect 8811 18871 8853 18880
rect 8715 17912 8757 17921
rect 8715 17872 8716 17912
rect 8756 17872 8757 17912
rect 8715 17863 8757 17872
rect 8764 17753 8804 17762
rect 8804 17713 8852 17744
rect 8764 17704 8852 17713
rect 8812 17240 8852 17704
rect 8908 17576 8948 17585
rect 8908 17417 8948 17536
rect 8907 17408 8949 17417
rect 8907 17368 8908 17408
rect 8948 17368 8949 17408
rect 8907 17359 8949 17368
rect 8908 17240 8948 17249
rect 8812 17200 8908 17240
rect 8908 17191 8948 17200
rect 8716 17072 8756 17081
rect 8620 17032 8716 17072
rect 8716 17023 8756 17032
rect 8523 16820 8565 16829
rect 8523 16780 8524 16820
rect 8564 16780 8565 16820
rect 8523 16771 8565 16780
rect 8523 16316 8565 16325
rect 8523 16276 8524 16316
rect 8564 16276 8565 16316
rect 8523 16267 8565 16276
rect 8524 16073 8564 16267
rect 8523 16064 8565 16073
rect 8523 16024 8524 16064
rect 8564 16024 8565 16064
rect 8523 16015 8565 16024
rect 8427 15728 8469 15737
rect 8427 15688 8428 15728
rect 8468 15688 8469 15728
rect 8427 15679 8469 15688
rect 8428 15560 8468 15569
rect 8332 15520 8428 15560
rect 8236 15436 8372 15476
rect 8140 14848 8276 14888
rect 8044 14671 8084 14680
rect 8140 14720 8180 14731
rect 8140 14645 8180 14680
rect 8139 14636 8181 14645
rect 8139 14596 8140 14636
rect 8180 14596 8181 14636
rect 8139 14587 8181 14596
rect 8236 14216 8276 14848
rect 8044 14176 8276 14216
rect 7660 14132 7700 14141
rect 7700 14092 7892 14132
rect 7660 14083 7700 14092
rect 7563 14048 7605 14057
rect 7468 14034 7508 14043
rect 7563 14008 7564 14048
rect 7604 14008 7605 14048
rect 7563 13999 7605 14008
rect 7468 13469 7508 13994
rect 7755 13796 7797 13805
rect 7755 13756 7756 13796
rect 7796 13756 7797 13796
rect 7755 13747 7797 13756
rect 7563 13712 7605 13721
rect 7563 13672 7564 13712
rect 7604 13672 7605 13712
rect 7563 13663 7605 13672
rect 7467 13460 7509 13469
rect 7467 13420 7468 13460
rect 7508 13420 7509 13460
rect 7467 13411 7509 13420
rect 7316 13168 7412 13208
rect 7276 13159 7316 13168
rect 7275 13040 7317 13049
rect 7275 13000 7276 13040
rect 7316 13000 7317 13040
rect 7275 12991 7317 13000
rect 7180 12522 7220 12531
rect 6891 12284 6933 12293
rect 6891 12244 6892 12284
rect 6932 12244 6933 12284
rect 6891 12235 6933 12244
rect 6892 11948 6932 11957
rect 7180 11948 7220 12482
rect 6932 11908 7220 11948
rect 6892 11899 6932 11908
rect 7084 11696 7124 11705
rect 7084 11537 7124 11656
rect 7083 11528 7125 11537
rect 7083 11488 7084 11528
rect 7124 11488 7125 11528
rect 7083 11479 7125 11488
rect 7276 11360 7316 12991
rect 6700 11320 6836 11360
rect 6892 11320 7316 11360
rect 7372 12620 7412 12629
rect 6603 9092 6645 9101
rect 6603 9052 6604 9092
rect 6644 9052 6645 9092
rect 6603 9043 6645 9052
rect 6507 8168 6549 8177
rect 6507 8128 6508 8168
rect 6548 8128 6549 8168
rect 6507 8119 6549 8128
rect 5932 7085 5972 7960
rect 6412 8000 6452 8009
rect 6412 7841 6452 7960
rect 6508 8000 6548 8009
rect 6123 7832 6165 7841
rect 6123 7792 6124 7832
rect 6164 7792 6165 7832
rect 6123 7783 6165 7792
rect 6411 7832 6453 7841
rect 6411 7792 6412 7832
rect 6452 7792 6453 7832
rect 6411 7783 6453 7792
rect 6124 7698 6164 7783
rect 6508 7757 6548 7960
rect 6700 7916 6740 11320
rect 6892 9596 6932 11320
rect 7275 11192 7317 11201
rect 7275 11152 7276 11192
rect 7316 11152 7317 11192
rect 7275 11143 7317 11152
rect 7276 11058 7316 11143
rect 7083 11024 7125 11033
rect 7083 10984 7084 11024
rect 7124 10984 7125 11024
rect 7083 10975 7125 10984
rect 7084 10890 7124 10975
rect 7083 10772 7125 10781
rect 7083 10732 7084 10772
rect 7124 10732 7125 10772
rect 7083 10723 7125 10732
rect 6987 9848 7029 9857
rect 6987 9808 6988 9848
rect 7028 9808 7029 9848
rect 6987 9799 7029 9808
rect 6604 7876 6740 7916
rect 6796 9556 6932 9596
rect 6507 7748 6549 7757
rect 6507 7708 6508 7748
rect 6548 7708 6549 7748
rect 6507 7699 6549 7708
rect 6508 7589 6548 7699
rect 6507 7580 6549 7589
rect 6507 7540 6508 7580
rect 6548 7540 6549 7580
rect 6507 7531 6549 7540
rect 6411 7496 6453 7505
rect 6411 7456 6412 7496
rect 6452 7456 6453 7496
rect 6411 7447 6453 7456
rect 6412 7160 6452 7447
rect 6412 7111 6452 7120
rect 5931 7076 5973 7085
rect 5931 7036 5932 7076
rect 5972 7036 5973 7076
rect 5931 7027 5973 7036
rect 6219 6824 6261 6833
rect 6219 6784 6220 6824
rect 6260 6784 6261 6824
rect 6219 6775 6261 6784
rect 5931 6488 5973 6497
rect 5931 6448 5932 6488
rect 5972 6448 5973 6488
rect 5931 6439 5973 6448
rect 6220 6488 6260 6775
rect 6220 6439 6260 6448
rect 5835 6152 5877 6161
rect 5835 6112 5836 6152
rect 5876 6112 5877 6152
rect 5835 6103 5877 6112
rect 5932 5405 5972 6439
rect 6604 6329 6644 7876
rect 6700 6474 6740 6483
rect 6603 6320 6645 6329
rect 6603 6280 6604 6320
rect 6644 6280 6645 6320
rect 6603 6271 6645 6280
rect 6315 6236 6357 6245
rect 6315 6196 6316 6236
rect 6356 6196 6357 6236
rect 6315 6187 6357 6196
rect 6316 5648 6356 6187
rect 6604 5900 6644 5909
rect 6700 5900 6740 6434
rect 6644 5860 6740 5900
rect 6604 5851 6644 5860
rect 6412 5648 6452 5657
rect 6316 5608 6412 5648
rect 5931 5396 5973 5405
rect 5931 5356 5932 5396
rect 5972 5356 5973 5396
rect 5931 5347 5973 5356
rect 6315 5396 6357 5405
rect 6315 5356 6316 5396
rect 6356 5356 6357 5396
rect 6315 5347 6357 5356
rect 5835 4220 5877 4229
rect 5835 4180 5836 4220
rect 5876 4180 5877 4220
rect 5835 4171 5877 4180
rect 5836 4086 5876 4171
rect 5932 4136 5972 4145
rect 5836 2792 5876 2801
rect 5836 2633 5876 2752
rect 5835 2624 5877 2633
rect 5835 2584 5836 2624
rect 5876 2584 5877 2624
rect 5835 2575 5877 2584
rect 5932 1457 5972 4096
rect 6123 3800 6165 3809
rect 6123 3760 6124 3800
rect 6164 3760 6165 3800
rect 6123 3751 6165 3760
rect 6124 2624 6164 3751
rect 6219 3464 6261 3473
rect 6219 3424 6220 3464
rect 6260 3424 6261 3464
rect 6219 3415 6261 3424
rect 6220 3221 6260 3415
rect 6316 3296 6356 5347
rect 6412 4640 6452 5608
rect 6796 5405 6836 9556
rect 6988 9521 7028 9799
rect 6987 9512 7029 9521
rect 6987 9472 6988 9512
rect 7028 9472 7029 9512
rect 6987 9463 7029 9472
rect 6892 9428 6932 9437
rect 6892 9269 6932 9388
rect 6988 9378 7028 9463
rect 6891 9260 6933 9269
rect 6891 9220 6892 9260
rect 6932 9220 6933 9260
rect 6891 9211 6933 9220
rect 6988 8000 7028 8009
rect 7084 8000 7124 10723
rect 7372 9680 7412 12580
rect 7467 12536 7509 12545
rect 7467 12496 7468 12536
rect 7508 12496 7509 12536
rect 7467 12487 7509 12496
rect 7468 10184 7508 12487
rect 7564 10361 7604 13663
rect 7659 12620 7701 12629
rect 7659 12580 7660 12620
rect 7700 12580 7701 12620
rect 7659 12571 7701 12580
rect 7660 12368 7700 12571
rect 7660 12319 7700 12328
rect 7756 12116 7796 13747
rect 7852 12629 7892 14092
rect 8044 13721 8084 14176
rect 8332 14132 8372 15436
rect 8236 14092 8372 14132
rect 8236 13880 8276 14092
rect 8428 14048 8468 15520
rect 8524 15560 8564 16015
rect 8524 15511 8564 15520
rect 9004 15560 9044 20056
rect 9196 20047 9236 20056
rect 9291 20012 9333 20021
rect 9291 19972 9292 20012
rect 9332 19972 9333 20012
rect 9291 19963 9333 19972
rect 9292 19878 9332 19963
rect 9195 19844 9237 19853
rect 9195 19804 9196 19844
rect 9236 19804 9237 19844
rect 9195 19795 9237 19804
rect 9099 18920 9141 18929
rect 9099 18880 9100 18920
rect 9140 18880 9141 18920
rect 9099 18871 9141 18880
rect 9100 17669 9140 18871
rect 9196 18173 9236 19795
rect 9291 18584 9333 18593
rect 9291 18544 9292 18584
rect 9332 18544 9333 18584
rect 9291 18535 9333 18544
rect 9195 18164 9237 18173
rect 9195 18124 9196 18164
rect 9236 18124 9237 18164
rect 9195 18115 9237 18124
rect 9195 17912 9237 17921
rect 9195 17872 9196 17912
rect 9236 17872 9237 17912
rect 9292 17912 9332 18535
rect 9388 18332 9428 21895
rect 9483 21020 9525 21029
rect 9483 20980 9484 21020
rect 9524 20980 9525 21020
rect 9483 20971 9525 20980
rect 9484 20886 9524 20971
rect 9483 19256 9525 19265
rect 9483 19216 9484 19256
rect 9524 19216 9525 19256
rect 9483 19207 9525 19216
rect 9484 18584 9524 19207
rect 9484 18535 9524 18544
rect 9388 18292 9524 18332
rect 9292 17872 9428 17912
rect 9195 17863 9237 17872
rect 9196 17744 9236 17863
rect 9196 17695 9236 17704
rect 9291 17744 9333 17753
rect 9291 17704 9292 17744
rect 9332 17704 9333 17744
rect 9291 17695 9333 17704
rect 9099 17660 9141 17669
rect 9099 17620 9100 17660
rect 9140 17620 9141 17660
rect 9099 17611 9141 17620
rect 9292 17610 9332 17695
rect 9099 17156 9141 17165
rect 9099 17116 9100 17156
rect 9140 17116 9141 17156
rect 9099 17107 9141 17116
rect 9100 16232 9140 17107
rect 9195 17072 9237 17081
rect 9195 17032 9196 17072
rect 9236 17032 9237 17072
rect 9195 17023 9237 17032
rect 9100 15569 9140 16192
rect 8619 15392 8661 15401
rect 8619 15352 8620 15392
rect 8660 15352 8661 15392
rect 8619 15343 8661 15352
rect 8620 14813 8660 15343
rect 8907 15140 8949 15149
rect 8907 15100 8908 15140
rect 8948 15100 8949 15140
rect 8907 15091 8949 15100
rect 8619 14804 8661 14813
rect 8619 14764 8620 14804
rect 8660 14764 8661 14804
rect 8619 14755 8661 14764
rect 8524 14720 8564 14729
rect 8524 14216 8564 14680
rect 8620 14670 8660 14755
rect 8811 14216 8853 14225
rect 8524 14176 8812 14216
rect 8852 14176 8853 14216
rect 8811 14167 8853 14176
rect 8140 13840 8276 13880
rect 8332 14008 8428 14048
rect 8043 13712 8085 13721
rect 8043 13672 8044 13712
rect 8084 13672 8085 13712
rect 8043 13663 8085 13672
rect 7851 12620 7893 12629
rect 7851 12580 7852 12620
rect 7892 12580 7893 12620
rect 7851 12571 7893 12580
rect 7947 12536 7989 12545
rect 7947 12496 7948 12536
rect 7988 12496 7989 12536
rect 7947 12487 7989 12496
rect 8044 12536 8084 12545
rect 7948 12402 7988 12487
rect 7660 12076 7796 12116
rect 7563 10352 7605 10361
rect 7563 10312 7564 10352
rect 7604 10312 7605 10352
rect 7563 10303 7605 10312
rect 7468 10135 7508 10144
rect 7563 10184 7605 10193
rect 7563 10144 7564 10184
rect 7604 10144 7605 10184
rect 7563 10135 7605 10144
rect 7660 10184 7700 12076
rect 8044 11360 8084 12496
rect 7756 11320 8084 11360
rect 7756 11192 7796 11320
rect 7756 11143 7796 11152
rect 7947 11024 7989 11033
rect 7947 10979 7948 11024
rect 7988 10979 7989 11024
rect 7947 10975 7989 10979
rect 7948 10889 7988 10975
rect 8140 10604 8180 13840
rect 8332 13049 8372 14008
rect 8428 13999 8468 14008
rect 8524 14048 8564 14057
rect 8716 14048 8756 14057
rect 8524 13553 8564 14008
rect 8620 14008 8716 14048
rect 8620 13637 8660 14008
rect 8716 13999 8756 14008
rect 8908 13880 8948 15091
rect 9004 14132 9044 15520
rect 9099 15560 9141 15569
rect 9099 15520 9100 15560
rect 9140 15520 9141 15560
rect 9099 15511 9141 15520
rect 9196 14897 9236 17023
rect 9388 16316 9428 17872
rect 9484 17501 9524 18292
rect 9580 18005 9620 22903
rect 9868 22700 9908 27691
rect 10059 27656 10101 27665
rect 10059 27616 10060 27656
rect 10100 27616 10101 27656
rect 10059 27607 10101 27616
rect 9963 24716 10005 24725
rect 9963 24676 9964 24716
rect 10004 24676 10005 24716
rect 9963 24667 10005 24676
rect 9964 24632 10004 24667
rect 9964 24581 10004 24592
rect 10060 24632 10100 27607
rect 10252 27245 10292 28288
rect 10540 27833 10580 29800
rect 10636 28412 10676 31396
rect 10828 30680 10868 32647
rect 10828 30631 10868 30640
rect 10924 29840 10964 33664
rect 11019 33704 11061 33713
rect 11019 33664 11020 33704
rect 11060 33664 11061 33704
rect 11019 33655 11061 33664
rect 11020 33570 11060 33655
rect 11019 31352 11061 31361
rect 11019 31312 11020 31352
rect 11060 31312 11061 31352
rect 11019 31303 11061 31312
rect 11116 31352 11156 31361
rect 10539 27824 10581 27833
rect 10539 27784 10540 27824
rect 10580 27784 10581 27824
rect 10539 27775 10581 27784
rect 10444 27656 10484 27665
rect 10251 27236 10293 27245
rect 10251 27196 10252 27236
rect 10292 27196 10293 27236
rect 10251 27187 10293 27196
rect 10348 27068 10388 27077
rect 10444 27068 10484 27616
rect 10539 27656 10581 27665
rect 10539 27616 10540 27656
rect 10580 27616 10581 27656
rect 10539 27607 10581 27616
rect 10540 27522 10580 27607
rect 10388 27028 10484 27068
rect 10348 27019 10388 27028
rect 10156 26816 10196 26827
rect 10156 26741 10196 26776
rect 10155 26732 10197 26741
rect 10155 26692 10156 26732
rect 10196 26692 10197 26732
rect 10155 26683 10197 26692
rect 10347 26732 10389 26741
rect 10347 26692 10348 26732
rect 10388 26692 10389 26732
rect 10347 26683 10389 26692
rect 10348 25304 10388 26683
rect 10443 26144 10485 26153
rect 10443 26104 10444 26144
rect 10484 26104 10485 26144
rect 10443 26095 10485 26104
rect 10444 26010 10484 26095
rect 10636 26060 10676 28372
rect 10828 29800 10924 29840
rect 10732 28328 10772 28337
rect 10732 27749 10772 28288
rect 10731 27740 10773 27749
rect 10731 27700 10732 27740
rect 10772 27700 10773 27740
rect 10731 27691 10773 27700
rect 10828 27646 10868 29800
rect 10924 29791 10964 29800
rect 11020 29924 11060 31303
rect 11116 31109 11156 31312
rect 11115 31100 11157 31109
rect 11115 31060 11116 31100
rect 11156 31060 11157 31100
rect 11115 31051 11157 31060
rect 11020 29000 11060 29884
rect 10540 26020 10676 26060
rect 10732 27606 10868 27646
rect 10924 28960 11060 29000
rect 10540 25892 10580 26020
rect 10348 25255 10388 25264
rect 10444 25852 10580 25892
rect 10635 25892 10677 25901
rect 10635 25852 10636 25892
rect 10676 25852 10677 25892
rect 10444 25136 10484 25852
rect 10635 25843 10677 25852
rect 10636 25758 10676 25843
rect 10539 25220 10581 25229
rect 10539 25180 10540 25220
rect 10580 25180 10581 25220
rect 10539 25171 10581 25180
rect 10060 22961 10100 24592
rect 10348 25096 10484 25136
rect 10155 24548 10197 24557
rect 10155 24508 10156 24548
rect 10196 24508 10197 24548
rect 10155 24499 10197 24508
rect 10059 22952 10101 22961
rect 10059 22912 10060 22952
rect 10100 22912 10101 22952
rect 10059 22903 10101 22912
rect 9868 22660 10100 22700
rect 9964 22280 10004 22289
rect 9676 22196 9716 22205
rect 9964 22196 10004 22240
rect 9716 22156 10004 22196
rect 10060 22280 10100 22660
rect 10156 22541 10196 24499
rect 10252 23792 10292 23801
rect 10252 23213 10292 23752
rect 10348 23540 10388 25096
rect 10540 25086 10580 25171
rect 10444 24548 10484 24559
rect 10732 24557 10772 27606
rect 10924 27572 10964 28960
rect 11212 28505 11252 35680
rect 11308 35393 11348 36520
rect 11404 35972 11444 37360
rect 11500 37351 11540 37360
rect 11692 37148 11732 38284
rect 11787 37904 11829 37913
rect 11787 37864 11788 37904
rect 11828 37864 11829 37904
rect 11787 37855 11829 37864
rect 11307 35384 11349 35393
rect 11307 35344 11308 35384
rect 11348 35344 11349 35384
rect 11307 35335 11349 35344
rect 11307 33704 11349 33713
rect 11307 33664 11308 33704
rect 11348 33664 11349 33704
rect 11307 33655 11349 33664
rect 11019 28496 11061 28505
rect 11019 28456 11020 28496
rect 11060 28456 11061 28496
rect 11019 28447 11061 28456
rect 11211 28496 11253 28505
rect 11211 28456 11212 28496
rect 11252 28456 11253 28496
rect 11211 28447 11253 28456
rect 11020 27656 11060 28447
rect 11211 28328 11253 28337
rect 11211 28288 11212 28328
rect 11252 28288 11253 28328
rect 11211 28279 11253 28288
rect 11212 27749 11252 28279
rect 11211 27740 11253 27749
rect 11211 27700 11212 27740
rect 11252 27700 11253 27740
rect 11211 27691 11253 27700
rect 11060 27646 11156 27656
rect 11060 27616 11252 27646
rect 11020 27607 11060 27616
rect 11116 27606 11252 27616
rect 10924 27329 10964 27532
rect 10923 27320 10965 27329
rect 10923 27280 10924 27320
rect 10964 27280 10965 27320
rect 10923 27271 10965 27280
rect 11115 27320 11157 27329
rect 11115 27280 11116 27320
rect 11156 27280 11157 27320
rect 11115 27271 11157 27280
rect 11019 27236 11061 27245
rect 11019 27196 11020 27236
rect 11060 27196 11061 27236
rect 11019 27187 11061 27196
rect 10827 26816 10869 26825
rect 10827 26776 10828 26816
rect 10868 26776 10869 26816
rect 10827 26767 10869 26776
rect 10828 26573 10868 26767
rect 10827 26564 10869 26573
rect 10827 26524 10828 26564
rect 10868 26524 10869 26564
rect 10827 26515 10869 26524
rect 10923 26396 10965 26405
rect 10923 26356 10924 26396
rect 10964 26356 10965 26396
rect 10923 26347 10965 26356
rect 10827 26312 10869 26321
rect 10827 26272 10828 26312
rect 10868 26272 10869 26312
rect 10827 26263 10869 26272
rect 10828 26144 10868 26263
rect 10828 26069 10868 26104
rect 10827 26060 10869 26069
rect 10827 26020 10828 26060
rect 10868 26020 10869 26060
rect 10827 26011 10869 26020
rect 10827 25892 10869 25901
rect 10827 25852 10828 25892
rect 10868 25852 10869 25892
rect 10827 25843 10869 25852
rect 10828 25304 10868 25843
rect 10924 25397 10964 26347
rect 10923 25388 10965 25397
rect 10923 25348 10924 25388
rect 10964 25348 10965 25388
rect 10923 25339 10965 25348
rect 10828 25255 10868 25264
rect 10924 25304 10964 25339
rect 10924 25253 10964 25264
rect 11020 25136 11060 27187
rect 10828 25096 11060 25136
rect 10444 24473 10484 24508
rect 10539 24548 10581 24557
rect 10539 24508 10540 24548
rect 10580 24508 10581 24548
rect 10539 24499 10581 24508
rect 10731 24548 10773 24557
rect 10731 24508 10732 24548
rect 10772 24508 10773 24548
rect 10731 24499 10773 24508
rect 10443 24464 10485 24473
rect 10443 24424 10444 24464
rect 10484 24424 10485 24464
rect 10443 24415 10485 24424
rect 10540 24414 10580 24499
rect 10444 23717 10484 23802
rect 10732 23801 10772 23886
rect 10731 23792 10773 23801
rect 10731 23751 10732 23792
rect 10772 23751 10773 23792
rect 10731 23743 10773 23751
rect 10828 23792 10868 25096
rect 11019 24632 11061 24641
rect 11019 24592 11020 24632
rect 11060 24592 11061 24632
rect 11019 24583 11061 24592
rect 11020 24498 11060 24583
rect 11116 23960 11156 27271
rect 11212 26405 11252 27606
rect 11211 26396 11253 26405
rect 11211 26356 11212 26396
rect 11252 26356 11253 26396
rect 11211 26347 11253 26356
rect 11308 25472 11348 33655
rect 11404 33041 11444 35932
rect 11500 37108 11732 37148
rect 11500 35477 11540 37108
rect 11595 36980 11637 36989
rect 11595 36940 11596 36980
rect 11636 36940 11637 36980
rect 11595 36931 11637 36940
rect 11596 36140 11636 36931
rect 11691 36728 11733 36737
rect 11691 36688 11692 36728
rect 11732 36688 11733 36728
rect 11691 36679 11733 36688
rect 11596 36091 11636 36100
rect 11499 35468 11541 35477
rect 11499 35428 11500 35468
rect 11540 35428 11541 35468
rect 11499 35419 11541 35428
rect 11499 34964 11541 34973
rect 11499 34924 11500 34964
rect 11540 34924 11541 34964
rect 11499 34915 11541 34924
rect 11500 33699 11540 34915
rect 11692 33956 11732 36679
rect 11788 36233 11828 37855
rect 11787 36224 11829 36233
rect 11787 36184 11788 36224
rect 11828 36184 11829 36224
rect 11787 36175 11829 36184
rect 11884 36056 11924 40174
rect 11980 39752 12020 40804
rect 12268 40424 12308 40433
rect 12460 40424 12500 41299
rect 12308 40384 12500 40424
rect 12268 40375 12308 40384
rect 12556 40340 12596 42928
rect 12651 41012 12693 41021
rect 12651 40972 12652 41012
rect 12692 40972 12693 41012
rect 12651 40963 12693 40972
rect 12364 40300 12596 40340
rect 12076 40256 12116 40265
rect 12267 40256 12309 40265
rect 12116 40216 12268 40256
rect 12308 40216 12309 40256
rect 12076 40207 12116 40216
rect 12267 40207 12309 40216
rect 12171 40088 12213 40097
rect 12171 40048 12172 40088
rect 12212 40048 12213 40088
rect 12171 40039 12213 40048
rect 12076 39752 12116 39761
rect 11980 39712 12076 39752
rect 12076 39703 12116 39712
rect 12076 38996 12116 39005
rect 11980 38956 12076 38996
rect 11980 37745 12020 38956
rect 12076 38947 12116 38956
rect 12076 38249 12116 38280
rect 12075 38240 12117 38249
rect 12075 38200 12076 38240
rect 12116 38200 12117 38240
rect 12075 38191 12117 38200
rect 12172 38240 12212 40039
rect 12364 39836 12404 40300
rect 12555 40172 12597 40181
rect 12555 40132 12556 40172
rect 12596 40132 12597 40172
rect 12555 40123 12597 40132
rect 12268 39796 12404 39836
rect 12268 38921 12308 39796
rect 12459 39752 12501 39761
rect 12459 39712 12460 39752
rect 12500 39712 12501 39752
rect 12459 39703 12501 39712
rect 12556 39747 12596 40123
rect 12363 39668 12405 39677
rect 12363 39628 12364 39668
rect 12404 39628 12405 39668
rect 12363 39619 12405 39628
rect 12267 38912 12309 38921
rect 12267 38872 12268 38912
rect 12308 38872 12309 38912
rect 12267 38863 12309 38872
rect 12267 38744 12309 38753
rect 12267 38704 12268 38744
rect 12308 38704 12309 38744
rect 12267 38695 12309 38704
rect 12268 38610 12308 38695
rect 12268 38501 12308 38503
rect 12267 38492 12309 38501
rect 12267 38452 12268 38492
rect 12308 38452 12309 38492
rect 12267 38443 12309 38452
rect 12268 38408 12308 38443
rect 12268 38359 12308 38368
rect 12268 38249 12308 38268
rect 12267 38240 12309 38249
rect 12172 38200 12268 38240
rect 12308 38200 12309 38240
rect 12076 38156 12116 38191
rect 12076 38081 12116 38116
rect 12075 38072 12117 38081
rect 12075 38032 12076 38072
rect 12116 38032 12117 38072
rect 12075 38023 12117 38032
rect 12172 37820 12212 38200
rect 12267 38191 12309 38200
rect 12172 37780 12308 37820
rect 11979 37736 12021 37745
rect 11979 37696 11980 37736
rect 12020 37696 12021 37736
rect 11979 37687 12021 37696
rect 12171 36812 12213 36821
rect 12171 36772 12172 36812
rect 12212 36772 12213 36812
rect 12171 36763 12213 36772
rect 11980 36686 12020 36695
rect 12172 36678 12212 36763
rect 12268 36737 12308 37780
rect 12267 36728 12309 36737
rect 12267 36688 12268 36728
rect 12308 36688 12309 36728
rect 12267 36679 12309 36688
rect 11980 36401 12020 36646
rect 11979 36392 12021 36401
rect 11979 36352 11980 36392
rect 12020 36352 12021 36392
rect 11979 36343 12021 36352
rect 12267 36392 12309 36401
rect 12267 36352 12268 36392
rect 12308 36352 12309 36392
rect 12267 36343 12309 36352
rect 11500 33650 11540 33659
rect 11596 33916 11732 33956
rect 11788 36016 11924 36056
rect 11403 33032 11445 33041
rect 11403 32992 11404 33032
rect 11444 32992 11445 33032
rect 11403 32983 11445 32992
rect 11404 32864 11444 32873
rect 11596 32864 11636 33916
rect 11692 33788 11732 33797
rect 11692 33629 11732 33748
rect 11691 33620 11733 33629
rect 11691 33580 11692 33620
rect 11732 33580 11733 33620
rect 11691 33571 11733 33580
rect 11404 31445 11444 32824
rect 11500 32824 11636 32864
rect 11403 31436 11445 31445
rect 11403 31396 11404 31436
rect 11444 31396 11445 31436
rect 11403 31387 11445 31396
rect 11404 31025 11444 31387
rect 11403 31016 11445 31025
rect 11403 30976 11404 31016
rect 11444 30976 11445 31016
rect 11403 30967 11445 30976
rect 11500 30269 11540 32824
rect 11596 32696 11636 32705
rect 11596 31366 11636 32656
rect 11788 31352 11828 36016
rect 11884 35888 11924 35897
rect 11884 32957 11924 35848
rect 12268 35216 12308 36343
rect 12364 36140 12404 39619
rect 12460 38501 12500 39703
rect 12556 39698 12596 39707
rect 12652 39005 12692 40963
rect 12748 40424 12788 42928
rect 12940 41021 12980 42928
rect 13035 42440 13077 42449
rect 13035 42400 13036 42440
rect 13076 42400 13077 42440
rect 13035 42391 13077 42400
rect 12939 41012 12981 41021
rect 12939 40972 12940 41012
rect 12980 40972 12981 41012
rect 12939 40963 12981 40972
rect 12748 40384 12884 40424
rect 12748 39845 12788 39930
rect 12747 39836 12789 39845
rect 12747 39796 12748 39836
rect 12788 39796 12789 39836
rect 12747 39787 12789 39796
rect 12844 39668 12884 40384
rect 13036 40340 13076 42391
rect 13132 40424 13172 42928
rect 13324 40517 13364 42928
rect 13516 41609 13556 42928
rect 13611 42860 13653 42869
rect 13611 42820 13612 42860
rect 13652 42820 13653 42860
rect 13611 42811 13653 42820
rect 13515 41600 13557 41609
rect 13515 41560 13516 41600
rect 13556 41560 13557 41600
rect 13515 41551 13557 41560
rect 13612 41516 13652 42811
rect 13708 42113 13748 42928
rect 13707 42104 13749 42113
rect 13707 42064 13708 42104
rect 13748 42064 13749 42104
rect 13707 42055 13749 42064
rect 13612 41476 13748 41516
rect 13420 41264 13460 41273
rect 13323 40508 13365 40517
rect 13323 40468 13324 40508
rect 13364 40468 13365 40508
rect 13323 40459 13365 40468
rect 13132 40384 13268 40424
rect 13036 40300 13172 40340
rect 13132 39920 13172 40300
rect 13132 39871 13172 39880
rect 13035 39836 13077 39845
rect 13035 39796 13036 39836
rect 13076 39796 13077 39836
rect 13035 39787 13077 39796
rect 12748 39628 12884 39668
rect 12940 39668 12980 39677
rect 12651 38996 12693 39005
rect 12651 38956 12652 38996
rect 12692 38956 12693 38996
rect 12651 38947 12693 38956
rect 12555 38912 12597 38921
rect 12555 38872 12556 38912
rect 12596 38872 12597 38912
rect 12555 38863 12597 38872
rect 12459 38492 12501 38501
rect 12459 38452 12460 38492
rect 12500 38452 12501 38492
rect 12459 38443 12501 38452
rect 12459 38240 12501 38249
rect 12459 38200 12460 38240
rect 12500 38200 12501 38240
rect 12459 38191 12501 38200
rect 12460 38156 12500 38191
rect 12460 38105 12500 38116
rect 12556 37913 12596 38863
rect 12651 38492 12693 38501
rect 12651 38452 12652 38492
rect 12692 38452 12693 38492
rect 12651 38443 12693 38452
rect 12652 38408 12692 38443
rect 12652 38357 12692 38368
rect 12555 37904 12597 37913
rect 12555 37864 12556 37904
rect 12596 37864 12597 37904
rect 12555 37855 12597 37864
rect 12556 37325 12596 37855
rect 12748 37820 12788 39628
rect 12940 39089 12980 39628
rect 12939 39080 12981 39089
rect 12939 39040 12940 39080
rect 12980 39040 12981 39080
rect 12939 39031 12981 39040
rect 13036 38828 13076 39787
rect 13228 39341 13268 40384
rect 13420 40097 13460 41224
rect 13612 41012 13652 41021
rect 13516 40424 13556 40433
rect 13419 40088 13461 40097
rect 13419 40048 13420 40088
rect 13460 40048 13461 40088
rect 13419 40039 13461 40048
rect 13324 39752 13364 39761
rect 13227 39332 13269 39341
rect 13227 39292 13228 39332
rect 13268 39292 13269 39332
rect 13227 39283 13269 39292
rect 13036 38788 13172 38828
rect 12843 38408 12885 38417
rect 12843 38368 12844 38408
rect 12884 38368 12885 38408
rect 12843 38359 12885 38368
rect 13035 38408 13077 38417
rect 13035 38368 13036 38408
rect 13076 38368 13077 38408
rect 13035 38359 13077 38368
rect 12844 38156 12884 38359
rect 12939 38324 12981 38333
rect 12939 38284 12940 38324
rect 12980 38284 12981 38324
rect 12939 38275 12981 38284
rect 12844 38107 12884 38116
rect 12940 37820 12980 38275
rect 13036 38274 13076 38359
rect 12652 37780 12788 37820
rect 12844 37780 12980 37820
rect 12555 37316 12597 37325
rect 12555 37276 12556 37316
rect 12596 37276 12597 37316
rect 12555 37267 12597 37276
rect 12459 36812 12501 36821
rect 12459 36772 12460 36812
rect 12500 36772 12501 36812
rect 12459 36763 12501 36772
rect 12460 36728 12500 36763
rect 12460 36677 12500 36688
rect 12556 36728 12596 36737
rect 12364 36091 12404 36100
rect 12268 35167 12308 35176
rect 12171 35132 12213 35141
rect 12171 35092 12172 35132
rect 12212 35092 12213 35132
rect 12171 35083 12213 35092
rect 12172 34964 12212 35083
rect 12363 35048 12405 35057
rect 12363 35008 12364 35048
rect 12404 35008 12405 35048
rect 12363 34999 12405 35008
rect 12267 34964 12309 34973
rect 12172 34924 12268 34964
rect 12308 34924 12309 34964
rect 12267 34915 12309 34924
rect 12268 34376 12308 34915
rect 11979 33788 12021 33797
rect 11979 33748 11980 33788
rect 12020 33748 12021 33788
rect 11979 33739 12021 33748
rect 11883 32948 11925 32957
rect 11883 32908 11884 32948
rect 11924 32908 11925 32948
rect 11883 32899 11925 32908
rect 11884 32814 11924 32899
rect 11980 32696 12020 33739
rect 12268 32864 12308 34336
rect 11596 31317 11636 31326
rect 11692 31312 11828 31352
rect 11884 32656 12020 32696
rect 12076 32824 12308 32864
rect 11692 30941 11732 31312
rect 11788 31184 11828 31193
rect 11884 31184 11924 32656
rect 11980 32192 12020 32201
rect 12076 32192 12116 32824
rect 12364 32705 12404 34999
rect 12460 34964 12500 34973
rect 12460 34385 12500 34924
rect 12459 34376 12501 34385
rect 12459 34336 12460 34376
rect 12500 34336 12501 34376
rect 12459 34327 12501 34336
rect 12460 34208 12500 34217
rect 12460 33704 12500 34168
rect 12460 33655 12500 33664
rect 12556 33704 12596 36688
rect 12652 35384 12692 37780
rect 12747 37568 12789 37577
rect 12747 37528 12748 37568
rect 12788 37528 12789 37568
rect 12747 37519 12789 37528
rect 12748 37400 12788 37519
rect 12748 36401 12788 37360
rect 12844 37064 12884 37780
rect 13132 37661 13172 38788
rect 13228 38156 13268 38165
rect 13131 37652 13173 37661
rect 13131 37612 13132 37652
rect 13172 37612 13173 37652
rect 13131 37603 13173 37612
rect 12940 37232 12980 37241
rect 12980 37192 13172 37232
rect 12940 37183 12980 37192
rect 12844 37024 13076 37064
rect 12843 36896 12885 36905
rect 12843 36856 12844 36896
rect 12884 36856 12885 36896
rect 12843 36847 12885 36856
rect 12747 36392 12789 36401
rect 12747 36352 12748 36392
rect 12788 36352 12789 36392
rect 12747 36343 12789 36352
rect 12652 35344 12788 35384
rect 12651 35216 12693 35225
rect 12651 35176 12652 35216
rect 12692 35176 12693 35216
rect 12651 35167 12693 35176
rect 12652 35082 12692 35167
rect 12748 34049 12788 35344
rect 12747 34040 12789 34049
rect 12747 34000 12748 34040
rect 12788 34000 12789 34040
rect 12747 33991 12789 34000
rect 12747 33704 12789 33713
rect 12596 33664 12748 33704
rect 12788 33664 12789 33704
rect 12556 33655 12596 33664
rect 12747 33655 12789 33664
rect 12651 32864 12693 32873
rect 12651 32824 12652 32864
rect 12692 32824 12693 32864
rect 12651 32815 12693 32824
rect 12652 32730 12692 32815
rect 12363 32696 12405 32705
rect 12363 32656 12364 32696
rect 12404 32656 12405 32696
rect 12363 32647 12405 32656
rect 12555 32696 12597 32705
rect 12555 32656 12556 32696
rect 12596 32656 12597 32696
rect 12555 32647 12597 32656
rect 12172 32276 12212 32285
rect 12212 32236 12500 32276
rect 12172 32227 12212 32236
rect 12020 32152 12116 32192
rect 12460 32192 12500 32236
rect 11980 31529 12020 32152
rect 12460 32143 12500 32152
rect 12556 32192 12596 32647
rect 12556 32117 12596 32152
rect 12555 32108 12597 32117
rect 12555 32068 12556 32108
rect 12596 32068 12597 32108
rect 12555 32059 12597 32068
rect 12459 31604 12501 31613
rect 12459 31564 12460 31604
rect 12500 31564 12501 31604
rect 12459 31555 12501 31564
rect 11979 31520 12021 31529
rect 11979 31480 11980 31520
rect 12020 31480 12021 31520
rect 11979 31471 12021 31480
rect 12363 31520 12405 31529
rect 12363 31480 12364 31520
rect 12404 31480 12405 31520
rect 12363 31471 12405 31480
rect 11828 31144 11924 31184
rect 11788 31135 11828 31144
rect 11691 30932 11733 30941
rect 11691 30892 11692 30932
rect 11732 30892 11733 30932
rect 11691 30883 11733 30892
rect 12075 30932 12117 30941
rect 12075 30892 12076 30932
rect 12116 30892 12117 30932
rect 12075 30883 12117 30892
rect 11499 30260 11541 30269
rect 11499 30220 11500 30260
rect 11540 30220 11541 30260
rect 11499 30211 11541 30220
rect 11500 29840 11540 29849
rect 11212 25432 11348 25472
rect 11404 29800 11500 29840
rect 11212 24296 11252 25432
rect 11404 25397 11444 29800
rect 11500 29791 11540 29800
rect 11692 29336 11732 30883
rect 12076 30680 12116 30883
rect 12076 30631 12116 30640
rect 12268 30428 12308 30437
rect 11980 30388 12268 30428
rect 11883 30008 11925 30017
rect 11883 29968 11884 30008
rect 11924 29968 11925 30008
rect 11883 29959 11925 29968
rect 11884 29513 11924 29959
rect 11980 29854 12020 30388
rect 12268 30379 12308 30388
rect 12171 29924 12213 29933
rect 12171 29884 12172 29924
rect 12212 29884 12213 29924
rect 12171 29875 12213 29884
rect 11980 29805 12020 29814
rect 12172 29756 12212 29875
rect 12172 29707 12212 29716
rect 11883 29504 11925 29513
rect 11883 29464 11884 29504
rect 11924 29464 11925 29504
rect 11883 29455 11925 29464
rect 11500 29296 11732 29336
rect 11500 27656 11540 29296
rect 11595 29168 11637 29177
rect 11595 29128 11596 29168
rect 11636 29128 11637 29168
rect 11595 29119 11637 29128
rect 11596 29034 11636 29119
rect 11884 29009 11924 29455
rect 11979 29420 12021 29429
rect 11979 29380 11980 29420
rect 12020 29380 12021 29420
rect 11979 29371 12021 29380
rect 11980 29168 12020 29371
rect 11691 29000 11733 29009
rect 11691 28960 11692 29000
rect 11732 28960 11733 29000
rect 11691 28951 11733 28960
rect 11883 29000 11925 29009
rect 11883 28960 11884 29000
rect 11924 28960 11925 29000
rect 11883 28951 11925 28960
rect 11692 28496 11732 28951
rect 11500 25649 11540 27616
rect 11596 28456 11732 28496
rect 11788 28916 11828 28925
rect 11596 25724 11636 28456
rect 11788 28412 11828 28876
rect 11740 28372 11828 28412
rect 11883 28412 11925 28421
rect 11883 28372 11884 28412
rect 11924 28372 11925 28412
rect 11740 28370 11780 28372
rect 11883 28363 11925 28372
rect 11740 28321 11780 28330
rect 11884 28244 11924 28363
rect 11884 28195 11924 28204
rect 11980 27740 12020 29128
rect 12075 29168 12117 29177
rect 12075 29128 12076 29168
rect 12116 29128 12117 29168
rect 12075 29119 12117 29128
rect 11788 27700 12020 27740
rect 11596 25684 11732 25724
rect 11499 25640 11541 25649
rect 11499 25600 11500 25640
rect 11540 25600 11636 25640
rect 11499 25591 11541 25600
rect 11403 25388 11445 25397
rect 11403 25348 11404 25388
rect 11444 25348 11445 25388
rect 11403 25339 11445 25348
rect 11308 25304 11348 25313
rect 11308 24473 11348 25264
rect 11404 25254 11444 25339
rect 11499 25220 11541 25229
rect 11499 25180 11500 25220
rect 11540 25180 11541 25220
rect 11499 25171 11541 25180
rect 11403 25136 11445 25145
rect 11403 25096 11404 25136
rect 11444 25096 11445 25136
rect 11403 25087 11445 25096
rect 11307 24464 11349 24473
rect 11307 24424 11308 24464
rect 11348 24424 11349 24464
rect 11307 24415 11349 24424
rect 11212 24256 11348 24296
rect 11020 23920 11156 23960
rect 10923 23876 10965 23885
rect 10923 23836 10924 23876
rect 10964 23836 10965 23876
rect 10923 23827 10965 23836
rect 10732 23742 10772 23743
rect 10443 23708 10485 23717
rect 10443 23668 10444 23708
rect 10484 23668 10485 23708
rect 10443 23659 10485 23668
rect 10348 23500 10676 23540
rect 10347 23372 10389 23381
rect 10347 23332 10348 23372
rect 10388 23332 10389 23372
rect 10347 23323 10389 23332
rect 10251 23204 10293 23213
rect 10251 23164 10252 23204
rect 10292 23164 10293 23204
rect 10251 23155 10293 23164
rect 10155 22532 10197 22541
rect 10155 22492 10156 22532
rect 10196 22492 10197 22532
rect 10155 22483 10197 22492
rect 10252 22289 10292 23155
rect 9676 22147 9716 22156
rect 9675 22028 9717 22037
rect 9675 21988 9676 22028
rect 9716 21988 9717 22028
rect 9675 21979 9717 21988
rect 9676 18593 9716 21979
rect 9867 21944 9909 21953
rect 9867 21904 9868 21944
rect 9908 21904 9909 21944
rect 9867 21895 9909 21904
rect 9771 21608 9813 21617
rect 9771 21568 9772 21608
rect 9812 21568 9813 21608
rect 9771 21559 9813 21568
rect 9868 21608 9908 21895
rect 9868 21559 9908 21568
rect 9772 20096 9812 21559
rect 9675 18584 9717 18593
rect 9675 18544 9676 18584
rect 9716 18544 9717 18584
rect 9675 18535 9717 18544
rect 9675 18332 9717 18341
rect 9675 18292 9676 18332
rect 9716 18292 9717 18332
rect 9675 18283 9717 18292
rect 9676 18198 9716 18283
rect 9579 17996 9621 18005
rect 9579 17956 9580 17996
rect 9620 17956 9621 17996
rect 9579 17947 9621 17956
rect 9675 17912 9717 17921
rect 9675 17872 9676 17912
rect 9716 17872 9717 17912
rect 9772 17912 9812 20056
rect 9868 18584 9908 18593
rect 9868 18257 9908 18544
rect 9867 18248 9909 18257
rect 9867 18208 9868 18248
rect 9908 18208 10004 18248
rect 9867 18199 9909 18208
rect 9772 17872 9908 17912
rect 9675 17863 9717 17872
rect 9676 17828 9716 17863
rect 9676 17777 9716 17788
rect 9772 17744 9812 17755
rect 9772 17669 9812 17704
rect 9771 17660 9813 17669
rect 9771 17620 9772 17660
rect 9812 17620 9813 17660
rect 9771 17611 9813 17620
rect 9483 17492 9525 17501
rect 9483 17452 9484 17492
rect 9524 17452 9525 17492
rect 9483 17443 9525 17452
rect 9484 16745 9524 17443
rect 9483 16736 9525 16745
rect 9483 16696 9484 16736
rect 9524 16696 9525 16736
rect 9483 16687 9525 16696
rect 9868 16661 9908 17872
rect 9964 17501 10004 18208
rect 9963 17492 10005 17501
rect 9963 17452 9964 17492
rect 10004 17452 10005 17492
rect 9963 17443 10005 17452
rect 9964 17081 10004 17166
rect 9963 17072 10005 17081
rect 9963 17032 9964 17072
rect 10004 17032 10005 17072
rect 9963 17023 10005 17032
rect 9867 16652 9909 16661
rect 9867 16612 9868 16652
rect 9908 16612 9909 16652
rect 9867 16603 9909 16612
rect 9867 16400 9909 16409
rect 9867 16360 9868 16400
rect 9908 16360 9909 16400
rect 9867 16351 9909 16360
rect 9483 16316 9525 16325
rect 9388 16276 9484 16316
rect 9524 16276 9525 16316
rect 9483 16267 9525 16276
rect 9484 16232 9524 16267
rect 9484 16181 9524 16192
rect 9292 16064 9332 16073
rect 9332 16024 9524 16064
rect 9292 16015 9332 16024
rect 9484 15555 9524 16024
rect 9484 15476 9524 15515
rect 9676 15644 9716 15653
rect 9484 15436 9620 15476
rect 9291 14972 9333 14981
rect 9291 14932 9292 14972
rect 9332 14932 9333 14972
rect 9291 14923 9333 14932
rect 9195 14888 9237 14897
rect 9195 14848 9196 14888
rect 9236 14848 9237 14888
rect 9195 14839 9237 14848
rect 9099 14804 9141 14813
rect 9099 14764 9100 14804
rect 9140 14764 9141 14804
rect 9099 14755 9141 14764
rect 9100 14720 9140 14755
rect 9292 14720 9332 14923
rect 9100 14669 9140 14680
rect 9196 14680 9332 14720
rect 9580 14734 9620 15436
rect 9676 14981 9716 15604
rect 9675 14972 9717 14981
rect 9675 14932 9676 14972
rect 9716 14932 9717 14972
rect 9675 14923 9717 14932
rect 9580 14685 9620 14694
rect 9099 14132 9141 14141
rect 9004 14092 9100 14132
rect 9140 14092 9141 14132
rect 9099 14083 9141 14092
rect 9196 14132 9236 14680
rect 9772 14552 9812 14561
rect 9772 14141 9812 14512
rect 9196 14083 9236 14092
rect 9291 14132 9333 14141
rect 9291 14092 9292 14132
rect 9332 14092 9333 14132
rect 9291 14083 9333 14092
rect 9771 14132 9813 14141
rect 9771 14092 9772 14132
rect 9812 14092 9813 14132
rect 9771 14083 9813 14092
rect 8908 13831 8948 13840
rect 8715 13796 8757 13805
rect 8715 13756 8716 13796
rect 8756 13756 8757 13796
rect 8715 13747 8757 13756
rect 8716 13662 8756 13747
rect 8907 13712 8949 13721
rect 8907 13672 8908 13712
rect 8948 13672 8949 13712
rect 8907 13663 8949 13672
rect 8619 13628 8661 13637
rect 8619 13588 8620 13628
rect 8660 13588 8661 13628
rect 8619 13579 8661 13588
rect 8716 13553 8756 13555
rect 8523 13544 8565 13553
rect 8523 13504 8524 13544
rect 8564 13504 8565 13544
rect 8523 13495 8565 13504
rect 8715 13544 8757 13553
rect 8715 13504 8716 13544
rect 8756 13504 8757 13544
rect 8715 13495 8757 13504
rect 8716 13460 8756 13495
rect 8716 13411 8756 13420
rect 8524 13208 8564 13217
rect 8428 13168 8524 13208
rect 8331 13040 8373 13049
rect 8331 13000 8332 13040
rect 8372 13000 8373 13040
rect 8331 12991 8373 13000
rect 8332 12536 8372 12545
rect 8236 12496 8332 12536
rect 8236 11201 8276 12496
rect 8332 12487 8372 12496
rect 8332 11696 8372 11705
rect 8428 11696 8468 13168
rect 8524 13159 8564 13168
rect 8908 13208 8948 13663
rect 8908 13159 8948 13168
rect 8523 13040 8565 13049
rect 8523 13000 8524 13040
rect 8564 13000 8565 13040
rect 8523 12991 8565 13000
rect 8716 13040 8756 13049
rect 8524 11948 8564 12991
rect 8716 12872 8756 13000
rect 8716 12832 8948 12872
rect 8811 12536 8853 12545
rect 8811 12496 8812 12536
rect 8852 12496 8853 12536
rect 8811 12487 8853 12496
rect 8812 12402 8852 12487
rect 8620 12284 8660 12293
rect 8620 12125 8660 12244
rect 8715 12200 8757 12209
rect 8715 12160 8716 12200
rect 8756 12160 8757 12200
rect 8715 12151 8757 12160
rect 8619 12116 8661 12125
rect 8619 12076 8620 12116
rect 8660 12076 8661 12116
rect 8619 12067 8661 12076
rect 8716 11948 8756 12151
rect 8524 11908 8660 11948
rect 8372 11656 8468 11696
rect 8332 11453 8372 11656
rect 8428 11572 8564 11612
rect 8331 11444 8373 11453
rect 8331 11404 8332 11444
rect 8372 11404 8373 11444
rect 8331 11395 8373 11404
rect 8428 11285 8468 11572
rect 8524 11528 8564 11572
rect 8524 11479 8564 11488
rect 8427 11276 8469 11285
rect 8427 11236 8428 11276
rect 8468 11236 8564 11276
rect 8427 11227 8469 11236
rect 8235 11192 8277 11201
rect 8235 11152 8236 11192
rect 8276 11152 8277 11192
rect 8235 11143 8277 11152
rect 8331 11024 8373 11033
rect 8331 10984 8332 11024
rect 8372 10984 8373 11024
rect 8331 10975 8373 10984
rect 8428 11024 8468 11033
rect 7852 10564 8180 10604
rect 7755 10268 7797 10277
rect 7755 10228 7756 10268
rect 7796 10228 7797 10268
rect 7755 10219 7797 10228
rect 7660 10135 7700 10144
rect 7756 10184 7796 10219
rect 7564 10050 7604 10135
rect 7756 10133 7796 10144
rect 7276 9640 7412 9680
rect 7179 9092 7221 9101
rect 7179 9052 7180 9092
rect 7220 9052 7221 9092
rect 7179 9043 7221 9052
rect 7028 7960 7124 8000
rect 7180 8672 7220 9043
rect 6988 7951 7028 7960
rect 6892 7916 6932 7925
rect 6892 7748 6932 7876
rect 6892 7708 7028 7748
rect 6891 7580 6933 7589
rect 6891 7540 6892 7580
rect 6932 7540 6933 7580
rect 6891 7531 6933 7540
rect 6892 6656 6932 7531
rect 6892 6607 6932 6616
rect 6988 6488 7028 7708
rect 7180 7253 7220 8632
rect 7179 7244 7221 7253
rect 7179 7204 7180 7244
rect 7220 7204 7221 7244
rect 7179 7195 7221 7204
rect 7180 6665 7220 7195
rect 7179 6656 7221 6665
rect 7179 6616 7180 6656
rect 7220 6616 7221 6656
rect 7179 6607 7221 6616
rect 7276 6572 7316 9640
rect 7467 9596 7509 9605
rect 7467 9556 7468 9596
rect 7508 9556 7509 9596
rect 7467 9547 7509 9556
rect 7755 9596 7797 9605
rect 7755 9556 7756 9596
rect 7796 9556 7797 9596
rect 7755 9547 7797 9556
rect 7372 9512 7412 9521
rect 7372 9344 7412 9472
rect 7468 9512 7508 9547
rect 7468 9461 7508 9472
rect 7756 9512 7796 9547
rect 7563 9344 7605 9353
rect 7372 9304 7564 9344
rect 7604 9304 7605 9344
rect 7563 9295 7605 9304
rect 7467 9092 7509 9101
rect 7467 9052 7468 9092
rect 7508 9052 7509 9092
rect 7467 9043 7509 9052
rect 7468 8000 7508 9043
rect 7468 7951 7508 7960
rect 7467 7748 7509 7757
rect 7467 7708 7468 7748
rect 7508 7708 7509 7748
rect 7467 7699 7509 7708
rect 7276 6532 7412 6572
rect 6892 6448 7028 6488
rect 7084 6488 7124 6497
rect 7124 6448 7316 6488
rect 6892 6161 6932 6448
rect 7084 6439 7124 6448
rect 7083 6320 7125 6329
rect 7083 6280 7084 6320
rect 7124 6280 7125 6320
rect 7083 6271 7125 6280
rect 6987 6236 7029 6245
rect 6987 6196 6988 6236
rect 7028 6196 7029 6236
rect 6987 6187 7029 6196
rect 6891 6152 6933 6161
rect 6891 6112 6892 6152
rect 6932 6112 6933 6152
rect 6891 6103 6933 6112
rect 6892 5909 6932 6103
rect 6891 5900 6933 5909
rect 6891 5860 6892 5900
rect 6932 5860 6933 5900
rect 6891 5851 6933 5860
rect 6988 5657 7028 6187
rect 7084 5909 7124 6271
rect 7180 6236 7220 6245
rect 7083 5900 7125 5909
rect 7083 5860 7084 5900
rect 7124 5860 7125 5900
rect 7083 5851 7125 5860
rect 6987 5648 7029 5657
rect 6987 5608 6988 5648
rect 7028 5608 7029 5648
rect 6987 5599 7029 5608
rect 6988 5514 7028 5599
rect 6795 5396 6837 5405
rect 6795 5356 6796 5396
rect 6836 5356 6837 5396
rect 6795 5347 6837 5356
rect 7180 5321 7220 6196
rect 6603 5312 6645 5321
rect 6603 5272 6604 5312
rect 6644 5272 6645 5312
rect 6603 5263 6645 5272
rect 7179 5312 7221 5321
rect 7179 5272 7180 5312
rect 7220 5272 7221 5312
rect 7179 5263 7221 5272
rect 6508 4976 6548 4985
rect 6508 4817 6548 4936
rect 6507 4808 6549 4817
rect 6507 4768 6508 4808
rect 6548 4768 6549 4808
rect 6507 4759 6549 4768
rect 6412 4600 6548 4640
rect 6508 4313 6548 4600
rect 6507 4304 6549 4313
rect 6507 4264 6508 4304
rect 6548 4264 6549 4304
rect 6507 4255 6549 4264
rect 6411 4136 6453 4145
rect 6411 4096 6412 4136
rect 6452 4096 6453 4136
rect 6411 4087 6453 4096
rect 6412 4002 6452 4087
rect 6508 3557 6548 4255
rect 6507 3548 6549 3557
rect 6507 3508 6508 3548
rect 6548 3508 6549 3548
rect 6507 3499 6549 3508
rect 6508 3464 6548 3499
rect 6604 3464 6644 5263
rect 7084 4976 7124 4985
rect 7084 4733 7124 4936
rect 7179 4976 7221 4985
rect 7179 4936 7180 4976
rect 7220 4936 7221 4976
rect 7179 4927 7221 4936
rect 7180 4842 7220 4927
rect 6699 4724 6741 4733
rect 6699 4684 6700 4724
rect 6740 4684 6741 4724
rect 6699 4675 6741 4684
rect 7083 4724 7125 4733
rect 7083 4684 7084 4724
rect 7124 4684 7125 4724
rect 7083 4675 7125 4684
rect 6700 4590 6740 4675
rect 7276 4313 7316 6448
rect 7372 4901 7412 6532
rect 7468 5573 7508 7699
rect 7467 5564 7509 5573
rect 7467 5524 7468 5564
rect 7508 5524 7509 5564
rect 7467 5515 7509 5524
rect 7371 4892 7413 4901
rect 7371 4852 7372 4892
rect 7412 4852 7413 4892
rect 7371 4843 7413 4852
rect 7371 4724 7413 4733
rect 7371 4684 7372 4724
rect 7412 4684 7413 4724
rect 7371 4675 7413 4684
rect 7275 4304 7317 4313
rect 7275 4264 7276 4304
rect 7316 4264 7317 4304
rect 7275 4255 7317 4264
rect 6892 4141 6932 4150
rect 6700 3632 6740 3641
rect 6892 3632 6932 4101
rect 7276 4136 7316 4145
rect 7372 4136 7412 4675
rect 7468 4481 7508 5515
rect 7564 4892 7604 9295
rect 7659 8420 7701 8429
rect 7659 8380 7660 8420
rect 7700 8380 7701 8420
rect 7659 8371 7701 8380
rect 7660 7328 7700 8371
rect 7756 7505 7796 9472
rect 7852 8429 7892 10564
rect 8235 10436 8277 10445
rect 8235 10396 8236 10436
rect 8276 10396 8277 10436
rect 8235 10387 8277 10396
rect 7948 10352 7988 10361
rect 7948 10193 7988 10312
rect 8043 10352 8085 10361
rect 8043 10312 8044 10352
rect 8084 10312 8085 10352
rect 8043 10303 8085 10312
rect 7947 10184 7989 10193
rect 7947 10144 7948 10184
rect 7988 10144 7989 10184
rect 7947 10135 7989 10144
rect 8044 9605 8084 10303
rect 8139 10268 8181 10277
rect 8139 10228 8140 10268
rect 8180 10228 8181 10268
rect 8139 10219 8181 10228
rect 8140 10184 8180 10219
rect 8140 10133 8180 10144
rect 8236 10184 8276 10387
rect 8043 9596 8085 9605
rect 8043 9556 8044 9596
rect 8084 9556 8085 9596
rect 8043 9547 8085 9556
rect 8236 8765 8276 10144
rect 8332 10184 8372 10975
rect 8428 10193 8468 10984
rect 8524 10277 8564 11236
rect 8523 10268 8565 10277
rect 8523 10228 8524 10268
rect 8564 10228 8565 10268
rect 8523 10219 8565 10228
rect 8332 10135 8372 10144
rect 8427 10184 8469 10193
rect 8427 10144 8428 10184
rect 8468 10144 8469 10184
rect 8427 10135 8469 10144
rect 8427 9596 8469 9605
rect 8427 9556 8428 9596
rect 8468 9556 8469 9596
rect 8427 9547 8469 9556
rect 8043 8756 8085 8765
rect 8043 8716 8044 8756
rect 8084 8716 8085 8756
rect 8043 8707 8085 8716
rect 8235 8756 8277 8765
rect 8235 8716 8236 8756
rect 8276 8716 8277 8756
rect 8235 8707 8277 8716
rect 7851 8420 7893 8429
rect 7851 8380 7852 8420
rect 7892 8380 7893 8420
rect 7851 8371 7893 8380
rect 7948 7986 7988 7995
rect 7755 7496 7797 7505
rect 7755 7456 7756 7496
rect 7796 7456 7797 7496
rect 7755 7447 7797 7456
rect 7852 7412 7892 7421
rect 7948 7412 7988 7946
rect 7892 7372 7988 7412
rect 7852 7363 7892 7372
rect 7660 7288 7796 7328
rect 7660 7160 7700 7171
rect 7660 7085 7700 7120
rect 7659 7076 7701 7085
rect 7659 7036 7660 7076
rect 7700 7036 7701 7076
rect 7659 7027 7701 7036
rect 7756 5237 7796 7288
rect 7755 5228 7797 5237
rect 7755 5188 7756 5228
rect 7796 5188 7797 5228
rect 7755 5179 7797 5188
rect 8044 4976 8084 8707
rect 8139 8084 8181 8093
rect 8139 8044 8140 8084
rect 8180 8044 8181 8084
rect 8139 8035 8181 8044
rect 8140 7950 8180 8035
rect 8236 7589 8276 8707
rect 8332 8672 8372 8681
rect 8332 8009 8372 8632
rect 8331 8000 8373 8009
rect 8331 7960 8332 8000
rect 8372 7960 8373 8000
rect 8331 7951 8373 7960
rect 8428 8000 8468 9547
rect 8523 9092 8565 9101
rect 8523 9052 8524 9092
rect 8564 9052 8565 9092
rect 8523 9043 8565 9052
rect 8235 7580 8277 7589
rect 8235 7540 8236 7580
rect 8276 7540 8277 7580
rect 8235 7531 8277 7540
rect 8332 7169 8372 7254
rect 8331 7160 8373 7169
rect 8331 7120 8332 7160
rect 8372 7120 8373 7160
rect 8331 7111 8373 7120
rect 8428 6992 8468 7960
rect 8524 7169 8564 9043
rect 8620 7589 8660 11908
rect 8716 11899 8756 11908
rect 8908 11780 8948 12832
rect 9003 12368 9045 12377
rect 9003 12328 9004 12368
rect 9044 12328 9045 12368
rect 9003 12319 9045 12328
rect 8716 11740 8948 11780
rect 8716 11696 8756 11740
rect 8716 11033 8756 11656
rect 9004 11696 9044 12319
rect 9004 11647 9044 11656
rect 9100 11528 9140 14083
rect 9292 14048 9332 14083
rect 9292 13997 9332 14008
rect 9579 14048 9621 14057
rect 9579 14008 9580 14048
rect 9620 14008 9621 14048
rect 9579 13999 9621 14008
rect 9580 13914 9620 13999
rect 9483 13712 9525 13721
rect 9483 13672 9484 13712
rect 9524 13672 9525 13712
rect 9483 13663 9525 13672
rect 9291 12536 9333 12545
rect 9291 12496 9292 12536
rect 9332 12496 9333 12536
rect 9291 12487 9333 12496
rect 9292 12209 9332 12487
rect 9291 12200 9333 12209
rect 9291 12160 9292 12200
rect 9332 12160 9333 12200
rect 9291 12151 9333 12160
rect 9195 11948 9237 11957
rect 9195 11908 9196 11948
rect 9236 11908 9237 11948
rect 9195 11899 9237 11908
rect 9196 11814 9236 11899
rect 9195 11696 9237 11705
rect 9195 11656 9196 11696
rect 9236 11656 9237 11696
rect 9195 11647 9237 11656
rect 9004 11488 9140 11528
rect 9004 11360 9044 11488
rect 9196 11369 9236 11647
rect 9292 11621 9332 12151
rect 9484 11957 9524 13663
rect 9579 13208 9621 13217
rect 9579 13168 9580 13208
rect 9620 13168 9621 13208
rect 9579 13159 9621 13168
rect 9580 12545 9620 13159
rect 9579 12536 9621 12545
rect 9579 12496 9580 12536
rect 9620 12496 9621 12536
rect 9579 12487 9621 12496
rect 9483 11948 9525 11957
rect 9483 11908 9484 11948
rect 9524 11908 9525 11948
rect 9483 11899 9525 11908
rect 9579 11864 9621 11873
rect 9868 11864 9908 16351
rect 10060 13553 10100 22240
rect 10251 22280 10293 22289
rect 10251 22240 10252 22280
rect 10292 22240 10293 22280
rect 10251 22231 10293 22240
rect 10348 21701 10388 23323
rect 10539 22364 10581 22373
rect 10539 22324 10540 22364
rect 10580 22324 10581 22364
rect 10539 22315 10581 22324
rect 10443 22280 10485 22289
rect 10443 22240 10444 22280
rect 10484 22240 10485 22280
rect 10443 22231 10485 22240
rect 10347 21692 10389 21701
rect 10347 21652 10348 21692
rect 10388 21652 10389 21692
rect 10347 21643 10389 21652
rect 10444 21356 10484 22231
rect 10540 22230 10580 22315
rect 10444 21316 10580 21356
rect 10155 20936 10197 20945
rect 10155 20896 10156 20936
rect 10196 20896 10197 20936
rect 10155 20887 10197 20896
rect 10156 19928 10196 20887
rect 10444 20180 10484 20189
rect 10300 20054 10340 20063
rect 10300 20012 10340 20014
rect 10300 19972 10388 20012
rect 10156 19888 10292 19928
rect 10155 19760 10197 19769
rect 10155 19720 10156 19760
rect 10196 19720 10197 19760
rect 10155 19711 10197 19720
rect 10156 19265 10196 19711
rect 10155 19256 10197 19265
rect 10155 19216 10156 19256
rect 10196 19216 10197 19256
rect 10155 19207 10197 19216
rect 10156 19122 10196 19207
rect 10252 17912 10292 19888
rect 10348 19508 10388 19972
rect 10444 19937 10484 20140
rect 10443 19928 10485 19937
rect 10443 19888 10444 19928
rect 10484 19888 10485 19928
rect 10443 19879 10485 19888
rect 10443 19676 10485 19685
rect 10443 19636 10444 19676
rect 10484 19636 10485 19676
rect 10443 19627 10485 19636
rect 10444 19517 10484 19627
rect 10348 19459 10388 19468
rect 10443 19508 10485 19517
rect 10443 19468 10444 19508
rect 10484 19468 10485 19508
rect 10443 19459 10485 19468
rect 10444 19340 10484 19459
rect 10156 17872 10292 17912
rect 10348 19300 10484 19340
rect 10059 13544 10101 13553
rect 10059 13504 10060 13544
rect 10100 13504 10101 13544
rect 10059 13495 10101 13504
rect 10156 13376 10196 17872
rect 10251 17744 10293 17753
rect 10251 17704 10252 17744
rect 10292 17704 10293 17744
rect 10251 17695 10293 17704
rect 10252 17610 10292 17695
rect 10251 14804 10293 14813
rect 10251 14764 10252 14804
rect 10292 14764 10293 14804
rect 10251 14755 10293 14764
rect 10060 13336 10196 13376
rect 10060 13133 10100 13336
rect 10156 13208 10196 13217
rect 10059 13124 10101 13133
rect 10059 13084 10060 13124
rect 10100 13084 10101 13124
rect 10059 13075 10101 13084
rect 10156 12713 10196 13168
rect 10155 12704 10197 12713
rect 10155 12664 10156 12704
rect 10196 12664 10197 12704
rect 10155 12655 10197 12664
rect 10059 12536 10101 12545
rect 10059 12496 10060 12536
rect 10100 12496 10101 12536
rect 10059 12487 10101 12496
rect 10060 12402 10100 12487
rect 10059 12116 10101 12125
rect 10059 12076 10060 12116
rect 10100 12076 10101 12116
rect 10059 12067 10101 12076
rect 9579 11824 9580 11864
rect 9620 11824 9621 11864
rect 9579 11815 9621 11824
rect 9772 11824 9908 11864
rect 9580 11696 9620 11815
rect 9580 11647 9620 11656
rect 9772 11621 9812 11824
rect 10060 11705 10100 12067
rect 9867 11696 9909 11705
rect 9867 11656 9868 11696
rect 9908 11656 9909 11696
rect 9867 11647 9909 11656
rect 10059 11696 10101 11705
rect 10059 11656 10060 11696
rect 10100 11656 10101 11696
rect 10059 11647 10101 11656
rect 10156 11696 10196 11705
rect 9291 11612 9333 11621
rect 9291 11572 9292 11612
rect 9332 11572 9333 11612
rect 9291 11563 9333 11572
rect 9484 11612 9524 11621
rect 8812 11320 9044 11360
rect 9195 11360 9237 11369
rect 9195 11320 9196 11360
rect 9236 11320 9237 11360
rect 8715 11024 8757 11033
rect 8715 10984 8716 11024
rect 8756 10984 8757 11024
rect 8715 10975 8757 10984
rect 8812 10445 8852 11320
rect 9195 11311 9237 11320
rect 9003 11192 9045 11201
rect 9003 11152 9004 11192
rect 9044 11152 9045 11192
rect 9003 11143 9045 11152
rect 8907 11024 8949 11033
rect 8907 10984 8908 11024
rect 8948 10984 8949 11024
rect 8907 10975 8949 10984
rect 8908 10890 8948 10975
rect 9004 10940 9044 11143
rect 8907 10772 8949 10781
rect 8907 10732 8908 10772
rect 8948 10732 8949 10772
rect 8907 10723 8949 10732
rect 8811 10436 8853 10445
rect 8811 10396 8812 10436
rect 8852 10396 8853 10436
rect 8811 10387 8853 10396
rect 8716 10184 8756 10195
rect 8716 10109 8756 10144
rect 8812 10184 8852 10193
rect 8908 10184 8948 10723
rect 9004 10529 9044 10900
rect 9003 10520 9045 10529
rect 9003 10480 9004 10520
rect 9044 10480 9045 10520
rect 9003 10471 9045 10480
rect 9195 10520 9237 10529
rect 9195 10480 9196 10520
rect 9236 10480 9237 10520
rect 9195 10471 9237 10480
rect 9196 10268 9236 10471
rect 9292 10445 9332 11563
rect 9484 11444 9524 11572
rect 9771 11612 9813 11621
rect 9771 11572 9772 11612
rect 9812 11572 9813 11612
rect 9771 11563 9813 11572
rect 9868 11562 9908 11647
rect 9484 11404 9812 11444
rect 9483 11276 9525 11285
rect 9483 11236 9484 11276
rect 9524 11236 9525 11276
rect 9483 11227 9525 11236
rect 9388 11024 9428 11033
rect 9388 10781 9428 10984
rect 9484 11024 9524 11227
rect 9772 11192 9812 11404
rect 9772 11143 9812 11152
rect 9868 11024 9908 11033
rect 9484 10975 9524 10984
rect 9676 10984 9868 11024
rect 9387 10772 9429 10781
rect 9387 10732 9388 10772
rect 9428 10732 9429 10772
rect 9387 10723 9429 10732
rect 9291 10436 9333 10445
rect 9291 10396 9292 10436
rect 9332 10396 9333 10436
rect 9291 10387 9333 10396
rect 9483 10436 9525 10445
rect 9483 10396 9484 10436
rect 9524 10396 9620 10436
rect 9483 10387 9525 10396
rect 9196 10219 9236 10228
rect 9291 10268 9333 10277
rect 9291 10228 9292 10268
rect 9332 10228 9333 10268
rect 9291 10219 9333 10228
rect 8852 10144 8948 10184
rect 8715 10100 8757 10109
rect 8715 10060 8716 10100
rect 8756 10060 8757 10100
rect 8715 10051 8757 10060
rect 8812 9932 8852 10144
rect 9195 10100 9237 10109
rect 9195 10060 9196 10100
rect 9236 10060 9237 10100
rect 9195 10051 9237 10060
rect 8716 9892 8852 9932
rect 8716 9353 8756 9892
rect 9003 9848 9045 9857
rect 9003 9808 9004 9848
rect 9044 9808 9045 9848
rect 9003 9799 9045 9808
rect 8907 9680 8949 9689
rect 8907 9640 8908 9680
rect 8948 9640 8949 9680
rect 8907 9631 8949 9640
rect 8715 9344 8757 9353
rect 8715 9304 8716 9344
rect 8756 9304 8757 9344
rect 8715 9295 8757 9304
rect 8619 7580 8661 7589
rect 8619 7540 8620 7580
rect 8660 7540 8661 7580
rect 8619 7531 8661 7540
rect 8523 7160 8565 7169
rect 8523 7120 8524 7160
rect 8564 7120 8565 7160
rect 8523 7111 8565 7120
rect 8332 6952 8468 6992
rect 8139 6824 8181 6833
rect 8139 6784 8140 6824
rect 8180 6784 8181 6824
rect 8139 6775 8181 6784
rect 8140 5144 8180 6775
rect 8332 5732 8372 6952
rect 8716 6488 8756 6497
rect 8428 5900 8468 5909
rect 8716 5900 8756 6448
rect 8812 6488 8852 6497
rect 8908 6488 8948 9631
rect 9004 9512 9044 9799
rect 9196 9605 9236 10051
rect 9195 9596 9237 9605
rect 9195 9556 9196 9596
rect 9236 9556 9237 9596
rect 9195 9547 9237 9556
rect 9004 9463 9044 9472
rect 9196 9462 9236 9547
rect 9292 9269 9332 10219
rect 9483 10016 9525 10025
rect 9483 9976 9484 10016
rect 9524 9976 9525 10016
rect 9483 9967 9525 9976
rect 9099 9260 9141 9269
rect 9099 9220 9100 9260
rect 9140 9220 9141 9260
rect 9099 9211 9141 9220
rect 9291 9260 9333 9269
rect 9291 9220 9292 9260
rect 9332 9220 9333 9260
rect 9291 9211 9333 9220
rect 8852 6448 8948 6488
rect 8812 6439 8852 6448
rect 8468 5860 8756 5900
rect 8428 5851 8468 5860
rect 8332 5692 8468 5732
rect 8235 5648 8277 5657
rect 8235 5608 8236 5648
rect 8276 5608 8277 5648
rect 8235 5599 8277 5608
rect 8236 5514 8276 5599
rect 8140 5104 8276 5144
rect 8140 4976 8180 4985
rect 8044 4936 8140 4976
rect 8140 4927 8180 4936
rect 7467 4472 7509 4481
rect 7467 4432 7468 4472
rect 7508 4432 7509 4472
rect 7467 4423 7509 4432
rect 7316 4096 7412 4136
rect 7276 4087 7316 4096
rect 7083 4052 7125 4061
rect 7083 4012 7084 4052
rect 7124 4012 7125 4052
rect 7083 4003 7125 4012
rect 7084 3918 7124 4003
rect 6740 3592 6932 3632
rect 7084 3632 7124 3641
rect 7124 3592 7508 3632
rect 6700 3583 6740 3592
rect 7084 3583 7124 3592
rect 6988 3464 7028 3473
rect 7179 3464 7221 3473
rect 6604 3424 6740 3464
rect 6508 3413 6548 3424
rect 6316 3256 6644 3296
rect 6219 3212 6261 3221
rect 6219 3172 6220 3212
rect 6260 3172 6261 3212
rect 6219 3163 6261 3172
rect 6124 2575 6164 2584
rect 6220 2624 6260 3163
rect 6507 2960 6549 2969
rect 6507 2920 6508 2960
rect 6548 2920 6549 2960
rect 6507 2911 6549 2920
rect 6220 2575 6260 2584
rect 6508 2624 6548 2911
rect 6220 1952 6260 1961
rect 6220 1793 6260 1912
rect 6315 1952 6357 1961
rect 6315 1912 6316 1952
rect 6356 1912 6357 1952
rect 6315 1903 6357 1912
rect 6219 1784 6261 1793
rect 6219 1744 6220 1784
rect 6260 1744 6261 1784
rect 6219 1735 6261 1744
rect 5931 1448 5973 1457
rect 5931 1408 5932 1448
rect 5972 1408 5973 1448
rect 5931 1399 5973 1408
rect 6027 1364 6069 1373
rect 6027 1324 6028 1364
rect 6068 1324 6069 1364
rect 6027 1315 6069 1324
rect 6028 1230 6068 1315
rect 6123 1280 6165 1289
rect 6123 1240 6124 1280
rect 6164 1240 6165 1280
rect 6123 1231 6165 1240
rect 6220 1280 6260 1289
rect 6316 1280 6356 1903
rect 6411 1868 6453 1877
rect 6411 1828 6412 1868
rect 6452 1828 6453 1868
rect 6411 1819 6453 1828
rect 6260 1240 6356 1280
rect 6412 1700 6452 1819
rect 6220 1231 6260 1240
rect 6124 1112 6164 1231
rect 6028 1072 6164 1112
rect 6316 1112 6356 1121
rect 6412 1112 6452 1660
rect 6508 1457 6548 2584
rect 6604 2036 6644 3256
rect 6700 2213 6740 3424
rect 7028 3424 7124 3464
rect 6988 3415 7028 3424
rect 6987 3296 7029 3305
rect 6987 3256 6988 3296
rect 7028 3256 7029 3296
rect 6987 3247 7029 3256
rect 6891 2876 6933 2885
rect 6891 2836 6892 2876
rect 6932 2836 6933 2876
rect 6891 2827 6933 2836
rect 6795 2792 6837 2801
rect 6795 2752 6796 2792
rect 6836 2752 6837 2792
rect 6795 2743 6837 2752
rect 6796 2624 6836 2743
rect 6796 2575 6836 2584
rect 6892 2624 6932 2827
rect 6892 2575 6932 2584
rect 6988 2456 7028 3247
rect 7084 2969 7124 3424
rect 7179 3424 7180 3464
rect 7220 3424 7221 3464
rect 7468 3464 7508 3592
rect 7564 3557 7604 4852
rect 7659 4892 7701 4901
rect 7659 4852 7660 4892
rect 7700 4852 7701 4892
rect 7659 4843 7701 4852
rect 7660 3893 7700 4843
rect 7947 4472 7989 4481
rect 7947 4432 7948 4472
rect 7988 4432 7989 4472
rect 7947 4423 7989 4432
rect 7948 4145 7988 4423
rect 7947 4136 7989 4145
rect 7947 4096 7948 4136
rect 7988 4096 7989 4136
rect 7947 4087 7989 4096
rect 7659 3884 7701 3893
rect 7659 3844 7660 3884
rect 7700 3844 7701 3884
rect 7659 3835 7701 3844
rect 7659 3632 7701 3641
rect 7659 3592 7660 3632
rect 7700 3592 7701 3632
rect 7659 3583 7701 3592
rect 7563 3548 7605 3557
rect 7563 3508 7564 3548
rect 7604 3508 7605 3548
rect 7563 3499 7605 3508
rect 7179 3415 7221 3424
rect 7276 3445 7316 3454
rect 7180 3330 7220 3415
rect 7468 3415 7508 3424
rect 7276 3053 7316 3405
rect 7564 3380 7604 3389
rect 7275 3044 7317 3053
rect 7275 3004 7276 3044
rect 7316 3004 7317 3044
rect 7275 2995 7317 3004
rect 7083 2960 7125 2969
rect 7083 2920 7084 2960
rect 7124 2920 7125 2960
rect 7083 2911 7125 2920
rect 7180 2633 7220 2718
rect 6988 2407 7028 2416
rect 7084 2624 7124 2633
rect 6891 2372 6933 2381
rect 6891 2332 6892 2372
rect 6932 2332 6933 2372
rect 6891 2323 6933 2332
rect 6699 2204 6741 2213
rect 6699 2164 6700 2204
rect 6740 2164 6741 2204
rect 6699 2155 6741 2164
rect 6604 1996 6740 2036
rect 6604 1868 6644 1877
rect 6604 1625 6644 1828
rect 6603 1616 6645 1625
rect 6603 1576 6604 1616
rect 6644 1576 6645 1616
rect 6603 1567 6645 1576
rect 6507 1448 6549 1457
rect 6507 1408 6508 1448
rect 6548 1408 6549 1448
rect 6507 1399 6549 1408
rect 6356 1072 6452 1112
rect 6507 1112 6549 1121
rect 6507 1072 6508 1112
rect 6548 1072 6549 1112
rect 5739 1028 5781 1037
rect 5739 988 5740 1028
rect 5780 988 5781 1028
rect 5739 979 5781 988
rect 5740 894 5780 979
rect 5835 692 5877 701
rect 5835 652 5836 692
rect 5876 652 5877 692
rect 5835 643 5877 652
rect 5643 524 5685 533
rect 5643 484 5644 524
rect 5684 484 5685 524
rect 5643 475 5685 484
rect 5644 80 5684 475
rect 5836 80 5876 643
rect 6028 80 6068 1072
rect 6316 1063 6356 1072
rect 6507 1063 6549 1072
rect 6604 1112 6644 1121
rect 6508 978 6548 1063
rect 6604 953 6644 1072
rect 6603 944 6645 953
rect 6603 904 6604 944
rect 6644 904 6645 944
rect 6603 895 6645 904
rect 6700 776 6740 1996
rect 6892 1784 6932 2323
rect 6988 1961 7028 2046
rect 6987 1952 7029 1961
rect 6987 1912 6988 1952
rect 7028 1912 7029 1952
rect 6987 1903 7029 1912
rect 6988 1784 7028 1793
rect 6892 1744 6988 1784
rect 6988 1735 7028 1744
rect 6796 1700 6836 1709
rect 6796 1289 6836 1660
rect 7084 1532 7124 2584
rect 7179 2624 7221 2633
rect 7179 2584 7180 2624
rect 7220 2584 7221 2624
rect 7179 2575 7221 2584
rect 7281 2624 7321 2633
rect 7281 2549 7321 2584
rect 7564 2549 7604 3340
rect 7660 3296 7700 3583
rect 7851 3548 7893 3557
rect 7851 3508 7852 3548
rect 7892 3508 7893 3548
rect 7851 3499 7893 3508
rect 7852 3464 7892 3499
rect 7852 3413 7892 3424
rect 7756 3380 7796 3391
rect 7756 3305 7796 3340
rect 7660 3247 7700 3256
rect 7755 3296 7797 3305
rect 7755 3256 7756 3296
rect 7796 3256 7797 3296
rect 7755 3247 7797 3256
rect 7948 3128 7988 4087
rect 8236 3716 8276 5104
rect 8236 3676 8372 3716
rect 8236 3590 8276 3599
rect 8139 3548 8181 3557
rect 8236 3548 8276 3550
rect 8139 3508 8140 3548
rect 8180 3508 8276 3548
rect 8139 3499 8181 3508
rect 8043 3464 8085 3473
rect 8043 3424 8044 3464
rect 8084 3424 8085 3464
rect 8043 3415 8085 3424
rect 8044 3330 8084 3415
rect 8140 3380 8180 3389
rect 8140 3212 8180 3340
rect 8332 3380 8372 3676
rect 8428 3641 8468 5692
rect 8523 5648 8565 5657
rect 8523 5608 8524 5648
rect 8564 5608 8565 5648
rect 8523 5599 8565 5608
rect 8716 5648 8756 5860
rect 8716 5599 8756 5608
rect 8812 5648 8852 5657
rect 8524 4817 8564 5599
rect 8812 5321 8852 5608
rect 8908 5489 8948 6448
rect 8907 5480 8949 5489
rect 8907 5440 8908 5480
rect 8948 5440 8949 5480
rect 8907 5431 8949 5440
rect 8811 5312 8853 5321
rect 8811 5272 8812 5312
rect 8852 5272 8853 5312
rect 8811 5263 8853 5272
rect 8812 5060 8852 5069
rect 8620 4962 8660 4971
rect 8523 4808 8565 4817
rect 8523 4768 8524 4808
rect 8564 4768 8565 4808
rect 8523 4759 8565 4768
rect 8524 4136 8564 4759
rect 8620 4388 8660 4922
rect 8716 4388 8756 4397
rect 8620 4348 8716 4388
rect 8716 4339 8756 4348
rect 8619 4220 8661 4229
rect 8619 4180 8620 4220
rect 8660 4180 8661 4220
rect 8619 4171 8661 4180
rect 8524 3893 8564 4096
rect 8523 3884 8565 3893
rect 8523 3844 8524 3884
rect 8564 3844 8565 3884
rect 8523 3835 8565 3844
rect 8427 3632 8469 3641
rect 8427 3592 8428 3632
rect 8468 3592 8469 3632
rect 8427 3583 8469 3592
rect 8428 3464 8468 3475
rect 8428 3389 8468 3424
rect 8620 3464 8660 4171
rect 8812 3809 8852 5020
rect 9003 4976 9045 4985
rect 9003 4936 9004 4976
rect 9044 4936 9045 4976
rect 9003 4927 9045 4936
rect 8907 4136 8949 4145
rect 8907 4096 8908 4136
rect 8948 4096 8949 4136
rect 8907 4087 8949 4096
rect 9004 4136 9044 4927
rect 9100 4817 9140 9211
rect 9291 8588 9333 8597
rect 9291 8548 9292 8588
rect 9332 8548 9333 8588
rect 9291 8539 9333 8548
rect 9195 7580 9237 7589
rect 9195 7540 9196 7580
rect 9236 7540 9237 7580
rect 9195 7531 9237 7540
rect 9196 6488 9236 7531
rect 9196 6439 9236 6448
rect 9292 6488 9332 8539
rect 9387 7412 9429 7421
rect 9387 7372 9388 7412
rect 9428 7372 9429 7412
rect 9387 7363 9429 7372
rect 9292 6439 9332 6448
rect 9195 5984 9237 5993
rect 9195 5944 9196 5984
rect 9236 5944 9237 5984
rect 9195 5935 9237 5944
rect 9196 5825 9236 5935
rect 9195 5816 9237 5825
rect 9195 5776 9196 5816
rect 9236 5776 9237 5816
rect 9195 5767 9237 5776
rect 9196 5732 9236 5767
rect 9196 5682 9236 5692
rect 9291 5732 9333 5741
rect 9291 5692 9292 5732
rect 9332 5692 9333 5732
rect 9291 5683 9333 5692
rect 9292 5598 9332 5683
rect 9291 5312 9333 5321
rect 9291 5272 9292 5312
rect 9332 5272 9333 5312
rect 9291 5263 9333 5272
rect 9292 4892 9332 5263
rect 9388 4976 9428 7363
rect 9484 5648 9524 9967
rect 9580 8672 9620 10396
rect 9676 9680 9716 10984
rect 9868 10975 9908 10984
rect 9964 11024 10004 11033
rect 9964 10445 10004 10984
rect 10060 11024 10100 11033
rect 9963 10436 10005 10445
rect 9963 10396 9964 10436
rect 10004 10396 10005 10436
rect 9963 10387 10005 10396
rect 9771 10184 9813 10193
rect 9771 10144 9772 10184
rect 9812 10144 9813 10184
rect 9771 10135 9813 10144
rect 9772 10050 9812 10135
rect 10060 9680 10100 10984
rect 10156 10613 10196 11656
rect 10252 11360 10292 14755
rect 10348 13301 10388 19300
rect 10443 17828 10485 17837
rect 10443 17788 10444 17828
rect 10484 17788 10485 17828
rect 10443 17779 10485 17788
rect 10444 16073 10484 17779
rect 10443 16064 10485 16073
rect 10443 16024 10444 16064
rect 10484 16024 10485 16064
rect 10443 16015 10485 16024
rect 10540 15896 10580 21316
rect 10444 15856 10580 15896
rect 10444 13385 10484 15856
rect 10539 15728 10581 15737
rect 10539 15688 10540 15728
rect 10580 15688 10581 15728
rect 10539 15679 10581 15688
rect 10540 13712 10580 15679
rect 10636 14813 10676 23500
rect 10731 23456 10773 23465
rect 10731 23416 10732 23456
rect 10772 23416 10773 23456
rect 10731 23407 10773 23416
rect 10732 23120 10772 23407
rect 10828 23381 10868 23752
rect 10827 23372 10869 23381
rect 10827 23332 10828 23372
rect 10868 23332 10869 23372
rect 10827 23323 10869 23332
rect 10772 23080 10868 23120
rect 10732 23071 10772 23080
rect 10731 20096 10773 20105
rect 10731 20056 10732 20096
rect 10772 20056 10773 20096
rect 10731 20047 10773 20056
rect 10732 19962 10772 20047
rect 10828 18845 10868 23080
rect 10827 18836 10869 18845
rect 10827 18796 10828 18836
rect 10868 18796 10869 18836
rect 10827 18787 10869 18796
rect 10731 18332 10773 18341
rect 10731 18292 10732 18332
rect 10772 18292 10773 18332
rect 10731 18283 10773 18292
rect 10732 17758 10772 18283
rect 10924 17837 10964 23827
rect 11020 23708 11060 23920
rect 11308 23885 11348 24256
rect 11307 23876 11349 23885
rect 11307 23836 11308 23876
rect 11348 23836 11349 23876
rect 11307 23827 11349 23836
rect 11116 23792 11252 23806
rect 11116 23766 11212 23792
rect 11116 23717 11156 23766
rect 11212 23743 11252 23752
rect 11308 23742 11348 23827
rect 11015 23668 11060 23708
rect 11115 23708 11157 23717
rect 11115 23668 11116 23708
rect 11156 23668 11157 23708
rect 11404 23708 11444 25087
rect 11500 24627 11540 25171
rect 11500 24578 11540 24587
rect 11596 23792 11636 25600
rect 11692 25229 11732 25684
rect 11691 25220 11733 25229
rect 11691 25180 11692 25220
rect 11732 25180 11733 25220
rect 11691 25171 11733 25180
rect 11691 25052 11733 25061
rect 11691 25012 11692 25052
rect 11732 25012 11733 25052
rect 11691 25003 11733 25012
rect 11692 24800 11732 25003
rect 11692 24751 11732 24760
rect 11788 23960 11828 27700
rect 11980 27642 12020 27651
rect 11980 26648 12020 27602
rect 12076 27413 12116 29119
rect 12172 27749 12212 27834
rect 12171 27740 12213 27749
rect 12171 27700 12172 27740
rect 12212 27700 12213 27740
rect 12171 27691 12213 27700
rect 12075 27404 12117 27413
rect 12075 27364 12076 27404
rect 12116 27364 12117 27404
rect 12075 27355 12117 27364
rect 12076 26825 12116 27355
rect 12075 26816 12117 26825
rect 12075 26776 12076 26816
rect 12116 26776 12117 26816
rect 12075 26767 12117 26776
rect 12268 26648 12308 26657
rect 11980 26608 12268 26648
rect 12268 26599 12308 26608
rect 11979 26480 12021 26489
rect 11979 26440 11980 26480
rect 12020 26440 12021 26480
rect 11979 26431 12021 26440
rect 11883 25640 11925 25649
rect 11883 25600 11884 25640
rect 11924 25600 11925 25640
rect 11883 25591 11925 25600
rect 11884 25304 11924 25591
rect 11884 25255 11924 25264
rect 11980 23960 12020 26431
rect 12075 26144 12117 26153
rect 12075 26104 12076 26144
rect 12116 26104 12117 26144
rect 12075 26095 12117 26104
rect 12076 26010 12116 26095
rect 12364 26060 12404 31471
rect 12460 30680 12500 31555
rect 12555 31352 12597 31361
rect 12555 31312 12556 31352
rect 12596 31312 12597 31352
rect 12555 31303 12597 31312
rect 12460 30631 12500 30640
rect 12459 30260 12501 30269
rect 12459 30220 12460 30260
rect 12500 30220 12501 30260
rect 12459 30211 12501 30220
rect 12460 29681 12500 30211
rect 12459 29672 12501 29681
rect 12459 29632 12460 29672
rect 12500 29632 12501 29672
rect 12459 29623 12501 29632
rect 12460 26312 12500 29623
rect 12556 26489 12596 31303
rect 12555 26480 12597 26489
rect 12555 26440 12556 26480
rect 12596 26440 12597 26480
rect 12555 26431 12597 26440
rect 12460 26272 12596 26312
rect 12172 26020 12404 26060
rect 12460 26144 12500 26153
rect 11788 23920 11924 23960
rect 11980 23920 12116 23960
rect 11788 23792 11828 23801
rect 11596 23752 11788 23792
rect 11788 23743 11828 23752
rect 11404 23668 11636 23708
rect 11015 23540 11055 23668
rect 11115 23659 11157 23668
rect 11015 23500 11060 23540
rect 11020 22448 11060 23500
rect 11403 23288 11445 23297
rect 11403 23248 11404 23288
rect 11444 23248 11445 23288
rect 11403 23239 11445 23248
rect 11020 22408 11252 22448
rect 11020 22293 11060 22302
rect 11020 21533 11060 22253
rect 11115 21608 11157 21617
rect 11115 21568 11116 21608
rect 11156 21568 11157 21608
rect 11115 21559 11157 21568
rect 11019 21524 11061 21533
rect 11019 21484 11020 21524
rect 11060 21484 11061 21524
rect 11019 21475 11061 21484
rect 11116 21474 11156 21559
rect 11020 20768 11060 20777
rect 11020 19685 11060 20728
rect 11019 19676 11061 19685
rect 11019 19636 11020 19676
rect 11060 19636 11061 19676
rect 11019 19627 11061 19636
rect 11212 19508 11252 22408
rect 11307 21860 11349 21869
rect 11307 21820 11308 21860
rect 11348 21820 11349 21860
rect 11307 21811 11349 21820
rect 11308 21776 11348 21811
rect 11308 21725 11348 21736
rect 11020 19468 11252 19508
rect 10923 17828 10965 17837
rect 10923 17788 10924 17828
rect 10964 17788 10965 17828
rect 10923 17779 10965 17788
rect 10732 17709 10772 17718
rect 10923 17576 10965 17585
rect 10923 17536 10924 17576
rect 10964 17536 10965 17576
rect 10923 17527 10965 17536
rect 10924 17442 10964 17527
rect 11020 16409 11060 19468
rect 11115 19256 11157 19265
rect 11115 19216 11116 19256
rect 11156 19216 11157 19256
rect 11115 19207 11157 19216
rect 11116 18584 11156 19207
rect 11211 18836 11253 18845
rect 11211 18796 11212 18836
rect 11252 18796 11253 18836
rect 11211 18787 11253 18796
rect 11019 16400 11061 16409
rect 11019 16360 11020 16400
rect 11060 16360 11061 16400
rect 11019 16351 11061 16360
rect 10732 16232 10772 16241
rect 11116 16232 11156 18544
rect 11212 18173 11252 18787
rect 11307 18668 11349 18677
rect 11307 18628 11308 18668
rect 11348 18628 11349 18668
rect 11307 18619 11349 18628
rect 11308 18534 11348 18619
rect 11211 18164 11253 18173
rect 11211 18124 11212 18164
rect 11252 18124 11253 18164
rect 11211 18115 11253 18124
rect 11404 17492 11444 23239
rect 11596 23129 11636 23668
rect 11787 23624 11829 23633
rect 11787 23584 11788 23624
rect 11828 23584 11829 23624
rect 11787 23575 11829 23584
rect 11595 23120 11637 23129
rect 11595 23080 11596 23120
rect 11636 23080 11637 23120
rect 11595 23071 11637 23080
rect 11500 22285 11540 22294
rect 11500 21869 11540 22245
rect 11499 21860 11541 21869
rect 11499 21820 11500 21860
rect 11540 21820 11541 21860
rect 11499 21811 11541 21820
rect 11596 19256 11636 23071
rect 11691 22196 11733 22205
rect 11691 22156 11692 22196
rect 11732 22156 11733 22196
rect 11691 22147 11733 22156
rect 11692 22062 11732 22147
rect 11691 19928 11733 19937
rect 11691 19888 11692 19928
rect 11732 19888 11733 19928
rect 11691 19879 11733 19888
rect 11692 19517 11732 19879
rect 11691 19508 11733 19517
rect 11691 19468 11692 19508
rect 11732 19468 11733 19508
rect 11691 19459 11733 19468
rect 11308 17452 11444 17492
rect 11500 19216 11596 19256
rect 11211 17156 11253 17165
rect 11211 17116 11212 17156
rect 11252 17116 11253 17156
rect 11211 17107 11253 17116
rect 11212 17072 11252 17107
rect 11308 17072 11348 17452
rect 11404 17249 11444 17334
rect 11403 17240 11445 17249
rect 11403 17200 11404 17240
rect 11444 17200 11445 17240
rect 11403 17191 11445 17200
rect 11308 17032 11444 17072
rect 11212 17021 11252 17032
rect 10772 16192 11156 16232
rect 10732 15392 10772 16192
rect 10924 16064 10964 16073
rect 10828 16024 10924 16064
rect 10828 15560 10868 16024
rect 10924 16015 10964 16024
rect 11404 15905 11444 17032
rect 11403 15896 11445 15905
rect 11403 15856 11404 15896
rect 11444 15856 11445 15896
rect 11403 15847 11445 15856
rect 11115 15728 11157 15737
rect 11115 15688 11116 15728
rect 11156 15688 11157 15728
rect 11115 15679 11157 15688
rect 10828 15511 10868 15520
rect 10923 15560 10965 15569
rect 10923 15520 10924 15560
rect 10964 15520 10965 15560
rect 10923 15511 10965 15520
rect 10924 15426 10964 15511
rect 10732 15352 10868 15392
rect 10828 15233 10868 15352
rect 10923 15308 10965 15317
rect 10923 15268 10924 15308
rect 10964 15268 10965 15308
rect 10923 15259 10965 15268
rect 10827 15224 10869 15233
rect 10827 15184 10828 15224
rect 10868 15184 10869 15224
rect 10827 15175 10869 15184
rect 10731 15140 10773 15149
rect 10731 15100 10732 15140
rect 10772 15100 10773 15140
rect 10731 15091 10773 15100
rect 10635 14804 10677 14813
rect 10635 14764 10636 14804
rect 10676 14764 10677 14804
rect 10635 14755 10677 14764
rect 10732 14720 10772 15091
rect 10732 14561 10772 14680
rect 10731 14552 10773 14561
rect 10731 14512 10732 14552
rect 10772 14512 10773 14552
rect 10731 14503 10773 14512
rect 10540 13672 10868 13712
rect 10731 13460 10773 13469
rect 10731 13420 10732 13460
rect 10772 13420 10773 13460
rect 10731 13411 10773 13420
rect 10443 13376 10485 13385
rect 10443 13336 10444 13376
rect 10484 13336 10485 13376
rect 10443 13327 10485 13336
rect 10347 13292 10389 13301
rect 10347 13252 10348 13292
rect 10388 13252 10389 13292
rect 10347 13243 10389 13252
rect 10636 13208 10676 13217
rect 10348 13124 10388 13133
rect 10636 13124 10676 13168
rect 10732 13208 10772 13411
rect 10732 13159 10772 13168
rect 10388 13084 10676 13124
rect 10348 13075 10388 13084
rect 10731 13040 10773 13049
rect 10731 13000 10732 13040
rect 10772 13000 10773 13040
rect 10731 12991 10773 13000
rect 10443 11864 10485 11873
rect 10443 11824 10444 11864
rect 10484 11824 10485 11864
rect 10443 11815 10485 11824
rect 10252 11320 10388 11360
rect 10155 10604 10197 10613
rect 10155 10564 10156 10604
rect 10196 10564 10197 10604
rect 10155 10555 10197 10564
rect 9676 9631 9716 9640
rect 9964 9640 10100 9680
rect 9867 9596 9909 9605
rect 9964 9596 10004 9640
rect 9867 9556 9868 9596
rect 9908 9556 10004 9596
rect 9867 9547 9909 9556
rect 9868 9512 9908 9547
rect 10060 9512 10100 9521
rect 9868 9462 9908 9472
rect 9964 9470 10004 9479
rect 9964 9260 10004 9430
rect 10060 9353 10100 9472
rect 10059 9344 10101 9353
rect 10059 9304 10060 9344
rect 10100 9304 10101 9344
rect 10059 9295 10101 9304
rect 9676 9220 10004 9260
rect 9676 8765 9716 9220
rect 9772 8840 9812 8849
rect 10060 8840 10100 9295
rect 9812 8800 10100 8840
rect 10156 8840 10196 10555
rect 10252 10189 10292 10198
rect 10252 9353 10292 10149
rect 10348 10109 10388 11320
rect 10347 10100 10389 10109
rect 10347 10060 10348 10100
rect 10388 10060 10389 10100
rect 10347 10051 10389 10060
rect 10444 10100 10484 11815
rect 10444 10051 10484 10060
rect 10540 11024 10580 11033
rect 10732 11024 10772 12991
rect 10828 12536 10868 13672
rect 10828 12041 10868 12496
rect 10827 12032 10869 12041
rect 10827 11992 10828 12032
rect 10868 11992 10869 12032
rect 10827 11983 10869 11992
rect 10924 11360 10964 15259
rect 11116 14384 11156 15679
rect 11211 15644 11253 15653
rect 11211 15604 11212 15644
rect 11252 15604 11253 15644
rect 11211 15595 11253 15604
rect 11212 14972 11252 15595
rect 11403 15560 11445 15569
rect 11403 15520 11404 15560
rect 11444 15520 11445 15560
rect 11403 15511 11445 15520
rect 11308 15476 11348 15485
rect 11308 15149 11348 15436
rect 11404 15426 11444 15511
rect 11307 15140 11349 15149
rect 11307 15100 11308 15140
rect 11348 15100 11349 15140
rect 11307 15091 11349 15100
rect 11212 14932 11348 14972
rect 11116 14344 11252 14384
rect 11020 14048 11060 14059
rect 11020 13973 11060 14008
rect 11212 13973 11252 14344
rect 11019 13964 11061 13973
rect 11019 13924 11020 13964
rect 11060 13924 11061 13964
rect 11019 13915 11061 13924
rect 11211 13964 11253 13973
rect 11211 13924 11212 13964
rect 11252 13924 11253 13964
rect 11211 13915 11253 13924
rect 11212 13292 11252 13915
rect 11212 13243 11252 13252
rect 11115 13208 11157 13217
rect 11115 13168 11116 13208
rect 11156 13168 11157 13208
rect 11115 13159 11157 13168
rect 11116 13074 11156 13159
rect 11115 12788 11157 12797
rect 11115 12748 11116 12788
rect 11156 12748 11157 12788
rect 11115 12739 11157 12748
rect 10924 11320 11060 11360
rect 10580 10984 10772 11024
rect 10540 9848 10580 10984
rect 10923 10688 10965 10697
rect 10923 10648 10924 10688
rect 10964 10648 10965 10688
rect 10923 10639 10965 10648
rect 10636 10445 10676 10530
rect 10635 10436 10677 10445
rect 10635 10396 10636 10436
rect 10676 10396 10677 10436
rect 10635 10387 10677 10396
rect 10924 10361 10964 10639
rect 10923 10352 10965 10361
rect 10923 10312 10924 10352
rect 10964 10312 10965 10352
rect 10923 10303 10965 10312
rect 10444 9808 10580 9848
rect 10636 10184 10676 10193
rect 10348 9521 10388 9606
rect 10347 9512 10389 9521
rect 10347 9472 10348 9512
rect 10388 9472 10389 9512
rect 10347 9463 10389 9472
rect 10251 9344 10293 9353
rect 10251 9304 10252 9344
rect 10292 9304 10293 9344
rect 10251 9295 10293 9304
rect 10156 8800 10388 8840
rect 9772 8791 9812 8800
rect 9675 8756 9717 8765
rect 9675 8716 9676 8756
rect 9716 8716 9717 8756
rect 9675 8707 9717 8716
rect 9580 8623 9620 8632
rect 10060 8672 10100 8681
rect 9868 8168 9908 8177
rect 10060 8168 10100 8632
rect 10156 8672 10196 8681
rect 10196 8632 10292 8672
rect 10156 8623 10196 8632
rect 10155 8504 10197 8513
rect 10155 8464 10156 8504
rect 10196 8464 10197 8504
rect 10155 8455 10197 8464
rect 9908 8128 10100 8168
rect 9868 8119 9908 8128
rect 9675 8000 9717 8009
rect 9675 7960 9676 8000
rect 9716 7960 9717 8000
rect 9675 7951 9717 7960
rect 10060 8000 10100 8009
rect 9676 7866 9716 7951
rect 10060 7757 10100 7960
rect 10059 7748 10101 7757
rect 10059 7708 10060 7748
rect 10100 7708 10101 7748
rect 10059 7699 10101 7708
rect 9963 7496 10005 7505
rect 9963 7456 9964 7496
rect 10004 7456 10005 7496
rect 9963 7447 10005 7456
rect 9964 7253 10004 7447
rect 9963 7244 10005 7253
rect 9963 7204 9964 7244
rect 10004 7204 10005 7244
rect 9963 7195 10005 7204
rect 9580 7160 9620 7169
rect 9964 7160 10004 7195
rect 9620 7120 9908 7160
rect 9580 7111 9620 7120
rect 9771 6992 9813 7001
rect 9771 6952 9772 6992
rect 9812 6952 9813 6992
rect 9771 6943 9813 6952
rect 9772 6858 9812 6943
rect 9771 6488 9813 6497
rect 9771 6448 9772 6488
rect 9812 6448 9813 6488
rect 9771 6439 9813 6448
rect 9772 6354 9812 6439
rect 9579 6152 9621 6161
rect 9579 6112 9580 6152
rect 9620 6112 9621 6152
rect 9579 6103 9621 6112
rect 9580 5909 9620 6103
rect 9579 5900 9621 5909
rect 9579 5860 9580 5900
rect 9620 5860 9621 5900
rect 9579 5851 9621 5860
rect 9772 5648 9812 5657
rect 9484 5608 9772 5648
rect 9772 5599 9812 5608
rect 9772 4976 9812 4985
rect 9388 4936 9772 4976
rect 9772 4927 9812 4936
rect 9292 4852 9428 4892
rect 9099 4808 9141 4817
rect 9099 4768 9100 4808
rect 9140 4768 9141 4808
rect 9099 4759 9141 4768
rect 8811 3800 8853 3809
rect 8811 3760 8812 3800
rect 8852 3760 8853 3800
rect 8811 3751 8853 3760
rect 8332 3331 8372 3340
rect 8427 3380 8469 3389
rect 8427 3340 8428 3380
rect 8468 3340 8469 3380
rect 8427 3331 8469 3340
rect 8140 3172 8564 3212
rect 7756 3088 7988 3128
rect 7660 2792 7700 2801
rect 7275 2540 7321 2549
rect 7275 2500 7276 2540
rect 7316 2500 7321 2540
rect 7563 2540 7605 2549
rect 7563 2500 7564 2540
rect 7604 2500 7605 2540
rect 7275 2491 7317 2500
rect 7563 2491 7605 2500
rect 7563 2372 7605 2381
rect 7563 2332 7564 2372
rect 7604 2332 7605 2372
rect 7563 2323 7605 2332
rect 7275 2288 7317 2297
rect 7275 2248 7276 2288
rect 7316 2248 7317 2288
rect 7275 2239 7317 2248
rect 7179 2204 7221 2213
rect 7179 2164 7180 2204
rect 7220 2164 7221 2204
rect 7179 2155 7221 2164
rect 7180 1961 7220 2155
rect 7179 1952 7221 1961
rect 7179 1912 7180 1952
rect 7220 1912 7221 1952
rect 7179 1903 7221 1912
rect 7276 1952 7316 2239
rect 7276 1903 7316 1912
rect 7180 1818 7220 1903
rect 6988 1492 7124 1532
rect 6891 1448 6933 1457
rect 6891 1408 6892 1448
rect 6932 1408 6933 1448
rect 6891 1399 6933 1408
rect 6795 1280 6837 1289
rect 6795 1240 6796 1280
rect 6836 1240 6837 1280
rect 6795 1231 6837 1240
rect 6892 1205 6932 1399
rect 6891 1196 6933 1205
rect 6891 1156 6892 1196
rect 6932 1156 6933 1196
rect 6891 1147 6933 1156
rect 6988 1028 7028 1492
rect 7083 1280 7125 1289
rect 7083 1240 7084 1280
rect 7124 1240 7125 1280
rect 7083 1231 7125 1240
rect 7084 1037 7124 1231
rect 7564 1196 7604 2323
rect 7660 2297 7700 2752
rect 7659 2288 7701 2297
rect 7659 2248 7660 2288
rect 7700 2248 7701 2288
rect 7659 2239 7701 2248
rect 7660 1952 7700 1961
rect 7660 1793 7700 1912
rect 7756 1952 7796 3088
rect 8331 2960 8373 2969
rect 8331 2920 8332 2960
rect 8372 2920 8373 2960
rect 8331 2911 8373 2920
rect 8139 2876 8181 2885
rect 8139 2836 8140 2876
rect 8180 2836 8181 2876
rect 8139 2827 8181 2836
rect 8043 2792 8085 2801
rect 8043 2752 8044 2792
rect 8084 2752 8085 2792
rect 8043 2743 8085 2752
rect 7947 2708 7989 2717
rect 7947 2668 7948 2708
rect 7988 2668 7989 2708
rect 7947 2659 7989 2668
rect 7948 2624 7988 2659
rect 7948 2573 7988 2584
rect 8044 2624 8084 2743
rect 8044 2575 8084 2584
rect 8043 2288 8085 2297
rect 8043 2248 8044 2288
rect 8084 2248 8085 2288
rect 8043 2239 8085 2248
rect 7756 1903 7796 1912
rect 7852 1952 7892 1963
rect 7852 1877 7892 1912
rect 7948 1952 7988 1961
rect 7851 1868 7893 1877
rect 7851 1828 7852 1868
rect 7892 1828 7893 1868
rect 7851 1819 7893 1828
rect 7659 1784 7701 1793
rect 7659 1744 7660 1784
rect 7700 1744 7701 1784
rect 7659 1735 7701 1744
rect 7660 1541 7700 1735
rect 7659 1532 7701 1541
rect 7659 1492 7660 1532
rect 7700 1492 7701 1532
rect 7659 1483 7701 1492
rect 7948 1457 7988 1912
rect 8044 1793 8084 2239
rect 8140 2204 8180 2827
rect 8332 2624 8372 2911
rect 8427 2876 8469 2885
rect 8427 2836 8428 2876
rect 8468 2836 8469 2876
rect 8524 2876 8564 3172
rect 8620 3137 8660 3424
rect 8715 3380 8757 3389
rect 8715 3340 8716 3380
rect 8756 3340 8757 3380
rect 8715 3331 8757 3340
rect 8908 3380 8948 4087
rect 9004 3977 9044 4096
rect 9003 3968 9045 3977
rect 9003 3928 9004 3968
rect 9044 3928 9045 3968
rect 9003 3919 9045 3928
rect 9003 3548 9045 3557
rect 9003 3508 9004 3548
rect 9044 3508 9045 3548
rect 9003 3499 9045 3508
rect 9291 3548 9333 3557
rect 9291 3508 9292 3548
rect 9332 3508 9333 3548
rect 9291 3499 9333 3508
rect 8908 3331 8948 3340
rect 9004 3464 9044 3499
rect 8716 3246 8756 3331
rect 8811 3296 8853 3305
rect 8811 3256 8812 3296
rect 8852 3256 8853 3296
rect 8811 3247 8853 3256
rect 8812 3162 8852 3247
rect 8619 3128 8661 3137
rect 8619 3088 8620 3128
rect 8660 3088 8661 3128
rect 8619 3079 8661 3088
rect 8716 2876 8756 2885
rect 9004 2876 9044 3424
rect 9196 3464 9236 3473
rect 9099 3128 9141 3137
rect 9099 3088 9100 3128
rect 9140 3088 9141 3128
rect 9099 3079 9141 3088
rect 8524 2836 8716 2876
rect 8427 2827 8469 2836
rect 8716 2827 8756 2836
rect 8812 2836 9044 2876
rect 8428 2717 8468 2827
rect 8427 2708 8469 2717
rect 8427 2668 8428 2708
rect 8468 2668 8469 2708
rect 8427 2659 8469 2668
rect 8716 2633 8756 2718
rect 8332 2540 8372 2584
rect 8715 2624 8757 2633
rect 8715 2584 8716 2624
rect 8756 2584 8757 2624
rect 8715 2575 8757 2584
rect 8332 2500 8660 2540
rect 8140 2164 8372 2204
rect 8332 2120 8372 2164
rect 8332 2071 8372 2080
rect 8620 2120 8660 2500
rect 8716 2297 8756 2575
rect 8715 2288 8757 2297
rect 8715 2248 8716 2288
rect 8756 2248 8757 2288
rect 8715 2239 8757 2248
rect 8620 2071 8660 2080
rect 8140 1952 8180 1961
rect 8043 1784 8085 1793
rect 8043 1744 8044 1784
rect 8084 1744 8085 1784
rect 8043 1735 8085 1744
rect 7947 1448 7989 1457
rect 7947 1408 7948 1448
rect 7988 1408 7989 1448
rect 7947 1399 7989 1408
rect 8140 1373 8180 1912
rect 8235 1952 8277 1961
rect 8235 1912 8236 1952
rect 8276 1912 8277 1952
rect 8235 1903 8277 1912
rect 8428 1941 8468 1963
rect 8236 1818 8276 1903
rect 8428 1877 8468 1901
rect 8716 1952 8756 1961
rect 8427 1868 8469 1877
rect 8427 1828 8428 1868
rect 8468 1828 8469 1868
rect 8427 1819 8469 1828
rect 8427 1532 8469 1541
rect 8427 1492 8428 1532
rect 8468 1492 8469 1532
rect 8427 1483 8469 1492
rect 8139 1364 8181 1373
rect 8139 1324 8140 1364
rect 8180 1324 8181 1364
rect 8139 1315 8181 1324
rect 7755 1280 7797 1289
rect 7755 1240 7756 1280
rect 7796 1240 7797 1280
rect 7755 1231 7797 1240
rect 8331 1280 8373 1289
rect 8331 1240 8332 1280
rect 8372 1240 8373 1280
rect 8331 1231 8373 1240
rect 7660 1196 7700 1205
rect 7564 1156 7660 1196
rect 7660 1147 7700 1156
rect 7371 1112 7413 1121
rect 7371 1072 7372 1112
rect 7412 1072 7413 1112
rect 7371 1063 7413 1072
rect 7468 1103 7513 1112
rect 7468 1063 7473 1103
rect 6796 988 7028 1028
rect 7083 1028 7125 1037
rect 7083 988 7084 1028
rect 7124 988 7125 1028
rect 6796 944 6836 988
rect 7083 979 7125 988
rect 7372 978 7412 1063
rect 7468 1054 7513 1063
rect 7468 1037 7508 1054
rect 7464 1028 7508 1037
rect 7464 988 7465 1028
rect 7505 988 7508 1028
rect 7464 979 7506 988
rect 6796 895 6836 904
rect 7179 944 7221 953
rect 7179 904 7180 944
rect 7220 904 7221 944
rect 7179 895 7221 904
rect 7180 810 7220 895
rect 6700 736 6836 776
rect 6411 440 6453 449
rect 6411 400 6412 440
rect 6452 400 6453 440
rect 6411 391 6453 400
rect 6219 104 6261 113
rect 6219 80 6220 104
rect 2036 64 2056 80
rect 1976 0 2056 64
rect 2168 0 2248 80
rect 2360 0 2440 80
rect 2552 0 2632 80
rect 2744 0 2824 80
rect 2936 0 3016 80
rect 3128 0 3208 80
rect 3320 0 3400 80
rect 3512 0 3592 80
rect 3704 0 3784 80
rect 3896 0 3976 80
rect 4088 0 4168 80
rect 4280 0 4360 80
rect 4472 0 4552 80
rect 4664 0 4744 80
rect 4856 0 4936 80
rect 5048 0 5128 80
rect 5240 0 5320 80
rect 5432 0 5512 80
rect 5624 0 5704 80
rect 5816 0 5896 80
rect 6008 0 6088 80
rect 6200 64 6220 80
rect 6260 80 6261 104
rect 6412 80 6452 391
rect 6603 272 6645 281
rect 6603 232 6604 272
rect 6644 232 6645 272
rect 6603 223 6645 232
rect 6604 80 6644 223
rect 6796 80 6836 736
rect 7563 692 7605 701
rect 7563 652 7564 692
rect 7604 652 7605 692
rect 7563 643 7605 652
rect 7371 524 7413 533
rect 7371 484 7372 524
rect 7412 484 7413 524
rect 7371 475 7413 484
rect 7179 356 7221 365
rect 7179 316 7180 356
rect 7220 316 7221 356
rect 7179 307 7221 316
rect 6987 272 7029 281
rect 6987 232 6988 272
rect 7028 232 7029 272
rect 6987 223 7029 232
rect 6988 80 7028 223
rect 7180 80 7220 307
rect 7372 80 7412 475
rect 7564 80 7604 643
rect 7756 80 7796 1231
rect 8043 1196 8085 1205
rect 8043 1156 8044 1196
rect 8084 1156 8085 1196
rect 8043 1147 8085 1156
rect 8044 1062 8084 1147
rect 7852 944 7892 953
rect 7852 701 7892 904
rect 7947 944 7989 953
rect 7947 904 7948 944
rect 7988 904 7989 944
rect 7947 895 7989 904
rect 8236 944 8276 953
rect 7851 692 7893 701
rect 7851 652 7852 692
rect 7892 652 7893 692
rect 7851 643 7893 652
rect 7948 80 7988 895
rect 8139 608 8181 617
rect 8139 568 8140 608
rect 8180 568 8181 608
rect 8139 559 8181 568
rect 8140 80 8180 559
rect 8236 533 8276 904
rect 8235 524 8277 533
rect 8235 484 8236 524
rect 8276 484 8277 524
rect 8235 475 8277 484
rect 8332 80 8372 1231
rect 8428 1196 8468 1483
rect 8716 1457 8756 1912
rect 8715 1448 8757 1457
rect 8715 1408 8716 1448
rect 8756 1408 8757 1448
rect 8715 1399 8757 1408
rect 8428 1147 8468 1156
rect 8812 1196 8852 2836
rect 9100 2633 9140 3079
rect 9196 2885 9236 3424
rect 9195 2876 9237 2885
rect 9195 2836 9196 2876
rect 9236 2836 9237 2876
rect 9195 2827 9237 2836
rect 9292 2792 9332 3499
rect 9292 2743 9332 2752
rect 9004 2624 9044 2633
rect 8907 2456 8949 2465
rect 8907 2416 8908 2456
rect 8948 2416 8949 2456
rect 8907 2407 8949 2416
rect 8908 2120 8948 2407
rect 8908 2071 8948 2080
rect 9004 1961 9044 2584
rect 9099 2624 9141 2633
rect 9099 2584 9100 2624
rect 9140 2584 9141 2624
rect 9099 2575 9141 2584
rect 9388 2540 9428 4852
rect 9868 4313 9908 7120
rect 9964 7110 10004 7120
rect 9867 4304 9909 4313
rect 9867 4264 9868 4304
rect 9908 4264 9909 4304
rect 9867 4255 9909 4264
rect 10059 4304 10101 4313
rect 10059 4264 10060 4304
rect 10100 4264 10101 4304
rect 10059 4255 10101 4264
rect 9579 3968 9621 3977
rect 9579 3928 9580 3968
rect 9620 3928 9621 3968
rect 9579 3919 9621 3928
rect 9483 3380 9525 3389
rect 9483 3340 9484 3380
rect 9524 3340 9525 3380
rect 9483 3331 9525 3340
rect 9484 2876 9524 3331
rect 9484 2827 9524 2836
rect 9292 2500 9428 2540
rect 9484 2624 9524 2633
rect 9196 2456 9236 2465
rect 9003 1952 9045 1961
rect 9003 1912 9004 1952
rect 9044 1912 9045 1952
rect 9003 1903 9045 1912
rect 9196 1868 9236 2416
rect 8907 1700 8949 1709
rect 8907 1660 8908 1700
rect 8948 1660 8949 1700
rect 8907 1651 8949 1660
rect 8812 1147 8852 1156
rect 8715 1028 8757 1037
rect 8715 988 8716 1028
rect 8756 988 8757 1028
rect 8715 979 8757 988
rect 8619 944 8661 953
rect 8619 904 8620 944
rect 8660 904 8661 944
rect 8619 895 8661 904
rect 8620 810 8660 895
rect 8523 776 8565 785
rect 8523 736 8524 776
rect 8564 736 8565 776
rect 8523 727 8565 736
rect 8524 80 8564 727
rect 8716 80 8756 979
rect 8908 80 8948 1651
rect 9196 1280 9236 1828
rect 9196 1231 9236 1240
rect 9099 1196 9141 1205
rect 9099 1156 9100 1196
rect 9140 1156 9141 1196
rect 9099 1147 9141 1156
rect 9100 1037 9140 1147
rect 9099 1028 9141 1037
rect 9099 988 9100 1028
rect 9140 988 9141 1028
rect 9099 979 9141 988
rect 9004 944 9044 953
rect 9004 365 9044 904
rect 9099 860 9141 869
rect 9099 820 9100 860
rect 9140 820 9141 860
rect 9099 811 9141 820
rect 9003 356 9045 365
rect 9003 316 9004 356
rect 9044 316 9045 356
rect 9003 307 9045 316
rect 9100 80 9140 811
rect 9292 785 9332 2500
rect 9484 1961 9524 2584
rect 9483 1952 9525 1961
rect 9483 1912 9484 1952
rect 9524 1912 9525 1952
rect 9483 1903 9525 1912
rect 9388 1700 9428 1709
rect 9388 1457 9428 1660
rect 9387 1448 9429 1457
rect 9387 1408 9388 1448
rect 9428 1408 9429 1448
rect 9387 1399 9429 1408
rect 9580 1196 9620 3919
rect 10060 3893 10100 4255
rect 10059 3884 10101 3893
rect 10059 3844 10060 3884
rect 10100 3844 10101 3884
rect 10059 3835 10101 3844
rect 9963 3632 10005 3641
rect 9963 3592 9964 3632
rect 10004 3592 10005 3632
rect 9963 3583 10005 3592
rect 9867 3044 9909 3053
rect 9867 3004 9868 3044
rect 9908 3004 9909 3044
rect 9867 2995 9909 3004
rect 9676 2633 9716 2718
rect 9675 2624 9717 2633
rect 9675 2584 9676 2624
rect 9716 2584 9717 2624
rect 9675 2575 9717 2584
rect 9868 2120 9908 2995
rect 9964 2624 10004 3583
rect 10060 2708 10100 3835
rect 10156 2885 10196 8455
rect 10252 8429 10292 8632
rect 10251 8420 10293 8429
rect 10251 8380 10252 8420
rect 10292 8380 10293 8420
rect 10251 8371 10293 8380
rect 10251 6992 10293 7001
rect 10251 6952 10252 6992
rect 10292 6952 10293 6992
rect 10251 6943 10293 6952
rect 10252 6483 10292 6943
rect 10252 5662 10292 6443
rect 10252 5613 10292 5622
rect 10348 5564 10388 8800
rect 10444 8513 10484 9808
rect 10540 9680 10580 9689
rect 10636 9680 10676 10144
rect 10580 9640 10676 9680
rect 10828 10184 10868 10193
rect 10540 9631 10580 9640
rect 10636 9512 10676 9521
rect 10828 9512 10868 10144
rect 10924 10184 10964 10195
rect 10924 10109 10964 10144
rect 10923 10100 10965 10109
rect 10923 10060 10924 10100
rect 10964 10060 10965 10100
rect 10923 10051 10965 10060
rect 10540 9472 10636 9512
rect 10676 9472 10868 9512
rect 10540 9353 10580 9472
rect 10636 9463 10676 9472
rect 10539 9344 10581 9353
rect 10539 9304 10540 9344
rect 10580 9304 10581 9344
rect 10539 9295 10581 9304
rect 10635 9260 10677 9269
rect 10635 9220 10636 9260
rect 10676 9220 10677 9260
rect 10635 9211 10677 9220
rect 10539 8756 10581 8765
rect 10539 8716 10540 8756
rect 10580 8716 10581 8756
rect 10539 8707 10581 8716
rect 10636 8756 10676 9211
rect 10636 8707 10676 8716
rect 10540 8622 10580 8707
rect 10443 8504 10485 8513
rect 10443 8464 10444 8504
rect 10484 8464 10485 8504
rect 10443 8455 10485 8464
rect 10731 7832 10773 7841
rect 10731 7792 10732 7832
rect 10772 7792 10773 7832
rect 10731 7783 10773 7792
rect 10635 7748 10677 7757
rect 10635 7708 10636 7748
rect 10676 7708 10677 7748
rect 10635 7699 10677 7708
rect 10444 6572 10484 6581
rect 10484 6532 10580 6572
rect 10444 6523 10484 6532
rect 10252 5524 10388 5564
rect 10252 4733 10292 5524
rect 10444 5480 10484 5489
rect 10348 5440 10444 5480
rect 10251 4724 10293 4733
rect 10251 4684 10252 4724
rect 10292 4684 10293 4724
rect 10251 4675 10293 4684
rect 10251 4304 10293 4313
rect 10251 4264 10252 4304
rect 10292 4264 10293 4304
rect 10251 4255 10293 4264
rect 10252 4136 10292 4255
rect 10252 4087 10292 4096
rect 10348 3968 10388 5440
rect 10444 5431 10484 5440
rect 10252 3928 10388 3968
rect 10444 3968 10484 3977
rect 10155 2876 10197 2885
rect 10155 2836 10156 2876
rect 10196 2836 10197 2876
rect 10155 2827 10197 2836
rect 10060 2668 10196 2708
rect 9964 2575 10004 2584
rect 10059 2540 10101 2549
rect 10059 2500 10060 2540
rect 10100 2500 10101 2540
rect 10059 2491 10101 2500
rect 9868 2071 9908 2080
rect 9675 2036 9717 2045
rect 9675 1996 9676 2036
rect 9716 1996 9717 2036
rect 9675 1987 9717 1996
rect 9580 1147 9620 1156
rect 9483 944 9525 953
rect 9483 904 9484 944
rect 9524 904 9525 944
rect 9483 895 9525 904
rect 9291 776 9333 785
rect 9291 736 9292 776
rect 9332 736 9333 776
rect 9291 727 9333 736
rect 9291 524 9333 533
rect 9291 484 9292 524
rect 9332 484 9333 524
rect 9291 475 9333 484
rect 9292 80 9332 475
rect 9484 80 9524 895
rect 9676 80 9716 1987
rect 9771 1952 9813 1961
rect 9771 1912 9772 1952
rect 9812 1912 9813 1952
rect 9771 1903 9813 1912
rect 10060 1952 10100 2491
rect 10156 2297 10196 2668
rect 10252 2624 10292 3928
rect 10347 3800 10389 3809
rect 10347 3760 10348 3800
rect 10388 3760 10389 3800
rect 10347 3751 10389 3760
rect 10348 3464 10388 3751
rect 10444 3641 10484 3928
rect 10443 3632 10485 3641
rect 10443 3592 10444 3632
rect 10484 3592 10485 3632
rect 10443 3583 10485 3592
rect 10444 3464 10484 3473
rect 10348 3424 10444 3464
rect 10444 3415 10484 3424
rect 10252 2575 10292 2584
rect 10348 2624 10388 2633
rect 10540 2624 10580 6532
rect 10636 4229 10676 7699
rect 10732 7589 10772 7783
rect 10731 7580 10773 7589
rect 10731 7540 10732 7580
rect 10772 7540 10773 7580
rect 10731 7531 10773 7540
rect 11020 5144 11060 11320
rect 11116 9521 11156 12739
rect 11308 11360 11348 14932
rect 11403 14888 11445 14897
rect 11403 14848 11404 14888
rect 11444 14848 11445 14888
rect 11403 14839 11445 14848
rect 11212 11320 11348 11360
rect 11404 11696 11444 14839
rect 11500 12125 11540 19216
rect 11596 19207 11636 19216
rect 11788 18593 11828 23575
rect 11884 22280 11924 23920
rect 12076 23717 12116 23920
rect 12075 23708 12117 23717
rect 12075 23668 12076 23708
rect 12116 23668 12117 23708
rect 12075 23659 12117 23668
rect 12172 23456 12212 26020
rect 12268 25892 12308 25901
rect 12308 25852 12404 25892
rect 12268 25843 12308 25852
rect 12267 25640 12309 25649
rect 12267 25600 12268 25640
rect 12308 25600 12309 25640
rect 12267 25591 12309 25600
rect 12268 24977 12308 25591
rect 12364 25318 12404 25852
rect 12460 25649 12500 26104
rect 12459 25640 12501 25649
rect 12459 25600 12460 25640
rect 12500 25600 12501 25640
rect 12459 25591 12501 25600
rect 12556 25304 12596 26272
rect 12651 25388 12693 25397
rect 12651 25348 12652 25388
rect 12692 25348 12693 25388
rect 12651 25339 12693 25348
rect 12364 25269 12404 25278
rect 12460 25264 12596 25304
rect 12267 24968 12309 24977
rect 12267 24928 12268 24968
rect 12308 24928 12309 24968
rect 12267 24919 12309 24928
rect 12460 24128 12500 25264
rect 12652 25220 12692 25339
rect 12556 25180 12692 25220
rect 12556 25136 12596 25180
rect 12556 25087 12596 25096
rect 12555 24968 12597 24977
rect 12555 24928 12556 24968
rect 12596 24928 12597 24968
rect 12555 24919 12597 24928
rect 12364 24088 12500 24128
rect 12076 23416 12212 23456
rect 12268 23797 12308 23806
rect 11979 23204 12021 23213
rect 11979 23164 11980 23204
rect 12020 23164 12021 23204
rect 11979 23155 12021 23164
rect 11595 18584 11637 18593
rect 11595 18544 11596 18584
rect 11636 18544 11637 18584
rect 11595 18535 11637 18544
rect 11692 18584 11732 18593
rect 11596 18450 11636 18535
rect 11692 18248 11732 18544
rect 11787 18584 11829 18593
rect 11787 18544 11788 18584
rect 11828 18544 11829 18584
rect 11787 18535 11829 18544
rect 11787 18248 11829 18257
rect 11692 18208 11788 18248
rect 11828 18208 11829 18248
rect 11787 18199 11829 18208
rect 11691 17240 11733 17249
rect 11691 17200 11692 17240
rect 11732 17200 11733 17240
rect 11691 17191 11733 17200
rect 11692 17072 11732 17191
rect 11692 17023 11732 17032
rect 11788 17072 11828 18199
rect 11788 16484 11828 17032
rect 11692 16444 11828 16484
rect 11595 15644 11637 15653
rect 11595 15604 11596 15644
rect 11636 15604 11637 15644
rect 11595 15595 11637 15604
rect 11596 12293 11636 15595
rect 11692 13553 11732 16444
rect 11884 16400 11924 22240
rect 11980 23120 12020 23155
rect 11980 21617 12020 23080
rect 11979 21608 12021 21617
rect 11979 21568 11980 21608
rect 12020 21568 12021 21608
rect 11979 21559 12021 21568
rect 12076 20768 12116 23416
rect 12172 23288 12212 23297
rect 12268 23288 12308 23757
rect 12212 23248 12308 23288
rect 12172 23239 12212 23248
rect 12364 23120 12404 24088
rect 12268 20768 12308 20777
rect 11980 20728 12268 20768
rect 11980 20096 12020 20728
rect 12268 20719 12308 20728
rect 12172 20264 12212 20273
rect 12172 20105 12212 20224
rect 11980 18332 12020 20056
rect 12171 20096 12213 20105
rect 12171 20056 12172 20096
rect 12212 20056 12213 20096
rect 12171 20047 12213 20056
rect 12172 20045 12212 20047
rect 12364 19853 12404 23080
rect 12460 23624 12500 23633
rect 12460 22625 12500 23584
rect 12459 22616 12501 22625
rect 12459 22576 12460 22616
rect 12500 22576 12501 22616
rect 12459 22567 12501 22576
rect 12556 21953 12596 24919
rect 12651 22532 12693 22541
rect 12651 22492 12652 22532
rect 12692 22492 12693 22532
rect 12651 22483 12693 22492
rect 12652 22121 12692 22483
rect 12651 22112 12693 22121
rect 12651 22072 12652 22112
rect 12692 22072 12693 22112
rect 12651 22063 12693 22072
rect 12555 21944 12597 21953
rect 12555 21904 12556 21944
rect 12596 21904 12597 21944
rect 12555 21895 12597 21904
rect 12459 21860 12501 21869
rect 12459 21820 12460 21860
rect 12500 21820 12501 21860
rect 12459 21811 12501 21820
rect 12460 21608 12500 21811
rect 12460 21559 12500 21568
rect 12748 21440 12788 33655
rect 12844 32201 12884 36847
rect 12940 36644 12980 36653
rect 12940 34469 12980 36604
rect 13036 36644 13076 37024
rect 13036 35309 13076 36604
rect 13132 35888 13172 37192
rect 13228 36056 13268 38116
rect 13324 37820 13364 39712
rect 13516 39584 13556 40384
rect 13612 39929 13652 40972
rect 13708 40676 13748 41476
rect 13803 41264 13845 41273
rect 13803 41224 13804 41264
rect 13844 41224 13845 41264
rect 13803 41215 13845 41224
rect 13708 40627 13748 40636
rect 13707 40088 13749 40097
rect 13707 40048 13708 40088
rect 13748 40048 13749 40088
rect 13707 40039 13749 40048
rect 13611 39920 13653 39929
rect 13611 39880 13612 39920
rect 13652 39880 13653 39920
rect 13611 39871 13653 39880
rect 13516 39544 13652 39584
rect 13515 39332 13557 39341
rect 13515 39292 13516 39332
rect 13556 39292 13557 39332
rect 13515 39283 13557 39292
rect 13419 39248 13461 39257
rect 13419 39208 13420 39248
rect 13460 39208 13461 39248
rect 13419 39199 13461 39208
rect 13420 38408 13460 39199
rect 13420 38359 13460 38368
rect 13324 37780 13460 37820
rect 13420 37493 13460 37780
rect 13419 37484 13461 37493
rect 13419 37444 13420 37484
rect 13460 37444 13461 37484
rect 13419 37435 13461 37444
rect 13323 37400 13365 37409
rect 13323 37360 13324 37400
rect 13364 37360 13365 37400
rect 13323 37351 13365 37360
rect 13324 36905 13364 37351
rect 13323 36896 13365 36905
rect 13323 36856 13324 36896
rect 13364 36856 13365 36896
rect 13323 36847 13365 36856
rect 13516 36728 13556 39283
rect 13612 38921 13652 39544
rect 13611 38912 13653 38921
rect 13611 38872 13612 38912
rect 13652 38872 13653 38912
rect 13611 38863 13653 38872
rect 13611 38240 13653 38249
rect 13611 38200 13612 38240
rect 13652 38200 13653 38240
rect 13611 38191 13653 38200
rect 13612 38106 13652 38191
rect 13708 37745 13748 40039
rect 13804 38912 13844 41215
rect 13900 41105 13940 42928
rect 14092 41189 14132 42928
rect 14091 41180 14133 41189
rect 14091 41140 14092 41180
rect 14132 41140 14133 41180
rect 14091 41131 14133 41140
rect 13899 41096 13941 41105
rect 13899 41056 13900 41096
rect 13940 41056 13941 41096
rect 13899 41047 13941 41056
rect 14284 40937 14324 42928
rect 14476 41273 14516 42928
rect 14571 42524 14613 42533
rect 14571 42484 14572 42524
rect 14612 42484 14613 42524
rect 14571 42475 14613 42484
rect 14475 41264 14517 41273
rect 14475 41224 14476 41264
rect 14516 41224 14517 41264
rect 14475 41215 14517 41224
rect 14283 40928 14325 40937
rect 14283 40888 14284 40928
rect 14324 40888 14325 40928
rect 14283 40879 14325 40888
rect 14187 40844 14229 40853
rect 14187 40804 14188 40844
rect 14228 40804 14229 40844
rect 14187 40795 14229 40804
rect 14091 40592 14133 40601
rect 14091 40552 14092 40592
rect 14132 40552 14133 40592
rect 14091 40543 14133 40552
rect 13900 40508 13940 40517
rect 13900 40349 13940 40468
rect 14092 40458 14132 40543
rect 13899 40340 13941 40349
rect 13899 40300 13900 40340
rect 13940 40300 13941 40340
rect 13899 40291 13941 40300
rect 14091 40172 14133 40181
rect 14091 40132 14092 40172
rect 14132 40132 14133 40172
rect 14091 40123 14133 40132
rect 14092 39509 14132 40123
rect 14091 39500 14133 39509
rect 14091 39460 14092 39500
rect 14132 39460 14133 39500
rect 14091 39451 14133 39460
rect 13844 38872 13940 38912
rect 13804 38863 13844 38872
rect 13803 38072 13845 38081
rect 13803 38032 13804 38072
rect 13844 38032 13845 38072
rect 13803 38023 13845 38032
rect 13707 37736 13749 37745
rect 13707 37696 13708 37736
rect 13748 37696 13749 37736
rect 13707 37687 13749 37696
rect 13708 37157 13748 37687
rect 13707 37148 13749 37157
rect 13707 37108 13708 37148
rect 13748 37108 13749 37148
rect 13707 37099 13749 37108
rect 13228 36016 13364 36056
rect 13132 35839 13172 35848
rect 13228 35888 13268 35897
rect 13035 35300 13077 35309
rect 13035 35260 13036 35300
rect 13076 35260 13077 35300
rect 13035 35251 13077 35260
rect 13228 34544 13268 35848
rect 13324 34889 13364 36016
rect 13516 35225 13556 36688
rect 13612 35888 13652 35897
rect 13515 35216 13557 35225
rect 13515 35176 13516 35216
rect 13556 35176 13557 35216
rect 13515 35167 13557 35176
rect 13323 34880 13365 34889
rect 13323 34840 13324 34880
rect 13364 34840 13365 34880
rect 13323 34831 13365 34840
rect 13228 34504 13460 34544
rect 12939 34460 12981 34469
rect 12939 34420 12940 34460
rect 12980 34420 12981 34460
rect 12939 34411 12981 34420
rect 12940 33620 12980 34411
rect 13323 34376 13365 34385
rect 13323 34336 13324 34376
rect 13364 34336 13365 34376
rect 13323 34327 13365 34336
rect 13420 34376 13460 34504
rect 13227 34292 13269 34301
rect 13227 34252 13228 34292
rect 13268 34252 13269 34292
rect 13227 34243 13269 34252
rect 12940 32285 12980 33580
rect 13036 33620 13076 33631
rect 13036 33545 13076 33580
rect 13035 33536 13077 33545
rect 13035 33496 13036 33536
rect 13076 33496 13077 33536
rect 13035 33487 13077 33496
rect 13035 32780 13077 32789
rect 13035 32740 13036 32780
rect 13076 32740 13077 32780
rect 13035 32731 13077 32740
rect 12939 32276 12981 32285
rect 12939 32236 12940 32276
rect 12980 32236 12981 32276
rect 12939 32227 12981 32236
rect 12843 32192 12885 32201
rect 12843 32152 12844 32192
rect 12884 32152 12885 32192
rect 12843 32143 12885 32152
rect 12940 32108 12980 32117
rect 12843 32024 12885 32033
rect 12843 31984 12844 32024
rect 12884 31984 12885 32024
rect 12843 31975 12885 31984
rect 12844 22373 12884 31975
rect 12940 31949 12980 32068
rect 13036 32108 13076 32731
rect 13036 32033 13076 32068
rect 13035 32024 13077 32033
rect 13035 31984 13036 32024
rect 13076 31984 13077 32024
rect 13035 31975 13077 31984
rect 12939 31940 12981 31949
rect 12939 31900 12940 31940
rect 12980 31900 12981 31940
rect 12939 31891 12981 31900
rect 12940 24632 12980 31891
rect 13228 31436 13268 34243
rect 13324 34242 13364 34327
rect 13323 34124 13365 34133
rect 13323 34084 13324 34124
rect 13364 34084 13365 34124
rect 13323 34075 13365 34084
rect 13324 32864 13364 34075
rect 13420 33713 13460 34336
rect 13516 34049 13556 35167
rect 13612 34469 13652 35848
rect 13708 35888 13748 35897
rect 13708 35309 13748 35848
rect 13707 35300 13749 35309
rect 13707 35260 13708 35300
rect 13748 35260 13749 35300
rect 13707 35251 13749 35260
rect 13611 34460 13653 34469
rect 13611 34420 13612 34460
rect 13652 34420 13653 34460
rect 13611 34411 13653 34420
rect 13708 34208 13748 35251
rect 13804 34721 13844 38023
rect 13900 37577 13940 38872
rect 13996 38744 14036 38753
rect 13899 37568 13941 37577
rect 13899 37528 13900 37568
rect 13940 37528 13941 37568
rect 13899 37519 13941 37528
rect 13899 37148 13941 37157
rect 13899 37108 13900 37148
rect 13940 37108 13941 37148
rect 13899 37099 13941 37108
rect 13900 35393 13940 37099
rect 13996 36723 14036 38704
rect 13996 36674 14036 36683
rect 13899 35384 13941 35393
rect 13899 35344 13900 35384
rect 13940 35344 13941 35384
rect 13899 35335 13941 35344
rect 13900 35216 13940 35225
rect 13900 34973 13940 35176
rect 14092 35132 14132 39451
rect 14188 37157 14228 40795
rect 14475 40592 14517 40601
rect 14475 40552 14476 40592
rect 14516 40552 14517 40592
rect 14475 40543 14517 40552
rect 14283 40508 14325 40517
rect 14283 40468 14284 40508
rect 14324 40468 14325 40508
rect 14283 40459 14325 40468
rect 14284 40374 14324 40459
rect 14476 40458 14516 40543
rect 14572 40340 14612 42475
rect 14668 41768 14708 42928
rect 14668 41728 14804 41768
rect 14667 41600 14709 41609
rect 14667 41560 14668 41600
rect 14708 41560 14709 41600
rect 14667 41551 14709 41560
rect 14668 40508 14708 41551
rect 14764 40517 14804 41728
rect 14860 41693 14900 42928
rect 15052 41777 15092 42928
rect 15051 41768 15093 41777
rect 15051 41728 15052 41768
rect 15092 41728 15093 41768
rect 15051 41719 15093 41728
rect 14859 41684 14901 41693
rect 14859 41644 14860 41684
rect 14900 41644 14901 41684
rect 14859 41635 14901 41644
rect 15244 41348 15284 42928
rect 15436 42281 15476 42928
rect 15435 42272 15477 42281
rect 15435 42232 15436 42272
rect 15476 42232 15477 42272
rect 15435 42223 15477 42232
rect 15435 42104 15477 42113
rect 15435 42064 15436 42104
rect 15476 42064 15477 42104
rect 15435 42055 15477 42064
rect 15244 41308 15380 41348
rect 15052 41264 15092 41273
rect 14956 41224 15052 41264
rect 14859 40592 14901 40601
rect 14859 40552 14860 40592
rect 14900 40552 14901 40592
rect 14859 40543 14901 40552
rect 14668 40459 14708 40468
rect 14763 40508 14805 40517
rect 14763 40468 14764 40508
rect 14804 40468 14805 40508
rect 14763 40459 14805 40468
rect 14860 40458 14900 40543
rect 14572 40300 14708 40340
rect 14283 39920 14325 39929
rect 14283 39880 14284 39920
rect 14324 39880 14325 39920
rect 14283 39871 14325 39880
rect 14284 37913 14324 39871
rect 14572 39845 14612 39876
rect 14571 39836 14613 39845
rect 14571 39796 14572 39836
rect 14612 39796 14613 39836
rect 14571 39787 14613 39796
rect 14572 39752 14612 39787
rect 14476 38996 14516 39005
rect 14476 38156 14516 38956
rect 14380 38116 14516 38156
rect 14283 37904 14325 37913
rect 14283 37864 14284 37904
rect 14324 37864 14325 37904
rect 14283 37855 14325 37864
rect 14187 37148 14229 37157
rect 14187 37108 14188 37148
rect 14228 37108 14229 37148
rect 14187 37099 14229 37108
rect 14187 36812 14229 36821
rect 14187 36772 14188 36812
rect 14228 36772 14229 36812
rect 14187 36763 14229 36772
rect 14188 36678 14228 36763
rect 14188 35888 14228 35897
rect 14228 35848 14324 35888
rect 14188 35839 14228 35848
rect 14284 35309 14324 35848
rect 14283 35300 14325 35309
rect 14380 35300 14420 38116
rect 14572 37577 14612 39712
rect 14668 39080 14708 40300
rect 14956 40181 14996 41224
rect 15052 41215 15092 41224
rect 15051 41096 15093 41105
rect 15051 41056 15052 41096
rect 15092 41056 15093 41096
rect 15051 41047 15093 41056
rect 15052 40508 15092 41047
rect 15244 41012 15284 41021
rect 15052 40459 15092 40468
rect 15148 40972 15244 41012
rect 15148 40349 15188 40972
rect 15244 40963 15284 40972
rect 15243 40592 15285 40601
rect 15243 40552 15244 40592
rect 15284 40552 15285 40592
rect 15243 40543 15285 40552
rect 15244 40458 15284 40543
rect 15147 40340 15189 40349
rect 15147 40300 15148 40340
rect 15188 40300 15189 40340
rect 15147 40291 15189 40300
rect 15340 40265 15380 41308
rect 15436 41180 15476 42055
rect 15628 41180 15668 42928
rect 15820 42113 15860 42928
rect 15819 42104 15861 42113
rect 15819 42064 15820 42104
rect 15860 42064 15861 42104
rect 15819 42055 15861 42064
rect 16012 41945 16052 42928
rect 16011 41936 16053 41945
rect 16011 41896 16012 41936
rect 16052 41896 16053 41936
rect 16011 41887 16053 41896
rect 16204 41348 16244 42928
rect 16299 42188 16341 42197
rect 16299 42148 16300 42188
rect 16340 42148 16341 42188
rect 16299 42139 16341 42148
rect 16300 41441 16340 42139
rect 16396 41609 16436 42928
rect 16588 42197 16628 42928
rect 16587 42188 16629 42197
rect 16587 42148 16588 42188
rect 16628 42148 16629 42188
rect 16587 42139 16629 42148
rect 16587 41684 16629 41693
rect 16587 41644 16588 41684
rect 16628 41644 16629 41684
rect 16587 41635 16629 41644
rect 16395 41600 16437 41609
rect 16395 41560 16396 41600
rect 16436 41560 16437 41600
rect 16395 41551 16437 41560
rect 16491 41516 16533 41525
rect 16491 41476 16492 41516
rect 16532 41476 16533 41516
rect 16491 41467 16533 41476
rect 16299 41432 16341 41441
rect 16299 41392 16300 41432
rect 16340 41392 16341 41432
rect 16299 41383 16341 41392
rect 16108 41308 16244 41348
rect 15819 41180 15861 41189
rect 15628 41140 15764 41180
rect 15436 41131 15476 41140
rect 15531 41096 15573 41105
rect 15531 41056 15532 41096
rect 15572 41056 15573 41096
rect 15531 41047 15573 41056
rect 15435 40928 15477 40937
rect 15435 40888 15436 40928
rect 15476 40888 15477 40928
rect 15435 40879 15477 40888
rect 15436 40508 15476 40879
rect 15436 40459 15476 40468
rect 15339 40256 15381 40265
rect 15339 40216 15340 40256
rect 15380 40216 15381 40256
rect 15339 40207 15381 40216
rect 14955 40172 14997 40181
rect 15532 40172 15572 41047
rect 15627 41012 15669 41021
rect 15627 40972 15628 41012
rect 15668 40972 15669 41012
rect 15627 40963 15669 40972
rect 15628 40878 15668 40963
rect 15628 40592 15668 40601
rect 15628 40433 15668 40552
rect 15627 40424 15669 40433
rect 15627 40384 15628 40424
rect 15668 40384 15669 40424
rect 15627 40375 15669 40384
rect 14955 40132 14956 40172
rect 14996 40132 14997 40172
rect 14955 40123 14997 40132
rect 15436 40132 15572 40172
rect 15244 39752 15284 39761
rect 15436 39752 15476 40132
rect 15531 40004 15573 40013
rect 15531 39964 15532 40004
rect 15572 39964 15573 40004
rect 15531 39955 15573 39964
rect 15148 39712 15244 39752
rect 15284 39712 15476 39752
rect 14764 39500 14804 39509
rect 14804 39460 14996 39500
rect 14764 39451 14804 39460
rect 14668 39031 14708 39040
rect 14956 38912 14996 39460
rect 14956 38863 14996 38872
rect 15052 38912 15092 38921
rect 15052 38492 15092 38872
rect 14956 38452 15092 38492
rect 14956 38249 14996 38452
rect 14860 38240 14900 38249
rect 14571 37568 14613 37577
rect 14860 37568 14900 38200
rect 14955 38240 14997 38249
rect 14955 38200 14956 38240
rect 14996 38200 14997 38240
rect 14955 38191 14997 38200
rect 15148 38156 15188 39712
rect 15244 39703 15284 39712
rect 15532 39089 15572 39955
rect 15724 39929 15764 41140
rect 15819 41140 15820 41180
rect 15860 41140 15861 41180
rect 15819 41131 15861 41140
rect 15820 41046 15860 41131
rect 16011 41012 16053 41021
rect 16011 40972 16012 41012
rect 16052 40972 16053 41012
rect 16011 40963 16053 40972
rect 16012 40878 16052 40963
rect 16011 40592 16053 40601
rect 16011 40552 16012 40592
rect 16052 40552 16053 40592
rect 16011 40543 16053 40552
rect 15820 40508 15860 40517
rect 15723 39920 15765 39929
rect 15723 39880 15724 39920
rect 15764 39880 15765 39920
rect 15723 39871 15765 39880
rect 15531 39080 15573 39089
rect 15531 39040 15532 39080
rect 15572 39040 15573 39080
rect 15531 39031 15573 39040
rect 15532 38996 15572 39031
rect 15532 38946 15572 38956
rect 15436 38912 15476 38921
rect 15436 38417 15476 38872
rect 15627 38744 15669 38753
rect 15627 38704 15628 38744
rect 15668 38704 15669 38744
rect 15627 38695 15669 38704
rect 15435 38408 15477 38417
rect 15435 38368 15436 38408
rect 15476 38368 15477 38408
rect 15435 38359 15477 38368
rect 15340 38240 15380 38249
rect 15148 38116 15284 38156
rect 15051 38072 15093 38081
rect 15051 38032 15052 38072
rect 15092 38032 15093 38072
rect 15051 38023 15093 38032
rect 15052 37938 15092 38023
rect 15147 37904 15189 37913
rect 15147 37864 15148 37904
rect 15188 37864 15189 37904
rect 15147 37855 15189 37864
rect 15051 37820 15093 37829
rect 15051 37780 15052 37820
rect 15092 37780 15093 37820
rect 15051 37771 15093 37780
rect 14571 37528 14572 37568
rect 14612 37528 14900 37568
rect 14571 37519 14613 37528
rect 14572 37400 14612 37519
rect 14476 36644 14516 36653
rect 14476 35309 14516 36604
rect 14572 35981 14612 37360
rect 14859 37316 14901 37325
rect 14859 37276 14860 37316
rect 14900 37276 14901 37316
rect 14859 37267 14901 37276
rect 14764 37232 14804 37241
rect 14667 36896 14709 36905
rect 14667 36856 14668 36896
rect 14708 36856 14709 36896
rect 14667 36847 14709 36856
rect 14668 36762 14708 36847
rect 14571 35972 14613 35981
rect 14764 35972 14804 37192
rect 14860 36644 14900 37267
rect 14955 36896 14997 36905
rect 14955 36856 14956 36896
rect 14996 36856 14997 36896
rect 14955 36847 14997 36856
rect 15052 36896 15092 37771
rect 15148 37745 15188 37855
rect 15244 37829 15284 38116
rect 15340 38081 15380 38200
rect 15435 38240 15477 38249
rect 15435 38200 15436 38240
rect 15476 38200 15477 38240
rect 15435 38191 15477 38200
rect 15339 38072 15381 38081
rect 15339 38032 15340 38072
rect 15380 38032 15381 38072
rect 15339 38023 15381 38032
rect 15243 37820 15285 37829
rect 15243 37780 15244 37820
rect 15284 37780 15285 37820
rect 15436 37820 15476 38191
rect 15628 37913 15668 38695
rect 15820 38576 15860 40468
rect 16012 40458 16052 40543
rect 15915 39080 15957 39089
rect 15915 39040 15916 39080
rect 15956 39040 15957 39080
rect 15915 39031 15957 39040
rect 15724 38536 15860 38576
rect 15627 37904 15669 37913
rect 15627 37864 15628 37904
rect 15668 37864 15669 37904
rect 15627 37855 15669 37864
rect 15436 37780 15572 37820
rect 15243 37771 15285 37780
rect 15147 37736 15189 37745
rect 15147 37696 15148 37736
rect 15188 37696 15189 37736
rect 15147 37687 15189 37696
rect 15052 36847 15092 36856
rect 14956 36728 14996 36847
rect 14956 36688 15092 36728
rect 14860 36595 14900 36604
rect 14955 36560 14997 36569
rect 14955 36520 14956 36560
rect 14996 36520 14997 36560
rect 14955 36511 14997 36520
rect 14571 35932 14572 35972
rect 14612 35932 14613 35972
rect 14571 35923 14613 35932
rect 14716 35932 14804 35972
rect 14956 35972 14996 36511
rect 15052 36140 15092 36688
rect 15052 36091 15092 36100
rect 14956 35932 15092 35972
rect 14716 35930 14756 35932
rect 14283 35260 14284 35300
rect 14324 35260 14325 35300
rect 14283 35251 14325 35260
rect 14379 35260 14420 35300
rect 14475 35300 14517 35309
rect 14475 35260 14476 35300
rect 14516 35260 14517 35300
rect 14379 35216 14419 35260
rect 14475 35251 14517 35260
rect 14379 35176 14420 35216
rect 13996 35092 14132 35132
rect 13899 34964 13941 34973
rect 13899 34924 13900 34964
rect 13940 34924 13941 34964
rect 13899 34915 13941 34924
rect 13803 34712 13845 34721
rect 13803 34672 13804 34712
rect 13844 34672 13845 34712
rect 13803 34663 13845 34672
rect 13803 34460 13845 34469
rect 13803 34420 13804 34460
rect 13844 34420 13845 34460
rect 13803 34411 13845 34420
rect 13804 34326 13844 34411
rect 13900 34376 13940 34385
rect 13900 34208 13940 34336
rect 13708 34168 13940 34208
rect 13515 34040 13557 34049
rect 13515 34000 13516 34040
rect 13556 34000 13557 34040
rect 13515 33991 13557 34000
rect 13419 33704 13461 33713
rect 13419 33664 13420 33704
rect 13460 33664 13461 33704
rect 13419 33655 13461 33664
rect 13516 33704 13556 33991
rect 13516 33655 13556 33664
rect 13804 33545 13844 34168
rect 13996 33788 14036 35092
rect 13900 33748 14036 33788
rect 14092 34964 14132 34973
rect 13419 33536 13461 33545
rect 13419 33496 13420 33536
rect 13460 33496 13461 33536
rect 13419 33487 13461 33496
rect 13803 33536 13845 33545
rect 13803 33496 13804 33536
rect 13844 33496 13845 33536
rect 13803 33487 13845 33496
rect 13324 31613 13364 32824
rect 13420 32024 13460 33487
rect 13515 33452 13557 33461
rect 13515 33412 13516 33452
rect 13556 33412 13557 33452
rect 13515 33403 13557 33412
rect 13516 32192 13556 33403
rect 13516 32143 13556 32152
rect 13420 31984 13556 32024
rect 13323 31604 13365 31613
rect 13323 31564 13324 31604
rect 13364 31564 13365 31604
rect 13323 31555 13365 31564
rect 13228 31396 13364 31436
rect 13228 29177 13268 29262
rect 13227 29168 13269 29177
rect 13227 29128 13228 29168
rect 13268 29128 13269 29168
rect 13227 29119 13269 29128
rect 13324 29000 13364 31396
rect 13228 28960 13364 29000
rect 13035 27656 13077 27665
rect 13035 27616 13036 27656
rect 13076 27616 13077 27656
rect 13035 27607 13077 27616
rect 13036 27522 13076 27607
rect 13131 26984 13173 26993
rect 13131 26944 13132 26984
rect 13172 26944 13173 26984
rect 13131 26935 13173 26944
rect 12940 24592 13076 24632
rect 12939 22700 12981 22709
rect 12939 22660 12940 22700
rect 12980 22660 12981 22700
rect 12939 22651 12981 22660
rect 12843 22364 12885 22373
rect 12843 22324 12844 22364
rect 12884 22324 12885 22364
rect 12843 22315 12885 22324
rect 12843 22112 12885 22121
rect 12843 22072 12844 22112
rect 12884 22072 12885 22112
rect 12843 22063 12885 22072
rect 12844 21608 12884 22063
rect 12940 21869 12980 22651
rect 12939 21860 12981 21869
rect 12939 21820 12940 21860
rect 12980 21820 12981 21860
rect 12939 21811 12981 21820
rect 12844 21559 12884 21568
rect 12940 21608 12980 21617
rect 12940 21440 12980 21568
rect 12748 21400 12980 21440
rect 12556 21356 12596 21365
rect 12460 20693 12500 20724
rect 12459 20684 12501 20693
rect 12459 20644 12460 20684
rect 12500 20644 12501 20684
rect 12459 20635 12501 20644
rect 12460 20600 12500 20635
rect 12460 20105 12500 20560
rect 12455 20096 12500 20105
rect 12495 20056 12500 20096
rect 12455 20047 12500 20056
rect 12556 20096 12596 21316
rect 12748 20777 12788 21400
rect 12652 20768 12692 20777
rect 12747 20768 12789 20777
rect 12692 20728 12748 20768
rect 12788 20728 12789 20768
rect 12652 20719 12692 20728
rect 12747 20719 12789 20728
rect 12844 20768 12884 20777
rect 12748 20600 12788 20609
rect 12556 20047 12596 20056
rect 12652 20096 12692 20107
rect 12748 20105 12788 20560
rect 12844 20189 12884 20728
rect 12940 20768 12980 20779
rect 12940 20693 12980 20728
rect 12939 20684 12981 20693
rect 12939 20644 12940 20684
rect 12980 20644 12981 20684
rect 12939 20635 12981 20644
rect 12843 20180 12885 20189
rect 12843 20140 12844 20180
rect 12884 20140 12885 20180
rect 12843 20131 12885 20140
rect 12363 19844 12405 19853
rect 12363 19804 12364 19844
rect 12404 19804 12405 19844
rect 12363 19795 12405 19804
rect 12460 19181 12500 20047
rect 12652 20021 12692 20056
rect 12747 20096 12789 20105
rect 12747 20056 12748 20096
rect 12788 20056 12789 20096
rect 12747 20047 12789 20056
rect 12844 20096 12884 20131
rect 12844 20047 12884 20056
rect 12939 20096 12981 20105
rect 12939 20056 12940 20096
rect 12980 20056 12981 20096
rect 12939 20047 12981 20056
rect 12651 20012 12693 20021
rect 12651 19972 12652 20012
rect 12692 19972 12693 20012
rect 12651 19963 12693 19972
rect 12940 19962 12980 20047
rect 12940 19844 12980 19853
rect 12652 19804 12940 19844
rect 12459 19172 12501 19181
rect 12459 19132 12460 19172
rect 12500 19132 12501 19172
rect 12459 19123 12501 19132
rect 12076 18628 12404 18668
rect 12076 18584 12116 18628
rect 12076 18535 12116 18544
rect 12172 18500 12212 18509
rect 11980 18292 12116 18332
rect 11979 16736 12021 16745
rect 11979 16696 11980 16736
rect 12020 16696 12021 16736
rect 11979 16687 12021 16696
rect 11788 16360 11924 16400
rect 11691 13544 11733 13553
rect 11691 13504 11692 13544
rect 11732 13504 11733 13544
rect 11691 13495 11733 13504
rect 11691 13376 11733 13385
rect 11691 13336 11692 13376
rect 11732 13336 11733 13376
rect 11691 13327 11733 13336
rect 11692 13207 11732 13327
rect 11692 13158 11732 13167
rect 11788 13040 11828 16360
rect 11884 16232 11924 16241
rect 11980 16232 12020 16687
rect 11924 16192 12020 16232
rect 11884 16183 11924 16192
rect 12076 15989 12116 18292
rect 12172 17660 12212 18460
rect 12172 17620 12308 17660
rect 12172 16988 12212 16997
rect 12172 16325 12212 16948
rect 12268 16988 12308 17620
rect 12268 16661 12308 16948
rect 12267 16652 12309 16661
rect 12267 16612 12268 16652
rect 12308 16612 12309 16652
rect 12267 16603 12309 16612
rect 12171 16316 12213 16325
rect 12171 16276 12172 16316
rect 12212 16276 12213 16316
rect 12171 16267 12213 16276
rect 12075 15980 12117 15989
rect 12075 15940 12076 15980
rect 12116 15940 12117 15980
rect 12075 15931 12117 15940
rect 11883 15896 11925 15905
rect 11883 15856 11884 15896
rect 11924 15856 11925 15896
rect 11883 15847 11925 15856
rect 11884 15560 11924 15847
rect 12172 15728 12212 16267
rect 12364 15737 12404 18628
rect 12652 18584 12692 19804
rect 12940 19795 12980 19804
rect 13036 19424 13076 24592
rect 13132 22541 13172 26935
rect 13228 26825 13268 28960
rect 13420 28916 13460 28925
rect 13324 28876 13420 28916
rect 13324 28328 13364 28876
rect 13420 28867 13460 28876
rect 13324 28279 13364 28288
rect 13419 28328 13461 28337
rect 13419 28288 13420 28328
rect 13460 28288 13461 28328
rect 13419 28279 13461 28288
rect 13420 28194 13460 28279
rect 13227 26816 13269 26825
rect 13227 26776 13228 26816
rect 13268 26776 13269 26816
rect 13227 26767 13269 26776
rect 13516 26228 13556 31984
rect 13803 31520 13845 31529
rect 13803 31480 13804 31520
rect 13844 31480 13845 31520
rect 13803 31471 13845 31480
rect 13804 31352 13844 31471
rect 13804 31303 13844 31312
rect 13707 30764 13749 30773
rect 13707 30724 13708 30764
rect 13748 30724 13749 30764
rect 13707 30715 13749 30724
rect 13611 30680 13653 30689
rect 13611 30640 13612 30680
rect 13652 30640 13653 30680
rect 13611 30631 13653 30640
rect 13708 30680 13748 30715
rect 13612 29168 13652 30631
rect 13708 30629 13748 30640
rect 13900 30596 13940 33748
rect 14092 33704 14132 34924
rect 14284 34964 14324 34973
rect 14284 34469 14324 34924
rect 14380 34889 14420 35176
rect 14476 35174 14516 35183
rect 14572 35174 14612 35923
rect 14716 35881 14756 35890
rect 14860 35720 14900 35729
rect 14900 35680 14996 35720
rect 14860 35671 14900 35680
rect 14667 35384 14709 35393
rect 14667 35344 14668 35384
rect 14708 35344 14709 35384
rect 14667 35335 14709 35344
rect 14516 35134 14612 35174
rect 14476 35125 14516 35134
rect 14379 34880 14421 34889
rect 14379 34840 14380 34880
rect 14420 34840 14421 34880
rect 14379 34831 14421 34840
rect 14283 34460 14325 34469
rect 14283 34420 14284 34460
rect 14324 34420 14325 34460
rect 14283 34411 14325 34420
rect 14380 34376 14420 34385
rect 14380 34049 14420 34336
rect 14379 34040 14421 34049
rect 14379 34000 14380 34040
rect 14420 34000 14421 34040
rect 14379 33991 14421 34000
rect 14188 33788 14228 33799
rect 14188 33713 14228 33748
rect 14044 33694 14132 33704
rect 14084 33664 14132 33694
rect 14187 33704 14229 33713
rect 14187 33664 14188 33704
rect 14228 33664 14229 33704
rect 14187 33655 14229 33664
rect 14475 33704 14517 33713
rect 14475 33664 14476 33704
rect 14516 33664 14517 33704
rect 14475 33655 14517 33664
rect 14044 33645 14084 33654
rect 14476 32696 14516 33655
rect 14668 33125 14708 35335
rect 14956 35309 14996 35680
rect 14955 35300 14997 35309
rect 14955 35260 14956 35300
rect 14996 35260 14997 35300
rect 14955 35251 14997 35260
rect 14763 34712 14805 34721
rect 14763 34672 14764 34712
rect 14804 34672 14805 34712
rect 14763 34663 14805 34672
rect 14764 34292 14804 34663
rect 14860 34469 14900 34485
rect 14859 34460 14901 34469
rect 14859 34420 14860 34460
rect 14900 34420 14901 34460
rect 14859 34411 14901 34420
rect 14860 34390 14900 34411
rect 14860 34341 14900 34350
rect 14764 34252 14900 34292
rect 14667 33116 14709 33125
rect 14667 33076 14668 33116
rect 14708 33076 14709 33116
rect 14667 33067 14709 33076
rect 14572 32873 14612 32958
rect 14667 32948 14709 32957
rect 14667 32908 14668 32948
rect 14708 32908 14709 32948
rect 14667 32899 14709 32908
rect 14571 32864 14613 32873
rect 14571 32824 14572 32864
rect 14612 32824 14613 32864
rect 14571 32815 14613 32824
rect 14476 32656 14612 32696
rect 14188 32276 14228 32285
rect 14188 32201 14228 32236
rect 14187 32192 14229 32201
rect 13996 32178 14036 32187
rect 14187 32152 14188 32192
rect 14228 32152 14229 32192
rect 14187 32143 14229 32152
rect 13996 31604 14036 32138
rect 13996 31555 14036 31564
rect 14091 31352 14133 31361
rect 14091 31312 14092 31352
rect 14132 31312 14133 31352
rect 14091 31303 14133 31312
rect 14092 30680 14132 31303
rect 14188 30932 14228 32143
rect 14572 31100 14612 32656
rect 14668 31277 14708 32899
rect 14860 32705 14900 34252
rect 14956 34217 14996 35251
rect 15052 34721 15092 35932
rect 15051 34712 15093 34721
rect 15051 34672 15052 34712
rect 15092 34672 15093 34712
rect 15051 34663 15093 34672
rect 15148 34376 15188 37687
rect 15435 37652 15477 37661
rect 15435 37612 15436 37652
rect 15476 37612 15477 37652
rect 15435 37603 15477 37612
rect 15436 37518 15476 37603
rect 15244 37484 15284 37493
rect 15244 37241 15284 37444
rect 15243 37232 15285 37241
rect 15243 37192 15244 37232
rect 15284 37192 15285 37232
rect 15243 37183 15285 37192
rect 15339 36896 15381 36905
rect 15339 36856 15340 36896
rect 15380 36856 15381 36896
rect 15339 36847 15381 36856
rect 15340 36728 15380 36847
rect 15532 36812 15572 37780
rect 15628 37400 15668 37409
rect 15628 37073 15668 37360
rect 15627 37064 15669 37073
rect 15627 37024 15628 37064
rect 15668 37024 15669 37064
rect 15627 37015 15669 37024
rect 15340 36679 15380 36688
rect 15436 36772 15572 36812
rect 15436 36728 15476 36772
rect 15436 36569 15476 36688
rect 15531 36644 15573 36653
rect 15531 36604 15532 36644
rect 15572 36604 15573 36644
rect 15531 36595 15573 36604
rect 15435 36560 15477 36569
rect 15435 36520 15436 36560
rect 15476 36520 15477 36560
rect 15435 36511 15477 36520
rect 15435 36392 15477 36401
rect 15435 36352 15436 36392
rect 15476 36352 15477 36392
rect 15435 36343 15477 36352
rect 15243 35972 15285 35981
rect 15243 35932 15244 35972
rect 15284 35932 15285 35972
rect 15243 35923 15285 35932
rect 15244 35888 15284 35923
rect 15244 35837 15284 35848
rect 15244 34376 15284 34385
rect 15148 34336 15244 34376
rect 15244 34327 15284 34336
rect 14955 34208 14997 34217
rect 14955 34168 14956 34208
rect 14996 34168 14997 34208
rect 14955 34159 14997 34168
rect 15052 34208 15092 34217
rect 15052 33965 15092 34168
rect 15147 34208 15189 34217
rect 15147 34168 15148 34208
rect 15188 34168 15189 34208
rect 15147 34159 15189 34168
rect 15051 33956 15093 33965
rect 15051 33916 15052 33956
rect 15092 33916 15093 33956
rect 15051 33907 15093 33916
rect 14764 32696 14804 32705
rect 14764 32192 14804 32656
rect 14859 32696 14901 32705
rect 14859 32656 14860 32696
rect 14900 32656 14901 32696
rect 14859 32647 14901 32656
rect 14764 32143 14804 32152
rect 14860 32192 14900 32203
rect 14860 32117 14900 32152
rect 14859 32108 14901 32117
rect 14859 32068 14860 32108
rect 14900 32068 14901 32108
rect 14859 32059 14901 32068
rect 14859 31352 14901 31361
rect 14859 31312 14860 31352
rect 14900 31312 14901 31352
rect 14859 31303 14901 31312
rect 14667 31268 14709 31277
rect 14667 31228 14668 31268
rect 14708 31228 14709 31268
rect 14667 31219 14709 31228
rect 14860 31218 14900 31303
rect 14572 31060 14708 31100
rect 14188 30892 14516 30932
rect 14187 30764 14229 30773
rect 14187 30724 14188 30764
rect 14228 30724 14229 30764
rect 14187 30715 14229 30724
rect 14092 30631 14132 30640
rect 13900 30556 14036 30596
rect 13996 30512 14036 30556
rect 13996 30472 14132 30512
rect 13900 30428 13940 30437
rect 13900 29840 13940 30388
rect 13900 29791 13940 29800
rect 13995 29840 14037 29849
rect 13995 29800 13996 29840
rect 14036 29800 14037 29840
rect 13995 29791 14037 29800
rect 13996 29588 14036 29791
rect 13804 29548 14036 29588
rect 13804 29261 13844 29548
rect 13899 29420 13941 29429
rect 13899 29380 13900 29420
rect 13940 29380 13941 29420
rect 13899 29371 13941 29380
rect 13803 29252 13845 29261
rect 13803 29212 13804 29252
rect 13844 29212 13845 29252
rect 13803 29203 13845 29212
rect 13612 26993 13652 29128
rect 13900 29000 13940 29371
rect 13995 29168 14037 29177
rect 13995 29128 13996 29168
rect 14036 29128 14037 29168
rect 13995 29119 14037 29128
rect 13996 29009 14036 29119
rect 13804 28960 13940 29000
rect 13995 29000 14037 29009
rect 13995 28960 13996 29000
rect 14036 28960 14037 29000
rect 13804 28328 13844 28960
rect 13995 28951 14037 28960
rect 13899 28496 13941 28505
rect 13899 28456 13900 28496
rect 13940 28456 13941 28496
rect 13899 28447 13941 28456
rect 13900 28412 13940 28447
rect 13900 28361 13940 28372
rect 13611 26984 13653 26993
rect 13611 26944 13612 26984
rect 13652 26944 13653 26984
rect 13611 26935 13653 26944
rect 13611 26816 13653 26825
rect 13611 26776 13612 26816
rect 13652 26776 13653 26816
rect 13611 26767 13653 26776
rect 13228 26188 13556 26228
rect 13228 22709 13268 26188
rect 13515 26060 13557 26069
rect 13515 26020 13516 26060
rect 13556 26020 13557 26060
rect 13515 26011 13557 26020
rect 13516 22952 13556 26011
rect 13612 24212 13652 26767
rect 13707 26144 13749 26153
rect 13707 26104 13708 26144
rect 13748 26104 13749 26144
rect 13707 26095 13749 26104
rect 13708 26010 13748 26095
rect 13804 26069 13844 28288
rect 13996 27824 14036 28951
rect 13900 27784 14036 27824
rect 13900 26405 13940 27784
rect 13995 27656 14037 27665
rect 14092 27656 14132 30472
rect 13995 27616 13996 27656
rect 14036 27616 14132 27656
rect 14188 27656 14228 30715
rect 14380 29840 14420 29849
rect 14380 29429 14420 29800
rect 14476 29840 14516 30892
rect 14379 29420 14421 29429
rect 14379 29380 14380 29420
rect 14420 29380 14421 29420
rect 14379 29371 14421 29380
rect 14379 28832 14421 28841
rect 14379 28792 14380 28832
rect 14420 28792 14421 28832
rect 14379 28783 14421 28792
rect 14380 28328 14420 28783
rect 14380 28279 14420 28288
rect 14476 27824 14516 29800
rect 14380 27784 14516 27824
rect 14668 27824 14708 31060
rect 14763 30596 14805 30605
rect 14763 30556 14764 30596
rect 14804 30556 14805 30596
rect 14763 30547 14805 30556
rect 14764 28244 14804 30547
rect 14955 30260 14997 30269
rect 14955 30220 14956 30260
rect 14996 30220 14997 30260
rect 14955 30211 14997 30220
rect 14956 30101 14996 30211
rect 14955 30092 14997 30101
rect 14955 30052 14956 30092
rect 14996 30052 14997 30092
rect 14955 30043 14997 30052
rect 14956 29840 14996 30043
rect 14956 29791 14996 29800
rect 14859 29420 14901 29429
rect 14859 29380 14860 29420
rect 14900 29380 14901 29420
rect 14859 29371 14901 29380
rect 14860 29168 14900 29371
rect 14860 29093 14900 29128
rect 14859 29084 14901 29093
rect 14859 29044 14860 29084
rect 14900 29044 14901 29084
rect 14859 29035 14901 29044
rect 14860 29004 14900 29035
rect 15052 28916 15092 28925
rect 14908 28370 14948 28379
rect 15052 28370 15092 28876
rect 14948 28330 15092 28370
rect 14908 28321 14948 28330
rect 15052 28244 15092 28253
rect 14764 28204 15052 28244
rect 15052 28195 15092 28204
rect 14668 27784 14996 27824
rect 14284 27656 14324 27665
rect 14188 27616 14284 27656
rect 13995 27607 14037 27616
rect 13899 26396 13941 26405
rect 13899 26356 13900 26396
rect 13940 26356 13941 26396
rect 13899 26347 13941 26356
rect 13900 26153 13940 26347
rect 13899 26144 13941 26153
rect 13899 26104 13900 26144
rect 13940 26104 13941 26144
rect 13899 26095 13941 26104
rect 13803 26060 13845 26069
rect 13803 26020 13804 26060
rect 13844 26020 13845 26060
rect 13803 26011 13845 26020
rect 13900 25892 13940 25901
rect 13708 25852 13900 25892
rect 13708 25304 13748 25852
rect 13900 25843 13940 25852
rect 13803 25472 13845 25481
rect 13803 25432 13804 25472
rect 13844 25432 13845 25472
rect 13803 25423 13845 25432
rect 13708 25255 13748 25264
rect 13804 25304 13844 25423
rect 13804 25255 13844 25264
rect 13900 24632 13940 24641
rect 13996 24632 14036 27607
rect 14284 27413 14324 27616
rect 14283 27404 14325 27413
rect 14283 27364 14284 27404
rect 14324 27364 14325 27404
rect 14283 27355 14325 27364
rect 14283 26984 14325 26993
rect 14283 26944 14284 26984
rect 14324 26944 14325 26984
rect 14283 26935 14325 26944
rect 14187 25304 14229 25313
rect 14187 25264 14188 25304
rect 14228 25264 14229 25304
rect 14187 25255 14229 25264
rect 14284 25304 14324 26935
rect 14188 25170 14228 25255
rect 14284 25229 14324 25264
rect 14283 25220 14325 25229
rect 14283 25180 14284 25220
rect 14324 25180 14325 25220
rect 14283 25171 14325 25180
rect 13940 24592 14036 24632
rect 13900 24583 13940 24592
rect 13612 24172 13748 24212
rect 13611 23204 13653 23213
rect 13611 23164 13612 23204
rect 13652 23164 13653 23204
rect 13611 23155 13653 23164
rect 13612 23120 13652 23155
rect 13612 23069 13652 23080
rect 13516 22912 13652 22952
rect 13227 22700 13269 22709
rect 13227 22660 13228 22700
rect 13268 22660 13269 22700
rect 13227 22651 13269 22660
rect 13131 22532 13173 22541
rect 13131 22492 13132 22532
rect 13172 22492 13173 22532
rect 13131 22483 13173 22492
rect 13515 22532 13557 22541
rect 13515 22492 13516 22532
rect 13556 22492 13557 22532
rect 13515 22483 13557 22492
rect 13131 22280 13173 22289
rect 13131 22240 13132 22280
rect 13172 22240 13173 22280
rect 13131 22231 13173 22240
rect 13516 22280 13556 22483
rect 13516 22231 13556 22240
rect 13132 22146 13172 22231
rect 13323 22112 13365 22121
rect 13323 22072 13324 22112
rect 13364 22072 13365 22112
rect 13323 22063 13365 22072
rect 13324 21978 13364 22063
rect 13323 21860 13365 21869
rect 13323 21820 13324 21860
rect 13364 21820 13365 21860
rect 13323 21811 13365 21820
rect 13324 21608 13364 21811
rect 13419 21692 13461 21701
rect 13419 21652 13420 21692
rect 13460 21652 13461 21692
rect 13419 21643 13461 21652
rect 13324 21559 13364 21568
rect 13420 21608 13460 21643
rect 13420 21557 13460 21568
rect 13227 20852 13269 20861
rect 13132 20812 13228 20852
rect 13268 20812 13269 20852
rect 13132 20768 13172 20812
rect 13227 20803 13269 20812
rect 13132 20719 13172 20728
rect 13419 20012 13461 20021
rect 13419 19972 13420 20012
rect 13460 19972 13461 20012
rect 13419 19963 13461 19972
rect 12459 18416 12501 18425
rect 12459 18376 12460 18416
rect 12500 18376 12501 18416
rect 12459 18367 12501 18376
rect 11884 15511 11924 15520
rect 11980 15688 12212 15728
rect 12363 15728 12405 15737
rect 12363 15688 12364 15728
rect 12404 15688 12405 15728
rect 11980 15392 12020 15688
rect 12363 15679 12405 15688
rect 11692 13000 11828 13040
rect 11884 15352 12020 15392
rect 12364 15546 12404 15555
rect 11595 12284 11637 12293
rect 11595 12244 11596 12284
rect 11636 12244 11637 12284
rect 11595 12235 11637 12244
rect 11499 12116 11541 12125
rect 11499 12076 11500 12116
rect 11540 12076 11541 12116
rect 11499 12067 11541 12076
rect 11596 12041 11636 12235
rect 11595 12032 11637 12041
rect 11595 11992 11596 12032
rect 11636 11992 11637 12032
rect 11595 11983 11637 11992
rect 11404 11360 11444 11656
rect 11596 11528 11636 11537
rect 11404 11320 11540 11360
rect 11115 9512 11157 9521
rect 11115 9472 11116 9512
rect 11156 9472 11157 9512
rect 11115 9463 11157 9472
rect 11212 9512 11252 11320
rect 11307 10604 11349 10613
rect 11307 10564 11308 10604
rect 11348 10564 11349 10604
rect 11307 10555 11349 10564
rect 11308 10277 11348 10555
rect 11403 10520 11445 10529
rect 11403 10480 11404 10520
rect 11444 10480 11445 10520
rect 11403 10471 11445 10480
rect 11307 10268 11349 10277
rect 11307 10228 11308 10268
rect 11348 10228 11349 10268
rect 11307 10219 11349 10228
rect 11404 10193 11444 10471
rect 11403 10184 11445 10193
rect 11403 10144 11404 10184
rect 11444 10144 11445 10184
rect 11403 10135 11445 10144
rect 11404 10050 11444 10135
rect 11500 10109 11540 11320
rect 11596 11033 11636 11488
rect 11595 11024 11637 11033
rect 11595 10984 11596 11024
rect 11636 10984 11637 11024
rect 11595 10975 11637 10984
rect 11499 10100 11541 10109
rect 11499 10060 11500 10100
rect 11540 10060 11541 10100
rect 11499 10051 11541 10060
rect 11115 9344 11157 9353
rect 11115 9304 11116 9344
rect 11156 9304 11157 9344
rect 11115 9295 11157 9304
rect 11116 8672 11156 9295
rect 11116 8623 11156 8632
rect 11212 8345 11252 9472
rect 11596 8677 11636 8686
rect 11211 8336 11253 8345
rect 11211 8296 11212 8336
rect 11252 8296 11253 8336
rect 11211 8287 11253 8296
rect 11500 8168 11540 8177
rect 11596 8168 11636 8637
rect 11540 8128 11636 8168
rect 11500 8119 11540 8128
rect 11692 8009 11732 13000
rect 11787 12116 11829 12125
rect 11787 12076 11788 12116
rect 11828 12076 11829 12116
rect 11787 12067 11829 12076
rect 11788 11537 11828 12067
rect 11884 11873 11924 15352
rect 11979 15224 12021 15233
rect 11979 15184 11980 15224
rect 12020 15184 12021 15224
rect 11979 15175 12021 15184
rect 11980 14720 12020 15175
rect 12172 14972 12212 14981
rect 12364 14972 12404 15506
rect 12460 14981 12500 18367
rect 12652 17072 12692 18544
rect 12748 19384 13076 19424
rect 12748 17240 12788 19384
rect 13228 19266 13268 19275
rect 12843 19256 12885 19265
rect 12843 19216 12844 19256
rect 12884 19216 12885 19256
rect 12843 19207 12885 19216
rect 13131 19247 13228 19256
rect 13131 19207 13132 19247
rect 13172 19226 13228 19247
rect 13324 19265 13364 19350
rect 13172 19216 13268 19226
rect 13323 19256 13365 19265
rect 13323 19216 13324 19256
rect 13364 19216 13365 19256
rect 13172 19207 13173 19216
rect 13323 19207 13365 19216
rect 12844 19122 12884 19207
rect 13131 19198 13173 19207
rect 12939 19088 12981 19097
rect 12939 19048 12940 19088
rect 12980 19048 12981 19088
rect 12939 19039 12981 19048
rect 13036 19088 13076 19097
rect 13227 19088 13269 19097
rect 13076 19048 13172 19088
rect 13036 19039 13076 19048
rect 12748 17200 12884 17240
rect 12748 17072 12788 17081
rect 12652 17032 12748 17072
rect 12748 17023 12788 17032
rect 12556 15728 12596 15737
rect 12651 15728 12693 15737
rect 12596 15688 12652 15728
rect 12692 15688 12693 15728
rect 12556 15679 12596 15688
rect 12651 15679 12693 15688
rect 12555 15560 12597 15569
rect 12555 15520 12556 15560
rect 12596 15520 12597 15560
rect 12555 15511 12597 15520
rect 12747 15560 12789 15569
rect 12747 15520 12748 15560
rect 12788 15520 12789 15560
rect 12747 15511 12789 15520
rect 12556 15401 12596 15511
rect 12748 15426 12788 15511
rect 12555 15392 12597 15401
rect 12555 15352 12556 15392
rect 12596 15352 12597 15392
rect 12555 15343 12597 15352
rect 12212 14932 12404 14972
rect 12459 14972 12501 14981
rect 12459 14932 12460 14972
rect 12500 14932 12501 14972
rect 12172 14923 12212 14932
rect 12459 14923 12501 14932
rect 12459 14720 12501 14729
rect 12020 14680 12116 14720
rect 11980 14671 12020 14680
rect 11979 13544 12021 13553
rect 11979 13504 11980 13544
rect 12020 13504 12021 13544
rect 11979 13495 12021 13504
rect 11883 11864 11925 11873
rect 11883 11824 11884 11864
rect 11924 11824 11925 11864
rect 11883 11815 11925 11824
rect 11884 11696 11924 11705
rect 11787 11528 11829 11537
rect 11787 11488 11788 11528
rect 11828 11488 11829 11528
rect 11787 11479 11829 11488
rect 11884 11369 11924 11656
rect 11980 11696 12020 13495
rect 12076 12713 12116 14680
rect 12459 14680 12460 14720
rect 12500 14680 12501 14720
rect 12459 14671 12501 14680
rect 12652 14720 12692 14729
rect 12267 14300 12309 14309
rect 12267 14260 12268 14300
rect 12308 14260 12309 14300
rect 12267 14251 12309 14260
rect 12268 14048 12308 14251
rect 12460 14216 12500 14671
rect 12652 14561 12692 14680
rect 12747 14720 12789 14729
rect 12747 14680 12748 14720
rect 12788 14680 12789 14720
rect 12747 14671 12789 14680
rect 12748 14586 12788 14671
rect 12651 14552 12693 14561
rect 12651 14512 12652 14552
rect 12692 14512 12693 14552
rect 12651 14503 12693 14512
rect 12844 14216 12884 17200
rect 12940 15737 12980 19039
rect 13035 18920 13077 18929
rect 13035 18880 13036 18920
rect 13076 18880 13077 18920
rect 13035 18871 13077 18880
rect 13036 16241 13076 18871
rect 13132 18579 13172 19048
rect 13227 19048 13228 19088
rect 13268 19048 13269 19088
rect 13420 19088 13460 19963
rect 13516 19844 13556 19853
rect 13516 19265 13556 19804
rect 13515 19256 13557 19265
rect 13515 19216 13516 19256
rect 13556 19216 13557 19256
rect 13515 19207 13557 19216
rect 13516 19088 13556 19097
rect 13420 19048 13516 19088
rect 13227 19039 13269 19048
rect 13516 19039 13556 19048
rect 13132 18530 13172 18539
rect 13228 17660 13268 19039
rect 13323 18752 13365 18761
rect 13323 18712 13324 18752
rect 13364 18712 13365 18752
rect 13323 18703 13365 18712
rect 13324 18618 13364 18703
rect 13515 18668 13557 18677
rect 13515 18628 13516 18668
rect 13556 18628 13557 18668
rect 13515 18619 13557 18628
rect 13516 18584 13556 18619
rect 13516 18533 13556 18544
rect 13228 17620 13364 17660
rect 13131 17156 13173 17165
rect 13131 17116 13132 17156
rect 13172 17116 13173 17156
rect 13131 17107 13173 17116
rect 13035 16232 13077 16241
rect 13035 16192 13036 16232
rect 13076 16192 13077 16232
rect 13035 16183 13077 16192
rect 13132 16232 13172 17107
rect 13228 17058 13268 17067
rect 13228 16484 13268 17018
rect 13324 16652 13364 17620
rect 13420 17240 13460 17249
rect 13460 17200 13556 17240
rect 13420 17191 13460 17200
rect 13324 16612 13460 16652
rect 13324 16484 13364 16493
rect 13228 16444 13324 16484
rect 13324 16435 13364 16444
rect 13132 16183 13172 16192
rect 12939 15728 12981 15737
rect 12939 15688 12940 15728
rect 12980 15688 12981 15728
rect 12939 15679 12981 15688
rect 13036 15569 13076 16183
rect 13035 15560 13077 15569
rect 13035 15520 13036 15560
rect 13076 15520 13077 15560
rect 13035 15511 13077 15520
rect 13420 15401 13460 16612
rect 13419 15392 13461 15401
rect 13419 15352 13420 15392
rect 13460 15352 13461 15392
rect 13419 15343 13461 15352
rect 13035 15140 13077 15149
rect 13035 15100 13036 15140
rect 13076 15100 13077 15140
rect 13035 15091 13077 15100
rect 12940 14897 12980 14982
rect 12939 14888 12981 14897
rect 12939 14848 12940 14888
rect 12980 14848 12981 14888
rect 12939 14839 12981 14848
rect 12940 14720 12980 14729
rect 12940 14225 12980 14680
rect 13036 14477 13076 15091
rect 13227 14720 13269 14729
rect 13227 14680 13228 14720
rect 13268 14680 13269 14720
rect 13227 14671 13269 14680
rect 13324 14720 13364 14729
rect 13035 14468 13077 14477
rect 13035 14428 13036 14468
rect 13076 14428 13077 14468
rect 13035 14419 13077 14428
rect 12500 14176 12692 14216
rect 12460 14167 12500 14176
rect 12171 13880 12213 13889
rect 12268 13880 12308 14008
rect 12171 13840 12172 13880
rect 12212 13840 12308 13880
rect 12363 13880 12405 13889
rect 12363 13840 12364 13880
rect 12404 13840 12405 13880
rect 12171 13831 12213 13840
rect 12363 13831 12405 13840
rect 12172 13217 12212 13226
rect 12172 13040 12212 13177
rect 12364 13124 12404 13831
rect 12459 13460 12501 13469
rect 12459 13420 12460 13460
rect 12500 13420 12501 13460
rect 12459 13411 12501 13420
rect 12364 13075 12404 13084
rect 12172 13000 12308 13040
rect 12171 12872 12213 12881
rect 12171 12832 12172 12872
rect 12212 12832 12213 12872
rect 12171 12823 12213 12832
rect 12075 12704 12117 12713
rect 12075 12664 12076 12704
rect 12116 12664 12117 12704
rect 12075 12655 12117 12664
rect 11980 11444 12020 11656
rect 12076 12536 12116 12655
rect 12076 11621 12116 12496
rect 12075 11612 12117 11621
rect 12075 11572 12076 11612
rect 12116 11572 12117 11612
rect 12075 11563 12117 11572
rect 11980 11404 12116 11444
rect 11883 11360 11925 11369
rect 11883 11320 11884 11360
rect 11924 11320 12020 11360
rect 11883 11311 11925 11320
rect 11883 11192 11925 11201
rect 11883 11152 11884 11192
rect 11924 11152 11925 11192
rect 11883 11143 11925 11152
rect 11980 11192 12020 11320
rect 11980 11143 12020 11152
rect 11787 11108 11829 11117
rect 11787 11068 11788 11108
rect 11828 11068 11829 11108
rect 11787 11059 11829 11068
rect 11788 11024 11828 11059
rect 11788 10973 11828 10984
rect 11787 8756 11829 8765
rect 11787 8716 11788 8756
rect 11828 8716 11829 8756
rect 11787 8707 11829 8716
rect 11788 8588 11828 8707
rect 11788 8539 11828 8548
rect 11211 8000 11253 8009
rect 11308 8000 11348 8009
rect 11211 7960 11212 8000
rect 11252 7960 11308 8000
rect 11211 7951 11253 7960
rect 11308 7757 11348 7960
rect 11691 8000 11733 8009
rect 11691 7960 11692 8000
rect 11732 7960 11733 8000
rect 11691 7951 11733 7960
rect 11692 7866 11732 7951
rect 11403 7832 11445 7841
rect 11403 7792 11404 7832
rect 11444 7792 11445 7832
rect 11403 7783 11445 7792
rect 11307 7748 11349 7757
rect 11307 7708 11308 7748
rect 11348 7708 11349 7748
rect 11307 7699 11349 7708
rect 11307 7580 11349 7589
rect 11307 7540 11308 7580
rect 11348 7540 11349 7580
rect 11307 7531 11349 7540
rect 11211 7412 11253 7421
rect 11211 7372 11212 7412
rect 11252 7372 11253 7412
rect 11211 7363 11253 7372
rect 11212 7160 11252 7363
rect 11212 7111 11252 7120
rect 11115 6572 11157 6581
rect 11115 6532 11116 6572
rect 11156 6532 11157 6572
rect 11115 6523 11157 6532
rect 10924 5104 11060 5144
rect 10635 4220 10677 4229
rect 10635 4180 10636 4220
rect 10676 4180 10677 4220
rect 10635 4171 10677 4180
rect 10636 3893 10676 4171
rect 10635 3884 10677 3893
rect 10635 3844 10636 3884
rect 10676 3844 10677 3884
rect 10635 3835 10677 3844
rect 10924 3557 10964 5104
rect 11020 4976 11060 4985
rect 11020 4901 11060 4936
rect 11019 4892 11061 4901
rect 11019 4852 11020 4892
rect 11060 4852 11061 4892
rect 11019 4843 11061 4852
rect 11020 3809 11060 4843
rect 11019 3800 11061 3809
rect 11019 3760 11020 3800
rect 11060 3760 11061 3800
rect 11019 3751 11061 3760
rect 11116 3557 11156 6523
rect 11212 6488 11252 6497
rect 11308 6488 11348 7531
rect 11404 7421 11444 7783
rect 11403 7412 11445 7421
rect 11403 7372 11404 7412
rect 11444 7372 11445 7412
rect 11403 7363 11445 7372
rect 11692 7160 11732 7169
rect 11404 7076 11444 7085
rect 11692 7076 11732 7120
rect 11444 7036 11732 7076
rect 11788 7160 11828 7169
rect 11404 7027 11444 7036
rect 11788 6665 11828 7120
rect 11403 6656 11445 6665
rect 11403 6616 11404 6656
rect 11444 6616 11445 6656
rect 11403 6607 11445 6616
rect 11787 6656 11829 6665
rect 11787 6616 11788 6656
rect 11828 6616 11829 6656
rect 11787 6607 11829 6616
rect 11252 6448 11348 6488
rect 11212 6439 11252 6448
rect 11404 5648 11444 6607
rect 11404 5599 11444 5608
rect 11403 4976 11445 4985
rect 11403 4936 11404 4976
rect 11444 4936 11445 4976
rect 11403 4927 11445 4936
rect 11404 4842 11444 4927
rect 11212 4724 11252 4733
rect 11252 4684 11444 4724
rect 11212 4675 11252 4684
rect 11404 4136 11444 4684
rect 11404 4087 11444 4096
rect 11500 4136 11540 4145
rect 11788 4136 11828 6607
rect 11884 4220 11924 11143
rect 12076 7412 12116 11404
rect 12172 11117 12212 12823
rect 12268 12704 12308 13000
rect 12268 12655 12308 12664
rect 12267 12536 12309 12545
rect 12267 12496 12268 12536
rect 12308 12496 12309 12536
rect 12267 12487 12309 12496
rect 12171 11108 12213 11117
rect 12171 11068 12172 11108
rect 12212 11068 12213 11108
rect 12171 11059 12213 11068
rect 11980 7372 12116 7412
rect 11980 4733 12020 7372
rect 12268 7328 12308 12487
rect 12460 12452 12500 13411
rect 12652 13208 12692 14176
rect 12748 14176 12884 14216
rect 12939 14216 12981 14225
rect 12939 14176 12940 14216
rect 12980 14176 12981 14216
rect 12748 13628 12788 14176
rect 12939 14167 12981 14176
rect 13228 14057 13268 14671
rect 12844 14048 12884 14057
rect 12844 13805 12884 14008
rect 13227 14048 13269 14057
rect 13227 14008 13228 14048
rect 13268 14008 13269 14048
rect 13227 13999 13269 14008
rect 12843 13796 12885 13805
rect 12843 13756 12844 13796
rect 12884 13756 12885 13796
rect 12843 13747 12885 13756
rect 12748 13588 12884 13628
rect 12747 13460 12789 13469
rect 12747 13420 12748 13460
rect 12788 13420 12789 13460
rect 12747 13411 12789 13420
rect 12652 13159 12692 13168
rect 12748 13208 12788 13411
rect 12748 13159 12788 13168
rect 12555 13124 12597 13133
rect 12555 13084 12556 13124
rect 12596 13084 12597 13124
rect 12555 13075 12597 13084
rect 12364 12412 12500 12452
rect 12364 11780 12404 12412
rect 12556 12041 12596 13075
rect 12844 12629 12884 13588
rect 13132 13208 13172 13219
rect 13132 13133 13172 13168
rect 13228 13208 13268 13217
rect 13131 13124 13173 13133
rect 13131 13084 13132 13124
rect 13172 13084 13173 13124
rect 13131 13075 13173 13084
rect 12843 12620 12885 12629
rect 12843 12580 12844 12620
rect 12884 12580 12885 12620
rect 12843 12571 12885 12580
rect 13131 12620 13173 12629
rect 13131 12580 13132 12620
rect 13172 12580 13173 12620
rect 13131 12571 13173 12580
rect 12940 12536 12980 12545
rect 12940 12452 12980 12496
rect 13035 12536 13077 12545
rect 13035 12496 13036 12536
rect 13076 12496 13077 12536
rect 13035 12487 13077 12496
rect 13132 12536 13172 12571
rect 12748 12412 12980 12452
rect 12555 12032 12597 12041
rect 12555 11992 12556 12032
rect 12596 11992 12597 12032
rect 12555 11983 12597 11992
rect 12364 11360 12404 11740
rect 12460 11780 12500 11789
rect 12556 11780 12596 11983
rect 12748 11789 12788 12412
rect 13036 12402 13076 12487
rect 13132 12485 13172 12496
rect 13228 12284 13268 13168
rect 13324 12545 13364 14680
rect 13419 14720 13461 14729
rect 13419 14680 13420 14720
rect 13460 14680 13461 14720
rect 13419 14671 13461 14680
rect 13420 14586 13460 14671
rect 13516 12704 13556 17200
rect 13612 15149 13652 22912
rect 13708 20861 13748 24172
rect 13900 23801 13940 23886
rect 13804 23792 13844 23801
rect 13804 23288 13844 23752
rect 13899 23792 13941 23801
rect 13899 23752 13900 23792
rect 13940 23752 13941 23792
rect 13899 23743 13941 23752
rect 13804 23239 13844 23248
rect 13900 21617 13940 21702
rect 13899 21608 13941 21617
rect 13899 21568 13900 21608
rect 13940 21568 13941 21608
rect 13899 21559 13941 21568
rect 13899 21356 13941 21365
rect 13899 21316 13900 21356
rect 13940 21316 13941 21356
rect 13899 21307 13941 21316
rect 13707 20852 13749 20861
rect 13707 20812 13708 20852
rect 13748 20812 13749 20852
rect 13707 20803 13749 20812
rect 13900 20180 13940 21307
rect 13708 20140 13940 20180
rect 13708 20096 13748 20140
rect 13708 19013 13748 20056
rect 13899 19256 13941 19265
rect 13899 19216 13900 19256
rect 13940 19216 13941 19256
rect 13899 19207 13941 19216
rect 13803 19172 13845 19181
rect 13803 19132 13804 19172
rect 13844 19132 13845 19172
rect 13803 19123 13845 19132
rect 13804 19038 13844 19123
rect 13900 19122 13940 19207
rect 13707 19004 13749 19013
rect 13707 18964 13708 19004
rect 13748 18964 13749 19004
rect 13707 18955 13749 18964
rect 13899 18836 13941 18845
rect 13899 18796 13900 18836
rect 13940 18796 13941 18836
rect 13899 18787 13941 18796
rect 13900 17912 13940 18787
rect 13996 18341 14036 24592
rect 14380 24548 14420 27784
rect 14571 27656 14613 27665
rect 14571 27616 14572 27656
rect 14612 27616 14613 27656
rect 14571 27607 14613 27616
rect 14764 27656 14804 27665
rect 14476 27404 14516 27413
rect 14476 27245 14516 27364
rect 14475 27236 14517 27245
rect 14475 27196 14476 27236
rect 14516 27196 14517 27236
rect 14475 27187 14517 27196
rect 14475 25304 14517 25313
rect 14475 25264 14476 25304
rect 14516 25264 14517 25304
rect 14475 25255 14517 25264
rect 14092 24508 14420 24548
rect 14092 19247 14132 24508
rect 14476 24464 14516 25255
rect 14284 24424 14516 24464
rect 14284 23792 14324 24424
rect 14379 24296 14421 24305
rect 14379 24256 14380 24296
rect 14420 24256 14421 24296
rect 14379 24247 14421 24256
rect 14380 23876 14420 24247
rect 14380 23827 14420 23836
rect 14284 20945 14324 23752
rect 14572 21860 14612 27607
rect 14764 27245 14804 27616
rect 14860 27656 14900 27665
rect 14763 27236 14805 27245
rect 14763 27196 14764 27236
rect 14804 27196 14805 27236
rect 14763 27187 14805 27196
rect 14860 26984 14900 27616
rect 14956 26993 14996 27784
rect 15148 27572 15188 34159
rect 15436 34049 15476 36343
rect 15532 34721 15572 36595
rect 15724 35384 15764 38536
rect 15819 38408 15861 38417
rect 15819 38368 15820 38408
rect 15860 38368 15861 38408
rect 15819 38359 15861 38368
rect 15820 38240 15860 38359
rect 15820 36644 15860 38200
rect 15916 38240 15956 39031
rect 16012 38912 16052 38923
rect 16012 38837 16052 38872
rect 16011 38828 16053 38837
rect 16011 38788 16012 38828
rect 16052 38788 16053 38828
rect 16011 38779 16053 38788
rect 15916 36653 15956 38200
rect 15820 35552 15860 36604
rect 15915 36644 15957 36653
rect 15915 36604 15916 36644
rect 15956 36604 15957 36644
rect 15915 36595 15957 36604
rect 15916 36510 15956 36595
rect 16011 36560 16053 36569
rect 16011 36520 16012 36560
rect 16052 36520 16053 36560
rect 16011 36511 16053 36520
rect 15820 35512 15956 35552
rect 15916 35393 15956 35512
rect 15915 35384 15957 35393
rect 15724 35344 15860 35384
rect 15627 35216 15669 35225
rect 15627 35176 15628 35216
rect 15668 35176 15669 35216
rect 15627 35167 15669 35176
rect 15724 35216 15764 35225
rect 15531 34712 15573 34721
rect 15531 34672 15532 34712
rect 15572 34672 15573 34712
rect 15531 34663 15573 34672
rect 15243 34040 15285 34049
rect 15243 34000 15244 34040
rect 15284 34000 15285 34040
rect 15243 33991 15285 34000
rect 15435 34040 15477 34049
rect 15435 34000 15436 34040
rect 15476 34000 15477 34040
rect 15435 33991 15477 34000
rect 15244 32192 15284 33991
rect 15532 33620 15572 33629
rect 15532 33545 15572 33580
rect 15339 33536 15381 33545
rect 15339 33496 15340 33536
rect 15380 33496 15381 33536
rect 15339 33487 15381 33496
rect 15531 33536 15573 33545
rect 15531 33496 15532 33536
rect 15572 33496 15573 33536
rect 15531 33487 15573 33496
rect 15340 33402 15380 33487
rect 15532 33485 15572 33487
rect 15435 33368 15477 33377
rect 15435 33328 15436 33368
rect 15476 33328 15477 33368
rect 15435 33319 15477 33328
rect 15436 32864 15476 33319
rect 15339 32528 15381 32537
rect 15339 32488 15340 32528
rect 15380 32488 15381 32528
rect 15339 32479 15381 32488
rect 15244 32143 15284 32152
rect 15340 32192 15380 32479
rect 15340 32143 15380 32152
rect 15339 30764 15381 30773
rect 15339 30724 15340 30764
rect 15380 30724 15381 30764
rect 15339 30715 15381 30724
rect 15340 30680 15380 30715
rect 15340 30629 15380 30640
rect 15436 30512 15476 32824
rect 15340 30472 15476 30512
rect 15628 30512 15668 35167
rect 15724 34805 15764 35176
rect 15820 34880 15860 35344
rect 15915 35344 15916 35384
rect 15956 35344 15957 35384
rect 15915 35335 15957 35344
rect 15915 35132 15957 35141
rect 15915 35092 15916 35132
rect 15956 35092 15957 35132
rect 15915 35083 15957 35092
rect 15916 34998 15956 35083
rect 15820 34840 15956 34880
rect 15723 34796 15765 34805
rect 15723 34756 15724 34796
rect 15764 34756 15765 34796
rect 15723 34747 15765 34756
rect 15819 34712 15861 34721
rect 15819 34672 15820 34712
rect 15860 34672 15861 34712
rect 15819 34663 15861 34672
rect 15723 34376 15765 34385
rect 15723 34336 15724 34376
rect 15764 34336 15765 34376
rect 15723 34327 15765 34336
rect 15724 33872 15764 34327
rect 15724 33823 15764 33832
rect 15723 33284 15765 33293
rect 15723 33244 15724 33284
rect 15764 33244 15765 33284
rect 15723 33235 15765 33244
rect 15724 31940 15764 33235
rect 15820 32789 15860 34663
rect 15819 32780 15861 32789
rect 15819 32740 15820 32780
rect 15860 32740 15861 32780
rect 15819 32731 15861 32740
rect 15819 32192 15861 32201
rect 15819 32152 15820 32192
rect 15860 32152 15861 32192
rect 15819 32143 15861 32152
rect 15820 32058 15860 32143
rect 15724 31900 15860 31940
rect 15724 30689 15764 30774
rect 15723 30680 15765 30689
rect 15723 30640 15724 30680
rect 15764 30640 15765 30680
rect 15723 30631 15765 30640
rect 15628 30472 15764 30512
rect 15243 29672 15285 29681
rect 15243 29632 15244 29672
rect 15284 29632 15285 29672
rect 15243 29623 15285 29632
rect 15244 29168 15284 29623
rect 15244 29119 15284 29128
rect 15243 28496 15285 28505
rect 15243 28456 15244 28496
rect 15284 28456 15285 28496
rect 15243 28447 15285 28456
rect 15244 28328 15284 28447
rect 15244 28279 15284 28288
rect 15340 28253 15380 30472
rect 15532 30428 15572 30437
rect 15532 29924 15572 30388
rect 15627 30176 15669 30185
rect 15627 30136 15628 30176
rect 15668 30136 15669 30176
rect 15627 30127 15669 30136
rect 15484 29884 15572 29924
rect 15484 29882 15524 29884
rect 15484 29833 15524 29842
rect 15628 29756 15668 30127
rect 15628 29707 15668 29716
rect 15435 29336 15477 29345
rect 15435 29296 15436 29336
rect 15476 29296 15477 29336
rect 15435 29287 15477 29296
rect 15339 28244 15381 28253
rect 15339 28204 15340 28244
rect 15380 28204 15381 28244
rect 15339 28195 15381 28204
rect 15340 27656 15380 27665
rect 15436 27656 15476 29287
rect 15531 28496 15573 28505
rect 15531 28456 15532 28496
rect 15572 28456 15573 28496
rect 15531 28447 15573 28456
rect 15380 27616 15476 27656
rect 15244 27572 15284 27581
rect 15148 27532 15244 27572
rect 14764 26944 14900 26984
rect 14955 26984 14997 26993
rect 14955 26944 14956 26984
rect 14996 26944 14997 26984
rect 14667 26480 14709 26489
rect 14667 26440 14668 26480
rect 14708 26440 14709 26480
rect 14667 26431 14709 26440
rect 14668 22373 14708 26431
rect 14764 25481 14804 26944
rect 14955 26935 14997 26944
rect 14860 26816 14900 26825
rect 14860 26405 14900 26776
rect 14955 26816 14997 26825
rect 14955 26776 14956 26816
rect 14996 26776 14997 26816
rect 14955 26767 14997 26776
rect 14859 26396 14901 26405
rect 14859 26356 14860 26396
rect 14900 26356 14901 26396
rect 14859 26347 14901 26356
rect 14859 26144 14901 26153
rect 14859 26104 14860 26144
rect 14900 26104 14901 26144
rect 14859 26095 14901 26104
rect 14860 25817 14900 26095
rect 14859 25808 14901 25817
rect 14859 25768 14860 25808
rect 14900 25768 14901 25808
rect 14859 25759 14901 25768
rect 14763 25472 14805 25481
rect 14763 25432 14764 25472
rect 14804 25432 14805 25472
rect 14763 25423 14805 25432
rect 14764 25304 14804 25313
rect 14956 25304 14996 26767
rect 15052 26648 15092 26657
rect 15052 25976 15092 26608
rect 15244 26321 15284 27532
rect 15340 27077 15380 27616
rect 15339 27068 15381 27077
rect 15339 27028 15340 27068
rect 15380 27028 15381 27068
rect 15339 27019 15381 27028
rect 15243 26312 15285 26321
rect 15243 26272 15244 26312
rect 15284 26272 15285 26312
rect 15243 26263 15285 26272
rect 15052 25936 15284 25976
rect 15051 25472 15093 25481
rect 15051 25432 15052 25472
rect 15092 25432 15093 25472
rect 15051 25423 15093 25432
rect 14804 25264 14996 25304
rect 14764 25255 14804 25264
rect 14763 24548 14805 24557
rect 14763 24508 14764 24548
rect 14804 24508 14805 24548
rect 14763 24499 14805 24508
rect 14764 23213 14804 24499
rect 14860 23792 14900 23803
rect 14860 23717 14900 23752
rect 14859 23708 14901 23717
rect 14859 23668 14860 23708
rect 14900 23668 14901 23708
rect 14859 23659 14901 23668
rect 14763 23204 14805 23213
rect 14763 23164 14764 23204
rect 14804 23164 14805 23204
rect 14763 23155 14805 23164
rect 14667 22364 14709 22373
rect 14667 22324 14668 22364
rect 14708 22324 14709 22364
rect 14667 22315 14709 22324
rect 14764 22301 14804 22375
rect 14763 22240 14764 22289
rect 14804 22240 14805 22289
rect 14763 22231 14805 22240
rect 14956 22112 14996 22121
rect 14859 21944 14901 21953
rect 14859 21904 14860 21944
rect 14900 21904 14901 21944
rect 14859 21895 14901 21904
rect 14476 21820 14612 21860
rect 14379 21608 14421 21617
rect 14379 21559 14380 21608
rect 14420 21559 14421 21608
rect 14380 21473 14420 21558
rect 14476 21365 14516 21820
rect 14572 21692 14612 21701
rect 14572 21533 14612 21652
rect 14860 21608 14900 21895
rect 14956 21617 14996 22072
rect 14860 21559 14900 21568
rect 14955 21608 14997 21617
rect 14955 21568 14956 21608
rect 14996 21568 14997 21608
rect 14955 21559 14997 21568
rect 14571 21524 14613 21533
rect 14571 21484 14572 21524
rect 14612 21484 14613 21524
rect 14571 21475 14613 21484
rect 14475 21356 14517 21365
rect 14475 21316 14476 21356
rect 14516 21316 14517 21356
rect 14475 21307 14517 21316
rect 14283 20936 14325 20945
rect 14283 20896 14284 20936
rect 14324 20896 14325 20936
rect 14283 20887 14325 20896
rect 14379 20768 14421 20777
rect 14860 20768 14900 20777
rect 14379 20728 14380 20768
rect 14420 20728 14516 20768
rect 14379 20719 14421 20728
rect 14283 20684 14325 20693
rect 14283 20644 14284 20684
rect 14324 20644 14325 20684
rect 14283 20635 14325 20644
rect 14284 19256 14324 20635
rect 14380 20634 14420 20719
rect 14476 19769 14516 20728
rect 14572 20684 14612 20693
rect 14860 20684 14900 20728
rect 14612 20644 14900 20684
rect 14956 20768 14996 20777
rect 15052 20768 15092 25423
rect 15244 25318 15284 25936
rect 15244 25269 15284 25278
rect 15435 25136 15477 25145
rect 15435 25096 15436 25136
rect 15476 25096 15477 25136
rect 15435 25087 15477 25096
rect 15436 25002 15476 25087
rect 15148 24641 15188 24726
rect 15147 24632 15189 24641
rect 15147 24592 15148 24632
rect 15188 24592 15189 24632
rect 15147 24583 15189 24592
rect 15340 24380 15380 24389
rect 15243 24044 15285 24053
rect 15243 24004 15244 24044
rect 15284 24004 15285 24044
rect 15243 23995 15285 24004
rect 15244 22280 15284 23995
rect 15340 23806 15380 24340
rect 15532 23969 15572 28447
rect 15627 26648 15669 26657
rect 15627 26608 15628 26648
rect 15668 26608 15669 26648
rect 15627 26599 15669 26608
rect 15628 24053 15668 26599
rect 15627 24044 15669 24053
rect 15627 24004 15628 24044
rect 15668 24004 15669 24044
rect 15724 24044 15764 30472
rect 15820 29261 15860 31900
rect 15819 29252 15861 29261
rect 15819 29212 15820 29252
rect 15860 29212 15861 29252
rect 15819 29203 15861 29212
rect 15820 27656 15860 27665
rect 15820 24305 15860 27616
rect 15916 24380 15956 34840
rect 16012 34385 16052 36511
rect 16108 35225 16148 41308
rect 16492 41264 16532 41467
rect 16300 41224 16532 41264
rect 16203 41180 16245 41189
rect 16203 41140 16204 41180
rect 16244 41140 16245 41180
rect 16203 41131 16245 41140
rect 16204 41046 16244 41131
rect 16203 40508 16245 40517
rect 16203 40468 16204 40508
rect 16244 40468 16245 40508
rect 16203 40459 16245 40468
rect 16204 40374 16244 40459
rect 16203 38996 16245 39005
rect 16203 38956 16204 38996
rect 16244 38956 16245 38996
rect 16203 38947 16245 38956
rect 16107 35216 16149 35225
rect 16107 35176 16108 35216
rect 16148 35176 16149 35216
rect 16107 35167 16149 35176
rect 16108 35048 16148 35057
rect 16204 35048 16244 38947
rect 16300 37661 16340 41224
rect 16491 41012 16533 41021
rect 16491 40972 16492 41012
rect 16532 40972 16533 41012
rect 16491 40963 16533 40972
rect 16395 40592 16437 40601
rect 16395 40552 16396 40592
rect 16436 40552 16437 40592
rect 16395 40543 16437 40552
rect 16396 40458 16436 40543
rect 16492 39845 16532 40963
rect 16588 40519 16628 41635
rect 16683 41264 16725 41273
rect 16683 41224 16684 41264
rect 16724 41224 16725 41264
rect 16683 41215 16725 41224
rect 16684 41130 16724 41215
rect 16588 40470 16628 40479
rect 16780 40424 16820 42928
rect 16972 41936 17012 42928
rect 16972 41896 17108 41936
rect 16971 41768 17013 41777
rect 16971 41728 16972 41768
rect 17012 41728 17013 41768
rect 16971 41719 17013 41728
rect 16972 40508 17012 41719
rect 16972 40459 17012 40468
rect 17068 40424 17108 41896
rect 17164 40685 17204 42928
rect 17356 42617 17396 42928
rect 17355 42608 17397 42617
rect 17355 42568 17356 42608
rect 17396 42568 17397 42608
rect 17355 42559 17397 42568
rect 17355 42356 17397 42365
rect 17355 42316 17356 42356
rect 17396 42316 17397 42356
rect 17355 42307 17397 42316
rect 17163 40676 17205 40685
rect 17163 40636 17164 40676
rect 17204 40636 17205 40676
rect 17163 40627 17205 40636
rect 17260 40508 17300 40517
rect 16780 40384 16906 40424
rect 17068 40384 17204 40424
rect 16780 40256 16820 40265
rect 16684 40216 16780 40256
rect 16866 40256 16906 40384
rect 17067 40256 17109 40265
rect 16866 40216 16916 40256
rect 16684 39845 16724 40216
rect 16780 40207 16820 40216
rect 16876 40088 16916 40216
rect 17067 40216 17068 40256
rect 17108 40216 17109 40256
rect 17067 40207 17109 40216
rect 16780 40048 16916 40088
rect 16491 39836 16533 39845
rect 16491 39796 16492 39836
rect 16532 39796 16533 39836
rect 16491 39787 16533 39796
rect 16683 39836 16725 39845
rect 16683 39796 16684 39836
rect 16724 39796 16725 39836
rect 16683 39787 16725 39796
rect 16492 39752 16532 39787
rect 16492 39702 16532 39712
rect 16684 39500 16724 39509
rect 16540 38921 16580 38930
rect 16684 38912 16724 39460
rect 16580 38881 16724 38912
rect 16540 38872 16724 38881
rect 16395 38828 16437 38837
rect 16395 38788 16396 38828
rect 16436 38788 16437 38828
rect 16395 38779 16437 38788
rect 16396 38240 16436 38779
rect 16299 37652 16341 37661
rect 16299 37612 16300 37652
rect 16340 37612 16341 37652
rect 16299 37603 16341 37612
rect 16299 37484 16341 37493
rect 16299 37444 16300 37484
rect 16340 37444 16341 37484
rect 16299 37435 16341 37444
rect 16148 35008 16244 35048
rect 16300 35132 16340 37435
rect 16108 34999 16148 35008
rect 16107 34880 16149 34889
rect 16107 34840 16108 34880
rect 16148 34840 16149 34880
rect 16107 34831 16149 34840
rect 16011 34376 16053 34385
rect 16011 34336 16012 34376
rect 16052 34336 16053 34376
rect 16011 34327 16053 34336
rect 16011 34208 16053 34217
rect 16011 34168 16012 34208
rect 16052 34168 16053 34208
rect 16011 34159 16053 34168
rect 16012 33704 16052 34159
rect 16012 33655 16052 33664
rect 16108 33704 16148 34831
rect 16011 32360 16053 32369
rect 16011 32320 16012 32360
rect 16052 32320 16053 32360
rect 16011 32311 16053 32320
rect 16012 27581 16052 32311
rect 16108 31949 16148 33664
rect 16203 33536 16245 33545
rect 16203 33496 16204 33536
rect 16244 33496 16245 33536
rect 16203 33487 16245 33496
rect 16107 31940 16149 31949
rect 16107 31900 16108 31940
rect 16148 31900 16149 31940
rect 16107 31891 16149 31900
rect 16108 31352 16148 31363
rect 16108 31277 16148 31312
rect 16107 31268 16149 31277
rect 16107 31228 16108 31268
rect 16148 31228 16149 31268
rect 16107 31219 16149 31228
rect 16108 30941 16148 31219
rect 16107 30932 16149 30941
rect 16107 30892 16108 30932
rect 16148 30892 16149 30932
rect 16107 30883 16149 30892
rect 16107 29924 16149 29933
rect 16107 29884 16108 29924
rect 16148 29884 16149 29924
rect 16107 29875 16149 29884
rect 16108 29790 16148 29875
rect 16011 27572 16053 27581
rect 16011 27532 16012 27572
rect 16052 27532 16053 27572
rect 16011 27523 16053 27532
rect 16012 25136 16052 27523
rect 16107 27404 16149 27413
rect 16107 27364 16108 27404
rect 16148 27364 16149 27404
rect 16107 27355 16149 27364
rect 16108 26144 16148 27355
rect 16108 25649 16148 26104
rect 16107 25640 16149 25649
rect 16107 25600 16108 25640
rect 16148 25600 16149 25640
rect 16107 25591 16149 25600
rect 16012 25096 16148 25136
rect 15916 24340 16052 24380
rect 15819 24296 15861 24305
rect 15819 24256 15820 24296
rect 15860 24256 15861 24296
rect 15819 24247 15861 24256
rect 15724 24004 15956 24044
rect 15627 23995 15669 24004
rect 15531 23960 15573 23969
rect 15531 23920 15532 23960
rect 15572 23920 15573 23960
rect 15531 23911 15573 23920
rect 15916 23960 15956 24004
rect 15916 23911 15956 23920
rect 15724 23876 15764 23885
rect 15340 23757 15380 23766
rect 15628 23836 15724 23876
rect 15532 23624 15572 23633
rect 15532 23045 15572 23584
rect 15531 23036 15573 23045
rect 15531 22996 15532 23036
rect 15572 22996 15573 23036
rect 15531 22987 15573 22996
rect 15531 22868 15573 22877
rect 15531 22828 15532 22868
rect 15572 22828 15573 22868
rect 15531 22819 15573 22828
rect 15244 22231 15284 22240
rect 15339 21272 15381 21281
rect 15339 21232 15340 21272
rect 15380 21232 15381 21272
rect 15339 21223 15381 21232
rect 15340 20852 15380 21223
rect 15340 20803 15380 20812
rect 14996 20728 15092 20768
rect 15436 20768 15476 20777
rect 14572 20635 14612 20644
rect 14956 20600 14996 20728
rect 14860 20560 14996 20600
rect 14475 19760 14517 19769
rect 14475 19720 14476 19760
rect 14516 19720 14517 19760
rect 14475 19711 14517 19720
rect 14092 19207 14228 19247
rect 14091 19088 14133 19097
rect 14091 19048 14092 19088
rect 14132 19048 14133 19088
rect 14091 19039 14133 19048
rect 14092 18954 14132 19039
rect 14188 18836 14228 19207
rect 14092 18796 14228 18836
rect 13995 18332 14037 18341
rect 13995 18292 13996 18332
rect 14036 18292 14037 18332
rect 13995 18283 14037 18292
rect 13900 17872 14036 17912
rect 13708 17744 13748 17753
rect 13708 17156 13748 17704
rect 13803 17744 13845 17753
rect 13803 17704 13804 17744
rect 13844 17704 13845 17744
rect 13803 17695 13845 17704
rect 13804 17610 13844 17695
rect 13996 17660 14036 17872
rect 13996 17611 14036 17620
rect 13708 17081 13748 17116
rect 13899 17156 13941 17165
rect 13899 17116 13900 17156
rect 13940 17116 13941 17156
rect 13899 17107 13941 17116
rect 13707 17072 13749 17081
rect 13707 17032 13708 17072
rect 13748 17032 13749 17072
rect 13707 17023 13749 17032
rect 13900 17072 13940 17107
rect 13900 17021 13940 17032
rect 13707 16820 13749 16829
rect 13707 16780 13708 16820
rect 13748 16780 13749 16820
rect 13707 16771 13749 16780
rect 13611 15140 13653 15149
rect 13611 15100 13612 15140
rect 13652 15100 13653 15140
rect 13611 15091 13653 15100
rect 13611 14720 13653 14729
rect 13611 14680 13612 14720
rect 13652 14680 13653 14720
rect 13611 14671 13653 14680
rect 13612 14552 13652 14671
rect 13612 14503 13652 14512
rect 13708 13376 13748 16771
rect 13995 15560 14037 15569
rect 13995 15520 13996 15560
rect 14036 15520 14037 15560
rect 13995 15511 14037 15520
rect 13996 15149 14036 15511
rect 13995 15140 14037 15149
rect 13995 15100 13996 15140
rect 14036 15100 14037 15140
rect 13995 15091 14037 15100
rect 13803 14972 13845 14981
rect 13803 14932 13804 14972
rect 13844 14932 13845 14972
rect 13803 14923 13845 14932
rect 13804 14838 13844 14923
rect 14092 14804 14132 18796
rect 14188 17753 14228 17762
rect 14188 17081 14228 17713
rect 14187 17072 14229 17081
rect 14187 17032 14188 17072
rect 14228 17032 14229 17072
rect 14187 17023 14229 17032
rect 14284 16661 14324 19216
rect 14379 19256 14421 19265
rect 14379 19216 14380 19256
rect 14420 19216 14421 19256
rect 14379 19207 14421 19216
rect 14380 19122 14420 19207
rect 14379 18332 14421 18341
rect 14379 18292 14380 18332
rect 14420 18292 14421 18332
rect 14379 18283 14421 18292
rect 14283 16652 14325 16661
rect 14283 16612 14284 16652
rect 14324 16612 14325 16652
rect 14283 16603 14325 16612
rect 14380 16484 14420 18283
rect 14284 16444 14420 16484
rect 14284 15653 14324 16444
rect 14476 15812 14516 19711
rect 14668 19256 14708 19267
rect 14668 19181 14708 19216
rect 14764 19256 14804 19265
rect 14667 19172 14709 19181
rect 14667 19132 14668 19172
rect 14708 19132 14709 19172
rect 14667 19123 14709 19132
rect 14572 19030 14612 19039
rect 14572 18845 14612 18990
rect 14667 19004 14709 19013
rect 14667 18964 14668 19004
rect 14708 18964 14709 19004
rect 14667 18955 14709 18964
rect 14571 18836 14613 18845
rect 14571 18796 14572 18836
rect 14612 18796 14613 18836
rect 14571 18787 14613 18796
rect 14668 18584 14708 18955
rect 14764 18761 14804 19216
rect 14763 18752 14805 18761
rect 14763 18712 14764 18752
rect 14804 18712 14805 18752
rect 14763 18703 14805 18712
rect 14764 18584 14804 18593
rect 14668 18544 14764 18584
rect 14571 17996 14613 18005
rect 14571 17956 14572 17996
rect 14612 17956 14613 17996
rect 14571 17947 14613 17956
rect 14380 15772 14516 15812
rect 14283 15644 14325 15653
rect 14283 15604 14284 15644
rect 14324 15604 14325 15644
rect 14283 15595 14325 15604
rect 14188 15308 14228 15317
rect 14228 15268 14324 15308
rect 14188 15259 14228 15268
rect 13996 14764 14132 14804
rect 14284 14804 14324 15268
rect 14380 14981 14420 15772
rect 14475 15644 14517 15653
rect 14475 15604 14476 15644
rect 14516 15604 14517 15644
rect 14475 15595 14517 15604
rect 14476 15560 14516 15595
rect 14476 15509 14516 15520
rect 14379 14972 14421 14981
rect 14379 14932 14380 14972
rect 14420 14932 14421 14972
rect 14379 14923 14421 14932
rect 14284 14764 14516 14804
rect 13803 14636 13845 14645
rect 13803 14596 13804 14636
rect 13844 14596 13845 14636
rect 13803 14587 13845 14596
rect 13420 12664 13556 12704
rect 13612 13336 13748 13376
rect 13323 12536 13365 12545
rect 13323 12496 13324 12536
rect 13364 12496 13365 12536
rect 13323 12487 13365 12496
rect 13420 12461 13460 12664
rect 13515 12536 13557 12545
rect 13515 12496 13516 12536
rect 13556 12496 13557 12536
rect 13515 12487 13557 12496
rect 13419 12452 13461 12461
rect 13419 12412 13420 12452
rect 13460 12412 13461 12452
rect 13419 12403 13461 12412
rect 12940 12244 13268 12284
rect 13324 12284 13364 12293
rect 12500 11740 12596 11780
rect 12747 11780 12789 11789
rect 12747 11740 12748 11780
rect 12788 11740 12789 11780
rect 12460 11731 12500 11740
rect 12747 11731 12789 11740
rect 12748 11453 12788 11731
rect 12940 11696 12980 12244
rect 13035 12032 13077 12041
rect 13035 11992 13036 12032
rect 13076 11992 13077 12032
rect 13035 11983 13077 11992
rect 13227 12032 13269 12041
rect 13227 11992 13228 12032
rect 13268 11992 13269 12032
rect 13227 11983 13269 11992
rect 12843 11528 12885 11537
rect 12843 11488 12844 11528
rect 12884 11488 12885 11528
rect 12843 11479 12885 11488
rect 12747 11444 12789 11453
rect 12747 11404 12748 11444
rect 12788 11404 12789 11444
rect 12747 11395 12789 11404
rect 12364 11320 12596 11360
rect 12363 11192 12405 11201
rect 12363 11152 12364 11192
rect 12404 11152 12405 11192
rect 12363 11143 12405 11152
rect 12364 9512 12404 11143
rect 12556 10940 12596 11320
rect 12748 11201 12788 11203
rect 12747 11192 12789 11201
rect 12747 11152 12748 11192
rect 12788 11152 12789 11192
rect 12747 11143 12789 11152
rect 12748 11108 12788 11143
rect 12748 11059 12788 11068
rect 12844 11024 12884 11479
rect 12844 10975 12884 10984
rect 12556 10900 12692 10940
rect 12459 10856 12501 10865
rect 12459 10816 12460 10856
rect 12500 10816 12501 10856
rect 12459 10807 12501 10816
rect 12460 10722 12500 10807
rect 12652 10772 12692 10900
rect 12843 10856 12885 10865
rect 12843 10816 12844 10856
rect 12884 10816 12885 10856
rect 12843 10807 12885 10816
rect 12652 10732 12788 10772
rect 12748 10268 12788 10732
rect 12844 10436 12884 10807
rect 12940 10613 12980 11656
rect 12939 10604 12981 10613
rect 12939 10564 12940 10604
rect 12980 10564 12981 10604
rect 12939 10555 12981 10564
rect 12844 10387 12884 10396
rect 12748 10228 12884 10268
rect 12652 10184 12692 10195
rect 12652 10109 12692 10144
rect 12651 10100 12693 10109
rect 12651 10060 12652 10100
rect 12692 10060 12693 10100
rect 12651 10051 12693 10060
rect 12555 9680 12597 9689
rect 12555 9640 12556 9680
rect 12596 9640 12597 9680
rect 12555 9631 12597 9640
rect 12460 9512 12500 9521
rect 12364 9472 12460 9512
rect 12460 9185 12500 9472
rect 12459 9176 12501 9185
rect 12459 9136 12460 9176
rect 12500 9136 12501 9176
rect 12459 9127 12501 9136
rect 12460 7841 12500 9127
rect 12459 7832 12501 7841
rect 12459 7792 12460 7832
rect 12500 7792 12501 7832
rect 12459 7783 12501 7792
rect 12556 7505 12596 9631
rect 12651 9596 12693 9605
rect 12651 9556 12652 9596
rect 12692 9556 12693 9596
rect 12651 9547 12693 9556
rect 12652 9462 12692 9547
rect 12747 9428 12789 9437
rect 12747 9388 12748 9428
rect 12788 9388 12789 9428
rect 12747 9379 12789 9388
rect 12555 7496 12597 7505
rect 12555 7456 12556 7496
rect 12596 7456 12597 7496
rect 12555 7447 12597 7456
rect 12076 7288 12308 7328
rect 11979 4724 12021 4733
rect 11979 4684 11980 4724
rect 12020 4684 12021 4724
rect 11979 4675 12021 4684
rect 11884 4171 11924 4180
rect 11540 4096 11828 4136
rect 11979 4136 12021 4145
rect 11979 4096 11980 4136
rect 12020 4096 12021 4136
rect 11500 4087 11540 4096
rect 11979 4087 12021 4096
rect 11980 4002 12020 4087
rect 10923 3548 10965 3557
rect 10923 3508 10924 3548
rect 10964 3508 10965 3548
rect 10923 3499 10965 3508
rect 11115 3548 11157 3557
rect 11115 3508 11116 3548
rect 11156 3508 11252 3548
rect 11115 3499 11157 3508
rect 11212 3464 11252 3508
rect 11212 3415 11252 3424
rect 11403 3464 11445 3473
rect 11403 3424 11404 3464
rect 11444 3424 11445 3464
rect 11403 3415 11445 3424
rect 10636 3212 10676 3221
rect 10676 3172 10964 3212
rect 10636 3163 10676 3172
rect 10388 2584 10580 2624
rect 10636 2792 10676 2801
rect 10348 2575 10388 2584
rect 10155 2288 10197 2297
rect 10155 2248 10156 2288
rect 10196 2248 10197 2288
rect 10155 2239 10197 2248
rect 10060 1903 10100 1912
rect 9772 1818 9812 1903
rect 10347 1868 10389 1877
rect 10347 1828 10348 1868
rect 10388 1828 10389 1868
rect 10347 1819 10389 1828
rect 10348 1734 10388 1819
rect 10540 1700 10580 1709
rect 10540 1289 10580 1660
rect 10539 1280 10581 1289
rect 10539 1240 10540 1280
rect 10580 1240 10581 1280
rect 10539 1231 10581 1240
rect 10636 1205 10676 2752
rect 10924 2624 10964 3172
rect 11404 2708 11444 3415
rect 11979 3044 12021 3053
rect 11979 3004 11980 3044
rect 12020 3004 12021 3044
rect 11979 2995 12021 3004
rect 11499 2792 11541 2801
rect 11499 2752 11500 2792
rect 11540 2752 11541 2792
rect 11499 2743 11541 2752
rect 11404 2659 11444 2668
rect 11500 2708 11540 2743
rect 11500 2657 11540 2668
rect 10924 2575 10964 2584
rect 11019 2624 11061 2633
rect 11019 2584 11020 2624
rect 11060 2584 11061 2624
rect 11019 2575 11061 2584
rect 11980 2624 12020 2995
rect 11980 2575 12020 2584
rect 11020 2490 11060 2575
rect 11211 2540 11253 2549
rect 11211 2500 11212 2540
rect 11252 2500 11253 2540
rect 11211 2491 11253 2500
rect 11212 2120 11252 2491
rect 11020 2080 11252 2120
rect 10731 1868 10773 1877
rect 10731 1828 10732 1868
rect 10772 1828 10773 1868
rect 10731 1819 10773 1828
rect 10732 1734 10772 1819
rect 10924 1700 10964 1709
rect 10924 1373 10964 1660
rect 10923 1364 10965 1373
rect 10923 1324 10924 1364
rect 10964 1324 10965 1364
rect 10923 1315 10965 1324
rect 9867 1196 9909 1205
rect 9964 1196 10004 1205
rect 9867 1156 9868 1196
rect 9908 1156 9964 1196
rect 9867 1147 9909 1156
rect 9964 1147 10004 1156
rect 10347 1196 10389 1205
rect 10347 1156 10348 1196
rect 10388 1156 10389 1196
rect 10347 1147 10389 1156
rect 10635 1196 10677 1205
rect 10635 1156 10636 1196
rect 10676 1156 10677 1196
rect 10635 1147 10677 1156
rect 10924 1196 10964 1205
rect 11020 1196 11060 2080
rect 11500 1952 11540 1961
rect 11115 1868 11157 1877
rect 11115 1828 11116 1868
rect 11156 1828 11157 1868
rect 11115 1819 11157 1828
rect 11116 1734 11156 1819
rect 11500 1793 11540 1912
rect 11499 1784 11541 1793
rect 11499 1744 11500 1784
rect 11540 1744 11541 1784
rect 11499 1735 11541 1744
rect 11307 1700 11349 1709
rect 11307 1660 11308 1700
rect 11348 1660 11349 1700
rect 11307 1651 11349 1660
rect 11308 1566 11348 1651
rect 11115 1448 11157 1457
rect 11115 1408 11116 1448
rect 11156 1408 11157 1448
rect 11115 1399 11157 1408
rect 10964 1156 11060 1196
rect 10924 1147 10964 1156
rect 10348 1062 10388 1147
rect 9772 944 9812 953
rect 10156 944 10196 953
rect 9812 904 10100 944
rect 9772 895 9812 904
rect 9867 608 9909 617
rect 9867 568 9868 608
rect 9908 568 9909 608
rect 9867 559 9909 568
rect 9868 80 9908 559
rect 10060 80 10100 904
rect 10156 449 10196 904
rect 10251 944 10293 953
rect 10251 904 10252 944
rect 10292 904 10293 944
rect 10251 895 10293 904
rect 10540 944 10580 953
rect 10155 440 10197 449
rect 10155 400 10156 440
rect 10196 400 10197 440
rect 10155 391 10197 400
rect 10252 80 10292 895
rect 10443 692 10485 701
rect 10443 652 10444 692
rect 10484 652 10485 692
rect 10443 643 10485 652
rect 10444 80 10484 643
rect 10540 533 10580 904
rect 10731 944 10773 953
rect 10731 904 10732 944
rect 10772 904 10773 944
rect 10731 895 10773 904
rect 10732 810 10772 895
rect 10827 860 10869 869
rect 10827 820 10828 860
rect 10868 820 10869 860
rect 11116 860 11156 1399
rect 11691 1280 11733 1289
rect 11691 1240 11692 1280
rect 11732 1240 11733 1280
rect 11691 1231 11733 1240
rect 11212 1196 11252 1205
rect 11212 1037 11252 1156
rect 11211 1028 11253 1037
rect 11211 988 11212 1028
rect 11252 988 11253 1028
rect 11211 979 11253 988
rect 11403 944 11445 953
rect 11403 904 11404 944
rect 11444 904 11445 944
rect 11403 895 11445 904
rect 11596 944 11636 953
rect 11116 820 11252 860
rect 10827 811 10869 820
rect 10539 524 10581 533
rect 10539 484 10540 524
rect 10580 484 10581 524
rect 10539 475 10581 484
rect 10635 104 10677 113
rect 10635 80 10636 104
rect 6260 64 6280 80
rect 6200 0 6280 64
rect 6392 0 6472 80
rect 6584 0 6664 80
rect 6776 0 6856 80
rect 6968 0 7048 80
rect 7160 0 7240 80
rect 7352 0 7432 80
rect 7544 0 7624 80
rect 7736 0 7816 80
rect 7928 0 8008 80
rect 8120 0 8200 80
rect 8312 0 8392 80
rect 8504 0 8584 80
rect 8696 0 8776 80
rect 8888 0 8968 80
rect 9080 0 9160 80
rect 9272 0 9352 80
rect 9464 0 9544 80
rect 9656 0 9736 80
rect 9848 0 9928 80
rect 10040 0 10120 80
rect 10232 0 10312 80
rect 10424 0 10504 80
rect 10616 64 10636 80
rect 10676 80 10677 104
rect 10828 80 10868 811
rect 11019 356 11061 365
rect 11019 316 11020 356
rect 11060 316 11061 356
rect 11019 307 11061 316
rect 11020 80 11060 307
rect 11212 80 11252 820
rect 11404 810 11444 895
rect 11596 617 11636 904
rect 11692 692 11732 1231
rect 11788 1196 11828 1205
rect 12076 1196 12116 7288
rect 12171 7160 12213 7169
rect 12171 7120 12172 7160
rect 12212 7120 12213 7160
rect 12171 7111 12213 7120
rect 12268 7160 12308 7169
rect 12748 7160 12788 9379
rect 12172 7026 12212 7111
rect 12268 6581 12308 7120
rect 12556 7120 12748 7160
rect 12459 7076 12501 7085
rect 12459 7036 12460 7076
rect 12500 7036 12501 7076
rect 12459 7027 12501 7036
rect 12267 6572 12309 6581
rect 12267 6532 12268 6572
rect 12308 6532 12309 6572
rect 12267 6523 12309 6532
rect 12268 4145 12308 6523
rect 12460 6488 12500 7027
rect 12363 5144 12405 5153
rect 12363 5104 12364 5144
rect 12404 5104 12405 5144
rect 12363 5095 12405 5104
rect 12267 4136 12309 4145
rect 12267 4096 12268 4136
rect 12308 4096 12309 4136
rect 12267 4087 12309 4096
rect 12364 3473 12404 5095
rect 12460 5069 12500 6448
rect 12459 5060 12501 5069
rect 12459 5020 12460 5060
rect 12500 5020 12501 5060
rect 12459 5011 12501 5020
rect 12556 4150 12596 7120
rect 12748 7111 12788 7120
rect 12844 6656 12884 10228
rect 13036 9689 13076 11983
rect 13228 11360 13268 11983
rect 13324 11705 13364 12244
rect 13323 11696 13365 11705
rect 13323 11656 13324 11696
rect 13364 11656 13365 11696
rect 13323 11647 13365 11656
rect 13420 11701 13460 11710
rect 13420 11621 13460 11661
rect 13419 11612 13461 11621
rect 13419 11572 13420 11612
rect 13460 11572 13461 11612
rect 13419 11563 13461 11572
rect 13516 11453 13556 12487
rect 13612 12461 13652 13336
rect 13708 13208 13748 13219
rect 13708 13133 13748 13168
rect 13707 13124 13749 13133
rect 13707 13084 13708 13124
rect 13748 13084 13749 13124
rect 13707 13075 13749 13084
rect 13611 12452 13653 12461
rect 13611 12412 13612 12452
rect 13652 12412 13653 12452
rect 13611 12403 13653 12412
rect 13612 12041 13652 12403
rect 13611 12032 13653 12041
rect 13611 11992 13612 12032
rect 13652 11992 13653 12032
rect 13611 11983 13653 11992
rect 13612 11537 13652 11622
rect 13611 11528 13653 11537
rect 13611 11488 13612 11528
rect 13652 11488 13653 11528
rect 13611 11479 13653 11488
rect 13515 11444 13557 11453
rect 13515 11404 13516 11444
rect 13556 11404 13557 11444
rect 13515 11395 13557 11404
rect 13419 11360 13461 11369
rect 13228 11320 13364 11360
rect 13131 11024 13173 11033
rect 13131 10984 13132 11024
rect 13172 10984 13173 11024
rect 13131 10975 13173 10984
rect 13132 10890 13172 10975
rect 13227 10772 13269 10781
rect 13227 10732 13228 10772
rect 13268 10732 13269 10772
rect 13227 10723 13269 10732
rect 13228 10529 13268 10723
rect 13227 10520 13269 10529
rect 13227 10480 13228 10520
rect 13268 10480 13269 10520
rect 13227 10471 13269 10480
rect 13131 10184 13173 10193
rect 13131 10144 13132 10184
rect 13172 10144 13173 10184
rect 13131 10135 13173 10144
rect 13228 10184 13268 10471
rect 13228 10135 13268 10144
rect 13035 9680 13077 9689
rect 13035 9640 13036 9680
rect 13076 9640 13077 9680
rect 13035 9631 13077 9640
rect 12939 9596 12981 9605
rect 12939 9556 12940 9596
rect 12980 9556 12981 9596
rect 12939 9547 12981 9556
rect 12940 9512 12980 9547
rect 12940 9461 12980 9472
rect 13036 9512 13076 9521
rect 13036 8840 13076 9472
rect 12940 8800 13076 8840
rect 12940 8504 12980 8800
rect 13036 8672 13076 8681
rect 13132 8672 13172 10135
rect 13076 8632 13172 8672
rect 13036 8623 13076 8632
rect 12940 8464 13076 8504
rect 12940 8000 12980 8009
rect 12940 7841 12980 7960
rect 12939 7832 12981 7841
rect 12939 7792 12940 7832
rect 12980 7792 12981 7832
rect 12939 7783 12981 7792
rect 13036 6740 13076 8464
rect 13132 7748 13172 7757
rect 13172 7708 13268 7748
rect 13132 7699 13172 7708
rect 13228 7174 13268 7708
rect 13228 7125 13268 7134
rect 13036 6700 13172 6740
rect 12844 6616 13076 6656
rect 12652 6572 12692 6581
rect 12692 6532 12980 6572
rect 12652 6523 12692 6532
rect 12940 6488 12980 6532
rect 12940 6439 12980 6448
rect 13036 6488 13076 6616
rect 13036 5741 13076 6448
rect 13035 5732 13077 5741
rect 13035 5692 13036 5732
rect 13076 5692 13077 5732
rect 13035 5683 13077 5692
rect 12652 5648 12692 5657
rect 12652 5069 12692 5608
rect 12844 5480 12884 5489
rect 12748 5440 12844 5480
rect 12651 5060 12693 5069
rect 12651 5020 12652 5060
rect 12692 5020 12693 5060
rect 12651 5011 12693 5020
rect 12459 4127 12596 4150
rect 12499 4110 12596 4127
rect 12652 4976 12692 5011
rect 12459 4061 12499 4087
rect 12459 4052 12501 4061
rect 12459 4012 12460 4052
rect 12500 4012 12501 4052
rect 12459 4003 12501 4012
rect 12652 3884 12692 4936
rect 12748 4808 12788 5440
rect 12844 5431 12884 5440
rect 13132 5312 13172 6700
rect 13227 5816 13269 5825
rect 13227 5776 13228 5816
rect 13268 5776 13269 5816
rect 13227 5767 13269 5776
rect 13228 5648 13268 5767
rect 13228 5489 13268 5608
rect 13227 5480 13269 5489
rect 13227 5440 13228 5480
rect 13268 5440 13269 5480
rect 13227 5431 13269 5440
rect 13132 5272 13268 5312
rect 12844 5060 12884 5069
rect 12884 5020 13172 5060
rect 12844 5011 12884 5020
rect 13132 4996 13172 5020
rect 13132 4947 13172 4956
rect 13228 4976 13268 5272
rect 13228 4901 13268 4936
rect 13035 4892 13077 4901
rect 13035 4852 13036 4892
rect 13076 4852 13077 4892
rect 13035 4843 13077 4852
rect 13227 4892 13269 4901
rect 13227 4852 13228 4892
rect 13268 4852 13269 4892
rect 13227 4843 13269 4852
rect 12748 4768 12980 4808
rect 12940 4150 12980 4768
rect 12940 4101 12980 4110
rect 12460 3844 12692 3884
rect 12843 3884 12885 3893
rect 12843 3844 12844 3884
rect 12884 3844 12885 3884
rect 12363 3464 12405 3473
rect 12363 3424 12364 3464
rect 12404 3424 12405 3464
rect 12363 3415 12405 3424
rect 12460 3464 12500 3844
rect 12843 3835 12885 3844
rect 12844 3473 12884 3835
rect 12460 3415 12500 3424
rect 12843 3464 12885 3473
rect 12843 3424 12844 3464
rect 12884 3424 12885 3464
rect 12843 3415 12885 3424
rect 12652 3212 12692 3221
rect 12556 3172 12652 3212
rect 12556 2708 12596 3172
rect 12652 3163 12692 3172
rect 12508 2668 12596 2708
rect 12508 2666 12548 2668
rect 12508 2617 12548 2626
rect 12652 2549 12692 2634
rect 12651 2540 12693 2549
rect 12651 2500 12652 2540
rect 12692 2500 12693 2540
rect 12651 2491 12693 2500
rect 12747 2288 12789 2297
rect 12747 2248 12748 2288
rect 12788 2248 12789 2288
rect 12747 2239 12789 2248
rect 12748 1952 12788 2239
rect 12651 1868 12693 1877
rect 12651 1828 12652 1868
rect 12692 1828 12693 1868
rect 12651 1819 12693 1828
rect 12363 1700 12405 1709
rect 12363 1660 12364 1700
rect 12404 1660 12405 1700
rect 12363 1651 12405 1660
rect 12171 1364 12213 1373
rect 12171 1324 12172 1364
rect 12212 1324 12213 1364
rect 12171 1315 12213 1324
rect 11828 1156 12116 1196
rect 11788 1147 11828 1156
rect 11979 944 12021 953
rect 11979 904 11980 944
rect 12020 904 12021 944
rect 11979 895 12021 904
rect 11692 652 11828 692
rect 11595 608 11637 617
rect 11595 568 11596 608
rect 11636 568 11637 608
rect 11595 559 11637 568
rect 11403 524 11445 533
rect 11403 484 11404 524
rect 11444 484 11445 524
rect 11403 475 11445 484
rect 11404 80 11444 475
rect 11595 440 11637 449
rect 11595 400 11596 440
rect 11636 400 11637 440
rect 11595 391 11637 400
rect 11596 80 11636 391
rect 11788 80 11828 652
rect 11980 80 12020 895
rect 12172 80 12212 1315
rect 12364 80 12404 1651
rect 12555 1280 12597 1289
rect 12555 1240 12556 1280
rect 12596 1240 12597 1280
rect 12555 1231 12597 1240
rect 12556 80 12596 1231
rect 12652 1037 12692 1819
rect 12748 1793 12788 1912
rect 12747 1784 12789 1793
rect 12747 1744 12748 1784
rect 12788 1744 12789 1784
rect 12747 1735 12789 1744
rect 12747 1112 12789 1121
rect 12747 1072 12748 1112
rect 12788 1072 12789 1112
rect 12844 1112 12884 3415
rect 13036 2633 13076 4843
rect 13227 4724 13269 4733
rect 13227 4684 13228 4724
rect 13268 4684 13269 4724
rect 13227 4675 13269 4684
rect 13131 3968 13173 3977
rect 13131 3928 13132 3968
rect 13172 3928 13173 3968
rect 13131 3919 13173 3928
rect 13132 3834 13172 3919
rect 13035 2624 13077 2633
rect 13035 2584 13036 2624
rect 13076 2584 13077 2624
rect 13035 2575 13077 2584
rect 13228 2540 13268 4675
rect 13324 4136 13364 11320
rect 13419 11320 13420 11360
rect 13460 11320 13461 11360
rect 13419 11311 13461 11320
rect 13420 11024 13460 11311
rect 13420 10975 13460 10984
rect 13708 11024 13748 13075
rect 13804 12713 13844 14587
rect 13996 13124 14036 14764
rect 14188 14720 14228 14729
rect 14476 14720 14516 14764
rect 14228 14680 14420 14720
rect 14188 14671 14228 14680
rect 14091 14636 14133 14645
rect 14091 14596 14092 14636
rect 14132 14596 14133 14636
rect 14091 14587 14133 14596
rect 14092 14502 14132 14587
rect 14091 14300 14133 14309
rect 14091 14260 14092 14300
rect 14132 14260 14133 14300
rect 14091 14251 14133 14260
rect 14283 14300 14325 14309
rect 14283 14260 14284 14300
rect 14324 14260 14325 14300
rect 14283 14251 14325 14260
rect 14092 14048 14132 14251
rect 14187 14216 14229 14225
rect 14187 14176 14188 14216
rect 14228 14176 14229 14216
rect 14187 14167 14229 14176
rect 14284 14216 14324 14251
rect 14092 13999 14132 14008
rect 14188 13721 14228 14167
rect 14284 14165 14324 14176
rect 14284 13796 14324 13805
rect 14187 13712 14229 13721
rect 14187 13672 14188 13712
rect 14228 13672 14229 13712
rect 14187 13663 14229 13672
rect 14284 13544 14324 13756
rect 14188 13504 14324 13544
rect 14188 13222 14228 13504
rect 14188 13173 14228 13182
rect 14380 13124 14420 14680
rect 14476 14671 14516 14680
rect 14475 14048 14517 14057
rect 14475 14008 14476 14048
rect 14516 14008 14517 14048
rect 14475 13999 14517 14008
rect 14476 13914 14516 13999
rect 14476 13796 14516 13807
rect 14476 13721 14516 13756
rect 14475 13712 14517 13721
rect 14475 13672 14476 13712
rect 14516 13672 14517 13712
rect 14475 13663 14517 13672
rect 13996 13084 14228 13124
rect 13803 12704 13845 12713
rect 13803 12664 13804 12704
rect 13844 12664 13845 12704
rect 13803 12655 13845 12664
rect 13804 12536 13844 12547
rect 13804 12461 13844 12496
rect 13803 12452 13845 12461
rect 13803 12412 13804 12452
rect 13844 12412 13845 12452
rect 13803 12403 13845 12412
rect 14091 12032 14133 12041
rect 14091 11992 14092 12032
rect 14132 11992 14133 12032
rect 14091 11983 14133 11992
rect 13995 11864 14037 11873
rect 13995 11824 13996 11864
rect 14036 11824 14037 11864
rect 13995 11815 14037 11824
rect 13996 11710 14036 11815
rect 13708 10975 13748 10984
rect 13804 11696 13844 11705
rect 13996 11661 14036 11670
rect 14092 11696 14132 11983
rect 13516 10940 13556 10949
rect 13516 10856 13556 10900
rect 13804 10856 13844 11656
rect 14092 11647 14132 11656
rect 13899 11528 13941 11537
rect 13899 11488 13900 11528
rect 13940 11488 13941 11528
rect 13899 11479 13941 11488
rect 13900 11394 13940 11479
rect 14091 11444 14133 11453
rect 14091 11404 14092 11444
rect 14132 11404 14133 11444
rect 14091 11395 14133 11404
rect 13516 10816 13844 10856
rect 14092 10613 14132 11395
rect 13707 10604 13749 10613
rect 13707 10564 13708 10604
rect 13748 10564 13749 10604
rect 13707 10555 13749 10564
rect 14091 10604 14133 10613
rect 14091 10564 14092 10604
rect 14132 10564 14133 10604
rect 14091 10555 14133 10564
rect 13515 10520 13557 10529
rect 13515 10480 13516 10520
rect 13556 10480 13557 10520
rect 13515 10471 13557 10480
rect 13516 9512 13556 10471
rect 13611 10100 13653 10109
rect 13611 10060 13612 10100
rect 13652 10060 13653 10100
rect 13611 10051 13653 10060
rect 13420 9428 13460 9437
rect 13420 7169 13460 9388
rect 13419 7160 13461 7169
rect 13419 7120 13420 7160
rect 13460 7120 13461 7160
rect 13419 7111 13461 7120
rect 13419 6992 13461 7001
rect 13419 6952 13420 6992
rect 13460 6952 13461 6992
rect 13419 6943 13461 6952
rect 13420 6858 13460 6943
rect 13420 6497 13460 6582
rect 13516 6572 13556 9472
rect 13612 6917 13652 10051
rect 13708 9185 13748 10555
rect 14092 9764 14132 10555
rect 14188 10529 14228 13084
rect 14380 13075 14420 13084
rect 14572 11873 14612 17947
rect 14667 17828 14709 17837
rect 14667 17788 14668 17828
rect 14708 17788 14709 17828
rect 14667 17779 14709 17788
rect 14668 17744 14708 17779
rect 14668 17693 14708 17704
rect 14764 17249 14804 18544
rect 14860 18509 14900 20560
rect 15243 20516 15285 20525
rect 15243 20476 15244 20516
rect 15284 20476 15285 20516
rect 15243 20467 15285 20476
rect 14956 20096 14996 20105
rect 14956 19937 14996 20056
rect 15148 20096 15188 20105
rect 14955 19928 14997 19937
rect 14955 19888 14956 19928
rect 14996 19888 14997 19928
rect 14955 19879 14997 19888
rect 15051 19844 15093 19853
rect 15051 19804 15052 19844
rect 15092 19804 15093 19844
rect 15051 19795 15093 19804
rect 15052 19508 15092 19795
rect 15052 19459 15092 19468
rect 15148 19340 15188 20056
rect 15244 20096 15284 20467
rect 15436 20441 15476 20728
rect 15435 20432 15477 20441
rect 15435 20392 15436 20432
rect 15476 20392 15477 20432
rect 15435 20383 15477 20392
rect 15244 19844 15284 20056
rect 15436 20264 15476 20273
rect 15244 19804 15380 19844
rect 15243 19676 15285 19685
rect 15243 19636 15244 19676
rect 15284 19636 15285 19676
rect 15243 19627 15285 19636
rect 15123 19300 15188 19340
rect 14955 19256 14997 19265
rect 15123 19256 15163 19300
rect 14955 19216 14956 19256
rect 14996 19216 15163 19256
rect 15244 19256 15284 19627
rect 14955 19207 14997 19216
rect 15244 19207 15284 19216
rect 14956 18752 14996 19207
rect 15147 19004 15189 19013
rect 15147 18964 15148 19004
rect 15188 18964 15189 19004
rect 15147 18955 15189 18964
rect 15051 18836 15093 18845
rect 15051 18796 15052 18836
rect 15092 18796 15093 18836
rect 15051 18787 15093 18796
rect 14956 18703 14996 18712
rect 14859 18500 14901 18509
rect 14859 18460 14860 18500
rect 14900 18460 14901 18500
rect 14859 18451 14901 18460
rect 14955 18332 14997 18341
rect 14955 18292 14956 18332
rect 14996 18292 14997 18332
rect 14955 18283 14997 18292
rect 14956 18198 14996 18283
rect 15052 17501 15092 18787
rect 15148 18584 15188 18955
rect 15148 18535 15188 18544
rect 15244 18584 15284 18593
rect 15244 18005 15284 18544
rect 15243 17996 15285 18005
rect 15243 17956 15244 17996
rect 15284 17956 15285 17996
rect 15243 17947 15285 17956
rect 15243 17828 15285 17837
rect 15243 17788 15244 17828
rect 15284 17788 15285 17828
rect 15243 17779 15285 17788
rect 15148 17744 15188 17753
rect 15051 17492 15093 17501
rect 15051 17452 15052 17492
rect 15092 17452 15093 17492
rect 15051 17443 15093 17452
rect 15148 17333 15188 17704
rect 15244 17694 15284 17779
rect 15340 17576 15380 19804
rect 15436 19424 15476 20224
rect 15532 19685 15572 22819
rect 15628 20189 15668 23836
rect 15724 23827 15764 23836
rect 16012 23708 16052 24340
rect 15724 23668 16052 23708
rect 16108 23792 16148 25096
rect 15627 20180 15669 20189
rect 15627 20140 15628 20180
rect 15668 20140 15669 20180
rect 15627 20131 15669 20140
rect 15724 19853 15764 23668
rect 16108 23624 16148 23752
rect 16012 23584 16148 23624
rect 15819 22700 15861 22709
rect 15819 22660 15820 22700
rect 15860 22660 15861 22700
rect 15819 22651 15861 22660
rect 15820 20525 15860 22651
rect 15915 20936 15957 20945
rect 15915 20896 15916 20936
rect 15956 20896 15957 20936
rect 15915 20887 15957 20896
rect 15916 20768 15956 20887
rect 15916 20719 15956 20728
rect 15819 20516 15861 20525
rect 15819 20476 15820 20516
rect 15860 20476 15861 20516
rect 15819 20467 15861 20476
rect 15820 20096 15860 20107
rect 15820 20021 15860 20056
rect 15915 20096 15957 20105
rect 15915 20056 15916 20096
rect 15956 20056 15957 20096
rect 15915 20047 15957 20056
rect 15819 20012 15861 20021
rect 15819 19972 15820 20012
rect 15860 19972 15861 20012
rect 15819 19963 15861 19972
rect 15723 19844 15765 19853
rect 15723 19804 15724 19844
rect 15764 19804 15765 19844
rect 15723 19795 15765 19804
rect 15531 19676 15573 19685
rect 15531 19636 15532 19676
rect 15572 19636 15573 19676
rect 15531 19627 15573 19636
rect 15436 19384 15572 19424
rect 15435 19088 15477 19097
rect 15435 19048 15436 19088
rect 15476 19048 15477 19088
rect 15435 19039 15477 19048
rect 15436 18584 15476 19039
rect 15436 18535 15476 18544
rect 15532 18584 15572 19384
rect 15820 18929 15860 19963
rect 15819 18920 15861 18929
rect 15819 18880 15820 18920
rect 15860 18880 15861 18920
rect 15819 18871 15861 18880
rect 15628 18761 15668 18846
rect 15627 18752 15669 18761
rect 15627 18712 15628 18752
rect 15668 18712 15669 18752
rect 15627 18703 15669 18712
rect 15819 18752 15861 18761
rect 15819 18712 15820 18752
rect 15860 18712 15861 18752
rect 15819 18703 15861 18712
rect 15633 18584 15673 18593
rect 15532 18535 15572 18544
rect 15628 18544 15633 18584
rect 15628 18535 15673 18544
rect 15628 18416 15668 18535
rect 15244 17536 15380 17576
rect 15436 18376 15668 18416
rect 14955 17324 14997 17333
rect 14955 17284 14956 17324
rect 14996 17284 14997 17324
rect 14955 17275 14997 17284
rect 15147 17324 15189 17333
rect 15147 17284 15148 17324
rect 15188 17284 15189 17324
rect 15147 17275 15189 17284
rect 14763 17240 14805 17249
rect 14763 17200 14764 17240
rect 14804 17200 14805 17240
rect 14763 17191 14805 17200
rect 14667 16652 14709 16661
rect 14667 16612 14668 16652
rect 14708 16612 14709 16652
rect 14667 16603 14709 16612
rect 14668 14477 14708 16603
rect 14956 16325 14996 17275
rect 15148 17165 15188 17196
rect 15147 17156 15189 17165
rect 15147 17116 15148 17156
rect 15188 17116 15189 17156
rect 15147 17107 15189 17116
rect 15148 17072 15188 17107
rect 14955 16316 14997 16325
rect 14955 16276 14956 16316
rect 14996 16276 14997 16316
rect 14955 16267 14997 16276
rect 14859 14888 14901 14897
rect 14859 14848 14860 14888
rect 14900 14848 14901 14888
rect 14859 14839 14901 14848
rect 14763 14804 14805 14813
rect 14763 14764 14764 14804
rect 14804 14764 14805 14804
rect 14763 14755 14805 14764
rect 14764 14720 14804 14755
rect 14667 14468 14709 14477
rect 14667 14428 14668 14468
rect 14708 14428 14709 14468
rect 14667 14419 14709 14428
rect 14764 14309 14804 14680
rect 14860 14720 14900 14839
rect 15052 14729 15092 14814
rect 14860 14671 14900 14680
rect 14948 14720 14996 14729
rect 14948 14680 14949 14720
rect 14948 14671 14996 14680
rect 15051 14720 15093 14729
rect 15051 14680 15052 14720
rect 15092 14680 15093 14720
rect 15051 14671 15093 14680
rect 14949 14592 14989 14671
rect 14859 14468 14901 14477
rect 14859 14428 14860 14468
rect 14900 14428 14901 14468
rect 15148 14468 15188 17032
rect 15244 14729 15284 17536
rect 15436 17240 15476 18376
rect 15723 18332 15765 18341
rect 15723 18292 15724 18332
rect 15764 18292 15765 18332
rect 15723 18283 15765 18292
rect 15627 18248 15669 18257
rect 15627 18208 15628 18248
rect 15668 18208 15669 18248
rect 15627 18199 15669 18208
rect 15628 17744 15668 18199
rect 15724 17837 15764 18283
rect 15723 17828 15765 17837
rect 15723 17788 15724 17828
rect 15764 17788 15765 17828
rect 15723 17779 15765 17788
rect 15628 17695 15668 17704
rect 15724 17744 15764 17779
rect 15724 17576 15764 17704
rect 15436 17191 15476 17200
rect 15532 17536 15764 17576
rect 15339 17072 15381 17081
rect 15339 17032 15340 17072
rect 15380 17032 15381 17072
rect 15339 17023 15381 17032
rect 15532 17072 15572 17536
rect 15532 17023 15572 17032
rect 15628 17072 15668 17081
rect 15820 17072 15860 18703
rect 15916 17240 15956 20047
rect 16012 18845 16052 23584
rect 16107 22280 16149 22289
rect 16107 22240 16108 22280
rect 16148 22240 16149 22280
rect 16107 22231 16149 22240
rect 16108 21608 16148 22231
rect 16108 21559 16148 21568
rect 16107 21440 16149 21449
rect 16107 21400 16108 21440
rect 16148 21400 16149 21440
rect 16107 21391 16149 21400
rect 16108 20861 16148 21391
rect 16107 20852 16149 20861
rect 16107 20812 16108 20852
rect 16148 20812 16149 20852
rect 16107 20803 16149 20812
rect 16204 20180 16244 33487
rect 16300 33293 16340 35092
rect 16396 36728 16436 38200
rect 16396 33620 16436 36688
rect 16684 38744 16724 38753
rect 16587 36644 16629 36653
rect 16587 36604 16588 36644
rect 16628 36604 16629 36644
rect 16587 36595 16629 36604
rect 16492 35888 16532 35899
rect 16492 35813 16532 35848
rect 16491 35804 16533 35813
rect 16491 35764 16492 35804
rect 16532 35764 16533 35804
rect 16491 35755 16533 35764
rect 16492 35048 16532 35057
rect 16588 35048 16628 36595
rect 16684 36317 16724 38704
rect 16683 36308 16725 36317
rect 16683 36268 16684 36308
rect 16724 36268 16725 36308
rect 16683 36259 16725 36268
rect 16683 36140 16725 36149
rect 16683 36100 16684 36140
rect 16724 36100 16725 36140
rect 16683 36091 16725 36100
rect 16684 36006 16724 36091
rect 16532 35008 16628 35048
rect 16684 35132 16724 35141
rect 16492 34999 16532 35008
rect 16684 34805 16724 35092
rect 16683 34796 16725 34805
rect 16683 34756 16684 34796
rect 16724 34756 16725 34796
rect 16683 34747 16725 34756
rect 16491 34376 16533 34385
rect 16491 34336 16492 34376
rect 16532 34336 16533 34376
rect 16491 34327 16533 34336
rect 16492 34242 16532 34327
rect 16683 34208 16725 34217
rect 16683 34168 16684 34208
rect 16724 34168 16725 34208
rect 16683 34159 16725 34168
rect 16684 34074 16724 34159
rect 16587 33956 16629 33965
rect 16587 33916 16588 33956
rect 16628 33916 16629 33956
rect 16587 33907 16629 33916
rect 16492 33620 16532 33629
rect 16396 33580 16492 33620
rect 16492 33461 16532 33580
rect 16588 33620 16628 33907
rect 16491 33452 16533 33461
rect 16491 33412 16492 33452
rect 16532 33412 16533 33452
rect 16491 33403 16533 33412
rect 16299 33284 16341 33293
rect 16299 33244 16300 33284
rect 16340 33244 16341 33284
rect 16299 33235 16341 33244
rect 16588 32873 16628 33580
rect 16587 32864 16629 32873
rect 16587 32824 16588 32864
rect 16628 32824 16629 32864
rect 16587 32815 16629 32824
rect 16684 32864 16724 32875
rect 16684 32789 16724 32824
rect 16683 32780 16725 32789
rect 16683 32740 16684 32780
rect 16724 32740 16725 32780
rect 16683 32731 16725 32740
rect 16491 32444 16533 32453
rect 16491 32404 16492 32444
rect 16532 32404 16533 32444
rect 16491 32395 16533 32404
rect 16492 32360 16532 32395
rect 16492 32309 16532 32320
rect 16300 32178 16340 32187
rect 16300 31604 16340 32138
rect 16684 32108 16724 32117
rect 16300 31555 16340 31564
rect 16588 32068 16684 32108
rect 16491 31436 16533 31445
rect 16491 31396 16492 31436
rect 16532 31396 16533 31436
rect 16491 31387 16533 31396
rect 16492 31352 16532 31387
rect 16492 31301 16532 31312
rect 16299 30008 16341 30017
rect 16299 29968 16300 30008
rect 16340 29968 16341 30008
rect 16299 29959 16341 29968
rect 16300 29874 16340 29959
rect 16492 29924 16532 29933
rect 16492 29429 16532 29884
rect 16491 29420 16533 29429
rect 16491 29380 16492 29420
rect 16532 29380 16533 29420
rect 16491 29371 16533 29380
rect 16588 29177 16628 32068
rect 16684 32059 16724 32068
rect 16684 30092 16724 30101
rect 16780 30092 16820 40048
rect 17068 39668 17108 40207
rect 17068 39619 17108 39628
rect 16875 39500 16917 39509
rect 16875 39460 16876 39500
rect 16916 39460 16917 39500
rect 16875 39451 16917 39460
rect 16876 39366 16916 39451
rect 17164 39257 17204 40384
rect 17260 39593 17300 40468
rect 17259 39584 17301 39593
rect 17259 39544 17260 39584
rect 17300 39544 17301 39584
rect 17259 39535 17301 39544
rect 17260 39450 17300 39535
rect 17163 39248 17205 39257
rect 17163 39208 17164 39248
rect 17204 39208 17205 39248
rect 17356 39248 17396 42307
rect 17451 41852 17493 41861
rect 17451 41812 17452 41852
rect 17492 41812 17493 41852
rect 17451 41803 17493 41812
rect 17452 40676 17492 41803
rect 17548 41693 17588 42928
rect 17740 41768 17780 42928
rect 17835 42272 17877 42281
rect 17835 42232 17836 42272
rect 17876 42232 17877 42272
rect 17835 42223 17877 42232
rect 17644 41728 17780 41768
rect 17547 41684 17589 41693
rect 17547 41644 17548 41684
rect 17588 41644 17589 41684
rect 17547 41635 17589 41644
rect 17644 40853 17684 41728
rect 17739 41600 17781 41609
rect 17739 41560 17740 41600
rect 17780 41560 17781 41600
rect 17739 41551 17781 41560
rect 17643 40844 17685 40853
rect 17643 40804 17644 40844
rect 17684 40804 17685 40844
rect 17643 40795 17685 40804
rect 17452 40627 17492 40636
rect 17644 40592 17684 40601
rect 17644 40433 17684 40552
rect 17643 40424 17685 40433
rect 17643 40384 17644 40424
rect 17684 40384 17685 40424
rect 17643 40375 17685 40384
rect 17740 40088 17780 41551
rect 17836 40508 17876 42223
rect 17932 41609 17972 42928
rect 18124 42029 18164 42928
rect 18219 42188 18261 42197
rect 18219 42148 18220 42188
rect 18260 42148 18261 42188
rect 18219 42139 18261 42148
rect 18123 42020 18165 42029
rect 18123 41980 18124 42020
rect 18164 41980 18165 42020
rect 18123 41971 18165 41980
rect 17931 41600 17973 41609
rect 17931 41560 17932 41600
rect 17972 41560 17973 41600
rect 17931 41551 17973 41560
rect 17836 40459 17876 40468
rect 17932 41264 17972 41273
rect 17835 40340 17877 40349
rect 17835 40300 17836 40340
rect 17876 40300 17877 40340
rect 17835 40291 17877 40300
rect 17644 40048 17780 40088
rect 17547 39920 17589 39929
rect 17547 39880 17548 39920
rect 17588 39880 17589 39920
rect 17547 39871 17589 39880
rect 17548 39786 17588 39871
rect 17356 39208 17492 39248
rect 17163 39199 17205 39208
rect 17452 39164 17492 39208
rect 17452 39115 17492 39124
rect 16971 39080 17013 39089
rect 16971 39040 16972 39080
rect 17012 39040 17013 39080
rect 16971 39031 17013 39040
rect 17644 39080 17684 40048
rect 17739 39668 17781 39677
rect 17739 39628 17740 39668
rect 17780 39628 17781 39668
rect 17739 39619 17781 39628
rect 17740 39534 17780 39619
rect 17836 39164 17876 40291
rect 17644 39031 17684 39040
rect 17740 39124 17876 39164
rect 16876 38996 16916 39005
rect 16876 38753 16916 38956
rect 16875 38744 16917 38753
rect 16875 38704 16876 38744
rect 16916 38704 16917 38744
rect 16875 38695 16917 38704
rect 16876 38226 16916 38235
rect 16876 37745 16916 38186
rect 16875 37736 16917 37745
rect 16875 37696 16876 37736
rect 16916 37696 16917 37736
rect 16875 37687 16917 37696
rect 16876 37400 16916 37409
rect 16876 37157 16916 37360
rect 16875 37148 16917 37157
rect 16875 37108 16876 37148
rect 16916 37108 16917 37148
rect 16875 37099 16917 37108
rect 16876 36714 16916 36723
rect 16876 36149 16916 36674
rect 16875 36140 16917 36149
rect 16875 36100 16876 36140
rect 16916 36100 16917 36140
rect 16875 36091 16917 36100
rect 16875 35972 16917 35981
rect 16875 35932 16876 35972
rect 16916 35932 16917 35972
rect 16875 35923 16917 35932
rect 16876 35888 16916 35923
rect 16876 35837 16916 35848
rect 16875 35468 16917 35477
rect 16875 35428 16876 35468
rect 16916 35428 16917 35468
rect 16875 35419 16917 35428
rect 16876 35048 16916 35419
rect 16876 34999 16916 35008
rect 16876 34376 16916 34387
rect 16876 34301 16916 34336
rect 16875 34292 16917 34301
rect 16875 34252 16876 34292
rect 16916 34252 16917 34292
rect 16875 34243 16917 34252
rect 16972 33125 17012 39031
rect 17260 38996 17300 39005
rect 17300 38956 17396 38996
rect 17260 38947 17300 38956
rect 17067 38744 17109 38753
rect 17067 38704 17068 38744
rect 17108 38704 17109 38744
rect 17067 38695 17109 38704
rect 17068 38610 17108 38695
rect 17068 38408 17108 38417
rect 17108 38368 17204 38408
rect 17068 38359 17108 38368
rect 17067 37736 17109 37745
rect 17067 37696 17068 37736
rect 17108 37696 17109 37736
rect 17067 37687 17109 37696
rect 17068 37652 17108 37687
rect 17068 37601 17108 37612
rect 17164 37493 17204 38368
rect 17356 38081 17396 38956
rect 17740 38753 17780 39124
rect 17836 38996 17876 39005
rect 17932 38996 17972 41224
rect 18124 41012 18164 41021
rect 18027 40508 18069 40517
rect 18027 40468 18028 40508
rect 18068 40468 18069 40508
rect 18027 40459 18069 40468
rect 18028 40374 18068 40459
rect 18028 39677 18068 39708
rect 18027 39668 18069 39677
rect 18027 39628 18028 39668
rect 18068 39628 18069 39668
rect 18027 39619 18069 39628
rect 18028 39584 18068 39619
rect 18028 39257 18068 39544
rect 18027 39248 18069 39257
rect 18027 39208 18028 39248
rect 18068 39208 18069 39248
rect 18027 39199 18069 39208
rect 18124 39173 18164 40972
rect 18220 40340 18260 42139
rect 18316 41684 18356 42928
rect 18316 41644 18452 41684
rect 18316 41096 18356 41105
rect 18316 40937 18356 41056
rect 18315 40928 18357 40937
rect 18315 40888 18316 40928
rect 18356 40888 18357 40928
rect 18315 40879 18357 40888
rect 18316 40676 18356 40685
rect 18412 40676 18452 41644
rect 18508 41609 18548 42928
rect 18700 42197 18740 42928
rect 18699 42188 18741 42197
rect 18699 42148 18700 42188
rect 18740 42148 18741 42188
rect 18699 42139 18741 42148
rect 18892 42113 18932 42928
rect 18603 42104 18645 42113
rect 18603 42064 18604 42104
rect 18644 42064 18645 42104
rect 18603 42055 18645 42064
rect 18891 42104 18933 42113
rect 18891 42064 18892 42104
rect 18932 42064 18933 42104
rect 18891 42055 18933 42064
rect 18507 41600 18549 41609
rect 18507 41560 18508 41600
rect 18548 41560 18549 41600
rect 18507 41551 18549 41560
rect 18604 41432 18644 42055
rect 18987 41936 19029 41945
rect 18987 41896 18988 41936
rect 19028 41896 19029 41936
rect 18987 41887 19029 41896
rect 18699 41684 18741 41693
rect 18699 41644 18700 41684
rect 18740 41644 18741 41684
rect 18699 41635 18741 41644
rect 18604 41383 18644 41392
rect 18507 40928 18549 40937
rect 18507 40888 18508 40928
rect 18548 40888 18549 40928
rect 18507 40879 18549 40888
rect 18356 40636 18452 40676
rect 18316 40627 18356 40636
rect 18508 40508 18548 40879
rect 18700 40844 18740 41635
rect 18988 41432 19028 41887
rect 19084 41861 19124 42928
rect 19083 41852 19125 41861
rect 19083 41812 19084 41852
rect 19124 41812 19125 41852
rect 19083 41803 19125 41812
rect 18988 41383 19028 41392
rect 18795 41348 18837 41357
rect 18795 41308 18796 41348
rect 18836 41308 18837 41348
rect 18795 41299 18837 41308
rect 18796 41180 18836 41299
rect 18796 41131 18836 41140
rect 19180 41180 19220 41189
rect 19180 41021 19220 41140
rect 19179 41012 19221 41021
rect 19179 40972 19180 41012
rect 19220 40972 19221 41012
rect 19179 40963 19221 40972
rect 18508 40459 18548 40468
rect 18604 40804 18740 40844
rect 18808 40844 19176 40853
rect 18848 40804 18890 40844
rect 18930 40804 18972 40844
rect 19012 40804 19054 40844
rect 19094 40804 19136 40844
rect 18220 40300 18548 40340
rect 18411 39920 18453 39929
rect 18411 39880 18412 39920
rect 18452 39880 18453 39920
rect 18411 39871 18453 39880
rect 18412 39786 18452 39871
rect 18220 39668 18260 39677
rect 18123 39164 18165 39173
rect 18123 39124 18124 39164
rect 18164 39124 18165 39164
rect 18123 39115 18165 39124
rect 17876 38956 17972 38996
rect 17739 38744 17781 38753
rect 17739 38704 17740 38744
rect 17780 38704 17781 38744
rect 17739 38695 17781 38704
rect 17836 38249 17876 38956
rect 18220 38753 18260 39628
rect 18508 39080 18548 40300
rect 18604 39920 18644 40804
rect 18808 40795 19176 40804
rect 19083 40676 19125 40685
rect 19276 40676 19316 42928
rect 19468 42533 19508 42928
rect 19467 42524 19509 42533
rect 19467 42484 19468 42524
rect 19508 42484 19509 42524
rect 19467 42475 19509 42484
rect 19467 42104 19509 42113
rect 19467 42064 19468 42104
rect 19508 42064 19509 42104
rect 19467 42055 19509 42064
rect 19371 41432 19413 41441
rect 19371 41392 19372 41432
rect 19412 41392 19413 41432
rect 19371 41383 19413 41392
rect 19372 41298 19412 41383
rect 19371 40760 19413 40769
rect 19371 40720 19372 40760
rect 19412 40720 19413 40760
rect 19371 40711 19413 40720
rect 19083 40636 19084 40676
rect 19124 40636 19125 40676
rect 19083 40627 19125 40636
rect 19180 40636 19316 40676
rect 18699 40592 18741 40601
rect 18699 40552 18700 40592
rect 18740 40552 18741 40592
rect 18699 40543 18741 40552
rect 18700 40458 18740 40543
rect 19084 40542 19124 40627
rect 18891 40508 18933 40517
rect 18891 40468 18892 40508
rect 18932 40468 18933 40508
rect 18891 40459 18933 40468
rect 18892 40374 18932 40459
rect 18699 40256 18741 40265
rect 18699 40216 18700 40256
rect 18740 40216 18741 40256
rect 18699 40207 18741 40216
rect 18604 39871 18644 39880
rect 18700 39164 18740 40207
rect 18987 40088 19029 40097
rect 18987 40048 18988 40088
rect 19028 40048 19029 40088
rect 18987 40039 19029 40048
rect 18988 39920 19028 40039
rect 19180 39929 19220 40636
rect 19372 40592 19412 40711
rect 19468 40676 19508 42055
rect 19851 42020 19893 42029
rect 19851 41980 19852 42020
rect 19892 41980 19893 42020
rect 19851 41971 19893 41980
rect 19563 41180 19605 41189
rect 19563 41140 19564 41180
rect 19604 41140 19605 41180
rect 19563 41131 19605 41140
rect 19756 41180 19796 41189
rect 19564 41046 19604 41131
rect 19756 41021 19796 41140
rect 19755 41012 19797 41021
rect 19755 40972 19756 41012
rect 19796 40972 19797 41012
rect 19755 40963 19797 40972
rect 19468 40627 19508 40636
rect 19852 40676 19892 41971
rect 20048 41600 20416 41609
rect 20088 41560 20130 41600
rect 20170 41560 20212 41600
rect 20252 41560 20294 41600
rect 20334 41560 20376 41600
rect 20048 41551 20416 41560
rect 19948 41012 19988 41021
rect 19948 40769 19988 40972
rect 19947 40760 19989 40769
rect 19947 40720 19948 40760
rect 19988 40720 19989 40760
rect 19947 40711 19989 40720
rect 19852 40627 19892 40636
rect 19276 40552 19412 40592
rect 19276 40508 19316 40552
rect 19276 40459 19316 40468
rect 19659 40508 19701 40517
rect 20044 40508 20084 40517
rect 19659 40468 19660 40508
rect 19700 40468 19701 40508
rect 19659 40459 19701 40468
rect 19948 40468 20044 40508
rect 19660 40374 19700 40459
rect 19755 40172 19797 40181
rect 19755 40132 19756 40172
rect 19796 40132 19797 40172
rect 19755 40123 19797 40132
rect 18988 39871 19028 39880
rect 19179 39920 19221 39929
rect 19179 39880 19180 39920
rect 19220 39880 19221 39920
rect 19179 39871 19221 39880
rect 18795 39668 18837 39677
rect 18795 39628 18796 39668
rect 18836 39628 18837 39668
rect 18795 39619 18837 39628
rect 19180 39668 19220 39677
rect 19372 39668 19412 39677
rect 19220 39628 19316 39668
rect 19180 39619 19220 39628
rect 18796 39534 18836 39619
rect 18808 39332 19176 39341
rect 18848 39292 18890 39332
rect 18930 39292 18972 39332
rect 19012 39292 19054 39332
rect 19094 39292 19136 39332
rect 18808 39283 19176 39292
rect 19276 39248 19316 39628
rect 19372 39425 19412 39628
rect 19756 39668 19796 40123
rect 19948 39677 19988 40468
rect 20044 40459 20084 40468
rect 20048 40088 20416 40097
rect 20088 40048 20130 40088
rect 20170 40048 20212 40088
rect 20252 40048 20294 40088
rect 20334 40048 20376 40088
rect 20048 40039 20416 40048
rect 21003 39752 21045 39761
rect 21003 39712 21004 39752
rect 21044 39712 21045 39752
rect 21003 39703 21045 39712
rect 19756 39619 19796 39628
rect 19947 39668 19989 39677
rect 19947 39628 19948 39668
rect 19988 39628 19989 39668
rect 19947 39619 19989 39628
rect 20139 39584 20181 39593
rect 20139 39544 20140 39584
rect 20180 39544 20181 39584
rect 20139 39535 20181 39544
rect 19563 39500 19605 39509
rect 19563 39460 19564 39500
rect 19604 39460 19605 39500
rect 19563 39451 19605 39460
rect 19948 39500 19988 39509
rect 19371 39416 19413 39425
rect 19371 39376 19372 39416
rect 19412 39376 19413 39416
rect 19371 39367 19413 39376
rect 19564 39366 19604 39451
rect 19276 39208 19412 39248
rect 19179 39164 19221 39173
rect 18700 39124 18836 39164
rect 18508 39031 18548 39040
rect 18700 38996 18740 39005
rect 18604 38956 18700 38996
rect 18219 38744 18261 38753
rect 18219 38704 18220 38744
rect 18260 38704 18261 38744
rect 18219 38695 18261 38704
rect 18220 38610 18260 38695
rect 18411 38324 18453 38333
rect 18411 38284 18412 38324
rect 18452 38284 18453 38324
rect 18411 38275 18453 38284
rect 17451 38240 17493 38249
rect 17835 38240 17877 38249
rect 17451 38200 17452 38240
rect 17492 38200 17588 38240
rect 17451 38191 17493 38200
rect 17452 38106 17492 38191
rect 17355 38072 17397 38081
rect 17355 38032 17356 38072
rect 17396 38032 17397 38072
rect 17355 38023 17397 38032
rect 17259 37988 17301 37997
rect 17259 37948 17260 37988
rect 17300 37948 17301 37988
rect 17259 37939 17301 37948
rect 17260 37854 17300 37939
rect 17355 37904 17397 37913
rect 17355 37864 17356 37904
rect 17396 37864 17397 37904
rect 17355 37855 17397 37864
rect 17163 37484 17205 37493
rect 17163 37444 17164 37484
rect 17204 37444 17205 37484
rect 17163 37435 17205 37444
rect 17260 37484 17300 37495
rect 17260 37409 17300 37444
rect 17259 37400 17301 37409
rect 17259 37360 17260 37400
rect 17300 37360 17301 37400
rect 17259 37351 17301 37360
rect 17067 36896 17109 36905
rect 17067 36856 17068 36896
rect 17108 36856 17109 36896
rect 17067 36847 17109 36856
rect 17068 36762 17108 36847
rect 17356 36653 17396 37855
rect 17451 37568 17493 37577
rect 17451 37528 17452 37568
rect 17492 37528 17493 37568
rect 17451 37519 17493 37528
rect 17452 37434 17492 37519
rect 17452 36728 17492 36737
rect 17548 36728 17588 38200
rect 17835 38200 17836 38240
rect 17876 38200 17877 38240
rect 17835 38191 17877 38200
rect 17739 37988 17781 37997
rect 17739 37948 17740 37988
rect 17780 37948 17781 37988
rect 17739 37939 17781 37948
rect 17740 37400 17780 37939
rect 18219 37484 18261 37493
rect 18219 37444 18220 37484
rect 18260 37444 18261 37484
rect 18219 37435 18261 37444
rect 17740 37351 17780 37360
rect 17835 37400 17877 37409
rect 17835 37360 17836 37400
rect 17876 37360 17877 37400
rect 17835 37351 17877 37360
rect 17836 37266 17876 37351
rect 18123 37148 18165 37157
rect 18123 37108 18124 37148
rect 18164 37108 18165 37148
rect 18123 37099 18165 37108
rect 17835 36896 17877 36905
rect 17835 36856 17836 36896
rect 17876 36856 17877 36896
rect 17835 36847 17877 36856
rect 17492 36688 17684 36728
rect 17452 36679 17492 36688
rect 17355 36644 17397 36653
rect 17355 36604 17356 36644
rect 17396 36604 17397 36644
rect 17355 36595 17397 36604
rect 17260 36476 17300 36485
rect 17300 36436 17588 36476
rect 17260 36427 17300 36436
rect 17451 36308 17493 36317
rect 17451 36268 17452 36308
rect 17492 36268 17493 36308
rect 17451 36259 17493 36268
rect 17067 35804 17109 35813
rect 17067 35764 17068 35804
rect 17108 35764 17109 35804
rect 17067 35755 17109 35764
rect 17068 35132 17108 35755
rect 17068 35057 17108 35092
rect 17067 35048 17109 35057
rect 17067 35008 17068 35048
rect 17108 35008 17109 35048
rect 17067 34999 17109 35008
rect 17259 35048 17301 35057
rect 17259 35008 17260 35048
rect 17300 35008 17301 35048
rect 17259 34999 17301 35008
rect 17260 34914 17300 34999
rect 17355 34544 17397 34553
rect 17355 34504 17356 34544
rect 17396 34504 17397 34544
rect 17355 34495 17397 34504
rect 17067 33704 17109 33713
rect 17067 33664 17068 33704
rect 17108 33664 17109 33704
rect 17067 33655 17109 33664
rect 17068 33570 17108 33655
rect 16971 33116 17013 33125
rect 16971 33076 16972 33116
rect 17012 33076 17013 33116
rect 16971 33067 17013 33076
rect 17356 33041 17396 34495
rect 17355 33032 17397 33041
rect 17355 32992 17356 33032
rect 17396 32992 17397 33032
rect 17355 32983 17397 32992
rect 17164 32864 17204 32873
rect 16972 32824 17164 32864
rect 16876 32780 16916 32789
rect 16972 32780 17012 32824
rect 17164 32815 17204 32824
rect 17260 32864 17300 32873
rect 17300 32824 17396 32864
rect 17260 32815 17300 32824
rect 16916 32740 17012 32780
rect 16876 32731 16916 32740
rect 17259 32612 17301 32621
rect 17259 32572 17260 32612
rect 17300 32572 17301 32612
rect 17259 32563 17301 32572
rect 16875 32360 16917 32369
rect 16875 32320 16876 32360
rect 16916 32320 16917 32360
rect 16875 32311 16917 32320
rect 17260 32360 17300 32563
rect 17260 32311 17300 32320
rect 16876 32226 16916 32311
rect 17068 32108 17108 32117
rect 17068 31361 17108 32068
rect 17067 31352 17109 31361
rect 17067 31312 17068 31352
rect 17108 31312 17109 31352
rect 17067 31303 17109 31312
rect 16971 30680 17013 30689
rect 16971 30640 16972 30680
rect 17012 30640 17013 30680
rect 16971 30631 17013 30640
rect 16724 30052 16820 30092
rect 16684 30043 16724 30052
rect 16492 29168 16532 29177
rect 16299 28916 16341 28925
rect 16299 28876 16300 28916
rect 16340 28876 16341 28916
rect 16299 28867 16341 28876
rect 16300 27651 16340 28867
rect 16492 28748 16532 29128
rect 16587 29168 16629 29177
rect 16587 29128 16588 29168
rect 16628 29128 16629 29168
rect 16972 29168 17012 30631
rect 17164 30428 17204 30437
rect 17164 29840 17204 30388
rect 17164 29791 17204 29800
rect 17259 29840 17301 29849
rect 17259 29800 17260 29840
rect 17300 29800 17301 29840
rect 17259 29791 17301 29800
rect 17260 29706 17300 29791
rect 17356 29345 17396 32824
rect 17452 32537 17492 36259
rect 17548 35216 17588 36436
rect 17644 35981 17684 36688
rect 17643 35972 17685 35981
rect 17643 35932 17644 35972
rect 17684 35932 17685 35972
rect 17643 35923 17685 35932
rect 17548 35167 17588 35176
rect 17643 35216 17685 35225
rect 17643 35176 17644 35216
rect 17684 35176 17685 35216
rect 17643 35167 17685 35176
rect 17644 35082 17684 35167
rect 17643 34712 17685 34721
rect 17643 34672 17644 34712
rect 17684 34672 17685 34712
rect 17643 34663 17685 34672
rect 17547 33704 17589 33713
rect 17547 33659 17548 33704
rect 17588 33659 17589 33704
rect 17547 33655 17589 33659
rect 17548 33569 17588 33655
rect 17644 33452 17684 34663
rect 17739 34460 17781 34469
rect 17739 34420 17740 34460
rect 17780 34420 17781 34460
rect 17739 34411 17781 34420
rect 17740 33872 17780 34411
rect 17740 33823 17780 33832
rect 17644 33412 17780 33452
rect 17740 32948 17780 33412
rect 17740 32873 17780 32908
rect 17547 32864 17589 32873
rect 17644 32864 17684 32873
rect 17547 32824 17548 32864
rect 17588 32824 17644 32864
rect 17547 32815 17589 32824
rect 17644 32815 17684 32824
rect 17739 32864 17781 32873
rect 17739 32824 17740 32864
rect 17780 32824 17781 32864
rect 17739 32815 17781 32824
rect 17451 32528 17493 32537
rect 17451 32488 17452 32528
rect 17492 32488 17493 32528
rect 17451 32479 17493 32488
rect 17451 32360 17493 32369
rect 17451 32320 17452 32360
rect 17492 32320 17493 32360
rect 17451 32311 17493 32320
rect 17452 32192 17492 32311
rect 17355 29336 17397 29345
rect 17355 29296 17356 29336
rect 17396 29296 17397 29336
rect 17355 29287 17397 29296
rect 17068 29168 17108 29177
rect 16972 29128 17068 29168
rect 16587 29119 16629 29128
rect 17068 29119 17108 29128
rect 17452 29000 17492 32152
rect 17164 28960 17492 29000
rect 16683 28916 16725 28925
rect 16683 28876 16684 28916
rect 16724 28876 16725 28916
rect 16683 28867 16725 28876
rect 16876 28916 16916 28925
rect 16684 28782 16724 28867
rect 16492 28708 16543 28748
rect 16503 28580 16543 28708
rect 16492 28540 16543 28580
rect 16492 28328 16532 28540
rect 16876 28505 16916 28876
rect 16875 28496 16917 28505
rect 16875 28456 16876 28496
rect 16916 28456 16917 28496
rect 16875 28447 16917 28456
rect 16395 28244 16437 28253
rect 16395 28204 16396 28244
rect 16436 28204 16437 28244
rect 16395 28195 16437 28204
rect 16300 27602 16340 27611
rect 16300 25901 16340 25986
rect 16299 25892 16341 25901
rect 16299 25852 16300 25892
rect 16340 25852 16341 25892
rect 16299 25843 16341 25852
rect 16299 25640 16341 25649
rect 16299 25600 16300 25640
rect 16340 25600 16341 25640
rect 16299 25591 16341 25600
rect 16300 24473 16340 25591
rect 16396 25304 16436 28195
rect 16492 28001 16532 28288
rect 17068 28412 17108 28421
rect 17068 28169 17108 28372
rect 16684 28160 16724 28169
rect 16588 28120 16684 28160
rect 16491 27992 16533 28001
rect 16491 27952 16492 27992
rect 16532 27952 16533 27992
rect 16491 27943 16533 27952
rect 16492 27740 16532 27751
rect 16492 27665 16532 27700
rect 16491 27656 16533 27665
rect 16491 27616 16492 27656
rect 16532 27616 16533 27656
rect 16491 27607 16533 27616
rect 16588 26816 16628 28120
rect 16684 28111 16724 28120
rect 17067 28160 17109 28169
rect 17067 28120 17068 28160
rect 17108 28120 17109 28160
rect 17067 28111 17109 28120
rect 16683 27908 16725 27917
rect 16683 27868 16684 27908
rect 16724 27868 16725 27908
rect 16683 27859 16725 27868
rect 17067 27908 17109 27917
rect 17067 27868 17068 27908
rect 17108 27868 17109 27908
rect 17067 27859 17109 27868
rect 16684 27656 16724 27859
rect 16724 27616 16820 27656
rect 16684 27607 16724 27616
rect 16588 26767 16628 26776
rect 16684 26816 16724 26825
rect 16684 26480 16724 26776
rect 16588 26440 16724 26480
rect 16491 25892 16533 25901
rect 16491 25852 16492 25892
rect 16532 25852 16533 25892
rect 16491 25843 16533 25852
rect 16299 24464 16341 24473
rect 16299 24424 16300 24464
rect 16340 24424 16341 24464
rect 16299 24415 16341 24424
rect 16396 22877 16436 25264
rect 16492 24632 16532 25843
rect 16492 24583 16532 24592
rect 16588 24632 16628 26440
rect 16491 24464 16533 24473
rect 16491 24424 16492 24464
rect 16532 24424 16533 24464
rect 16491 24415 16533 24424
rect 16395 22868 16437 22877
rect 16395 22828 16396 22868
rect 16436 22828 16437 22868
rect 16395 22819 16437 22828
rect 16492 22700 16532 24415
rect 16396 22660 16532 22700
rect 16300 21449 16340 21534
rect 16299 21440 16341 21449
rect 16299 21400 16300 21440
rect 16340 21400 16341 21440
rect 16299 21391 16341 21400
rect 16396 21020 16436 22660
rect 16491 22532 16533 22541
rect 16491 22492 16492 22532
rect 16532 22492 16533 22532
rect 16491 22483 16533 22492
rect 16300 20980 16436 21020
rect 16492 22280 16532 22483
rect 16300 20684 16340 20980
rect 16396 20861 16436 20877
rect 16395 20852 16437 20861
rect 16395 20812 16396 20852
rect 16436 20812 16437 20852
rect 16395 20803 16437 20812
rect 16396 20782 16436 20803
rect 16396 20733 16436 20742
rect 16300 20644 16436 20684
rect 16108 20140 16244 20180
rect 16011 18836 16053 18845
rect 16011 18796 16012 18836
rect 16052 18796 16053 18836
rect 16011 18787 16053 18796
rect 16011 18584 16053 18593
rect 16011 18544 16012 18584
rect 16052 18544 16053 18584
rect 16011 18535 16053 18544
rect 16012 18257 16052 18535
rect 16011 18248 16053 18257
rect 16011 18208 16012 18248
rect 16052 18208 16053 18248
rect 16011 18199 16053 18208
rect 16011 17996 16053 18005
rect 16011 17956 16012 17996
rect 16052 17956 16053 17996
rect 16011 17947 16053 17956
rect 16012 17862 16052 17947
rect 16011 17744 16053 17753
rect 16011 17704 16012 17744
rect 16052 17704 16053 17744
rect 16011 17695 16053 17704
rect 16012 17610 16052 17695
rect 15916 17200 16052 17240
rect 15668 17032 15860 17072
rect 15916 17072 15956 17081
rect 15340 16938 15380 17023
rect 15628 16652 15668 17032
rect 15916 16745 15956 17032
rect 15915 16736 15957 16745
rect 15915 16696 15916 16736
rect 15956 16696 15957 16736
rect 15915 16687 15957 16696
rect 15436 16612 15668 16652
rect 15436 16232 15476 16612
rect 15627 16484 15669 16493
rect 15627 16444 15628 16484
rect 15668 16444 15669 16484
rect 15627 16435 15669 16444
rect 15339 15056 15381 15065
rect 15339 15016 15340 15056
rect 15380 15016 15381 15056
rect 15339 15007 15381 15016
rect 15243 14720 15285 14729
rect 15243 14680 15244 14720
rect 15284 14680 15285 14720
rect 15243 14671 15285 14680
rect 15340 14720 15380 15007
rect 15340 14671 15380 14680
rect 15148 14428 15380 14468
rect 14859 14419 14901 14428
rect 14763 14300 14805 14309
rect 14763 14260 14764 14300
rect 14804 14260 14805 14300
rect 14763 14251 14805 14260
rect 14667 14048 14709 14057
rect 14667 14008 14668 14048
rect 14708 14008 14709 14048
rect 14667 13999 14709 14008
rect 14764 14048 14804 14059
rect 14668 13460 14708 13999
rect 14764 13973 14804 14008
rect 14763 13964 14805 13973
rect 14763 13924 14764 13964
rect 14804 13924 14805 13964
rect 14763 13915 14805 13924
rect 14668 13411 14708 13420
rect 14763 13208 14805 13217
rect 14763 13168 14764 13208
rect 14804 13168 14805 13208
rect 14763 13159 14805 13168
rect 14764 13074 14804 13159
rect 14860 12041 14900 14419
rect 14955 14216 14997 14225
rect 14955 14176 14956 14216
rect 14996 14176 14997 14216
rect 14955 14167 14997 14176
rect 14956 14048 14996 14167
rect 14956 13999 14996 14008
rect 14955 13880 14997 13889
rect 14955 13840 14956 13880
rect 14996 13840 14997 13880
rect 14955 13831 14997 13840
rect 14859 12032 14901 12041
rect 14859 11992 14860 12032
rect 14900 11992 14901 12032
rect 14859 11983 14901 11992
rect 14571 11864 14613 11873
rect 14571 11824 14572 11864
rect 14612 11824 14613 11864
rect 14571 11815 14613 11824
rect 14859 11864 14901 11873
rect 14859 11824 14860 11864
rect 14900 11824 14901 11864
rect 14859 11815 14901 11824
rect 14284 11696 14324 11707
rect 14284 11621 14324 11656
rect 14380 11696 14420 11705
rect 14283 11612 14325 11621
rect 14283 11572 14284 11612
rect 14324 11572 14325 11612
rect 14283 11563 14325 11572
rect 14380 11537 14420 11656
rect 14475 11696 14517 11705
rect 14475 11656 14476 11696
rect 14516 11656 14517 11696
rect 14475 11647 14517 11656
rect 14476 11562 14516 11647
rect 14379 11528 14421 11537
rect 14379 11488 14380 11528
rect 14420 11488 14421 11528
rect 14379 11479 14421 11488
rect 14572 11528 14612 11537
rect 14475 11444 14517 11453
rect 14475 11404 14476 11444
rect 14516 11404 14517 11444
rect 14475 11395 14517 11404
rect 14187 10520 14229 10529
rect 14187 10480 14188 10520
rect 14228 10480 14229 10520
rect 14187 10471 14229 10480
rect 14476 10352 14516 11395
rect 14572 11201 14612 11488
rect 14571 11192 14613 11201
rect 14571 11152 14572 11192
rect 14612 11152 14613 11192
rect 14571 11143 14613 11152
rect 14571 10688 14613 10697
rect 14571 10648 14572 10688
rect 14612 10648 14613 10688
rect 14571 10639 14613 10648
rect 14380 10312 14516 10352
rect 14092 9724 14228 9764
rect 13803 9680 13845 9689
rect 13803 9640 13804 9680
rect 13844 9640 13845 9680
rect 13803 9631 13845 9640
rect 13707 9176 13749 9185
rect 13707 9136 13708 9176
rect 13748 9136 13749 9176
rect 13707 9127 13749 9136
rect 13611 6908 13653 6917
rect 13611 6868 13612 6908
rect 13652 6868 13653 6908
rect 13611 6859 13653 6868
rect 13804 6833 13844 9631
rect 13996 9512 14036 9521
rect 13996 8429 14036 9472
rect 14091 9428 14133 9437
rect 14091 9388 14092 9428
rect 14132 9388 14133 9428
rect 14091 9379 14133 9388
rect 13995 8420 14037 8429
rect 13995 8380 13996 8420
rect 14036 8380 14037 8420
rect 13995 8371 14037 8380
rect 13900 8009 13940 8094
rect 13899 8000 13941 8009
rect 13899 7960 13900 8000
rect 13940 7960 14036 8000
rect 13899 7951 13941 7960
rect 13899 7832 13941 7841
rect 13899 7792 13900 7832
rect 13940 7792 13941 7832
rect 13899 7783 13941 7792
rect 13803 6824 13845 6833
rect 13803 6784 13804 6824
rect 13844 6784 13845 6824
rect 13803 6775 13845 6784
rect 13516 6532 13748 6572
rect 13419 6488 13461 6497
rect 13419 6448 13420 6488
rect 13460 6448 13461 6488
rect 13419 6439 13461 6448
rect 13516 6404 13556 6413
rect 13516 6320 13556 6364
rect 13420 6280 13556 6320
rect 13420 5993 13460 6280
rect 13419 5984 13461 5993
rect 13419 5944 13420 5984
rect 13460 5944 13461 5984
rect 13419 5935 13461 5944
rect 13611 5984 13653 5993
rect 13611 5944 13612 5984
rect 13652 5944 13653 5984
rect 13611 5935 13653 5944
rect 13419 5732 13461 5741
rect 13419 5692 13420 5732
rect 13460 5692 13461 5732
rect 13419 5683 13461 5692
rect 13324 4087 13364 4096
rect 13420 3893 13460 5683
rect 13612 4976 13652 5935
rect 13708 5573 13748 6532
rect 13804 6497 13844 6775
rect 13803 6488 13845 6497
rect 13803 6448 13804 6488
rect 13844 6448 13845 6488
rect 13803 6439 13845 6448
rect 13707 5564 13749 5573
rect 13707 5524 13708 5564
rect 13748 5524 13749 5564
rect 13707 5515 13749 5524
rect 13612 4927 13652 4936
rect 13708 4976 13748 5515
rect 13708 4927 13748 4936
rect 13707 3968 13749 3977
rect 13707 3928 13708 3968
rect 13748 3928 13749 3968
rect 13707 3919 13749 3928
rect 13419 3884 13461 3893
rect 13419 3844 13420 3884
rect 13460 3844 13461 3884
rect 13419 3835 13461 3844
rect 13228 2500 13364 2540
rect 12940 2036 12980 2045
rect 12980 1996 13268 2036
rect 12940 1987 12980 1996
rect 13228 1952 13268 1996
rect 13228 1903 13268 1912
rect 13324 1952 13364 2500
rect 13419 2204 13461 2213
rect 13419 2164 13420 2204
rect 13460 2164 13461 2204
rect 13419 2155 13461 2164
rect 13228 1112 13268 1121
rect 12844 1072 13228 1112
rect 12747 1063 12789 1072
rect 13228 1063 13268 1072
rect 12651 1028 12693 1037
rect 12651 988 12652 1028
rect 12692 988 12693 1028
rect 12651 979 12693 988
rect 12748 80 12788 1063
rect 13324 953 13364 1912
rect 13323 944 13365 953
rect 13323 904 13324 944
rect 13364 904 13365 944
rect 13323 895 13365 904
rect 13420 869 13460 2155
rect 13708 1952 13748 3919
rect 13900 2540 13940 7783
rect 13996 7421 14036 7960
rect 14092 7673 14132 9379
rect 14188 8597 14228 9724
rect 14284 8672 14324 8681
rect 14187 8588 14229 8597
rect 14187 8548 14188 8588
rect 14228 8548 14229 8588
rect 14187 8539 14229 8548
rect 14187 8420 14229 8429
rect 14187 8380 14188 8420
rect 14228 8380 14229 8420
rect 14187 8371 14229 8380
rect 14091 7664 14133 7673
rect 14091 7624 14092 7664
rect 14132 7624 14133 7664
rect 14091 7615 14133 7624
rect 13995 7412 14037 7421
rect 13995 7372 13996 7412
rect 14036 7372 14037 7412
rect 13995 7363 14037 7372
rect 14091 7328 14133 7337
rect 14091 7288 14092 7328
rect 14132 7288 14133 7328
rect 14091 7279 14133 7288
rect 13995 7076 14037 7085
rect 13995 7036 13996 7076
rect 14036 7036 14037 7076
rect 13995 7027 14037 7036
rect 13996 6488 14036 7027
rect 13996 6439 14036 6448
rect 14092 3800 14132 7279
rect 14188 4976 14228 8371
rect 14284 7841 14324 8632
rect 14283 7832 14325 7841
rect 14283 7792 14284 7832
rect 14324 7792 14325 7832
rect 14283 7783 14325 7792
rect 14283 7160 14325 7169
rect 14283 7120 14284 7160
rect 14324 7120 14325 7160
rect 14283 7111 14325 7120
rect 14284 7026 14324 7111
rect 14380 6656 14420 10312
rect 14476 10184 14516 10193
rect 14476 9773 14516 10144
rect 14475 9764 14517 9773
rect 14475 9724 14476 9764
rect 14516 9724 14517 9764
rect 14475 9715 14517 9724
rect 14476 9596 14516 9715
rect 14572 9680 14612 10639
rect 14667 10100 14709 10109
rect 14667 10060 14668 10100
rect 14708 10060 14709 10100
rect 14667 10051 14709 10060
rect 14668 9966 14708 10051
rect 14668 9680 14708 9689
rect 14572 9640 14668 9680
rect 14668 9631 14708 9640
rect 14476 9556 14612 9596
rect 14476 9498 14516 9507
rect 14476 8924 14516 9458
rect 14476 8875 14516 8884
rect 14475 8588 14517 8597
rect 14475 8548 14476 8588
rect 14516 8548 14517 8588
rect 14475 8539 14517 8548
rect 14476 7337 14516 8539
rect 14475 7328 14517 7337
rect 14475 7288 14476 7328
rect 14516 7288 14517 7328
rect 14475 7279 14517 7288
rect 14572 6740 14612 9556
rect 14860 9512 14900 11815
rect 14956 11453 14996 13831
rect 15147 13544 15189 13553
rect 15147 13504 15148 13544
rect 15188 13504 15189 13544
rect 15147 13495 15189 13504
rect 15051 13208 15093 13217
rect 15051 13168 15052 13208
rect 15092 13168 15093 13208
rect 15051 13159 15093 13168
rect 15148 13208 15188 13495
rect 15148 13159 15188 13168
rect 15243 13208 15285 13217
rect 15243 13168 15244 13208
rect 15284 13168 15285 13208
rect 15243 13159 15285 13168
rect 15052 13074 15092 13159
rect 15051 12956 15093 12965
rect 15051 12916 15052 12956
rect 15092 12916 15093 12956
rect 15051 12907 15093 12916
rect 15052 12536 15092 12907
rect 15244 12620 15284 13159
rect 15244 12571 15284 12580
rect 15092 12496 15188 12536
rect 15052 12487 15092 12496
rect 15051 12116 15093 12125
rect 15051 12076 15052 12116
rect 15092 12076 15093 12116
rect 15051 12067 15093 12076
rect 15052 11696 15092 12067
rect 15148 11705 15188 12496
rect 15052 11647 15092 11656
rect 15147 11696 15189 11705
rect 15147 11656 15148 11696
rect 15188 11656 15189 11696
rect 15147 11647 15189 11656
rect 14955 11444 14997 11453
rect 14955 11404 14956 11444
rect 14996 11404 14997 11444
rect 14955 11395 14997 11404
rect 15147 10688 15189 10697
rect 15147 10648 15148 10688
rect 15188 10648 15189 10688
rect 15147 10639 15189 10648
rect 15148 10277 15188 10639
rect 15147 10268 15189 10277
rect 15147 10228 15148 10268
rect 15188 10228 15189 10268
rect 15147 10219 15189 10228
rect 14956 10184 14996 10193
rect 14956 10109 14996 10144
rect 15052 10184 15092 10195
rect 15052 10109 15092 10144
rect 14948 10100 14996 10109
rect 14948 10060 14949 10100
rect 14989 10060 14996 10100
rect 15051 10100 15093 10109
rect 15051 10060 15052 10100
rect 15092 10060 15093 10100
rect 14948 10051 14990 10060
rect 15051 10051 15093 10060
rect 14860 9463 14900 9472
rect 15148 9512 15188 10219
rect 15148 9463 15188 9472
rect 14859 9344 14901 9353
rect 15340 9344 15380 14428
rect 15436 13964 15476 16192
rect 15531 16232 15573 16241
rect 15531 16192 15532 16232
rect 15572 16192 15573 16232
rect 15531 16183 15573 16192
rect 15532 16098 15572 16183
rect 15628 16148 15668 16435
rect 15916 16400 15956 16409
rect 15724 16360 15916 16400
rect 15724 16232 15764 16360
rect 15916 16351 15956 16360
rect 15724 16183 15764 16192
rect 15915 16232 15957 16241
rect 15915 16192 15916 16232
rect 15956 16192 15957 16232
rect 15915 16183 15957 16192
rect 15628 16099 15668 16108
rect 15916 15728 15956 16183
rect 15916 15569 15956 15688
rect 15723 15560 15765 15569
rect 15723 15520 15724 15560
rect 15764 15520 15765 15560
rect 15723 15511 15765 15520
rect 15915 15560 15957 15569
rect 15915 15520 15916 15560
rect 15956 15520 15957 15560
rect 15915 15511 15957 15520
rect 15724 15426 15764 15511
rect 15723 14972 15765 14981
rect 15723 14932 15724 14972
rect 15764 14932 15765 14972
rect 15723 14923 15765 14932
rect 15627 14552 15669 14561
rect 15627 14512 15628 14552
rect 15668 14512 15669 14552
rect 15627 14503 15669 14512
rect 15436 13924 15572 13964
rect 15435 13628 15477 13637
rect 15435 13588 15436 13628
rect 15476 13588 15477 13628
rect 15435 13579 15477 13588
rect 15436 12620 15476 13579
rect 15532 13469 15572 13924
rect 15531 13460 15573 13469
rect 15531 13420 15532 13460
rect 15572 13420 15573 13460
rect 15531 13411 15573 13420
rect 15628 13292 15668 14503
rect 15628 13243 15668 13252
rect 15532 13208 15572 13217
rect 15532 13133 15572 13168
rect 15531 13124 15573 13133
rect 15531 13084 15532 13124
rect 15572 13084 15573 13124
rect 15531 13075 15573 13084
rect 15532 12788 15572 13075
rect 15724 12965 15764 14923
rect 15819 13880 15861 13889
rect 15819 13840 15820 13880
rect 15860 13840 15861 13880
rect 15819 13831 15861 13840
rect 15723 12956 15765 12965
rect 15723 12916 15724 12956
rect 15764 12916 15765 12956
rect 15723 12907 15765 12916
rect 15532 12748 15764 12788
rect 15532 12620 15572 12629
rect 15436 12580 15532 12620
rect 15532 12571 15572 12580
rect 15627 12536 15669 12545
rect 15627 12496 15628 12536
rect 15668 12496 15669 12536
rect 15627 12487 15669 12496
rect 15628 12402 15668 12487
rect 15531 11864 15573 11873
rect 15531 11824 15532 11864
rect 15572 11824 15573 11864
rect 15531 11815 15573 11824
rect 15435 10520 15477 10529
rect 15435 10480 15436 10520
rect 15476 10480 15477 10520
rect 15435 10471 15477 10480
rect 15436 10268 15476 10471
rect 15436 10219 15476 10228
rect 15532 10184 15572 11815
rect 15724 11789 15764 12748
rect 15820 12536 15860 13831
rect 15915 13376 15957 13385
rect 15915 13336 15916 13376
rect 15956 13336 15957 13376
rect 15915 13327 15957 13336
rect 15820 12487 15860 12496
rect 15916 12536 15956 13327
rect 15916 12487 15956 12496
rect 16012 12368 16052 17200
rect 16108 13880 16148 20140
rect 16203 19928 16245 19937
rect 16203 19888 16204 19928
rect 16244 19888 16245 19928
rect 16203 19879 16245 19888
rect 16204 18005 16244 19879
rect 16299 18920 16341 18929
rect 16299 18880 16300 18920
rect 16340 18880 16341 18920
rect 16299 18871 16341 18880
rect 16203 17996 16245 18005
rect 16203 17956 16204 17996
rect 16244 17956 16245 17996
rect 16300 17996 16340 18871
rect 16300 17956 16344 17996
rect 16203 17947 16245 17956
rect 16304 17858 16344 17956
rect 16203 17828 16245 17837
rect 16203 17788 16204 17828
rect 16244 17788 16245 17828
rect 16203 17779 16245 17788
rect 16300 17788 16344 17858
rect 16204 17744 16244 17779
rect 16204 17693 16244 17704
rect 16300 17763 16340 17788
rect 16300 17660 16340 17723
rect 16396 17744 16436 20644
rect 16492 19265 16532 22240
rect 16588 21944 16628 24592
rect 16780 23549 16820 27616
rect 17068 26816 17108 27859
rect 17164 27656 17204 28960
rect 17548 28748 17588 32815
rect 17740 32784 17780 32815
rect 17836 32696 17876 36847
rect 18027 36812 18069 36821
rect 18027 36772 18028 36812
rect 18068 36772 18069 36812
rect 18027 36763 18069 36772
rect 17931 35972 17973 35981
rect 17931 35932 17932 35972
rect 17972 35932 17973 35972
rect 17931 35923 17973 35932
rect 17932 32789 17972 35923
rect 18028 35216 18068 36763
rect 18124 35888 18164 37099
rect 18124 35561 18164 35848
rect 18123 35552 18165 35561
rect 18123 35512 18124 35552
rect 18164 35512 18165 35552
rect 18123 35503 18165 35512
rect 18123 35300 18165 35309
rect 18123 35260 18124 35300
rect 18164 35260 18165 35300
rect 18123 35251 18165 35260
rect 18028 34721 18068 35176
rect 18124 35216 18164 35251
rect 18124 35165 18164 35176
rect 18027 34712 18069 34721
rect 18027 34672 18028 34712
rect 18068 34672 18069 34712
rect 18027 34663 18069 34672
rect 18220 34544 18260 37435
rect 18316 37400 18356 37409
rect 18316 36905 18356 37360
rect 18315 36896 18357 36905
rect 18315 36856 18316 36896
rect 18356 36856 18357 36896
rect 18315 36847 18357 36856
rect 18315 36476 18357 36485
rect 18315 36436 18316 36476
rect 18356 36436 18357 36476
rect 18315 36427 18357 36436
rect 18316 35888 18356 36427
rect 18412 36401 18452 38275
rect 18507 37652 18549 37661
rect 18507 37612 18508 37652
rect 18548 37612 18549 37652
rect 18507 37603 18549 37612
rect 18508 37409 18548 37603
rect 18507 37400 18549 37409
rect 18507 37360 18508 37400
rect 18548 37360 18549 37400
rect 18507 37351 18549 37360
rect 18411 36392 18453 36401
rect 18411 36352 18412 36392
rect 18452 36352 18453 36392
rect 18411 36343 18453 36352
rect 18316 35813 18356 35848
rect 18315 35804 18357 35813
rect 18315 35764 18316 35804
rect 18356 35764 18357 35804
rect 18315 35755 18357 35764
rect 18028 34504 18260 34544
rect 18028 33368 18068 34504
rect 18123 34376 18165 34385
rect 18123 34336 18124 34376
rect 18164 34336 18165 34376
rect 18123 34327 18165 34336
rect 18124 34242 18164 34327
rect 18316 34208 18356 34217
rect 18316 33713 18356 34168
rect 18315 33704 18357 33713
rect 18315 33664 18316 33704
rect 18356 33664 18357 33704
rect 18315 33655 18357 33664
rect 18219 33620 18261 33629
rect 18219 33580 18220 33620
rect 18260 33580 18261 33620
rect 18219 33571 18261 33580
rect 18220 33486 18260 33571
rect 18411 33452 18453 33461
rect 18411 33412 18412 33452
rect 18452 33412 18453 33452
rect 18411 33403 18453 33412
rect 18028 33328 18356 33368
rect 18027 32864 18069 32873
rect 18220 32864 18260 32873
rect 18027 32824 18028 32864
rect 18068 32824 18069 32864
rect 18027 32815 18069 32824
rect 18124 32824 18220 32864
rect 17931 32780 17973 32789
rect 17931 32740 17932 32780
rect 17972 32740 17973 32780
rect 17931 32731 17973 32740
rect 17644 32656 17876 32696
rect 17644 29924 17684 32656
rect 17740 31361 17780 31446
rect 17739 31352 17781 31361
rect 17739 31312 17740 31352
rect 17780 31312 17781 31352
rect 17739 31303 17781 31312
rect 17932 31184 17972 31193
rect 17740 31144 17932 31184
rect 17740 30680 17780 31144
rect 17932 31135 17972 31144
rect 18028 31016 18068 32815
rect 17932 30976 18068 31016
rect 17740 30631 17780 30640
rect 17836 30680 17876 30689
rect 17644 29000 17684 29884
rect 17739 29840 17781 29849
rect 17836 29840 17876 30640
rect 17739 29800 17740 29840
rect 17780 29800 17876 29840
rect 17739 29791 17781 29800
rect 17740 29706 17780 29791
rect 17644 28960 17780 29000
rect 17356 28708 17588 28748
rect 17260 28160 17300 28169
rect 17260 27833 17300 28120
rect 17259 27824 17301 27833
rect 17259 27784 17260 27824
rect 17300 27784 17301 27824
rect 17259 27775 17301 27784
rect 17164 27616 17300 27656
rect 17163 26900 17205 26909
rect 17163 26860 17164 26900
rect 17204 26860 17205 26900
rect 17163 26851 17205 26860
rect 17068 25304 17108 26776
rect 16876 25264 17108 25304
rect 16779 23540 16821 23549
rect 16779 23500 16780 23540
rect 16820 23500 16821 23540
rect 16779 23491 16821 23500
rect 16876 22709 16916 25264
rect 16972 24548 17012 24557
rect 16875 22700 16917 22709
rect 16875 22660 16876 22700
rect 16916 22660 16917 22700
rect 16875 22651 16917 22660
rect 16972 22289 17012 24508
rect 17068 24548 17108 24559
rect 17068 24473 17108 24508
rect 17067 24464 17109 24473
rect 17067 24424 17068 24464
rect 17108 24424 17109 24464
rect 17067 24415 17109 24424
rect 17164 24128 17204 26851
rect 17260 26153 17300 27616
rect 17259 26144 17301 26153
rect 17259 26104 17260 26144
rect 17300 26104 17301 26144
rect 17259 26095 17301 26104
rect 17260 24809 17300 26095
rect 17259 24800 17301 24809
rect 17259 24760 17260 24800
rect 17300 24760 17301 24800
rect 17259 24751 17301 24760
rect 17356 24473 17396 28708
rect 17547 28496 17589 28505
rect 17547 28456 17548 28496
rect 17588 28456 17589 28496
rect 17547 28447 17589 28456
rect 17548 28328 17588 28447
rect 17548 28279 17588 28288
rect 17644 28328 17684 28337
rect 17451 27404 17493 27413
rect 17451 27364 17452 27404
rect 17492 27364 17493 27404
rect 17451 27355 17493 27364
rect 17452 26144 17492 27355
rect 17644 26984 17684 28288
rect 17452 26095 17492 26104
rect 17548 26944 17684 26984
rect 17548 26144 17588 26944
rect 17643 26816 17685 26825
rect 17643 26776 17644 26816
rect 17684 26776 17685 26816
rect 17643 26767 17685 26776
rect 17644 26682 17684 26767
rect 17548 25136 17588 26104
rect 17643 25640 17685 25649
rect 17643 25600 17644 25640
rect 17684 25600 17685 25640
rect 17643 25591 17685 25600
rect 17644 25481 17684 25591
rect 17643 25472 17685 25481
rect 17643 25432 17644 25472
rect 17684 25432 17685 25472
rect 17643 25423 17685 25432
rect 17644 25304 17684 25423
rect 17644 25255 17684 25264
rect 17548 25096 17684 25136
rect 17547 24632 17589 24641
rect 17547 24592 17548 24632
rect 17588 24592 17589 24632
rect 17547 24583 17589 24592
rect 17451 24548 17493 24557
rect 17451 24508 17452 24548
rect 17492 24508 17493 24548
rect 17451 24499 17493 24508
rect 17355 24464 17397 24473
rect 17355 24424 17356 24464
rect 17396 24424 17397 24464
rect 17355 24415 17397 24424
rect 17068 24088 17204 24128
rect 16971 22280 17013 22289
rect 16971 22240 16972 22280
rect 17012 22240 17013 22280
rect 16971 22231 17013 22240
rect 16684 22112 16724 22121
rect 16724 22072 17012 22112
rect 16684 22063 16724 22072
rect 16588 21904 16820 21944
rect 16587 20852 16629 20861
rect 16587 20812 16588 20852
rect 16628 20812 16629 20852
rect 16587 20803 16629 20812
rect 16588 20684 16628 20803
rect 16588 20635 16628 20644
rect 16780 19769 16820 21904
rect 16972 21608 17012 22072
rect 16972 21559 17012 21568
rect 17068 21608 17108 24088
rect 17163 23960 17205 23969
rect 17163 23920 17164 23960
rect 17204 23920 17205 23960
rect 17163 23911 17205 23920
rect 17068 20441 17108 21568
rect 17164 22280 17204 23911
rect 17356 23792 17396 23801
rect 17452 23792 17492 24499
rect 17548 24305 17588 24583
rect 17547 24296 17589 24305
rect 17547 24256 17548 24296
rect 17588 24256 17589 24296
rect 17547 24247 17589 24256
rect 17644 23969 17684 25096
rect 17740 24464 17780 28960
rect 17835 28916 17877 28925
rect 17835 28876 17836 28916
rect 17876 28876 17877 28916
rect 17835 28867 17877 28876
rect 17836 26825 17876 28867
rect 17932 27917 17972 30976
rect 18027 30680 18069 30689
rect 18027 30640 18028 30680
rect 18068 30640 18069 30680
rect 18027 30631 18069 30640
rect 18028 28337 18068 30631
rect 18124 29924 18164 32824
rect 18220 32815 18260 32824
rect 18219 32528 18261 32537
rect 18219 32488 18220 32528
rect 18260 32488 18261 32528
rect 18219 32479 18261 32488
rect 18220 30680 18260 32479
rect 18316 30689 18356 33328
rect 18412 33318 18452 33403
rect 18412 31352 18452 31361
rect 18412 30857 18452 31312
rect 18411 30848 18453 30857
rect 18411 30808 18412 30848
rect 18452 30808 18453 30848
rect 18411 30799 18453 30808
rect 18220 30008 18260 30640
rect 18315 30680 18357 30689
rect 18315 30640 18316 30680
rect 18356 30640 18357 30680
rect 18315 30631 18357 30640
rect 18316 30546 18356 30631
rect 18220 29968 18356 30008
rect 18124 29884 18259 29924
rect 18124 28589 18164 29884
rect 18219 29882 18259 29884
rect 18219 29833 18259 29842
rect 18316 29756 18356 29968
rect 18220 29716 18356 29756
rect 18123 28580 18165 28589
rect 18123 28540 18124 28580
rect 18164 28540 18165 28580
rect 18123 28531 18165 28540
rect 18027 28328 18069 28337
rect 18027 28288 18028 28328
rect 18068 28288 18069 28328
rect 18027 28279 18069 28288
rect 18124 28328 18164 28339
rect 18028 28194 18068 28279
rect 18124 28253 18164 28288
rect 18123 28244 18165 28253
rect 18123 28204 18124 28244
rect 18164 28204 18165 28244
rect 18123 28195 18165 28204
rect 18027 27992 18069 28001
rect 18027 27952 18028 27992
rect 18068 27952 18069 27992
rect 18027 27943 18069 27952
rect 17931 27908 17973 27917
rect 17931 27868 17932 27908
rect 17972 27868 17973 27908
rect 17931 27859 17973 27868
rect 18028 27740 18068 27943
rect 17932 27700 18068 27740
rect 17932 27656 17972 27700
rect 17835 26816 17877 26825
rect 17835 26776 17836 26816
rect 17876 26776 17877 26816
rect 17835 26767 17877 26776
rect 17836 26489 17876 26767
rect 17835 26480 17877 26489
rect 17835 26440 17836 26480
rect 17876 26440 17877 26480
rect 17835 26431 17877 26440
rect 17932 26405 17972 27616
rect 18123 27404 18165 27413
rect 18123 27364 18124 27404
rect 18164 27364 18165 27404
rect 18123 27355 18165 27364
rect 18124 27270 18164 27355
rect 18220 26984 18260 29716
rect 18315 29504 18357 29513
rect 18315 29464 18316 29504
rect 18356 29464 18357 29504
rect 18315 29455 18357 29464
rect 18316 29168 18356 29455
rect 18508 29345 18548 37351
rect 18604 35384 18644 38956
rect 18700 38947 18740 38956
rect 18699 38828 18741 38837
rect 18699 38788 18700 38828
rect 18740 38788 18741 38828
rect 18699 38779 18741 38788
rect 18700 38240 18740 38779
rect 18796 38417 18836 39124
rect 19179 39124 19180 39164
rect 19220 39124 19221 39164
rect 19179 39115 19221 39124
rect 18988 38753 19028 38838
rect 18987 38744 19029 38753
rect 18987 38704 18988 38744
rect 19028 38704 19029 38744
rect 18987 38695 19029 38704
rect 19180 38660 19220 39115
rect 19276 38996 19316 39005
rect 19276 38837 19316 38956
rect 19275 38828 19317 38837
rect 19275 38788 19276 38828
rect 19316 38788 19317 38828
rect 19275 38779 19317 38788
rect 19372 38753 19412 39208
rect 19660 38996 19700 39005
rect 19564 38956 19660 38996
rect 19371 38744 19413 38753
rect 19371 38704 19372 38744
rect 19412 38704 19413 38744
rect 19371 38695 19413 38704
rect 19468 38744 19508 38753
rect 19180 38620 19316 38660
rect 18987 38576 19029 38585
rect 18987 38536 18988 38576
rect 19028 38536 19029 38576
rect 18987 38527 19029 38536
rect 18795 38408 18837 38417
rect 18795 38368 18796 38408
rect 18836 38368 18837 38408
rect 18795 38359 18837 38368
rect 18700 37073 18740 38200
rect 18988 38156 19028 38527
rect 19180 38408 19220 38417
rect 18988 38107 19028 38116
rect 19084 38368 19180 38408
rect 19084 37997 19124 38368
rect 19180 38359 19220 38368
rect 19083 37988 19125 37997
rect 19083 37948 19084 37988
rect 19124 37948 19125 37988
rect 19083 37939 19125 37948
rect 18808 37820 19176 37829
rect 18848 37780 18890 37820
rect 18930 37780 18972 37820
rect 19012 37780 19054 37820
rect 19094 37780 19136 37820
rect 18808 37771 19176 37780
rect 18891 37484 18933 37493
rect 18891 37444 18892 37484
rect 18932 37444 18933 37484
rect 18891 37435 18933 37444
rect 18795 37400 18837 37409
rect 18795 37360 18796 37400
rect 18836 37360 18837 37400
rect 18795 37351 18837 37360
rect 18796 37266 18836 37351
rect 18699 37064 18741 37073
rect 18699 37024 18700 37064
rect 18740 37024 18741 37064
rect 18699 37015 18741 37024
rect 18700 36728 18740 36737
rect 18700 36401 18740 36688
rect 18892 36485 18932 37435
rect 19276 37414 19316 38620
rect 19468 38417 19508 38704
rect 19467 38408 19509 38417
rect 19467 38368 19468 38408
rect 19508 38368 19509 38408
rect 19467 38359 19509 38368
rect 19371 38324 19413 38333
rect 19371 38284 19372 38324
rect 19412 38284 19413 38324
rect 19371 38275 19413 38284
rect 19372 38156 19412 38275
rect 19564 38156 19604 38956
rect 19660 38947 19700 38956
rect 19948 38753 19988 39460
rect 20140 39450 20180 39535
rect 20044 38996 20084 39007
rect 20044 38921 20084 38956
rect 20043 38912 20085 38921
rect 20043 38872 20044 38912
rect 20084 38872 20085 38912
rect 20043 38863 20085 38872
rect 19852 38744 19892 38753
rect 19372 38107 19412 38116
rect 19468 38116 19604 38156
rect 19659 38157 19701 38165
rect 19756 38157 19796 38165
rect 19659 38156 19796 38157
rect 19659 38116 19660 38156
rect 19700 38117 19756 38156
rect 19700 38116 19701 38117
rect 19746 38116 19756 38117
rect 19371 37988 19413 37997
rect 19371 37948 19372 37988
rect 19412 37948 19413 37988
rect 19371 37939 19413 37948
rect 19276 37365 19316 37374
rect 19372 37148 19412 37939
rect 19468 37316 19508 38116
rect 19659 38107 19701 38116
rect 19756 38107 19796 38116
rect 19564 37988 19604 37997
rect 19564 37904 19604 37948
rect 19659 37904 19701 37913
rect 19564 37864 19660 37904
rect 19700 37864 19701 37904
rect 19659 37855 19701 37864
rect 19660 37484 19700 37493
rect 19468 37267 19508 37276
rect 19564 37444 19660 37484
rect 19564 37157 19604 37444
rect 19660 37435 19700 37444
rect 19852 37409 19892 38704
rect 19947 38744 19989 38753
rect 19947 38704 19948 38744
rect 19988 38704 19989 38744
rect 19947 38695 19989 38704
rect 20236 38744 20276 38753
rect 20276 38704 20564 38744
rect 20236 38695 20276 38704
rect 20048 38576 20416 38585
rect 20088 38536 20130 38576
rect 20170 38536 20212 38576
rect 20252 38536 20294 38576
rect 20334 38536 20376 38576
rect 20048 38527 20416 38536
rect 20139 38324 20181 38333
rect 20139 38284 20140 38324
rect 20180 38284 20181 38324
rect 20139 38275 20181 38284
rect 20140 38190 20180 38275
rect 19947 37988 19989 37997
rect 19947 37948 19948 37988
rect 19988 37948 19989 37988
rect 19947 37939 19989 37948
rect 19948 37854 19988 37939
rect 20524 37745 20564 38704
rect 21004 38669 21044 39703
rect 21003 38660 21045 38669
rect 21003 38620 21004 38660
rect 21044 38620 21045 38660
rect 21003 38611 21045 38620
rect 20907 37988 20949 37997
rect 20907 37948 20908 37988
rect 20948 37948 20949 37988
rect 20907 37939 20949 37948
rect 20619 37904 20661 37913
rect 20619 37864 20620 37904
rect 20660 37864 20661 37904
rect 20619 37855 20661 37864
rect 20523 37736 20565 37745
rect 20523 37696 20524 37736
rect 20564 37696 20565 37736
rect 20523 37687 20565 37696
rect 20043 37484 20085 37493
rect 20043 37444 20044 37484
rect 20084 37444 20085 37484
rect 20043 37435 20085 37444
rect 19851 37400 19893 37409
rect 19851 37360 19852 37400
rect 19892 37360 19893 37400
rect 19851 37351 19893 37360
rect 20044 37350 20084 37435
rect 19659 37316 19701 37325
rect 19659 37276 19660 37316
rect 19700 37276 19701 37316
rect 19659 37267 19701 37276
rect 19563 37148 19605 37157
rect 19372 37108 19508 37148
rect 19179 36896 19221 36905
rect 19179 36856 19180 36896
rect 19220 36856 19221 36896
rect 19179 36847 19221 36856
rect 19180 36762 19220 36847
rect 19468 36737 19508 37108
rect 19563 37108 19564 37148
rect 19604 37108 19605 37148
rect 19563 37099 19605 37108
rect 19563 36896 19605 36905
rect 19563 36856 19564 36896
rect 19604 36856 19605 36896
rect 19563 36847 19605 36856
rect 19564 36762 19604 36847
rect 19467 36728 19509 36737
rect 19467 36688 19468 36728
rect 19508 36688 19509 36728
rect 19467 36679 19509 36688
rect 18988 36644 19028 36653
rect 19371 36644 19413 36653
rect 19028 36604 19316 36644
rect 18988 36595 19028 36604
rect 18891 36476 18933 36485
rect 18891 36436 18892 36476
rect 18932 36436 18933 36476
rect 18891 36427 18933 36436
rect 18699 36392 18741 36401
rect 18699 36352 18700 36392
rect 18740 36352 18741 36392
rect 18699 36343 18741 36352
rect 18808 36308 19176 36317
rect 18848 36268 18890 36308
rect 18930 36268 18972 36308
rect 19012 36268 19054 36308
rect 19094 36268 19136 36308
rect 18808 36259 19176 36268
rect 19276 35897 19316 36604
rect 19371 36604 19372 36644
rect 19412 36604 19413 36644
rect 19371 36595 19413 36604
rect 19372 36510 19412 36595
rect 19563 35972 19605 35981
rect 19563 35932 19564 35972
rect 19604 35932 19605 35972
rect 19563 35923 19605 35932
rect 19275 35888 19317 35897
rect 19275 35848 19276 35888
rect 19316 35848 19317 35888
rect 19275 35839 19317 35848
rect 19564 35888 19604 35923
rect 19564 35837 19604 35848
rect 19083 35720 19125 35729
rect 19083 35680 19084 35720
rect 19124 35680 19125 35720
rect 19083 35671 19125 35680
rect 18604 35344 18740 35384
rect 18603 35216 18645 35225
rect 18603 35176 18604 35216
rect 18644 35176 18645 35216
rect 18603 35167 18645 35176
rect 18604 35082 18644 35167
rect 18603 34460 18645 34469
rect 18603 34420 18604 34460
rect 18644 34420 18645 34460
rect 18603 34411 18645 34420
rect 18604 34326 18644 34411
rect 18700 34385 18740 35344
rect 19084 35211 19124 35671
rect 19275 35300 19317 35309
rect 19275 35260 19276 35300
rect 19316 35260 19317 35300
rect 19275 35251 19317 35260
rect 19084 35162 19124 35171
rect 19276 35166 19316 35251
rect 19467 35132 19509 35141
rect 19660 35132 19700 37267
rect 19852 37232 19892 37241
rect 20236 37232 20276 37241
rect 19892 37192 19988 37232
rect 19852 37183 19892 37192
rect 19948 36728 19988 37192
rect 20276 37192 20564 37232
rect 20236 37183 20276 37192
rect 20048 37064 20416 37073
rect 20088 37024 20130 37064
rect 20170 37024 20212 37064
rect 20252 37024 20294 37064
rect 20334 37024 20376 37064
rect 20048 37015 20416 37024
rect 19948 36688 20084 36728
rect 19756 36644 19796 36653
rect 19796 36604 19892 36644
rect 19756 36595 19796 36604
rect 19755 35720 19797 35729
rect 19755 35680 19756 35720
rect 19796 35680 19797 35720
rect 19755 35671 19797 35680
rect 19756 35586 19796 35671
rect 19852 35309 19892 36604
rect 19947 36560 19989 36569
rect 19947 36520 19948 36560
rect 19988 36520 19989 36560
rect 19947 36511 19989 36520
rect 19948 36426 19988 36511
rect 19947 35972 19989 35981
rect 19947 35932 19948 35972
rect 19988 35932 19989 35972
rect 19947 35923 19989 35932
rect 19948 35838 19988 35923
rect 20044 35720 20084 36688
rect 20524 35897 20564 37192
rect 20620 36065 20660 37855
rect 20715 37400 20757 37409
rect 20715 37360 20716 37400
rect 20756 37360 20757 37400
rect 20715 37351 20757 37360
rect 20619 36056 20661 36065
rect 20619 36016 20620 36056
rect 20660 36016 20661 36056
rect 20619 36007 20661 36016
rect 20523 35888 20565 35897
rect 20523 35848 20524 35888
rect 20564 35848 20565 35888
rect 20523 35839 20565 35848
rect 19948 35680 20084 35720
rect 20140 35720 20180 35729
rect 20180 35680 20660 35720
rect 19948 35393 19988 35680
rect 20140 35671 20180 35680
rect 20048 35552 20416 35561
rect 20088 35512 20130 35552
rect 20170 35512 20212 35552
rect 20252 35512 20294 35552
rect 20334 35512 20376 35552
rect 20048 35503 20416 35512
rect 19947 35384 19989 35393
rect 19947 35344 19948 35384
rect 19988 35344 19989 35384
rect 19947 35335 19989 35344
rect 19851 35300 19893 35309
rect 19851 35260 19852 35300
rect 19892 35260 19893 35300
rect 19851 35251 19893 35260
rect 19947 35216 19989 35225
rect 19947 35176 19948 35216
rect 19988 35176 19989 35216
rect 19947 35167 19989 35176
rect 19467 35092 19468 35132
rect 19508 35092 19509 35132
rect 19467 35083 19509 35092
rect 19564 35092 19700 35132
rect 19852 35132 19892 35141
rect 19468 34998 19508 35083
rect 19564 34880 19604 35092
rect 19468 34840 19604 34880
rect 19660 34964 19700 34973
rect 18808 34796 19176 34805
rect 18848 34756 18890 34796
rect 18930 34756 18972 34796
rect 19012 34756 19054 34796
rect 19094 34756 19136 34796
rect 18808 34747 19176 34756
rect 18988 34460 19028 34469
rect 18892 34420 18988 34460
rect 18699 34376 18741 34385
rect 18699 34336 18700 34376
rect 18740 34336 18741 34376
rect 18699 34327 18741 34336
rect 18795 34208 18837 34217
rect 18795 34168 18796 34208
rect 18836 34168 18837 34208
rect 18795 34159 18837 34168
rect 18796 34074 18836 34159
rect 18604 33620 18644 33629
rect 18604 33116 18644 33580
rect 18796 33461 18836 33546
rect 18892 33545 18932 34420
rect 18988 34411 19028 34420
rect 19372 34460 19412 34469
rect 19180 34208 19220 34217
rect 19220 34168 19316 34208
rect 19180 34159 19220 34168
rect 18987 33620 19029 33629
rect 18987 33580 18988 33620
rect 19028 33580 19029 33620
rect 18987 33571 19029 33580
rect 18891 33536 18933 33545
rect 18891 33496 18892 33536
rect 18932 33496 18933 33536
rect 18891 33487 18933 33496
rect 18988 33486 19028 33571
rect 19180 33545 19220 33630
rect 19179 33536 19221 33545
rect 19179 33496 19180 33536
rect 19220 33496 19221 33536
rect 19179 33487 19221 33496
rect 19276 33461 19316 34168
rect 19372 34133 19412 34420
rect 19371 34124 19413 34133
rect 19371 34084 19372 34124
rect 19412 34084 19413 34124
rect 19371 34075 19413 34084
rect 19371 33788 19413 33797
rect 19371 33748 19372 33788
rect 19412 33748 19413 33788
rect 19371 33739 19413 33748
rect 19372 33620 19412 33739
rect 19372 33571 19412 33580
rect 18795 33452 18837 33461
rect 18795 33412 18796 33452
rect 18836 33412 18837 33452
rect 18795 33403 18837 33412
rect 19275 33452 19317 33461
rect 19275 33412 19276 33452
rect 19316 33412 19317 33452
rect 19275 33403 19317 33412
rect 18808 33284 19176 33293
rect 19468 33284 19508 34840
rect 19563 34208 19605 34217
rect 19563 34168 19564 34208
rect 19604 34168 19605 34208
rect 19563 34159 19605 34168
rect 19564 34074 19604 34159
rect 19660 33713 19700 34924
rect 19852 34637 19892 35092
rect 19851 34628 19893 34637
rect 19851 34588 19852 34628
rect 19892 34588 19893 34628
rect 19851 34579 19893 34588
rect 19755 34544 19797 34553
rect 19755 34504 19756 34544
rect 19796 34504 19797 34544
rect 19755 34495 19797 34504
rect 19756 34460 19796 34495
rect 19756 34409 19796 34420
rect 19948 34376 19988 35167
rect 19852 34336 19988 34376
rect 20044 34964 20084 34973
rect 19852 33881 19892 34336
rect 20044 34217 20084 34924
rect 20620 34385 20660 35680
rect 20619 34376 20661 34385
rect 20619 34336 20620 34376
rect 20660 34336 20661 34376
rect 20619 34327 20661 34336
rect 19948 34208 19988 34217
rect 19851 33872 19893 33881
rect 19851 33832 19852 33872
rect 19892 33832 19893 33872
rect 19851 33823 19893 33832
rect 19659 33704 19701 33713
rect 19659 33664 19660 33704
rect 19700 33664 19701 33704
rect 19659 33655 19701 33664
rect 19756 33620 19796 33629
rect 19948 33620 19988 34168
rect 20043 34208 20085 34217
rect 20043 34168 20044 34208
rect 20084 34168 20085 34208
rect 20043 34159 20085 34168
rect 20048 34040 20416 34049
rect 20088 34000 20130 34040
rect 20170 34000 20212 34040
rect 20252 34000 20294 34040
rect 20334 34000 20376 34040
rect 20048 33991 20416 34000
rect 19796 33580 19892 33620
rect 19948 33580 20084 33620
rect 19756 33571 19796 33580
rect 19564 33452 19604 33461
rect 19604 33412 19700 33452
rect 19564 33403 19604 33412
rect 18848 33244 18890 33284
rect 18930 33244 18972 33284
rect 19012 33244 19054 33284
rect 19094 33244 19136 33284
rect 18808 33235 19176 33244
rect 19276 33244 19508 33284
rect 18604 33076 18932 33116
rect 18748 32873 18788 32882
rect 18788 32833 18836 32864
rect 18748 32824 18836 32833
rect 18603 32780 18645 32789
rect 18603 32740 18604 32780
rect 18644 32740 18645 32780
rect 18603 32731 18645 32740
rect 18604 32192 18644 32731
rect 18796 32360 18836 32824
rect 18892 32780 18932 33076
rect 18892 32731 18932 32740
rect 18892 32360 18932 32369
rect 18796 32320 18892 32360
rect 18892 32311 18932 32320
rect 18700 32192 18740 32201
rect 18604 32152 18700 32192
rect 18604 31361 18644 32152
rect 18700 32143 18740 32152
rect 18808 31772 19176 31781
rect 18848 31732 18890 31772
rect 18930 31732 18972 31772
rect 19012 31732 19054 31772
rect 19094 31732 19136 31772
rect 18808 31723 19176 31732
rect 19276 31529 19316 33244
rect 19564 33125 19604 33210
rect 19660 33209 19700 33412
rect 19659 33200 19701 33209
rect 19659 33160 19660 33200
rect 19700 33160 19701 33200
rect 19659 33151 19701 33160
rect 19563 33116 19605 33125
rect 19563 33076 19564 33116
rect 19604 33076 19605 33116
rect 19563 33067 19605 33076
rect 19371 32948 19413 32957
rect 19756 32948 19796 32957
rect 19371 32908 19372 32948
rect 19412 32908 19413 32948
rect 19371 32899 19413 32908
rect 19468 32908 19756 32948
rect 19372 32814 19412 32899
rect 19372 32108 19412 32117
rect 19275 31520 19317 31529
rect 19275 31480 19276 31520
rect 19316 31480 19317 31520
rect 19275 31471 19317 31480
rect 18603 31352 18645 31361
rect 18603 31312 18604 31352
rect 18644 31312 18645 31352
rect 18603 31303 18645 31312
rect 19372 31268 19412 32068
rect 19180 31228 19412 31268
rect 18795 30680 18837 30689
rect 18795 30640 18796 30680
rect 18836 30640 18837 30680
rect 18795 30631 18837 30640
rect 18796 30546 18836 30631
rect 19180 30512 19220 31228
rect 19468 30848 19508 32908
rect 19756 32899 19796 32908
rect 19852 32453 19892 33580
rect 19947 33452 19989 33461
rect 19947 33412 19948 33452
rect 19988 33412 19989 33452
rect 19947 33403 19989 33412
rect 19948 33318 19988 33403
rect 20044 33041 20084 33580
rect 19948 33032 19988 33041
rect 19948 32789 19988 32992
rect 20043 33032 20085 33041
rect 20043 32992 20044 33032
rect 20084 32992 20085 33032
rect 20043 32983 20085 32992
rect 19947 32780 19989 32789
rect 19947 32740 19948 32780
rect 19988 32740 19989 32780
rect 19947 32731 19989 32740
rect 20048 32528 20416 32537
rect 20088 32488 20130 32528
rect 20170 32488 20212 32528
rect 20252 32488 20294 32528
rect 20334 32488 20376 32528
rect 20048 32479 20416 32488
rect 19851 32444 19893 32453
rect 19851 32404 19852 32444
rect 19892 32404 19893 32444
rect 19851 32395 19893 32404
rect 19756 32108 19796 32117
rect 19563 31940 19605 31949
rect 19563 31900 19564 31940
rect 19604 31900 19605 31940
rect 19563 31891 19605 31900
rect 19564 31806 19604 31891
rect 19564 31361 19604 31446
rect 19563 31352 19605 31361
rect 19660 31352 19700 31361
rect 19563 31312 19564 31352
rect 19604 31312 19660 31352
rect 19563 31303 19605 31312
rect 19660 31303 19700 31312
rect 19468 30799 19508 30808
rect 19275 30764 19317 30773
rect 19275 30724 19276 30764
rect 19316 30724 19317 30764
rect 19275 30715 19317 30724
rect 19276 30675 19316 30715
rect 19276 30626 19316 30635
rect 19180 30472 19316 30512
rect 18808 30260 19176 30269
rect 18848 30220 18890 30260
rect 18930 30220 18972 30260
rect 19012 30220 19054 30260
rect 19094 30220 19136 30260
rect 18808 30211 19176 30220
rect 18795 30092 18837 30101
rect 18795 30052 18796 30092
rect 18836 30052 18837 30092
rect 18795 30043 18837 30052
rect 18700 29845 18740 29854
rect 18700 29345 18740 29805
rect 18507 29336 18549 29345
rect 18507 29296 18508 29336
rect 18548 29296 18549 29336
rect 18507 29287 18549 29296
rect 18699 29336 18741 29345
rect 18699 29296 18700 29336
rect 18740 29296 18741 29336
rect 18699 29287 18741 29296
rect 18316 29119 18356 29128
rect 18507 29168 18549 29177
rect 18507 29128 18508 29168
rect 18548 29128 18549 29168
rect 18507 29119 18549 29128
rect 18508 29034 18548 29119
rect 18796 29000 18836 30043
rect 18892 29756 18932 29765
rect 19276 29756 19316 30472
rect 19564 30269 19604 31303
rect 19660 30596 19700 30605
rect 19563 30260 19605 30269
rect 19563 30220 19564 30260
rect 19604 30220 19605 30260
rect 19563 30211 19605 30220
rect 18932 29716 19316 29756
rect 19372 29924 19412 29933
rect 18892 29707 18932 29716
rect 19372 29000 19412 29884
rect 19564 29672 19604 29681
rect 19564 29093 19604 29632
rect 19660 29597 19700 30556
rect 19756 30185 19796 32068
rect 20716 32033 20756 37351
rect 20908 36401 20948 37939
rect 21291 36896 21333 36905
rect 21291 36856 21292 36896
rect 21332 36856 21333 36896
rect 21291 36847 21333 36856
rect 20907 36392 20949 36401
rect 20907 36352 20908 36392
rect 20948 36352 20949 36392
rect 20907 36343 20949 36352
rect 21292 34721 21332 36847
rect 21387 35888 21429 35897
rect 21387 35848 21388 35888
rect 21428 35848 21429 35888
rect 21387 35839 21429 35848
rect 21388 35729 21428 35839
rect 21387 35720 21429 35729
rect 21387 35680 21388 35720
rect 21428 35680 21429 35720
rect 21387 35671 21429 35680
rect 21291 34712 21333 34721
rect 21291 34672 21292 34712
rect 21332 34672 21333 34712
rect 21291 34663 21333 34672
rect 20811 33536 20853 33545
rect 20811 33496 20812 33536
rect 20852 33496 20853 33536
rect 20811 33487 20853 33496
rect 20715 32024 20757 32033
rect 20715 31984 20716 32024
rect 20756 31984 20757 32024
rect 20715 31975 20757 31984
rect 19948 31940 19988 31949
rect 19852 31900 19948 31940
rect 19852 31361 19892 31900
rect 19948 31891 19988 31900
rect 20812 31697 20852 33487
rect 21195 33284 21237 33293
rect 21195 33244 21196 33284
rect 21236 33244 21237 33284
rect 21195 33235 21237 33244
rect 21099 31940 21141 31949
rect 21099 31900 21100 31940
rect 21140 31900 21141 31940
rect 21099 31891 21141 31900
rect 20811 31688 20853 31697
rect 20811 31648 20812 31688
rect 20852 31648 20853 31688
rect 20811 31639 20853 31648
rect 20044 31436 20084 31445
rect 19851 31352 19893 31361
rect 19851 31312 19852 31352
rect 19892 31312 19893 31352
rect 19851 31303 19893 31312
rect 20044 31193 20084 31396
rect 19852 31184 19892 31193
rect 19852 30773 19892 31144
rect 20043 31184 20085 31193
rect 20043 31144 20044 31184
rect 20084 31144 20085 31184
rect 20043 31135 20085 31144
rect 20236 31184 20276 31193
rect 20276 31144 20756 31184
rect 20236 31135 20276 31144
rect 20048 31016 20416 31025
rect 20088 30976 20130 31016
rect 20170 30976 20212 31016
rect 20252 30976 20294 31016
rect 20334 30976 20376 31016
rect 20048 30967 20416 30976
rect 19851 30764 19893 30773
rect 19851 30724 19852 30764
rect 19892 30724 19893 30764
rect 19851 30715 19893 30724
rect 20043 30596 20085 30605
rect 20043 30556 20044 30596
rect 20084 30556 20085 30596
rect 20043 30547 20085 30556
rect 20044 30462 20084 30547
rect 19852 30428 19892 30437
rect 19755 30176 19797 30185
rect 19755 30136 19756 30176
rect 19796 30136 19797 30176
rect 19755 30127 19797 30136
rect 19755 29924 19797 29933
rect 19755 29884 19756 29924
rect 19796 29884 19797 29924
rect 19755 29875 19797 29884
rect 19756 29790 19796 29875
rect 19659 29588 19701 29597
rect 19659 29548 19660 29588
rect 19700 29548 19701 29588
rect 19659 29539 19701 29548
rect 19756 29168 19796 29177
rect 19563 29084 19605 29093
rect 19563 29044 19564 29084
rect 19604 29044 19605 29084
rect 19563 29035 19605 29044
rect 18700 28960 18836 29000
rect 19276 28960 19412 29000
rect 18604 28328 18644 28337
rect 18700 28328 18740 28960
rect 18808 28748 19176 28757
rect 18848 28708 18890 28748
rect 18930 28708 18972 28748
rect 19012 28708 19054 28748
rect 19094 28708 19136 28748
rect 18808 28699 19176 28708
rect 18795 28580 18837 28589
rect 18795 28540 18796 28580
rect 18836 28540 18837 28580
rect 18795 28531 18837 28540
rect 18644 28288 18740 28328
rect 18316 27656 18356 27667
rect 18316 27581 18356 27616
rect 18315 27572 18357 27581
rect 18315 27532 18316 27572
rect 18356 27532 18357 27572
rect 18315 27523 18357 27532
rect 18508 26984 18548 26993
rect 18028 26944 18260 26984
rect 18316 26944 18508 26984
rect 17931 26396 17973 26405
rect 17931 26356 17932 26396
rect 17972 26356 17973 26396
rect 17931 26347 17973 26356
rect 17931 26060 17973 26069
rect 17931 26020 17932 26060
rect 17972 26020 17973 26060
rect 17931 26011 17973 26020
rect 18028 26060 18068 26944
rect 18172 26825 18212 26834
rect 18316 26825 18356 26944
rect 18508 26935 18548 26944
rect 18212 26785 18356 26825
rect 18172 26776 18212 26785
rect 18315 26648 18357 26657
rect 18315 26608 18316 26648
rect 18356 26608 18357 26648
rect 18315 26599 18357 26608
rect 18316 26514 18356 26599
rect 18411 26564 18453 26573
rect 18411 26524 18412 26564
rect 18452 26524 18453 26564
rect 18411 26515 18453 26524
rect 18219 26480 18261 26489
rect 18219 26440 18220 26480
rect 18260 26440 18261 26480
rect 18219 26431 18261 26440
rect 18068 26020 18164 26060
rect 18028 26011 18068 26020
rect 17932 25926 17972 26011
rect 18028 25313 18068 25398
rect 18027 25304 18069 25313
rect 18027 25264 18028 25304
rect 18068 25264 18069 25304
rect 18027 25255 18069 25264
rect 17836 25136 17876 25145
rect 17876 25096 18068 25136
rect 17836 25087 17876 25096
rect 18028 24627 18068 25096
rect 18028 24578 18068 24587
rect 17740 24424 18068 24464
rect 17643 23960 17685 23969
rect 17643 23920 17644 23960
rect 17684 23920 17685 23960
rect 17643 23911 17685 23920
rect 17931 23876 17973 23885
rect 17931 23836 17932 23876
rect 17972 23836 17973 23876
rect 17931 23827 17973 23836
rect 17836 23792 17876 23801
rect 17396 23752 17492 23792
rect 17356 23743 17396 23752
rect 17452 22541 17492 23752
rect 17548 23752 17836 23792
rect 17548 23708 17588 23752
rect 17836 23743 17876 23752
rect 17932 23792 17972 23827
rect 17932 23741 17972 23752
rect 17548 23659 17588 23668
rect 18028 23624 18068 24424
rect 18124 24380 18164 26020
rect 18220 24884 18260 26431
rect 18315 26396 18357 26405
rect 18315 26356 18316 26396
rect 18356 26356 18357 26396
rect 18315 26347 18357 26356
rect 18316 25481 18356 26347
rect 18315 25472 18357 25481
rect 18315 25432 18316 25472
rect 18356 25432 18357 25472
rect 18315 25423 18357 25432
rect 18220 24844 18356 24884
rect 18220 24716 18260 24725
rect 18220 24557 18260 24676
rect 18219 24548 18261 24557
rect 18219 24508 18220 24548
rect 18260 24508 18261 24548
rect 18219 24499 18261 24508
rect 18124 24340 18260 24380
rect 18123 23960 18165 23969
rect 18123 23920 18124 23960
rect 18164 23920 18165 23960
rect 18123 23911 18165 23920
rect 17932 23584 18068 23624
rect 17739 23456 17781 23465
rect 17739 23416 17740 23456
rect 17780 23416 17781 23456
rect 17739 23407 17781 23416
rect 17451 22532 17493 22541
rect 17451 22492 17452 22532
rect 17492 22492 17493 22532
rect 17451 22483 17493 22492
rect 17164 20693 17204 22240
rect 17451 22280 17493 22289
rect 17451 22240 17452 22280
rect 17492 22240 17493 22280
rect 17451 22231 17493 22240
rect 17452 21617 17492 22231
rect 17451 21608 17493 21617
rect 17451 21568 17452 21608
rect 17492 21568 17493 21608
rect 17451 21559 17493 21568
rect 17452 21474 17492 21559
rect 17548 21524 17588 21533
rect 17548 21449 17588 21484
rect 17547 21440 17589 21449
rect 17547 21400 17548 21440
rect 17588 21400 17589 21440
rect 17547 21391 17589 21400
rect 17548 21281 17588 21391
rect 17547 21272 17589 21281
rect 17547 21232 17548 21272
rect 17588 21232 17589 21272
rect 17547 21223 17589 21232
rect 17548 20768 17588 20777
rect 17163 20684 17205 20693
rect 17163 20644 17164 20684
rect 17204 20644 17205 20684
rect 17163 20635 17205 20644
rect 17067 20432 17109 20441
rect 17067 20392 17068 20432
rect 17108 20392 17109 20432
rect 17067 20383 17109 20392
rect 17260 20273 17300 20358
rect 17548 20273 17588 20728
rect 17643 20768 17685 20777
rect 17643 20728 17644 20768
rect 17684 20728 17685 20768
rect 17643 20719 17685 20728
rect 17644 20634 17684 20719
rect 17643 20348 17685 20357
rect 17643 20308 17644 20348
rect 17684 20308 17685 20348
rect 17643 20299 17685 20308
rect 17259 20264 17301 20273
rect 17259 20224 17260 20264
rect 17300 20224 17301 20264
rect 17259 20215 17301 20224
rect 17547 20264 17589 20273
rect 17547 20224 17548 20264
rect 17588 20224 17589 20264
rect 17547 20215 17589 20224
rect 17068 20096 17108 20105
rect 17108 20056 17204 20096
rect 17068 20047 17108 20056
rect 16779 19760 16821 19769
rect 16779 19720 16780 19760
rect 16820 19720 16821 19760
rect 16779 19711 16821 19720
rect 17067 19760 17109 19769
rect 17067 19720 17068 19760
rect 17108 19720 17109 19760
rect 17067 19711 17109 19720
rect 16587 19592 16629 19601
rect 16587 19552 16588 19592
rect 16628 19552 16629 19592
rect 16587 19543 16629 19552
rect 16491 19256 16533 19265
rect 16491 19216 16492 19256
rect 16532 19216 16533 19256
rect 16491 19207 16533 19216
rect 16492 19122 16532 19207
rect 16588 19097 16628 19543
rect 16972 19256 17012 19265
rect 16684 19172 16724 19181
rect 16972 19172 17012 19216
rect 17068 19256 17108 19711
rect 17164 19265 17204 20056
rect 17547 19424 17589 19433
rect 17547 19384 17548 19424
rect 17588 19384 17589 19424
rect 17547 19375 17589 19384
rect 17548 19340 17588 19375
rect 17548 19289 17588 19300
rect 17068 19207 17108 19216
rect 17163 19256 17205 19265
rect 17163 19216 17164 19256
rect 17204 19216 17205 19256
rect 17163 19207 17205 19216
rect 17452 19256 17492 19265
rect 16724 19132 17012 19172
rect 16684 19123 16724 19132
rect 16587 19088 16629 19097
rect 16587 19048 16588 19088
rect 16628 19048 16629 19088
rect 16587 19039 16629 19048
rect 17067 19088 17109 19097
rect 17067 19048 17068 19088
rect 17108 19048 17109 19088
rect 17067 19039 17109 19048
rect 16971 18416 17013 18425
rect 16971 18376 16972 18416
rect 17012 18376 17013 18416
rect 16971 18367 17013 18376
rect 16683 17996 16725 18005
rect 16683 17956 16684 17996
rect 16724 17956 16725 17996
rect 16683 17947 16725 17956
rect 16396 17704 16532 17744
rect 16291 17620 16340 17660
rect 16291 17576 16331 17620
rect 16291 17536 16340 17576
rect 16300 16409 16340 17536
rect 16492 16661 16532 17704
rect 16684 17081 16724 17947
rect 16779 17912 16821 17921
rect 16779 17872 16780 17912
rect 16820 17872 16821 17912
rect 16779 17863 16821 17872
rect 16683 17072 16725 17081
rect 16683 17032 16684 17072
rect 16724 17032 16725 17072
rect 16683 17023 16725 17032
rect 16491 16652 16533 16661
rect 16491 16612 16492 16652
rect 16532 16612 16533 16652
rect 16491 16603 16533 16612
rect 16684 16409 16724 17023
rect 16299 16400 16341 16409
rect 16299 16360 16300 16400
rect 16340 16360 16341 16400
rect 16299 16351 16341 16360
rect 16491 16400 16533 16409
rect 16683 16400 16725 16409
rect 16491 16360 16492 16400
rect 16532 16360 16628 16400
rect 16491 16351 16533 16360
rect 16203 16316 16245 16325
rect 16203 16276 16204 16316
rect 16244 16276 16245 16316
rect 16203 16267 16245 16276
rect 16204 16232 16244 16267
rect 16204 15989 16244 16192
rect 16491 16232 16533 16241
rect 16491 16192 16492 16232
rect 16532 16192 16533 16232
rect 16491 16183 16533 16192
rect 16588 16232 16628 16360
rect 16683 16360 16684 16400
rect 16724 16360 16725 16400
rect 16683 16351 16725 16360
rect 16588 16183 16628 16192
rect 16683 16232 16725 16241
rect 16683 16192 16684 16232
rect 16724 16192 16725 16232
rect 16683 16183 16725 16192
rect 16492 16098 16532 16183
rect 16684 16098 16724 16183
rect 16587 16064 16629 16073
rect 16587 16024 16588 16064
rect 16628 16024 16629 16064
rect 16587 16015 16629 16024
rect 16203 15980 16245 15989
rect 16203 15940 16204 15980
rect 16244 15940 16245 15980
rect 16203 15931 16245 15940
rect 16203 15560 16245 15569
rect 16203 15520 16204 15560
rect 16244 15520 16245 15560
rect 16203 15511 16245 15520
rect 16300 15560 16340 15571
rect 16588 15569 16628 16015
rect 16683 15644 16725 15653
rect 16683 15604 16684 15644
rect 16724 15604 16725 15644
rect 16683 15595 16725 15604
rect 16204 15426 16244 15511
rect 16300 15485 16340 15520
rect 16587 15560 16629 15569
rect 16587 15520 16588 15560
rect 16628 15520 16629 15560
rect 16587 15511 16629 15520
rect 16299 15476 16341 15485
rect 16299 15436 16300 15476
rect 16340 15436 16341 15476
rect 16299 15427 16341 15436
rect 16300 15149 16340 15427
rect 16299 15140 16341 15149
rect 16299 15100 16300 15140
rect 16340 15100 16341 15140
rect 16299 15091 16341 15100
rect 16203 14972 16245 14981
rect 16203 14932 16204 14972
rect 16244 14932 16245 14972
rect 16203 14923 16245 14932
rect 16204 14048 16244 14923
rect 16588 14720 16628 15511
rect 16684 15476 16724 15595
rect 16780 15560 16820 17863
rect 16875 16652 16917 16661
rect 16875 16612 16876 16652
rect 16916 16612 16917 16652
rect 16875 16603 16917 16612
rect 16876 16484 16916 16603
rect 16876 16435 16916 16444
rect 16875 16232 16917 16241
rect 16875 16192 16876 16232
rect 16916 16192 16917 16232
rect 16875 16183 16917 16192
rect 16780 15485 16820 15520
rect 16684 15233 16724 15436
rect 16779 15476 16821 15485
rect 16779 15436 16780 15476
rect 16820 15436 16821 15476
rect 16779 15427 16821 15436
rect 16780 15396 16820 15427
rect 16683 15224 16725 15233
rect 16683 15184 16684 15224
rect 16724 15184 16725 15224
rect 16683 15175 16725 15184
rect 16780 14972 16820 14981
rect 16876 14972 16916 16183
rect 16820 14932 16916 14972
rect 16780 14923 16820 14932
rect 16588 14671 16628 14680
rect 16972 14561 17012 18367
rect 17068 16904 17108 19039
rect 17164 18584 17204 19207
rect 17452 18929 17492 19216
rect 17451 18920 17493 18929
rect 17451 18880 17452 18920
rect 17492 18880 17493 18920
rect 17451 18871 17493 18880
rect 17451 18668 17493 18677
rect 17451 18628 17452 18668
rect 17492 18628 17493 18668
rect 17451 18619 17493 18628
rect 17260 18584 17300 18593
rect 17164 18544 17260 18584
rect 17164 17753 17204 18544
rect 17260 18535 17300 18544
rect 17452 18534 17492 18619
rect 17259 18332 17301 18341
rect 17259 18292 17260 18332
rect 17300 18292 17301 18332
rect 17259 18283 17301 18292
rect 17163 17744 17205 17753
rect 17163 17704 17164 17744
rect 17204 17704 17205 17744
rect 17163 17695 17205 17704
rect 17260 17744 17300 18283
rect 17260 17695 17300 17704
rect 17644 17333 17684 20299
rect 17740 20105 17780 23407
rect 17739 20096 17781 20105
rect 17739 20056 17740 20096
rect 17780 20056 17781 20096
rect 17739 20047 17781 20056
rect 17740 19013 17780 20047
rect 17739 19004 17781 19013
rect 17739 18964 17740 19004
rect 17780 18964 17781 19004
rect 17739 18955 17781 18964
rect 17739 18668 17781 18677
rect 17739 18628 17740 18668
rect 17780 18628 17781 18668
rect 17739 18619 17781 18628
rect 17740 18584 17780 18619
rect 17740 18533 17780 18544
rect 17835 18584 17877 18593
rect 17835 18544 17836 18584
rect 17876 18544 17877 18584
rect 17835 18535 17877 18544
rect 17836 18450 17876 18535
rect 17643 17324 17685 17333
rect 17643 17284 17644 17324
rect 17684 17284 17685 17324
rect 17643 17275 17685 17284
rect 17164 17081 17204 17166
rect 17548 17156 17588 17165
rect 17260 17116 17548 17156
rect 17163 17072 17205 17081
rect 17163 17032 17164 17072
rect 17204 17032 17205 17072
rect 17163 17023 17205 17032
rect 17068 16864 17204 16904
rect 17067 16400 17109 16409
rect 17067 16360 17068 16400
rect 17108 16360 17109 16400
rect 17067 16351 17109 16360
rect 17068 16266 17108 16351
rect 16683 14552 16725 14561
rect 16683 14512 16684 14552
rect 16724 14512 16725 14552
rect 16683 14503 16725 14512
rect 16971 14552 17013 14561
rect 16971 14512 16972 14552
rect 17012 14512 17013 14552
rect 16971 14503 17013 14512
rect 16684 14069 16724 14503
rect 16204 13999 16244 14008
rect 16588 14048 16628 14057
rect 16684 14020 16724 14029
rect 16780 14048 16820 14057
rect 16396 13880 16436 13889
rect 16108 13840 16244 13880
rect 16107 13460 16149 13469
rect 16107 13420 16108 13460
rect 16148 13420 16149 13460
rect 16107 13411 16149 13420
rect 16108 13208 16148 13411
rect 16108 13159 16148 13168
rect 16108 12536 16148 12547
rect 16108 12461 16148 12496
rect 16107 12452 16149 12461
rect 16107 12412 16108 12452
rect 16148 12412 16149 12452
rect 16107 12403 16149 12412
rect 15916 12328 16052 12368
rect 15819 12200 15861 12209
rect 15819 12160 15820 12200
rect 15860 12160 15861 12200
rect 15819 12151 15861 12160
rect 15723 11780 15765 11789
rect 15723 11740 15724 11780
rect 15764 11740 15765 11780
rect 15723 11731 15765 11740
rect 15723 11276 15765 11285
rect 15723 11236 15724 11276
rect 15764 11236 15765 11276
rect 15723 11227 15765 11236
rect 15724 10613 15764 11227
rect 15723 10604 15765 10613
rect 15723 10564 15724 10604
rect 15764 10564 15765 10604
rect 15723 10555 15765 10564
rect 15724 10277 15764 10555
rect 15723 10268 15765 10277
rect 15723 10228 15724 10268
rect 15764 10228 15765 10268
rect 15723 10219 15765 10228
rect 15532 9941 15572 10144
rect 15531 9932 15573 9941
rect 15531 9892 15532 9932
rect 15572 9892 15573 9932
rect 15531 9883 15573 9892
rect 15723 9848 15765 9857
rect 15723 9808 15724 9848
rect 15764 9808 15765 9848
rect 15723 9799 15765 9808
rect 14859 9304 14860 9344
rect 14900 9304 14901 9344
rect 14859 9295 14901 9304
rect 15148 9304 15380 9344
rect 14763 8672 14805 8681
rect 14763 8632 14764 8672
rect 14804 8632 14805 8672
rect 14763 8623 14805 8632
rect 14764 8538 14804 8623
rect 14572 6700 14804 6740
rect 14188 4927 14228 4936
rect 14284 6616 14420 6656
rect 14284 3884 14324 6616
rect 14668 6572 14708 6581
rect 14380 6532 14668 6572
rect 14380 3968 14420 6532
rect 14668 6523 14708 6532
rect 14524 6446 14564 6455
rect 14524 6404 14564 6406
rect 14524 6364 14708 6404
rect 14668 5900 14708 6364
rect 14668 5851 14708 5860
rect 14476 5648 14516 5657
rect 14764 5648 14804 6700
rect 14516 5608 14804 5648
rect 14476 5599 14516 5608
rect 14572 5069 14612 5608
rect 14860 5480 14900 9295
rect 14955 9260 14997 9269
rect 14955 9220 14956 9260
rect 14996 9220 14997 9260
rect 14955 9211 14997 9220
rect 14956 9126 14996 9211
rect 14955 9008 14997 9017
rect 14955 8968 14956 9008
rect 14996 8968 14997 9008
rect 14955 8959 14997 8968
rect 14956 8840 14996 8959
rect 14956 8791 14996 8800
rect 14955 8672 14997 8681
rect 14955 8632 14956 8672
rect 14996 8632 14997 8672
rect 14955 8623 14997 8632
rect 15052 8672 15092 8681
rect 14956 8538 14996 8623
rect 15052 8513 15092 8632
rect 15148 8597 15188 9304
rect 15627 9260 15669 9269
rect 15627 9220 15628 9260
rect 15668 9220 15669 9260
rect 15627 9211 15669 9220
rect 15339 9008 15381 9017
rect 15339 8968 15340 9008
rect 15380 8968 15381 9008
rect 15339 8959 15381 8968
rect 15340 8840 15380 8959
rect 15244 8800 15380 8840
rect 15244 8672 15284 8800
rect 15244 8623 15284 8632
rect 15339 8672 15381 8681
rect 15339 8632 15340 8672
rect 15380 8632 15381 8672
rect 15339 8623 15381 8632
rect 15532 8672 15572 8681
rect 15147 8588 15189 8597
rect 15147 8548 15148 8588
rect 15188 8548 15189 8588
rect 15147 8539 15189 8548
rect 15051 8504 15093 8513
rect 15051 8464 15052 8504
rect 15092 8464 15093 8504
rect 15051 8455 15093 8464
rect 15148 8168 15188 8539
rect 15052 8128 15188 8168
rect 15340 8168 15380 8623
rect 15436 8504 15476 8515
rect 15436 8429 15476 8464
rect 15435 8420 15477 8429
rect 15435 8380 15436 8420
rect 15476 8380 15477 8420
rect 15435 8371 15477 8380
rect 15532 8177 15572 8632
rect 15628 8672 15668 9211
rect 15724 8840 15764 9799
rect 15820 9680 15860 12151
rect 15916 9857 15956 12328
rect 16108 12284 16148 12293
rect 16011 12200 16053 12209
rect 16011 12160 16012 12200
rect 16052 12160 16053 12200
rect 16011 12151 16053 12160
rect 16012 10697 16052 12151
rect 16011 10688 16053 10697
rect 16011 10648 16012 10688
rect 16052 10648 16053 10688
rect 16011 10639 16053 10648
rect 16011 10268 16053 10277
rect 16011 10228 16012 10268
rect 16052 10228 16053 10268
rect 16011 10219 16053 10228
rect 16012 10184 16052 10219
rect 16012 10133 16052 10144
rect 16011 9932 16053 9941
rect 16011 9892 16012 9932
rect 16052 9892 16053 9932
rect 16011 9883 16053 9892
rect 15915 9848 15957 9857
rect 15915 9808 15916 9848
rect 15956 9808 15957 9848
rect 15915 9799 15957 9808
rect 15820 9640 15956 9680
rect 15724 8800 15860 8840
rect 15628 8623 15668 8632
rect 15729 8672 15769 8681
rect 15729 8513 15769 8632
rect 15728 8504 15770 8513
rect 15724 8464 15729 8504
rect 15769 8464 15770 8504
rect 15724 8455 15770 8464
rect 15052 7832 15092 8128
rect 15340 8119 15380 8128
rect 15531 8168 15573 8177
rect 15531 8128 15532 8168
rect 15572 8128 15573 8168
rect 15531 8119 15573 8128
rect 15148 8000 15188 8009
rect 15531 8000 15573 8009
rect 15188 7960 15380 8000
rect 15148 7951 15188 7960
rect 15052 7792 15188 7832
rect 15148 6245 15188 7792
rect 15340 6824 15380 7960
rect 15531 7960 15532 8000
rect 15572 7960 15573 8000
rect 15531 7951 15573 7960
rect 15532 7866 15572 7951
rect 15724 7673 15764 8455
rect 15723 7664 15765 7673
rect 15723 7624 15724 7664
rect 15764 7624 15765 7664
rect 15723 7615 15765 7624
rect 15724 7412 15764 7615
rect 15724 7363 15764 7372
rect 15532 7160 15572 7169
rect 15532 6824 15572 7120
rect 15340 6784 15572 6824
rect 15147 6236 15189 6245
rect 15147 6196 15148 6236
rect 15188 6196 15189 6236
rect 15147 6187 15189 6196
rect 15147 6068 15189 6077
rect 15147 6028 15148 6068
rect 15188 6028 15189 6068
rect 15147 6019 15189 6028
rect 14955 5732 14997 5741
rect 14955 5692 14956 5732
rect 14996 5692 14997 5732
rect 14955 5683 14997 5692
rect 14956 5648 14996 5683
rect 14956 5597 14996 5608
rect 15052 5648 15092 5657
rect 14860 5440 14996 5480
rect 14571 5060 14613 5069
rect 14571 5020 14572 5060
rect 14612 5020 14613 5060
rect 14571 5011 14613 5020
rect 14860 5060 14900 5069
rect 14572 4136 14612 5011
rect 14668 4962 14708 4971
rect 14668 4556 14708 4922
rect 14668 4516 14804 4556
rect 14667 4388 14709 4397
rect 14667 4348 14668 4388
rect 14708 4348 14709 4388
rect 14667 4339 14709 4348
rect 14764 4388 14804 4516
rect 14764 4339 14804 4348
rect 14572 4087 14612 4096
rect 14380 3928 14612 3968
rect 14284 3844 14516 3884
rect 14092 3760 14324 3800
rect 14187 3464 14229 3473
rect 14187 3424 14188 3464
rect 14228 3424 14229 3464
rect 14187 3415 14229 3424
rect 14188 3330 14228 3415
rect 13996 2708 14036 2717
rect 14187 2708 14229 2717
rect 14036 2668 14132 2708
rect 13996 2659 14036 2668
rect 13900 2500 14036 2540
rect 13804 2456 13844 2465
rect 13804 2213 13844 2416
rect 13803 2204 13845 2213
rect 13803 2164 13804 2204
rect 13844 2164 13845 2204
rect 13803 2155 13845 2164
rect 13708 1903 13748 1912
rect 13804 1877 13844 1962
rect 13803 1868 13845 1877
rect 13803 1828 13804 1868
rect 13844 1828 13845 1868
rect 13803 1819 13845 1828
rect 13996 1373 14036 2500
rect 14092 2213 14132 2668
rect 14187 2668 14188 2708
rect 14228 2668 14229 2708
rect 14187 2659 14229 2668
rect 14188 2574 14228 2659
rect 14091 2204 14133 2213
rect 14091 2164 14092 2204
rect 14132 2164 14133 2204
rect 14091 2155 14133 2164
rect 14284 1952 14324 3760
rect 14380 2456 14420 2465
rect 14380 1961 14420 2416
rect 14284 1903 14324 1912
rect 14379 1952 14421 1961
rect 14379 1912 14380 1952
rect 14420 1912 14421 1952
rect 14379 1903 14421 1912
rect 14187 1784 14229 1793
rect 14187 1744 14188 1784
rect 14228 1744 14229 1784
rect 14187 1735 14229 1744
rect 13995 1364 14037 1373
rect 13995 1324 13996 1364
rect 14036 1324 14037 1364
rect 13995 1315 14037 1324
rect 14188 1112 14228 1735
rect 14476 1280 14516 3844
rect 14572 1541 14612 3928
rect 14668 2624 14708 4339
rect 14860 2633 14900 5020
rect 14956 4733 14996 5440
rect 15052 5144 15092 5608
rect 15148 5648 15188 6019
rect 15148 5599 15188 5608
rect 15244 5648 15284 5657
rect 15244 5321 15284 5608
rect 15243 5312 15285 5321
rect 15243 5272 15244 5312
rect 15284 5272 15285 5312
rect 15243 5263 15285 5272
rect 15052 5104 15188 5144
rect 15051 4976 15093 4985
rect 15051 4936 15052 4976
rect 15092 4936 15093 4976
rect 15051 4927 15093 4936
rect 15052 4842 15092 4927
rect 14955 4724 14997 4733
rect 14955 4684 14956 4724
rect 14996 4684 14997 4724
rect 14955 4675 14997 4684
rect 15148 4145 15188 5104
rect 15147 4136 15189 4145
rect 15147 4096 15148 4136
rect 15188 4096 15189 4136
rect 15147 4087 15189 4096
rect 15340 3725 15380 6784
rect 15820 6749 15860 8800
rect 15916 8009 15956 9640
rect 15915 8000 15957 8009
rect 15915 7960 15916 8000
rect 15956 7960 15957 8000
rect 15915 7951 15957 7960
rect 15915 7664 15957 7673
rect 15915 7624 15916 7664
rect 15956 7624 15957 7664
rect 15915 7615 15957 7624
rect 15916 7160 15956 7615
rect 15916 7111 15956 7120
rect 16012 7160 16052 9883
rect 16012 7111 16052 7120
rect 15819 6740 15861 6749
rect 15819 6700 15820 6740
rect 15860 6700 15861 6740
rect 15819 6691 15861 6700
rect 15916 6497 15956 6582
rect 15724 6488 15764 6497
rect 15915 6488 15957 6497
rect 15764 6448 15860 6488
rect 15724 6439 15764 6448
rect 15627 6320 15669 6329
rect 15627 6280 15628 6320
rect 15668 6280 15669 6320
rect 15820 6320 15860 6448
rect 15915 6448 15916 6488
rect 15956 6448 15957 6488
rect 15915 6439 15957 6448
rect 16012 6488 16052 6497
rect 15820 6280 15956 6320
rect 15627 6271 15669 6280
rect 15435 6236 15477 6245
rect 15435 6196 15436 6236
rect 15476 6196 15477 6236
rect 15435 6187 15477 6196
rect 15436 5648 15476 6187
rect 15628 6068 15668 6271
rect 15724 6236 15764 6245
rect 15764 6196 15860 6236
rect 15724 6187 15764 6196
rect 15628 6028 15764 6068
rect 15628 5825 15668 5910
rect 15627 5816 15669 5825
rect 15627 5776 15628 5816
rect 15668 5776 15669 5816
rect 15627 5767 15669 5776
rect 15532 5732 15572 5741
rect 15532 5648 15572 5692
rect 15724 5732 15764 6028
rect 15724 5683 15764 5692
rect 15627 5648 15669 5657
rect 15532 5608 15628 5648
rect 15668 5608 15669 5648
rect 15436 5599 15476 5608
rect 15627 5599 15669 5608
rect 15820 5648 15860 6196
rect 15820 5599 15860 5608
rect 15627 5312 15669 5321
rect 15627 5272 15628 5312
rect 15668 5272 15669 5312
rect 15627 5263 15669 5272
rect 15531 5228 15573 5237
rect 15531 5188 15532 5228
rect 15572 5188 15573 5228
rect 15531 5179 15573 5188
rect 15435 4976 15477 4985
rect 15435 4936 15436 4976
rect 15476 4936 15477 4976
rect 15435 4927 15477 4936
rect 15436 3809 15476 4927
rect 15435 3800 15477 3809
rect 15435 3760 15436 3800
rect 15476 3760 15477 3800
rect 15435 3751 15477 3760
rect 15339 3716 15381 3725
rect 15339 3676 15340 3716
rect 15380 3676 15381 3716
rect 15339 3667 15381 3676
rect 15340 2801 15380 3667
rect 15436 3464 15476 3751
rect 15436 3415 15476 3424
rect 15435 3212 15477 3221
rect 15435 3172 15436 3212
rect 15476 3172 15477 3212
rect 15435 3163 15477 3172
rect 15339 2792 15381 2801
rect 15339 2752 15340 2792
rect 15380 2752 15381 2792
rect 15339 2743 15381 2752
rect 14764 2624 14804 2633
rect 14668 2584 14764 2624
rect 14764 2575 14804 2584
rect 14859 2624 14901 2633
rect 14859 2584 14860 2624
rect 14900 2584 14901 2624
rect 14859 2575 14901 2584
rect 14859 2456 14901 2465
rect 14859 2416 14860 2456
rect 14900 2416 14901 2456
rect 14859 2407 14901 2416
rect 14764 1938 14804 1947
rect 14571 1532 14613 1541
rect 14571 1492 14572 1532
rect 14612 1492 14613 1532
rect 14571 1483 14613 1492
rect 14668 1364 14708 1373
rect 14764 1364 14804 1898
rect 14860 1625 14900 2407
rect 15243 2372 15285 2381
rect 15243 2332 15244 2372
rect 15284 2332 15285 2372
rect 15243 2323 15285 2332
rect 14955 2204 14997 2213
rect 14955 2164 14956 2204
rect 14996 2164 14997 2204
rect 14955 2155 14997 2164
rect 14956 2120 14996 2155
rect 14956 2069 14996 2080
rect 14955 1952 14997 1961
rect 14955 1912 14956 1952
rect 14996 1912 14997 1952
rect 14955 1903 14997 1912
rect 15244 1952 15284 2323
rect 15244 1903 15284 1912
rect 14859 1616 14901 1625
rect 14859 1576 14860 1616
rect 14900 1576 14901 1616
rect 14859 1567 14901 1576
rect 14708 1324 14804 1364
rect 14668 1315 14708 1324
rect 14476 1240 14612 1280
rect 14572 1196 14612 1240
rect 14859 1196 14901 1205
rect 14572 1156 14708 1196
rect 14476 1112 14516 1121
rect 14188 1072 14476 1112
rect 14476 1063 14516 1072
rect 13515 1028 13557 1037
rect 13515 988 13516 1028
rect 13556 988 13557 1028
rect 13515 979 13557 988
rect 13419 860 13461 869
rect 13419 820 13420 860
rect 13460 820 13461 860
rect 13419 811 13461 820
rect 13323 608 13365 617
rect 13323 568 13324 608
rect 13364 568 13365 608
rect 13323 559 13365 568
rect 13131 524 13173 533
rect 13131 484 13132 524
rect 13172 484 13173 524
rect 13131 475 13173 484
rect 12939 440 12981 449
rect 12939 400 12940 440
rect 12980 400 12981 440
rect 12939 391 12981 400
rect 12940 80 12980 391
rect 13132 80 13172 475
rect 13324 80 13364 559
rect 13516 80 13556 979
rect 14283 860 14325 869
rect 14283 820 14284 860
rect 14324 820 14325 860
rect 14283 811 14325 820
rect 14475 860 14517 869
rect 14475 820 14476 860
rect 14516 820 14517 860
rect 14475 811 14517 820
rect 13707 776 13749 785
rect 13707 736 13708 776
rect 13748 736 13749 776
rect 13707 727 13749 736
rect 13708 80 13748 727
rect 14091 356 14133 365
rect 14091 316 14092 356
rect 14132 316 14133 356
rect 14091 307 14133 316
rect 13899 272 13941 281
rect 13899 232 13900 272
rect 13940 232 13941 272
rect 13899 223 13941 232
rect 13900 80 13940 223
rect 14092 80 14132 307
rect 14284 80 14324 811
rect 14476 80 14516 811
rect 14668 80 14708 1156
rect 14859 1156 14860 1196
rect 14900 1156 14901 1196
rect 14859 1147 14901 1156
rect 14860 1062 14900 1147
rect 14859 944 14901 953
rect 14859 904 14860 944
rect 14900 904 14901 944
rect 14859 895 14901 904
rect 14860 80 14900 895
rect 14956 776 14996 1903
rect 15052 944 15092 953
rect 15339 944 15381 953
rect 15092 904 15284 944
rect 15052 895 15092 904
rect 14956 736 15092 776
rect 15052 80 15092 736
rect 15244 80 15284 904
rect 15339 904 15340 944
rect 15380 904 15381 944
rect 15339 895 15381 904
rect 15340 810 15380 895
rect 15436 80 15476 3163
rect 15532 2540 15572 5179
rect 15628 3632 15668 5263
rect 15916 4397 15956 6280
rect 16012 6068 16052 6448
rect 16009 6028 16052 6068
rect 16009 5825 16049 6028
rect 16009 5816 16052 5825
rect 16009 5776 16012 5816
rect 16012 5767 16052 5776
rect 15915 4388 15957 4397
rect 15915 4348 15916 4388
rect 15956 4348 15957 4388
rect 15915 4339 15957 4348
rect 15915 4136 15957 4145
rect 15915 4096 15916 4136
rect 15956 4096 15957 4136
rect 15915 4087 15957 4096
rect 15723 3800 15765 3809
rect 15723 3760 15724 3800
rect 15764 3760 15765 3800
rect 15723 3751 15765 3760
rect 15628 3583 15668 3592
rect 15724 2633 15764 3751
rect 15819 3212 15861 3221
rect 15819 3172 15820 3212
rect 15860 3172 15861 3212
rect 15819 3163 15861 3172
rect 15820 3078 15860 3163
rect 15916 2876 15956 4087
rect 16012 3380 16052 3389
rect 16108 3380 16148 12244
rect 16204 11528 16244 13840
rect 16436 13840 16532 13880
rect 16396 13831 16436 13840
rect 16492 13133 16532 13840
rect 16588 13301 16628 14008
rect 16683 13964 16725 13973
rect 16683 13924 16684 13964
rect 16724 13924 16725 13964
rect 16683 13915 16725 13924
rect 16587 13292 16629 13301
rect 16587 13252 16588 13292
rect 16628 13252 16629 13292
rect 16587 13243 16629 13252
rect 16588 13213 16628 13243
rect 16491 13124 16533 13133
rect 16491 13084 16492 13124
rect 16532 13084 16533 13124
rect 16491 13075 16533 13084
rect 16396 12536 16436 12545
rect 16588 12536 16628 13173
rect 16436 12496 16628 12536
rect 16684 12536 16724 13915
rect 16780 13217 16820 14008
rect 16876 14048 16916 14057
rect 17068 14048 17108 14057
rect 16779 13208 16821 13217
rect 16779 13168 16780 13208
rect 16820 13168 16821 13208
rect 16876 13208 16916 14008
rect 16972 14008 17068 14048
rect 16972 13637 17012 14008
rect 17068 13999 17108 14008
rect 17164 13973 17204 16864
rect 17260 16148 17300 17116
rect 17548 17107 17588 17116
rect 17740 17072 17780 17081
rect 17644 17030 17684 17039
rect 17644 16988 17684 16990
rect 17548 16948 17684 16988
rect 17356 16820 17396 16829
rect 17356 16325 17396 16780
rect 17548 16661 17588 16948
rect 17547 16652 17589 16661
rect 17547 16612 17548 16652
rect 17588 16612 17589 16652
rect 17547 16603 17589 16612
rect 17740 16493 17780 17032
rect 17836 17072 17876 17081
rect 17739 16484 17781 16493
rect 17739 16444 17740 16484
rect 17780 16444 17781 16484
rect 17739 16435 17781 16444
rect 17355 16316 17397 16325
rect 17355 16276 17356 16316
rect 17396 16276 17397 16316
rect 17355 16267 17397 16276
rect 17739 16316 17781 16325
rect 17739 16276 17740 16316
rect 17780 16276 17781 16316
rect 17739 16267 17781 16276
rect 17452 16232 17492 16241
rect 17356 16148 17396 16157
rect 17260 16108 17356 16148
rect 17356 16099 17396 16108
rect 17452 15737 17492 16192
rect 17740 16232 17780 16267
rect 17836 16241 17876 17032
rect 17740 16181 17780 16192
rect 17835 16232 17877 16241
rect 17835 16192 17836 16232
rect 17876 16192 17877 16232
rect 17835 16183 17877 16192
rect 17451 15728 17493 15737
rect 17451 15688 17452 15728
rect 17492 15688 17493 15728
rect 17451 15679 17493 15688
rect 17259 15560 17301 15569
rect 17836 15560 17876 16183
rect 17932 15896 17972 23584
rect 18028 21608 18068 21617
rect 18124 21608 18164 23911
rect 18068 21568 18164 21608
rect 18028 20945 18068 21568
rect 18123 21020 18165 21029
rect 18123 20980 18124 21020
rect 18164 20980 18165 21020
rect 18123 20971 18165 20980
rect 18027 20936 18069 20945
rect 18027 20896 18028 20936
rect 18068 20896 18069 20936
rect 18027 20887 18069 20896
rect 18124 20852 18164 20971
rect 18124 20803 18164 20812
rect 18027 20768 18069 20777
rect 18027 20728 18028 20768
rect 18068 20728 18069 20768
rect 18027 20719 18069 20728
rect 18028 20357 18068 20719
rect 18220 20600 18260 24340
rect 18316 23969 18356 24844
rect 18412 24641 18452 26515
rect 18507 26144 18549 26153
rect 18507 26104 18508 26144
rect 18548 26104 18549 26144
rect 18507 26095 18549 26104
rect 18508 24893 18548 26095
rect 18507 24884 18549 24893
rect 18507 24844 18508 24884
rect 18548 24844 18549 24884
rect 18507 24835 18549 24844
rect 18604 24716 18644 28288
rect 18796 27404 18836 28531
rect 19276 28496 19316 28960
rect 19756 28496 19796 29128
rect 19852 28589 19892 30388
rect 20235 30428 20277 30437
rect 20235 30388 20236 30428
rect 20276 30388 20277 30428
rect 20235 30379 20277 30388
rect 20236 30294 20276 30379
rect 19947 29672 19989 29681
rect 19947 29632 19948 29672
rect 19988 29632 19989 29672
rect 19947 29623 19989 29632
rect 19948 29538 19988 29623
rect 20048 29504 20416 29513
rect 20088 29464 20130 29504
rect 20170 29464 20212 29504
rect 20252 29464 20294 29504
rect 20334 29464 20376 29504
rect 20048 29455 20416 29464
rect 19947 29336 19989 29345
rect 19947 29296 19948 29336
rect 19988 29296 19989 29336
rect 19947 29287 19989 29296
rect 19948 29202 19988 29287
rect 20716 29000 20756 31144
rect 20811 29672 20853 29681
rect 20811 29632 20812 29672
rect 20852 29632 20853 29672
rect 20811 29623 20853 29632
rect 20620 28960 20756 29000
rect 19851 28580 19893 28589
rect 19851 28540 19852 28580
rect 19892 28540 19893 28580
rect 19851 28531 19893 28540
rect 18988 28456 19316 28496
rect 19564 28456 19796 28496
rect 18988 27665 19028 28456
rect 19468 28412 19508 28421
rect 19132 28337 19172 28346
rect 19172 28297 19220 28328
rect 19132 28288 19220 28297
rect 19180 27917 19220 28288
rect 19275 28160 19317 28169
rect 19275 28120 19276 28160
rect 19316 28120 19317 28160
rect 19275 28111 19317 28120
rect 19276 28026 19316 28111
rect 19179 27908 19221 27917
rect 19179 27868 19180 27908
rect 19220 27868 19221 27908
rect 19179 27859 19221 27868
rect 19468 27749 19508 28372
rect 19467 27740 19509 27749
rect 19467 27700 19468 27740
rect 19508 27700 19509 27740
rect 19467 27691 19509 27700
rect 18987 27656 19029 27665
rect 18987 27616 18988 27656
rect 19028 27616 19029 27656
rect 18987 27607 19029 27616
rect 19564 27656 19604 28456
rect 19852 28412 19892 28421
rect 19756 28372 19852 28412
rect 19659 28160 19701 28169
rect 19659 28120 19660 28160
rect 19700 28120 19701 28160
rect 19659 28111 19701 28120
rect 19660 28026 19700 28111
rect 19756 28085 19796 28372
rect 19852 28363 19892 28372
rect 20044 28160 20084 28169
rect 19852 28120 20044 28160
rect 19755 28076 19797 28085
rect 19755 28036 19756 28076
rect 19796 28036 19797 28076
rect 19755 28027 19797 28036
rect 19755 27908 19797 27917
rect 19755 27868 19756 27908
rect 19796 27868 19797 27908
rect 19755 27859 19797 27868
rect 19756 27824 19796 27859
rect 19756 27773 19796 27784
rect 19659 27740 19701 27749
rect 19659 27700 19660 27740
rect 19700 27700 19701 27740
rect 19659 27691 19701 27700
rect 18700 27364 18836 27404
rect 18700 26984 18740 27364
rect 18808 27236 19176 27245
rect 18848 27196 18890 27236
rect 18930 27196 18972 27236
rect 19012 27196 19054 27236
rect 19094 27196 19136 27236
rect 18808 27187 19176 27196
rect 18700 26944 18836 26984
rect 18700 26816 18740 26825
rect 18700 26405 18740 26776
rect 18699 26396 18741 26405
rect 18699 26356 18700 26396
rect 18740 26356 18741 26396
rect 18699 26347 18741 26356
rect 18796 26153 18836 26944
rect 19564 26405 19604 27616
rect 19563 26396 19605 26405
rect 19563 26356 19564 26396
rect 19604 26356 19605 26396
rect 19563 26347 19605 26356
rect 19180 26228 19220 26237
rect 18892 26188 19180 26228
rect 18795 26144 18837 26153
rect 18795 26104 18796 26144
rect 18836 26104 18837 26144
rect 18795 26095 18837 26104
rect 18892 25892 18932 26188
rect 19180 26179 19220 26188
rect 19036 26102 19076 26111
rect 19036 26060 19076 26062
rect 19372 26060 19412 26069
rect 19036 26020 19316 26060
rect 18508 24676 18644 24716
rect 18700 25852 18932 25892
rect 18411 24632 18453 24641
rect 18411 24592 18412 24632
rect 18452 24592 18453 24632
rect 18411 24583 18453 24592
rect 18315 23960 18357 23969
rect 18315 23920 18316 23960
rect 18356 23920 18357 23960
rect 18315 23911 18357 23920
rect 18412 23876 18452 24583
rect 18315 23792 18357 23801
rect 18315 23752 18316 23792
rect 18356 23752 18357 23792
rect 18315 23743 18357 23752
rect 18316 23658 18356 23743
rect 18316 23129 18356 23214
rect 18315 23120 18357 23129
rect 18315 23080 18316 23120
rect 18356 23080 18357 23120
rect 18315 23071 18357 23080
rect 18412 22700 18452 23836
rect 18508 23801 18548 24676
rect 18604 24548 18644 24557
rect 18700 24548 18740 25852
rect 18808 25724 19176 25733
rect 18848 25684 18890 25724
rect 18930 25684 18972 25724
rect 19012 25684 19054 25724
rect 19094 25684 19136 25724
rect 18808 25675 19176 25684
rect 19276 25556 19316 26020
rect 19372 25733 19412 26020
rect 19564 25892 19604 25901
rect 19371 25724 19413 25733
rect 19371 25684 19372 25724
rect 19412 25684 19413 25724
rect 19371 25675 19413 25684
rect 19468 25556 19508 25565
rect 19276 25516 19468 25556
rect 19468 25507 19508 25516
rect 19179 25472 19221 25481
rect 19179 25432 19180 25472
rect 19220 25432 19316 25472
rect 19179 25423 19221 25432
rect 19276 25304 19316 25432
rect 19276 25255 19316 25264
rect 18795 25220 18837 25229
rect 18795 25180 18796 25220
rect 18836 25180 18837 25220
rect 18795 25171 18837 25180
rect 18796 24800 18836 25171
rect 19371 25136 19413 25145
rect 19371 25096 19372 25136
rect 19412 25096 19413 25136
rect 19371 25087 19413 25096
rect 18796 24751 18836 24760
rect 18795 24632 18837 24641
rect 18795 24592 18796 24632
rect 18836 24592 18837 24632
rect 18795 24583 18837 24592
rect 18644 24508 18740 24548
rect 18604 24499 18644 24508
rect 18796 24380 18836 24583
rect 18987 24548 19029 24557
rect 18987 24508 18988 24548
rect 19028 24508 19029 24548
rect 18987 24499 19029 24508
rect 19372 24548 19412 25087
rect 19564 25061 19604 25852
rect 19660 25556 19700 27691
rect 19852 26321 19892 28120
rect 20044 28111 20084 28120
rect 20048 27992 20416 28001
rect 20088 27952 20130 27992
rect 20170 27952 20212 27992
rect 20252 27952 20294 27992
rect 20334 27952 20376 27992
rect 20048 27943 20416 27952
rect 19948 27572 19988 27581
rect 19988 27532 20084 27572
rect 19948 27523 19988 27532
rect 19948 26816 19988 26827
rect 19948 26741 19988 26776
rect 19947 26732 19989 26741
rect 19947 26692 19948 26732
rect 19988 26692 19989 26732
rect 19947 26683 19989 26692
rect 20044 26657 20084 27532
rect 20140 27404 20180 27413
rect 20180 27364 20564 27404
rect 20140 27355 20180 27364
rect 20043 26648 20085 26657
rect 20043 26608 20044 26648
rect 20084 26608 20085 26648
rect 20043 26599 20085 26608
rect 20048 26480 20416 26489
rect 20088 26440 20130 26480
rect 20170 26440 20212 26480
rect 20252 26440 20294 26480
rect 20334 26440 20376 26480
rect 20048 26431 20416 26440
rect 19851 26312 19893 26321
rect 19851 26272 19852 26312
rect 19892 26272 19893 26312
rect 19851 26263 19893 26272
rect 19755 26228 19797 26237
rect 19755 26188 19756 26228
rect 19796 26188 19797 26228
rect 19755 26179 19797 26188
rect 19756 26060 19796 26179
rect 19756 26011 19796 26020
rect 19948 25892 19988 25901
rect 19660 25516 19796 25556
rect 19659 25388 19701 25397
rect 19659 25348 19660 25388
rect 19700 25348 19701 25388
rect 19659 25339 19701 25348
rect 19660 25254 19700 25339
rect 19563 25052 19605 25061
rect 19563 25012 19564 25052
rect 19604 25012 19605 25052
rect 19563 25003 19605 25012
rect 19756 24800 19796 25516
rect 19851 25472 19893 25481
rect 19851 25432 19852 25472
rect 19892 25432 19893 25472
rect 19851 25423 19893 25432
rect 19852 25338 19892 25423
rect 19851 24968 19893 24977
rect 19851 24928 19852 24968
rect 19892 24928 19893 24968
rect 19851 24919 19893 24928
rect 19372 24499 19412 24508
rect 19468 24760 19796 24800
rect 18988 24414 19028 24499
rect 19180 24389 19220 24474
rect 18700 24340 18836 24380
rect 19179 24380 19221 24389
rect 19179 24340 19180 24380
rect 19220 24340 19221 24380
rect 18507 23792 18549 23801
rect 18507 23752 18508 23792
rect 18548 23752 18549 23792
rect 18507 23743 18549 23752
rect 18124 20560 18260 20600
rect 18316 22660 18452 22700
rect 18027 20348 18069 20357
rect 18027 20308 18028 20348
rect 18068 20308 18069 20348
rect 18027 20299 18069 20308
rect 18027 19256 18069 19265
rect 18027 19216 18028 19256
rect 18068 19216 18069 19256
rect 18027 19207 18069 19216
rect 18028 19122 18068 19207
rect 18027 17576 18069 17585
rect 18027 17536 18028 17576
rect 18068 17536 18069 17576
rect 18027 17527 18069 17536
rect 18028 16988 18068 17527
rect 18028 16939 18068 16948
rect 17932 15856 18068 15896
rect 17931 15728 17973 15737
rect 17931 15688 17932 15728
rect 17972 15688 17973 15728
rect 17931 15679 17973 15688
rect 17932 15594 17972 15679
rect 17259 15520 17260 15560
rect 17300 15520 17301 15560
rect 17259 15511 17301 15520
rect 17788 15550 17876 15560
rect 17260 15426 17300 15511
rect 17828 15520 17876 15550
rect 17788 15501 17828 15510
rect 17835 15056 17877 15065
rect 17835 15016 17836 15056
rect 17876 15016 17877 15056
rect 17835 15007 17877 15016
rect 17644 14720 17684 14729
rect 17644 14141 17684 14680
rect 17739 14468 17781 14477
rect 17739 14428 17740 14468
rect 17780 14428 17781 14468
rect 17739 14419 17781 14428
rect 17643 14132 17685 14141
rect 17643 14092 17644 14132
rect 17684 14092 17685 14132
rect 17643 14083 17685 14092
rect 17259 14048 17301 14057
rect 17259 14008 17260 14048
rect 17300 14008 17301 14048
rect 17259 13999 17301 14008
rect 17356 14048 17396 14057
rect 17396 14008 17492 14048
rect 17356 13999 17396 14008
rect 17163 13964 17205 13973
rect 17163 13924 17164 13964
rect 17204 13924 17205 13964
rect 17163 13915 17205 13924
rect 17260 13914 17300 13999
rect 17067 13880 17109 13889
rect 17067 13840 17068 13880
rect 17108 13840 17109 13880
rect 17067 13831 17109 13840
rect 17068 13746 17108 13831
rect 16971 13628 17013 13637
rect 16971 13588 16972 13628
rect 17012 13588 17013 13628
rect 16971 13579 17013 13588
rect 16972 13385 17012 13470
rect 16971 13376 17013 13385
rect 16971 13336 16972 13376
rect 17012 13336 17013 13376
rect 16971 13327 17013 13336
rect 17356 13301 17396 13346
rect 17355 13292 17397 13301
rect 17355 13252 17356 13292
rect 17396 13252 17397 13292
rect 17355 13251 17397 13252
rect 17355 13243 17356 13251
rect 17260 13208 17300 13217
rect 16876 13168 17260 13208
rect 17396 13243 17397 13251
rect 17356 13202 17396 13211
rect 16779 13159 16821 13168
rect 17260 13159 17300 13168
rect 17452 13124 17492 14008
rect 16780 13082 16820 13091
rect 16780 13040 16820 13042
rect 17356 13084 17492 13124
rect 16780 13000 17300 13040
rect 17067 12872 17109 12881
rect 17067 12832 17068 12872
rect 17108 12832 17109 12872
rect 17067 12823 17109 12832
rect 16396 12487 16436 12496
rect 16492 11948 16532 12496
rect 16684 12487 16724 12496
rect 16780 12536 16820 12545
rect 16780 12041 16820 12496
rect 17068 12368 17108 12823
rect 17260 12536 17300 13000
rect 17356 12881 17396 13084
rect 17452 12982 17492 12991
rect 17355 12872 17397 12881
rect 17355 12832 17356 12872
rect 17396 12832 17397 12872
rect 17452 12872 17492 12942
rect 17452 12832 17588 12872
rect 17355 12823 17397 12832
rect 17548 12620 17588 12832
rect 17644 12620 17684 12629
rect 17548 12580 17644 12620
rect 17644 12571 17684 12580
rect 17260 12487 17300 12496
rect 17451 12536 17493 12545
rect 17451 12496 17452 12536
rect 17492 12496 17493 12536
rect 17451 12487 17493 12496
rect 17740 12536 17780 14419
rect 17836 13208 17876 15007
rect 17836 13159 17876 13168
rect 17835 13040 17877 13049
rect 17835 13000 17836 13040
rect 17876 13000 17877 13040
rect 17835 12991 17877 13000
rect 17355 12452 17397 12461
rect 17355 12412 17356 12452
rect 17396 12412 17397 12452
rect 17355 12403 17397 12412
rect 17068 12319 17108 12328
rect 17356 12318 17396 12403
rect 17452 12402 17492 12487
rect 16779 12032 16821 12041
rect 16779 11992 16780 12032
rect 16820 11992 16821 12032
rect 16779 11983 16821 11992
rect 16492 11899 16532 11908
rect 16875 11948 16917 11957
rect 16875 11908 16876 11948
rect 16916 11908 16917 11948
rect 16875 11899 16917 11908
rect 16300 11705 16340 11790
rect 16299 11696 16341 11705
rect 16299 11656 16300 11696
rect 16340 11656 16341 11696
rect 16299 11647 16341 11656
rect 16779 11696 16821 11705
rect 16779 11656 16780 11696
rect 16820 11656 16821 11696
rect 16779 11647 16821 11656
rect 16876 11696 16916 11899
rect 16876 11647 16916 11656
rect 16204 11488 16340 11528
rect 16204 8672 16244 8681
rect 16204 8345 16244 8632
rect 16203 8336 16245 8345
rect 16203 8296 16204 8336
rect 16244 8296 16245 8336
rect 16203 8287 16245 8296
rect 16203 8168 16245 8177
rect 16203 8128 16204 8168
rect 16244 8128 16245 8168
rect 16203 8119 16245 8128
rect 16204 6992 16244 8119
rect 16300 7673 16340 11488
rect 16683 10688 16725 10697
rect 16683 10648 16684 10688
rect 16724 10648 16725 10688
rect 16683 10639 16725 10648
rect 16540 10193 16580 10202
rect 16580 10153 16628 10184
rect 16540 10144 16628 10153
rect 16491 9932 16533 9941
rect 16491 9892 16492 9932
rect 16532 9892 16533 9932
rect 16491 9883 16533 9892
rect 16395 9764 16437 9773
rect 16395 9724 16396 9764
rect 16436 9724 16437 9764
rect 16395 9715 16437 9724
rect 16396 9512 16436 9715
rect 16396 9463 16436 9472
rect 16492 8840 16532 9883
rect 16588 9680 16628 10144
rect 16684 10100 16724 10639
rect 16684 10051 16724 10060
rect 16588 9631 16628 9640
rect 16396 8800 16532 8840
rect 16299 7664 16341 7673
rect 16299 7624 16300 7664
rect 16340 7624 16341 7664
rect 16299 7615 16341 7624
rect 16396 7160 16436 8800
rect 16780 8000 16820 11647
rect 17740 11621 17780 12496
rect 17739 11612 17781 11621
rect 17739 11572 17740 11612
rect 17780 11572 17781 11612
rect 17739 11563 17781 11572
rect 16875 11528 16917 11537
rect 16875 11488 16876 11528
rect 16916 11488 16917 11528
rect 16875 11479 16917 11488
rect 16683 7580 16725 7589
rect 16683 7540 16684 7580
rect 16724 7540 16725 7580
rect 16683 7531 16725 7540
rect 16396 7085 16436 7120
rect 16684 7160 16724 7531
rect 16780 7328 16820 7960
rect 16876 7841 16916 11479
rect 17836 11444 17876 12991
rect 17932 12536 17972 12545
rect 17932 12209 17972 12496
rect 18028 12536 18068 15856
rect 18124 13049 18164 20560
rect 18219 20096 18261 20105
rect 18219 20056 18220 20096
rect 18260 20056 18261 20096
rect 18219 20047 18261 20056
rect 18220 19962 18260 20047
rect 18316 18929 18356 22660
rect 18411 22532 18453 22541
rect 18411 22492 18412 22532
rect 18452 22492 18453 22532
rect 18411 22483 18453 22492
rect 18412 22280 18452 22483
rect 18412 22231 18452 22240
rect 18604 22112 18644 22121
rect 18604 21608 18644 22072
rect 18700 21860 18740 24340
rect 19179 24331 19221 24340
rect 18808 24212 19176 24221
rect 18848 24172 18890 24212
rect 18930 24172 18972 24212
rect 19012 24172 19054 24212
rect 19094 24172 19136 24212
rect 18808 24163 19176 24172
rect 19468 23960 19508 24760
rect 19852 24716 19892 24919
rect 19756 24676 19892 24716
rect 19756 24545 19796 24676
rect 19948 24548 19988 25852
rect 20524 25649 20564 27364
rect 20620 27329 20660 28960
rect 20812 28328 20852 29623
rect 20907 29084 20949 29093
rect 20907 29044 20908 29084
rect 20948 29044 20949 29084
rect 20907 29035 20949 29044
rect 20908 28412 20948 29035
rect 20908 28372 21044 28412
rect 20812 28288 20948 28328
rect 20715 28160 20757 28169
rect 20715 28120 20716 28160
rect 20756 28120 20757 28160
rect 20715 28111 20757 28120
rect 20619 27320 20661 27329
rect 20619 27280 20620 27320
rect 20660 27280 20661 27320
rect 20619 27271 20661 27280
rect 20716 25985 20756 28111
rect 20811 27824 20853 27833
rect 20811 27784 20812 27824
rect 20852 27784 20853 27824
rect 20811 27775 20853 27784
rect 20812 26657 20852 27775
rect 20908 27665 20948 28288
rect 20907 27656 20949 27665
rect 20907 27616 20908 27656
rect 20948 27616 20949 27656
rect 20907 27607 20949 27616
rect 21004 26993 21044 28372
rect 21100 28001 21140 31891
rect 21196 29681 21236 33235
rect 21291 30428 21333 30437
rect 21291 30388 21292 30428
rect 21332 30388 21333 30428
rect 21291 30379 21333 30388
rect 21195 29672 21237 29681
rect 21195 29632 21196 29672
rect 21236 29632 21237 29672
rect 21195 29623 21237 29632
rect 21195 28580 21237 28589
rect 21195 28540 21196 28580
rect 21236 28540 21237 28580
rect 21195 28531 21237 28540
rect 21099 27992 21141 28001
rect 21099 27952 21100 27992
rect 21140 27952 21141 27992
rect 21099 27943 21141 27952
rect 21003 26984 21045 26993
rect 21003 26944 21004 26984
rect 21044 26944 21045 26984
rect 21003 26935 21045 26944
rect 20811 26648 20853 26657
rect 21196 26648 21236 28531
rect 20811 26608 20812 26648
rect 20852 26608 20853 26648
rect 20811 26599 20853 26608
rect 21004 26608 21236 26648
rect 20715 25976 20757 25985
rect 20715 25936 20716 25976
rect 20756 25936 20757 25976
rect 20715 25927 20757 25936
rect 20523 25640 20565 25649
rect 20523 25600 20524 25640
rect 20564 25600 20565 25640
rect 20523 25591 20565 25600
rect 20811 25472 20853 25481
rect 20811 25432 20812 25472
rect 20852 25432 20853 25472
rect 20811 25423 20853 25432
rect 20044 25388 20084 25397
rect 20044 25145 20084 25348
rect 20043 25136 20085 25145
rect 20043 25096 20044 25136
rect 20084 25096 20085 25136
rect 20043 25087 20085 25096
rect 20236 25136 20276 25145
rect 20276 25096 20564 25136
rect 20236 25087 20276 25096
rect 20048 24968 20416 24977
rect 20088 24928 20130 24968
rect 20170 24928 20212 24968
rect 20252 24928 20294 24968
rect 20334 24928 20376 24968
rect 20048 24919 20416 24928
rect 20524 24641 20564 25096
rect 20523 24632 20565 24641
rect 20523 24592 20524 24632
rect 20564 24592 20565 24632
rect 20523 24583 20565 24592
rect 19948 24508 20084 24548
rect 19756 24496 19796 24505
rect 19564 24380 19604 24389
rect 19948 24380 19988 24389
rect 19604 24340 19892 24380
rect 19564 24331 19604 24340
rect 19276 23920 19508 23960
rect 18891 23792 18933 23801
rect 18891 23752 18892 23792
rect 18932 23752 18933 23792
rect 18891 23743 18933 23752
rect 18892 23658 18932 23743
rect 19276 23456 19316 23920
rect 19420 23801 19460 23810
rect 19460 23761 19796 23792
rect 19420 23752 19796 23761
rect 19564 23624 19604 23633
rect 19276 23416 19508 23456
rect 19275 23288 19317 23297
rect 19275 23248 19276 23288
rect 19316 23248 19317 23288
rect 19275 23239 19317 23248
rect 18808 22700 19176 22709
rect 18848 22660 18890 22700
rect 18930 22660 18972 22700
rect 19012 22660 19054 22700
rect 19094 22660 19136 22700
rect 18808 22651 19176 22660
rect 18988 22364 19028 22373
rect 19276 22364 19316 23239
rect 19028 22324 19316 22364
rect 19372 22364 19412 22373
rect 18988 22315 19028 22324
rect 19372 22205 19412 22324
rect 19371 22196 19413 22205
rect 19371 22156 19372 22196
rect 19412 22156 19413 22196
rect 19371 22147 19413 22156
rect 19180 22112 19220 22121
rect 19084 22072 19180 22112
rect 18700 21820 18836 21860
rect 18699 21692 18741 21701
rect 18699 21652 18700 21692
rect 18740 21652 18741 21692
rect 18699 21643 18741 21652
rect 18556 21598 18644 21608
rect 18596 21568 18644 21598
rect 18700 21558 18740 21643
rect 18556 21549 18596 21558
rect 18796 21449 18836 21820
rect 18987 21776 19029 21785
rect 18987 21736 18988 21776
rect 19028 21736 19029 21776
rect 18987 21727 19029 21736
rect 18988 21524 19028 21727
rect 18988 21475 19028 21484
rect 18507 21440 18549 21449
rect 18507 21400 18508 21440
rect 18548 21400 18549 21440
rect 18507 21391 18549 21400
rect 18795 21440 18837 21449
rect 18795 21400 18796 21440
rect 18836 21400 18837 21440
rect 18795 21391 18837 21400
rect 18411 20936 18453 20945
rect 18411 20896 18412 20936
rect 18452 20896 18453 20936
rect 18411 20887 18453 20896
rect 18315 18920 18357 18929
rect 18220 18880 18316 18920
rect 18356 18880 18357 18920
rect 18220 18584 18260 18880
rect 18315 18871 18357 18880
rect 18220 17837 18260 18544
rect 18315 18500 18357 18509
rect 18315 18460 18316 18500
rect 18356 18460 18357 18500
rect 18315 18451 18357 18460
rect 18316 18366 18356 18451
rect 18315 18164 18357 18173
rect 18315 18124 18316 18164
rect 18356 18124 18357 18164
rect 18315 18115 18357 18124
rect 18219 17828 18261 17837
rect 18219 17788 18220 17828
rect 18260 17788 18261 17828
rect 18219 17779 18261 17788
rect 18316 17165 18356 18115
rect 18412 17240 18452 20887
rect 18508 20777 18548 21391
rect 19084 21365 19124 22072
rect 19180 22063 19220 22072
rect 19468 21860 19508 23416
rect 19564 23297 19604 23584
rect 19659 23624 19701 23633
rect 19659 23584 19660 23624
rect 19700 23584 19701 23624
rect 19659 23575 19701 23584
rect 19563 23288 19605 23297
rect 19563 23248 19564 23288
rect 19604 23248 19605 23288
rect 19563 23239 19605 23248
rect 19564 23120 19604 23129
rect 19564 22541 19604 23080
rect 19563 22532 19605 22541
rect 19563 22492 19564 22532
rect 19604 22492 19605 22532
rect 19563 22483 19605 22492
rect 19660 22457 19700 23575
rect 19756 23288 19796 23752
rect 19756 23239 19796 23248
rect 19852 22961 19892 24340
rect 19948 23633 19988 24340
rect 20044 23717 20084 24508
rect 20043 23708 20085 23717
rect 20043 23668 20044 23708
rect 20084 23668 20085 23708
rect 20043 23659 20085 23668
rect 19947 23624 19989 23633
rect 19947 23584 19948 23624
rect 19988 23584 19989 23624
rect 19947 23575 19989 23584
rect 20048 23456 20416 23465
rect 20088 23416 20130 23456
rect 20170 23416 20212 23456
rect 20252 23416 20294 23456
rect 20334 23416 20376 23456
rect 20048 23407 20416 23416
rect 20043 23288 20085 23297
rect 20043 23248 20044 23288
rect 20084 23248 20085 23288
rect 20043 23239 20085 23248
rect 19947 23036 19989 23045
rect 19947 22996 19948 23036
rect 19988 22996 19989 23036
rect 19947 22987 19989 22996
rect 19851 22952 19893 22961
rect 19851 22912 19852 22952
rect 19892 22912 19893 22952
rect 19851 22903 19893 22912
rect 19948 22902 19988 22987
rect 19755 22616 19797 22625
rect 19755 22576 19756 22616
rect 19796 22576 19797 22616
rect 19755 22567 19797 22576
rect 19659 22448 19701 22457
rect 19659 22408 19660 22448
rect 19700 22408 19701 22448
rect 19659 22399 19701 22408
rect 19756 22364 19796 22567
rect 19948 22532 19988 22541
rect 20044 22532 20084 23239
rect 20140 22868 20180 22877
rect 20140 22541 20180 22828
rect 19988 22492 20084 22532
rect 20139 22532 20181 22541
rect 20139 22492 20140 22532
rect 20180 22492 20181 22532
rect 19948 22483 19988 22492
rect 20139 22483 20181 22492
rect 19756 22315 19796 22324
rect 19563 22112 19605 22121
rect 19563 22072 19564 22112
rect 19604 22072 19605 22112
rect 19563 22063 19605 22072
rect 19564 21978 19604 22063
rect 20048 21944 20416 21953
rect 20088 21904 20130 21944
rect 20170 21904 20212 21944
rect 20252 21904 20294 21944
rect 20334 21904 20376 21944
rect 20048 21895 20416 21904
rect 19468 21820 19796 21860
rect 19467 21692 19509 21701
rect 19467 21652 19468 21692
rect 19508 21652 19509 21692
rect 19467 21643 19509 21652
rect 19371 21524 19413 21533
rect 19371 21484 19372 21524
rect 19412 21484 19413 21524
rect 19371 21475 19413 21484
rect 19372 21390 19412 21475
rect 19083 21356 19125 21365
rect 19083 21316 19084 21356
rect 19124 21316 19125 21356
rect 19083 21307 19125 21316
rect 19180 21356 19220 21365
rect 19220 21316 19316 21356
rect 19180 21307 19220 21316
rect 18808 21188 19176 21197
rect 18848 21148 18890 21188
rect 18930 21148 18972 21188
rect 19012 21148 19054 21188
rect 19094 21148 19136 21188
rect 18808 21139 19176 21148
rect 19276 20945 19316 21316
rect 18603 20936 18645 20945
rect 18603 20896 18604 20936
rect 18644 20896 18645 20936
rect 18603 20887 18645 20896
rect 19275 20936 19317 20945
rect 19275 20896 19276 20936
rect 19316 20896 19317 20936
rect 19275 20887 19317 20896
rect 18507 20768 18549 20777
rect 18507 20728 18508 20768
rect 18548 20728 18549 20768
rect 18507 20719 18549 20728
rect 18604 20768 18644 20887
rect 19468 20852 19508 21643
rect 19563 21440 19605 21449
rect 19563 21400 19564 21440
rect 19604 21400 19605 21440
rect 19563 21391 19605 21400
rect 19564 21306 19604 21391
rect 19468 20803 19508 20812
rect 19132 20777 19172 20786
rect 19172 20737 19412 20768
rect 19132 20728 19412 20737
rect 18604 20719 18644 20728
rect 19275 20600 19317 20609
rect 19275 20560 19276 20600
rect 19316 20560 19317 20600
rect 19275 20551 19317 20560
rect 19276 20466 19316 20551
rect 19372 20348 19412 20728
rect 19660 20600 19700 20609
rect 19660 20357 19700 20560
rect 19659 20348 19701 20357
rect 19372 20308 19604 20348
rect 19564 20180 19604 20308
rect 19659 20308 19660 20348
rect 19700 20308 19701 20348
rect 19659 20299 19701 20308
rect 19660 20180 19700 20189
rect 19564 20140 19660 20180
rect 19660 20131 19700 20140
rect 19467 20096 19509 20105
rect 19467 20056 19468 20096
rect 19508 20056 19509 20096
rect 19467 20047 19509 20056
rect 19468 19962 19508 20047
rect 18808 19676 19176 19685
rect 18848 19636 18890 19676
rect 18930 19636 18972 19676
rect 19012 19636 19054 19676
rect 19094 19636 19136 19676
rect 18808 19627 19176 19636
rect 19563 19592 19605 19601
rect 19563 19552 19564 19592
rect 19604 19552 19605 19592
rect 19563 19543 19605 19552
rect 18987 19508 19029 19517
rect 18987 19468 18988 19508
rect 19028 19468 19029 19508
rect 18987 19459 19029 19468
rect 19564 19508 19604 19543
rect 19756 19508 19796 21820
rect 19851 20852 19893 20861
rect 19851 20812 19852 20852
rect 19892 20812 19893 20852
rect 19851 20803 19893 20812
rect 19852 20718 19892 20803
rect 20812 20609 20852 25423
rect 20907 22532 20949 22541
rect 20907 22492 20908 22532
rect 20948 22492 20949 22532
rect 20907 22483 20949 22492
rect 20908 21617 20948 22483
rect 20907 21608 20949 21617
rect 20907 21568 20908 21608
rect 20948 21568 20949 21608
rect 20907 21559 20949 21568
rect 19851 20600 19893 20609
rect 20044 20600 20084 20609
rect 19851 20560 19852 20600
rect 19892 20560 19893 20600
rect 19851 20551 19893 20560
rect 19948 20560 20044 20600
rect 19852 20012 19892 20551
rect 19852 19963 19892 19972
rect 18988 19340 19028 19459
rect 19564 19457 19604 19468
rect 19660 19468 19796 19508
rect 18988 19291 19028 19300
rect 19371 19340 19413 19349
rect 19371 19300 19372 19340
rect 19412 19300 19413 19340
rect 19371 19291 19413 19300
rect 18556 19265 18596 19274
rect 18596 19256 18634 19265
rect 18795 19256 18837 19265
rect 18596 19225 18644 19256
rect 18556 19216 18644 19225
rect 18604 17996 18644 19216
rect 18795 19216 18796 19256
rect 18836 19216 18837 19256
rect 18795 19207 18837 19216
rect 18699 19172 18741 19181
rect 18699 19132 18700 19172
rect 18740 19132 18741 19172
rect 18699 19123 18741 19132
rect 18700 19038 18740 19123
rect 18796 18593 18836 19207
rect 19372 19206 19412 19291
rect 19180 19088 19220 19097
rect 18795 18584 18837 18593
rect 18795 18544 18796 18584
rect 18836 18544 18837 18584
rect 18795 18535 18837 18544
rect 18796 18450 18836 18535
rect 19180 18341 19220 19048
rect 19660 19004 19700 19468
rect 19756 19340 19796 19349
rect 19756 19181 19796 19300
rect 19948 19256 19988 20560
rect 20044 20551 20084 20560
rect 20811 20600 20853 20609
rect 20811 20560 20812 20600
rect 20852 20560 20853 20600
rect 20811 20551 20853 20560
rect 20048 20432 20416 20441
rect 20088 20392 20130 20432
rect 20170 20392 20212 20432
rect 20252 20392 20294 20432
rect 20334 20392 20376 20432
rect 20048 20383 20416 20392
rect 21004 20180 21044 26608
rect 21292 22625 21332 30379
rect 21291 22616 21333 22625
rect 21291 22576 21292 22616
rect 21332 22576 21333 22616
rect 21291 22567 21333 22576
rect 21099 21440 21141 21449
rect 21099 21400 21100 21440
rect 21140 21400 21141 21440
rect 21099 21391 21141 21400
rect 20908 20140 21044 20180
rect 20043 19928 20085 19937
rect 20043 19888 20044 19928
rect 20084 19888 20085 19928
rect 20043 19879 20085 19888
rect 20044 19794 20084 19879
rect 19852 19216 19988 19256
rect 20619 19256 20661 19265
rect 20619 19216 20620 19256
rect 20660 19216 20661 19256
rect 19755 19172 19797 19181
rect 19755 19132 19756 19172
rect 19796 19132 19797 19172
rect 19755 19123 19797 19132
rect 19660 18964 19796 19004
rect 19468 18668 19508 18677
rect 19508 18628 19700 18668
rect 19468 18619 19508 18628
rect 19276 18570 19316 18579
rect 19179 18332 19221 18341
rect 19179 18292 19180 18332
rect 19220 18292 19221 18332
rect 19179 18283 19221 18292
rect 18808 18164 19176 18173
rect 18848 18124 18890 18164
rect 18930 18124 18972 18164
rect 19012 18124 19054 18164
rect 19094 18124 19136 18164
rect 18808 18115 19176 18124
rect 18700 17996 18740 18005
rect 18604 17956 18700 17996
rect 18700 17947 18740 17956
rect 18795 17996 18837 18005
rect 18795 17956 18796 17996
rect 18836 17956 18837 17996
rect 18795 17947 18837 17956
rect 18507 17912 18549 17921
rect 18507 17872 18508 17912
rect 18548 17872 18549 17912
rect 18507 17863 18549 17872
rect 18508 17753 18548 17863
rect 18507 17744 18549 17753
rect 18507 17704 18508 17744
rect 18548 17704 18549 17744
rect 18507 17695 18549 17704
rect 18412 17200 18548 17240
rect 18315 17156 18357 17165
rect 18315 17116 18316 17156
rect 18356 17116 18357 17156
rect 18315 17107 18357 17116
rect 18412 17030 18452 17039
rect 18315 16988 18357 16997
rect 18412 16988 18452 16990
rect 18315 16948 18316 16988
rect 18356 16948 18452 16988
rect 18315 16939 18357 16948
rect 18220 16820 18260 16829
rect 18260 16780 18356 16820
rect 18220 16771 18260 16780
rect 18219 16652 18261 16661
rect 18219 16612 18220 16652
rect 18260 16612 18261 16652
rect 18219 16603 18261 16612
rect 18220 16232 18260 16603
rect 18316 16241 18356 16780
rect 18220 16183 18260 16192
rect 18315 16232 18357 16241
rect 18315 16192 18316 16232
rect 18356 16192 18357 16232
rect 18315 16183 18357 16192
rect 18508 15728 18548 17200
rect 18796 16829 18836 17947
rect 19083 17912 19125 17921
rect 19083 17872 19084 17912
rect 19124 17872 19125 17912
rect 19083 17863 19125 17872
rect 19084 17778 19124 17863
rect 19276 17249 19316 18530
rect 19660 18500 19700 18628
rect 19660 18451 19700 18460
rect 19756 17912 19796 18964
rect 19852 18836 19892 19216
rect 20619 19207 20661 19216
rect 19947 19088 19989 19097
rect 19947 19048 19948 19088
rect 19988 19048 19989 19088
rect 19947 19039 19989 19048
rect 19948 18954 19988 19039
rect 20048 18920 20416 18929
rect 20088 18880 20130 18920
rect 20170 18880 20212 18920
rect 20252 18880 20294 18920
rect 20334 18880 20376 18920
rect 20048 18871 20416 18880
rect 19852 18796 19988 18836
rect 19851 18584 19893 18593
rect 19851 18544 19852 18584
rect 19892 18544 19893 18584
rect 19851 18535 19893 18544
rect 19852 18416 19892 18535
rect 19852 18367 19892 18376
rect 19564 17872 19796 17912
rect 19467 17744 19509 17753
rect 19467 17704 19468 17744
rect 19508 17704 19509 17744
rect 19467 17695 19509 17704
rect 19372 17660 19412 17669
rect 19275 17240 19317 17249
rect 19275 17200 19276 17240
rect 19316 17200 19317 17240
rect 19275 17191 19317 17200
rect 18795 16820 18837 16829
rect 18795 16780 18796 16820
rect 18836 16780 18837 16820
rect 18795 16771 18837 16780
rect 18808 16652 19176 16661
rect 18848 16612 18890 16652
rect 18930 16612 18972 16652
rect 19012 16612 19054 16652
rect 19094 16612 19136 16652
rect 18808 16603 19176 16612
rect 19372 16073 19412 17620
rect 19468 17610 19508 17695
rect 19468 16232 19508 16241
rect 19564 16232 19604 17872
rect 19756 17744 19796 17753
rect 19659 17660 19701 17669
rect 19659 17620 19660 17660
rect 19700 17620 19701 17660
rect 19659 17611 19701 17620
rect 19660 17072 19700 17611
rect 19660 17023 19700 17032
rect 19660 16400 19700 16409
rect 19756 16400 19796 17704
rect 19948 17669 19988 18796
rect 20044 18500 20084 18509
rect 20044 18089 20084 18460
rect 20236 18332 20276 18341
rect 20043 18080 20085 18089
rect 20043 18040 20044 18080
rect 20084 18040 20085 18080
rect 20043 18031 20085 18040
rect 20236 17921 20276 18292
rect 20235 17912 20277 17921
rect 20235 17872 20236 17912
rect 20276 17872 20277 17912
rect 20235 17863 20277 17872
rect 20523 17744 20565 17753
rect 20523 17704 20524 17744
rect 20564 17704 20565 17744
rect 20523 17695 20565 17704
rect 19947 17660 19989 17669
rect 19947 17620 19948 17660
rect 19988 17620 19989 17660
rect 19947 17611 19989 17620
rect 19947 17408 19989 17417
rect 19947 17368 19948 17408
rect 19988 17368 19989 17408
rect 19947 17359 19989 17368
rect 20048 17408 20416 17417
rect 20088 17368 20130 17408
rect 20170 17368 20212 17408
rect 20252 17368 20294 17408
rect 20334 17368 20376 17408
rect 20048 17359 20416 17368
rect 19851 17240 19893 17249
rect 19851 17200 19852 17240
rect 19892 17200 19893 17240
rect 19851 17191 19893 17200
rect 19852 17106 19892 17191
rect 19948 16988 19988 17359
rect 20044 16988 20084 16997
rect 19948 16948 20044 16988
rect 20044 16939 20084 16948
rect 20235 16904 20277 16913
rect 20235 16864 20236 16904
rect 20276 16864 20277 16904
rect 20235 16855 20277 16864
rect 20236 16770 20276 16855
rect 19700 16360 19796 16400
rect 19660 16351 19700 16360
rect 19948 16232 19988 16241
rect 19508 16192 19604 16232
rect 19756 16192 19948 16232
rect 19371 16064 19413 16073
rect 19371 16024 19372 16064
rect 19412 16024 19413 16064
rect 19371 16015 19413 16024
rect 18412 15688 18548 15728
rect 19083 15728 19125 15737
rect 19083 15688 19084 15728
rect 19124 15688 19125 15728
rect 18219 15392 18261 15401
rect 18219 15352 18220 15392
rect 18260 15352 18261 15392
rect 18219 15343 18261 15352
rect 18220 14048 18260 15343
rect 18412 14477 18452 15688
rect 19083 15679 19125 15688
rect 18987 15644 19029 15653
rect 18987 15604 18988 15644
rect 19028 15604 19029 15644
rect 18987 15595 19029 15604
rect 18508 15560 18548 15569
rect 18508 14981 18548 15520
rect 18604 15560 18644 15569
rect 18604 15149 18644 15520
rect 18988 15560 19028 15595
rect 18988 15509 19028 15520
rect 19084 15485 19124 15679
rect 19468 15546 19508 16192
rect 19659 16148 19701 16157
rect 19659 16108 19660 16148
rect 19700 16108 19701 16148
rect 19659 16099 19701 16108
rect 19276 15506 19508 15546
rect 19563 15560 19605 15569
rect 19563 15520 19564 15560
rect 19604 15520 19605 15560
rect 19563 15511 19605 15520
rect 19083 15476 19125 15485
rect 19083 15436 19084 15476
rect 19124 15436 19125 15476
rect 19083 15427 19125 15436
rect 19084 15342 19124 15427
rect 18603 15140 18645 15149
rect 18603 15100 18604 15140
rect 18644 15100 18645 15140
rect 18603 15091 18645 15100
rect 18808 15140 19176 15149
rect 18848 15100 18890 15140
rect 18930 15100 18972 15140
rect 19012 15100 19054 15140
rect 19094 15100 19136 15140
rect 18808 15091 19176 15100
rect 18507 14972 18549 14981
rect 18507 14932 18508 14972
rect 18548 14932 18549 14972
rect 18507 14923 18549 14932
rect 19083 14972 19125 14981
rect 19276 14972 19316 15506
rect 19564 15426 19604 15511
rect 19563 15224 19605 15233
rect 19660 15224 19700 16099
rect 19563 15184 19564 15224
rect 19604 15184 19700 15224
rect 19563 15175 19605 15184
rect 19083 14932 19084 14972
rect 19124 14932 19125 14972
rect 19083 14923 19125 14932
rect 19180 14932 19316 14972
rect 19371 14972 19413 14981
rect 19371 14932 19372 14972
rect 19412 14932 19413 14972
rect 18411 14468 18453 14477
rect 18411 14428 18412 14468
rect 18452 14428 18453 14468
rect 18411 14419 18453 14428
rect 18411 14216 18453 14225
rect 18411 14176 18412 14216
rect 18452 14176 18453 14216
rect 18411 14167 18453 14176
rect 18412 14082 18452 14167
rect 18220 13301 18260 14008
rect 18508 14048 18548 14923
rect 19084 14838 19124 14923
rect 18892 14720 18932 14729
rect 19180 14720 19220 14932
rect 19371 14923 19413 14932
rect 18932 14680 19220 14720
rect 19372 14720 19412 14923
rect 18603 14636 18645 14645
rect 18603 14596 18604 14636
rect 18644 14596 18645 14636
rect 18603 14587 18645 14596
rect 18604 14477 18644 14587
rect 18603 14468 18645 14477
rect 18603 14428 18604 14468
rect 18644 14428 18645 14468
rect 18603 14419 18645 14428
rect 18699 14384 18741 14393
rect 18699 14344 18700 14384
rect 18740 14344 18741 14384
rect 18699 14335 18741 14344
rect 18508 13999 18548 14008
rect 18700 14048 18740 14335
rect 18892 14057 18932 14680
rect 19372 14671 19412 14680
rect 19467 14720 19509 14729
rect 19467 14680 19468 14720
rect 19508 14680 19509 14720
rect 19467 14671 19509 14680
rect 19564 14720 19604 15175
rect 19756 14972 19796 16192
rect 19948 16183 19988 16192
rect 20044 16232 20084 16241
rect 19851 16064 19893 16073
rect 20044 16064 20084 16192
rect 20140 16211 20180 16220
rect 20140 16073 20180 16171
rect 19851 16024 19852 16064
rect 19892 16024 19893 16064
rect 19851 16015 19893 16024
rect 19948 16024 20084 16064
rect 20139 16064 20181 16073
rect 20139 16024 20140 16064
rect 20180 16024 20181 16064
rect 19852 15930 19892 16015
rect 19851 15728 19893 15737
rect 19851 15688 19852 15728
rect 19892 15688 19893 15728
rect 19851 15679 19893 15688
rect 19852 15485 19892 15679
rect 19851 15476 19893 15485
rect 19851 15436 19852 15476
rect 19892 15436 19893 15476
rect 19851 15427 19893 15436
rect 19756 14923 19796 14932
rect 19948 14972 19988 16024
rect 20139 16015 20181 16024
rect 20048 15896 20416 15905
rect 20088 15856 20130 15896
rect 20170 15856 20212 15896
rect 20252 15856 20294 15896
rect 20334 15856 20376 15896
rect 20048 15847 20416 15856
rect 20236 15728 20276 15737
rect 20524 15728 20564 17695
rect 20276 15688 20564 15728
rect 20236 15679 20276 15688
rect 20620 15644 20660 19207
rect 20908 16577 20948 20140
rect 21100 17249 21140 21391
rect 21291 18836 21333 18845
rect 21291 18796 21292 18836
rect 21332 18796 21333 18836
rect 21291 18787 21333 18796
rect 21099 17240 21141 17249
rect 21099 17200 21100 17240
rect 21140 17200 21141 17240
rect 21099 17191 21141 17200
rect 20907 16568 20949 16577
rect 20907 16528 20908 16568
rect 20948 16528 20949 16568
rect 20907 16519 20949 16528
rect 20524 15604 20660 15644
rect 20044 15546 20084 15555
rect 20044 15233 20084 15506
rect 20043 15224 20085 15233
rect 20043 15184 20044 15224
rect 20084 15184 20085 15224
rect 20043 15175 20085 15184
rect 19948 14923 19988 14932
rect 20139 14972 20181 14981
rect 20139 14932 20140 14972
rect 20180 14932 20181 14972
rect 20139 14923 20181 14932
rect 20140 14734 20180 14923
rect 19468 14586 19508 14671
rect 19564 14141 19604 14680
rect 19948 14720 19988 14729
rect 20140 14685 20180 14694
rect 20236 14720 20276 14729
rect 19948 14225 19988 14680
rect 20236 14561 20276 14680
rect 20235 14552 20277 14561
rect 20235 14512 20236 14552
rect 20276 14512 20277 14552
rect 20235 14503 20277 14512
rect 20048 14384 20416 14393
rect 20088 14344 20130 14384
rect 20170 14344 20212 14384
rect 20252 14344 20294 14384
rect 20334 14344 20376 14384
rect 20048 14335 20416 14344
rect 19947 14216 19989 14225
rect 19947 14176 19948 14216
rect 19988 14176 19989 14216
rect 19947 14167 19989 14176
rect 19563 14132 19605 14141
rect 19563 14092 19564 14132
rect 19604 14092 19605 14132
rect 19563 14083 19605 14092
rect 20139 14132 20181 14141
rect 20139 14092 20140 14132
rect 20180 14092 20181 14132
rect 20139 14083 20181 14092
rect 18700 13999 18740 14008
rect 18891 14048 18933 14057
rect 18891 14008 18892 14048
rect 18932 14008 18933 14048
rect 18891 13999 18933 14008
rect 19947 14048 19989 14057
rect 19947 14008 19948 14048
rect 19988 14008 19989 14048
rect 19947 13999 19989 14008
rect 18808 13628 19176 13637
rect 18848 13588 18890 13628
rect 18930 13588 18972 13628
rect 19012 13588 19054 13628
rect 19094 13588 19136 13628
rect 18808 13579 19176 13588
rect 18219 13292 18261 13301
rect 18219 13252 18220 13292
rect 18260 13252 18261 13292
rect 18219 13243 18261 13252
rect 18603 13208 18645 13217
rect 19084 13208 19124 13217
rect 18603 13168 18604 13208
rect 18644 13168 18645 13208
rect 18603 13159 18645 13168
rect 18988 13168 19084 13208
rect 18123 13040 18165 13049
rect 18123 13000 18124 13040
rect 18164 13000 18165 13040
rect 18123 12991 18165 13000
rect 17931 12200 17973 12209
rect 17931 12160 17932 12200
rect 17972 12160 17973 12200
rect 17931 12151 17973 12160
rect 18028 11948 18068 12496
rect 18124 12536 18164 12545
rect 18124 12032 18164 12496
rect 18219 12536 18261 12545
rect 18219 12496 18220 12536
rect 18260 12496 18261 12536
rect 18219 12487 18261 12496
rect 18412 12536 18452 12545
rect 18220 12402 18260 12487
rect 18412 12293 18452 12496
rect 18411 12284 18453 12293
rect 18411 12244 18412 12284
rect 18452 12244 18453 12284
rect 18411 12235 18453 12244
rect 18124 11992 18548 12032
rect 18508 11948 18548 11992
rect 18028 11908 18260 11948
rect 18123 11696 18165 11705
rect 18123 11656 18124 11696
rect 18164 11656 18165 11696
rect 18123 11647 18165 11656
rect 18124 11562 18164 11647
rect 17740 11404 17876 11444
rect 17740 11360 17780 11404
rect 17644 11320 17780 11360
rect 17355 11108 17397 11117
rect 17355 11068 17356 11108
rect 17396 11068 17397 11108
rect 17355 11059 17397 11068
rect 17356 10277 17396 11059
rect 17355 10268 17397 10277
rect 17355 10228 17356 10268
rect 17396 10228 17397 10268
rect 17355 10219 17397 10228
rect 17164 9521 17204 9606
rect 16972 9512 17012 9521
rect 16972 8933 17012 9472
rect 17068 9512 17108 9521
rect 17068 9353 17108 9472
rect 17163 9512 17205 9521
rect 17163 9472 17164 9512
rect 17204 9472 17205 9512
rect 17163 9463 17205 9472
rect 17260 9512 17300 9521
rect 17067 9344 17109 9353
rect 17067 9304 17068 9344
rect 17108 9304 17109 9344
rect 17067 9295 17109 9304
rect 17260 9017 17300 9472
rect 17259 9008 17301 9017
rect 17259 8968 17260 9008
rect 17300 8968 17301 9008
rect 17259 8959 17301 8968
rect 16971 8924 17013 8933
rect 16971 8884 16972 8924
rect 17012 8884 17013 8924
rect 16971 8875 17013 8884
rect 17356 8672 17396 10219
rect 17451 10184 17493 10193
rect 17451 10144 17452 10184
rect 17492 10144 17493 10184
rect 17451 10135 17493 10144
rect 17452 10050 17492 10135
rect 17644 10100 17684 11320
rect 17739 11192 17781 11201
rect 17739 11152 17740 11192
rect 17780 11152 17781 11192
rect 17739 11143 17781 11152
rect 17548 10060 17684 10100
rect 17740 11024 17780 11143
rect 18027 11108 18069 11117
rect 18027 11068 18028 11108
rect 18068 11068 18069 11108
rect 18027 11059 18069 11068
rect 17548 9521 17588 10060
rect 17740 9941 17780 10984
rect 17835 11024 17877 11033
rect 17835 10984 17836 11024
rect 17876 10984 17877 11024
rect 17835 10975 17877 10984
rect 18028 11024 18068 11059
rect 17836 10890 17876 10975
rect 18028 10973 18068 10984
rect 17931 10940 17973 10949
rect 17931 10900 17932 10940
rect 17972 10900 17973 10940
rect 17931 10891 17973 10900
rect 17932 10613 17972 10891
rect 18027 10856 18069 10865
rect 18027 10816 18028 10856
rect 18068 10816 18069 10856
rect 18027 10807 18069 10816
rect 18028 10722 18068 10807
rect 18220 10688 18260 11908
rect 18508 11899 18548 11908
rect 18315 11612 18357 11621
rect 18315 11572 18316 11612
rect 18356 11572 18357 11612
rect 18315 11563 18357 11572
rect 18316 11024 18356 11563
rect 18316 10975 18356 10984
rect 18412 11024 18452 11033
rect 18220 10648 18356 10688
rect 17931 10604 17973 10613
rect 17931 10564 17932 10604
rect 17972 10564 17973 10604
rect 17931 10555 17973 10564
rect 18219 10520 18261 10529
rect 18219 10480 18220 10520
rect 18260 10480 18261 10520
rect 18219 10471 18261 10480
rect 18123 10268 18165 10277
rect 18123 10228 18124 10268
rect 18164 10228 18165 10268
rect 18123 10219 18165 10228
rect 18124 10109 18164 10219
rect 18123 10100 18165 10109
rect 18123 10060 18124 10100
rect 18164 10060 18165 10100
rect 18123 10051 18165 10060
rect 17739 9932 17781 9941
rect 17739 9892 17740 9932
rect 17780 9892 17781 9932
rect 17739 9883 17781 9892
rect 17740 9689 17780 9883
rect 17739 9680 17781 9689
rect 17739 9640 17740 9680
rect 17780 9640 17781 9680
rect 17739 9631 17781 9640
rect 18028 9605 18068 9636
rect 17643 9596 17685 9605
rect 17643 9556 17644 9596
rect 17684 9556 17685 9596
rect 17643 9547 17685 9556
rect 18027 9596 18069 9605
rect 18027 9556 18028 9596
rect 18068 9556 18069 9596
rect 18027 9547 18069 9556
rect 17547 9512 17589 9521
rect 17547 9472 17548 9512
rect 17588 9472 17589 9512
rect 17547 9463 17589 9472
rect 17644 9512 17684 9547
rect 17644 9461 17684 9472
rect 18028 9512 18068 9547
rect 17451 9344 17493 9353
rect 17451 9304 17452 9344
rect 17492 9304 17493 9344
rect 17451 9295 17493 9304
rect 17643 9344 17685 9353
rect 17643 9304 17644 9344
rect 17684 9304 17685 9344
rect 17643 9295 17685 9304
rect 17452 9210 17492 9295
rect 17644 9210 17684 9295
rect 17739 9260 17781 9269
rect 17739 9220 17740 9260
rect 17780 9220 17781 9260
rect 17739 9211 17781 9220
rect 17451 8672 17493 8681
rect 17356 8632 17452 8672
rect 17492 8632 17493 8672
rect 17451 8623 17493 8632
rect 17452 8538 17492 8623
rect 17644 8504 17684 8513
rect 17644 8009 17684 8464
rect 17643 8000 17685 8009
rect 17643 7960 17644 8000
rect 17684 7960 17685 8000
rect 17643 7951 17685 7960
rect 16875 7832 16917 7841
rect 16875 7792 16876 7832
rect 16916 7792 16917 7832
rect 16875 7783 16917 7792
rect 16971 7748 17013 7757
rect 16971 7708 16972 7748
rect 17012 7708 17013 7748
rect 16971 7699 17013 7708
rect 16972 7614 17012 7699
rect 16780 7288 17012 7328
rect 16684 7111 16724 7120
rect 16395 7076 16437 7085
rect 16395 7036 16396 7076
rect 16436 7036 16437 7076
rect 16395 7027 16437 7036
rect 16396 7025 16436 7027
rect 16204 6943 16244 6952
rect 16492 6992 16532 7001
rect 16532 6952 16724 6992
rect 16492 6943 16532 6952
rect 16684 6714 16724 6952
rect 16684 6665 16724 6674
rect 16492 6488 16532 6497
rect 16300 6448 16492 6488
rect 16203 6236 16245 6245
rect 16203 6196 16204 6236
rect 16244 6196 16245 6236
rect 16203 6187 16245 6196
rect 16204 6102 16244 6187
rect 16300 5741 16340 6448
rect 16492 6439 16532 6448
rect 16588 6488 16628 6497
rect 16876 6488 16916 6497
rect 16628 6448 16724 6488
rect 16588 6439 16628 6448
rect 16587 6236 16629 6245
rect 16587 6196 16588 6236
rect 16628 6196 16629 6236
rect 16587 6187 16629 6196
rect 16395 5984 16437 5993
rect 16395 5944 16396 5984
rect 16436 5944 16437 5984
rect 16395 5935 16437 5944
rect 16299 5732 16341 5741
rect 16299 5692 16300 5732
rect 16340 5692 16341 5732
rect 16299 5683 16341 5692
rect 16396 5648 16436 5935
rect 16396 5599 16436 5608
rect 16299 5564 16341 5573
rect 16204 5524 16300 5564
rect 16340 5524 16341 5564
rect 16204 4649 16244 5524
rect 16299 5515 16341 5524
rect 16300 5430 16340 5515
rect 16491 5228 16533 5237
rect 16491 5188 16492 5228
rect 16532 5188 16533 5228
rect 16491 5179 16533 5188
rect 16492 5060 16532 5179
rect 16396 5020 16492 5060
rect 16299 4976 16341 4985
rect 16299 4936 16300 4976
rect 16340 4936 16341 4976
rect 16299 4927 16341 4936
rect 16300 4842 16340 4927
rect 16203 4640 16245 4649
rect 16203 4600 16204 4640
rect 16244 4600 16245 4640
rect 16203 4591 16245 4600
rect 16299 4388 16341 4397
rect 16299 4348 16300 4388
rect 16340 4348 16341 4388
rect 16299 4339 16341 4348
rect 16300 4254 16340 4339
rect 16396 4136 16436 5020
rect 16492 5011 16532 5020
rect 16588 4388 16628 6187
rect 16684 5741 16724 6448
rect 16780 6448 16876 6488
rect 16683 5732 16725 5741
rect 16683 5692 16684 5732
rect 16724 5692 16725 5732
rect 16683 5683 16725 5692
rect 16684 5648 16724 5683
rect 16684 5321 16724 5608
rect 16683 5312 16725 5321
rect 16683 5272 16684 5312
rect 16724 5272 16725 5312
rect 16683 5263 16725 5272
rect 16684 4976 16724 5263
rect 16780 5237 16820 6448
rect 16876 6439 16916 6448
rect 16875 6320 16917 6329
rect 16875 6280 16876 6320
rect 16916 6280 16917 6320
rect 16875 6271 16917 6280
rect 16876 6186 16916 6271
rect 16972 6068 17012 7288
rect 17067 6488 17109 6497
rect 17067 6448 17068 6488
rect 17108 6448 17109 6488
rect 17067 6439 17109 6448
rect 17164 6488 17204 6497
rect 17068 6245 17108 6439
rect 17067 6236 17109 6245
rect 17067 6196 17068 6236
rect 17108 6196 17109 6236
rect 17067 6187 17109 6196
rect 16876 6028 17012 6068
rect 16779 5228 16821 5237
rect 16779 5188 16780 5228
rect 16820 5188 16821 5228
rect 16779 5179 16821 5188
rect 16780 4976 16820 4985
rect 16684 4936 16780 4976
rect 16780 4927 16820 4936
rect 16876 4808 16916 6028
rect 16972 5816 17012 5825
rect 16972 5657 17012 5776
rect 16971 5648 17013 5657
rect 16971 5608 16972 5648
rect 17012 5608 17013 5648
rect 16971 5599 17013 5608
rect 17164 5396 17204 6448
rect 17644 6488 17684 6497
rect 17644 5825 17684 6448
rect 17740 6488 17780 9211
rect 17836 8672 17876 8683
rect 17836 8597 17876 8632
rect 17931 8672 17973 8681
rect 17931 8632 17932 8672
rect 17972 8632 17973 8672
rect 17931 8623 17973 8632
rect 17835 8588 17877 8597
rect 17835 8548 17836 8588
rect 17876 8548 17877 8588
rect 17835 8539 17877 8548
rect 17932 7160 17972 8623
rect 18028 8261 18068 9472
rect 18124 9512 18164 10051
rect 18124 8345 18164 9472
rect 18123 8336 18165 8345
rect 18123 8296 18124 8336
rect 18164 8296 18165 8336
rect 18123 8287 18165 8296
rect 18027 8252 18069 8261
rect 18027 8212 18028 8252
rect 18068 8212 18069 8252
rect 18027 8203 18069 8212
rect 18220 8084 18260 10471
rect 18316 8597 18356 10648
rect 18412 10277 18452 10984
rect 18507 10856 18549 10865
rect 18604 10856 18644 13159
rect 18988 12461 19028 13168
rect 19084 13159 19124 13168
rect 19563 13208 19605 13217
rect 19563 13168 19564 13208
rect 19604 13168 19605 13208
rect 19563 13159 19605 13168
rect 19660 13208 19700 13217
rect 19564 13074 19604 13159
rect 19276 13040 19316 13049
rect 19468 13040 19508 13049
rect 18987 12452 19029 12461
rect 18987 12412 18988 12452
rect 19028 12412 19029 12452
rect 18987 12403 19029 12412
rect 18699 12200 18741 12209
rect 18699 12160 18700 12200
rect 18740 12160 18741 12200
rect 18699 12151 18741 12160
rect 18700 11873 18740 12151
rect 18808 12116 19176 12125
rect 18848 12076 18890 12116
rect 18930 12076 18972 12116
rect 19012 12076 19054 12116
rect 19094 12076 19136 12116
rect 18808 12067 19176 12076
rect 18699 11864 18741 11873
rect 18699 11824 18700 11864
rect 18740 11824 18741 11864
rect 18699 11815 18741 11824
rect 19084 11864 19124 11873
rect 18700 11696 18740 11707
rect 19084 11705 19124 11824
rect 19276 11705 19316 13000
rect 19372 13000 19468 13040
rect 18700 11621 18740 11656
rect 19083 11696 19125 11705
rect 19083 11656 19084 11696
rect 19124 11656 19125 11696
rect 19083 11647 19125 11656
rect 19275 11696 19317 11705
rect 19275 11656 19276 11696
rect 19316 11656 19317 11696
rect 19275 11647 19317 11656
rect 19372 11696 19412 13000
rect 19468 12991 19508 13000
rect 19660 12704 19700 13168
rect 19564 12664 19700 12704
rect 19756 13208 19796 13217
rect 19756 12704 19796 13168
rect 19852 12704 19892 12713
rect 19756 12664 19852 12704
rect 19564 12545 19604 12664
rect 19852 12655 19892 12664
rect 19563 12536 19605 12545
rect 19563 12496 19564 12536
rect 19604 12496 19605 12536
rect 19563 12487 19605 12496
rect 19660 12536 19700 12545
rect 19660 12461 19700 12496
rect 19948 12461 19988 13999
rect 20140 13998 20180 14083
rect 20048 12872 20416 12881
rect 20088 12832 20130 12872
rect 20170 12832 20212 12872
rect 20252 12832 20294 12872
rect 20334 12832 20376 12872
rect 20048 12823 20416 12832
rect 19659 12452 19701 12461
rect 19659 12412 19660 12452
rect 19700 12412 19701 12452
rect 19659 12403 19701 12412
rect 19947 12452 19989 12461
rect 19947 12412 19948 12452
rect 19988 12412 19989 12452
rect 19947 12403 19989 12412
rect 19660 12041 19700 12403
rect 19852 12284 19892 12293
rect 19659 12032 19701 12041
rect 19659 11992 19660 12032
rect 19700 11992 19701 12032
rect 19659 11983 19701 11992
rect 19372 11647 19412 11656
rect 19468 11696 19508 11705
rect 18699 11612 18741 11621
rect 18699 11572 18700 11612
rect 18740 11572 18741 11612
rect 18699 11563 18741 11572
rect 19468 11201 19508 11656
rect 19755 11696 19797 11705
rect 19755 11656 19756 11696
rect 19796 11656 19797 11696
rect 19755 11647 19797 11656
rect 19756 11562 19796 11647
rect 19467 11192 19509 11201
rect 19467 11152 19468 11192
rect 19508 11152 19509 11192
rect 19467 11143 19509 11152
rect 18796 10949 18836 11034
rect 19852 11033 19892 12244
rect 20140 11864 20180 11873
rect 19948 11824 20140 11864
rect 19948 11117 19988 11824
rect 20140 11815 20180 11824
rect 20043 11696 20085 11705
rect 20043 11656 20044 11696
rect 20084 11656 20085 11696
rect 20043 11647 20085 11656
rect 20044 11562 20084 11647
rect 20048 11360 20416 11369
rect 20088 11320 20130 11360
rect 20170 11320 20212 11360
rect 20252 11320 20294 11360
rect 20334 11320 20376 11360
rect 20048 11311 20416 11320
rect 20043 11192 20085 11201
rect 20043 11152 20044 11192
rect 20084 11152 20085 11192
rect 20043 11143 20085 11152
rect 19947 11108 19989 11117
rect 19947 11068 19948 11108
rect 19988 11068 19989 11108
rect 19947 11059 19989 11068
rect 20044 11058 20084 11143
rect 19372 11024 19412 11033
rect 18795 10940 18837 10949
rect 18795 10900 18796 10940
rect 18836 10900 18837 10940
rect 18795 10891 18837 10900
rect 18892 10940 18932 10949
rect 18507 10816 18508 10856
rect 18548 10816 18644 10856
rect 18507 10807 18549 10816
rect 18892 10772 18932 10900
rect 18604 10732 18932 10772
rect 18507 10604 18549 10613
rect 18507 10564 18508 10604
rect 18548 10564 18549 10604
rect 18507 10555 18549 10564
rect 18411 10268 18453 10277
rect 18411 10228 18412 10268
rect 18452 10228 18453 10268
rect 18411 10219 18453 10228
rect 18508 9437 18548 10555
rect 18507 9428 18549 9437
rect 18507 9388 18508 9428
rect 18548 9388 18549 9428
rect 18507 9379 18549 9388
rect 18604 9428 18644 10732
rect 18808 10604 19176 10613
rect 18848 10564 18890 10604
rect 18930 10564 18972 10604
rect 19012 10564 19054 10604
rect 19094 10564 19136 10604
rect 18808 10555 19176 10564
rect 19372 10436 19412 10984
rect 19851 11024 19893 11033
rect 19851 10979 19852 11024
rect 19892 10979 19893 11024
rect 19851 10975 19893 10979
rect 19852 10889 19892 10975
rect 19372 10396 19892 10436
rect 19083 10352 19125 10361
rect 19083 10312 19084 10352
rect 19124 10312 19125 10352
rect 19083 10303 19125 10312
rect 19276 10312 19796 10352
rect 19084 10218 19124 10303
rect 18699 10184 18741 10193
rect 18699 10144 18700 10184
rect 18740 10144 18741 10184
rect 18699 10135 18741 10144
rect 18700 10050 18740 10135
rect 18891 10100 18933 10109
rect 18891 10060 18892 10100
rect 18932 10060 18933 10100
rect 18891 10051 18933 10060
rect 18892 9966 18932 10051
rect 19083 9512 19125 9521
rect 19083 9472 19084 9512
rect 19124 9472 19125 9512
rect 19083 9463 19125 9472
rect 18644 9388 18740 9428
rect 18604 9379 18644 9388
rect 18603 9008 18645 9017
rect 18603 8968 18604 9008
rect 18644 8968 18645 9008
rect 18603 8959 18645 8968
rect 18315 8588 18357 8597
rect 18315 8548 18316 8588
rect 18356 8548 18357 8588
rect 18315 8539 18357 8548
rect 18604 8168 18644 8959
rect 18604 8119 18644 8128
rect 18124 8044 18260 8084
rect 17932 7111 17972 7120
rect 18028 8000 18068 8009
rect 18028 7916 18068 7960
rect 18124 7916 18164 8044
rect 18316 8000 18356 8009
rect 18316 7916 18356 7960
rect 18507 8000 18549 8009
rect 18507 7960 18508 8000
rect 18548 7960 18549 8000
rect 18507 7951 18549 7960
rect 18028 7876 18164 7916
rect 18220 7876 18356 7916
rect 17740 6245 17780 6448
rect 17835 6488 17877 6497
rect 17835 6448 17836 6488
rect 17876 6448 17877 6488
rect 17835 6439 17877 6448
rect 18028 6483 18068 7876
rect 18124 7076 18164 7085
rect 18220 7076 18260 7876
rect 18508 7866 18548 7951
rect 18316 7748 18356 7757
rect 18356 7708 18548 7748
rect 18316 7699 18356 7708
rect 18315 7412 18357 7421
rect 18315 7372 18316 7412
rect 18356 7372 18357 7412
rect 18315 7363 18357 7372
rect 18316 7160 18356 7363
rect 18316 7111 18356 7120
rect 18164 7036 18260 7076
rect 18124 7027 18164 7036
rect 18220 6488 18260 7036
rect 18411 6740 18453 6749
rect 18411 6700 18412 6740
rect 18452 6700 18453 6740
rect 18411 6691 18453 6700
rect 18316 6488 18356 6497
rect 18028 6443 18164 6483
rect 18220 6448 18316 6488
rect 17836 6354 17876 6439
rect 17931 6404 17973 6413
rect 17931 6364 17932 6404
rect 17972 6364 17973 6404
rect 17931 6355 17973 6364
rect 17739 6236 17781 6245
rect 17739 6196 17740 6236
rect 17780 6196 17781 6236
rect 17739 6187 17781 6196
rect 17643 5816 17685 5825
rect 17356 5741 17396 5786
rect 17643 5776 17644 5816
rect 17684 5776 17685 5816
rect 17643 5767 17685 5776
rect 17355 5732 17397 5741
rect 17355 5692 17356 5732
rect 17396 5692 17397 5732
rect 17355 5691 17397 5692
rect 17355 5683 17356 5691
rect 17259 5648 17301 5657
rect 17259 5608 17260 5648
rect 17300 5608 17301 5648
rect 17396 5683 17397 5691
rect 17932 5693 17972 6355
rect 18027 6320 18069 6329
rect 18027 6280 18028 6320
rect 18068 6280 18069 6320
rect 18027 6271 18069 6280
rect 18028 6186 18068 6271
rect 18027 5984 18069 5993
rect 18027 5944 18028 5984
rect 18068 5944 18069 5984
rect 18027 5935 18069 5944
rect 17356 5642 17396 5651
rect 17643 5648 17685 5657
rect 17740 5656 17780 5665
rect 17259 5599 17301 5608
rect 17643 5608 17644 5648
rect 17684 5608 17685 5648
rect 17643 5599 17685 5608
rect 17732 5616 17740 5656
rect 17732 5607 17780 5616
rect 17836 5648 17876 5657
rect 17876 5608 17877 5648
rect 17932 5644 17972 5653
rect 17260 5514 17300 5599
rect 17644 5514 17684 5599
rect 17452 5422 17492 5431
rect 17732 5422 17772 5607
rect 17836 5599 17877 5608
rect 17837 5564 17877 5599
rect 17931 5564 17973 5573
rect 17837 5524 17932 5564
rect 17972 5524 17973 5564
rect 17931 5515 17973 5524
rect 17164 5356 17300 5396
rect 17492 5382 17588 5422
rect 17452 5373 17492 5382
rect 17067 4976 17109 4985
rect 17067 4936 17068 4976
rect 17108 4936 17109 4976
rect 17067 4927 17109 4936
rect 17164 4934 17204 4943
rect 17068 4842 17108 4927
rect 17163 4894 17164 4901
rect 17204 4894 17205 4901
rect 17163 4892 17205 4894
rect 17163 4852 17164 4892
rect 17204 4852 17205 4892
rect 17163 4843 17205 4852
rect 16588 4339 16628 4348
rect 16684 4768 16916 4808
rect 17164 4799 17204 4843
rect 17260 4808 17300 5356
rect 17452 4808 17492 4817
rect 17260 4768 17452 4808
rect 16684 4313 16724 4768
rect 17452 4759 17492 4768
rect 17548 4724 17588 5382
rect 17644 5382 17772 5422
rect 17644 5069 17684 5382
rect 17643 5060 17685 5069
rect 17643 5020 17644 5060
rect 17684 5020 17685 5060
rect 17643 5011 17685 5020
rect 17739 4976 17781 4985
rect 17739 4936 17740 4976
rect 17780 4936 17781 4976
rect 17739 4927 17781 4936
rect 17931 4976 17973 4985
rect 17931 4936 17932 4976
rect 17972 4936 17973 4976
rect 17931 4927 17973 4936
rect 17740 4842 17780 4927
rect 17932 4733 17972 4927
rect 17644 4724 17684 4733
rect 17548 4684 17644 4724
rect 17355 4640 17397 4649
rect 17355 4600 17356 4640
rect 17396 4600 17397 4640
rect 17355 4591 17397 4600
rect 16683 4304 16725 4313
rect 16683 4264 16684 4304
rect 16724 4264 16725 4304
rect 16683 4255 16725 4264
rect 16396 4087 16436 4096
rect 16683 4136 16725 4145
rect 16683 4096 16684 4136
rect 16724 4096 16725 4136
rect 16683 4087 16725 4096
rect 16971 4136 17013 4145
rect 16971 4096 16972 4136
rect 17012 4096 17013 4136
rect 16971 4087 17013 4096
rect 17259 4136 17301 4145
rect 17259 4096 17260 4136
rect 17300 4096 17301 4136
rect 17259 4087 17301 4096
rect 17356 4136 17396 4591
rect 17356 4087 17396 4096
rect 16684 4002 16724 4087
rect 16203 3716 16245 3725
rect 16203 3676 16204 3716
rect 16244 3676 16245 3716
rect 16203 3667 16245 3676
rect 16875 3716 16917 3725
rect 16875 3676 16876 3716
rect 16916 3676 16917 3716
rect 16875 3667 16917 3676
rect 16204 3506 16244 3667
rect 16204 3457 16244 3466
rect 16588 3464 16628 3473
rect 16052 3340 16148 3380
rect 16300 3380 16340 3389
rect 16012 3331 16052 3340
rect 16300 3305 16340 3340
rect 16492 3380 16532 3389
rect 16299 3296 16341 3305
rect 16299 3256 16300 3296
rect 16340 3256 16341 3296
rect 16299 3247 16341 3256
rect 16396 3296 16436 3305
rect 16300 3245 16340 3247
rect 16204 2876 16244 2885
rect 15916 2836 16204 2876
rect 16204 2827 16244 2836
rect 15819 2792 15861 2801
rect 15819 2752 15820 2792
rect 15860 2752 15861 2792
rect 15819 2743 15861 2752
rect 15723 2624 15765 2633
rect 15723 2584 15724 2624
rect 15764 2584 15765 2624
rect 15723 2575 15765 2584
rect 15532 2500 15668 2540
rect 15531 1196 15573 1205
rect 15531 1156 15532 1196
rect 15572 1156 15573 1196
rect 15531 1147 15573 1156
rect 15532 1062 15572 1147
rect 15628 80 15668 2500
rect 15723 2288 15765 2297
rect 15723 2248 15724 2288
rect 15764 2248 15765 2288
rect 15723 2239 15765 2248
rect 15724 1112 15764 2239
rect 15724 1063 15764 1072
rect 15820 80 15860 2743
rect 16012 2633 16052 2718
rect 16011 2624 16053 2633
rect 16396 2624 16436 3256
rect 16492 2969 16532 3340
rect 16588 3053 16628 3424
rect 16779 3296 16821 3305
rect 16779 3256 16780 3296
rect 16820 3256 16821 3296
rect 16779 3247 16821 3256
rect 16780 3162 16820 3247
rect 16587 3044 16629 3053
rect 16587 3004 16588 3044
rect 16628 3004 16629 3044
rect 16587 2995 16629 3004
rect 16491 2960 16533 2969
rect 16491 2920 16492 2960
rect 16532 2920 16533 2960
rect 16491 2911 16533 2920
rect 16491 2792 16533 2801
rect 16491 2752 16492 2792
rect 16532 2752 16533 2792
rect 16491 2743 16533 2752
rect 16011 2584 16012 2624
rect 16052 2584 16148 2624
rect 16011 2575 16053 2584
rect 16011 1700 16053 1709
rect 16011 1660 16012 1700
rect 16052 1660 16053 1700
rect 16011 1651 16053 1660
rect 16012 80 16052 1651
rect 16108 785 16148 2584
rect 16300 2584 16436 2624
rect 16492 2624 16532 2743
rect 16300 1784 16340 2584
rect 16492 2575 16532 2584
rect 16588 2624 16628 2635
rect 16684 2633 16724 2718
rect 16588 2549 16628 2584
rect 16683 2624 16725 2633
rect 16683 2584 16684 2624
rect 16724 2584 16725 2624
rect 16683 2575 16725 2584
rect 16587 2540 16629 2549
rect 16587 2500 16588 2540
rect 16628 2500 16629 2540
rect 16587 2491 16629 2500
rect 16396 2456 16436 2465
rect 16396 1961 16436 2416
rect 16491 2456 16533 2465
rect 16491 2416 16492 2456
rect 16532 2416 16533 2456
rect 16491 2407 16533 2416
rect 16395 1952 16437 1961
rect 16395 1912 16396 1952
rect 16436 1912 16437 1952
rect 16395 1903 16437 1912
rect 16492 1952 16532 2407
rect 16587 2372 16629 2381
rect 16587 2332 16588 2372
rect 16628 2332 16629 2372
rect 16587 2323 16629 2332
rect 16492 1793 16532 1912
rect 16491 1784 16533 1793
rect 16300 1744 16436 1784
rect 16203 1448 16245 1457
rect 16203 1408 16204 1448
rect 16244 1408 16245 1448
rect 16203 1399 16245 1408
rect 16107 776 16149 785
rect 16107 736 16108 776
rect 16148 736 16149 776
rect 16107 727 16149 736
rect 16204 80 16244 1399
rect 16396 1205 16436 1744
rect 16491 1744 16492 1784
rect 16532 1744 16533 1784
rect 16491 1735 16533 1744
rect 16395 1196 16437 1205
rect 16395 1156 16396 1196
rect 16436 1156 16437 1196
rect 16395 1147 16437 1156
rect 16395 1028 16437 1037
rect 16395 988 16396 1028
rect 16436 988 16437 1028
rect 16395 979 16437 988
rect 16396 80 16436 979
rect 16588 80 16628 2323
rect 16779 1868 16821 1877
rect 16779 1828 16780 1868
rect 16820 1828 16821 1868
rect 16779 1819 16821 1828
rect 16684 1700 16724 1709
rect 16780 1700 16820 1819
rect 16876 1784 16916 3667
rect 16972 3473 17012 4087
rect 17260 4002 17300 4087
rect 17548 3884 17588 4684
rect 17644 4675 17684 4684
rect 17931 4724 17973 4733
rect 17931 4684 17932 4724
rect 17972 4684 17973 4724
rect 17931 4675 17973 4684
rect 17644 4304 17684 4313
rect 17684 4264 17876 4304
rect 17644 4255 17684 4264
rect 17739 4136 17781 4145
rect 17739 4096 17740 4136
rect 17780 4096 17781 4136
rect 17739 4087 17781 4096
rect 17260 3844 17588 3884
rect 17067 3716 17109 3725
rect 17067 3676 17068 3716
rect 17108 3676 17109 3716
rect 17067 3667 17109 3676
rect 17260 3690 17300 3844
rect 16971 3464 17013 3473
rect 16971 3424 16972 3464
rect 17012 3424 17013 3464
rect 16971 3415 17013 3424
rect 17068 3464 17108 3667
rect 17355 3716 17397 3725
rect 17355 3676 17356 3716
rect 17396 3676 17492 3716
rect 17355 3667 17397 3676
rect 17260 3641 17300 3650
rect 17452 3632 17492 3676
rect 17452 3583 17492 3592
rect 17548 3464 17588 3473
rect 17068 3415 17108 3424
rect 17164 3422 17204 3431
rect 16972 3296 17012 3415
rect 17164 3296 17204 3382
rect 16972 3256 17204 3296
rect 17355 3296 17397 3305
rect 17355 3256 17356 3296
rect 17396 3256 17397 3296
rect 16972 2633 17012 3256
rect 17355 3247 17397 3256
rect 16971 2624 17013 2633
rect 16971 2584 16972 2624
rect 17012 2584 17013 2624
rect 16971 2575 17013 2584
rect 17259 2624 17301 2633
rect 17259 2584 17260 2624
rect 17300 2584 17301 2624
rect 17259 2575 17301 2584
rect 17356 2624 17396 3247
rect 17548 3044 17588 3424
rect 17643 3464 17685 3473
rect 17643 3424 17644 3464
rect 17684 3424 17685 3464
rect 17643 3415 17685 3424
rect 17740 3464 17780 4087
rect 17740 3415 17780 3424
rect 17644 3330 17684 3415
rect 17452 3004 17588 3044
rect 17452 2801 17492 3004
rect 17836 2960 17876 4264
rect 18028 3977 18068 5935
rect 18124 4145 18164 6443
rect 18316 6320 18356 6448
rect 18412 6488 18452 6691
rect 18412 6439 18452 6448
rect 18316 6280 18452 6320
rect 18412 5825 18452 6280
rect 18411 5816 18453 5825
rect 18411 5776 18412 5816
rect 18452 5776 18453 5816
rect 18411 5767 18453 5776
rect 18316 5648 18356 5657
rect 18316 5489 18356 5608
rect 18315 5480 18357 5489
rect 18315 5440 18316 5480
rect 18356 5440 18357 5480
rect 18315 5431 18357 5440
rect 18412 5018 18452 5767
rect 18316 4976 18356 4985
rect 18412 4969 18452 4978
rect 18508 4976 18548 7708
rect 18700 6413 18740 9388
rect 19084 9378 19124 9463
rect 18808 9092 19176 9101
rect 18848 9052 18890 9092
rect 18930 9052 18972 9092
rect 19012 9052 19054 9092
rect 19094 9052 19136 9092
rect 18808 9043 19176 9052
rect 19276 8840 19316 10312
rect 19468 10228 19700 10268
rect 19468 10184 19508 10228
rect 19468 10135 19508 10144
rect 19276 8791 19316 8800
rect 19372 10100 19412 10109
rect 19083 8672 19125 8681
rect 19083 8632 19084 8672
rect 19124 8632 19125 8672
rect 19083 8623 19125 8632
rect 19084 8093 19124 8623
rect 19372 8504 19412 10060
rect 19563 10100 19605 10109
rect 19563 10060 19564 10100
rect 19604 10060 19605 10100
rect 19563 10051 19605 10060
rect 19564 9507 19604 10051
rect 19660 9680 19700 10228
rect 19756 10184 19796 10312
rect 19756 10135 19796 10144
rect 19756 9680 19796 9689
rect 19660 9640 19756 9680
rect 19756 9631 19796 9640
rect 19852 9521 19892 10396
rect 19947 10100 19989 10109
rect 19947 10060 19948 10100
rect 19988 10060 19989 10100
rect 19947 10051 19989 10060
rect 19948 9680 19988 10051
rect 20048 9848 20416 9857
rect 20088 9808 20130 9848
rect 20170 9808 20212 9848
rect 20252 9808 20294 9848
rect 20334 9808 20376 9848
rect 20048 9799 20416 9808
rect 20235 9680 20277 9689
rect 19948 9640 20180 9680
rect 19564 9428 19604 9467
rect 19851 9512 19893 9521
rect 19851 9472 19852 9512
rect 19892 9472 19893 9512
rect 19851 9463 19893 9472
rect 19948 9512 19988 9521
rect 20140 9518 20180 9640
rect 20235 9640 20236 9680
rect 20276 9640 20277 9680
rect 20235 9631 20277 9640
rect 19988 9472 20084 9512
rect 19948 9463 19988 9472
rect 19468 9388 19604 9428
rect 19468 8672 19508 9388
rect 19948 9260 19988 9269
rect 19660 9220 19948 9260
rect 19563 8924 19605 8933
rect 19563 8884 19564 8924
rect 19604 8884 19605 8924
rect 19563 8875 19605 8884
rect 19468 8623 19508 8632
rect 19564 8672 19604 8875
rect 19564 8623 19604 8632
rect 19660 8672 19700 9220
rect 19948 9211 19988 9220
rect 20044 9017 20084 9472
rect 20140 9469 20180 9478
rect 20236 9512 20276 9631
rect 20236 9463 20276 9472
rect 20043 9008 20085 9017
rect 20043 8968 20044 9008
rect 20084 8968 20085 9008
rect 20043 8959 20085 8968
rect 20524 8924 20564 15604
rect 20619 13544 20661 13553
rect 20619 13504 20620 13544
rect 20660 13504 20661 13544
rect 20619 13495 20661 13504
rect 20140 8884 20564 8924
rect 20140 8840 20180 8884
rect 20140 8791 20180 8800
rect 19947 8756 19989 8765
rect 19947 8716 19948 8756
rect 19988 8716 19989 8756
rect 19947 8707 19989 8716
rect 19660 8623 19700 8632
rect 19948 8622 19988 8707
rect 19756 8504 19796 8513
rect 19372 8464 19756 8504
rect 19756 8455 19796 8464
rect 20048 8336 20416 8345
rect 20088 8296 20130 8336
rect 20170 8296 20212 8336
rect 20252 8296 20294 8336
rect 20334 8296 20376 8336
rect 20048 8287 20416 8296
rect 19468 8212 19988 8252
rect 19275 8168 19317 8177
rect 19275 8128 19276 8168
rect 19316 8128 19317 8168
rect 19275 8119 19317 8128
rect 19083 8084 19125 8093
rect 19083 8044 19084 8084
rect 19124 8044 19125 8084
rect 19083 8035 19125 8044
rect 19084 7757 19124 7842
rect 19083 7748 19125 7757
rect 19083 7708 19084 7748
rect 19124 7708 19125 7748
rect 19083 7699 19125 7708
rect 18808 7580 19176 7589
rect 18848 7540 18890 7580
rect 18930 7540 18972 7580
rect 19012 7540 19054 7580
rect 19094 7540 19136 7580
rect 18808 7531 19176 7540
rect 18987 6740 19029 6749
rect 18987 6700 18988 6740
rect 19028 6700 19029 6740
rect 18987 6691 19029 6700
rect 18795 6656 18837 6665
rect 18795 6616 18796 6656
rect 18836 6616 18837 6656
rect 18795 6607 18837 6616
rect 18699 6404 18741 6413
rect 18699 6364 18700 6404
rect 18740 6364 18741 6404
rect 18699 6355 18741 6364
rect 18796 6404 18836 6607
rect 18891 6572 18933 6581
rect 18891 6532 18892 6572
rect 18932 6532 18933 6572
rect 18891 6523 18933 6532
rect 18796 6236 18836 6364
rect 18892 6488 18932 6523
rect 18892 6245 18932 6448
rect 18988 6413 19028 6691
rect 19276 6488 19316 8119
rect 19371 8000 19413 8009
rect 19371 7960 19372 8000
rect 19412 7960 19413 8000
rect 19371 7951 19413 7960
rect 19468 8000 19508 8212
rect 19563 8084 19605 8093
rect 19563 8044 19564 8084
rect 19604 8044 19605 8084
rect 19563 8035 19605 8044
rect 19468 7951 19508 7960
rect 19372 7866 19412 7951
rect 19564 7160 19604 8035
rect 19756 8000 19796 8009
rect 19756 7412 19796 7960
rect 19756 7363 19796 7372
rect 19372 6488 19412 6497
rect 19276 6448 19372 6488
rect 18987 6404 19029 6413
rect 18987 6364 18988 6404
rect 19028 6364 19029 6404
rect 18987 6355 19029 6364
rect 18700 6196 18836 6236
rect 18891 6236 18933 6245
rect 18891 6196 18892 6236
rect 18932 6196 18933 6236
rect 18604 4976 18644 4985
rect 18508 4936 18604 4976
rect 18316 4892 18356 4936
rect 18604 4927 18644 4936
rect 18316 4852 18452 4892
rect 18412 4649 18452 4852
rect 18603 4724 18645 4733
rect 18603 4684 18604 4724
rect 18644 4684 18645 4724
rect 18603 4675 18645 4684
rect 18411 4640 18453 4649
rect 18411 4600 18412 4640
rect 18452 4600 18453 4640
rect 18411 4591 18453 4600
rect 18604 4590 18644 4675
rect 18123 4136 18165 4145
rect 18123 4096 18124 4136
rect 18164 4096 18165 4136
rect 18123 4087 18165 4096
rect 18508 4136 18548 4145
rect 18027 3968 18069 3977
rect 18027 3928 18028 3968
rect 18068 3928 18069 3968
rect 18027 3919 18069 3928
rect 18027 3632 18069 3641
rect 18027 3592 18028 3632
rect 18068 3592 18069 3632
rect 18027 3583 18069 3592
rect 17548 2920 17876 2960
rect 17451 2792 17493 2801
rect 17451 2752 17452 2792
rect 17492 2752 17493 2792
rect 17451 2743 17493 2752
rect 17356 2575 17396 2584
rect 16972 2213 17012 2575
rect 17260 2490 17300 2575
rect 16971 2204 17013 2213
rect 16971 2164 16972 2204
rect 17012 2164 17013 2204
rect 16971 2155 17013 2164
rect 17259 2204 17301 2213
rect 17259 2164 17260 2204
rect 17300 2164 17301 2204
rect 17259 2155 17301 2164
rect 17163 1952 17205 1961
rect 17163 1912 17164 1952
rect 17204 1912 17205 1952
rect 17163 1903 17205 1912
rect 17260 1952 17300 2155
rect 17260 1903 17300 1912
rect 17356 2124 17396 2133
rect 17164 1818 17204 1903
rect 16876 1735 16916 1744
rect 17259 1784 17301 1793
rect 17259 1744 17260 1784
rect 17300 1744 17301 1784
rect 17259 1735 17301 1744
rect 16724 1660 16820 1700
rect 16684 1651 16724 1660
rect 17260 1373 17300 1735
rect 16683 1364 16725 1373
rect 16683 1324 16684 1364
rect 16724 1324 16725 1364
rect 16683 1315 16725 1324
rect 16971 1364 17013 1373
rect 16971 1324 16972 1364
rect 17012 1324 17013 1364
rect 16971 1315 17013 1324
rect 17259 1364 17301 1373
rect 17259 1324 17260 1364
rect 17300 1324 17301 1364
rect 17259 1315 17301 1324
rect 17356 1364 17396 2084
rect 17452 1448 17492 2743
rect 17548 1952 17588 2920
rect 17644 2792 17684 2801
rect 17684 2752 17876 2792
rect 17644 2743 17684 2752
rect 17836 2624 17876 2752
rect 17836 2575 17876 2584
rect 17932 2624 17972 2633
rect 17932 2120 17972 2584
rect 18028 2213 18068 3583
rect 18411 3548 18453 3557
rect 18411 3508 18412 3548
rect 18452 3508 18453 3548
rect 18411 3499 18453 3508
rect 18123 3464 18165 3473
rect 18123 3424 18124 3464
rect 18164 3424 18165 3464
rect 18123 3415 18165 3424
rect 18124 3330 18164 3415
rect 18219 3044 18261 3053
rect 18219 3004 18220 3044
rect 18260 3004 18261 3044
rect 18219 2995 18261 3004
rect 18123 2960 18165 2969
rect 18123 2920 18124 2960
rect 18164 2920 18165 2960
rect 18123 2911 18165 2920
rect 18124 2876 18164 2911
rect 18124 2825 18164 2836
rect 18124 2624 18164 2633
rect 18027 2204 18069 2213
rect 18027 2164 18028 2204
rect 18068 2164 18069 2204
rect 18027 2155 18069 2164
rect 17548 1903 17588 1912
rect 17644 2080 17972 2120
rect 17644 1952 17684 2080
rect 17644 1903 17684 1912
rect 17452 1408 17684 1448
rect 17356 1315 17396 1324
rect 16684 533 16724 1315
rect 16779 1280 16821 1289
rect 16779 1240 16780 1280
rect 16820 1240 16821 1280
rect 16779 1231 16821 1240
rect 16683 524 16725 533
rect 16683 484 16684 524
rect 16724 484 16725 524
rect 16683 475 16725 484
rect 16780 80 16820 1231
rect 16972 1112 17012 1315
rect 17164 1280 17204 1289
rect 17164 1121 17204 1240
rect 17547 1280 17589 1289
rect 17547 1240 17548 1280
rect 17588 1240 17589 1280
rect 17547 1231 17589 1240
rect 16972 80 17012 1072
rect 17163 1112 17205 1121
rect 17163 1072 17164 1112
rect 17204 1072 17205 1112
rect 17163 1063 17205 1072
rect 17452 1112 17492 1121
rect 17452 869 17492 1072
rect 17451 860 17493 869
rect 17451 820 17452 860
rect 17492 820 17493 860
rect 17451 811 17493 820
rect 17163 776 17205 785
rect 17163 736 17164 776
rect 17204 736 17205 776
rect 17163 727 17205 736
rect 17164 80 17204 727
rect 17355 524 17397 533
rect 17355 484 17356 524
rect 17396 484 17397 524
rect 17355 475 17397 484
rect 17356 80 17396 475
rect 17548 80 17588 1231
rect 17644 1121 17684 1408
rect 17740 1364 17780 2080
rect 18124 1961 18164 2584
rect 17836 1952 17876 1961
rect 18028 1952 18068 1961
rect 17876 1912 18028 1952
rect 17836 1903 17876 1912
rect 18028 1903 18068 1912
rect 18123 1952 18165 1961
rect 18123 1912 18124 1952
rect 18164 1912 18165 1952
rect 18123 1903 18165 1912
rect 17836 1784 17876 1793
rect 18220 1784 18260 2995
rect 18315 2876 18357 2885
rect 18315 2836 18316 2876
rect 18356 2836 18357 2876
rect 18315 2827 18357 2836
rect 17876 1744 18260 1784
rect 17836 1735 17876 1744
rect 17931 1532 17973 1541
rect 17931 1492 17932 1532
rect 17972 1492 17973 1532
rect 17931 1483 17973 1492
rect 17740 1315 17780 1324
rect 17643 1112 17685 1121
rect 17643 1072 17644 1112
rect 17684 1072 17685 1112
rect 17643 1063 17685 1072
rect 17644 978 17684 1063
rect 17739 944 17781 953
rect 17739 904 17740 944
rect 17780 904 17781 944
rect 17739 895 17781 904
rect 17740 80 17780 895
rect 17932 80 17972 1483
rect 18124 1112 18164 1121
rect 18316 1112 18356 2827
rect 18412 1952 18452 3499
rect 18508 2717 18548 4096
rect 18604 4136 18644 4145
rect 18700 4136 18740 6196
rect 18891 6187 18933 6196
rect 18808 6068 19176 6077
rect 18848 6028 18890 6068
rect 18930 6028 18972 6068
rect 19012 6028 19054 6068
rect 19094 6028 19136 6068
rect 18808 6019 19176 6028
rect 19083 4976 19125 4985
rect 19083 4936 19084 4976
rect 19124 4936 19125 4976
rect 19083 4927 19125 4936
rect 19084 4808 19124 4927
rect 19084 4759 19124 4768
rect 18808 4556 19176 4565
rect 18848 4516 18890 4556
rect 18930 4516 18972 4556
rect 19012 4516 19054 4556
rect 19094 4516 19136 4556
rect 18808 4507 19176 4516
rect 18795 4388 18837 4397
rect 19276 4388 19316 6448
rect 19372 6439 19412 6448
rect 19564 5648 19604 7120
rect 19948 6656 19988 8212
rect 20523 8000 20565 8009
rect 20523 7960 20524 8000
rect 20564 7960 20565 8000
rect 20523 7951 20565 7960
rect 20048 6824 20416 6833
rect 20088 6784 20130 6824
rect 20170 6784 20212 6824
rect 20252 6784 20294 6824
rect 20334 6784 20376 6824
rect 20048 6775 20416 6784
rect 20044 6656 20084 6665
rect 19948 6616 20044 6656
rect 20044 6607 20084 6616
rect 19851 6488 19893 6497
rect 19851 6443 19852 6488
rect 19892 6443 19893 6488
rect 19851 6439 19893 6443
rect 19659 6236 19701 6245
rect 19659 6196 19660 6236
rect 19700 6196 19701 6236
rect 19659 6187 19701 6196
rect 19372 4976 19412 4985
rect 19372 4565 19412 4936
rect 19467 4976 19509 4985
rect 19467 4936 19468 4976
rect 19508 4936 19509 4976
rect 19467 4927 19509 4936
rect 19468 4842 19508 4927
rect 19371 4556 19413 4565
rect 19371 4516 19372 4556
rect 19412 4516 19413 4556
rect 19371 4507 19413 4516
rect 18795 4348 18796 4388
rect 18836 4348 18837 4388
rect 18795 4339 18837 4348
rect 18988 4348 19316 4388
rect 18644 4096 18740 4136
rect 18604 2885 18644 4096
rect 18796 3212 18836 4339
rect 18988 4220 19028 4348
rect 19564 4304 19604 5608
rect 19660 5489 19700 6187
rect 19756 5900 19796 5909
rect 19852 5900 19892 6439
rect 20235 6320 20277 6329
rect 20235 6280 20236 6320
rect 20276 6280 20277 6320
rect 20235 6271 20277 6280
rect 20236 6068 20276 6271
rect 20140 6028 20276 6068
rect 19796 5860 19988 5900
rect 19756 5851 19796 5860
rect 19948 5648 19988 5860
rect 20140 5690 20180 6028
rect 20524 5900 20564 7951
rect 20620 7001 20660 13495
rect 21292 11201 21332 18787
rect 21387 15392 21429 15401
rect 21387 15352 21388 15392
rect 21428 15352 21429 15392
rect 21387 15343 21429 15352
rect 21291 11192 21333 11201
rect 21291 11152 21292 11192
rect 21332 11152 21333 11192
rect 21291 11143 21333 11152
rect 21388 7841 21428 15343
rect 21387 7832 21429 7841
rect 21387 7792 21388 7832
rect 21428 7792 21429 7832
rect 21387 7783 21429 7792
rect 20619 6992 20661 7001
rect 20619 6952 20620 6992
rect 20660 6952 20661 6992
rect 20619 6943 20661 6952
rect 19948 5599 19988 5608
rect 20044 5648 20084 5657
rect 20140 5641 20180 5650
rect 20236 5860 20564 5900
rect 20236 5648 20276 5860
rect 19659 5480 19701 5489
rect 20044 5480 20084 5608
rect 20236 5599 20276 5608
rect 19659 5440 19660 5480
rect 19700 5440 19701 5480
rect 19659 5431 19701 5440
rect 19948 5440 20084 5480
rect 19468 4264 19604 4304
rect 18988 4171 19028 4180
rect 19083 4220 19125 4229
rect 19468 4220 19508 4264
rect 19660 4229 19700 5431
rect 19756 4976 19796 4985
rect 19083 4180 19084 4220
rect 19124 4180 19125 4220
rect 19083 4171 19125 4180
rect 19372 4180 19508 4220
rect 19659 4220 19701 4229
rect 19659 4180 19660 4220
rect 19700 4180 19701 4220
rect 19084 4086 19124 4171
rect 19372 3464 19412 4180
rect 19659 4171 19701 4180
rect 19563 4136 19605 4145
rect 19563 4096 19564 4136
rect 19604 4096 19605 4136
rect 19563 4087 19605 4096
rect 19467 4052 19509 4061
rect 19467 4012 19468 4052
rect 19508 4012 19509 4052
rect 19467 4003 19509 4012
rect 19468 3464 19508 4003
rect 19564 4002 19604 4087
rect 19564 3632 19604 3641
rect 19756 3632 19796 4936
rect 19948 4733 19988 5440
rect 20048 5312 20416 5321
rect 20088 5272 20130 5312
rect 20170 5272 20212 5312
rect 20252 5272 20294 5312
rect 20334 5272 20376 5312
rect 20048 5263 20416 5272
rect 20235 4976 20277 4985
rect 20235 4936 20236 4976
rect 20276 4936 20277 4976
rect 20235 4927 20277 4936
rect 19947 4724 19989 4733
rect 19947 4684 19948 4724
rect 19988 4684 19989 4724
rect 19947 4675 19989 4684
rect 20044 4141 20084 4150
rect 20044 3968 20084 4101
rect 20236 4052 20276 4927
rect 20236 4003 20276 4012
rect 19604 3592 19796 3632
rect 19948 3928 20084 3968
rect 19564 3583 19604 3592
rect 19948 3548 19988 3928
rect 20048 3800 20416 3809
rect 20088 3760 20130 3800
rect 20170 3760 20212 3800
rect 20252 3760 20294 3800
rect 20334 3760 20376 3800
rect 20048 3751 20416 3760
rect 19852 3508 20084 3548
rect 19756 3464 19796 3473
rect 19468 3424 19756 3464
rect 19372 3380 19412 3424
rect 19756 3415 19796 3424
rect 19372 3340 19508 3380
rect 18700 3172 18836 3212
rect 18603 2876 18645 2885
rect 18603 2836 18604 2876
rect 18644 2836 18645 2876
rect 18700 2876 18740 3172
rect 19275 3128 19317 3137
rect 19275 3088 19276 3128
rect 19316 3088 19317 3128
rect 19275 3079 19317 3088
rect 18808 3044 19176 3053
rect 18848 3004 18890 3044
rect 18930 3004 18972 3044
rect 19012 3004 19054 3044
rect 19094 3004 19136 3044
rect 18808 2995 19176 3004
rect 18700 2836 18836 2876
rect 18603 2827 18645 2836
rect 18507 2708 18549 2717
rect 18507 2668 18508 2708
rect 18548 2668 18549 2708
rect 18507 2659 18549 2668
rect 18508 2624 18548 2659
rect 18604 2633 18644 2718
rect 18508 2574 18548 2584
rect 18603 2624 18645 2633
rect 18603 2584 18604 2624
rect 18644 2584 18645 2624
rect 18603 2575 18645 2584
rect 18700 2624 18740 2633
rect 18700 2456 18740 2584
rect 18796 2624 18836 2836
rect 18796 2575 18836 2584
rect 18988 2792 19028 2801
rect 18988 2540 19028 2752
rect 19179 2708 19221 2717
rect 19179 2668 19180 2708
rect 19220 2668 19221 2708
rect 19179 2659 19221 2668
rect 19180 2624 19220 2659
rect 19180 2573 19220 2584
rect 19276 2624 19316 3079
rect 19372 2633 19412 2718
rect 19276 2575 19316 2584
rect 19371 2624 19413 2633
rect 19371 2584 19372 2624
rect 19412 2584 19413 2624
rect 19371 2575 19413 2584
rect 18892 2500 19028 2540
rect 18892 2456 18932 2500
rect 18700 2416 18932 2456
rect 18507 2204 18549 2213
rect 18507 2164 18508 2204
rect 18548 2164 18549 2204
rect 18507 2155 18549 2164
rect 18412 1903 18452 1912
rect 18164 1072 18356 1112
rect 18124 1063 18164 1072
rect 18508 1028 18548 2155
rect 19275 1616 19317 1625
rect 19275 1576 19276 1616
rect 19316 1576 19317 1616
rect 19275 1567 19317 1576
rect 18808 1532 19176 1541
rect 18848 1492 18890 1532
rect 18930 1492 18972 1532
rect 19012 1492 19054 1532
rect 19094 1492 19136 1532
rect 18808 1483 19176 1492
rect 18699 1280 18741 1289
rect 18699 1240 18700 1280
rect 18740 1240 18741 1280
rect 18699 1231 18741 1240
rect 18316 988 18548 1028
rect 18123 944 18165 953
rect 18123 904 18124 944
rect 18164 904 18165 944
rect 18123 895 18165 904
rect 18124 80 18164 895
rect 18316 80 18356 988
rect 18507 608 18549 617
rect 18507 568 18508 608
rect 18548 568 18549 608
rect 18507 559 18549 568
rect 18508 80 18548 559
rect 18700 80 18740 1231
rect 18891 944 18933 953
rect 18891 904 18892 944
rect 18932 904 18933 944
rect 18891 895 18933 904
rect 18892 80 18932 895
rect 19083 272 19125 281
rect 19083 232 19084 272
rect 19124 232 19125 272
rect 19083 223 19125 232
rect 19084 80 19124 223
rect 19276 80 19316 1567
rect 19468 1457 19508 3340
rect 19659 3296 19701 3305
rect 19659 3256 19660 3296
rect 19700 3256 19701 3296
rect 19659 3247 19701 3256
rect 19563 2708 19605 2717
rect 19563 2668 19564 2708
rect 19604 2668 19605 2708
rect 19563 2659 19605 2668
rect 19467 1448 19509 1457
rect 19467 1408 19468 1448
rect 19508 1408 19509 1448
rect 19467 1399 19509 1408
rect 19467 1280 19509 1289
rect 19467 1240 19468 1280
rect 19508 1240 19509 1280
rect 19467 1231 19509 1240
rect 19564 1280 19604 2659
rect 19660 2624 19700 3247
rect 19852 3044 19892 3508
rect 20044 3464 20084 3508
rect 20044 3415 20084 3424
rect 19756 3004 19892 3044
rect 19948 3380 19988 3389
rect 19756 2633 19796 3004
rect 19660 2575 19700 2584
rect 19755 2624 19797 2633
rect 19755 2584 19756 2624
rect 19796 2584 19797 2624
rect 19755 2575 19797 2584
rect 19756 2120 19796 2575
rect 19852 2549 19892 2634
rect 19948 2624 19988 3340
rect 19948 2575 19988 2584
rect 19851 2540 19893 2549
rect 19851 2500 19852 2540
rect 19892 2500 19893 2540
rect 19851 2491 19893 2500
rect 20048 2288 20416 2297
rect 20088 2248 20130 2288
rect 20170 2248 20212 2288
rect 20252 2248 20294 2288
rect 20334 2248 20376 2288
rect 20048 2239 20416 2248
rect 19852 2120 19892 2129
rect 19756 2080 19852 2120
rect 19852 2071 19892 2080
rect 19947 2036 19989 2045
rect 19947 1996 19948 2036
rect 19988 1996 19989 2036
rect 19947 1987 19989 1996
rect 19564 1231 19604 1240
rect 19660 1952 19700 1961
rect 19372 1112 19412 1123
rect 19372 1037 19412 1072
rect 19371 1028 19413 1037
rect 19371 988 19372 1028
rect 19412 988 19413 1028
rect 19371 979 19413 988
rect 19468 80 19508 1231
rect 19660 1037 19700 1912
rect 19948 1457 19988 1987
rect 19947 1448 19989 1457
rect 19947 1408 19948 1448
rect 19988 1408 19989 1448
rect 19947 1399 19989 1408
rect 19659 1028 19701 1037
rect 19659 988 19660 1028
rect 19700 988 19701 1028
rect 19659 979 19701 988
rect 20048 776 20416 785
rect 20088 736 20130 776
rect 20170 736 20212 776
rect 20252 736 20294 776
rect 20334 736 20376 776
rect 20048 727 20416 736
rect 10676 64 10696 80
rect 10616 0 10696 64
rect 10808 0 10888 80
rect 11000 0 11080 80
rect 11192 0 11272 80
rect 11384 0 11464 80
rect 11576 0 11656 80
rect 11768 0 11848 80
rect 11960 0 12040 80
rect 12152 0 12232 80
rect 12344 0 12424 80
rect 12536 0 12616 80
rect 12728 0 12808 80
rect 12920 0 13000 80
rect 13112 0 13192 80
rect 13304 0 13384 80
rect 13496 0 13576 80
rect 13688 0 13768 80
rect 13880 0 13960 80
rect 14072 0 14152 80
rect 14264 0 14344 80
rect 14456 0 14536 80
rect 14648 0 14728 80
rect 14840 0 14920 80
rect 15032 0 15112 80
rect 15224 0 15304 80
rect 15416 0 15496 80
rect 15608 0 15688 80
rect 15800 0 15880 80
rect 15992 0 16072 80
rect 16184 0 16264 80
rect 16376 0 16456 80
rect 16568 0 16648 80
rect 16760 0 16840 80
rect 16952 0 17032 80
rect 17144 0 17224 80
rect 17336 0 17416 80
rect 17528 0 17608 80
rect 17720 0 17800 80
rect 17912 0 17992 80
rect 18104 0 18184 80
rect 18296 0 18376 80
rect 18488 0 18568 80
rect 18680 0 18760 80
rect 18872 0 18952 80
rect 19064 0 19144 80
rect 19256 0 19336 80
rect 19448 0 19528 80
<< via2 >>
rect 1420 40972 1460 41012
rect 1324 40552 1364 40592
rect 1516 40552 1556 40592
rect 844 38116 884 38156
rect 844 28204 884 28244
rect 76 26692 116 26732
rect 76 26440 116 26480
rect 172 25768 212 25808
rect 76 17872 116 17912
rect 556 19384 596 19424
rect 268 18460 308 18500
rect 172 13840 212 13880
rect 76 6028 116 6068
rect 460 17620 500 17660
rect 364 14008 404 14048
rect 364 4264 404 4304
rect 268 3256 308 3296
rect 652 18292 692 18332
rect 556 11236 596 11276
rect 1420 39544 1460 39584
rect 1324 38956 1364 38996
rect 1516 38872 1556 38912
rect 1036 38452 1076 38492
rect 1228 38116 1268 38156
rect 1036 21064 1076 21104
rect 1420 38368 1460 38408
rect 1708 42484 1748 42524
rect 1804 41224 1844 41264
rect 1708 39712 1748 39752
rect 1708 38872 1748 38912
rect 1804 38704 1844 38744
rect 1612 37864 1652 37904
rect 1516 37696 1556 37736
rect 1420 37528 1460 37568
rect 1612 37444 1652 37484
rect 1324 36772 1364 36812
rect 1324 36604 1364 36644
rect 1324 35932 1364 35972
rect 1612 37024 1652 37064
rect 1516 36940 1556 36980
rect 1804 37612 1844 37652
rect 2092 40636 2132 40676
rect 2092 39964 2132 40004
rect 1996 38620 2036 38660
rect 2092 38284 2132 38324
rect 2284 40888 2324 40928
rect 1996 37192 2036 37232
rect 1900 37024 1940 37064
rect 1900 36856 1940 36896
rect 1708 36436 1748 36476
rect 1708 36016 1748 36056
rect 1228 34336 1268 34376
rect 1420 35092 1460 35132
rect 1612 35008 1652 35048
rect 1516 34924 1556 34964
rect 1612 33916 1652 33956
rect 1420 33580 1460 33620
rect 1324 32908 1364 32948
rect 1324 31312 1364 31352
rect 1324 29800 1364 29840
rect 1228 26776 1268 26816
rect 1228 24592 1268 24632
rect 1228 23752 1268 23792
rect 1516 33160 1556 33200
rect 1516 32824 1556 32864
rect 1900 35344 1940 35384
rect 1996 35176 2036 35216
rect 1804 33916 1844 33956
rect 1900 33832 1940 33872
rect 2188 37948 2228 37988
rect 2284 37612 2324 37652
rect 2284 37024 2324 37064
rect 2188 35680 2228 35720
rect 2092 35008 2132 35048
rect 2092 34504 2132 34544
rect 1900 33160 1940 33200
rect 1708 32908 1748 32948
rect 1612 32740 1652 32780
rect 1900 32740 1940 32780
rect 1516 29800 1556 29840
rect 1804 31060 1844 31100
rect 1804 29296 1844 29336
rect 1708 27196 1748 27236
rect 1708 27028 1748 27068
rect 1516 25936 1556 25976
rect 1420 25432 1460 25472
rect 2572 42820 2612 42860
rect 2764 40720 2804 40760
rect 2668 40384 2708 40424
rect 2476 38620 2516 38660
rect 2476 38032 2516 38072
rect 2668 37612 2708 37652
rect 2572 37360 2612 37400
rect 2668 37276 2708 37316
rect 2380 36940 2420 36980
rect 2380 36688 2420 36728
rect 2764 36772 2804 36812
rect 2764 35932 2804 35972
rect 2469 35260 2509 35300
rect 2476 33916 2516 33956
rect 2476 33412 2516 33452
rect 2380 33160 2420 33200
rect 2284 32992 2324 33032
rect 3052 40804 3092 40844
rect 2956 40468 2996 40508
rect 3148 40384 3188 40424
rect 3436 41224 3476 41264
rect 4108 42232 4148 42272
rect 3916 42148 3956 42188
rect 4108 41728 4148 41768
rect 3724 40972 3764 41012
rect 3688 40804 3728 40844
rect 3770 40804 3810 40844
rect 3852 40804 3892 40844
rect 3934 40804 3974 40844
rect 4016 40804 4056 40844
rect 3532 40720 3572 40760
rect 4492 42064 4532 42104
rect 4876 42484 4916 42524
rect 5260 41896 5300 41936
rect 4928 41560 4968 41600
rect 5010 41560 5050 41600
rect 5092 41560 5132 41600
rect 5174 41560 5214 41600
rect 5256 41560 5296 41600
rect 4300 40888 4340 40928
rect 3244 40300 3284 40340
rect 3340 40216 3380 40256
rect 3340 39796 3380 39836
rect 3052 38368 3092 38408
rect 2956 38284 2996 38324
rect 3052 38032 3092 38072
rect 3148 37780 3188 37820
rect 2956 37276 2996 37316
rect 3052 35260 3092 35300
rect 2956 35092 2996 35132
rect 3052 33496 3092 33536
rect 2956 32992 2996 33032
rect 2860 32404 2900 32444
rect 2668 32152 2708 32192
rect 3340 38452 3380 38492
rect 3340 38284 3380 38324
rect 3532 40552 3572 40592
rect 3628 40468 3668 40508
rect 4012 40300 4052 40340
rect 3820 39460 3860 39500
rect 4108 39628 4148 39668
rect 4492 39628 4532 39668
rect 4396 39544 4436 39584
rect 3688 39292 3728 39332
rect 3770 39292 3810 39332
rect 3852 39292 3892 39332
rect 3934 39292 3974 39332
rect 4016 39292 4056 39332
rect 4012 39124 4052 39164
rect 3688 37780 3728 37820
rect 3770 37780 3810 37820
rect 3852 37780 3892 37820
rect 3934 37780 3974 37820
rect 4016 37780 4056 37820
rect 3916 37612 3956 37652
rect 3340 35848 3380 35888
rect 3340 34588 3380 34628
rect 4396 39376 4436 39416
rect 4204 38452 4244 38492
rect 4204 37360 4244 37400
rect 3820 36856 3860 36896
rect 3688 36268 3728 36308
rect 3770 36268 3810 36308
rect 3852 36268 3892 36308
rect 3934 36268 3974 36308
rect 4016 36268 4056 36308
rect 4012 36100 4052 36140
rect 3820 36016 3860 36056
rect 3628 35932 3668 35972
rect 4204 36772 4244 36812
rect 4492 37696 4532 37736
rect 4492 37192 4532 37232
rect 4684 40384 4724 40424
rect 5260 40972 5300 41012
rect 5356 40720 5396 40760
rect 5356 40384 5396 40424
rect 4928 40048 4968 40088
rect 5010 40048 5050 40088
rect 5092 40048 5132 40088
rect 5174 40048 5214 40088
rect 5256 40048 5296 40088
rect 5260 39880 5300 39920
rect 4972 39796 5012 39836
rect 4972 39124 5012 39164
rect 5260 38704 5300 38744
rect 5356 38620 5396 38660
rect 4928 38536 4968 38576
rect 5010 38536 5050 38576
rect 5092 38536 5132 38576
rect 5174 38536 5214 38576
rect 5256 38536 5296 38576
rect 5644 41896 5684 41936
rect 5548 40804 5588 40844
rect 5548 40300 5588 40340
rect 5548 40048 5588 40088
rect 4876 37696 4916 37736
rect 4684 37612 4724 37652
rect 5356 37780 5396 37820
rect 5740 40552 5780 40592
rect 5644 39880 5684 39920
rect 5644 39712 5684 39752
rect 6220 42568 6260 42608
rect 6220 41644 6260 41684
rect 6124 40972 6164 41012
rect 6124 40720 6164 40760
rect 5836 40384 5876 40424
rect 5932 40048 5972 40088
rect 5836 39460 5876 39500
rect 5932 38872 5972 38912
rect 5836 38620 5876 38660
rect 4876 37528 4916 37568
rect 5260 37444 5300 37484
rect 4928 37024 4968 37064
rect 5010 37024 5050 37064
rect 5092 37024 5132 37064
rect 5174 37024 5214 37064
rect 5256 37024 5296 37064
rect 4972 36856 5012 36896
rect 4300 36016 4340 36056
rect 3532 35092 3572 35132
rect 4012 35176 4052 35216
rect 4108 35008 4148 35048
rect 3628 34924 3668 34964
rect 3688 34756 3728 34796
rect 3770 34756 3810 34796
rect 3852 34756 3892 34796
rect 3934 34756 3974 34796
rect 4016 34756 4056 34796
rect 3436 34504 3476 34544
rect 3916 34420 3956 34460
rect 3340 34336 3380 34376
rect 3532 34168 3572 34208
rect 3436 34084 3476 34124
rect 3628 33916 3668 33956
rect 3148 32824 3188 32864
rect 3340 32572 3380 32612
rect 2572 31816 2612 31856
rect 2476 31648 2516 31688
rect 2188 31312 2228 31352
rect 2476 31312 2516 31352
rect 2092 31060 2132 31100
rect 2188 30892 2228 30932
rect 2380 30640 2420 30680
rect 1900 28876 1940 28916
rect 2572 30640 2612 30680
rect 2860 31816 2900 31856
rect 3052 31144 3092 31184
rect 2956 30640 2996 30680
rect 2476 30136 2516 30176
rect 2668 30136 2708 30176
rect 2284 30052 2324 30092
rect 2476 29800 2516 29840
rect 2860 30052 2900 30092
rect 4204 33664 4244 33704
rect 4204 33328 4244 33368
rect 3688 33244 3728 33284
rect 3770 33244 3810 33284
rect 3852 33244 3892 33284
rect 3934 33244 3974 33284
rect 4016 33244 4056 33284
rect 4012 33076 4052 33116
rect 3724 32572 3764 32612
rect 3532 32068 3572 32108
rect 3916 32068 3956 32108
rect 3688 31732 3728 31772
rect 3770 31732 3810 31772
rect 3852 31732 3892 31772
rect 3934 31732 3974 31772
rect 4016 31732 4056 31772
rect 3532 31648 3572 31688
rect 3436 31144 3476 31184
rect 3340 30976 3380 31016
rect 3436 30892 3476 30932
rect 3340 30136 3380 30176
rect 3345 29800 3385 29840
rect 2764 29212 2804 29252
rect 2764 28372 2804 28412
rect 1996 27616 2036 27656
rect 2188 27616 2228 27656
rect 1804 26776 1844 26816
rect 1612 25012 1652 25052
rect 1516 24592 1556 24632
rect 1612 23920 1652 23960
rect 1420 23836 1460 23876
rect 1420 23080 1460 23120
rect 1516 21988 1556 22028
rect 1900 24592 1940 24632
rect 1804 23584 1844 23624
rect 1804 21904 1844 21944
rect 1324 19384 1364 19424
rect 1420 17452 1460 17492
rect 1324 17116 1364 17156
rect 1132 16360 1172 16400
rect 1324 15520 1364 15560
rect 1324 15016 1364 15056
rect 1708 16612 1748 16652
rect 1612 14092 1652 14132
rect 1516 13924 1556 13964
rect 940 13084 980 13124
rect 1324 11824 1364 11864
rect 1420 11488 1460 11528
rect 1228 10984 1268 11024
rect 1324 10900 1364 10940
rect 1228 10144 1268 10184
rect 1324 7792 1364 7832
rect 652 7288 692 7328
rect 1324 7204 1364 7244
rect 1324 7036 1364 7076
rect 1324 4684 1364 4724
rect 1324 4264 1364 4304
rect 1708 13840 1748 13880
rect 1612 11068 1652 11108
rect 1612 10228 1652 10268
rect 1612 9724 1652 9764
rect 1516 6532 1556 6572
rect 1516 6028 1556 6068
rect 1420 3172 1460 3212
rect 1900 19384 1940 19424
rect 1900 18712 1940 18752
rect 1900 15520 1940 15560
rect 1900 10900 1940 10940
rect 1804 8800 1844 8840
rect 2188 27196 2228 27236
rect 2092 25012 2132 25052
rect 2572 27616 2612 27656
rect 2476 27112 2516 27152
rect 2668 27112 2708 27152
rect 2476 26776 2516 26816
rect 2380 24928 2420 24968
rect 3148 29632 3188 29672
rect 4492 35680 4532 35720
rect 4492 35092 4532 35132
rect 4492 34420 4532 34460
rect 4972 35848 5012 35888
rect 4780 35680 4820 35720
rect 4684 35512 4724 35552
rect 4928 35512 4968 35552
rect 5010 35512 5050 35552
rect 5092 35512 5132 35552
rect 5174 35512 5214 35552
rect 5256 35512 5296 35552
rect 4588 34252 4628 34292
rect 4780 35344 4820 35384
rect 4972 35344 5012 35384
rect 4396 34000 4436 34040
rect 4396 32320 4436 32360
rect 4300 31480 4340 31520
rect 4492 32152 4532 32192
rect 3916 30472 3956 30512
rect 4396 31060 4436 31100
rect 4108 30892 4148 30932
rect 4684 32992 4724 33032
rect 4928 34000 4968 34040
rect 5010 34000 5050 34040
rect 5092 34000 5132 34040
rect 5174 34000 5214 34040
rect 5256 34000 5296 34040
rect 5260 32824 5300 32864
rect 4928 32488 4968 32528
rect 5010 32488 5050 32528
rect 5092 32488 5132 32528
rect 5174 32488 5214 32528
rect 5256 32488 5296 32528
rect 5452 35680 5492 35720
rect 5644 35260 5684 35300
rect 5548 34924 5588 34964
rect 5740 34840 5780 34880
rect 5740 34672 5780 34712
rect 5836 34504 5876 34544
rect 6412 40552 6452 40592
rect 6316 40384 6356 40424
rect 6316 39712 6356 39752
rect 6508 40300 6548 40340
rect 6412 39040 6452 39080
rect 6412 38788 6452 38828
rect 6316 38284 6356 38324
rect 6700 40384 6740 40424
rect 6604 38368 6644 38408
rect 6124 37612 6164 37652
rect 6508 37444 6548 37484
rect 6508 36520 6548 36560
rect 6988 40468 7028 40508
rect 6988 39208 7028 39248
rect 6796 39124 6836 39164
rect 6892 38368 6932 38408
rect 6796 37024 6836 37064
rect 6700 36520 6740 36560
rect 6604 35848 6644 35888
rect 6316 35260 6356 35300
rect 6220 35176 6260 35216
rect 6124 34756 6164 34796
rect 5740 34336 5780 34376
rect 5644 34252 5684 34292
rect 5548 34000 5588 34040
rect 5644 33916 5684 33956
rect 5452 33328 5492 33368
rect 5452 32908 5492 32948
rect 5356 32236 5396 32276
rect 4972 32152 5012 32192
rect 4780 32068 4820 32108
rect 4684 31060 4724 31100
rect 3688 30220 3728 30260
rect 3770 30220 3810 30260
rect 3852 30220 3892 30260
rect 3934 30220 3974 30260
rect 4016 30220 4056 30260
rect 3628 29800 3668 29840
rect 3532 29212 3572 29252
rect 3916 29632 3956 29672
rect 3820 29380 3860 29420
rect 3340 28372 3380 28412
rect 2956 28288 2996 28328
rect 3052 27532 3092 27572
rect 2860 27196 2900 27236
rect 3340 28120 3380 28160
rect 3688 28708 3728 28748
rect 3770 28708 3810 28748
rect 3852 28708 3892 28748
rect 3934 28708 3974 28748
rect 4016 28708 4056 28748
rect 3628 28288 3668 28328
rect 4396 30388 4436 30428
rect 4204 29548 4244 29588
rect 3148 26860 3188 26900
rect 2860 26776 2900 26816
rect 2860 26440 2900 26480
rect 3436 27700 3476 27740
rect 3532 27616 3572 27656
rect 4012 28120 4052 28160
rect 3916 27700 3956 27740
rect 3688 27196 3728 27236
rect 3770 27196 3810 27236
rect 3852 27196 3892 27236
rect 3934 27196 3974 27236
rect 4016 27196 4056 27236
rect 3340 26188 3380 26228
rect 3436 26104 3476 26144
rect 3148 25516 3188 25556
rect 3340 25516 3380 25556
rect 3052 25348 3092 25388
rect 2764 24760 2804 24800
rect 3148 24760 3188 24800
rect 3436 24760 3476 24800
rect 2380 23920 2420 23960
rect 2668 24340 2708 24380
rect 2956 24592 2996 24632
rect 2956 24340 2996 24380
rect 2956 23836 2996 23876
rect 3340 23837 3380 23876
rect 3340 23836 3380 23837
rect 2284 23584 2324 23624
rect 2188 21652 2228 21692
rect 2092 19552 2132 19592
rect 2092 19216 2132 19256
rect 2188 18712 2228 18752
rect 2188 18544 2228 18584
rect 2092 14092 2132 14132
rect 2092 13840 2132 13880
rect 2284 17536 2324 17576
rect 2284 17116 2324 17156
rect 2284 15352 2324 15392
rect 2764 23752 2804 23792
rect 3052 23752 3092 23792
rect 3628 26188 3668 26228
rect 3916 26020 3956 26060
rect 3820 25852 3860 25892
rect 4108 26440 4148 26480
rect 4492 26776 4532 26816
rect 4300 26188 4340 26228
rect 3688 25684 3728 25724
rect 3770 25684 3810 25724
rect 3852 25684 3892 25724
rect 3934 25684 3974 25724
rect 4016 25684 4056 25724
rect 3724 25348 3764 25388
rect 3820 25264 3860 25304
rect 3688 24172 3728 24212
rect 3770 24172 3810 24212
rect 3852 24172 3892 24212
rect 3934 24172 3974 24212
rect 4016 24172 4056 24212
rect 4396 25852 4436 25892
rect 4204 25768 4244 25808
rect 2476 23500 2516 23540
rect 3148 23584 3188 23624
rect 3532 23584 3572 23624
rect 3340 23332 3380 23372
rect 2476 19216 2516 19256
rect 2860 23164 2900 23204
rect 3244 23164 3284 23204
rect 3532 23164 3572 23204
rect 2764 22240 2804 22280
rect 2860 22156 2900 22196
rect 2956 22072 2996 22112
rect 3052 20644 3092 20684
rect 3148 20644 3188 20684
rect 2668 19468 2708 19508
rect 2764 19216 2804 19256
rect 2572 18544 2612 18584
rect 2572 17452 2612 17492
rect 3340 20056 3380 20096
rect 3244 19972 3284 20012
rect 2956 19888 2996 19928
rect 3244 19720 3284 19760
rect 3340 19552 3380 19592
rect 3244 18880 3284 18920
rect 3820 23416 3860 23456
rect 3724 23164 3764 23204
rect 4012 23836 4052 23876
rect 4108 23584 4148 23624
rect 3724 22996 3764 23036
rect 3628 22912 3668 22952
rect 4108 22828 4148 22868
rect 3688 22660 3728 22700
rect 3770 22660 3810 22700
rect 3852 22660 3892 22700
rect 3934 22660 3974 22700
rect 4016 22660 4056 22700
rect 3628 21568 3668 21608
rect 4012 21568 4052 21608
rect 3688 21148 3728 21188
rect 3770 21148 3810 21188
rect 3852 21148 3892 21188
rect 3934 21148 3974 21188
rect 4016 21148 4056 21188
rect 6028 34336 6068 34376
rect 5932 34084 5972 34124
rect 5932 33916 5972 33956
rect 5644 32992 5684 33032
rect 5644 32824 5684 32864
rect 5548 31480 5588 31520
rect 4928 30976 4968 31016
rect 5010 30976 5050 31016
rect 5092 30976 5132 31016
rect 5174 30976 5214 31016
rect 5256 30976 5296 31016
rect 4876 30808 4916 30848
rect 4780 30640 4820 30680
rect 4972 30640 5012 30680
rect 4972 30388 5012 30428
rect 5452 31144 5492 31184
rect 4928 29464 4968 29504
rect 5010 29464 5050 29504
rect 5092 29464 5132 29504
rect 5174 29464 5214 29504
rect 5256 29464 5296 29504
rect 4780 29380 4820 29420
rect 5356 29380 5396 29420
rect 4684 28540 4724 28580
rect 5068 29212 5108 29252
rect 5740 32656 5780 32696
rect 5644 30472 5684 30512
rect 5644 30220 5684 30260
rect 5548 29044 5588 29084
rect 5452 28960 5492 29000
rect 6028 33664 6068 33704
rect 6220 33244 6260 33284
rect 6124 32740 6164 32780
rect 6028 31984 6068 32024
rect 6028 31480 6068 31520
rect 5932 31312 5972 31352
rect 6220 32320 6260 32360
rect 6124 31312 6164 31352
rect 6028 31144 6068 31184
rect 5740 30052 5780 30092
rect 5356 28372 5396 28412
rect 5356 28204 5396 28244
rect 4928 27952 4968 27992
rect 5010 27952 5050 27992
rect 5092 27952 5132 27992
rect 5174 27952 5214 27992
rect 5256 27952 5296 27992
rect 4780 27028 4820 27068
rect 4780 26776 4820 26816
rect 4684 26440 4724 26480
rect 4928 26440 4968 26480
rect 5010 26440 5050 26480
rect 5092 26440 5132 26480
rect 5174 26440 5214 26480
rect 5256 26440 5296 26480
rect 5548 27028 5588 27068
rect 4876 26188 4916 26228
rect 5068 26188 5108 26228
rect 5452 26020 5492 26060
rect 5452 25348 5492 25388
rect 4928 24928 4968 24968
rect 5010 24928 5050 24968
rect 5092 24928 5132 24968
rect 5174 24928 5214 24968
rect 5256 24928 5296 24968
rect 5740 26776 5780 26816
rect 5932 28876 5972 28916
rect 5932 28288 5972 28328
rect 6412 34756 6452 34796
rect 6412 34336 6452 34376
rect 6508 33328 6548 33368
rect 7084 38704 7124 38744
rect 7084 38116 7124 38156
rect 7084 37276 7124 37316
rect 7372 41728 7412 41768
rect 7756 41644 7796 41684
rect 7564 41224 7604 41264
rect 7276 40552 7316 40592
rect 7660 40384 7700 40424
rect 8044 41140 8084 41180
rect 7948 40720 7988 40760
rect 7756 40132 7796 40172
rect 7660 40048 7700 40088
rect 7372 39460 7412 39500
rect 7756 38872 7796 38912
rect 8524 40552 8564 40592
rect 8236 40048 8276 40088
rect 8428 39460 8468 39500
rect 8044 39376 8084 39416
rect 8140 39040 8180 39080
rect 8332 39040 8372 39080
rect 7948 38872 7988 38912
rect 7276 38200 7316 38240
rect 7276 37192 7316 37232
rect 7372 36856 7412 36896
rect 7276 36772 7316 36812
rect 6988 36688 7028 36728
rect 6892 36520 6932 36560
rect 7276 36520 7316 36560
rect 6892 34084 6932 34124
rect 6796 33664 6836 33704
rect 7276 35764 7316 35804
rect 7852 38536 7892 38576
rect 8044 37612 8084 37652
rect 7660 37276 7700 37316
rect 7564 36016 7604 36056
rect 7660 35680 7700 35720
rect 7564 35512 7604 35552
rect 7468 35428 7508 35468
rect 7948 37360 7988 37400
rect 7852 37276 7892 37316
rect 8428 38872 8468 38912
rect 8332 38452 8372 38492
rect 8332 37612 8372 37652
rect 8716 40636 8756 40676
rect 8620 40048 8660 40088
rect 8620 38368 8660 38408
rect 8524 37780 8564 37820
rect 8908 38956 8948 38996
rect 9196 40216 9236 40256
rect 8812 38032 8852 38072
rect 9100 38872 9140 38912
rect 8140 37360 8180 37400
rect 7948 35848 7988 35888
rect 8044 35680 8084 35720
rect 7852 35596 7892 35636
rect 7372 35176 7412 35216
rect 7276 35008 7316 35048
rect 7468 35008 7508 35048
rect 7276 34756 7316 34796
rect 7756 34924 7796 34964
rect 7756 34588 7796 34628
rect 8044 34336 8084 34376
rect 7564 34168 7604 34208
rect 7276 33244 7316 33284
rect 6892 32908 6932 32948
rect 8620 37276 8660 37316
rect 8236 36772 8276 36812
rect 8236 35764 8276 35804
rect 8236 35512 8276 35552
rect 8620 36856 8660 36896
rect 9388 41224 9428 41264
rect 9388 39460 9428 39500
rect 9388 38704 9428 38744
rect 9292 38284 9332 38324
rect 9388 38032 9428 38072
rect 8908 37024 8948 37064
rect 8524 36772 8564 36812
rect 7756 33580 7796 33620
rect 7756 32992 7796 33032
rect 7276 32908 7316 32948
rect 7084 32824 7124 32864
rect 7372 32740 7412 32780
rect 6796 32488 6836 32528
rect 6508 32152 6548 32192
rect 6316 31228 6356 31268
rect 6316 30892 6356 30932
rect 6892 32236 6932 32276
rect 6700 32152 6740 32192
rect 6604 31564 6644 31604
rect 6604 31396 6644 31436
rect 7180 32488 7220 32528
rect 7084 32152 7124 32192
rect 6892 31480 6932 31520
rect 7084 31480 7124 31520
rect 6892 31060 6932 31100
rect 6796 30808 6836 30848
rect 7852 32824 7892 32864
rect 8044 32992 8084 33032
rect 7564 31480 7604 31520
rect 8428 34420 8468 34460
rect 8236 33664 8276 33704
rect 8332 33580 8372 33620
rect 8236 32740 8276 32780
rect 8140 32320 8180 32360
rect 8140 32152 8180 32192
rect 8428 32320 8468 32360
rect 7948 31648 7988 31688
rect 7756 31480 7796 31520
rect 8044 31480 8084 31520
rect 7660 31396 7700 31436
rect 8236 31396 8276 31436
rect 7180 31144 7220 31184
rect 6220 30220 6260 30260
rect 6220 30052 6260 30092
rect 6124 29128 6164 29168
rect 6316 29968 6356 30008
rect 6412 29800 6452 29840
rect 6316 29716 6356 29756
rect 6220 27784 6260 27824
rect 5932 27028 5972 27068
rect 5932 26692 5972 26732
rect 5836 26608 5876 26648
rect 5644 25264 5684 25304
rect 5452 24844 5492 24884
rect 4876 24004 4916 24044
rect 4300 23668 4340 23708
rect 4492 23752 4532 23792
rect 4396 23332 4436 23372
rect 4588 23584 4628 23624
rect 4492 23248 4532 23288
rect 5740 24004 5780 24044
rect 5164 23752 5204 23792
rect 5068 23668 5108 23708
rect 5644 23752 5684 23792
rect 4972 23584 5012 23624
rect 4928 23416 4968 23456
rect 5010 23416 5050 23456
rect 5092 23416 5132 23456
rect 5174 23416 5214 23456
rect 5256 23416 5296 23456
rect 5452 23584 5492 23624
rect 5644 23416 5684 23456
rect 4780 23248 4820 23288
rect 4492 22912 4532 22952
rect 4300 22240 4340 22280
rect 4780 22912 4820 22952
rect 4972 22240 5012 22280
rect 5356 23080 5396 23120
rect 5164 22912 5204 22952
rect 5548 22912 5588 22952
rect 5452 22240 5492 22280
rect 5356 22156 5396 22196
rect 4928 21904 4968 21944
rect 5010 21904 5050 21944
rect 5092 21904 5132 21944
rect 5174 21904 5214 21944
rect 5256 21904 5296 21944
rect 5260 21736 5300 21776
rect 4684 21484 4724 21524
rect 4108 20896 4148 20936
rect 3628 20644 3668 20684
rect 4300 20980 4340 21020
rect 3532 20224 3572 20264
rect 4108 19972 4148 20012
rect 3916 19888 3956 19928
rect 3820 19804 3860 19844
rect 3688 19636 3728 19676
rect 3770 19636 3810 19676
rect 3852 19636 3892 19676
rect 3934 19636 3974 19676
rect 4016 19636 4056 19676
rect 3820 19300 3860 19340
rect 3916 19216 3956 19256
rect 3340 18628 3380 18668
rect 3244 18544 3284 18584
rect 2860 17368 2900 17408
rect 2476 17032 2516 17072
rect 2860 16948 2900 16988
rect 2476 15436 2516 15476
rect 2764 16192 2804 16232
rect 2860 16024 2900 16064
rect 2860 15268 2900 15308
rect 2380 15016 2420 15056
rect 3148 18208 3188 18248
rect 3052 17368 3092 17408
rect 3052 17200 3092 17240
rect 3052 16780 3092 16820
rect 3052 16024 3092 16064
rect 3052 15520 3092 15560
rect 3340 17200 3380 17240
rect 3340 16948 3380 16988
rect 3340 16444 3380 16484
rect 4108 18796 4148 18836
rect 4204 18712 4244 18752
rect 3532 18208 3572 18248
rect 3688 18124 3728 18164
rect 3770 18124 3810 18164
rect 3852 18124 3892 18164
rect 3934 18124 3974 18164
rect 4016 18124 4056 18164
rect 3532 17116 3572 17156
rect 3820 17032 3860 17072
rect 3532 16612 3572 16652
rect 3688 16612 3728 16652
rect 3770 16612 3810 16652
rect 3852 16612 3892 16652
rect 3934 16612 3974 16652
rect 4016 16612 4056 16652
rect 3628 16444 3668 16484
rect 5452 21316 5492 21356
rect 5644 22744 5684 22784
rect 5644 22576 5684 22616
rect 5836 23752 5876 23792
rect 6220 27532 6260 27572
rect 6124 26692 6164 26732
rect 6124 26524 6164 26564
rect 7372 30640 7412 30680
rect 8332 31144 8372 31184
rect 7372 29968 7412 30008
rect 7852 29968 7892 30008
rect 7468 29884 7508 29924
rect 7276 29800 7316 29840
rect 6700 28372 6740 28412
rect 6508 26860 6548 26900
rect 6316 26440 6356 26480
rect 6220 26104 6260 26144
rect 6124 25096 6164 25136
rect 6028 23668 6068 23708
rect 6028 23416 6068 23456
rect 6220 24928 6260 24968
rect 6892 29212 6932 29252
rect 6796 27532 6836 27572
rect 6988 29128 7028 29168
rect 7756 28372 7796 28412
rect 6988 27616 7028 27656
rect 6892 27448 6932 27488
rect 6700 26776 6740 26816
rect 6700 26524 6740 26564
rect 7084 27028 7124 27068
rect 7660 27616 7700 27656
rect 7276 27448 7316 27488
rect 7468 27364 7508 27404
rect 7372 26524 7412 26564
rect 6796 26104 6836 26144
rect 7084 26104 7124 26144
rect 6604 25936 6644 25976
rect 6796 25852 6836 25892
rect 6700 24592 6740 24632
rect 6508 23752 6548 23792
rect 6124 23248 6164 23288
rect 5740 21736 5780 21776
rect 5644 21652 5684 21692
rect 5740 21568 5780 21608
rect 5548 20980 5588 21020
rect 4684 20812 4724 20852
rect 5068 20728 5108 20768
rect 4684 20308 4724 20348
rect 4396 20056 4436 20096
rect 4588 19972 4628 20012
rect 4492 19888 4532 19928
rect 4396 19300 4436 19340
rect 4492 19216 4532 19256
rect 4928 20392 4968 20432
rect 5010 20392 5050 20432
rect 5092 20392 5132 20432
rect 5174 20392 5214 20432
rect 5256 20392 5296 20432
rect 5356 20056 5396 20096
rect 5260 19888 5300 19928
rect 5356 19216 5396 19256
rect 4928 18880 4968 18920
rect 5010 18880 5050 18920
rect 5092 18880 5132 18920
rect 5174 18880 5214 18920
rect 5256 18880 5296 18920
rect 5164 18712 5204 18752
rect 5548 18460 5588 18500
rect 5260 17872 5300 17912
rect 4928 17368 4968 17408
rect 5010 17368 5050 17408
rect 5092 17368 5132 17408
rect 5174 17368 5214 17408
rect 5256 17368 5296 17408
rect 3820 16444 3860 16484
rect 3436 16360 3476 16400
rect 3340 16192 3380 16232
rect 2956 15100 2996 15140
rect 3148 15352 3188 15392
rect 3244 14848 3284 14888
rect 2668 14512 2708 14552
rect 2764 14344 2804 14384
rect 3148 14596 3188 14636
rect 3244 14344 3284 14384
rect 3916 16276 3956 16316
rect 3820 15520 3860 15560
rect 4492 16360 4532 16400
rect 4396 16024 4436 16064
rect 4300 15772 4340 15812
rect 4204 15688 4244 15728
rect 4108 15520 4148 15560
rect 4588 15772 4628 15812
rect 3436 15436 3476 15476
rect 4492 15352 4532 15392
rect 3628 15268 3668 15308
rect 4108 15268 4148 15308
rect 3688 15100 3728 15140
rect 3770 15100 3810 15140
rect 3852 15100 3892 15140
rect 3934 15100 3974 15140
rect 4016 15100 4056 15140
rect 4108 14764 4148 14804
rect 3820 14596 3860 14636
rect 3532 14512 3572 14552
rect 3532 14344 3572 14384
rect 2956 14176 2996 14216
rect 3340 14176 3380 14216
rect 2860 13840 2900 13880
rect 2572 13084 2612 13124
rect 2284 12580 2324 12620
rect 2476 12496 2516 12536
rect 2764 12580 2804 12620
rect 2284 12328 2324 12368
rect 2188 10984 2228 11024
rect 2476 11656 2516 11696
rect 2668 11236 2708 11276
rect 2572 10732 2612 10772
rect 2092 10144 2132 10184
rect 2476 10228 2516 10268
rect 2284 10144 2324 10184
rect 2188 9556 2228 9596
rect 1996 7960 2036 8000
rect 1996 7792 2036 7832
rect 1804 6952 1844 6992
rect 1900 5440 1940 5480
rect 2188 7960 2228 8000
rect 2092 7456 2132 7496
rect 2092 5944 2132 5984
rect 1996 4600 2036 4640
rect 1996 3676 2036 3716
rect 1612 3088 1652 3128
rect 460 2752 500 2792
rect 1612 2584 1652 2624
rect 1708 2500 1748 2540
rect 1324 1912 1364 1952
rect 1804 1660 1844 1700
rect 1804 1492 1844 1532
rect 2476 9388 2516 9428
rect 2668 10564 2708 10604
rect 2860 10060 2900 10100
rect 3244 13756 3284 13796
rect 3340 13672 3380 13712
rect 3916 14176 3956 14216
rect 4396 14512 4436 14552
rect 4108 13924 4148 13964
rect 3688 13588 3728 13628
rect 3770 13588 3810 13628
rect 3852 13588 3892 13628
rect 3934 13588 3974 13628
rect 4016 13588 4056 13628
rect 3724 13168 3764 13208
rect 3532 12496 3572 12536
rect 4108 13168 4148 13208
rect 4396 13840 4436 13880
rect 3916 12496 3956 12536
rect 3820 12244 3860 12284
rect 3244 12076 3284 12116
rect 3688 12076 3728 12116
rect 3770 12076 3810 12116
rect 3852 12076 3892 12116
rect 3934 12076 3974 12116
rect 4016 12076 4056 12116
rect 3052 11152 3092 11192
rect 3052 10396 3092 10436
rect 2956 9472 2996 9512
rect 2764 9388 2804 9428
rect 3724 11152 3764 11192
rect 3724 10816 3764 10856
rect 3820 10732 3860 10772
rect 3688 10564 3728 10604
rect 3770 10564 3810 10604
rect 3852 10564 3892 10604
rect 3934 10564 3974 10604
rect 4016 10564 4056 10604
rect 4588 14176 4628 14216
rect 4492 12160 4532 12200
rect 4780 17032 4820 17072
rect 4780 16780 4820 16820
rect 5260 16360 5300 16400
rect 5164 16192 5204 16232
rect 5068 16108 5108 16148
rect 4928 15856 4968 15896
rect 5010 15856 5050 15896
rect 5092 15856 5132 15896
rect 5174 15856 5214 15896
rect 5256 15856 5296 15896
rect 4780 15520 4820 15560
rect 4684 14092 4724 14132
rect 4588 11320 4628 11360
rect 4300 11236 4340 11276
rect 4492 10984 4532 11024
rect 3436 10060 3476 10100
rect 3532 9976 3572 10016
rect 4108 10144 4148 10184
rect 4396 10816 4436 10856
rect 4492 10732 4532 10772
rect 4396 10396 4436 10436
rect 3340 9472 3380 9512
rect 3148 9220 3188 9260
rect 2668 8884 2708 8924
rect 3052 8800 3092 8840
rect 3052 8548 3092 8588
rect 2956 8464 2996 8504
rect 2668 7960 2708 8000
rect 2572 7540 2612 7580
rect 2572 7372 2612 7412
rect 2860 7876 2900 7916
rect 2764 7708 2804 7748
rect 2476 7120 2516 7160
rect 2380 6448 2420 6488
rect 2668 6616 2708 6656
rect 3532 9472 3572 9512
rect 3436 9388 3476 9428
rect 4108 9388 4148 9428
rect 3688 9052 3728 9092
rect 3770 9052 3810 9092
rect 3852 9052 3892 9092
rect 3934 9052 3974 9092
rect 4016 9052 4056 9092
rect 3532 8884 3572 8924
rect 3820 8884 3860 8924
rect 3340 8548 3380 8588
rect 3436 8128 3476 8168
rect 3052 7120 3092 7160
rect 3148 6448 3188 6488
rect 2572 6280 2612 6320
rect 2284 5020 2324 5060
rect 3052 6280 3092 6320
rect 3244 6280 3284 6320
rect 2764 5608 2804 5648
rect 2476 5440 2516 5480
rect 2188 4768 2228 4808
rect 2668 4768 2708 4808
rect 2188 3172 2228 3212
rect 2092 1492 2132 1532
rect 1900 232 1940 272
rect 1996 64 2036 104
rect 2284 3088 2324 3128
rect 2668 3928 2708 3968
rect 2668 2836 2708 2876
rect 2855 4936 2860 4976
rect 2860 4936 2895 4976
rect 2956 4936 2996 4976
rect 2860 4768 2900 4808
rect 2860 3928 2900 3968
rect 2956 3844 2996 3884
rect 2956 1828 2996 1868
rect 3148 5776 3188 5816
rect 3148 5440 3188 5480
rect 3148 4768 3188 4808
rect 3436 7624 3476 7664
rect 3436 7120 3476 7160
rect 4684 10732 4724 10772
rect 4588 9472 4628 9512
rect 4684 9388 4724 9428
rect 4492 9136 4532 9176
rect 4204 8716 4244 8756
rect 4876 15352 4916 15392
rect 4928 14344 4968 14384
rect 5010 14344 5050 14384
rect 5092 14344 5132 14384
rect 5174 14344 5214 14384
rect 5256 14344 5296 14384
rect 4928 12832 4968 12872
rect 5010 12832 5050 12872
rect 5092 12832 5132 12872
rect 5174 12832 5214 12872
rect 5256 12832 5296 12872
rect 5452 16276 5492 16316
rect 6700 23332 6740 23372
rect 6316 23164 6356 23204
rect 6604 23164 6644 23204
rect 5932 22996 5972 23036
rect 6316 22912 6356 22952
rect 6028 22828 6068 22868
rect 6220 22324 6260 22364
rect 6220 22156 6260 22196
rect 6124 21316 6164 21356
rect 5932 20644 5972 20684
rect 6028 18292 6068 18332
rect 5932 18208 5972 18248
rect 6028 17872 6068 17912
rect 5548 16192 5588 16232
rect 5740 15436 5780 15476
rect 5644 14848 5684 14888
rect 5740 14596 5780 14636
rect 5548 13840 5588 13880
rect 5644 13168 5684 13208
rect 5452 12832 5492 12872
rect 5164 12244 5204 12284
rect 6028 14260 6068 14300
rect 6028 14008 6068 14048
rect 5836 13840 5876 13880
rect 5452 11992 5492 12032
rect 4928 11320 4968 11360
rect 5010 11320 5050 11360
rect 5092 11320 5132 11360
rect 5174 11320 5214 11360
rect 5256 11320 5296 11360
rect 4972 11152 5012 11192
rect 4876 10984 4916 11024
rect 5164 10984 5204 11024
rect 5068 10816 5108 10856
rect 6220 16108 6260 16148
rect 6220 15604 6260 15644
rect 6220 13840 6260 13880
rect 5932 12496 5972 12536
rect 5836 11824 5876 11864
rect 5932 11740 5972 11780
rect 4928 9808 4968 9848
rect 5010 9808 5050 9848
rect 5092 9808 5132 9848
rect 5174 9808 5214 9848
rect 5256 9808 5296 9848
rect 5356 9808 5396 9848
rect 5356 9556 5396 9596
rect 5548 9556 5588 9596
rect 5356 9136 5396 9176
rect 4108 8632 4148 8672
rect 4492 8632 4532 8672
rect 4012 8548 4052 8588
rect 4204 8464 4244 8504
rect 4396 8128 4436 8168
rect 4204 7876 4244 7916
rect 3724 7792 3764 7832
rect 4108 7708 4148 7748
rect 3688 7540 3728 7580
rect 3770 7540 3810 7580
rect 3852 7540 3892 7580
rect 3934 7540 3974 7580
rect 4016 7540 4056 7580
rect 3532 6616 3572 6656
rect 3436 6532 3476 6572
rect 4396 7456 4436 7496
rect 4300 7204 4340 7244
rect 4108 6196 4148 6236
rect 4300 6196 4340 6236
rect 3688 6028 3728 6068
rect 3770 6028 3810 6068
rect 3852 6028 3892 6068
rect 3934 6028 3974 6068
rect 4016 6028 4056 6068
rect 3340 5860 3380 5900
rect 3724 5860 3764 5900
rect 3628 5692 3668 5732
rect 4108 5524 4148 5564
rect 4684 7960 4724 8000
rect 5356 8632 5396 8672
rect 4876 8464 4916 8504
rect 4928 8296 4968 8336
rect 5010 8296 5050 8336
rect 5092 8296 5132 8336
rect 5174 8296 5214 8336
rect 5256 8296 5296 8336
rect 4780 7540 4820 7580
rect 4588 7372 4628 7412
rect 4780 6952 4820 6992
rect 4928 6784 4968 6824
rect 5010 6784 5050 6824
rect 5092 6784 5132 6824
rect 5174 6784 5214 6824
rect 5256 6784 5296 6824
rect 4588 6280 4628 6320
rect 4684 6196 4724 6236
rect 5260 6364 5300 6404
rect 4396 5356 4436 5396
rect 4300 5104 4340 5144
rect 3340 5020 3380 5060
rect 4204 5020 4244 5060
rect 3244 4180 3284 4220
rect 3148 4096 3188 4136
rect 3148 3592 3188 3632
rect 4780 5608 4820 5648
rect 5164 5608 5204 5648
rect 4684 5356 4724 5396
rect 4492 4936 4532 4976
rect 4396 4852 4436 4892
rect 4108 4768 4148 4808
rect 3688 4516 3728 4556
rect 3770 4516 3810 4556
rect 3852 4516 3892 4556
rect 3934 4516 3974 4556
rect 4016 4516 4056 4556
rect 3532 4264 3572 4304
rect 3436 2836 3476 2876
rect 4108 4180 4148 4220
rect 3628 3424 3668 3464
rect 3724 3340 3764 3380
rect 3688 3004 3728 3044
rect 3770 3004 3810 3044
rect 3852 3004 3892 3044
rect 3934 3004 3974 3044
rect 4016 3004 4056 3044
rect 3916 2668 3956 2708
rect 3148 1660 3188 1700
rect 3340 1576 3380 1616
rect 3532 1744 3572 1784
rect 4108 1744 4148 1784
rect 3688 1492 3728 1532
rect 3770 1492 3810 1532
rect 3852 1492 3892 1532
rect 3934 1492 3974 1532
rect 4016 1492 4056 1532
rect 2572 736 2612 776
rect 2764 904 2804 944
rect 2668 652 2708 692
rect 3340 1240 3380 1280
rect 3724 1240 3764 1280
rect 3532 988 3572 1028
rect 3916 1156 3956 1196
rect 4588 4180 4628 4220
rect 4492 4096 4532 4136
rect 4928 5272 4968 5312
rect 5010 5272 5050 5312
rect 5092 5272 5132 5312
rect 5174 5272 5214 5312
rect 5256 5272 5296 5312
rect 4780 5020 4820 5060
rect 5452 8464 5492 8504
rect 5548 8044 5588 8084
rect 5452 6196 5492 6236
rect 5260 4600 5300 4640
rect 4972 4264 5012 4304
rect 4780 4012 4820 4052
rect 5452 4264 5492 4304
rect 5356 4012 5396 4052
rect 5260 3928 5300 3968
rect 5356 3844 5396 3884
rect 4928 3760 4968 3800
rect 5010 3760 5050 3800
rect 5092 3760 5132 3800
rect 5174 3760 5214 3800
rect 5256 3760 5296 3800
rect 4684 3592 4724 3632
rect 5068 3596 5108 3632
rect 5068 3592 5108 3596
rect 4588 3508 4628 3548
rect 4876 3256 4916 3296
rect 4972 2836 5012 2876
rect 5260 2836 5300 2876
rect 5740 9640 5780 9680
rect 5932 9136 5972 9176
rect 6220 12832 6260 12872
rect 6124 12496 6164 12536
rect 6124 12244 6164 12284
rect 5644 7708 5684 7748
rect 5644 6448 5684 6488
rect 4928 2248 4968 2288
rect 5010 2248 5050 2288
rect 5092 2248 5132 2288
rect 5174 2248 5214 2288
rect 5256 2248 5296 2288
rect 4780 2080 4820 2120
rect 4780 1912 4820 1952
rect 4972 1912 5012 1952
rect 5644 1996 5684 2036
rect 5356 1744 5396 1784
rect 4972 1492 5012 1532
rect 4876 1408 4916 1448
rect 4204 1072 4244 1112
rect 4780 1072 4820 1112
rect 4492 988 4532 1028
rect 4108 904 4148 944
rect 4300 568 4340 608
rect 5452 1240 5492 1280
rect 5068 1072 5108 1112
rect 4588 904 4628 944
rect 5356 904 5396 944
rect 4928 736 4968 776
rect 5010 736 5050 776
rect 5092 736 5132 776
rect 5174 736 5214 776
rect 5256 736 5296 776
rect 4876 568 4916 608
rect 5260 568 5300 608
rect 5068 484 5108 524
rect 5644 1156 5684 1196
rect 7276 26440 7316 26480
rect 7180 25264 7220 25304
rect 7180 24592 7220 24632
rect 6892 23752 6932 23792
rect 7564 27028 7604 27068
rect 7660 26440 7700 26480
rect 7564 25264 7604 25304
rect 7084 23584 7124 23624
rect 6892 23416 6932 23456
rect 6988 23164 7028 23204
rect 6892 22660 6932 22700
rect 7084 22996 7124 23036
rect 7180 22828 7220 22868
rect 7084 22660 7124 22700
rect 7276 22240 7316 22280
rect 6892 21736 6932 21776
rect 7084 21736 7124 21776
rect 6796 20812 6836 20852
rect 6700 20728 6740 20768
rect 6604 20644 6644 20684
rect 7180 20812 7220 20852
rect 6796 20056 6836 20096
rect 6988 19720 7028 19760
rect 6988 19468 7028 19508
rect 6412 19216 6452 19256
rect 7564 23584 7604 23624
rect 7468 22912 7508 22952
rect 7660 23080 7700 23120
rect 8044 29884 8084 29924
rect 7948 28540 7988 28580
rect 8428 29968 8468 30008
rect 8236 29800 8276 29840
rect 8812 36688 8852 36728
rect 8716 36520 8756 36560
rect 8716 36016 8756 36056
rect 8620 33664 8660 33704
rect 8620 32152 8660 32192
rect 8908 36436 8948 36476
rect 9868 41560 9908 41600
rect 10060 41560 10100 41600
rect 9964 41224 10004 41264
rect 9772 40468 9812 40508
rect 9772 40300 9812 40340
rect 9676 40216 9716 40256
rect 9580 39880 9620 39920
rect 10060 40804 10100 40844
rect 9580 38200 9620 38240
rect 10252 40636 10292 40676
rect 10252 40216 10292 40256
rect 10156 40132 10196 40172
rect 10444 40804 10484 40844
rect 10444 40636 10484 40676
rect 10924 40636 10964 40676
rect 10540 40468 10580 40508
rect 10732 40384 10772 40424
rect 11788 42568 11828 42608
rect 11404 41560 11444 41600
rect 11596 41560 11636 41600
rect 11308 41392 11348 41432
rect 11596 41224 11636 41264
rect 11404 41140 11444 41180
rect 10732 40132 10772 40172
rect 11020 40132 11060 40172
rect 10252 39544 10292 39584
rect 10060 38788 10100 38828
rect 10060 38200 10100 38240
rect 9100 35512 9140 35552
rect 9772 37360 9812 37400
rect 9004 35260 9044 35300
rect 9292 35260 9332 35300
rect 8908 35092 8948 35132
rect 9484 36436 9524 36476
rect 9580 35428 9620 35468
rect 9004 35008 9044 35048
rect 8908 34672 8948 34712
rect 8908 34168 8948 34208
rect 8716 31312 8756 31352
rect 8620 31228 8660 31268
rect 8716 31060 8756 31100
rect 8812 30892 8852 30932
rect 8236 28288 8276 28328
rect 8044 27364 8084 27404
rect 7852 26440 7892 26480
rect 7852 25096 7892 25136
rect 7852 24592 7892 24632
rect 7852 24340 7892 24380
rect 8140 25936 8180 25976
rect 8140 25264 8180 25304
rect 8332 26440 8372 26480
rect 8332 25936 8372 25976
rect 8236 24760 8276 24800
rect 8236 24592 8276 24632
rect 7756 22576 7796 22616
rect 7756 22324 7796 22364
rect 7660 22240 7700 22280
rect 8140 23584 8180 23624
rect 8332 23584 8372 23624
rect 8716 28792 8756 28832
rect 8716 27700 8756 27740
rect 9004 29128 9044 29168
rect 8908 28624 8948 28664
rect 8908 28456 8948 28496
rect 9772 36688 9812 36728
rect 9772 36520 9812 36560
rect 10060 37360 10100 37400
rect 10060 37024 10100 37064
rect 9964 36520 10004 36560
rect 10636 39208 10676 39248
rect 10924 39880 10964 39920
rect 11020 39124 11060 39164
rect 10828 39040 10868 39080
rect 10540 38200 10580 38240
rect 10444 38116 10484 38156
rect 10156 36856 10196 36896
rect 10060 36352 10100 36392
rect 9964 35848 10004 35888
rect 9868 35680 9908 35720
rect 10060 35680 10100 35720
rect 9484 34084 9524 34124
rect 9676 34168 9716 34208
rect 9580 33832 9620 33872
rect 9292 32824 9332 32864
rect 9196 32152 9236 32192
rect 9100 28540 9140 28580
rect 9484 31144 9524 31184
rect 10156 33412 10196 33452
rect 10444 36772 10484 36812
rect 10348 36688 10388 36728
rect 10540 36436 10580 36476
rect 10732 38200 10772 38240
rect 10732 37948 10772 37988
rect 10732 37696 10772 37736
rect 11116 37528 11156 37568
rect 10828 37024 10868 37064
rect 11020 36940 11060 36980
rect 10732 36520 10772 36560
rect 10636 35176 10676 35216
rect 10348 34756 10388 34796
rect 10252 33244 10292 33284
rect 10060 33160 10100 33200
rect 9772 32908 9812 32948
rect 9868 32824 9908 32864
rect 11020 36436 11060 36476
rect 10828 34924 10868 34964
rect 10636 34084 10676 34124
rect 10444 33664 10484 33704
rect 12172 41392 12212 41432
rect 12172 41224 12212 41264
rect 11980 41140 12020 41180
rect 11596 41056 11636 41096
rect 12460 41308 12500 41348
rect 11596 40300 11636 40340
rect 11788 39964 11828 40004
rect 11596 39628 11636 39668
rect 11500 39208 11540 39248
rect 11404 38620 11444 38660
rect 11404 38116 11444 38156
rect 11308 36772 11348 36812
rect 11116 34504 11156 34544
rect 11020 34168 11060 34208
rect 11116 33748 11156 33788
rect 10444 33412 10484 33452
rect 10156 32824 10196 32864
rect 9868 31396 9908 31436
rect 10060 29800 10100 29840
rect 9580 29128 9620 29168
rect 9964 29128 10004 29168
rect 9484 28624 9524 28664
rect 9388 28540 9428 28580
rect 9196 28456 9236 28496
rect 9292 28036 9332 28076
rect 9292 27532 9332 27572
rect 9196 27364 9236 27404
rect 9100 26944 9140 26984
rect 8620 26020 8660 26060
rect 8716 25852 8756 25892
rect 8716 25600 8756 25640
rect 8812 25516 8852 25556
rect 9004 26272 9044 26312
rect 8908 23836 8948 23876
rect 9004 23752 9044 23792
rect 8524 23668 8564 23708
rect 8716 23584 8756 23624
rect 8140 22996 8180 23036
rect 7948 22576 7988 22616
rect 8140 22408 8180 22448
rect 8620 23248 8660 23288
rect 8332 23164 8372 23204
rect 10636 33328 10676 33368
rect 10828 32656 10868 32696
rect 10732 31564 10772 31604
rect 10540 31312 10580 31352
rect 10444 30976 10484 31016
rect 10444 29968 10484 30008
rect 10348 29296 10388 29336
rect 10348 29044 10388 29084
rect 10252 28456 10292 28496
rect 9868 27700 9908 27740
rect 9484 26944 9524 26984
rect 9484 26692 9524 26732
rect 9484 26524 9524 26564
rect 9676 24676 9716 24716
rect 9580 24340 9620 24380
rect 9292 23584 9332 23624
rect 9196 23164 9236 23204
rect 8812 23080 8852 23120
rect 9292 23080 9332 23120
rect 8524 22744 8564 22784
rect 8428 22660 8468 22700
rect 8428 22492 8468 22532
rect 7468 21736 7508 21776
rect 7564 21400 7604 21440
rect 7372 20308 7412 20348
rect 7276 19720 7316 19760
rect 6508 17704 6548 17744
rect 6508 15940 6548 15980
rect 6508 15520 6548 15560
rect 6412 14764 6452 14804
rect 6508 14092 6548 14132
rect 7660 20140 7700 20180
rect 7948 21568 7988 21608
rect 8044 21316 8084 21356
rect 8140 20812 8180 20852
rect 8044 20728 8084 20768
rect 8140 20644 8180 20684
rect 7756 19972 7796 20012
rect 8044 20476 8084 20516
rect 7852 19300 7892 19340
rect 7180 18040 7220 18080
rect 7276 17788 7316 17828
rect 6988 17704 7028 17744
rect 7468 18208 7508 18248
rect 7756 18460 7796 18500
rect 7756 17620 7796 17660
rect 7948 17620 7988 17660
rect 6796 16948 6836 16988
rect 6700 16360 6740 16400
rect 6700 16024 6740 16064
rect 6604 13756 6644 13796
rect 6604 13588 6644 13628
rect 6508 13252 6548 13292
rect 6412 12496 6452 12536
rect 6316 10984 6356 11024
rect 6412 8716 6452 8756
rect 6220 8548 6260 8588
rect 7180 16192 7220 16232
rect 7372 16948 7412 16988
rect 7377 16360 7417 16400
rect 7852 16192 7892 16232
rect 7084 16024 7124 16064
rect 6988 15772 7028 15812
rect 6892 15688 6932 15728
rect 6796 15016 6836 15056
rect 6700 12244 6740 12284
rect 6892 14848 6932 14888
rect 6988 14008 7028 14048
rect 7084 13420 7124 13460
rect 8044 17536 8084 17576
rect 8044 17032 8084 17072
rect 8044 16360 8084 16400
rect 7948 15688 7988 15728
rect 7468 15520 7508 15560
rect 7468 14848 7508 14888
rect 8332 21400 8372 21440
rect 8236 20476 8276 20516
rect 8620 21904 8660 21944
rect 8524 21568 8564 21608
rect 8620 21316 8660 21356
rect 9196 22324 9236 22364
rect 9292 22240 9332 22280
rect 9196 21904 9236 21944
rect 9004 20980 9044 21020
rect 8716 20644 8756 20684
rect 8236 20056 8276 20096
rect 8620 20056 8660 20096
rect 8236 18544 8276 18584
rect 8236 17956 8276 17996
rect 8428 19888 8468 19928
rect 8716 19888 8756 19928
rect 8620 19216 8660 19256
rect 8524 19048 8564 19088
rect 8428 18544 8468 18584
rect 8524 17116 8564 17156
rect 9484 23416 9524 23456
rect 9772 23248 9812 23288
rect 9676 23080 9716 23120
rect 9484 22996 9524 23036
rect 9580 22912 9620 22952
rect 9484 22240 9524 22280
rect 9388 21904 9428 21944
rect 9292 21820 9332 21860
rect 9196 21736 9236 21776
rect 8908 20056 8948 20096
rect 8908 19636 8948 19676
rect 8812 18880 8852 18920
rect 8716 17872 8756 17912
rect 8908 17368 8948 17408
rect 8524 16780 8564 16820
rect 8524 16276 8564 16316
rect 8524 16024 8564 16064
rect 8428 15688 8468 15728
rect 8140 14596 8180 14636
rect 7564 14008 7604 14048
rect 7756 13756 7796 13796
rect 7564 13672 7604 13712
rect 7468 13420 7508 13460
rect 7276 13000 7316 13040
rect 6892 12244 6932 12284
rect 7084 11488 7124 11528
rect 6604 9052 6644 9092
rect 6508 8128 6548 8168
rect 6124 7792 6164 7832
rect 6412 7792 6452 7832
rect 7276 11152 7316 11192
rect 7084 10984 7124 11024
rect 7084 10732 7124 10772
rect 6988 9808 7028 9848
rect 6508 7708 6548 7748
rect 6508 7540 6548 7580
rect 6412 7456 6452 7496
rect 5932 7036 5972 7076
rect 6220 6784 6260 6824
rect 5932 6448 5972 6488
rect 5836 6112 5876 6152
rect 6604 6280 6644 6320
rect 6316 6196 6356 6236
rect 5932 5356 5972 5396
rect 6316 5356 6356 5396
rect 5836 4180 5876 4220
rect 5836 2584 5876 2624
rect 6124 3760 6164 3800
rect 6220 3424 6260 3464
rect 6988 9472 7028 9512
rect 6892 9220 6932 9260
rect 7468 12496 7508 12536
rect 7660 12580 7700 12620
rect 9292 19972 9332 20012
rect 9196 19804 9236 19844
rect 9100 18880 9140 18920
rect 9292 18544 9332 18584
rect 9196 18124 9236 18164
rect 9196 17872 9236 17912
rect 9484 20980 9524 21020
rect 9484 19216 9524 19256
rect 9292 17704 9332 17744
rect 9100 17620 9140 17660
rect 9100 17116 9140 17156
rect 9196 17032 9236 17072
rect 8620 15352 8660 15392
rect 8908 15100 8948 15140
rect 8620 14764 8660 14804
rect 8812 14176 8852 14216
rect 8044 13672 8084 13712
rect 7852 12580 7892 12620
rect 7948 12496 7988 12536
rect 7564 10312 7604 10352
rect 7564 10144 7604 10184
rect 7948 11019 7988 11024
rect 7948 10984 7988 11019
rect 9100 15520 9140 15560
rect 10060 27616 10100 27656
rect 9964 24676 10004 24716
rect 11020 33664 11060 33704
rect 11020 31312 11060 31352
rect 10540 27784 10580 27824
rect 10252 27196 10292 27236
rect 10540 27616 10580 27656
rect 10156 26692 10196 26732
rect 10348 26692 10388 26732
rect 10444 26104 10484 26144
rect 10732 27700 10772 27740
rect 11116 31060 11156 31100
rect 10636 25852 10676 25892
rect 10540 25180 10580 25220
rect 10156 24508 10196 24548
rect 10060 22912 10100 22952
rect 11788 37864 11828 37904
rect 11308 35344 11348 35384
rect 11308 33664 11348 33704
rect 11020 28456 11060 28496
rect 11212 28456 11252 28496
rect 11212 28288 11252 28328
rect 11212 27700 11252 27740
rect 10924 27280 10964 27320
rect 11116 27280 11156 27320
rect 11020 27196 11060 27236
rect 10828 26776 10868 26816
rect 10828 26524 10868 26564
rect 10924 26356 10964 26396
rect 10828 26272 10868 26312
rect 10828 26020 10868 26060
rect 10828 25852 10868 25892
rect 10924 25348 10964 25388
rect 10540 24508 10580 24548
rect 10732 24508 10772 24548
rect 10444 24424 10484 24464
rect 10732 23791 10772 23792
rect 10732 23752 10772 23791
rect 11020 24592 11060 24632
rect 11212 26356 11252 26396
rect 11596 36940 11636 36980
rect 11692 36688 11732 36728
rect 11500 35428 11540 35468
rect 11500 34924 11540 34964
rect 11788 36184 11828 36224
rect 12652 40972 12692 41012
rect 12268 40216 12308 40256
rect 12172 40048 12212 40088
rect 12076 38200 12116 38240
rect 12556 40132 12596 40172
rect 12460 39712 12500 39752
rect 12364 39628 12404 39668
rect 12268 38872 12308 38912
rect 12268 38704 12308 38744
rect 12268 38452 12308 38492
rect 12268 38200 12308 38240
rect 12076 38032 12116 38072
rect 11980 37696 12020 37736
rect 12172 36772 12212 36812
rect 12268 36688 12308 36728
rect 11980 36352 12020 36392
rect 12268 36352 12308 36392
rect 11404 32992 11444 33032
rect 11692 33580 11732 33620
rect 11404 31396 11444 31436
rect 11404 30976 11444 31016
rect 13036 42400 13076 42440
rect 12940 40972 12980 41012
rect 12748 39796 12788 39836
rect 13612 42820 13652 42860
rect 13516 41560 13556 41600
rect 13708 42064 13748 42104
rect 13324 40468 13364 40508
rect 13036 39796 13076 39836
rect 12652 38956 12692 38996
rect 12556 38872 12596 38912
rect 12460 38452 12500 38492
rect 12460 38200 12500 38240
rect 12652 38452 12692 38492
rect 12556 37864 12596 37904
rect 12940 39040 12980 39080
rect 13420 40048 13460 40088
rect 13228 39292 13268 39332
rect 12844 38368 12884 38408
rect 13036 38368 13076 38408
rect 12940 38284 12980 38324
rect 12556 37276 12596 37316
rect 12460 36772 12500 36812
rect 12172 35092 12212 35132
rect 12364 35008 12404 35048
rect 12268 34924 12308 34964
rect 11980 33748 12020 33788
rect 11884 32908 11924 32948
rect 12460 34336 12500 34376
rect 12748 37528 12788 37568
rect 13132 37612 13172 37652
rect 12844 36856 12884 36896
rect 12748 36352 12788 36392
rect 12652 35176 12692 35216
rect 12748 34000 12788 34040
rect 12748 33664 12788 33704
rect 12652 32824 12692 32864
rect 12364 32656 12404 32696
rect 12556 32656 12596 32696
rect 12556 32068 12596 32108
rect 12460 31564 12500 31604
rect 11980 31480 12020 31520
rect 12364 31480 12404 31520
rect 11692 30892 11732 30932
rect 12076 30892 12116 30932
rect 11500 30220 11540 30260
rect 11884 29968 11924 30008
rect 12172 29884 12212 29924
rect 11884 29464 11924 29504
rect 11596 29128 11636 29168
rect 11980 29380 12020 29420
rect 11692 28960 11732 29000
rect 11884 28960 11924 29000
rect 11884 28372 11924 28412
rect 12076 29128 12116 29168
rect 11500 25600 11540 25640
rect 11404 25348 11444 25388
rect 11500 25180 11540 25220
rect 11404 25096 11444 25136
rect 11308 24424 11348 24464
rect 10924 23836 10964 23876
rect 10444 23668 10484 23708
rect 10348 23332 10388 23372
rect 10252 23164 10292 23204
rect 10156 22492 10196 22532
rect 9676 21988 9716 22028
rect 9868 21904 9908 21944
rect 9772 21568 9812 21608
rect 9676 18544 9716 18584
rect 9676 18292 9716 18332
rect 9580 17956 9620 17996
rect 9676 17872 9716 17912
rect 9868 18208 9908 18248
rect 9772 17620 9812 17660
rect 9484 17452 9524 17492
rect 9484 16696 9524 16736
rect 9964 17452 10004 17492
rect 9964 17032 10004 17072
rect 9868 16612 9908 16652
rect 9868 16360 9908 16400
rect 9484 16276 9524 16316
rect 9292 14932 9332 14972
rect 9196 14848 9236 14888
rect 9100 14764 9140 14804
rect 9676 14932 9716 14972
rect 9100 14092 9140 14132
rect 9292 14092 9332 14132
rect 9772 14092 9812 14132
rect 8716 13756 8756 13796
rect 8908 13672 8948 13712
rect 8620 13588 8660 13628
rect 8524 13504 8564 13544
rect 8716 13504 8756 13544
rect 8332 13000 8372 13040
rect 8524 13000 8564 13040
rect 8812 12496 8852 12536
rect 8716 12160 8756 12200
rect 8620 12076 8660 12116
rect 8332 11404 8372 11444
rect 8428 11236 8468 11276
rect 8236 11152 8276 11192
rect 8332 10984 8372 11024
rect 7756 10228 7796 10268
rect 7180 9052 7220 9092
rect 6892 7540 6932 7580
rect 7180 7204 7220 7244
rect 7180 6616 7220 6656
rect 7468 9556 7508 9596
rect 7756 9556 7796 9596
rect 7564 9304 7604 9344
rect 7468 9052 7508 9092
rect 7468 7708 7508 7748
rect 7084 6280 7124 6320
rect 6988 6196 7028 6236
rect 6892 6112 6932 6152
rect 6892 5860 6932 5900
rect 7084 5860 7124 5900
rect 6988 5608 7028 5648
rect 6796 5356 6836 5396
rect 6604 5272 6644 5312
rect 7180 5272 7220 5312
rect 6508 4768 6548 4808
rect 6508 4264 6548 4304
rect 6412 4096 6452 4136
rect 6508 3508 6548 3548
rect 7180 4936 7220 4976
rect 6700 4684 6740 4724
rect 7084 4684 7124 4724
rect 7468 5524 7508 5564
rect 7372 4852 7412 4892
rect 7372 4684 7412 4724
rect 7276 4264 7316 4304
rect 7660 8380 7700 8420
rect 8236 10396 8276 10436
rect 8044 10312 8084 10352
rect 7948 10144 7988 10184
rect 8140 10228 8180 10268
rect 8044 9556 8084 9596
rect 8524 10228 8564 10268
rect 8428 10144 8468 10184
rect 8428 9556 8468 9596
rect 8044 8716 8084 8756
rect 8236 8716 8276 8756
rect 7852 8380 7892 8420
rect 7756 7456 7796 7496
rect 7660 7036 7700 7076
rect 7756 5188 7796 5228
rect 8140 8044 8180 8084
rect 8332 7960 8372 8000
rect 8524 9052 8564 9092
rect 8236 7540 8276 7580
rect 8332 7120 8372 7160
rect 9004 12328 9044 12368
rect 9580 14008 9620 14048
rect 9484 13672 9524 13712
rect 9292 12496 9332 12536
rect 9292 12160 9332 12200
rect 9196 11908 9236 11948
rect 9196 11656 9236 11696
rect 9580 13168 9620 13208
rect 9580 12496 9620 12536
rect 9484 11908 9524 11948
rect 10252 22240 10292 22280
rect 10540 22324 10580 22364
rect 10444 22240 10484 22280
rect 10348 21652 10388 21692
rect 10156 20896 10196 20936
rect 10156 19720 10196 19760
rect 10156 19216 10196 19256
rect 10444 19888 10484 19928
rect 10444 19636 10484 19676
rect 10444 19468 10484 19508
rect 10060 13504 10100 13544
rect 10252 17704 10292 17744
rect 10252 14764 10292 14804
rect 10060 13084 10100 13124
rect 10156 12664 10196 12704
rect 10060 12496 10100 12536
rect 10060 12076 10100 12116
rect 9580 11824 9620 11864
rect 9868 11656 9908 11696
rect 10060 11656 10100 11696
rect 9292 11572 9332 11612
rect 9196 11320 9236 11360
rect 8716 10984 8756 11024
rect 9004 11152 9044 11192
rect 8908 10984 8948 11024
rect 8908 10732 8948 10772
rect 8812 10396 8852 10436
rect 9004 10480 9044 10520
rect 9196 10480 9236 10520
rect 9772 11572 9812 11612
rect 9484 11236 9524 11276
rect 9388 10732 9428 10772
rect 9292 10396 9332 10436
rect 9484 10396 9524 10436
rect 9292 10228 9332 10268
rect 8716 10060 8756 10100
rect 9196 10060 9236 10100
rect 9004 9808 9044 9848
rect 8908 9640 8948 9680
rect 8716 9304 8756 9344
rect 8620 7540 8660 7580
rect 8524 7120 8564 7160
rect 8140 6784 8180 6824
rect 9196 9556 9236 9596
rect 9484 9976 9524 10016
rect 9100 9220 9140 9260
rect 9292 9220 9332 9260
rect 8236 5608 8276 5648
rect 7468 4432 7508 4472
rect 7084 4012 7124 4052
rect 6220 3172 6260 3212
rect 6508 2920 6548 2960
rect 6316 1912 6356 1952
rect 6220 1744 6260 1784
rect 5932 1408 5972 1448
rect 6028 1324 6068 1364
rect 6124 1240 6164 1280
rect 6412 1828 6452 1868
rect 6988 3256 7028 3296
rect 6892 2836 6932 2876
rect 6796 2752 6836 2792
rect 7180 3424 7220 3464
rect 7660 4852 7700 4892
rect 7948 4432 7988 4472
rect 7948 4096 7988 4136
rect 7660 3844 7700 3884
rect 7660 3592 7700 3632
rect 7564 3508 7604 3548
rect 7276 3004 7316 3044
rect 7084 2920 7124 2960
rect 6892 2332 6932 2372
rect 6700 2164 6740 2204
rect 6604 1576 6644 1616
rect 6508 1408 6548 1448
rect 6508 1072 6548 1112
rect 5740 988 5780 1028
rect 5836 652 5876 692
rect 5644 484 5684 524
rect 6604 904 6644 944
rect 6988 1912 7028 1952
rect 7180 2584 7220 2624
rect 7852 3508 7892 3548
rect 7756 3256 7796 3296
rect 8140 3508 8180 3548
rect 8044 3424 8084 3464
rect 8524 5608 8564 5648
rect 8908 5440 8948 5480
rect 8812 5272 8852 5312
rect 8524 4768 8564 4808
rect 8620 4180 8660 4220
rect 8524 3844 8564 3884
rect 8428 3592 8468 3632
rect 9004 4936 9044 4976
rect 8908 4096 8948 4136
rect 9292 8548 9332 8588
rect 9196 7540 9236 7580
rect 9388 7372 9428 7412
rect 9196 5944 9236 5984
rect 9196 5776 9236 5816
rect 9292 5692 9332 5732
rect 9292 5272 9332 5312
rect 9964 10396 10004 10436
rect 9772 10144 9812 10184
rect 10444 17788 10484 17828
rect 10444 16024 10484 16064
rect 10540 15688 10580 15728
rect 10732 23416 10772 23456
rect 10828 23332 10868 23372
rect 10732 20056 10772 20096
rect 10828 18796 10868 18836
rect 10732 18292 10772 18332
rect 11308 23836 11348 23876
rect 11116 23668 11156 23708
rect 11692 25180 11732 25220
rect 11692 25012 11732 25052
rect 12172 27700 12212 27740
rect 12076 27364 12116 27404
rect 12076 26776 12116 26816
rect 11980 26440 12020 26480
rect 11884 25600 11924 25640
rect 12076 26104 12116 26144
rect 12556 31312 12596 31352
rect 12460 30220 12500 30260
rect 12460 29632 12500 29672
rect 12556 26440 12596 26480
rect 11404 23248 11444 23288
rect 11116 21568 11156 21608
rect 11020 21484 11060 21524
rect 11020 19636 11060 19676
rect 11308 21820 11348 21860
rect 10924 17788 10964 17828
rect 10924 17536 10964 17576
rect 11116 19216 11156 19256
rect 11212 18796 11252 18836
rect 11020 16360 11060 16400
rect 11308 18628 11348 18668
rect 11212 18124 11252 18164
rect 11788 23584 11828 23624
rect 11596 23080 11636 23120
rect 11500 21820 11540 21860
rect 11692 22156 11732 22196
rect 11692 19888 11732 19928
rect 11692 19468 11732 19508
rect 11212 17116 11252 17156
rect 11404 17200 11444 17240
rect 11404 15856 11444 15896
rect 11116 15688 11156 15728
rect 10924 15520 10964 15560
rect 10924 15268 10964 15308
rect 10828 15184 10868 15224
rect 10732 15100 10772 15140
rect 10636 14764 10676 14804
rect 10732 14512 10772 14552
rect 10732 13420 10772 13460
rect 10444 13336 10484 13376
rect 10348 13252 10388 13292
rect 10732 13000 10772 13040
rect 10444 11824 10484 11864
rect 10156 10564 10196 10604
rect 9868 9556 9908 9596
rect 10060 9304 10100 9344
rect 10348 10060 10388 10100
rect 10828 11992 10868 12032
rect 11212 15604 11252 15644
rect 11404 15520 11444 15560
rect 11308 15100 11348 15140
rect 11020 13924 11060 13964
rect 11212 13924 11252 13964
rect 11116 13168 11156 13208
rect 11116 12748 11156 12788
rect 10924 10648 10964 10688
rect 10636 10396 10676 10436
rect 10924 10312 10964 10352
rect 10348 9472 10388 9512
rect 10252 9304 10292 9344
rect 9676 8716 9716 8756
rect 10156 8464 10196 8504
rect 9676 7960 9716 8000
rect 10060 7708 10100 7748
rect 9964 7456 10004 7496
rect 9964 7204 10004 7244
rect 9772 6952 9812 6992
rect 9772 6448 9812 6488
rect 9580 6112 9620 6152
rect 9580 5860 9620 5900
rect 9100 4768 9140 4808
rect 8812 3760 8852 3800
rect 8428 3340 8468 3380
rect 7276 2500 7316 2540
rect 7564 2500 7604 2540
rect 7564 2332 7604 2372
rect 7276 2248 7316 2288
rect 7180 2164 7220 2204
rect 7180 1912 7220 1952
rect 6892 1408 6932 1448
rect 6796 1240 6836 1280
rect 6892 1156 6932 1196
rect 7084 1240 7124 1280
rect 7660 2248 7700 2288
rect 8332 2920 8372 2960
rect 8140 2836 8180 2876
rect 8044 2752 8084 2792
rect 7948 2668 7988 2708
rect 8044 2248 8084 2288
rect 7852 1828 7892 1868
rect 7660 1744 7700 1784
rect 7660 1492 7700 1532
rect 8428 2836 8468 2876
rect 8716 3340 8756 3380
rect 9004 3928 9044 3968
rect 9004 3508 9044 3548
rect 9292 3508 9332 3548
rect 8812 3256 8852 3296
rect 8620 3088 8660 3128
rect 9100 3088 9140 3128
rect 8428 2668 8468 2708
rect 8716 2584 8756 2624
rect 8716 2248 8756 2288
rect 8044 1744 8084 1784
rect 7948 1408 7988 1448
rect 8236 1912 8276 1952
rect 8428 1828 8468 1868
rect 8428 1492 8468 1532
rect 8140 1324 8180 1364
rect 7756 1240 7796 1280
rect 8332 1240 8372 1280
rect 7372 1072 7412 1112
rect 7084 988 7124 1028
rect 7465 988 7505 1028
rect 7180 904 7220 944
rect 6412 400 6452 440
rect 6220 64 6260 104
rect 6604 232 6644 272
rect 7564 652 7604 692
rect 7372 484 7412 524
rect 7180 316 7220 356
rect 6988 232 7028 272
rect 8044 1156 8084 1196
rect 7948 904 7988 944
rect 7852 652 7892 692
rect 8140 568 8180 608
rect 8236 484 8276 524
rect 8716 1408 8756 1448
rect 9196 2836 9236 2876
rect 8908 2416 8948 2456
rect 9100 2584 9140 2624
rect 9868 4264 9908 4304
rect 10060 4264 10100 4304
rect 9580 3928 9620 3968
rect 9484 3340 9524 3380
rect 9004 1912 9044 1952
rect 8908 1660 8948 1700
rect 8716 988 8756 1028
rect 8620 904 8660 944
rect 8524 736 8564 776
rect 9100 1156 9140 1196
rect 9100 988 9140 1028
rect 9100 820 9140 860
rect 9004 316 9044 356
rect 9484 1912 9524 1952
rect 9388 1408 9428 1448
rect 10060 3844 10100 3884
rect 9964 3592 10004 3632
rect 9868 3004 9908 3044
rect 9676 2584 9716 2624
rect 10252 8380 10292 8420
rect 10252 6952 10292 6992
rect 10924 10060 10964 10100
rect 10540 9304 10580 9344
rect 10636 9220 10676 9260
rect 10540 8716 10580 8756
rect 10444 8464 10484 8504
rect 10732 7792 10772 7832
rect 10636 7708 10676 7748
rect 10252 4684 10292 4724
rect 10252 4264 10292 4304
rect 10156 2836 10196 2876
rect 10060 2500 10100 2540
rect 9676 1996 9716 2036
rect 9484 904 9524 944
rect 9292 736 9332 776
rect 9292 484 9332 524
rect 9772 1912 9812 1952
rect 10348 3760 10388 3800
rect 10444 3592 10484 3632
rect 10732 7540 10772 7580
rect 11404 14848 11444 14888
rect 12076 23668 12116 23708
rect 12268 25600 12308 25640
rect 12460 25600 12500 25640
rect 12652 25348 12692 25388
rect 12268 24928 12308 24968
rect 12556 24928 12596 24968
rect 11980 23164 12020 23204
rect 11596 18544 11636 18584
rect 11788 18544 11828 18584
rect 11788 18208 11828 18248
rect 11692 17200 11732 17240
rect 11596 15604 11636 15644
rect 11980 21568 12020 21608
rect 12172 20056 12212 20096
rect 12460 22576 12500 22616
rect 12652 22492 12692 22532
rect 12652 22072 12692 22112
rect 12556 21904 12596 21944
rect 12460 21820 12500 21860
rect 13804 41224 13844 41264
rect 13708 40048 13748 40088
rect 13612 39880 13652 39920
rect 13516 39292 13556 39332
rect 13420 39208 13460 39248
rect 13420 37444 13460 37484
rect 13324 37360 13364 37400
rect 13324 36856 13364 36896
rect 13612 38872 13652 38912
rect 13612 38200 13652 38240
rect 14092 41140 14132 41180
rect 13900 41056 13940 41096
rect 14572 42484 14612 42524
rect 14476 41224 14516 41264
rect 14284 40888 14324 40928
rect 14188 40804 14228 40844
rect 14092 40552 14132 40592
rect 13900 40300 13940 40340
rect 14092 40132 14132 40172
rect 14092 39460 14132 39500
rect 13804 38032 13844 38072
rect 13708 37696 13748 37736
rect 13708 37108 13748 37148
rect 13036 35260 13076 35300
rect 13516 35176 13556 35216
rect 13324 34840 13364 34880
rect 12940 34420 12980 34460
rect 13324 34336 13364 34376
rect 13228 34252 13268 34292
rect 13036 33496 13076 33536
rect 13036 32740 13076 32780
rect 12940 32236 12980 32276
rect 12844 32152 12884 32192
rect 12844 31984 12884 32024
rect 13036 31984 13076 32024
rect 12940 31900 12980 31940
rect 13324 34084 13364 34124
rect 13708 35260 13748 35300
rect 13612 34420 13652 34460
rect 13900 37528 13940 37568
rect 13900 37108 13940 37148
rect 13900 35344 13940 35384
rect 14476 40552 14516 40592
rect 14284 40468 14324 40508
rect 14668 41560 14708 41600
rect 15052 41728 15092 41768
rect 14860 41644 14900 41684
rect 15436 42232 15476 42272
rect 15436 42064 15476 42104
rect 14860 40552 14900 40592
rect 14764 40468 14804 40508
rect 14284 39880 14324 39920
rect 14572 39796 14612 39836
rect 14284 37864 14324 37904
rect 14188 37108 14228 37148
rect 14188 36772 14228 36812
rect 15052 41056 15092 41096
rect 15244 40552 15284 40592
rect 15148 40300 15188 40340
rect 15820 42064 15860 42104
rect 16012 41896 16052 41936
rect 16300 42148 16340 42188
rect 16588 42148 16628 42188
rect 16588 41644 16628 41684
rect 16396 41560 16436 41600
rect 16492 41476 16532 41516
rect 16300 41392 16340 41432
rect 15532 41056 15572 41096
rect 15436 40888 15476 40928
rect 15340 40216 15380 40256
rect 15628 40972 15668 41012
rect 15628 40384 15668 40424
rect 14956 40132 14996 40172
rect 15532 39964 15572 40004
rect 14956 38200 14996 38240
rect 15820 41140 15860 41180
rect 16012 40972 16052 41012
rect 16012 40552 16052 40592
rect 15724 39880 15764 39920
rect 15532 39040 15572 39080
rect 15628 38704 15668 38744
rect 15436 38368 15476 38408
rect 15052 38032 15092 38072
rect 15148 37864 15188 37904
rect 15052 37780 15092 37820
rect 14572 37528 14612 37568
rect 14860 37276 14900 37316
rect 14668 36856 14708 36896
rect 14956 36856 14996 36896
rect 15436 38200 15476 38240
rect 15340 38032 15380 38072
rect 15244 37780 15284 37820
rect 15916 39040 15956 39080
rect 15628 37864 15668 37904
rect 15148 37696 15188 37736
rect 14956 36520 14996 36560
rect 14572 35932 14612 35972
rect 14284 35260 14324 35300
rect 14476 35260 14516 35300
rect 13900 34924 13940 34964
rect 13804 34672 13844 34712
rect 13804 34420 13844 34460
rect 13516 34000 13556 34040
rect 13420 33664 13460 33704
rect 13420 33496 13460 33536
rect 13804 33496 13844 33536
rect 13516 33412 13556 33452
rect 13324 31564 13364 31604
rect 13228 29128 13268 29168
rect 13036 27616 13076 27656
rect 13132 26944 13172 26984
rect 12940 22660 12980 22700
rect 12844 22324 12884 22364
rect 12844 22072 12884 22112
rect 12940 21820 12980 21860
rect 12460 20644 12500 20684
rect 12748 20728 12788 20768
rect 12940 20644 12980 20684
rect 12844 20140 12884 20180
rect 12364 19804 12404 19844
rect 12748 20056 12788 20096
rect 12940 20056 12980 20096
rect 12652 19972 12692 20012
rect 12460 19132 12500 19172
rect 11980 16696 12020 16736
rect 11692 13504 11732 13544
rect 11692 13336 11732 13376
rect 12268 16612 12308 16652
rect 12172 16276 12212 16316
rect 12076 15940 12116 15980
rect 11884 15856 11924 15896
rect 13420 28288 13460 28328
rect 13228 26776 13268 26816
rect 13804 31480 13844 31520
rect 13708 30724 13748 30764
rect 13612 30640 13652 30680
rect 14668 35344 14708 35384
rect 14380 34840 14420 34880
rect 14284 34420 14324 34460
rect 14380 34000 14420 34040
rect 14188 33664 14228 33704
rect 14476 33664 14516 33704
rect 14956 35260 14996 35300
rect 14764 34672 14804 34712
rect 14860 34420 14900 34460
rect 14668 33076 14708 33116
rect 14668 32908 14708 32948
rect 14572 32824 14612 32864
rect 14188 32152 14228 32192
rect 14092 31312 14132 31352
rect 15052 34672 15092 34712
rect 15436 37612 15476 37652
rect 15244 37192 15284 37232
rect 15340 36856 15380 36896
rect 15628 37024 15668 37064
rect 15532 36604 15572 36644
rect 15436 36520 15476 36560
rect 15436 36352 15476 36392
rect 15244 35932 15284 35972
rect 14956 34168 14996 34208
rect 15148 34168 15188 34208
rect 15052 33916 15092 33956
rect 14860 32656 14900 32696
rect 14860 32068 14900 32108
rect 14860 31312 14900 31352
rect 14668 31228 14708 31268
rect 14188 30724 14228 30764
rect 13996 29800 14036 29840
rect 13900 29380 13940 29420
rect 13804 29212 13844 29252
rect 13996 29128 14036 29168
rect 13996 28960 14036 29000
rect 13900 28456 13940 28496
rect 13612 26944 13652 26984
rect 13612 26776 13652 26816
rect 13516 26020 13556 26060
rect 13708 26104 13748 26144
rect 13996 27616 14036 27656
rect 14380 29380 14420 29420
rect 14380 28792 14420 28832
rect 14764 30556 14804 30596
rect 14956 30220 14996 30260
rect 14956 30052 14996 30092
rect 14860 29380 14900 29420
rect 14860 29044 14900 29084
rect 13900 26356 13940 26396
rect 13900 26104 13940 26144
rect 13804 26020 13844 26060
rect 13804 25432 13844 25472
rect 14284 27364 14324 27404
rect 14284 26944 14324 26984
rect 14188 25264 14228 25304
rect 14284 25180 14324 25220
rect 13612 23164 13652 23204
rect 13228 22660 13268 22700
rect 13132 22492 13172 22532
rect 13516 22492 13556 22532
rect 13132 22240 13172 22280
rect 13324 22072 13364 22112
rect 13324 21820 13364 21860
rect 13420 21652 13460 21692
rect 13228 20812 13268 20852
rect 13420 19972 13460 20012
rect 12460 18376 12500 18416
rect 12364 15688 12404 15728
rect 11596 12244 11636 12284
rect 11500 12076 11540 12116
rect 11596 11992 11636 12032
rect 11116 9472 11156 9512
rect 11308 10564 11348 10604
rect 11404 10480 11444 10520
rect 11308 10228 11348 10268
rect 11404 10144 11444 10184
rect 11596 10984 11636 11024
rect 11500 10060 11540 10100
rect 11116 9304 11156 9344
rect 11212 8296 11252 8336
rect 11788 12076 11828 12116
rect 11980 15184 12020 15224
rect 12844 19216 12884 19256
rect 13132 19207 13172 19247
rect 13324 19216 13364 19256
rect 12940 19048 12980 19088
rect 12652 15688 12692 15728
rect 12556 15520 12596 15560
rect 12748 15520 12788 15560
rect 12556 15352 12596 15392
rect 12460 14932 12500 14972
rect 11980 13504 12020 13544
rect 11884 11824 11924 11864
rect 11788 11488 11828 11528
rect 12460 14680 12500 14720
rect 12268 14260 12308 14300
rect 12748 14680 12788 14720
rect 12652 14512 12692 14552
rect 13036 18880 13076 18920
rect 13228 19048 13268 19088
rect 13516 19216 13556 19256
rect 13324 18712 13364 18752
rect 13516 18628 13556 18668
rect 13132 17116 13172 17156
rect 13036 16192 13076 16232
rect 12940 15688 12980 15728
rect 13036 15520 13076 15560
rect 13420 15352 13460 15392
rect 13036 15100 13076 15140
rect 12940 14848 12980 14888
rect 13228 14680 13268 14720
rect 13036 14428 13076 14468
rect 12172 13840 12212 13880
rect 12364 13840 12404 13880
rect 12460 13420 12500 13460
rect 12172 12832 12212 12872
rect 12076 12664 12116 12704
rect 12076 11572 12116 11612
rect 11884 11320 11924 11360
rect 11884 11152 11924 11192
rect 11788 11068 11828 11108
rect 11788 8716 11828 8756
rect 11212 7960 11252 8000
rect 11692 7960 11732 8000
rect 11404 7792 11444 7832
rect 11308 7708 11348 7748
rect 11308 7540 11348 7580
rect 11212 7372 11252 7412
rect 11116 6532 11156 6572
rect 10636 4180 10676 4220
rect 10636 3844 10676 3884
rect 11020 4852 11060 4892
rect 11020 3760 11060 3800
rect 11404 7372 11444 7412
rect 11404 6616 11444 6656
rect 11788 6616 11828 6656
rect 11404 4936 11444 4976
rect 12268 12496 12308 12536
rect 12172 11068 12212 11108
rect 12940 14176 12980 14216
rect 13228 14008 13268 14048
rect 12844 13756 12884 13796
rect 12748 13420 12788 13460
rect 12556 13084 12596 13124
rect 13132 13084 13172 13124
rect 12844 12580 12884 12620
rect 13132 12580 13172 12620
rect 13036 12496 13076 12536
rect 12556 11992 12596 12032
rect 13420 14680 13460 14720
rect 13900 23752 13940 23792
rect 13900 21568 13940 21608
rect 13900 21316 13940 21356
rect 13708 20812 13748 20852
rect 13900 19216 13940 19256
rect 13804 19132 13844 19172
rect 13708 18964 13748 19004
rect 13900 18796 13940 18836
rect 14572 27616 14612 27656
rect 14476 27196 14516 27236
rect 14476 25264 14516 25304
rect 14380 24256 14420 24296
rect 14764 27196 14804 27236
rect 15820 38368 15860 38408
rect 16012 38788 16052 38828
rect 15916 36604 15956 36644
rect 16012 36520 16052 36560
rect 15628 35176 15668 35216
rect 15532 34672 15572 34712
rect 15244 34000 15284 34040
rect 15436 34000 15476 34040
rect 15340 33496 15380 33536
rect 15532 33496 15572 33536
rect 15436 33328 15476 33368
rect 15340 32488 15380 32528
rect 15340 30724 15380 30764
rect 15916 35344 15956 35384
rect 15916 35092 15956 35132
rect 15724 34756 15764 34796
rect 15820 34672 15860 34712
rect 15724 34336 15764 34376
rect 15724 33244 15764 33284
rect 15820 32740 15860 32780
rect 15820 32152 15860 32192
rect 15724 30640 15764 30680
rect 15244 29632 15284 29672
rect 15244 28456 15284 28496
rect 15628 30136 15668 30176
rect 15436 29296 15476 29336
rect 15340 28204 15380 28244
rect 15532 28456 15572 28496
rect 14956 26944 14996 26984
rect 14668 26440 14708 26480
rect 14956 26776 14996 26816
rect 14860 26356 14900 26396
rect 14860 26104 14900 26144
rect 14860 25768 14900 25808
rect 14764 25432 14804 25472
rect 15340 27028 15380 27068
rect 15244 26272 15284 26312
rect 15052 25432 15092 25472
rect 14764 24508 14804 24548
rect 14860 23668 14900 23708
rect 14764 23164 14804 23204
rect 14668 22324 14708 22364
rect 14764 22261 14804 22280
rect 14764 22240 14804 22261
rect 14860 21904 14900 21944
rect 14380 21598 14420 21608
rect 14380 21568 14420 21598
rect 14956 21568 14996 21608
rect 14572 21484 14612 21524
rect 14476 21316 14516 21356
rect 14284 20896 14324 20936
rect 14380 20728 14420 20768
rect 14284 20644 14324 20684
rect 15436 25096 15476 25136
rect 15148 24592 15188 24632
rect 15244 24004 15284 24044
rect 15628 26608 15668 26648
rect 15628 24004 15668 24044
rect 15820 29212 15860 29252
rect 16204 41140 16244 41180
rect 16204 40468 16244 40508
rect 16204 38956 16244 38996
rect 16108 35176 16148 35216
rect 16492 40972 16532 41012
rect 16396 40552 16436 40592
rect 16684 41224 16724 41264
rect 16972 41728 17012 41768
rect 17356 42568 17396 42608
rect 17356 42316 17396 42356
rect 17164 40636 17204 40676
rect 17068 40216 17108 40256
rect 16492 39796 16532 39836
rect 16684 39796 16724 39836
rect 16396 38788 16436 38828
rect 16300 37612 16340 37652
rect 16300 37444 16340 37484
rect 16108 34840 16148 34880
rect 16012 34336 16052 34376
rect 16012 34168 16052 34208
rect 16012 32320 16052 32360
rect 16204 33496 16244 33536
rect 16108 31900 16148 31940
rect 16108 31228 16148 31268
rect 16108 30892 16148 30932
rect 16108 29884 16148 29924
rect 16012 27532 16052 27572
rect 16108 27364 16148 27404
rect 16108 25600 16148 25640
rect 15820 24256 15860 24296
rect 15532 23920 15572 23960
rect 15532 22996 15572 23036
rect 15532 22828 15572 22868
rect 15340 21232 15380 21272
rect 14476 19720 14516 19760
rect 14092 19048 14132 19088
rect 13996 18292 14036 18332
rect 13804 17704 13844 17744
rect 13900 17116 13940 17156
rect 13708 17032 13748 17072
rect 13708 16780 13748 16820
rect 13612 15100 13652 15140
rect 13612 14680 13652 14720
rect 13996 15520 14036 15560
rect 13996 15100 14036 15140
rect 13804 14932 13844 14972
rect 14188 17032 14228 17072
rect 14380 19216 14420 19256
rect 14380 18292 14420 18332
rect 14284 16612 14324 16652
rect 14668 19132 14708 19172
rect 14668 18964 14708 19004
rect 14572 18796 14612 18836
rect 14764 18712 14804 18752
rect 14572 17956 14612 17996
rect 14284 15604 14324 15644
rect 14476 15604 14516 15644
rect 14380 14932 14420 14972
rect 13804 14596 13844 14636
rect 13324 12496 13364 12536
rect 13516 12496 13556 12536
rect 13420 12412 13460 12452
rect 12748 11740 12788 11780
rect 13036 11992 13076 12032
rect 13228 11992 13268 12032
rect 12844 11488 12884 11528
rect 12748 11404 12788 11444
rect 12364 11152 12404 11192
rect 12748 11152 12788 11192
rect 12460 10816 12500 10856
rect 12844 10816 12884 10856
rect 12940 10564 12980 10604
rect 12652 10060 12692 10100
rect 12556 9640 12596 9680
rect 12460 9136 12500 9176
rect 12460 7792 12500 7832
rect 12652 9556 12692 9596
rect 12748 9388 12788 9428
rect 12556 7456 12596 7496
rect 11980 4684 12020 4724
rect 11980 4096 12020 4136
rect 10924 3508 10964 3548
rect 11116 3508 11156 3548
rect 11404 3424 11444 3464
rect 10156 2248 10196 2288
rect 10348 1828 10388 1868
rect 10540 1240 10580 1280
rect 11980 3004 12020 3044
rect 11500 2752 11540 2792
rect 11020 2584 11060 2624
rect 11212 2500 11252 2540
rect 10732 1828 10772 1868
rect 10924 1324 10964 1364
rect 9868 1156 9908 1196
rect 10348 1156 10388 1196
rect 10636 1156 10676 1196
rect 11116 1828 11156 1868
rect 11500 1744 11540 1784
rect 11308 1660 11348 1700
rect 11116 1408 11156 1448
rect 9868 568 9908 608
rect 10252 904 10292 944
rect 10156 400 10196 440
rect 10444 652 10484 692
rect 10732 904 10772 944
rect 10828 820 10868 860
rect 11692 1240 11732 1280
rect 11212 988 11252 1028
rect 11404 904 11444 944
rect 10540 484 10580 524
rect 10636 64 10676 104
rect 11020 316 11060 356
rect 12172 7120 12212 7160
rect 12460 7036 12500 7076
rect 12268 6532 12308 6572
rect 12364 5104 12404 5144
rect 12268 4096 12308 4136
rect 12460 5020 12500 5060
rect 13324 11656 13364 11696
rect 13420 11572 13460 11612
rect 13708 13084 13748 13124
rect 13612 12412 13652 12452
rect 13612 11992 13652 12032
rect 13612 11488 13652 11528
rect 13516 11404 13556 11444
rect 13132 10984 13172 11024
rect 13228 10732 13268 10772
rect 13228 10480 13268 10520
rect 13132 10144 13172 10184
rect 13036 9640 13076 9680
rect 12940 9556 12980 9596
rect 12940 7792 12980 7832
rect 13036 5692 13076 5732
rect 12652 5020 12692 5060
rect 12460 4012 12500 4052
rect 13228 5776 13268 5816
rect 13228 5440 13268 5480
rect 13036 4852 13076 4892
rect 13228 4852 13268 4892
rect 12844 3844 12884 3884
rect 12364 3424 12404 3464
rect 12844 3424 12884 3464
rect 12652 2500 12692 2540
rect 12748 2248 12788 2288
rect 12652 1828 12692 1868
rect 12364 1660 12404 1700
rect 12172 1324 12212 1364
rect 11980 904 12020 944
rect 11596 568 11636 608
rect 11404 484 11444 524
rect 11596 400 11636 440
rect 12556 1240 12596 1280
rect 12748 1744 12788 1784
rect 12748 1072 12788 1112
rect 13228 4684 13268 4724
rect 13132 3928 13172 3968
rect 13036 2584 13076 2624
rect 13420 11320 13460 11360
rect 14092 14596 14132 14636
rect 14092 14260 14132 14300
rect 14284 14260 14324 14300
rect 14188 14176 14228 14216
rect 14188 13672 14228 13712
rect 14476 14008 14516 14048
rect 14476 13672 14516 13712
rect 13804 12664 13844 12704
rect 13804 12412 13844 12452
rect 14092 11992 14132 12032
rect 13996 11824 14036 11864
rect 13900 11488 13940 11528
rect 14092 11404 14132 11444
rect 13708 10564 13748 10604
rect 14092 10564 14132 10604
rect 13516 10480 13556 10520
rect 13612 10060 13652 10100
rect 13420 7120 13460 7160
rect 13420 6952 13460 6992
rect 14668 17788 14708 17828
rect 15244 20476 15284 20516
rect 14956 19888 14996 19928
rect 15052 19804 15092 19844
rect 15436 20392 15476 20432
rect 15244 19636 15284 19676
rect 14956 19216 14996 19256
rect 15148 18964 15188 19004
rect 15052 18796 15092 18836
rect 14860 18460 14900 18500
rect 14956 18292 14996 18332
rect 15244 17956 15284 17996
rect 15244 17788 15284 17828
rect 15052 17452 15092 17492
rect 15628 20140 15668 20180
rect 15820 22660 15860 22700
rect 15916 20896 15956 20936
rect 15820 20476 15860 20516
rect 15916 20056 15956 20096
rect 15820 19972 15860 20012
rect 15724 19804 15764 19844
rect 15532 19636 15572 19676
rect 15436 19048 15476 19088
rect 15820 18880 15860 18920
rect 15628 18712 15668 18752
rect 15820 18712 15860 18752
rect 14956 17284 14996 17324
rect 15148 17284 15188 17324
rect 14764 17200 14804 17240
rect 14668 16612 14708 16652
rect 15148 17116 15188 17156
rect 14956 16276 14996 16316
rect 14860 14848 14900 14888
rect 14764 14764 14804 14804
rect 14668 14428 14708 14468
rect 14949 14680 14956 14720
rect 14956 14680 14989 14720
rect 15052 14680 15092 14720
rect 14860 14428 14900 14468
rect 15724 18292 15764 18332
rect 15628 18208 15668 18248
rect 15724 17788 15764 17828
rect 15340 17032 15380 17072
rect 16108 22240 16148 22280
rect 16108 21400 16148 21440
rect 16108 20812 16148 20852
rect 16588 36604 16628 36644
rect 16492 35764 16532 35804
rect 16684 36268 16724 36308
rect 16684 36100 16724 36140
rect 16684 34756 16724 34796
rect 16492 34336 16532 34376
rect 16684 34168 16724 34208
rect 16588 33916 16628 33956
rect 16492 33412 16532 33452
rect 16300 33244 16340 33284
rect 16588 32824 16628 32864
rect 16684 32740 16724 32780
rect 16492 32404 16532 32444
rect 16492 31396 16532 31436
rect 16300 29968 16340 30008
rect 16492 29380 16532 29420
rect 16876 39460 16916 39500
rect 17260 39544 17300 39584
rect 17164 39208 17204 39248
rect 17452 41812 17492 41852
rect 17836 42232 17876 42272
rect 17548 41644 17588 41684
rect 17740 41560 17780 41600
rect 17644 40804 17684 40844
rect 17644 40384 17684 40424
rect 18220 42148 18260 42188
rect 18124 41980 18164 42020
rect 17932 41560 17972 41600
rect 17836 40300 17876 40340
rect 17548 39880 17588 39920
rect 16972 39040 17012 39080
rect 17740 39628 17780 39668
rect 16876 38704 16916 38744
rect 16876 37696 16916 37736
rect 16876 37108 16916 37148
rect 16876 36100 16916 36140
rect 16876 35932 16916 35972
rect 16876 35428 16916 35468
rect 16876 34252 16916 34292
rect 17068 38704 17108 38744
rect 17068 37696 17108 37736
rect 18028 40468 18068 40508
rect 18028 39628 18068 39668
rect 18028 39208 18068 39248
rect 18316 40888 18356 40928
rect 18700 42148 18740 42188
rect 18604 42064 18644 42104
rect 18892 42064 18932 42104
rect 18508 41560 18548 41600
rect 18988 41896 19028 41936
rect 18700 41644 18740 41684
rect 18508 40888 18548 40928
rect 19084 41812 19124 41852
rect 18796 41308 18836 41348
rect 19180 40972 19220 41012
rect 18808 40804 18848 40844
rect 18890 40804 18930 40844
rect 18972 40804 19012 40844
rect 19054 40804 19094 40844
rect 19136 40804 19176 40844
rect 18412 39880 18452 39920
rect 18124 39124 18164 39164
rect 17740 38704 17780 38744
rect 19468 42484 19508 42524
rect 19468 42064 19508 42104
rect 19372 41392 19412 41432
rect 19372 40720 19412 40760
rect 19084 40636 19124 40676
rect 18700 40552 18740 40592
rect 18892 40468 18932 40508
rect 18700 40216 18740 40256
rect 18988 40048 19028 40088
rect 19852 41980 19892 42020
rect 19564 41140 19604 41180
rect 19756 40972 19796 41012
rect 20048 41560 20088 41600
rect 20130 41560 20170 41600
rect 20212 41560 20252 41600
rect 20294 41560 20334 41600
rect 20376 41560 20416 41600
rect 19948 40720 19988 40760
rect 19660 40468 19700 40508
rect 19756 40132 19796 40172
rect 19180 39880 19220 39920
rect 18796 39628 18836 39668
rect 18808 39292 18848 39332
rect 18890 39292 18930 39332
rect 18972 39292 19012 39332
rect 19054 39292 19094 39332
rect 19136 39292 19176 39332
rect 20048 40048 20088 40088
rect 20130 40048 20170 40088
rect 20212 40048 20252 40088
rect 20294 40048 20334 40088
rect 20376 40048 20416 40088
rect 21004 39712 21044 39752
rect 19948 39628 19988 39668
rect 20140 39544 20180 39584
rect 19564 39460 19604 39500
rect 19372 39376 19412 39416
rect 18220 38704 18260 38744
rect 18412 38284 18452 38324
rect 17452 38200 17492 38240
rect 17356 38032 17396 38072
rect 17260 37948 17300 37988
rect 17356 37864 17396 37904
rect 17164 37444 17204 37484
rect 17260 37360 17300 37400
rect 17068 36856 17108 36896
rect 17452 37528 17492 37568
rect 17836 38200 17876 38240
rect 17740 37948 17780 37988
rect 18220 37444 18260 37484
rect 17836 37360 17876 37400
rect 18124 37108 18164 37148
rect 17836 36856 17876 36896
rect 17356 36604 17396 36644
rect 17452 36268 17492 36308
rect 17068 35764 17108 35804
rect 17068 35008 17108 35048
rect 17260 35008 17300 35048
rect 17356 34504 17396 34544
rect 17068 33664 17108 33704
rect 16972 33076 17012 33116
rect 17356 32992 17396 33032
rect 17260 32572 17300 32612
rect 16876 32320 16916 32360
rect 17068 31312 17108 31352
rect 16972 30640 17012 30680
rect 16300 28876 16340 28916
rect 16588 29128 16628 29168
rect 17260 29800 17300 29840
rect 17644 35932 17684 35972
rect 17644 35176 17684 35216
rect 17644 34672 17684 34712
rect 17548 33699 17588 33704
rect 17548 33664 17588 33699
rect 17740 34420 17780 34460
rect 17548 32824 17588 32864
rect 17740 32824 17780 32864
rect 17452 32488 17492 32528
rect 17452 32320 17492 32360
rect 17356 29296 17396 29336
rect 16684 28876 16724 28916
rect 16876 28456 16916 28496
rect 16396 28204 16436 28244
rect 16300 25852 16340 25892
rect 16300 25600 16340 25640
rect 16492 27952 16532 27992
rect 16492 27616 16532 27656
rect 17068 28120 17108 28160
rect 16684 27868 16724 27908
rect 17068 27868 17108 27908
rect 16492 25852 16532 25892
rect 16300 24424 16340 24464
rect 16492 24424 16532 24464
rect 16396 22828 16436 22868
rect 16300 21400 16340 21440
rect 16492 22492 16532 22532
rect 16396 20812 16436 20852
rect 16012 18796 16052 18836
rect 16012 18544 16052 18584
rect 16012 18208 16052 18248
rect 16012 17956 16052 17996
rect 16012 17704 16052 17744
rect 15916 16696 15956 16736
rect 15628 16444 15668 16484
rect 15340 15016 15380 15056
rect 15244 14680 15284 14720
rect 14764 14260 14804 14300
rect 14668 14008 14708 14048
rect 14764 13924 14804 13964
rect 14764 13168 14804 13208
rect 14956 14176 14996 14216
rect 14956 13840 14996 13880
rect 14860 11992 14900 12032
rect 14572 11824 14612 11864
rect 14860 11824 14900 11864
rect 14284 11572 14324 11612
rect 14476 11656 14516 11696
rect 14380 11488 14420 11528
rect 14476 11404 14516 11444
rect 14188 10480 14228 10520
rect 14572 11152 14612 11192
rect 14572 10648 14612 10688
rect 13804 9640 13844 9680
rect 13708 9136 13748 9176
rect 13612 6868 13652 6908
rect 14092 9388 14132 9428
rect 13996 8380 14036 8420
rect 13900 7960 13940 8000
rect 13900 7792 13940 7832
rect 13804 6784 13844 6824
rect 13420 6448 13460 6488
rect 13420 5944 13460 5984
rect 13612 5944 13652 5984
rect 13420 5692 13460 5732
rect 13804 6448 13844 6488
rect 13708 5524 13748 5564
rect 13708 3928 13748 3968
rect 13420 3844 13460 3884
rect 13420 2164 13460 2204
rect 12652 988 12692 1028
rect 13324 904 13364 944
rect 14188 8548 14228 8588
rect 14188 8380 14228 8420
rect 14092 7624 14132 7664
rect 13996 7372 14036 7412
rect 14092 7288 14132 7328
rect 13996 7036 14036 7076
rect 14284 7792 14324 7832
rect 14284 7120 14324 7160
rect 14476 9724 14516 9764
rect 14668 10060 14708 10100
rect 14476 8548 14516 8588
rect 14476 7288 14516 7328
rect 15148 13504 15188 13544
rect 15052 13168 15092 13208
rect 15244 13168 15284 13208
rect 15052 12916 15092 12956
rect 15052 12076 15092 12116
rect 15148 11656 15188 11696
rect 14956 11404 14996 11444
rect 15148 10648 15188 10688
rect 15148 10228 15188 10268
rect 14949 10060 14989 10100
rect 15052 10060 15092 10100
rect 15532 16192 15572 16232
rect 15916 16192 15956 16232
rect 15724 15520 15764 15560
rect 15916 15520 15956 15560
rect 15724 14932 15764 14972
rect 15628 14512 15668 14552
rect 15436 13588 15476 13628
rect 15532 13420 15572 13460
rect 15532 13084 15572 13124
rect 15820 13840 15860 13880
rect 15724 12916 15764 12956
rect 15628 12496 15668 12536
rect 15532 11824 15572 11864
rect 15436 10480 15476 10520
rect 15916 13336 15956 13376
rect 16204 19888 16244 19928
rect 16300 18880 16340 18920
rect 16204 17956 16244 17996
rect 16204 17788 16244 17828
rect 18028 36772 18068 36812
rect 17932 35932 17972 35972
rect 18124 35512 18164 35552
rect 18124 35260 18164 35300
rect 18028 34672 18068 34712
rect 18316 36856 18356 36896
rect 18316 36436 18356 36476
rect 18508 37612 18548 37652
rect 18508 37360 18548 37400
rect 18412 36352 18452 36392
rect 18316 35764 18356 35804
rect 18124 34336 18164 34376
rect 18316 33664 18356 33704
rect 18220 33580 18260 33620
rect 18412 33412 18452 33452
rect 18028 32824 18068 32864
rect 17932 32740 17972 32780
rect 17740 31312 17780 31352
rect 17740 29800 17780 29840
rect 17260 27784 17300 27824
rect 17164 26860 17204 26900
rect 16780 23500 16820 23540
rect 16876 22660 16916 22700
rect 17068 24424 17108 24464
rect 17260 26104 17300 26144
rect 17260 24760 17300 24800
rect 17548 28456 17588 28496
rect 17452 27364 17492 27404
rect 17644 26776 17684 26816
rect 17644 25600 17684 25640
rect 17644 25432 17684 25472
rect 17548 24592 17588 24632
rect 17452 24508 17492 24548
rect 17356 24424 17396 24464
rect 16972 22240 17012 22280
rect 16588 20812 16628 20852
rect 17164 23920 17204 23960
rect 17548 24256 17588 24296
rect 17836 28876 17876 28916
rect 18028 30640 18068 30680
rect 18220 32488 18260 32528
rect 18412 30808 18452 30848
rect 18316 30640 18356 30680
rect 18124 28540 18164 28580
rect 18028 28288 18068 28328
rect 18124 28204 18164 28244
rect 18028 27952 18068 27992
rect 17932 27868 17972 27908
rect 17836 26776 17876 26816
rect 17836 26440 17876 26480
rect 18124 27364 18164 27404
rect 18316 29464 18356 29504
rect 18700 38788 18740 38828
rect 19180 39124 19220 39164
rect 18988 38704 19028 38744
rect 19276 38788 19316 38828
rect 19372 38704 19412 38744
rect 18988 38536 19028 38576
rect 18796 38368 18836 38408
rect 19084 37948 19124 37988
rect 18808 37780 18848 37820
rect 18890 37780 18930 37820
rect 18972 37780 19012 37820
rect 19054 37780 19094 37820
rect 19136 37780 19176 37820
rect 18892 37444 18932 37484
rect 18796 37360 18836 37400
rect 18700 37024 18740 37064
rect 19468 38368 19508 38408
rect 19372 38284 19412 38324
rect 20044 38872 20084 38912
rect 19660 38116 19700 38156
rect 19372 37948 19412 37988
rect 19660 37864 19700 37904
rect 19948 38704 19988 38744
rect 20048 38536 20088 38576
rect 20130 38536 20170 38576
rect 20212 38536 20252 38576
rect 20294 38536 20334 38576
rect 20376 38536 20416 38576
rect 20140 38284 20180 38324
rect 19948 37948 19988 37988
rect 21004 38620 21044 38660
rect 20908 37948 20948 37988
rect 20620 37864 20660 37904
rect 20524 37696 20564 37736
rect 20044 37444 20084 37484
rect 19852 37360 19892 37400
rect 19660 37276 19700 37316
rect 19180 36856 19220 36896
rect 19564 37108 19604 37148
rect 19564 36856 19604 36896
rect 19468 36688 19508 36728
rect 18892 36436 18932 36476
rect 18700 36352 18740 36392
rect 18808 36268 18848 36308
rect 18890 36268 18930 36308
rect 18972 36268 19012 36308
rect 19054 36268 19094 36308
rect 19136 36268 19176 36308
rect 19372 36604 19412 36644
rect 19564 35932 19604 35972
rect 19276 35848 19316 35888
rect 19084 35680 19124 35720
rect 18604 35176 18644 35216
rect 18604 34420 18644 34460
rect 19276 35260 19316 35300
rect 20048 37024 20088 37064
rect 20130 37024 20170 37064
rect 20212 37024 20252 37064
rect 20294 37024 20334 37064
rect 20376 37024 20416 37064
rect 19756 35680 19796 35720
rect 19948 36520 19988 36560
rect 19948 35932 19988 35972
rect 20716 37360 20756 37400
rect 20620 36016 20660 36056
rect 20524 35848 20564 35888
rect 20048 35512 20088 35552
rect 20130 35512 20170 35552
rect 20212 35512 20252 35552
rect 20294 35512 20334 35552
rect 20376 35512 20416 35552
rect 19948 35344 19988 35384
rect 19852 35260 19892 35300
rect 19948 35176 19988 35216
rect 19468 35092 19508 35132
rect 18808 34756 18848 34796
rect 18890 34756 18930 34796
rect 18972 34756 19012 34796
rect 19054 34756 19094 34796
rect 19136 34756 19176 34796
rect 18700 34336 18740 34376
rect 18796 34168 18836 34208
rect 18988 33580 19028 33620
rect 18892 33496 18932 33536
rect 19180 33496 19220 33536
rect 19372 34084 19412 34124
rect 19372 33748 19412 33788
rect 18796 33412 18836 33452
rect 19276 33412 19316 33452
rect 19564 34168 19604 34208
rect 19852 34588 19892 34628
rect 19756 34504 19796 34544
rect 20620 34336 20660 34376
rect 19852 33832 19892 33872
rect 19660 33664 19700 33704
rect 20044 34168 20084 34208
rect 20048 34000 20088 34040
rect 20130 34000 20170 34040
rect 20212 34000 20252 34040
rect 20294 34000 20334 34040
rect 20376 34000 20416 34040
rect 18808 33244 18848 33284
rect 18890 33244 18930 33284
rect 18972 33244 19012 33284
rect 19054 33244 19094 33284
rect 19136 33244 19176 33284
rect 18604 32740 18644 32780
rect 18808 31732 18848 31772
rect 18890 31732 18930 31772
rect 18972 31732 19012 31772
rect 19054 31732 19094 31772
rect 19136 31732 19176 31772
rect 19660 33160 19700 33200
rect 19564 33076 19604 33116
rect 19372 32908 19412 32948
rect 19276 31480 19316 31520
rect 18604 31312 18644 31352
rect 18796 30640 18836 30680
rect 19948 33412 19988 33452
rect 20044 32992 20084 33032
rect 19948 32740 19988 32780
rect 20048 32488 20088 32528
rect 20130 32488 20170 32528
rect 20212 32488 20252 32528
rect 20294 32488 20334 32528
rect 20376 32488 20416 32528
rect 19852 32404 19892 32444
rect 19564 31900 19604 31940
rect 19564 31312 19604 31352
rect 19276 30724 19316 30764
rect 18808 30220 18848 30260
rect 18890 30220 18930 30260
rect 18972 30220 19012 30260
rect 19054 30220 19094 30260
rect 19136 30220 19176 30260
rect 18796 30052 18836 30092
rect 18508 29296 18548 29336
rect 18700 29296 18740 29336
rect 18508 29128 18548 29168
rect 19564 30220 19604 30260
rect 21292 36856 21332 36896
rect 20908 36352 20948 36392
rect 21388 35848 21428 35888
rect 21388 35680 21428 35720
rect 21292 34672 21332 34712
rect 20812 33496 20852 33536
rect 20716 31984 20756 32024
rect 21196 33244 21236 33284
rect 21100 31900 21140 31940
rect 20812 31648 20852 31688
rect 19852 31312 19892 31352
rect 20044 31144 20084 31184
rect 20048 30976 20088 31016
rect 20130 30976 20170 31016
rect 20212 30976 20252 31016
rect 20294 30976 20334 31016
rect 20376 30976 20416 31016
rect 19852 30724 19892 30764
rect 20044 30556 20084 30596
rect 19756 30136 19796 30176
rect 19756 29884 19796 29924
rect 19660 29548 19700 29588
rect 19564 29044 19604 29084
rect 18808 28708 18848 28748
rect 18890 28708 18930 28748
rect 18972 28708 19012 28748
rect 19054 28708 19094 28748
rect 19136 28708 19176 28748
rect 18796 28540 18836 28580
rect 18316 27532 18356 27572
rect 17932 26356 17972 26396
rect 17932 26020 17972 26060
rect 18316 26608 18356 26648
rect 18412 26524 18452 26564
rect 18220 26440 18260 26480
rect 18028 25264 18068 25304
rect 17644 23920 17684 23960
rect 17932 23836 17972 23876
rect 18316 26356 18356 26396
rect 18316 25432 18356 25472
rect 18220 24508 18260 24548
rect 18124 23920 18164 23960
rect 17740 23416 17780 23456
rect 17452 22492 17492 22532
rect 17452 22240 17492 22280
rect 17452 21568 17492 21608
rect 17548 21400 17588 21440
rect 17548 21232 17588 21272
rect 17164 20644 17204 20684
rect 17068 20392 17108 20432
rect 17644 20728 17684 20768
rect 17644 20308 17684 20348
rect 17260 20224 17300 20264
rect 17548 20224 17588 20264
rect 16780 19720 16820 19760
rect 17068 19720 17108 19760
rect 16588 19552 16628 19592
rect 16492 19216 16532 19256
rect 17548 19384 17588 19424
rect 17164 19216 17204 19256
rect 16588 19048 16628 19088
rect 17068 19048 17108 19088
rect 16972 18376 17012 18416
rect 16684 17956 16724 17996
rect 16780 17872 16820 17912
rect 16684 17032 16724 17072
rect 16492 16612 16532 16652
rect 16300 16360 16340 16400
rect 16492 16360 16532 16400
rect 16204 16276 16244 16316
rect 16492 16192 16532 16232
rect 16684 16360 16724 16400
rect 16684 16192 16724 16232
rect 16588 16024 16628 16064
rect 16204 15940 16244 15980
rect 16204 15520 16244 15560
rect 16684 15604 16724 15644
rect 16588 15520 16628 15560
rect 16300 15436 16340 15476
rect 16300 15100 16340 15140
rect 16204 14932 16244 14972
rect 16876 16612 16916 16652
rect 16876 16192 16916 16232
rect 16780 15436 16820 15476
rect 16684 15184 16724 15224
rect 17452 18880 17492 18920
rect 17452 18628 17492 18668
rect 17260 18292 17300 18332
rect 17164 17704 17204 17744
rect 17740 20056 17780 20096
rect 17740 18964 17780 19004
rect 17740 18628 17780 18668
rect 17836 18544 17876 18584
rect 17644 17284 17684 17324
rect 17164 17032 17204 17072
rect 17068 16360 17108 16400
rect 16684 14512 16724 14552
rect 16972 14512 17012 14552
rect 16108 13420 16148 13460
rect 16108 12412 16148 12452
rect 15820 12160 15860 12200
rect 15724 11740 15764 11780
rect 15724 11236 15764 11276
rect 15724 10564 15764 10604
rect 15724 10228 15764 10268
rect 15532 9892 15572 9932
rect 15724 9808 15764 9848
rect 14860 9304 14900 9344
rect 14764 8632 14804 8672
rect 14956 9220 14996 9260
rect 14956 8968 14996 9008
rect 14956 8632 14996 8672
rect 15628 9220 15668 9260
rect 15340 8968 15380 9008
rect 15340 8632 15380 8672
rect 15148 8548 15188 8588
rect 15052 8464 15092 8504
rect 15436 8380 15476 8420
rect 16012 12160 16052 12200
rect 16012 10648 16052 10688
rect 16012 10228 16052 10268
rect 16012 9892 16052 9932
rect 15916 9808 15956 9848
rect 15729 8464 15769 8504
rect 15532 8128 15572 8168
rect 15532 7960 15572 8000
rect 15724 7624 15764 7664
rect 15148 6196 15188 6236
rect 15148 6028 15188 6068
rect 14956 5692 14996 5732
rect 14572 5020 14612 5060
rect 14668 4348 14708 4388
rect 14188 3424 14228 3464
rect 13804 2164 13844 2204
rect 13804 1828 13844 1868
rect 14188 2668 14228 2708
rect 14092 2164 14132 2204
rect 14380 1912 14420 1952
rect 14188 1744 14228 1784
rect 13996 1324 14036 1364
rect 15244 5272 15284 5312
rect 15052 4936 15092 4976
rect 14956 4684 14996 4724
rect 15148 4096 15188 4136
rect 15916 7960 15956 8000
rect 15916 7624 15956 7664
rect 15820 6700 15860 6740
rect 15628 6280 15668 6320
rect 15916 6448 15956 6488
rect 15436 6196 15476 6236
rect 15628 5776 15668 5816
rect 15628 5608 15668 5648
rect 15628 5272 15668 5312
rect 15532 5188 15572 5228
rect 15436 4936 15476 4976
rect 15436 3760 15476 3800
rect 15340 3676 15380 3716
rect 15436 3172 15476 3212
rect 15340 2752 15380 2792
rect 14860 2584 14900 2624
rect 14860 2416 14900 2456
rect 14572 1492 14612 1532
rect 15244 2332 15284 2372
rect 14956 2164 14996 2204
rect 14956 1912 14996 1952
rect 14860 1576 14900 1616
rect 13516 988 13556 1028
rect 13420 820 13460 860
rect 13324 568 13364 608
rect 13132 484 13172 524
rect 12940 400 12980 440
rect 14284 820 14324 860
rect 14476 820 14516 860
rect 13708 736 13748 776
rect 14092 316 14132 356
rect 13900 232 13940 272
rect 14860 1156 14900 1196
rect 14860 904 14900 944
rect 15340 904 15380 944
rect 15916 4348 15956 4388
rect 15916 4096 15956 4136
rect 15724 3760 15764 3800
rect 15820 3172 15860 3212
rect 16684 13924 16724 13964
rect 16588 13252 16628 13292
rect 16492 13084 16532 13124
rect 16780 13168 16820 13208
rect 17548 16612 17588 16652
rect 17740 16444 17780 16484
rect 17356 16276 17396 16316
rect 17740 16276 17780 16316
rect 17836 16192 17876 16232
rect 17452 15688 17492 15728
rect 18124 20980 18164 21020
rect 18028 20896 18068 20936
rect 18028 20728 18068 20768
rect 18508 26104 18548 26144
rect 18508 24844 18548 24884
rect 20236 30388 20276 30428
rect 19948 29632 19988 29672
rect 20048 29464 20088 29504
rect 20130 29464 20170 29504
rect 20212 29464 20252 29504
rect 20294 29464 20334 29504
rect 20376 29464 20416 29504
rect 19948 29296 19988 29336
rect 20812 29632 20852 29672
rect 19852 28540 19892 28580
rect 19276 28120 19316 28160
rect 19180 27868 19220 27908
rect 19468 27700 19508 27740
rect 18988 27616 19028 27656
rect 19660 28120 19700 28160
rect 19756 28036 19796 28076
rect 19756 27868 19796 27908
rect 19660 27700 19700 27740
rect 18808 27196 18848 27236
rect 18890 27196 18930 27236
rect 18972 27196 19012 27236
rect 19054 27196 19094 27236
rect 19136 27196 19176 27236
rect 18700 26356 18740 26396
rect 19564 26356 19604 26396
rect 18796 26104 18836 26144
rect 18412 24592 18452 24632
rect 18316 23920 18356 23960
rect 18316 23752 18356 23792
rect 18316 23080 18356 23120
rect 18808 25684 18848 25724
rect 18890 25684 18930 25724
rect 18972 25684 19012 25724
rect 19054 25684 19094 25724
rect 19136 25684 19176 25724
rect 19372 25684 19412 25724
rect 19180 25432 19220 25472
rect 18796 25180 18836 25220
rect 19372 25096 19412 25136
rect 18796 24592 18836 24632
rect 18988 24508 19028 24548
rect 20048 27952 20088 27992
rect 20130 27952 20170 27992
rect 20212 27952 20252 27992
rect 20294 27952 20334 27992
rect 20376 27952 20416 27992
rect 19948 26692 19988 26732
rect 20044 26608 20084 26648
rect 20048 26440 20088 26480
rect 20130 26440 20170 26480
rect 20212 26440 20252 26480
rect 20294 26440 20334 26480
rect 20376 26440 20416 26480
rect 19852 26272 19892 26312
rect 19756 26188 19796 26228
rect 19660 25348 19700 25388
rect 19564 25012 19604 25052
rect 19852 25432 19892 25472
rect 19852 24928 19892 24968
rect 19180 24340 19220 24380
rect 18508 23752 18548 23792
rect 18028 20308 18068 20348
rect 18028 19216 18068 19256
rect 18028 17536 18068 17576
rect 17932 15688 17972 15728
rect 17260 15520 17300 15560
rect 17836 15016 17876 15056
rect 17740 14428 17780 14468
rect 17644 14092 17684 14132
rect 17260 14008 17300 14048
rect 17164 13924 17204 13964
rect 17068 13840 17108 13880
rect 16972 13588 17012 13628
rect 16972 13336 17012 13376
rect 17356 13252 17396 13292
rect 17068 12832 17108 12872
rect 17356 12832 17396 12872
rect 17452 12496 17492 12536
rect 17836 13000 17876 13040
rect 17356 12412 17396 12452
rect 16780 11992 16820 12032
rect 16876 11908 16916 11948
rect 16300 11656 16340 11696
rect 16780 11656 16820 11696
rect 16204 8296 16244 8336
rect 16204 8128 16244 8168
rect 16684 10648 16724 10688
rect 16492 9892 16532 9932
rect 16396 9724 16436 9764
rect 16300 7624 16340 7664
rect 17740 11572 17780 11612
rect 16876 11488 16916 11528
rect 16684 7540 16724 7580
rect 18220 20056 18260 20096
rect 18412 22492 18452 22532
rect 18808 24172 18848 24212
rect 18890 24172 18930 24212
rect 18972 24172 19012 24212
rect 19054 24172 19094 24212
rect 19136 24172 19176 24212
rect 20908 29044 20948 29084
rect 20716 28120 20756 28160
rect 20620 27280 20660 27320
rect 20812 27784 20852 27824
rect 20908 27616 20948 27656
rect 21292 30388 21332 30428
rect 21196 29632 21236 29672
rect 21196 28540 21236 28580
rect 21100 27952 21140 27992
rect 21004 26944 21044 26984
rect 20812 26608 20852 26648
rect 20716 25936 20756 25976
rect 20524 25600 20564 25640
rect 20812 25432 20852 25472
rect 20044 25096 20084 25136
rect 20048 24928 20088 24968
rect 20130 24928 20170 24968
rect 20212 24928 20252 24968
rect 20294 24928 20334 24968
rect 20376 24928 20416 24968
rect 20524 24592 20564 24632
rect 18892 23752 18932 23792
rect 19276 23248 19316 23288
rect 18808 22660 18848 22700
rect 18890 22660 18930 22700
rect 18972 22660 19012 22700
rect 19054 22660 19094 22700
rect 19136 22660 19176 22700
rect 19372 22156 19412 22196
rect 18700 21652 18740 21692
rect 18988 21736 19028 21776
rect 18508 21400 18548 21440
rect 18796 21400 18836 21440
rect 18412 20896 18452 20936
rect 18316 18880 18356 18920
rect 18316 18460 18356 18500
rect 18316 18124 18356 18164
rect 18220 17788 18260 17828
rect 19660 23584 19700 23624
rect 19564 23248 19604 23288
rect 19564 22492 19604 22532
rect 20044 23668 20084 23708
rect 19948 23584 19988 23624
rect 20048 23416 20088 23456
rect 20130 23416 20170 23456
rect 20212 23416 20252 23456
rect 20294 23416 20334 23456
rect 20376 23416 20416 23456
rect 20044 23248 20084 23288
rect 19948 22996 19988 23036
rect 19852 22912 19892 22952
rect 19756 22576 19796 22616
rect 19660 22408 19700 22448
rect 20140 22492 20180 22532
rect 19564 22072 19604 22112
rect 20048 21904 20088 21944
rect 20130 21904 20170 21944
rect 20212 21904 20252 21944
rect 20294 21904 20334 21944
rect 20376 21904 20416 21944
rect 19468 21652 19508 21692
rect 19372 21484 19412 21524
rect 19084 21316 19124 21356
rect 18808 21148 18848 21188
rect 18890 21148 18930 21188
rect 18972 21148 19012 21188
rect 19054 21148 19094 21188
rect 19136 21148 19176 21188
rect 18604 20896 18644 20936
rect 19276 20896 19316 20936
rect 18508 20728 18548 20768
rect 19564 21400 19604 21440
rect 19276 20560 19316 20600
rect 19660 20308 19700 20348
rect 19468 20056 19508 20096
rect 18808 19636 18848 19676
rect 18890 19636 18930 19676
rect 18972 19636 19012 19676
rect 19054 19636 19094 19676
rect 19136 19636 19176 19676
rect 19564 19552 19604 19592
rect 18988 19468 19028 19508
rect 19852 20812 19892 20852
rect 20908 22492 20948 22532
rect 20908 21568 20948 21608
rect 19852 20560 19892 20600
rect 19372 19300 19412 19340
rect 18796 19216 18836 19256
rect 18700 19132 18740 19172
rect 18796 18544 18836 18584
rect 20812 20560 20852 20600
rect 20048 20392 20088 20432
rect 20130 20392 20170 20432
rect 20212 20392 20252 20432
rect 20294 20392 20334 20432
rect 20376 20392 20416 20432
rect 21292 22576 21332 22616
rect 21100 21400 21140 21440
rect 20044 19888 20084 19928
rect 20620 19216 20660 19256
rect 19756 19132 19796 19172
rect 19180 18292 19220 18332
rect 18808 18124 18848 18164
rect 18890 18124 18930 18164
rect 18972 18124 19012 18164
rect 19054 18124 19094 18164
rect 19136 18124 19176 18164
rect 18796 17956 18836 17996
rect 18508 17872 18548 17912
rect 18508 17704 18548 17744
rect 18316 17116 18356 17156
rect 18316 16948 18356 16988
rect 18220 16612 18260 16652
rect 18316 16192 18356 16232
rect 19084 17872 19124 17912
rect 19948 19048 19988 19088
rect 20048 18880 20088 18920
rect 20130 18880 20170 18920
rect 20212 18880 20252 18920
rect 20294 18880 20334 18920
rect 20376 18880 20416 18920
rect 19852 18544 19892 18584
rect 19468 17704 19508 17744
rect 19276 17200 19316 17240
rect 18796 16780 18836 16820
rect 18808 16612 18848 16652
rect 18890 16612 18930 16652
rect 18972 16612 19012 16652
rect 19054 16612 19094 16652
rect 19136 16612 19176 16652
rect 19660 17620 19700 17660
rect 20044 18040 20084 18080
rect 20236 17872 20276 17912
rect 20524 17704 20564 17744
rect 19948 17620 19988 17660
rect 19948 17368 19988 17408
rect 20048 17368 20088 17408
rect 20130 17368 20170 17408
rect 20212 17368 20252 17408
rect 20294 17368 20334 17408
rect 20376 17368 20416 17408
rect 19852 17200 19892 17240
rect 20236 16864 20276 16904
rect 19372 16024 19412 16064
rect 19084 15688 19124 15728
rect 18220 15352 18260 15392
rect 18988 15604 19028 15644
rect 19660 16108 19700 16148
rect 19564 15520 19604 15560
rect 19084 15436 19124 15476
rect 18604 15100 18644 15140
rect 18808 15100 18848 15140
rect 18890 15100 18930 15140
rect 18972 15100 19012 15140
rect 19054 15100 19094 15140
rect 19136 15100 19176 15140
rect 18508 14932 18548 14972
rect 19564 15184 19604 15224
rect 19084 14932 19124 14972
rect 19372 14932 19412 14972
rect 18412 14428 18452 14468
rect 18412 14176 18452 14216
rect 18604 14596 18644 14636
rect 18604 14428 18644 14468
rect 18700 14344 18740 14384
rect 19468 14680 19508 14720
rect 19852 16024 19892 16064
rect 20140 16024 20180 16064
rect 19852 15688 19892 15728
rect 19852 15436 19892 15476
rect 20048 15856 20088 15896
rect 20130 15856 20170 15896
rect 20212 15856 20252 15896
rect 20294 15856 20334 15896
rect 20376 15856 20416 15896
rect 21292 18796 21332 18836
rect 21100 17200 21140 17240
rect 20908 16528 20948 16568
rect 20044 15184 20084 15224
rect 20140 14932 20180 14972
rect 20236 14512 20276 14552
rect 20048 14344 20088 14384
rect 20130 14344 20170 14384
rect 20212 14344 20252 14384
rect 20294 14344 20334 14384
rect 20376 14344 20416 14384
rect 19948 14176 19988 14216
rect 19564 14092 19604 14132
rect 20140 14092 20180 14132
rect 18892 14008 18932 14048
rect 19948 14008 19988 14048
rect 18808 13588 18848 13628
rect 18890 13588 18930 13628
rect 18972 13588 19012 13628
rect 19054 13588 19094 13628
rect 19136 13588 19176 13628
rect 18220 13252 18260 13292
rect 18604 13168 18644 13208
rect 18124 13000 18164 13040
rect 17932 12160 17972 12200
rect 18220 12496 18260 12536
rect 18412 12244 18452 12284
rect 18124 11656 18164 11696
rect 17356 11068 17396 11108
rect 17356 10228 17396 10268
rect 17164 9472 17204 9512
rect 17068 9304 17108 9344
rect 17260 8968 17300 9008
rect 16972 8884 17012 8924
rect 17452 10144 17492 10184
rect 17740 11152 17780 11192
rect 18028 11068 18068 11108
rect 17836 10984 17876 11024
rect 17932 10900 17972 10940
rect 18028 10816 18068 10856
rect 18316 11572 18356 11612
rect 17932 10564 17972 10604
rect 18220 10480 18260 10520
rect 18124 10228 18164 10268
rect 18124 10060 18164 10100
rect 17740 9892 17780 9932
rect 17740 9640 17780 9680
rect 17644 9556 17684 9596
rect 18028 9556 18068 9596
rect 17548 9472 17588 9512
rect 17452 9304 17492 9344
rect 17644 9304 17684 9344
rect 17740 9220 17780 9260
rect 17452 8632 17492 8672
rect 17644 7960 17684 8000
rect 16876 7792 16916 7832
rect 16972 7708 17012 7748
rect 16396 7036 16436 7076
rect 16204 6196 16244 6236
rect 16588 6196 16628 6236
rect 16396 5944 16436 5984
rect 16300 5692 16340 5732
rect 16300 5524 16340 5564
rect 16492 5188 16532 5228
rect 16300 4936 16340 4976
rect 16204 4600 16244 4640
rect 16300 4348 16340 4388
rect 16684 5692 16724 5732
rect 16684 5272 16724 5312
rect 16876 6280 16916 6320
rect 17068 6448 17108 6488
rect 17068 6196 17108 6236
rect 16780 5188 16820 5228
rect 16972 5608 17012 5648
rect 17932 8632 17972 8672
rect 17836 8548 17876 8588
rect 18124 8296 18164 8336
rect 18028 8212 18068 8252
rect 19564 13168 19604 13208
rect 18988 12412 19028 12452
rect 18700 12160 18740 12200
rect 18808 12076 18848 12116
rect 18890 12076 18930 12116
rect 18972 12076 19012 12116
rect 19054 12076 19094 12116
rect 19136 12076 19176 12116
rect 18700 11824 18740 11864
rect 19084 11656 19124 11696
rect 19276 11656 19316 11696
rect 19564 12496 19604 12536
rect 20048 12832 20088 12872
rect 20130 12832 20170 12872
rect 20212 12832 20252 12872
rect 20294 12832 20334 12872
rect 20376 12832 20416 12872
rect 19660 12412 19700 12452
rect 19948 12412 19988 12452
rect 19660 11992 19700 12032
rect 18700 11572 18740 11612
rect 19756 11656 19796 11696
rect 19468 11152 19508 11192
rect 20044 11656 20084 11696
rect 20048 11320 20088 11360
rect 20130 11320 20170 11360
rect 20212 11320 20252 11360
rect 20294 11320 20334 11360
rect 20376 11320 20416 11360
rect 20044 11152 20084 11192
rect 19948 11068 19988 11108
rect 18796 10900 18836 10940
rect 18508 10816 18548 10856
rect 18508 10564 18548 10604
rect 18412 10228 18452 10268
rect 18508 9388 18548 9428
rect 18808 10564 18848 10604
rect 18890 10564 18930 10604
rect 18972 10564 19012 10604
rect 19054 10564 19094 10604
rect 19136 10564 19176 10604
rect 19852 11019 19892 11024
rect 19852 10984 19892 11019
rect 19084 10312 19124 10352
rect 18700 10144 18740 10184
rect 18892 10060 18932 10100
rect 19084 9472 19124 9512
rect 18604 8968 18644 9008
rect 18316 8548 18356 8588
rect 18508 7960 18548 8000
rect 17836 6448 17876 6488
rect 18316 7372 18356 7412
rect 18412 6700 18452 6740
rect 17932 6364 17972 6404
rect 17740 6196 17780 6236
rect 17644 5776 17684 5816
rect 17356 5692 17396 5732
rect 17260 5608 17300 5648
rect 18028 6280 18068 6320
rect 18028 5944 18068 5984
rect 17644 5608 17684 5648
rect 17932 5524 17972 5564
rect 17068 4936 17108 4976
rect 17164 4852 17204 4892
rect 17644 5020 17684 5060
rect 17740 4936 17780 4976
rect 17932 4936 17972 4976
rect 17356 4600 17396 4640
rect 16684 4264 16724 4304
rect 16684 4096 16724 4136
rect 16972 4096 17012 4136
rect 17260 4096 17300 4136
rect 16204 3676 16244 3716
rect 16876 3676 16916 3716
rect 16300 3256 16340 3296
rect 15820 2752 15860 2792
rect 15724 2584 15764 2624
rect 15532 1156 15572 1196
rect 15724 2248 15764 2288
rect 16780 3256 16820 3296
rect 16588 3004 16628 3044
rect 16492 2920 16532 2960
rect 16492 2752 16532 2792
rect 16012 2584 16052 2624
rect 16012 1660 16052 1700
rect 16684 2584 16724 2624
rect 16588 2500 16628 2540
rect 16492 2416 16532 2456
rect 16396 1912 16436 1952
rect 16588 2332 16628 2372
rect 16204 1408 16244 1448
rect 16108 736 16148 776
rect 16492 1744 16532 1784
rect 16396 1156 16436 1196
rect 16396 988 16436 1028
rect 16780 1828 16820 1868
rect 17932 4684 17972 4724
rect 17740 4096 17780 4136
rect 17068 3676 17108 3716
rect 16972 3424 17012 3464
rect 17356 3676 17396 3716
rect 17356 3256 17396 3296
rect 16972 2584 17012 2624
rect 17260 2584 17300 2624
rect 17644 3424 17684 3464
rect 18412 5776 18452 5816
rect 18316 5440 18356 5480
rect 18808 9052 18848 9092
rect 18890 9052 18930 9092
rect 18972 9052 19012 9092
rect 19054 9052 19094 9092
rect 19136 9052 19176 9092
rect 19084 8632 19124 8672
rect 19564 10060 19604 10100
rect 19948 10060 19988 10100
rect 20048 9808 20088 9848
rect 20130 9808 20170 9848
rect 20212 9808 20252 9848
rect 20294 9808 20334 9848
rect 20376 9808 20416 9848
rect 19852 9472 19892 9512
rect 20236 9640 20276 9680
rect 19564 8884 19604 8924
rect 20044 8968 20084 9008
rect 20620 13504 20660 13544
rect 19948 8716 19988 8756
rect 20048 8296 20088 8336
rect 20130 8296 20170 8336
rect 20212 8296 20252 8336
rect 20294 8296 20334 8336
rect 20376 8296 20416 8336
rect 19276 8128 19316 8168
rect 19084 8044 19124 8084
rect 19084 7708 19124 7748
rect 18808 7540 18848 7580
rect 18890 7540 18930 7580
rect 18972 7540 19012 7580
rect 19054 7540 19094 7580
rect 19136 7540 19176 7580
rect 18988 6700 19028 6740
rect 18796 6616 18836 6656
rect 18700 6364 18740 6404
rect 18892 6532 18932 6572
rect 19372 7960 19412 8000
rect 19564 8044 19604 8084
rect 18988 6364 19028 6404
rect 18892 6196 18932 6236
rect 18604 4684 18644 4724
rect 18412 4600 18452 4640
rect 18124 4096 18164 4136
rect 18028 3928 18068 3968
rect 18028 3592 18068 3632
rect 17452 2752 17492 2792
rect 16972 2164 17012 2204
rect 17260 2164 17300 2204
rect 17164 1912 17204 1952
rect 17260 1744 17300 1784
rect 16684 1324 16724 1364
rect 16972 1324 17012 1364
rect 17260 1324 17300 1364
rect 18412 3508 18452 3548
rect 18124 3424 18164 3464
rect 18220 3004 18260 3044
rect 18124 2920 18164 2960
rect 18028 2164 18068 2204
rect 16780 1240 16820 1280
rect 16684 484 16724 524
rect 17548 1240 17588 1280
rect 17164 1072 17204 1112
rect 17452 820 17492 860
rect 17164 736 17204 776
rect 17356 484 17396 524
rect 18124 1912 18164 1952
rect 18316 2836 18356 2876
rect 17932 1492 17972 1532
rect 17644 1072 17684 1112
rect 17740 904 17780 944
rect 18808 6028 18848 6068
rect 18890 6028 18930 6068
rect 18972 6028 19012 6068
rect 19054 6028 19094 6068
rect 19136 6028 19176 6068
rect 19084 4936 19124 4976
rect 18808 4516 18848 4556
rect 18890 4516 18930 4556
rect 18972 4516 19012 4556
rect 19054 4516 19094 4556
rect 19136 4516 19176 4556
rect 20524 7960 20564 8000
rect 20048 6784 20088 6824
rect 20130 6784 20170 6824
rect 20212 6784 20252 6824
rect 20294 6784 20334 6824
rect 20376 6784 20416 6824
rect 19852 6483 19892 6488
rect 19852 6448 19892 6483
rect 19660 6196 19700 6236
rect 19468 4936 19508 4976
rect 19372 4516 19412 4556
rect 18796 4348 18836 4388
rect 20236 6280 20276 6320
rect 21388 15352 21428 15392
rect 21292 11152 21332 11192
rect 21388 7792 21428 7832
rect 20620 6952 20660 6992
rect 19660 5440 19700 5480
rect 19084 4180 19124 4220
rect 19660 4180 19700 4220
rect 19564 4096 19604 4136
rect 19468 4012 19508 4052
rect 20048 5272 20088 5312
rect 20130 5272 20170 5312
rect 20212 5272 20252 5312
rect 20294 5272 20334 5312
rect 20376 5272 20416 5312
rect 20236 4936 20276 4976
rect 19948 4684 19988 4724
rect 20048 3760 20088 3800
rect 20130 3760 20170 3800
rect 20212 3760 20252 3800
rect 20294 3760 20334 3800
rect 20376 3760 20416 3800
rect 18604 2836 18644 2876
rect 19276 3088 19316 3128
rect 18808 3004 18848 3044
rect 18890 3004 18930 3044
rect 18972 3004 19012 3044
rect 19054 3004 19094 3044
rect 19136 3004 19176 3044
rect 18508 2668 18548 2708
rect 18604 2584 18644 2624
rect 19180 2668 19220 2708
rect 19372 2584 19412 2624
rect 18508 2164 18548 2204
rect 19276 1576 19316 1616
rect 18808 1492 18848 1532
rect 18890 1492 18930 1532
rect 18972 1492 19012 1532
rect 19054 1492 19094 1532
rect 19136 1492 19176 1532
rect 18700 1240 18740 1280
rect 18124 904 18164 944
rect 18508 568 18548 608
rect 18892 904 18932 944
rect 19084 232 19124 272
rect 19660 3256 19700 3296
rect 19564 2668 19604 2708
rect 19468 1408 19508 1448
rect 19468 1240 19508 1280
rect 19756 2584 19796 2624
rect 19852 2500 19892 2540
rect 20048 2248 20088 2288
rect 20130 2248 20170 2288
rect 20212 2248 20252 2288
rect 20294 2248 20334 2288
rect 20376 2248 20416 2288
rect 19948 1996 19988 2036
rect 19372 988 19412 1028
rect 19948 1408 19988 1448
rect 19660 988 19700 1028
rect 20048 736 20088 776
rect 20130 736 20170 776
rect 20212 736 20252 776
rect 20294 736 20334 776
rect 20376 736 20416 776
<< metal3 >>
rect 2563 42820 2572 42860
rect 2612 42820 13612 42860
rect 13652 42820 13661 42860
rect 20611 42776 20669 42777
rect 21424 42776 21504 42796
rect 20611 42736 20620 42776
rect 20660 42736 21504 42776
rect 20611 42735 20669 42736
rect 21424 42716 21504 42736
rect 4099 42608 4157 42609
rect 11779 42608 11837 42609
rect 4099 42568 4108 42608
rect 4148 42568 6220 42608
rect 6260 42568 6269 42608
rect 11694 42568 11788 42608
rect 11828 42568 11837 42608
rect 4099 42567 4157 42568
rect 11779 42567 11837 42568
rect 14659 42608 14717 42609
rect 14659 42568 14668 42608
rect 14708 42568 17356 42608
rect 17396 42568 17405 42608
rect 14659 42567 14717 42568
rect 1699 42484 1708 42524
rect 1748 42484 4876 42524
rect 4916 42484 4925 42524
rect 14563 42484 14572 42524
rect 14612 42484 19468 42524
rect 19508 42484 19517 42524
rect 21424 42440 21504 42460
rect 13027 42400 13036 42440
rect 13076 42400 21504 42440
rect 21424 42380 21504 42400
rect 17347 42316 17356 42356
rect 17396 42316 20180 42356
rect 1891 42272 1949 42273
rect 1891 42232 1900 42272
rect 1940 42232 4108 42272
rect 4148 42232 4157 42272
rect 15427 42232 15436 42272
rect 15476 42232 17836 42272
rect 17876 42232 17885 42272
rect 1891 42231 1949 42232
rect 18691 42188 18749 42189
rect 3907 42148 3916 42188
rect 3956 42148 16300 42188
rect 16340 42148 16349 42188
rect 16579 42148 16588 42188
rect 16628 42148 18220 42188
rect 18260 42148 18269 42188
rect 18606 42148 18700 42188
rect 18740 42148 18749 42188
rect 18691 42147 18749 42148
rect 1507 42104 1565 42105
rect 20140 42104 20180 42316
rect 21424 42104 21504 42124
rect 1507 42064 1516 42104
rect 1556 42064 4492 42104
rect 4532 42064 4541 42104
rect 13699 42064 13708 42104
rect 13748 42064 15436 42104
rect 15476 42064 15485 42104
rect 15811 42064 15820 42104
rect 15860 42064 18604 42104
rect 18644 42064 18653 42104
rect 18883 42064 18892 42104
rect 18932 42064 19468 42104
rect 19508 42064 19517 42104
rect 20140 42064 21504 42104
rect 1507 42063 1565 42064
rect 21424 42044 21504 42064
rect 18115 41980 18124 42020
rect 18164 41980 19852 42020
rect 19892 41980 19901 42020
rect 5251 41896 5260 41936
rect 5300 41896 5644 41936
rect 5684 41896 5693 41936
rect 16003 41896 16012 41936
rect 16052 41896 18988 41936
rect 19028 41896 19037 41936
rect 17443 41812 17452 41852
rect 17492 41812 19084 41852
rect 19124 41812 19133 41852
rect 21424 41768 21504 41788
rect 4099 41728 4108 41768
rect 4148 41728 7372 41768
rect 7412 41728 7421 41768
rect 15043 41728 15052 41768
rect 15092 41728 16972 41768
rect 17012 41728 17021 41768
rect 20140 41728 21504 41768
rect 20140 41684 20180 41728
rect 21424 41708 21504 41728
rect 6211 41644 6220 41684
rect 6260 41644 7756 41684
rect 7796 41644 7805 41684
rect 14851 41644 14860 41684
rect 14900 41644 16588 41684
rect 16628 41644 16637 41684
rect 17539 41644 17548 41684
rect 17588 41644 18700 41684
rect 18740 41644 18749 41684
rect 18796 41644 20180 41684
rect 9859 41600 9917 41601
rect 4919 41560 4928 41600
rect 4968 41560 5010 41600
rect 5050 41560 5092 41600
rect 5132 41560 5174 41600
rect 5214 41560 5256 41600
rect 5296 41560 5305 41600
rect 9774 41560 9868 41600
rect 9908 41560 9917 41600
rect 9859 41559 9917 41560
rect 10051 41600 10109 41601
rect 11395 41600 11453 41601
rect 11587 41600 11645 41601
rect 17923 41600 17981 41601
rect 18499 41600 18557 41601
rect 18796 41600 18836 41644
rect 10051 41560 10060 41600
rect 10100 41560 10194 41600
rect 11395 41560 11404 41600
rect 11444 41560 11538 41600
rect 11587 41560 11596 41600
rect 11636 41560 11730 41600
rect 13507 41560 13516 41600
rect 13556 41560 14668 41600
rect 14708 41560 14717 41600
rect 16387 41560 16396 41600
rect 16436 41560 17740 41600
rect 17780 41560 17789 41600
rect 17923 41560 17932 41600
rect 17972 41560 18066 41600
rect 18414 41560 18508 41600
rect 18548 41560 18557 41600
rect 10051 41559 10109 41560
rect 11395 41559 11453 41560
rect 11587 41559 11645 41560
rect 17923 41559 17981 41560
rect 18499 41559 18557 41560
rect 18604 41560 18836 41600
rect 20039 41560 20048 41600
rect 20088 41560 20130 41600
rect 20170 41560 20212 41600
rect 20252 41560 20294 41600
rect 20334 41560 20376 41600
rect 20416 41560 20425 41600
rect 18604 41516 18644 41560
rect 16483 41476 16492 41516
rect 16532 41476 18644 41516
rect 20803 41432 20861 41433
rect 21424 41432 21504 41452
rect 11299 41392 11308 41432
rect 11348 41392 12172 41432
rect 12212 41392 12221 41432
rect 16291 41392 16300 41432
rect 16340 41392 19372 41432
rect 19412 41392 19421 41432
rect 20803 41392 20812 41432
rect 20852 41392 21504 41432
rect 20803 41391 20861 41392
rect 21424 41372 21504 41392
rect 11596 41308 12460 41348
rect 12500 41308 18796 41348
rect 18836 41308 18845 41348
rect 1795 41264 1853 41265
rect 1710 41224 1804 41264
rect 1844 41224 1853 41264
rect 1795 41223 1853 41224
rect 2755 41264 2813 41265
rect 11596 41264 11636 41308
rect 16675 41264 16733 41265
rect 2755 41224 2764 41264
rect 2804 41224 3436 41264
rect 3476 41224 7564 41264
rect 7604 41224 7613 41264
rect 9379 41224 9388 41264
rect 9428 41224 9964 41264
rect 10004 41224 11596 41264
rect 11636 41224 11645 41264
rect 12163 41224 12172 41264
rect 12212 41224 13804 41264
rect 13844 41224 13853 41264
rect 14467 41224 14476 41264
rect 14516 41224 16244 41264
rect 16590 41224 16684 41264
rect 16724 41224 16733 41264
rect 2755 41223 2813 41224
rect 7564 41096 7604 41224
rect 8035 41180 8093 41181
rect 16204 41180 16244 41224
rect 16675 41223 16733 41224
rect 19747 41180 19805 41181
rect 7950 41140 8044 41180
rect 8084 41140 8093 41180
rect 11395 41140 11404 41180
rect 11444 41140 11980 41180
rect 12020 41140 12029 41180
rect 14083 41140 14092 41180
rect 14132 41140 15820 41180
rect 15860 41140 15869 41180
rect 16195 41140 16204 41180
rect 16244 41140 16253 41180
rect 19555 41140 19564 41180
rect 19604 41140 19756 41180
rect 19796 41140 19805 41180
rect 8035 41139 8093 41140
rect 19747 41139 19805 41140
rect 19843 41096 19901 41097
rect 21424 41096 21504 41116
rect 7564 41056 11596 41096
rect 11636 41056 11645 41096
rect 13891 41056 13900 41096
rect 13940 41056 15052 41096
rect 15092 41056 15101 41096
rect 15148 41056 15380 41096
rect 15523 41056 15532 41096
rect 15572 41056 19796 41096
rect 13315 41012 13373 41013
rect 15148 41012 15188 41056
rect 1411 40972 1420 41012
rect 1460 40972 3724 41012
rect 3764 40972 3773 41012
rect 5251 40972 5260 41012
rect 5300 40972 6124 41012
rect 6164 40972 6173 41012
rect 12643 40972 12652 41012
rect 12692 40972 12940 41012
rect 12980 40972 12989 41012
rect 13315 40972 13324 41012
rect 13364 40972 15188 41012
rect 15340 41012 15380 41056
rect 15619 41012 15677 41013
rect 16003 41012 16061 41013
rect 19756 41012 19796 41056
rect 19843 41056 19852 41096
rect 19892 41056 21504 41096
rect 19843 41055 19901 41056
rect 21424 41036 21504 41056
rect 15340 40972 15572 41012
rect 13315 40971 13373 40972
rect 15532 40928 15572 40972
rect 15619 40972 15628 41012
rect 15668 40972 15762 41012
rect 15918 40972 16012 41012
rect 16052 40972 16061 41012
rect 16483 40972 16492 41012
rect 16532 40972 19180 41012
rect 19220 40972 19229 41012
rect 19747 40972 19756 41012
rect 19796 40972 19805 41012
rect 15619 40971 15677 40972
rect 16003 40971 16061 40972
rect 2275 40888 2284 40928
rect 2324 40888 4300 40928
rect 4340 40888 4349 40928
rect 14275 40888 14284 40928
rect 14324 40888 15436 40928
rect 15476 40888 15485 40928
rect 15532 40888 18316 40928
rect 18356 40888 18508 40928
rect 18548 40888 18557 40928
rect 3043 40844 3101 40845
rect 4195 40844 4253 40845
rect 17635 40844 17693 40845
rect 2958 40804 3052 40844
rect 3092 40804 3101 40844
rect 3679 40804 3688 40844
rect 3728 40804 3770 40844
rect 3810 40804 3852 40844
rect 3892 40804 3934 40844
rect 3974 40804 4016 40844
rect 4056 40804 4065 40844
rect 4195 40804 4204 40844
rect 4244 40804 5548 40844
rect 5588 40804 5597 40844
rect 10051 40804 10060 40844
rect 10100 40804 10444 40844
rect 10484 40804 10493 40844
rect 14179 40804 14188 40844
rect 14228 40804 17396 40844
rect 17550 40804 17644 40844
rect 17684 40804 17693 40844
rect 18799 40804 18808 40844
rect 18848 40804 18890 40844
rect 18930 40804 18972 40844
rect 19012 40804 19054 40844
rect 19094 40804 19136 40844
rect 19176 40804 19185 40844
rect 3043 40803 3101 40804
rect 4195 40803 4253 40804
rect 17356 40760 17396 40804
rect 17635 40803 17693 40804
rect 21424 40760 21504 40780
rect 2755 40720 2764 40760
rect 2804 40720 3532 40760
rect 3572 40720 3581 40760
rect 5347 40720 5356 40760
rect 5396 40720 6124 40760
rect 6164 40720 6173 40760
rect 7939 40720 7948 40760
rect 7988 40720 11360 40760
rect 17356 40720 19372 40760
rect 19412 40720 19421 40760
rect 19939 40720 19948 40760
rect 19988 40720 21504 40760
rect 10915 40676 10973 40677
rect 2083 40636 2092 40676
rect 2132 40636 8716 40676
rect 8756 40636 8765 40676
rect 10243 40636 10252 40676
rect 10292 40636 10444 40676
rect 10484 40636 10493 40676
rect 10830 40636 10924 40676
rect 10964 40636 10973 40676
rect 11320 40676 11360 40720
rect 21424 40700 21504 40720
rect 11320 40636 16532 40676
rect 17155 40636 17164 40676
rect 17204 40636 19084 40676
rect 19124 40636 19133 40676
rect 10915 40635 10973 40636
rect 3331 40592 3389 40593
rect 14083 40592 14141 40593
rect 14467 40592 14525 40593
rect 14851 40592 14909 40593
rect 1315 40552 1324 40592
rect 1364 40552 1516 40592
rect 1556 40552 3340 40592
rect 3380 40552 3389 40592
rect 3523 40552 3532 40592
rect 3572 40552 5740 40592
rect 5780 40552 5789 40592
rect 6403 40552 6412 40592
rect 6452 40552 7276 40592
rect 7316 40552 7325 40592
rect 8515 40552 8524 40592
rect 8564 40552 11360 40592
rect 13998 40552 14092 40592
rect 14132 40552 14141 40592
rect 14382 40552 14476 40592
rect 14516 40552 14525 40592
rect 14766 40552 14860 40592
rect 14900 40552 14909 40592
rect 3331 40551 3389 40552
rect 2947 40468 2956 40508
rect 2996 40468 3572 40508
rect 3619 40468 3628 40508
rect 3668 40468 6988 40508
rect 7028 40468 7037 40508
rect 9763 40468 9772 40508
rect 9812 40468 10540 40508
rect 10580 40468 10589 40508
rect 3532 40424 3572 40468
rect 5827 40424 5885 40425
rect 10819 40424 10877 40425
rect 2659 40384 2668 40424
rect 2708 40384 3148 40424
rect 3188 40384 3197 40424
rect 3532 40384 4684 40424
rect 4724 40384 5356 40424
rect 5396 40384 5405 40424
rect 5742 40384 5836 40424
rect 5876 40384 5885 40424
rect 6307 40384 6316 40424
rect 6356 40384 6700 40424
rect 6740 40384 7660 40424
rect 7700 40384 7709 40424
rect 10723 40384 10732 40424
rect 10772 40384 10828 40424
rect 10868 40384 10877 40424
rect 11320 40424 11360 40552
rect 14083 40551 14141 40552
rect 14467 40551 14525 40552
rect 14851 40551 14909 40552
rect 15139 40592 15197 40593
rect 15811 40592 15869 40593
rect 16387 40592 16445 40593
rect 15139 40552 15148 40592
rect 15188 40552 15244 40592
rect 15284 40552 15293 40592
rect 15811 40552 15820 40592
rect 15860 40552 16012 40592
rect 16052 40552 16061 40592
rect 16302 40552 16396 40592
rect 16436 40552 16445 40592
rect 16492 40592 16532 40636
rect 16492 40552 18700 40592
rect 18740 40552 18749 40592
rect 18796 40552 19700 40592
rect 15139 40551 15197 40552
rect 15811 40551 15869 40552
rect 16387 40551 16445 40552
rect 18796 40508 18836 40552
rect 19660 40509 19700 40552
rect 13315 40468 13324 40508
rect 13364 40468 14284 40508
rect 14324 40468 14333 40508
rect 14755 40468 14764 40508
rect 14804 40468 16204 40508
rect 16244 40468 16253 40508
rect 18019 40468 18028 40508
rect 18068 40468 18836 40508
rect 18883 40508 18941 40509
rect 19651 40508 19709 40509
rect 18883 40468 18892 40508
rect 18932 40468 19026 40508
rect 19566 40468 19660 40508
rect 19700 40468 19709 40508
rect 18883 40467 18941 40468
rect 19651 40467 19709 40468
rect 21424 40424 21504 40444
rect 11320 40384 15628 40424
rect 15668 40384 15677 40424
rect 15724 40384 17644 40424
rect 17684 40384 17693 40424
rect 17740 40384 21504 40424
rect 5827 40383 5885 40384
rect 10819 40383 10877 40384
rect 9763 40340 9821 40341
rect 14947 40340 15005 40341
rect 15235 40340 15293 40341
rect 3235 40300 3244 40340
rect 3284 40300 4012 40340
rect 4052 40300 4061 40340
rect 5539 40300 5548 40340
rect 5588 40300 6508 40340
rect 6548 40300 6557 40340
rect 9763 40300 9772 40340
rect 9812 40300 9906 40340
rect 11587 40300 11596 40340
rect 11636 40300 12212 40340
rect 13891 40300 13900 40340
rect 13940 40300 14956 40340
rect 14996 40300 15005 40340
rect 15139 40300 15148 40340
rect 15188 40300 15244 40340
rect 15284 40300 15293 40340
rect 9763 40299 9821 40300
rect 3043 40256 3101 40257
rect 10243 40256 10301 40257
rect 3043 40216 3052 40256
rect 3092 40216 3340 40256
rect 3380 40216 3389 40256
rect 9187 40216 9196 40256
rect 9236 40216 9676 40256
rect 9716 40216 9725 40256
rect 10158 40216 10252 40256
rect 10292 40216 10301 40256
rect 3043 40215 3101 40216
rect 10243 40215 10301 40216
rect 7747 40132 7756 40172
rect 7796 40132 10156 40172
rect 10196 40132 10205 40172
rect 10723 40132 10732 40172
rect 10772 40132 11020 40172
rect 11060 40132 11069 40172
rect 0 40088 80 40108
rect 3139 40088 3197 40089
rect 12172 40088 12212 40300
rect 14947 40299 15005 40300
rect 15235 40299 15293 40300
rect 15619 40340 15677 40341
rect 15724 40340 15764 40384
rect 15619 40300 15628 40340
rect 15668 40300 15764 40340
rect 17347 40340 17405 40341
rect 17740 40340 17780 40384
rect 21424 40364 21504 40384
rect 19843 40340 19901 40341
rect 17347 40300 17356 40340
rect 17396 40300 17780 40340
rect 17827 40300 17836 40340
rect 17876 40300 19852 40340
rect 19892 40300 19901 40340
rect 15619 40299 15677 40300
rect 17347 40299 17405 40300
rect 19843 40299 19901 40300
rect 18691 40256 18749 40257
rect 12259 40216 12268 40256
rect 12308 40216 12596 40256
rect 15331 40216 15340 40256
rect 15380 40216 17068 40256
rect 17108 40216 17117 40256
rect 18606 40216 18700 40256
rect 18740 40216 18749 40256
rect 12556 40172 12596 40216
rect 18691 40215 18749 40216
rect 12547 40132 12556 40172
rect 12596 40132 12605 40172
rect 14083 40132 14092 40172
rect 14132 40132 14956 40172
rect 14996 40132 19756 40172
rect 19796 40132 19805 40172
rect 17923 40088 17981 40089
rect 21424 40088 21504 40108
rect 0 40048 3148 40088
rect 3188 40048 3197 40088
rect 4919 40048 4928 40088
rect 4968 40048 5010 40088
rect 5050 40048 5092 40088
rect 5132 40048 5174 40088
rect 5214 40048 5256 40088
rect 5296 40048 5305 40088
rect 5539 40048 5548 40088
rect 5588 40048 5932 40088
rect 5972 40048 5981 40088
rect 7651 40048 7660 40088
rect 7700 40048 8236 40088
rect 8276 40048 8285 40088
rect 8611 40048 8620 40088
rect 8660 40048 12116 40088
rect 12163 40048 12172 40088
rect 12212 40048 12221 40088
rect 13411 40048 13420 40088
rect 13460 40048 13708 40088
rect 13748 40048 13757 40088
rect 17923 40048 17932 40088
rect 17972 40048 18988 40088
rect 19028 40048 19037 40088
rect 20039 40048 20048 40088
rect 20088 40048 20130 40088
rect 20170 40048 20212 40088
rect 20252 40048 20294 40088
rect 20334 40048 20376 40088
rect 20416 40048 20425 40088
rect 20812 40048 21504 40088
rect 0 40028 80 40048
rect 3139 40047 3197 40048
rect 12076 40004 12116 40048
rect 17923 40047 17981 40048
rect 20812 40004 20852 40048
rect 21424 40028 21504 40048
rect 2083 39964 2092 40004
rect 2132 39964 11788 40004
rect 11828 39964 11837 40004
rect 12076 39964 15532 40004
rect 15572 39964 15581 40004
rect 15628 39964 20852 40004
rect 15628 39920 15668 39964
rect 5251 39880 5260 39920
rect 5300 39880 5644 39920
rect 5684 39880 5693 39920
rect 9571 39880 9580 39920
rect 9620 39880 10924 39920
rect 10964 39880 10973 39920
rect 11320 39880 13612 39920
rect 13652 39880 13661 39920
rect 14275 39880 14284 39920
rect 14324 39880 15668 39920
rect 15715 39880 15724 39920
rect 15764 39880 17548 39920
rect 17588 39880 17597 39920
rect 18403 39880 18412 39920
rect 18452 39880 19180 39920
rect 19220 39880 19229 39920
rect 11320 39836 11360 39880
rect 17155 39836 17213 39837
rect 3331 39796 3340 39836
rect 3380 39796 3389 39836
rect 4963 39796 4972 39836
rect 5012 39796 11360 39836
rect 12739 39796 12748 39836
rect 12788 39796 13036 39836
rect 13076 39796 13085 39836
rect 14563 39796 14572 39836
rect 14612 39796 16492 39836
rect 16532 39796 16541 39836
rect 16675 39796 16684 39836
rect 16724 39796 17164 39836
rect 17204 39796 17213 39836
rect 1603 39752 1661 39753
rect 3340 39752 3380 39796
rect 17155 39795 17213 39796
rect 20803 39752 20861 39753
rect 21424 39752 21504 39772
rect 1603 39712 1612 39752
rect 1652 39712 1708 39752
rect 1748 39712 1757 39752
rect 3340 39712 5644 39752
rect 5684 39712 6316 39752
rect 6356 39712 6365 39752
rect 6412 39712 12308 39752
rect 12451 39712 12460 39752
rect 12500 39712 20812 39752
rect 20852 39712 20861 39752
rect 20995 39712 21004 39752
rect 21044 39712 21504 39752
rect 1603 39711 1661 39712
rect 6412 39668 6452 39712
rect 4099 39628 4108 39668
rect 4148 39628 4492 39668
rect 4532 39628 6452 39668
rect 10915 39668 10973 39669
rect 11107 39668 11165 39669
rect 10915 39628 10924 39668
rect 10964 39628 11116 39668
rect 11156 39628 11596 39668
rect 11636 39628 11645 39668
rect 10915 39627 10973 39628
rect 11107 39627 11165 39628
rect 0 39584 80 39604
rect 2467 39584 2525 39585
rect 0 39544 1420 39584
rect 1460 39544 1469 39584
rect 2467 39544 2476 39584
rect 2516 39544 4396 39584
rect 4436 39544 10252 39584
rect 10292 39544 11360 39584
rect 0 39524 80 39544
rect 2467 39543 2525 39544
rect 3811 39460 3820 39500
rect 3860 39460 4148 39500
rect 5827 39460 5836 39500
rect 5876 39460 7372 39500
rect 7412 39460 7421 39500
rect 8419 39460 8428 39500
rect 8468 39460 9388 39500
rect 9428 39460 9437 39500
rect 4108 39332 4148 39460
rect 11320 39416 11360 39544
rect 12268 39500 12308 39712
rect 20803 39711 20861 39712
rect 21424 39692 21504 39712
rect 12355 39628 12364 39668
rect 12404 39628 17740 39668
rect 17780 39628 17789 39668
rect 18019 39628 18028 39668
rect 18068 39628 18796 39668
rect 18836 39628 18845 39668
rect 19939 39628 19948 39668
rect 19988 39628 20028 39668
rect 12355 39584 12413 39585
rect 17251 39584 17309 39585
rect 19948 39584 19988 39628
rect 12355 39544 12364 39584
rect 12404 39544 17108 39584
rect 17166 39544 17260 39584
rect 17300 39544 17309 39584
rect 12355 39543 12413 39544
rect 16867 39500 16925 39501
rect 12268 39460 14092 39500
rect 14132 39460 14141 39500
rect 16782 39460 16876 39500
rect 16916 39460 16925 39500
rect 17068 39500 17108 39544
rect 17251 39543 17309 39544
rect 19468 39544 20140 39584
rect 20180 39544 20189 39584
rect 19468 39500 19508 39544
rect 17068 39460 19508 39500
rect 19555 39460 19564 39500
rect 19604 39460 20180 39500
rect 16867 39459 16925 39460
rect 20140 39416 20180 39460
rect 21424 39416 21504 39436
rect 4387 39376 4396 39416
rect 4436 39376 8044 39416
rect 8084 39376 8093 39416
rect 11320 39376 19372 39416
rect 19412 39376 19421 39416
rect 20140 39376 21504 39416
rect 21424 39356 21504 39376
rect 12931 39332 12989 39333
rect 3679 39292 3688 39332
rect 3728 39292 3770 39332
rect 3810 39292 3852 39332
rect 3892 39292 3934 39332
rect 3974 39292 4016 39332
rect 4056 39292 4065 39332
rect 4108 39292 12940 39332
rect 12980 39292 12989 39332
rect 13219 39292 13228 39332
rect 13268 39292 13516 39332
rect 13556 39292 13565 39332
rect 18799 39292 18808 39332
rect 18848 39292 18890 39332
rect 18930 39292 18972 39332
rect 19012 39292 19054 39332
rect 19094 39292 19136 39332
rect 19176 39292 19185 39332
rect 12931 39291 12989 39292
rect 8899 39248 8957 39249
rect 2500 39208 6988 39248
rect 7028 39208 7037 39248
rect 8899 39208 8908 39248
rect 8948 39208 10636 39248
rect 10676 39208 11500 39248
rect 11540 39208 11549 39248
rect 13411 39208 13420 39248
rect 13460 39208 17164 39248
rect 17204 39208 17213 39248
rect 18019 39208 18028 39248
rect 18068 39208 18077 39248
rect 0 39080 80 39100
rect 2500 39080 2540 39208
rect 8899 39207 8957 39208
rect 11779 39164 11837 39165
rect 4003 39124 4012 39164
rect 4052 39124 4972 39164
rect 5012 39124 5021 39164
rect 6220 39124 6796 39164
rect 6836 39124 6845 39164
rect 11011 39124 11020 39164
rect 11060 39124 11788 39164
rect 11828 39124 11837 39164
rect 0 39040 2540 39080
rect 0 39020 80 39040
rect 1411 38996 1469 38997
rect 6220 38996 6260 39124
rect 11779 39123 11837 39124
rect 13507 39164 13565 39165
rect 18028 39164 18068 39208
rect 13507 39124 13516 39164
rect 13556 39124 18068 39164
rect 18115 39124 18124 39164
rect 18164 39124 19180 39164
rect 19220 39124 19229 39164
rect 13507 39123 13565 39124
rect 21424 39080 21504 39100
rect 6403 39040 6412 39080
rect 6452 39040 8140 39080
rect 8180 39040 8332 39080
rect 8372 39040 8381 39080
rect 10819 39040 10828 39080
rect 10868 39040 12940 39080
rect 12980 39040 12989 39080
rect 15523 39040 15532 39080
rect 15572 39040 15916 39080
rect 15956 39040 15965 39080
rect 16963 39040 16972 39080
rect 17012 39040 21504 39080
rect 21424 39020 21504 39040
rect 17635 38996 17693 38997
rect 1315 38956 1324 38996
rect 1364 38956 1420 38996
rect 1460 38956 1469 38996
rect 1411 38955 1469 38956
rect 1516 38956 6260 38996
rect 8899 38956 8908 38996
rect 8948 38956 12652 38996
rect 12692 38956 12701 38996
rect 16195 38956 16204 38996
rect 16244 38956 17644 38996
rect 17684 38956 17693 38996
rect 1516 38912 1556 38956
rect 17635 38955 17693 38956
rect 1699 38912 1757 38913
rect 14179 38912 14237 38913
rect 16675 38912 16733 38913
rect 1507 38872 1516 38912
rect 1556 38872 1565 38912
rect 1614 38872 1708 38912
rect 1748 38872 1757 38912
rect 5923 38872 5932 38912
rect 5972 38872 7756 38912
rect 7796 38872 7948 38912
rect 7988 38872 7997 38912
rect 8419 38872 8428 38912
rect 8468 38872 9100 38912
rect 9140 38872 9149 38912
rect 12259 38872 12268 38912
rect 12308 38872 12317 38912
rect 12547 38872 12556 38912
rect 12596 38872 13612 38912
rect 13652 38872 13661 38912
rect 14179 38872 14188 38912
rect 14228 38872 16684 38912
rect 16724 38872 20044 38912
rect 20084 38872 20093 38912
rect 1699 38871 1757 38872
rect 8428 38828 8468 38872
rect 11203 38828 11261 38829
rect 6403 38788 6412 38828
rect 6452 38788 8468 38828
rect 10051 38788 10060 38828
rect 10100 38788 11212 38828
rect 11252 38788 11261 38828
rect 12268 38828 12308 38872
rect 14179 38871 14237 38872
rect 16675 38871 16733 38872
rect 12268 38788 16012 38828
rect 16052 38788 16396 38828
rect 16436 38788 16445 38828
rect 18691 38788 18700 38828
rect 18740 38788 19276 38828
rect 19316 38788 19325 38828
rect 11203 38787 11261 38788
rect 18211 38744 18269 38745
rect 18979 38744 19037 38745
rect 21424 38744 21504 38764
rect 1795 38704 1804 38744
rect 1844 38704 5260 38744
rect 5300 38704 5309 38744
rect 7075 38704 7084 38744
rect 7124 38704 9388 38744
rect 9428 38704 9437 38744
rect 12259 38704 12268 38744
rect 12308 38704 12317 38744
rect 15619 38704 15628 38744
rect 15668 38704 16876 38744
rect 16916 38704 16925 38744
rect 17059 38704 17068 38744
rect 17108 38704 17740 38744
rect 17780 38704 17789 38744
rect 18126 38704 18220 38744
rect 18260 38704 18269 38744
rect 18894 38704 18988 38744
rect 19028 38704 19372 38744
rect 19412 38704 19421 38744
rect 19939 38704 19948 38744
rect 19988 38704 21504 38744
rect 2083 38660 2141 38661
rect 12268 38660 12308 38704
rect 18211 38703 18269 38704
rect 18979 38703 19037 38704
rect 21424 38684 21504 38704
rect 1987 38620 1996 38660
rect 2036 38620 2092 38660
rect 2132 38620 2141 38660
rect 2467 38620 2476 38660
rect 2516 38620 5356 38660
rect 5396 38620 5405 38660
rect 5827 38620 5836 38660
rect 5876 38620 11404 38660
rect 11444 38620 11453 38660
rect 12268 38620 21004 38660
rect 21044 38620 21053 38660
rect 2083 38619 2141 38620
rect 0 38576 80 38596
rect 8611 38576 8669 38577
rect 0 38536 4148 38576
rect 4919 38536 4928 38576
rect 4968 38536 5010 38576
rect 5050 38536 5092 38576
rect 5132 38536 5174 38576
rect 5214 38536 5256 38576
rect 5296 38536 5305 38576
rect 7843 38536 7852 38576
rect 7892 38536 8620 38576
rect 8660 38536 18988 38576
rect 19028 38536 19037 38576
rect 20039 38536 20048 38576
rect 20088 38536 20130 38576
rect 20170 38536 20212 38576
rect 20252 38536 20294 38576
rect 20334 38536 20376 38576
rect 20416 38536 20425 38576
rect 0 38516 80 38536
rect 1027 38452 1036 38492
rect 1076 38452 3340 38492
rect 3380 38452 3389 38492
rect 1411 38368 1420 38408
rect 1460 38368 3052 38408
rect 3092 38368 3101 38408
rect 2083 38284 2092 38324
rect 2132 38284 2516 38324
rect 2947 38284 2956 38324
rect 2996 38284 3340 38324
rect 3380 38284 3389 38324
rect 835 38116 844 38156
rect 884 38116 1228 38156
rect 1268 38116 1277 38156
rect 0 38072 80 38092
rect 1795 38072 1853 38073
rect 2476 38072 2516 38284
rect 4108 38240 4148 38536
rect 8611 38535 8669 38536
rect 4195 38452 4204 38492
rect 4244 38452 8332 38492
rect 8372 38452 8381 38492
rect 12259 38452 12268 38492
rect 12308 38452 12460 38492
rect 12500 38452 12509 38492
rect 12643 38452 12652 38492
rect 12692 38452 20180 38492
rect 12643 38408 12701 38409
rect 12835 38408 12893 38409
rect 20140 38408 20180 38452
rect 21424 38408 21504 38428
rect 6595 38368 6604 38408
rect 6644 38368 6892 38408
rect 6932 38368 6941 38408
rect 8611 38368 8620 38408
rect 8660 38368 12652 38408
rect 12692 38368 12701 38408
rect 12750 38368 12844 38408
rect 12884 38368 12893 38408
rect 13027 38368 13036 38408
rect 13076 38368 13085 38408
rect 15427 38368 15436 38408
rect 15476 38368 15820 38408
rect 15860 38368 15869 38408
rect 15916 38368 18796 38408
rect 18836 38368 18845 38408
rect 19459 38368 19468 38408
rect 19508 38368 19517 38408
rect 20140 38368 21504 38408
rect 12643 38367 12701 38368
rect 12835 38367 12893 38368
rect 13036 38324 13076 38368
rect 15916 38324 15956 38368
rect 6307 38284 6316 38324
rect 6356 38284 6396 38324
rect 9283 38284 9292 38324
rect 9332 38284 12940 38324
rect 12980 38284 12989 38324
rect 13036 38284 15956 38324
rect 18403 38284 18412 38324
rect 18452 38284 19372 38324
rect 19412 38284 19421 38324
rect 6316 38240 6356 38284
rect 9571 38240 9629 38241
rect 10339 38240 10397 38241
rect 12643 38240 12701 38241
rect 14179 38240 14237 38241
rect 19468 38240 19508 38368
rect 21424 38348 21504 38368
rect 20131 38324 20189 38325
rect 20131 38284 20140 38324
rect 20180 38284 20274 38324
rect 20131 38283 20189 38284
rect 4108 38200 7276 38240
rect 7316 38200 7325 38240
rect 9486 38200 9580 38240
rect 9620 38200 10060 38240
rect 10100 38200 10109 38240
rect 10339 38200 10348 38240
rect 10388 38200 10540 38240
rect 10580 38200 10589 38240
rect 10723 38200 10732 38240
rect 10772 38200 12076 38240
rect 12116 38200 12125 38240
rect 12259 38200 12268 38240
rect 12308 38200 12460 38240
rect 12500 38200 12509 38240
rect 12643 38200 12652 38240
rect 12692 38200 13612 38240
rect 13652 38200 14188 38240
rect 14228 38200 14237 38240
rect 14947 38200 14956 38240
rect 14996 38200 15436 38240
rect 15476 38200 15485 38240
rect 17443 38200 17452 38240
rect 17492 38200 17836 38240
rect 17876 38200 17885 38240
rect 19468 38200 21428 38240
rect 9571 38199 9629 38200
rect 10339 38199 10397 38200
rect 12643 38199 12701 38200
rect 14179 38199 14237 38200
rect 7363 38156 7421 38157
rect 7075 38116 7084 38156
rect 7124 38116 7372 38156
rect 7412 38116 7421 38156
rect 7363 38115 7421 38116
rect 8419 38156 8477 38157
rect 8419 38116 8428 38156
rect 8468 38116 10444 38156
rect 10484 38116 10493 38156
rect 10540 38116 10868 38156
rect 11395 38116 11404 38156
rect 11444 38116 19660 38156
rect 19700 38116 19709 38156
rect 8419 38115 8477 38116
rect 10540 38072 10580 38116
rect 0 38032 1804 38072
rect 1844 38032 1853 38072
rect 2467 38032 2476 38072
rect 2516 38032 2525 38072
rect 3043 38032 3052 38072
rect 3092 38032 8812 38072
rect 8852 38032 8861 38072
rect 9379 38032 9388 38072
rect 9428 38032 10580 38072
rect 0 38012 80 38032
rect 1795 38031 1853 38032
rect 4195 37988 4253 37989
rect 10828 37988 10868 38116
rect 21388 38092 21428 38200
rect 12067 38032 12076 38072
rect 12116 38032 13804 38072
rect 13844 38032 13853 38072
rect 15043 38032 15052 38072
rect 15092 38032 15340 38072
rect 15380 38032 15389 38072
rect 17068 38032 17356 38072
rect 17396 38032 17405 38072
rect 21388 38032 21504 38092
rect 17068 37988 17108 38032
rect 21424 38012 21504 38032
rect 2179 37948 2188 37988
rect 2228 37948 4204 37988
rect 4244 37948 4253 37988
rect 4195 37947 4253 37948
rect 4300 37948 10732 37988
rect 10772 37948 10781 37988
rect 10828 37948 17108 37988
rect 17251 37948 17260 37988
rect 17300 37948 17740 37988
rect 17780 37948 17789 37988
rect 19075 37948 19084 37988
rect 19124 37948 19372 37988
rect 19412 37948 19421 37988
rect 19939 37948 19948 37988
rect 19988 37948 20908 37988
rect 20948 37948 20957 37988
rect 2563 37904 2621 37905
rect 4300 37904 4340 37948
rect 11203 37904 11261 37905
rect 17347 37904 17405 37905
rect 1603 37864 1612 37904
rect 1652 37864 2572 37904
rect 2612 37864 2621 37904
rect 2563 37863 2621 37864
rect 2668 37864 4340 37904
rect 8140 37864 11212 37904
rect 11252 37864 11261 37904
rect 11779 37864 11788 37904
rect 11828 37864 12556 37904
rect 12596 37864 12605 37904
rect 14275 37864 14284 37904
rect 14324 37864 15092 37904
rect 15139 37864 15148 37904
rect 15188 37864 15628 37904
rect 15668 37864 15677 37904
rect 17262 37864 17356 37904
rect 17396 37864 17405 37904
rect 19651 37864 19660 37904
rect 19700 37864 20620 37904
rect 20660 37864 20669 37904
rect 1795 37820 1853 37821
rect 2668 37820 2708 37864
rect 1795 37780 1804 37820
rect 1844 37780 2708 37820
rect 3108 37780 3148 37820
rect 3188 37780 3197 37820
rect 3679 37780 3688 37820
rect 3728 37780 3770 37820
rect 3810 37780 3852 37820
rect 3892 37780 3934 37820
rect 3974 37780 4016 37820
rect 4056 37780 4065 37820
rect 5316 37780 5356 37820
rect 5396 37780 5405 37820
rect 1795 37779 1853 37780
rect 2467 37736 2525 37737
rect 1507 37696 1516 37736
rect 1556 37696 2476 37736
rect 2516 37696 2525 37736
rect 3148 37736 3188 37780
rect 5356 37736 5396 37780
rect 8140 37736 8180 37864
rect 11203 37863 11261 37864
rect 15052 37820 15092 37864
rect 17347 37863 17405 37864
rect 8515 37780 8524 37820
rect 8564 37780 8660 37820
rect 15043 37780 15052 37820
rect 15092 37780 15101 37820
rect 15204 37780 15244 37820
rect 15284 37780 15293 37820
rect 18799 37780 18808 37820
rect 18848 37780 18890 37820
rect 18930 37780 18972 37820
rect 19012 37780 19054 37820
rect 19094 37780 19136 37820
rect 19176 37780 19185 37820
rect 3148 37696 3956 37736
rect 4483 37696 4492 37736
rect 4532 37696 4876 37736
rect 4916 37696 4925 37736
rect 5356 37696 8180 37736
rect 8323 37736 8381 37737
rect 8620 37736 8660 37780
rect 15244 37736 15284 37780
rect 15715 37736 15773 37737
rect 21424 37736 21504 37756
rect 8323 37696 8332 37736
rect 8372 37696 10732 37736
rect 10772 37696 11980 37736
rect 12020 37696 12029 37736
rect 13699 37696 13708 37736
rect 13748 37696 15148 37736
rect 15188 37696 15197 37736
rect 15244 37696 15724 37736
rect 15764 37696 15773 37736
rect 16867 37696 16876 37736
rect 16916 37696 17068 37736
rect 17108 37696 17117 37736
rect 20515 37696 20524 37736
rect 20564 37696 21504 37736
rect 2467 37695 2525 37696
rect 3916 37652 3956 37696
rect 8323 37695 8381 37696
rect 15715 37695 15773 37696
rect 21424 37676 21504 37696
rect 1795 37612 1804 37652
rect 1844 37612 2284 37652
rect 2324 37612 2333 37652
rect 2380 37612 2668 37652
rect 2708 37612 2717 37652
rect 3907 37612 3916 37652
rect 3956 37612 3965 37652
rect 4675 37612 4684 37652
rect 4724 37612 6124 37652
rect 6164 37612 6173 37652
rect 8035 37612 8044 37652
rect 8084 37612 8332 37652
rect 8372 37612 8381 37652
rect 13123 37612 13132 37652
rect 13172 37612 14708 37652
rect 15427 37612 15436 37652
rect 15476 37612 16300 37652
rect 16340 37612 16349 37652
rect 16396 37612 18508 37652
rect 18548 37612 18557 37652
rect 0 37568 80 37588
rect 2380 37568 2420 37612
rect 0 37528 212 37568
rect 1411 37528 1420 37568
rect 1460 37528 2420 37568
rect 2467 37568 2525 37569
rect 14668 37568 14708 37612
rect 16396 37568 16436 37612
rect 2467 37528 2476 37568
rect 2516 37528 4876 37568
rect 4916 37528 11116 37568
rect 11156 37528 11165 37568
rect 12739 37528 12748 37568
rect 12788 37528 13900 37568
rect 13940 37528 14572 37568
rect 14612 37528 14621 37568
rect 14668 37528 16436 37568
rect 17443 37528 17452 37568
rect 17492 37528 21332 37568
rect 0 37508 80 37528
rect 172 37400 212 37528
rect 2467 37527 2525 37528
rect 2755 37484 2813 37485
rect 1603 37444 1612 37484
rect 1652 37444 2764 37484
rect 2804 37444 2813 37484
rect 5251 37444 5260 37484
rect 5300 37444 5309 37484
rect 6499 37444 6508 37484
rect 6548 37444 13420 37484
rect 13460 37444 16300 37484
rect 16340 37444 16349 37484
rect 17155 37444 17164 37484
rect 17204 37444 18220 37484
rect 18260 37444 18269 37484
rect 18883 37444 18892 37484
rect 18932 37444 20044 37484
rect 20084 37444 20093 37484
rect 2755 37443 2813 37444
rect 20 37360 212 37400
rect 643 37400 701 37401
rect 2371 37400 2429 37401
rect 643 37360 652 37400
rect 692 37360 2380 37400
rect 2420 37360 2429 37400
rect 20 37232 60 37360
rect 643 37359 701 37360
rect 2371 37359 2429 37360
rect 2563 37400 2621 37401
rect 4195 37400 4253 37401
rect 2563 37360 2572 37400
rect 2612 37360 2706 37400
rect 4110 37360 4204 37400
rect 4244 37360 4253 37400
rect 5260 37400 5300 37444
rect 7555 37400 7613 37401
rect 18115 37400 18173 37401
rect 21292 37400 21332 37528
rect 21424 37400 21504 37420
rect 5260 37360 7564 37400
rect 7604 37360 7613 37400
rect 7939 37360 7948 37400
rect 7988 37360 8140 37400
rect 8180 37360 8189 37400
rect 9763 37360 9772 37400
rect 9812 37360 10060 37400
rect 10100 37360 10109 37400
rect 13315 37360 13324 37400
rect 13364 37360 17260 37400
rect 17300 37360 17309 37400
rect 17827 37360 17836 37400
rect 17876 37360 18124 37400
rect 18164 37360 18173 37400
rect 18499 37360 18508 37400
rect 18548 37360 18796 37400
rect 18836 37360 18845 37400
rect 19843 37360 19852 37400
rect 19892 37360 20716 37400
rect 20756 37360 20765 37400
rect 21292 37360 21504 37400
rect 2563 37359 2621 37360
rect 4195 37359 4253 37360
rect 7555 37359 7613 37360
rect 18115 37359 18173 37360
rect 21424 37340 21504 37360
rect 1219 37316 1277 37317
rect 8323 37316 8381 37317
rect 19651 37316 19709 37317
rect 1219 37276 1228 37316
rect 1268 37276 2540 37316
rect 2659 37276 2668 37316
rect 2708 37276 2956 37316
rect 2996 37276 3005 37316
rect 7075 37276 7084 37316
rect 7124 37276 7660 37316
rect 7700 37276 7709 37316
rect 7843 37276 7852 37316
rect 7892 37276 8332 37316
rect 8372 37276 8381 37316
rect 8611 37276 8620 37316
rect 8660 37276 11360 37316
rect 12547 37276 12556 37316
rect 12596 37276 14860 37316
rect 14900 37276 14909 37316
rect 19566 37276 19660 37316
rect 19700 37276 19709 37316
rect 1219 37275 1277 37276
rect 1987 37232 2045 37233
rect 20 37192 1844 37232
rect 1902 37192 1996 37232
rect 2036 37192 2045 37232
rect 2500 37232 2540 37276
rect 8323 37275 8381 37276
rect 6883 37232 6941 37233
rect 11320 37232 11360 37276
rect 19651 37275 19709 37276
rect 2500 37192 4492 37232
rect 4532 37192 4541 37232
rect 6883 37192 6892 37232
rect 6932 37192 7276 37232
rect 7316 37192 7325 37232
rect 11320 37192 15244 37232
rect 15284 37192 15293 37232
rect 1804 37148 1844 37192
rect 1987 37191 2045 37192
rect 6883 37191 6941 37192
rect 9187 37148 9245 37149
rect 1804 37108 2036 37148
rect 0 37064 80 37084
rect 163 37064 221 37065
rect 1996 37064 2036 37108
rect 2500 37108 9196 37148
rect 9236 37108 9245 37148
rect 2500 37064 2540 37108
rect 9187 37107 9245 37108
rect 9379 37148 9437 37149
rect 16291 37148 16349 37149
rect 9379 37108 9388 37148
rect 9428 37108 13708 37148
rect 13748 37108 13757 37148
rect 13891 37108 13900 37148
rect 13940 37108 14188 37148
rect 14228 37108 14237 37148
rect 16291 37108 16300 37148
rect 16340 37108 16876 37148
rect 16916 37108 16925 37148
rect 18115 37108 18124 37148
rect 18164 37108 19564 37148
rect 19604 37108 19613 37148
rect 9379 37107 9437 37108
rect 16291 37107 16349 37108
rect 21424 37064 21504 37084
rect 0 37024 172 37064
rect 212 37024 221 37064
rect 1603 37024 1612 37064
rect 1652 37024 1900 37064
rect 1940 37024 1949 37064
rect 1996 37024 2284 37064
rect 2324 37024 2540 37064
rect 4919 37024 4928 37064
rect 4968 37024 5010 37064
rect 5050 37024 5092 37064
rect 5132 37024 5174 37064
rect 5214 37024 5256 37064
rect 5296 37024 5305 37064
rect 6787 37024 6796 37064
rect 6836 37024 8908 37064
rect 8948 37024 10060 37064
rect 10100 37024 10109 37064
rect 10819 37024 10828 37064
rect 10868 37024 10877 37064
rect 11320 37024 15628 37064
rect 15668 37024 18700 37064
rect 18740 37024 18749 37064
rect 20039 37024 20048 37064
rect 20088 37024 20130 37064
rect 20170 37024 20212 37064
rect 20252 37024 20294 37064
rect 20334 37024 20376 37064
rect 20416 37024 20425 37064
rect 20812 37024 21504 37064
rect 0 37004 80 37024
rect 163 37023 221 37024
rect 10828 36980 10868 37024
rect 1507 36940 1516 36980
rect 1556 36940 2380 36980
rect 2420 36940 2429 36980
rect 2476 36940 11020 36980
rect 11060 36940 11069 36980
rect 2476 36897 2516 36940
rect 2467 36896 2525 36897
rect 1891 36856 1900 36896
rect 1940 36856 2420 36896
rect 2275 36812 2333 36813
rect 1315 36772 1324 36812
rect 1364 36772 2284 36812
rect 2324 36772 2333 36812
rect 2380 36812 2420 36856
rect 2467 36856 2476 36896
rect 2516 36856 2525 36896
rect 2467 36855 2525 36856
rect 3523 36896 3581 36897
rect 4972 36896 5012 36940
rect 11320 36896 11360 37024
rect 20812 36980 20852 37024
rect 21424 37004 21504 37024
rect 11587 36940 11596 36980
rect 11636 36940 20852 36980
rect 14659 36896 14717 36897
rect 3523 36856 3532 36896
rect 3572 36856 3820 36896
rect 3860 36856 3869 36896
rect 4963 36856 4972 36896
rect 5012 36856 5021 36896
rect 7363 36856 7372 36896
rect 7412 36856 8620 36896
rect 8660 36856 8669 36896
rect 10147 36856 10156 36896
rect 10196 36856 11360 36896
rect 12835 36856 12844 36896
rect 12884 36856 13324 36896
rect 13364 36856 13373 36896
rect 14574 36856 14668 36896
rect 14708 36856 14717 36896
rect 14947 36856 14956 36896
rect 14996 36856 15340 36896
rect 15380 36856 15389 36896
rect 17059 36856 17068 36896
rect 17108 36856 17836 36896
rect 17876 36856 18316 36896
rect 18356 36856 18365 36896
rect 19171 36856 19180 36896
rect 19220 36856 19229 36896
rect 19555 36856 19564 36896
rect 19604 36856 21292 36896
rect 21332 36856 21341 36896
rect 3523 36855 3581 36856
rect 14659 36855 14717 36856
rect 19180 36812 19220 36856
rect 20995 36812 21053 36813
rect 2380 36772 2764 36812
rect 2804 36772 2813 36812
rect 4195 36772 4204 36812
rect 4244 36772 7276 36812
rect 7316 36772 7325 36812
rect 8227 36772 8236 36812
rect 8276 36772 8524 36812
rect 8564 36772 8573 36812
rect 10435 36772 10444 36812
rect 10484 36772 11308 36812
rect 11348 36772 11357 36812
rect 12163 36772 12172 36812
rect 12212 36772 12460 36812
rect 12500 36772 12509 36812
rect 14179 36772 14188 36812
rect 14228 36772 18028 36812
rect 18068 36772 18077 36812
rect 19180 36772 21004 36812
rect 21044 36772 21053 36812
rect 2275 36771 2333 36772
rect 20995 36771 21053 36772
rect 5827 36728 5885 36729
rect 12643 36728 12701 36729
rect 21424 36728 21504 36748
rect 2371 36688 2380 36728
rect 2420 36688 5836 36728
rect 5876 36688 5885 36728
rect 6979 36688 6988 36728
rect 7028 36688 8812 36728
rect 8852 36688 8861 36728
rect 9763 36688 9772 36728
rect 9812 36688 10348 36728
rect 10388 36688 10397 36728
rect 11683 36688 11692 36728
rect 11732 36688 12268 36728
rect 12308 36688 12317 36728
rect 12643 36688 12652 36728
rect 12692 36688 19412 36728
rect 19459 36688 19468 36728
rect 19508 36688 21504 36728
rect 5827 36687 5885 36688
rect 12643 36687 12701 36688
rect 11971 36644 12029 36645
rect 19372 36644 19412 36688
rect 21424 36668 21504 36688
rect 1315 36604 1324 36644
rect 1364 36604 11980 36644
rect 12020 36604 12029 36644
rect 15523 36604 15532 36644
rect 15572 36604 15916 36644
rect 15956 36604 15965 36644
rect 16579 36604 16588 36644
rect 16628 36604 17356 36644
rect 17396 36604 17405 36644
rect 19363 36604 19372 36644
rect 19412 36604 19421 36644
rect 11971 36603 12029 36604
rect 0 36560 80 36580
rect 6691 36560 6749 36561
rect 18499 36560 18557 36561
rect 21187 36560 21245 36561
rect 0 36520 6508 36560
rect 6548 36520 6557 36560
rect 6606 36520 6700 36560
rect 6740 36520 6892 36560
rect 6932 36520 6941 36560
rect 7267 36520 7276 36560
rect 7316 36520 8716 36560
rect 8756 36520 9772 36560
rect 9812 36520 9821 36560
rect 9955 36520 9964 36560
rect 10004 36520 10732 36560
rect 10772 36520 10781 36560
rect 14947 36520 14956 36560
rect 14996 36520 15436 36560
rect 15476 36520 15485 36560
rect 16003 36520 16012 36560
rect 16052 36520 18508 36560
rect 18548 36520 18557 36560
rect 19939 36520 19948 36560
rect 19988 36520 21196 36560
rect 21236 36520 21245 36560
rect 0 36500 80 36520
rect 6691 36519 6749 36520
rect 18499 36519 18557 36520
rect 21187 36519 21245 36520
rect 931 36476 989 36477
rect 931 36436 940 36476
rect 980 36436 1708 36476
rect 1748 36436 1757 36476
rect 8899 36436 8908 36476
rect 8948 36436 9484 36476
rect 9524 36436 9533 36476
rect 10531 36436 10540 36476
rect 10580 36436 11020 36476
rect 11060 36436 11069 36476
rect 18307 36436 18316 36476
rect 18356 36436 18892 36476
rect 18932 36436 18941 36476
rect 931 36435 989 36436
rect 21424 36392 21504 36412
rect 10051 36352 10060 36392
rect 10100 36352 11980 36392
rect 12020 36352 12268 36392
rect 12308 36352 12748 36392
rect 12788 36352 12797 36392
rect 15427 36352 15436 36392
rect 15476 36352 18412 36392
rect 18452 36352 18700 36392
rect 18740 36352 18749 36392
rect 20899 36352 20908 36392
rect 20948 36352 21504 36392
rect 21424 36332 21504 36352
rect 3679 36268 3688 36308
rect 3728 36268 3770 36308
rect 3810 36268 3852 36308
rect 3892 36268 3934 36308
rect 3974 36268 4016 36308
rect 4056 36268 4065 36308
rect 16675 36268 16684 36308
rect 16724 36268 17452 36308
rect 17492 36268 17501 36308
rect 18799 36268 18808 36308
rect 18848 36268 18890 36308
rect 18930 36268 18972 36308
rect 19012 36268 19054 36308
rect 19094 36268 19136 36308
rect 19176 36268 19185 36308
rect 2500 36184 11788 36224
rect 11828 36184 11837 36224
rect 0 36056 80 36076
rect 2500 36056 2540 36184
rect 4099 36140 4157 36141
rect 4003 36100 4012 36140
rect 4052 36100 4108 36140
rect 4148 36100 4157 36140
rect 16675 36100 16684 36140
rect 16724 36100 16876 36140
rect 16916 36100 16925 36140
rect 4099 36099 4157 36100
rect 0 36016 1708 36056
rect 1748 36016 2540 36056
rect 3523 36056 3581 36057
rect 21424 36056 21504 36076
rect 3523 36016 3532 36056
rect 3572 36016 3820 36056
rect 3860 36016 4300 36056
rect 4340 36016 4349 36056
rect 7555 36016 7564 36056
rect 7604 36016 8716 36056
rect 8756 36016 8765 36056
rect 20611 36016 20620 36056
rect 20660 36016 21504 36056
rect 0 35996 80 36016
rect 3523 36015 3581 36016
rect 21424 35996 21504 36016
rect 8803 35972 8861 35973
rect 16291 35972 16349 35973
rect 19939 35972 19997 35973
rect 1315 35932 1324 35972
rect 1364 35932 2764 35972
rect 2804 35932 2813 35972
rect 3619 35932 3628 35972
rect 3668 35932 8812 35972
rect 8852 35932 8861 35972
rect 14563 35932 14572 35972
rect 14612 35932 15244 35972
rect 15284 35932 16300 35972
rect 16340 35932 16876 35972
rect 16916 35932 16925 35972
rect 17635 35932 17644 35972
rect 17684 35932 17932 35972
rect 17972 35932 19564 35972
rect 19604 35932 19613 35972
rect 19854 35932 19948 35972
rect 19988 35932 19997 35972
rect 8803 35931 8861 35932
rect 16291 35931 16349 35932
rect 19939 35931 19997 35932
rect 6595 35888 6653 35889
rect 9667 35888 9725 35889
rect 3331 35848 3340 35888
rect 3380 35848 4972 35888
rect 5012 35848 5021 35888
rect 6510 35848 6604 35888
rect 6644 35848 7948 35888
rect 7988 35848 7997 35888
rect 9667 35848 9676 35888
rect 9716 35848 9964 35888
rect 10004 35848 10013 35888
rect 11320 35848 19276 35888
rect 19316 35848 19325 35888
rect 20515 35848 20524 35888
rect 20564 35848 21388 35888
rect 21428 35848 21437 35888
rect 4972 35804 5012 35848
rect 6595 35847 6653 35848
rect 9667 35847 9725 35848
rect 11320 35804 11360 35848
rect 18211 35804 18269 35805
rect 4972 35764 7276 35804
rect 7316 35764 7325 35804
rect 8227 35764 8236 35804
rect 8276 35764 11360 35804
rect 16483 35764 16492 35804
rect 16532 35764 17068 35804
rect 17108 35764 17117 35804
rect 18211 35764 18220 35804
rect 18260 35764 18316 35804
rect 18356 35764 18365 35804
rect 18211 35763 18269 35764
rect 2179 35720 2237 35721
rect 4483 35720 4541 35721
rect 8995 35720 9053 35721
rect 21424 35720 21504 35740
rect 2094 35680 2188 35720
rect 2228 35680 2237 35720
rect 4398 35680 4492 35720
rect 4532 35680 4541 35720
rect 4771 35680 4780 35720
rect 4820 35680 5452 35720
rect 5492 35680 5501 35720
rect 7651 35680 7660 35720
rect 7700 35680 8044 35720
rect 8084 35680 8093 35720
rect 8995 35680 9004 35720
rect 9044 35680 9868 35720
rect 9908 35680 10060 35720
rect 10100 35680 10109 35720
rect 19075 35680 19084 35720
rect 19124 35680 19756 35720
rect 19796 35680 19805 35720
rect 21379 35680 21388 35720
rect 21428 35680 21504 35720
rect 2179 35679 2237 35680
rect 4483 35679 4541 35680
rect 8995 35679 9053 35680
rect 21424 35660 21504 35680
rect 4684 35596 7852 35636
rect 7892 35596 7901 35636
rect 0 35552 80 35572
rect 4684 35552 4724 35596
rect 16483 35552 16541 35553
rect 0 35512 4684 35552
rect 4724 35512 4733 35552
rect 4919 35512 4928 35552
rect 4968 35512 5010 35552
rect 5050 35512 5092 35552
rect 5132 35512 5174 35552
rect 5214 35512 5256 35552
rect 5296 35512 5305 35552
rect 7555 35512 7564 35552
rect 7604 35512 8236 35552
rect 8276 35512 8285 35552
rect 9091 35512 9100 35552
rect 9140 35512 16492 35552
rect 16532 35512 18124 35552
rect 18164 35512 18173 35552
rect 20039 35512 20048 35552
rect 20088 35512 20130 35552
rect 20170 35512 20212 35552
rect 20252 35512 20294 35552
rect 20334 35512 20376 35552
rect 20416 35512 20425 35552
rect 0 35492 80 35512
rect 16483 35511 16541 35512
rect 7459 35468 7517 35469
rect 9571 35468 9629 35469
rect 14755 35468 14813 35469
rect 20611 35468 20669 35469
rect 7374 35428 7468 35468
rect 7508 35428 7517 35468
rect 9486 35428 9580 35468
rect 9620 35428 9629 35468
rect 11491 35428 11500 35468
rect 11540 35428 14764 35468
rect 14804 35428 16820 35468
rect 16867 35428 16876 35468
rect 16916 35428 20620 35468
rect 20660 35428 20669 35468
rect 7459 35427 7517 35428
rect 9571 35427 9629 35428
rect 14755 35427 14813 35428
rect 16099 35384 16157 35385
rect 1891 35344 1900 35384
rect 1940 35344 4780 35384
rect 4820 35344 4829 35384
rect 4963 35344 4972 35384
rect 5012 35344 11308 35384
rect 11348 35344 11357 35384
rect 13891 35344 13900 35384
rect 13940 35344 14668 35384
rect 14708 35344 14717 35384
rect 15907 35344 15916 35384
rect 15956 35344 16108 35384
rect 16148 35344 16157 35384
rect 16780 35384 16820 35428
rect 20611 35427 20669 35428
rect 21424 35384 21504 35404
rect 16780 35344 18644 35384
rect 19939 35344 19948 35384
rect 19988 35344 21504 35384
rect 16099 35343 16157 35344
rect 8707 35300 8765 35301
rect 9283 35300 9341 35301
rect 2460 35260 2469 35300
rect 2509 35260 3052 35300
rect 3092 35260 3101 35300
rect 5635 35260 5644 35300
rect 5684 35260 6316 35300
rect 6356 35260 6365 35300
rect 8707 35260 8716 35300
rect 8756 35260 9004 35300
rect 9044 35260 9053 35300
rect 9198 35260 9292 35300
rect 9332 35260 9341 35300
rect 13027 35260 13036 35300
rect 13076 35260 13708 35300
rect 13748 35260 13757 35300
rect 14275 35260 14284 35300
rect 14324 35260 14333 35300
rect 14467 35260 14476 35300
rect 14516 35260 14525 35300
rect 14947 35260 14956 35300
rect 14996 35260 18124 35300
rect 18164 35260 18173 35300
rect 8707 35259 8765 35260
rect 9283 35259 9341 35260
rect 2563 35216 2621 35217
rect 1987 35176 1996 35216
rect 2036 35176 2572 35216
rect 2612 35176 2621 35216
rect 2563 35175 2621 35176
rect 2755 35216 2813 35217
rect 12643 35216 12701 35217
rect 14284 35216 14324 35260
rect 2755 35176 2764 35216
rect 2804 35176 4012 35216
rect 4052 35176 4061 35216
rect 6211 35176 6220 35216
rect 6260 35176 7372 35216
rect 7412 35176 10636 35216
rect 10676 35176 10685 35216
rect 12558 35176 12652 35216
rect 12692 35176 12701 35216
rect 13507 35176 13516 35216
rect 13556 35176 14324 35216
rect 2755 35175 2813 35176
rect 12643 35175 12701 35176
rect 739 35132 797 35133
rect 12835 35132 12893 35133
rect 14476 35132 14516 35260
rect 17635 35216 17693 35217
rect 18604 35216 18644 35344
rect 21424 35324 21504 35344
rect 19267 35260 19276 35300
rect 19316 35260 19852 35300
rect 19892 35260 19901 35300
rect 19939 35216 19997 35217
rect 15619 35176 15628 35216
rect 15668 35176 16108 35216
rect 16148 35176 16157 35216
rect 17550 35176 17644 35216
rect 17684 35176 17693 35216
rect 18595 35176 18604 35216
rect 18644 35176 18653 35216
rect 19854 35176 19948 35216
rect 19988 35176 19997 35216
rect 17635 35175 17693 35176
rect 19939 35175 19997 35176
rect 15907 35132 15965 35133
rect 739 35092 748 35132
rect 788 35092 1420 35132
rect 1460 35092 1469 35132
rect 2947 35092 2956 35132
rect 2996 35092 3532 35132
rect 3572 35092 3581 35132
rect 4483 35092 4492 35132
rect 4532 35092 8908 35132
rect 8948 35092 8957 35132
rect 9004 35092 12172 35132
rect 12212 35092 12221 35132
rect 12835 35092 12844 35132
rect 12884 35092 14516 35132
rect 15822 35092 15916 35132
rect 15956 35092 15965 35132
rect 739 35091 797 35092
rect 0 35048 80 35068
rect 8707 35048 8765 35049
rect 9004 35048 9044 35092
rect 12835 35091 12893 35092
rect 15907 35091 15965 35092
rect 16012 35092 19468 35132
rect 19508 35092 19517 35132
rect 16012 35048 16052 35092
rect 17059 35048 17117 35049
rect 21424 35048 21504 35068
rect 0 35008 1556 35048
rect 1603 35008 1612 35048
rect 1652 35008 2092 35048
rect 2132 35008 2141 35048
rect 4099 35008 4108 35048
rect 4148 35008 5972 35048
rect 7267 35008 7276 35048
rect 7316 35008 7468 35048
rect 7508 35008 8716 35048
rect 8756 35008 8765 35048
rect 8995 35008 9004 35048
rect 9044 35008 9053 35048
rect 12355 35008 12364 35048
rect 12404 35008 16052 35048
rect 16974 35008 17068 35048
rect 17108 35008 17117 35048
rect 17251 35008 17260 35048
rect 17300 35008 21504 35048
rect 0 34988 80 35008
rect 1516 34964 1556 35008
rect 5932 34964 5972 35008
rect 8707 35007 8765 35008
rect 17059 35007 17117 35008
rect 21424 34988 21504 35008
rect 1507 34924 1516 34964
rect 1556 34924 1565 34964
rect 3619 34924 3628 34964
rect 3668 34924 5548 34964
rect 5588 34924 5597 34964
rect 5932 34924 7756 34964
rect 7796 34924 7805 34964
rect 10819 34924 10828 34964
rect 10868 34924 11500 34964
rect 11540 34924 11549 34964
rect 12259 34924 12268 34964
rect 12308 34924 13900 34964
rect 13940 34924 13949 34964
rect 1123 34880 1181 34881
rect 13027 34880 13085 34881
rect 14659 34880 14717 34881
rect 16099 34880 16157 34881
rect 1123 34840 1132 34880
rect 1172 34840 5740 34880
rect 5780 34840 5789 34880
rect 6220 34840 11360 34880
rect 1123 34839 1181 34840
rect 6220 34796 6260 34840
rect 11320 34796 11360 34840
rect 13027 34840 13036 34880
rect 13076 34840 13324 34880
rect 13364 34840 13373 34880
rect 14371 34840 14380 34880
rect 14420 34840 14668 34880
rect 14708 34840 14717 34880
rect 16014 34840 16108 34880
rect 16148 34840 16157 34880
rect 13027 34839 13085 34840
rect 14659 34839 14717 34840
rect 16099 34839 16157 34840
rect 3679 34756 3688 34796
rect 3728 34756 3770 34796
rect 3810 34756 3852 34796
rect 3892 34756 3934 34796
rect 3974 34756 4016 34796
rect 4056 34756 4065 34796
rect 5644 34756 6124 34796
rect 6164 34756 6260 34796
rect 6403 34756 6412 34796
rect 6452 34756 7276 34796
rect 7316 34756 7325 34796
rect 7372 34756 10348 34796
rect 10388 34756 10397 34796
rect 11320 34756 15724 34796
rect 15764 34756 16684 34796
rect 16724 34756 16733 34796
rect 18799 34756 18808 34796
rect 18848 34756 18890 34796
rect 18930 34756 18972 34796
rect 19012 34756 19054 34796
rect 19094 34756 19136 34796
rect 19176 34756 19185 34796
rect 3139 34712 3197 34713
rect 5644 34712 5684 34756
rect 7372 34712 7412 34756
rect 9379 34712 9437 34713
rect 13795 34712 13853 34713
rect 21424 34712 21504 34732
rect 3139 34672 3148 34712
rect 3188 34672 5684 34712
rect 5731 34672 5740 34712
rect 5780 34672 7412 34712
rect 8899 34672 8908 34712
rect 8948 34672 9388 34712
rect 9428 34672 9437 34712
rect 13710 34672 13804 34712
rect 13844 34672 13853 34712
rect 14755 34672 14764 34712
rect 14804 34672 15052 34712
rect 15092 34672 15101 34712
rect 15523 34672 15532 34712
rect 15572 34672 15820 34712
rect 15860 34672 15869 34712
rect 17635 34672 17644 34712
rect 17684 34672 18028 34712
rect 18068 34672 18077 34712
rect 21283 34672 21292 34712
rect 21332 34672 21504 34712
rect 3139 34671 3197 34672
rect 9379 34671 9437 34672
rect 13795 34671 13853 34672
rect 21424 34652 21504 34672
rect 2659 34628 2717 34629
rect 2659 34588 2668 34628
rect 2708 34588 3340 34628
rect 3380 34588 3389 34628
rect 7747 34588 7756 34628
rect 7796 34588 19852 34628
rect 19892 34588 19901 34628
rect 2659 34587 2717 34588
rect 0 34544 80 34564
rect 2083 34544 2141 34545
rect 0 34504 2092 34544
rect 2132 34504 2141 34544
rect 3427 34504 3436 34544
rect 3476 34504 5836 34544
rect 5876 34504 5885 34544
rect 0 34484 80 34504
rect 2083 34503 2141 34504
rect 6595 34460 6653 34461
rect 3907 34420 3916 34460
rect 3956 34420 4492 34460
rect 4532 34420 4541 34460
rect 6595 34420 6604 34460
rect 6644 34420 8428 34460
rect 8468 34420 8477 34460
rect 6595 34419 6653 34420
rect 1123 34376 1181 34377
rect 8131 34376 8189 34377
rect 1123 34336 1132 34376
rect 1172 34336 1228 34376
rect 1268 34336 1277 34376
rect 3331 34336 3340 34376
rect 3380 34336 5740 34376
rect 5780 34336 5789 34376
rect 6019 34336 6028 34376
rect 6068 34336 6412 34376
rect 6452 34336 6461 34376
rect 8035 34336 8044 34376
rect 8084 34336 8140 34376
rect 8180 34336 8189 34376
rect 1123 34335 1181 34336
rect 6028 34292 6068 34336
rect 8131 34335 8189 34336
rect 2500 34252 4588 34292
rect 4628 34252 4637 34292
rect 5635 34252 5644 34292
rect 5684 34252 6068 34292
rect 2500 34124 2540 34252
rect 8908 34208 8948 34588
rect 11107 34504 11116 34544
rect 11156 34504 17356 34544
rect 17396 34504 19756 34544
rect 19796 34504 19805 34544
rect 12931 34420 12940 34460
rect 12980 34420 13612 34460
rect 13652 34420 13804 34460
rect 13844 34420 13853 34460
rect 14275 34420 14284 34460
rect 14324 34420 14860 34460
rect 14900 34420 14909 34460
rect 17731 34420 17740 34460
rect 17780 34420 18604 34460
rect 18644 34420 18653 34460
rect 16771 34376 16829 34377
rect 21424 34376 21504 34396
rect 12451 34336 12460 34376
rect 12500 34336 13324 34376
rect 13364 34336 13373 34376
rect 15715 34336 15724 34376
rect 15764 34336 16012 34376
rect 16052 34336 16061 34376
rect 16483 34336 16492 34376
rect 16532 34336 16780 34376
rect 16820 34336 18124 34376
rect 18164 34336 18700 34376
rect 18740 34336 18749 34376
rect 20611 34336 20620 34376
rect 20660 34336 21504 34376
rect 16771 34335 16829 34336
rect 21424 34316 21504 34336
rect 13795 34292 13853 34293
rect 13219 34252 13228 34292
rect 13268 34252 13804 34292
rect 13844 34252 16876 34292
rect 16916 34252 16925 34292
rect 13795 34251 13853 34252
rect 18499 34208 18557 34209
rect 19555 34208 19613 34209
rect 3523 34168 3532 34208
rect 3572 34168 7564 34208
rect 7604 34168 7613 34208
rect 8899 34168 8908 34208
rect 8948 34168 8957 34208
rect 9667 34168 9676 34208
rect 9716 34168 11020 34208
rect 11060 34168 11069 34208
rect 14947 34168 14956 34208
rect 14996 34168 15148 34208
rect 15188 34168 15197 34208
rect 16003 34168 16012 34208
rect 16052 34168 16684 34208
rect 16724 34168 16733 34208
rect 18499 34168 18508 34208
rect 18548 34168 18796 34208
rect 18836 34168 18845 34208
rect 19470 34168 19564 34208
rect 19604 34168 19613 34208
rect 20035 34168 20044 34208
rect 20084 34168 21332 34208
rect 18499 34167 18557 34168
rect 19555 34167 19613 34168
rect 1228 34084 2540 34124
rect 3427 34084 3436 34124
rect 3476 34084 5932 34124
rect 5972 34084 6892 34124
rect 6932 34084 6941 34124
rect 9475 34084 9484 34124
rect 9524 34084 10636 34124
rect 10676 34084 10685 34124
rect 13315 34084 13324 34124
rect 13364 34084 19372 34124
rect 19412 34084 19421 34124
rect 0 34040 80 34060
rect 1228 34040 1268 34084
rect 10435 34040 10493 34041
rect 15427 34040 15485 34041
rect 21292 34040 21332 34168
rect 21424 34040 21504 34060
rect 0 34000 1268 34040
rect 1324 34000 4396 34040
rect 4436 34000 4445 34040
rect 4919 34000 4928 34040
rect 4968 34000 5010 34040
rect 5050 34000 5092 34040
rect 5132 34000 5174 34040
rect 5214 34000 5256 34040
rect 5296 34000 5305 34040
rect 5539 34000 5548 34040
rect 5588 34000 5972 34040
rect 0 33980 80 34000
rect 1027 33956 1085 33957
rect 1324 33956 1364 34000
rect 2467 33956 2525 33957
rect 5932 33956 5972 34000
rect 10435 34000 10444 34040
rect 10484 34000 12748 34040
rect 12788 34000 12797 34040
rect 13507 34000 13516 34040
rect 13556 34000 14380 34040
rect 14420 34000 15244 34040
rect 15284 34000 15293 34040
rect 15427 34000 15436 34040
rect 15476 34000 15570 34040
rect 20039 34000 20048 34040
rect 20088 34000 20130 34040
rect 20170 34000 20212 34040
rect 20252 34000 20294 34040
rect 20334 34000 20376 34040
rect 20416 34000 20425 34040
rect 21292 34000 21504 34040
rect 10435 33999 10493 34000
rect 15427 33999 15485 34000
rect 21424 33980 21504 34000
rect 1027 33916 1036 33956
rect 1076 33916 1364 33956
rect 1603 33916 1612 33956
rect 1652 33916 1804 33956
rect 1844 33916 1853 33956
rect 2382 33916 2476 33956
rect 2516 33916 2525 33956
rect 3619 33916 3628 33956
rect 3668 33916 5644 33956
rect 5684 33916 5693 33956
rect 5923 33916 5932 33956
rect 5972 33916 5981 33956
rect 15043 33916 15052 33956
rect 15092 33916 16588 33956
rect 16628 33916 16637 33956
rect 1027 33915 1085 33916
rect 2467 33915 2525 33916
rect 1891 33832 1900 33872
rect 1940 33832 9580 33872
rect 9620 33832 9629 33872
rect 11320 33832 19852 33872
rect 19892 33832 19901 33872
rect 11320 33788 11360 33832
rect 5452 33748 11116 33788
rect 11156 33748 11360 33788
rect 11971 33748 11980 33788
rect 12020 33748 19372 33788
rect 19412 33748 19421 33788
rect 5452 33705 5492 33748
rect 5443 33704 5501 33705
rect 8227 33704 8285 33705
rect 10435 33704 10493 33705
rect 21424 33704 21504 33724
rect 4195 33664 4204 33704
rect 4244 33664 5452 33704
rect 5492 33664 5501 33704
rect 6019 33664 6028 33704
rect 6068 33664 6796 33704
rect 6836 33664 6845 33704
rect 8142 33664 8236 33704
rect 8276 33664 8620 33704
rect 8660 33664 8669 33704
rect 10350 33664 10444 33704
rect 10484 33664 10493 33704
rect 11011 33664 11020 33704
rect 11060 33664 11308 33704
rect 11348 33664 11357 33704
rect 12739 33664 12748 33704
rect 12788 33664 13420 33704
rect 13460 33664 13469 33704
rect 14179 33664 14188 33704
rect 14228 33664 14476 33704
rect 14516 33664 17068 33704
rect 17108 33664 17117 33704
rect 17539 33664 17548 33704
rect 17588 33664 18316 33704
rect 18356 33664 18365 33704
rect 19651 33664 19660 33704
rect 19700 33664 21504 33704
rect 5443 33663 5501 33664
rect 835 33620 893 33621
rect 4675 33620 4733 33621
rect 6028 33620 6068 33664
rect 8227 33663 8285 33664
rect 10435 33663 10493 33664
rect 835 33580 844 33620
rect 884 33580 1420 33620
rect 1460 33580 1469 33620
rect 4675 33580 4684 33620
rect 4724 33580 6068 33620
rect 7747 33580 7756 33620
rect 7796 33580 8332 33620
rect 8372 33580 8381 33620
rect 835 33579 893 33580
rect 4675 33579 4733 33580
rect 0 33536 80 33556
rect 2851 33536 2909 33537
rect 10444 33536 10484 33663
rect 21424 33644 21504 33664
rect 18595 33620 18653 33621
rect 11683 33580 11692 33620
rect 11732 33580 18220 33620
rect 18260 33580 18269 33620
rect 18595 33580 18604 33620
rect 18644 33580 18988 33620
rect 19028 33580 19037 33620
rect 18595 33579 18653 33580
rect 0 33496 2860 33536
rect 2900 33496 2909 33536
rect 3043 33496 3052 33536
rect 3092 33496 10484 33536
rect 13027 33496 13036 33536
rect 13076 33496 13420 33536
rect 13460 33496 13804 33536
rect 13844 33496 13853 33536
rect 15331 33496 15340 33536
rect 15380 33496 15532 33536
rect 15572 33496 16204 33536
rect 16244 33496 16253 33536
rect 17620 33496 18892 33536
rect 18932 33496 18941 33536
rect 19171 33496 19180 33536
rect 19220 33496 20812 33536
rect 20852 33496 20861 33536
rect 0 33476 80 33496
rect 2851 33495 2909 33496
rect 2467 33452 2525 33453
rect 2382 33412 2476 33452
rect 2516 33412 2525 33452
rect 2467 33411 2525 33412
rect 9283 33452 9341 33453
rect 9283 33412 9292 33452
rect 9332 33412 9341 33452
rect 10147 33412 10156 33452
rect 10196 33412 10444 33452
rect 10484 33412 10493 33452
rect 13507 33412 13516 33452
rect 13556 33412 16492 33452
rect 16532 33412 16541 33452
rect 9283 33411 9341 33412
rect 9292 33368 9332 33411
rect 12643 33368 12701 33369
rect 17620 33368 17660 33496
rect 18403 33452 18461 33453
rect 20803 33452 20861 33453
rect 18318 33412 18412 33452
rect 18452 33412 18461 33452
rect 18787 33412 18796 33452
rect 18836 33412 18845 33452
rect 19267 33412 19276 33452
rect 19316 33412 19700 33452
rect 19939 33412 19948 33452
rect 19988 33412 20812 33452
rect 20852 33412 20861 33452
rect 18403 33411 18461 33412
rect 4195 33328 4204 33368
rect 4244 33328 5452 33368
rect 5492 33328 6508 33368
rect 6548 33328 6557 33368
rect 9292 33328 10636 33368
rect 10676 33328 10685 33368
rect 11320 33328 12652 33368
rect 12692 33328 12701 33368
rect 15427 33328 15436 33368
rect 15476 33328 17660 33368
rect 18796 33368 18836 33412
rect 19660 33368 19700 33412
rect 20803 33411 20861 33412
rect 21424 33368 21504 33388
rect 18796 33328 19508 33368
rect 19660 33328 21504 33368
rect 6211 33284 6269 33285
rect 3679 33244 3688 33284
rect 3728 33244 3770 33284
rect 3810 33244 3852 33284
rect 3892 33244 3934 33284
rect 3974 33244 4016 33284
rect 4056 33244 4065 33284
rect 6126 33244 6220 33284
rect 6260 33244 6269 33284
rect 6211 33243 6269 33244
rect 7171 33284 7229 33285
rect 9283 33284 9341 33285
rect 7171 33244 7180 33284
rect 7220 33244 7276 33284
rect 7316 33244 7325 33284
rect 9283 33244 9292 33284
rect 9332 33244 10252 33284
rect 10292 33244 10301 33284
rect 7171 33243 7229 33244
rect 9283 33243 9341 33244
rect 1507 33200 1565 33201
rect 1891 33200 1949 33201
rect 5827 33200 5885 33201
rect 1422 33160 1516 33200
rect 1556 33160 1565 33200
rect 1806 33160 1900 33200
rect 1940 33160 1949 33200
rect 2371 33160 2380 33200
rect 2420 33160 5836 33200
rect 5876 33160 10060 33200
rect 10100 33160 10109 33200
rect 1507 33159 1565 33160
rect 1891 33159 1949 33160
rect 5827 33159 5885 33160
rect 11320 33116 11360 33328
rect 12643 33327 12701 33328
rect 19468 33284 19508 33328
rect 21424 33308 21504 33328
rect 15715 33244 15724 33284
rect 15764 33244 16300 33284
rect 16340 33244 16349 33284
rect 18799 33244 18808 33284
rect 18848 33244 18890 33284
rect 18930 33244 18972 33284
rect 19012 33244 19054 33284
rect 19094 33244 19136 33284
rect 19176 33244 19185 33284
rect 19468 33244 21196 33284
rect 21236 33244 21245 33284
rect 19843 33200 19901 33201
rect 19651 33160 19660 33200
rect 19700 33160 19852 33200
rect 19892 33160 19901 33200
rect 19843 33159 19901 33160
rect 1228 33076 3956 33116
rect 4003 33076 4012 33116
rect 4052 33076 11360 33116
rect 14563 33116 14621 33117
rect 16963 33116 17021 33117
rect 19651 33116 19709 33117
rect 14563 33076 14572 33116
rect 14612 33076 14668 33116
rect 14708 33076 14717 33116
rect 16878 33076 16972 33116
rect 17012 33076 17021 33116
rect 19555 33076 19564 33116
rect 19604 33076 19660 33116
rect 19700 33076 19709 33116
rect 0 33032 80 33052
rect 1228 33032 1268 33076
rect 3916 33032 3956 33076
rect 0 32992 1268 33032
rect 2275 32992 2284 33032
rect 2324 32992 2956 33032
rect 2996 32992 3005 33032
rect 3916 32992 4684 33032
rect 4724 32992 4733 33032
rect 0 32972 80 32992
rect 1315 32948 1373 32949
rect 2563 32948 2621 32949
rect 3715 32948 3773 32949
rect 5452 32948 5492 33076
rect 14563 33075 14621 33076
rect 16963 33075 17021 33076
rect 19651 33075 19709 33076
rect 17443 33032 17501 33033
rect 21424 33032 21504 33052
rect 5635 32992 5644 33032
rect 5684 32992 7756 33032
rect 7796 32992 7805 33032
rect 8035 32992 8044 33032
rect 8084 32992 11404 33032
rect 11444 32992 11453 33032
rect 17347 32992 17356 33032
rect 17396 32992 17452 33032
rect 17492 32992 17501 33032
rect 20035 32992 20044 33032
rect 20084 32992 21504 33032
rect 17443 32991 17501 32992
rect 21424 32972 21504 32992
rect 1230 32908 1324 32948
rect 1364 32908 1373 32948
rect 1699 32908 1708 32948
rect 1748 32908 2572 32948
rect 2612 32908 3724 32948
rect 3764 32908 3773 32948
rect 5443 32908 5452 32948
rect 5492 32908 5501 32948
rect 6883 32908 6892 32948
rect 6932 32908 7276 32948
rect 7316 32908 7325 32948
rect 9763 32908 9772 32948
rect 9812 32908 11884 32948
rect 11924 32908 11933 32948
rect 14659 32908 14668 32948
rect 14708 32908 19372 32948
rect 19412 32908 19421 32948
rect 1315 32907 1373 32908
rect 2563 32907 2621 32908
rect 3715 32907 3773 32908
rect 1795 32864 1853 32865
rect 4195 32864 4253 32865
rect 10147 32864 10205 32865
rect 12643 32864 12701 32865
rect 1507 32824 1516 32864
rect 1556 32824 1804 32864
rect 1844 32824 1853 32864
rect 3139 32824 3148 32864
rect 3188 32824 4204 32864
rect 4244 32824 4253 32864
rect 5251 32824 5260 32864
rect 5300 32824 5644 32864
rect 5684 32824 5693 32864
rect 7075 32824 7084 32864
rect 7124 32824 7852 32864
rect 7892 32824 7901 32864
rect 9283 32824 9292 32864
rect 9332 32824 9868 32864
rect 9908 32824 9917 32864
rect 10062 32824 10156 32864
rect 10196 32824 10205 32864
rect 12558 32824 12652 32864
rect 12692 32824 12701 32864
rect 14563 32824 14572 32864
rect 14612 32824 16436 32864
rect 16579 32824 16588 32864
rect 16628 32824 17548 32864
rect 17588 32824 17597 32864
rect 17731 32824 17740 32864
rect 17780 32824 18028 32864
rect 18068 32824 18077 32864
rect 1795 32823 1853 32824
rect 4195 32823 4253 32824
rect 10147 32823 10205 32824
rect 12643 32823 12701 32824
rect 4291 32780 4349 32781
rect 7075 32780 7133 32781
rect 16396 32780 16436 32824
rect 19939 32780 19997 32781
rect 1603 32740 1612 32780
rect 1652 32740 1900 32780
rect 1940 32740 1949 32780
rect 4291 32740 4300 32780
rect 4340 32740 6124 32780
rect 6164 32740 7084 32780
rect 7124 32740 7133 32780
rect 7363 32740 7372 32780
rect 7412 32740 8236 32780
rect 8276 32740 8285 32780
rect 13027 32740 13036 32780
rect 13076 32740 15820 32780
rect 15860 32740 15869 32780
rect 16396 32740 16684 32780
rect 16724 32740 17932 32780
rect 17972 32740 18604 32780
rect 18644 32740 18653 32780
rect 19854 32740 19948 32780
rect 19988 32740 19997 32780
rect 4291 32739 4349 32740
rect 7075 32739 7133 32740
rect 19939 32739 19997 32740
rect 6211 32696 6269 32697
rect 21424 32696 21504 32716
rect 5731 32656 5740 32696
rect 5780 32656 6220 32696
rect 6260 32656 10828 32696
rect 10868 32656 12364 32696
rect 12404 32656 12413 32696
rect 12547 32656 12556 32696
rect 12596 32656 14860 32696
rect 14900 32656 14909 32696
rect 17260 32656 21504 32696
rect 6211 32655 6269 32656
rect 8611 32612 8669 32613
rect 17260 32612 17300 32656
rect 21424 32636 21504 32656
rect 3331 32572 3340 32612
rect 3380 32572 3724 32612
rect 3764 32572 8620 32612
rect 8660 32572 8669 32612
rect 17251 32572 17260 32612
rect 17300 32572 17309 32612
rect 8611 32571 8669 32572
rect 0 32528 80 32548
rect 0 32488 2540 32528
rect 4919 32488 4928 32528
rect 4968 32488 5010 32528
rect 5050 32488 5092 32528
rect 5132 32488 5174 32528
rect 5214 32488 5256 32528
rect 5296 32488 5305 32528
rect 6787 32488 6796 32528
rect 6836 32488 7180 32528
rect 7220 32488 7229 32528
rect 15331 32488 15340 32528
rect 15380 32488 17452 32528
rect 17492 32488 18220 32528
rect 18260 32488 18269 32528
rect 20039 32488 20048 32528
rect 20088 32488 20130 32528
rect 20170 32488 20212 32528
rect 20252 32488 20294 32528
rect 20334 32488 20376 32528
rect 20416 32488 20425 32528
rect 0 32468 80 32488
rect 2500 32444 2540 32488
rect 2500 32404 2860 32444
rect 2900 32404 8468 32444
rect 16483 32404 16492 32444
rect 16532 32404 19852 32444
rect 19892 32404 19901 32444
rect 8428 32360 8468 32404
rect 16963 32360 17021 32361
rect 17443 32360 17501 32361
rect 4387 32320 4396 32360
rect 4436 32320 6220 32360
rect 6260 32320 6269 32360
rect 6892 32320 8140 32360
rect 8180 32320 8189 32360
rect 8419 32320 8428 32360
rect 8468 32320 16012 32360
rect 16052 32320 16061 32360
rect 16867 32320 16876 32360
rect 16916 32320 16972 32360
rect 17012 32320 17021 32360
rect 17358 32320 17452 32360
rect 17492 32320 17501 32360
rect 2467 32276 2525 32277
rect 6892 32276 6932 32320
rect 16963 32319 17021 32320
rect 17443 32319 17501 32320
rect 19555 32360 19613 32361
rect 21424 32360 21504 32380
rect 19555 32320 19564 32360
rect 19604 32320 21504 32360
rect 19555 32319 19613 32320
rect 21424 32300 21504 32320
rect 2467 32236 2476 32276
rect 2516 32236 5356 32276
rect 5396 32236 5405 32276
rect 6883 32236 6892 32276
rect 6932 32236 6941 32276
rect 12931 32236 12940 32276
rect 12980 32236 12989 32276
rect 2467 32235 2525 32236
rect 4675 32192 4733 32193
rect 2659 32152 2668 32192
rect 2708 32152 4492 32192
rect 4532 32152 4541 32192
rect 4675 32152 4684 32192
rect 4724 32152 4972 32192
rect 5012 32152 5021 32192
rect 6499 32152 6508 32192
rect 6548 32152 6700 32192
rect 6740 32152 6749 32192
rect 4675 32151 4733 32152
rect 6892 32108 6932 32236
rect 8611 32192 8669 32193
rect 7075 32152 7084 32192
rect 7124 32152 8140 32192
rect 8180 32152 8189 32192
rect 8526 32152 8620 32192
rect 8660 32152 9196 32192
rect 9236 32152 9245 32192
rect 11320 32152 12844 32192
rect 12884 32152 12893 32192
rect 8611 32151 8669 32152
rect 3523 32068 3532 32108
rect 3572 32068 3916 32108
rect 3956 32068 4780 32108
rect 4820 32068 6932 32108
rect 0 32024 80 32044
rect 11320 32024 11360 32152
rect 12259 32108 12317 32109
rect 12940 32108 12980 32236
rect 14179 32152 14188 32192
rect 14228 32152 15820 32192
rect 15860 32152 15869 32192
rect 13603 32108 13661 32109
rect 12259 32068 12268 32108
rect 12308 32068 12556 32108
rect 12596 32068 12605 32108
rect 12940 32068 13612 32108
rect 13652 32068 14860 32108
rect 14900 32068 14909 32108
rect 12259 32067 12317 32068
rect 13603 32067 13661 32068
rect 21424 32024 21504 32044
rect 0 31984 6028 32024
rect 6068 31984 11360 32024
rect 12835 31984 12844 32024
rect 12884 31984 13036 32024
rect 13076 31984 13085 32024
rect 20707 31984 20716 32024
rect 20756 31984 21504 32024
rect 0 31964 80 31984
rect 21424 31964 21504 31984
rect 12931 31900 12940 31940
rect 12980 31900 16108 31940
rect 16148 31900 16157 31940
rect 19555 31900 19564 31940
rect 19604 31900 21100 31940
rect 21140 31900 21149 31940
rect 2563 31816 2572 31856
rect 2612 31816 2860 31856
rect 2900 31816 2909 31856
rect 3679 31732 3688 31772
rect 3728 31732 3770 31772
rect 3810 31732 3852 31772
rect 3892 31732 3934 31772
rect 3974 31732 4016 31772
rect 4056 31732 4065 31772
rect 18799 31732 18808 31772
rect 18848 31732 18890 31772
rect 18930 31732 18972 31772
rect 19012 31732 19054 31772
rect 19094 31732 19136 31772
rect 19176 31732 19185 31772
rect 7747 31688 7805 31689
rect 21424 31688 21504 31708
rect 2467 31648 2476 31688
rect 2516 31648 3532 31688
rect 3572 31648 3581 31688
rect 6508 31648 7756 31688
rect 7796 31648 7948 31688
rect 7988 31648 7997 31688
rect 20803 31648 20812 31688
rect 20852 31648 21504 31688
rect 6508 31604 6548 31648
rect 7747 31647 7805 31648
rect 21424 31628 21504 31648
rect 7075 31604 7133 31605
rect 10627 31604 10685 31605
rect 2284 31564 6548 31604
rect 6595 31564 6604 31604
rect 6644 31564 6653 31604
rect 7075 31564 7084 31604
rect 7124 31564 8276 31604
rect 0 31520 80 31540
rect 2284 31520 2324 31564
rect 0 31480 2324 31520
rect 2371 31520 2429 31521
rect 6604 31520 6644 31564
rect 7075 31563 7133 31564
rect 2371 31480 2380 31520
rect 2420 31480 4300 31520
rect 4340 31480 4349 31520
rect 5539 31480 5548 31520
rect 5588 31480 6028 31520
rect 6068 31480 6077 31520
rect 6604 31480 6892 31520
rect 6932 31480 6941 31520
rect 7075 31480 7084 31520
rect 7124 31480 7564 31520
rect 7604 31480 7613 31520
rect 7747 31480 7756 31520
rect 7796 31480 8044 31520
rect 8084 31480 8093 31520
rect 0 31460 80 31480
rect 2371 31479 2429 31480
rect 6595 31396 6604 31436
rect 6644 31396 7660 31436
rect 7700 31396 7709 31436
rect 2659 31352 2717 31353
rect 6979 31352 7037 31353
rect 1315 31312 1324 31352
rect 1364 31312 2188 31352
rect 2228 31312 2237 31352
rect 2467 31312 2476 31352
rect 2516 31312 2668 31352
rect 2708 31312 2717 31352
rect 5923 31312 5932 31352
rect 5972 31312 5981 31352
rect 6115 31312 6124 31352
rect 6164 31312 6988 31352
rect 7028 31312 7037 31352
rect 2659 31311 2717 31312
rect 5932 31184 5972 31312
rect 6979 31311 7037 31312
rect 7948 31268 7988 31480
rect 8236 31436 8276 31564
rect 10627 31564 10636 31604
rect 10676 31564 10732 31604
rect 10772 31564 12460 31604
rect 12500 31564 13324 31604
rect 13364 31564 13373 31604
rect 19756 31564 19988 31604
rect 10627 31563 10685 31564
rect 19756 31520 19796 31564
rect 11971 31480 11980 31520
rect 12020 31480 12364 31520
rect 12404 31480 13804 31520
rect 13844 31480 13853 31520
rect 19267 31480 19276 31520
rect 19316 31480 19796 31520
rect 19843 31520 19901 31521
rect 19843 31480 19852 31520
rect 19892 31480 19901 31520
rect 19948 31520 19988 31564
rect 20515 31520 20573 31521
rect 19948 31480 20524 31520
rect 20564 31480 20573 31520
rect 19843 31479 19901 31480
rect 20515 31479 20573 31480
rect 16483 31436 16541 31437
rect 8227 31396 8236 31436
rect 8276 31396 8285 31436
rect 9859 31396 9868 31436
rect 9908 31396 11404 31436
rect 11444 31396 11453 31436
rect 16398 31396 16492 31436
rect 16532 31396 16541 31436
rect 19852 31436 19892 31479
rect 19852 31396 20180 31436
rect 16483 31395 16541 31396
rect 19843 31352 19901 31353
rect 8707 31312 8716 31352
rect 8756 31312 10540 31352
rect 10580 31312 11020 31352
rect 11060 31312 11069 31352
rect 12547 31312 12556 31352
rect 12596 31312 14092 31352
rect 14132 31312 14860 31352
rect 14900 31312 17068 31352
rect 17108 31312 17117 31352
rect 17731 31312 17740 31352
rect 17780 31312 18604 31352
rect 18644 31312 19564 31352
rect 19604 31312 19613 31352
rect 19758 31312 19852 31352
rect 19892 31312 19901 31352
rect 20140 31352 20180 31396
rect 21424 31352 21504 31372
rect 20140 31312 21504 31352
rect 17740 31268 17780 31312
rect 19843 31311 19901 31312
rect 21424 31292 21504 31312
rect 6307 31228 6316 31268
rect 6356 31228 7988 31268
rect 8611 31228 8620 31268
rect 8660 31228 14668 31268
rect 14708 31228 14717 31268
rect 16099 31228 16108 31268
rect 16148 31228 17780 31268
rect 18595 31184 18653 31185
rect 3043 31144 3052 31184
rect 3092 31144 3436 31184
rect 3476 31144 5452 31184
rect 5492 31144 5501 31184
rect 5932 31144 6028 31184
rect 6068 31144 7180 31184
rect 7220 31144 8332 31184
rect 8372 31144 8381 31184
rect 9475 31144 9484 31184
rect 9524 31144 18604 31184
rect 18644 31144 18653 31184
rect 18595 31143 18653 31144
rect 19267 31184 19325 31185
rect 19267 31144 19276 31184
rect 19316 31144 20044 31184
rect 20084 31144 20093 31184
rect 19267 31143 19325 31144
rect 1795 31060 1804 31100
rect 1844 31060 2092 31100
rect 2132 31060 2141 31100
rect 4387 31060 4396 31100
rect 4436 31060 4684 31100
rect 4724 31060 5396 31100
rect 6883 31060 6892 31100
rect 6932 31060 8716 31100
rect 8756 31060 11116 31100
rect 11156 31060 11165 31100
rect 0 31016 80 31036
rect 5356 31016 5396 31060
rect 21187 31016 21245 31017
rect 21424 31016 21504 31036
rect 0 30976 3340 31016
rect 3380 30976 3389 31016
rect 4919 30976 4928 31016
rect 4968 30976 5010 31016
rect 5050 30976 5092 31016
rect 5132 30976 5174 31016
rect 5214 30976 5256 31016
rect 5296 30976 5305 31016
rect 5356 30976 10444 31016
rect 10484 30976 10493 31016
rect 11395 30976 11404 31016
rect 11444 30976 12116 31016
rect 20039 30976 20048 31016
rect 20088 30976 20130 31016
rect 20170 30976 20212 31016
rect 20252 30976 20294 31016
rect 20334 30976 20376 31016
rect 20416 30976 20425 31016
rect 21187 30976 21196 31016
rect 21236 30976 21504 31016
rect 0 30956 80 30976
rect 12076 30932 12116 30976
rect 21187 30975 21245 30976
rect 21424 30956 21504 30976
rect 2179 30892 2188 30932
rect 2228 30892 3436 30932
rect 3476 30892 3485 30932
rect 4099 30892 4108 30932
rect 4148 30892 6316 30932
rect 6356 30892 6365 30932
rect 8803 30892 8812 30932
rect 8852 30892 11692 30932
rect 11732 30892 11741 30932
rect 12067 30892 12076 30932
rect 12116 30892 16108 30932
rect 16148 30892 16157 30932
rect 4771 30848 4829 30849
rect 7459 30848 7517 30849
rect 16675 30848 16733 30849
rect 17059 30848 17117 30849
rect 4752 30808 4780 30848
rect 4820 30808 4876 30848
rect 4916 30808 6796 30848
rect 6836 30808 6845 30848
rect 7459 30808 7468 30848
rect 7508 30808 16684 30848
rect 16724 30808 17068 30848
rect 17108 30808 18412 30848
rect 18452 30808 18461 30848
rect 4771 30807 4829 30808
rect 7459 30807 7517 30808
rect 16675 30807 16733 30808
rect 17059 30807 17117 30808
rect 13699 30724 13708 30764
rect 13748 30724 14188 30764
rect 14228 30724 15340 30764
rect 15380 30724 16820 30764
rect 19267 30724 19276 30764
rect 19316 30724 19852 30764
rect 19892 30724 19901 30764
rect 16780 30681 16820 30724
rect 7267 30680 7325 30681
rect 15715 30680 15773 30681
rect 2371 30640 2380 30680
rect 2420 30640 2572 30680
rect 2612 30640 2956 30680
rect 2996 30640 3005 30680
rect 4771 30640 4780 30680
rect 4820 30640 4972 30680
rect 5012 30640 5021 30680
rect 7267 30640 7276 30680
rect 7316 30640 7372 30680
rect 7412 30640 7421 30680
rect 13603 30640 13612 30680
rect 13652 30640 15724 30680
rect 15764 30640 15773 30680
rect 7267 30639 7325 30640
rect 15715 30639 15773 30640
rect 16771 30680 16829 30681
rect 18595 30680 18653 30681
rect 19939 30680 19997 30681
rect 21424 30680 21504 30700
rect 16771 30640 16780 30680
rect 16820 30640 16972 30680
rect 17012 30640 17021 30680
rect 18019 30640 18028 30680
rect 18068 30640 18316 30680
rect 18356 30640 18365 30680
rect 18595 30640 18604 30680
rect 18644 30640 18796 30680
rect 18836 30640 18845 30680
rect 19939 30640 19948 30680
rect 19988 30640 21504 30680
rect 16771 30639 16829 30640
rect 18595 30639 18653 30640
rect 19939 30639 19997 30640
rect 21424 30620 21504 30640
rect 14755 30556 14764 30596
rect 14804 30556 20044 30596
rect 20084 30556 20093 30596
rect 0 30512 80 30532
rect 1123 30512 1181 30513
rect 14563 30512 14621 30513
rect 0 30472 1132 30512
rect 1172 30472 1181 30512
rect 3907 30472 3916 30512
rect 3956 30472 5644 30512
rect 5684 30472 14572 30512
rect 14612 30472 14621 30512
rect 0 30452 80 30472
rect 1123 30471 1181 30472
rect 14563 30471 14621 30472
rect 4387 30388 4396 30428
rect 4436 30388 4972 30428
rect 5012 30388 5021 30428
rect 20227 30388 20236 30428
rect 20276 30388 21292 30428
rect 21332 30388 21341 30428
rect 19651 30344 19709 30345
rect 21424 30344 21504 30364
rect 19651 30304 19660 30344
rect 19700 30304 21504 30344
rect 19651 30303 19709 30304
rect 21424 30284 21504 30304
rect 1699 30260 1757 30261
rect 14755 30260 14813 30261
rect 19939 30260 19997 30261
rect 1699 30220 1708 30260
rect 1748 30220 3572 30260
rect 3679 30220 3688 30260
rect 3728 30220 3770 30260
rect 3810 30220 3852 30260
rect 3892 30220 3934 30260
rect 3974 30220 4016 30260
rect 4056 30220 4065 30260
rect 5635 30220 5644 30260
rect 5684 30220 6220 30260
rect 6260 30220 6269 30260
rect 11491 30220 11500 30260
rect 11540 30220 12460 30260
rect 12500 30220 12509 30260
rect 14755 30220 14764 30260
rect 14804 30220 14956 30260
rect 14996 30220 15005 30260
rect 18799 30220 18808 30260
rect 18848 30220 18890 30260
rect 18930 30220 18972 30260
rect 19012 30220 19054 30260
rect 19094 30220 19136 30260
rect 19176 30220 19185 30260
rect 19555 30220 19564 30260
rect 19604 30220 19948 30260
rect 19988 30220 19997 30260
rect 1699 30219 1757 30220
rect 3532 30176 3572 30220
rect 5644 30176 5684 30220
rect 14755 30219 14813 30220
rect 19939 30219 19997 30220
rect 2467 30136 2476 30176
rect 2516 30136 2668 30176
rect 2708 30136 3340 30176
rect 3380 30136 3389 30176
rect 3532 30136 5684 30176
rect 15619 30136 15628 30176
rect 15668 30136 19756 30176
rect 19796 30136 19805 30176
rect 2275 30052 2284 30092
rect 2324 30052 2860 30092
rect 2900 30052 2909 30092
rect 5731 30052 5740 30092
rect 5780 30052 6220 30092
rect 6260 30052 6269 30092
rect 14947 30052 14956 30092
rect 14996 30052 18796 30092
rect 18836 30052 18845 30092
rect 0 30008 80 30028
rect 21424 30008 21504 30028
rect 0 29968 6316 30008
rect 6356 29968 6365 30008
rect 7363 29968 7372 30008
rect 7412 29968 7852 30008
rect 7892 29968 8428 30008
rect 8468 29968 8477 30008
rect 10435 29968 10444 30008
rect 10484 29968 11884 30008
rect 11924 29968 11933 30008
rect 16291 29968 16300 30008
rect 16340 29968 21504 30008
rect 0 29948 80 29968
rect 21424 29948 21504 29968
rect 7075 29924 7133 29925
rect 17731 29924 17789 29925
rect 7075 29884 7084 29924
rect 7124 29884 7468 29924
rect 7508 29884 8044 29924
rect 8084 29884 8093 29924
rect 12163 29884 12172 29924
rect 12212 29884 16108 29924
rect 16148 29884 16157 29924
rect 17731 29884 17740 29924
rect 17780 29884 19756 29924
rect 19796 29884 19805 29924
rect 7075 29883 7133 29884
rect 17731 29883 17789 29884
rect 2659 29840 2717 29841
rect 17539 29840 17597 29841
rect 17827 29840 17885 29841
rect 1315 29800 1324 29840
rect 1364 29800 1516 29840
rect 1556 29800 1565 29840
rect 2467 29800 2476 29840
rect 2516 29800 2668 29840
rect 2708 29800 2717 29840
rect 3336 29800 3345 29840
rect 3385 29800 3628 29840
rect 3668 29800 3677 29840
rect 6403 29800 6412 29840
rect 6452 29800 7276 29840
rect 7316 29800 8236 29840
rect 8276 29800 10060 29840
rect 10100 29800 10109 29840
rect 13987 29800 13996 29840
rect 14036 29800 17260 29840
rect 17300 29800 17548 29840
rect 17588 29800 17597 29840
rect 17731 29800 17740 29840
rect 17780 29800 17836 29840
rect 17876 29800 17885 29840
rect 2659 29799 2717 29800
rect 17539 29799 17597 29800
rect 17827 29799 17885 29800
rect 7171 29756 7229 29757
rect 15427 29756 15485 29757
rect 6307 29716 6316 29756
rect 6356 29716 7180 29756
rect 7220 29716 15436 29756
rect 15476 29716 15485 29756
rect 7171 29715 7229 29716
rect 15427 29715 15485 29716
rect 21424 29672 21504 29692
rect 3139 29632 3148 29672
rect 3188 29632 3916 29672
rect 3956 29632 3965 29672
rect 12451 29632 12460 29672
rect 12500 29632 15244 29672
rect 15284 29632 15293 29672
rect 19939 29632 19948 29672
rect 19988 29632 20812 29672
rect 20852 29632 20861 29672
rect 21187 29632 21196 29672
rect 21236 29632 21504 29672
rect 21424 29612 21504 29632
rect 4195 29548 4204 29588
rect 4244 29548 19660 29588
rect 19700 29548 19709 29588
rect 0 29504 80 29524
rect 1699 29504 1757 29505
rect 0 29464 1708 29504
rect 1748 29464 1757 29504
rect 4919 29464 4928 29504
rect 4968 29464 5010 29504
rect 5050 29464 5092 29504
rect 5132 29464 5174 29504
rect 5214 29464 5256 29504
rect 5296 29464 5305 29504
rect 11875 29464 11884 29504
rect 11924 29464 18316 29504
rect 18356 29464 18365 29504
rect 20039 29464 20048 29504
rect 20088 29464 20130 29504
rect 20170 29464 20212 29504
rect 20252 29464 20294 29504
rect 20334 29464 20376 29504
rect 20416 29464 20425 29504
rect 0 29444 80 29464
rect 1699 29463 1757 29464
rect 3811 29380 3820 29420
rect 3860 29380 4780 29420
rect 4820 29380 4829 29420
rect 5347 29380 5356 29420
rect 5396 29380 11924 29420
rect 11971 29380 11980 29420
rect 12020 29380 12980 29420
rect 13891 29380 13900 29420
rect 13940 29380 14380 29420
rect 14420 29380 14429 29420
rect 14851 29380 14860 29420
rect 14900 29380 16492 29420
rect 16532 29380 16541 29420
rect 11884 29336 11924 29380
rect 12835 29336 12893 29337
rect 1795 29296 1804 29336
rect 1844 29296 10348 29336
rect 10388 29296 10397 29336
rect 11884 29296 12844 29336
rect 12884 29296 12893 29336
rect 12940 29336 12980 29380
rect 18307 29336 18365 29337
rect 20803 29336 20861 29337
rect 21424 29336 21504 29356
rect 12940 29296 14228 29336
rect 15427 29296 15436 29336
rect 15476 29296 17356 29336
rect 17396 29296 17405 29336
rect 18307 29296 18316 29336
rect 18356 29296 18508 29336
rect 18548 29296 18557 29336
rect 18691 29296 18700 29336
rect 18740 29296 19948 29336
rect 19988 29296 19997 29336
rect 20803 29296 20812 29336
rect 20852 29296 21504 29336
rect 12835 29295 12893 29296
rect 5443 29252 5501 29253
rect 14188 29252 14228 29296
rect 18307 29295 18365 29296
rect 20803 29295 20861 29296
rect 21424 29276 21504 29296
rect 2755 29212 2764 29252
rect 2804 29212 3532 29252
rect 3572 29212 5068 29252
rect 5108 29212 5117 29252
rect 5443 29212 5452 29252
rect 5492 29212 6836 29252
rect 6883 29212 6892 29252
rect 6932 29212 13804 29252
rect 13844 29212 13853 29252
rect 14188 29212 15820 29252
rect 15860 29212 18548 29252
rect 5443 29211 5501 29212
rect 6796 29168 6836 29212
rect 18508 29168 18548 29212
rect 2500 29128 6124 29168
rect 6164 29128 6173 29168
rect 6796 29128 6988 29168
rect 7028 29128 7037 29168
rect 8995 29128 9004 29168
rect 9044 29128 9580 29168
rect 9620 29128 9964 29168
rect 10004 29128 11596 29168
rect 11636 29128 12076 29168
rect 12116 29128 12125 29168
rect 13219 29128 13228 29168
rect 13268 29128 13996 29168
rect 14036 29128 14045 29168
rect 14092 29128 16588 29168
rect 16628 29128 16637 29168
rect 18499 29128 18508 29168
rect 18548 29128 18557 29168
rect 2275 29084 2333 29085
rect 2500 29084 2540 29128
rect 14092 29084 14132 29128
rect 460 29044 2228 29084
rect 0 29000 80 29020
rect 460 29000 500 29044
rect 0 28960 500 29000
rect 2188 29000 2228 29044
rect 2275 29044 2284 29084
rect 2324 29044 2540 29084
rect 2668 29044 5492 29084
rect 5539 29044 5548 29084
rect 5588 29044 5780 29084
rect 10339 29044 10348 29084
rect 10388 29044 14132 29084
rect 14476 29044 14860 29084
rect 14900 29044 14909 29084
rect 19555 29044 19564 29084
rect 19604 29044 20908 29084
rect 20948 29044 20957 29084
rect 2275 29043 2333 29044
rect 2668 29000 2708 29044
rect 5452 29000 5492 29044
rect 2188 28960 2708 29000
rect 5412 28960 5452 29000
rect 5492 28960 5501 29000
rect 0 28940 80 28960
rect 5740 28916 5780 29044
rect 14476 29000 14516 29044
rect 11683 28960 11692 29000
rect 11732 28960 11884 29000
rect 11924 28960 11933 29000
rect 13987 28960 13996 29000
rect 14036 28960 14516 29000
rect 20995 29000 21053 29001
rect 21424 29000 21504 29020
rect 20995 28960 21004 29000
rect 21044 28960 21504 29000
rect 20995 28959 21053 28960
rect 21424 28940 21504 28960
rect 18307 28916 18365 28917
rect 1891 28876 1900 28916
rect 1940 28876 2540 28916
rect 5740 28876 5932 28916
rect 5972 28876 5981 28916
rect 16291 28876 16300 28916
rect 16340 28876 16684 28916
rect 16724 28876 16733 28916
rect 16876 28876 17836 28916
rect 17876 28876 18316 28916
rect 18356 28876 18365 28916
rect 2500 28832 2540 28876
rect 16876 28832 16916 28876
rect 18307 28875 18365 28876
rect 2500 28792 8716 28832
rect 8756 28792 8765 28832
rect 14371 28792 14380 28832
rect 14420 28792 16916 28832
rect 6691 28748 6749 28749
rect 11491 28748 11549 28749
rect 3679 28708 3688 28748
rect 3728 28708 3770 28748
rect 3810 28708 3852 28748
rect 3892 28708 3934 28748
rect 3974 28708 4016 28748
rect 4056 28708 4065 28748
rect 6691 28708 6700 28748
rect 6740 28708 11500 28748
rect 11540 28708 11549 28748
rect 18799 28708 18808 28748
rect 18848 28708 18890 28748
rect 18930 28708 18972 28748
rect 19012 28708 19054 28748
rect 19094 28708 19136 28748
rect 19176 28708 19185 28748
rect 6691 28707 6749 28708
rect 11491 28707 11549 28708
rect 18403 28664 18461 28665
rect 21424 28664 21504 28684
rect 8899 28624 8908 28664
rect 8948 28624 9484 28664
rect 9524 28624 9533 28664
rect 18403 28624 18412 28664
rect 18452 28624 21504 28664
rect 18403 28623 18461 28624
rect 21424 28604 21504 28624
rect 4675 28540 4684 28580
rect 4724 28540 7948 28580
rect 7988 28540 7997 28580
rect 9091 28540 9100 28580
rect 9140 28540 9388 28580
rect 9428 28540 9437 28580
rect 13900 28540 18124 28580
rect 18164 28540 18796 28580
rect 18836 28540 18845 28580
rect 19843 28540 19852 28580
rect 19892 28540 21196 28580
rect 21236 28540 21245 28580
rect 0 28496 80 28516
rect 7459 28496 7517 28497
rect 0 28456 7468 28496
rect 7508 28456 7517 28496
rect 0 28436 80 28456
rect 7459 28455 7517 28456
rect 7747 28412 7805 28413
rect 2755 28372 2764 28412
rect 2804 28372 3340 28412
rect 3380 28372 3389 28412
rect 5347 28372 5356 28412
rect 5396 28372 6700 28412
rect 6740 28372 6749 28412
rect 7662 28372 7756 28412
rect 7796 28372 7805 28412
rect 7948 28412 7988 28540
rect 13900 28496 13940 28540
rect 15427 28496 15485 28497
rect 8899 28456 8908 28496
rect 8948 28456 9196 28496
rect 9236 28456 9245 28496
rect 10243 28456 10252 28496
rect 10292 28456 11020 28496
rect 11060 28456 11069 28496
rect 11203 28456 11212 28496
rect 11252 28456 13900 28496
rect 13940 28456 13949 28496
rect 15235 28456 15244 28496
rect 15284 28456 15436 28496
rect 15476 28456 15532 28496
rect 15572 28456 15600 28496
rect 16867 28456 16876 28496
rect 16916 28456 17548 28496
rect 17588 28456 17597 28496
rect 15427 28455 15485 28456
rect 19267 28412 19325 28413
rect 7948 28372 11252 28412
rect 11875 28372 11884 28412
rect 11924 28372 19276 28412
rect 19316 28372 19325 28412
rect 2947 28288 2956 28328
rect 2996 28288 3628 28328
rect 3668 28288 3677 28328
rect 835 28204 844 28244
rect 884 28204 5356 28244
rect 5396 28204 5405 28244
rect 3331 28120 3340 28160
rect 3380 28120 4012 28160
rect 4052 28120 4061 28160
rect 5452 28076 5492 28372
rect 7747 28371 7805 28372
rect 11212 28328 11252 28372
rect 19267 28371 19325 28372
rect 17827 28328 17885 28329
rect 18019 28328 18077 28329
rect 5923 28288 5932 28328
rect 5972 28288 8236 28328
rect 8276 28288 8285 28328
rect 11203 28288 11212 28328
rect 11252 28288 11261 28328
rect 13411 28288 13420 28328
rect 13460 28288 17836 28328
rect 17876 28288 17885 28328
rect 17934 28288 18028 28328
rect 18068 28288 18077 28328
rect 17827 28287 17885 28288
rect 18019 28287 18077 28288
rect 18499 28328 18557 28329
rect 21424 28328 21504 28348
rect 18499 28288 18508 28328
rect 18548 28288 21504 28328
rect 18499 28287 18557 28288
rect 21424 28268 21504 28288
rect 18115 28244 18173 28245
rect 18307 28244 18365 28245
rect 15331 28204 15340 28244
rect 15380 28204 16396 28244
rect 16436 28204 16445 28244
rect 18030 28204 18124 28244
rect 18164 28204 18316 28244
rect 18356 28204 18365 28244
rect 18115 28203 18173 28204
rect 18307 28203 18365 28204
rect 17059 28120 17068 28160
rect 17108 28120 19276 28160
rect 19316 28120 19325 28160
rect 19651 28120 19660 28160
rect 19700 28120 20716 28160
rect 20756 28120 20765 28160
rect 2500 28036 5492 28076
rect 9283 28036 9292 28076
rect 9332 28036 19756 28076
rect 19796 28036 19805 28076
rect 0 27992 80 28012
rect 2500 27992 2540 28036
rect 21424 27992 21504 28012
rect 0 27952 2540 27992
rect 4919 27952 4928 27992
rect 4968 27952 5010 27992
rect 5050 27952 5092 27992
rect 5132 27952 5174 27992
rect 5214 27952 5256 27992
rect 5296 27952 5305 27992
rect 16483 27952 16492 27992
rect 16532 27952 18028 27992
rect 18068 27952 18077 27992
rect 20039 27952 20048 27992
rect 20088 27952 20130 27992
rect 20170 27952 20212 27992
rect 20252 27952 20294 27992
rect 20334 27952 20376 27992
rect 20416 27952 20425 27992
rect 21091 27952 21100 27992
rect 21140 27952 21504 27992
rect 0 27932 80 27952
rect 21424 27932 21504 27952
rect 16675 27908 16733 27909
rect 16590 27868 16684 27908
rect 16724 27868 16733 27908
rect 17059 27868 17068 27908
rect 17108 27868 17932 27908
rect 17972 27868 17981 27908
rect 19171 27868 19180 27908
rect 19220 27868 19756 27908
rect 19796 27868 19805 27908
rect 16675 27867 16733 27868
rect 6211 27824 6269 27825
rect 6126 27784 6220 27824
rect 6260 27784 6269 27824
rect 10531 27784 10540 27824
rect 10580 27784 10620 27824
rect 17251 27784 17260 27824
rect 17300 27784 20812 27824
rect 20852 27784 20861 27824
rect 6211 27783 6269 27784
rect 3139 27740 3197 27741
rect 7171 27740 7229 27741
rect 10540 27740 10580 27784
rect 11011 27740 11069 27741
rect 19939 27740 19997 27741
rect 3139 27700 3148 27740
rect 3188 27700 3436 27740
rect 3476 27700 3485 27740
rect 3907 27700 3916 27740
rect 3956 27700 7180 27740
rect 7220 27700 7229 27740
rect 8707 27700 8716 27740
rect 8756 27700 9332 27740
rect 9859 27700 9868 27740
rect 9908 27700 10732 27740
rect 10772 27700 10781 27740
rect 11011 27700 11020 27740
rect 11060 27700 11212 27740
rect 11252 27700 11261 27740
rect 12163 27700 12172 27740
rect 12212 27700 19468 27740
rect 19508 27700 19517 27740
rect 19651 27700 19660 27740
rect 19700 27700 19948 27740
rect 19988 27700 19997 27740
rect 3139 27699 3197 27700
rect 7171 27699 7229 27700
rect 1987 27616 1996 27656
rect 2036 27616 2188 27656
rect 2228 27616 2572 27656
rect 2612 27616 2621 27656
rect 3523 27616 3532 27656
rect 3572 27616 6988 27656
rect 7028 27616 7660 27656
rect 7700 27616 7709 27656
rect 3043 27572 3101 27573
rect 9292 27572 9332 27700
rect 11011 27699 11069 27700
rect 19939 27699 19997 27700
rect 14563 27656 14621 27657
rect 21424 27656 21504 27676
rect 10051 27616 10060 27656
rect 10100 27616 10540 27656
rect 10580 27616 10589 27656
rect 13027 27616 13036 27656
rect 13076 27616 13996 27656
rect 14036 27616 14045 27656
rect 14478 27616 14572 27656
rect 14612 27616 14621 27656
rect 16483 27616 16492 27656
rect 16532 27616 18988 27656
rect 19028 27616 19037 27656
rect 20899 27616 20908 27656
rect 20948 27616 21504 27656
rect 14563 27615 14621 27616
rect 21424 27596 21504 27616
rect 2958 27532 3052 27572
rect 3092 27532 6164 27572
rect 6211 27532 6220 27572
rect 6260 27532 6796 27572
rect 6836 27532 6845 27572
rect 9283 27532 9292 27572
rect 9332 27532 9341 27572
rect 16003 27532 16012 27572
rect 16052 27532 18316 27572
rect 18356 27532 18365 27572
rect 3043 27531 3101 27532
rect 0 27488 80 27508
rect 5347 27488 5405 27489
rect 0 27448 5356 27488
rect 5396 27448 5405 27488
rect 6124 27488 6164 27532
rect 17731 27488 17789 27489
rect 6124 27448 6892 27488
rect 6932 27448 6941 27488
rect 7267 27448 7276 27488
rect 7316 27448 17740 27488
rect 17780 27448 17789 27488
rect 0 27428 80 27448
rect 5347 27447 5405 27448
rect 17731 27447 17789 27448
rect 10147 27404 10205 27405
rect 7459 27364 7468 27404
rect 7508 27364 8044 27404
rect 8084 27364 8093 27404
rect 9187 27364 9196 27404
rect 9236 27364 10156 27404
rect 10196 27364 10205 27404
rect 12067 27364 12076 27404
rect 12116 27364 14284 27404
rect 14324 27364 16108 27404
rect 16148 27364 16157 27404
rect 17443 27364 17452 27404
rect 17492 27364 18124 27404
rect 18164 27364 18173 27404
rect 10147 27363 10205 27364
rect 21424 27320 21504 27340
rect 10915 27280 10924 27320
rect 10964 27280 11116 27320
rect 11156 27280 11165 27320
rect 20611 27280 20620 27320
rect 20660 27280 21504 27320
rect 21424 27260 21504 27280
rect 1699 27196 1708 27236
rect 1748 27196 2188 27236
rect 2228 27196 2860 27236
rect 2900 27196 2909 27236
rect 3679 27196 3688 27236
rect 3728 27196 3770 27236
rect 3810 27196 3852 27236
rect 3892 27196 3934 27236
rect 3974 27196 4016 27236
rect 4056 27196 4065 27236
rect 10243 27196 10252 27236
rect 10292 27196 11020 27236
rect 11060 27196 11069 27236
rect 14467 27196 14476 27236
rect 14516 27196 14764 27236
rect 14804 27196 14813 27236
rect 18799 27196 18808 27236
rect 18848 27196 18890 27236
rect 18930 27196 18972 27236
rect 19012 27196 19054 27236
rect 19094 27196 19136 27236
rect 19176 27196 19185 27236
rect 2467 27112 2476 27152
rect 2516 27112 2668 27152
rect 2708 27112 2717 27152
rect 13891 27068 13949 27069
rect 1699 27028 1708 27068
rect 1748 27028 4780 27068
rect 4820 27028 4829 27068
rect 5539 27028 5548 27068
rect 5588 27028 5932 27068
rect 5972 27028 5981 27068
rect 7075 27028 7084 27068
rect 7124 27028 7564 27068
rect 7604 27028 7613 27068
rect 13891 27028 13900 27068
rect 13940 27028 15340 27068
rect 15380 27028 15389 27068
rect 13891 27027 13949 27028
rect 0 26984 80 27004
rect 21424 26984 21504 27004
rect 0 26944 9100 26984
rect 9140 26944 9484 26984
rect 9524 26944 9533 26984
rect 13123 26944 13132 26984
rect 13172 26944 13612 26984
rect 13652 26944 13661 26984
rect 14275 26944 14284 26984
rect 14324 26944 14956 26984
rect 14996 26944 15005 26984
rect 20995 26944 21004 26984
rect 21044 26944 21504 26984
rect 0 26924 80 26944
rect 21424 26924 21504 26944
rect 17635 26900 17693 26901
rect 2500 26860 3148 26900
rect 3188 26860 6508 26900
rect 6548 26860 6557 26900
rect 17155 26860 17164 26900
rect 17204 26860 17644 26900
rect 17684 26860 17693 26900
rect 2500 26816 2540 26860
rect 17635 26859 17693 26860
rect 10147 26816 10205 26817
rect 1219 26776 1228 26816
rect 1268 26776 1804 26816
rect 1844 26776 1853 26816
rect 2467 26776 2476 26816
rect 2516 26776 2540 26816
rect 2851 26776 2860 26816
rect 2900 26776 4492 26816
rect 4532 26776 4541 26816
rect 4771 26776 4780 26816
rect 4820 26776 4829 26816
rect 5731 26776 5740 26816
rect 5780 26776 6700 26816
rect 6740 26776 6749 26816
rect 10147 26776 10156 26816
rect 10196 26776 10828 26816
rect 10868 26776 10877 26816
rect 12067 26776 12076 26816
rect 12116 26776 12125 26816
rect 13219 26776 13228 26816
rect 13268 26776 13612 26816
rect 13652 26776 13661 26816
rect 14947 26776 14956 26816
rect 14996 26776 17644 26816
rect 17684 26776 17836 26816
rect 17876 26776 17885 26816
rect 4780 26732 4820 26776
rect 10147 26775 10205 26776
rect 12076 26732 12116 26776
rect 18211 26732 18269 26733
rect 67 26692 76 26732
rect 116 26692 2540 26732
rect 4780 26692 5932 26732
rect 5972 26692 6124 26732
rect 6164 26692 6173 26732
rect 9475 26692 9484 26732
rect 9524 26692 10156 26732
rect 10196 26692 10348 26732
rect 10388 26692 12116 26732
rect 15628 26692 18220 26732
rect 18260 26692 19948 26732
rect 19988 26692 19997 26732
rect 2500 26564 2540 26692
rect 15628 26648 15668 26692
rect 18211 26691 18269 26692
rect 21424 26648 21504 26668
rect 5827 26608 5836 26648
rect 5876 26608 15628 26648
rect 15668 26608 15677 26648
rect 18307 26608 18316 26648
rect 18356 26608 20044 26648
rect 20084 26608 20093 26648
rect 20803 26608 20812 26648
rect 20852 26608 21504 26648
rect 21424 26588 21504 26608
rect 6211 26564 6269 26565
rect 18595 26564 18653 26565
rect 2500 26524 6124 26564
rect 6164 26524 6220 26564
rect 6260 26524 6269 26564
rect 6691 26524 6700 26564
rect 6740 26524 7372 26564
rect 7412 26524 9484 26564
rect 9524 26524 9533 26564
rect 10819 26524 10828 26564
rect 10868 26524 11360 26564
rect 18403 26524 18412 26564
rect 18452 26524 18604 26564
rect 18644 26524 18653 26564
rect 6211 26523 6269 26524
rect 0 26480 80 26500
rect 8332 26480 8372 26524
rect 0 26440 76 26480
rect 116 26440 125 26480
rect 2851 26440 2860 26480
rect 2900 26440 4108 26480
rect 4148 26440 4684 26480
rect 4724 26440 4733 26480
rect 4919 26440 4928 26480
rect 4968 26440 5010 26480
rect 5050 26440 5092 26480
rect 5132 26440 5174 26480
rect 5214 26440 5256 26480
rect 5296 26440 5305 26480
rect 6307 26440 6316 26480
rect 6356 26440 7276 26480
rect 7316 26440 7325 26480
rect 7651 26440 7660 26480
rect 7700 26440 7852 26480
rect 7892 26440 7901 26480
rect 8323 26440 8332 26480
rect 8372 26440 8381 26480
rect 0 26420 80 26440
rect 10915 26356 10924 26396
rect 10964 26356 11212 26396
rect 11252 26356 11261 26396
rect 11320 26312 11360 26524
rect 18595 26523 18653 26524
rect 14659 26480 14717 26481
rect 11971 26440 11980 26480
rect 12020 26440 12556 26480
rect 12596 26440 12605 26480
rect 14574 26440 14668 26480
rect 14708 26440 14717 26480
rect 17827 26440 17836 26480
rect 17876 26440 18220 26480
rect 18260 26440 18269 26480
rect 20039 26440 20048 26480
rect 20088 26440 20130 26480
rect 20170 26440 20212 26480
rect 20252 26440 20294 26480
rect 20334 26440 20376 26480
rect 20416 26440 20425 26480
rect 14659 26439 14717 26440
rect 13891 26356 13900 26396
rect 13940 26356 14860 26396
rect 14900 26356 14909 26396
rect 17923 26356 17932 26396
rect 17972 26356 18316 26396
rect 18356 26356 18700 26396
rect 18740 26356 19564 26396
rect 19604 26356 19613 26396
rect 14563 26312 14621 26313
rect 8995 26272 9004 26312
rect 9044 26272 10828 26312
rect 10868 26272 10877 26312
rect 11320 26272 14572 26312
rect 14612 26272 14621 26312
rect 14563 26271 14621 26272
rect 14755 26312 14813 26313
rect 21424 26312 21504 26332
rect 14755 26272 14764 26312
rect 14804 26272 15244 26312
rect 15284 26272 15293 26312
rect 19843 26272 19852 26312
rect 19892 26272 21504 26312
rect 14755 26271 14813 26272
rect 21424 26252 21504 26272
rect 3235 26228 3293 26229
rect 4099 26228 4157 26229
rect 3235 26188 3244 26228
rect 3284 26188 3340 26228
rect 3380 26188 3389 26228
rect 3619 26188 3628 26228
rect 3668 26188 4108 26228
rect 4148 26188 4157 26228
rect 4291 26188 4300 26228
rect 4340 26188 4876 26228
rect 4916 26188 4925 26228
rect 5059 26188 5068 26228
rect 5108 26188 19756 26228
rect 19796 26188 19805 26228
rect 3235 26187 3293 26188
rect 4099 26187 4157 26188
rect 6691 26144 6749 26145
rect 13795 26144 13853 26145
rect 3427 26104 3436 26144
rect 3476 26104 6220 26144
rect 6260 26104 6269 26144
rect 6691 26104 6700 26144
rect 6740 26104 6796 26144
rect 6836 26104 7084 26144
rect 7124 26104 7133 26144
rect 10435 26104 10444 26144
rect 10484 26104 12076 26144
rect 12116 26104 13708 26144
rect 13748 26104 13804 26144
rect 13844 26104 13900 26144
rect 13940 26104 13968 26144
rect 14851 26104 14860 26144
rect 14900 26104 17260 26144
rect 17300 26104 17309 26144
rect 18499 26104 18508 26144
rect 18548 26104 18796 26144
rect 18836 26104 18845 26144
rect 6691 26103 6749 26104
rect 13795 26103 13853 26104
rect 4291 26060 4349 26061
rect 3907 26020 3916 26060
rect 3956 26020 4300 26060
rect 4340 26020 4349 26060
rect 4291 26019 4349 26020
rect 5347 26060 5405 26061
rect 11875 26060 11933 26061
rect 17731 26060 17789 26061
rect 5347 26020 5356 26060
rect 5396 26020 5452 26060
rect 5492 26020 5501 26060
rect 8611 26020 8620 26060
rect 8660 26020 8669 26060
rect 10819 26020 10828 26060
rect 10868 26020 11884 26060
rect 11924 26020 11933 26060
rect 13507 26020 13516 26060
rect 13556 26020 13804 26060
rect 13844 26020 13853 26060
rect 17731 26020 17740 26060
rect 17780 26020 17932 26060
rect 17972 26020 17981 26060
rect 5347 26019 5405 26020
rect 0 25976 80 25996
rect 1603 25976 1661 25977
rect 4300 25976 4340 26019
rect 8620 25976 8660 26020
rect 11875 26019 11933 26020
rect 17731 26019 17789 26020
rect 21424 25976 21504 25996
rect 0 25936 1516 25976
rect 1556 25936 1612 25976
rect 1652 25936 1680 25976
rect 4300 25936 6604 25976
rect 6644 25936 8140 25976
rect 8180 25936 8189 25976
rect 8323 25936 8332 25976
rect 8372 25936 8660 25976
rect 20707 25936 20716 25976
rect 20756 25936 21504 25976
rect 0 25916 80 25936
rect 1603 25935 1661 25936
rect 21424 25916 21504 25936
rect 3811 25852 3820 25892
rect 3860 25852 3869 25892
rect 4387 25852 4396 25892
rect 4436 25852 6796 25892
rect 6836 25852 8716 25892
rect 8756 25852 8765 25892
rect 10627 25852 10636 25892
rect 10676 25852 10828 25892
rect 10868 25852 10877 25892
rect 16291 25852 16300 25892
rect 16340 25852 16492 25892
rect 16532 25852 16541 25892
rect 3820 25808 3860 25852
rect 163 25768 172 25808
rect 212 25768 4204 25808
rect 4244 25768 4253 25808
rect 6892 25768 14860 25808
rect 14900 25768 14909 25808
rect 3679 25684 3688 25724
rect 3728 25684 3770 25724
rect 3810 25684 3852 25724
rect 3892 25684 3934 25724
rect 3974 25684 4016 25724
rect 4056 25684 4065 25724
rect 3139 25516 3148 25556
rect 3188 25516 3340 25556
rect 3380 25516 3389 25556
rect 0 25472 80 25492
rect 6892 25472 6932 25768
rect 16483 25724 16541 25725
rect 0 25432 1420 25472
rect 1460 25432 6932 25472
rect 8332 25684 16492 25724
rect 16532 25684 16541 25724
rect 18799 25684 18808 25724
rect 18848 25684 18890 25724
rect 18930 25684 18972 25724
rect 19012 25684 19054 25724
rect 19094 25684 19136 25724
rect 19176 25684 19185 25724
rect 19363 25684 19372 25724
rect 19412 25684 19421 25724
rect 0 25412 80 25432
rect 8332 25388 8372 25684
rect 16483 25683 16541 25684
rect 8707 25600 8716 25640
rect 8756 25600 11500 25640
rect 11540 25600 11884 25640
rect 11924 25600 11933 25640
rect 12259 25600 12268 25640
rect 12308 25600 12460 25640
rect 12500 25600 12509 25640
rect 16099 25600 16108 25640
rect 16148 25600 16300 25640
rect 16340 25600 17644 25640
rect 17684 25600 17693 25640
rect 19372 25556 19412 25684
rect 21424 25640 21504 25660
rect 20515 25600 20524 25640
rect 20564 25600 21504 25640
rect 21424 25580 21504 25600
rect 8803 25516 8812 25556
rect 8852 25516 19412 25556
rect 3043 25348 3052 25388
rect 3092 25348 3724 25388
rect 3764 25348 3773 25388
rect 5443 25348 5452 25388
rect 5492 25348 8372 25388
rect 8800 25432 11360 25472
rect 13795 25432 13804 25472
rect 13844 25432 14764 25472
rect 14804 25432 15052 25472
rect 15092 25432 15101 25472
rect 17635 25432 17644 25472
rect 17684 25432 18316 25472
rect 18356 25432 19180 25472
rect 19220 25432 19229 25472
rect 19843 25432 19852 25472
rect 19892 25432 20812 25472
rect 20852 25432 20861 25472
rect 6211 25304 6269 25305
rect 3811 25264 3820 25304
rect 3860 25264 5644 25304
rect 5684 25264 6220 25304
rect 6260 25264 6269 25304
rect 6211 25263 6269 25264
rect 6499 25304 6557 25305
rect 7939 25304 7997 25305
rect 8800 25304 8840 25432
rect 11320 25388 11360 25432
rect 6499 25264 6508 25304
rect 6548 25264 7180 25304
rect 7220 25264 7229 25304
rect 7555 25264 7564 25304
rect 7604 25264 7948 25304
rect 7988 25264 7997 25304
rect 8131 25264 8140 25304
rect 8180 25264 8840 25304
rect 9292 25348 10924 25388
rect 10964 25348 10973 25388
rect 11320 25348 11404 25388
rect 11444 25348 11453 25388
rect 12643 25348 12652 25388
rect 12692 25348 19660 25388
rect 19700 25348 19709 25388
rect 6499 25263 6557 25264
rect 7939 25263 7997 25264
rect 6019 25220 6077 25221
rect 9292 25220 9332 25348
rect 16579 25304 16637 25305
rect 21424 25304 21504 25324
rect 14179 25264 14188 25304
rect 14228 25264 14476 25304
rect 14516 25264 14525 25304
rect 16579 25264 16588 25304
rect 16628 25264 18028 25304
rect 18068 25264 18077 25304
rect 20140 25264 21504 25304
rect 16579 25263 16637 25264
rect 14275 25220 14333 25221
rect 20140 25220 20180 25264
rect 21424 25244 21504 25264
rect 6019 25180 6028 25220
rect 6068 25180 9332 25220
rect 10531 25180 10540 25220
rect 10580 25180 11500 25220
rect 11540 25180 11549 25220
rect 11596 25180 11692 25220
rect 11732 25180 11741 25220
rect 14190 25180 14284 25220
rect 14324 25180 14333 25220
rect 18787 25180 18796 25220
rect 18836 25180 20180 25220
rect 6019 25179 6077 25180
rect 11596 25136 11636 25180
rect 14275 25179 14333 25180
rect 6115 25096 6124 25136
rect 6164 25096 7852 25136
rect 7892 25096 7901 25136
rect 11395 25096 11404 25136
rect 11444 25096 11636 25136
rect 15427 25096 15436 25136
rect 15476 25096 19372 25136
rect 19412 25096 19421 25136
rect 19468 25096 20044 25136
rect 20084 25096 20093 25136
rect 19468 25052 19508 25096
rect 1603 25012 1612 25052
rect 1652 25012 2092 25052
rect 2132 25012 2141 25052
rect 11683 25012 11692 25052
rect 11732 25012 19508 25052
rect 19555 25012 19564 25052
rect 19604 25012 20852 25052
rect 0 24968 80 24988
rect 6403 24968 6461 24969
rect 16483 24968 16541 24969
rect 20812 24968 20852 25012
rect 21424 24968 21504 24988
rect 0 24928 2380 24968
rect 2420 24928 2429 24968
rect 4919 24928 4928 24968
rect 4968 24928 5010 24968
rect 5050 24928 5092 24968
rect 5132 24928 5174 24968
rect 5214 24928 5256 24968
rect 5296 24928 5305 24968
rect 6211 24928 6220 24968
rect 6260 24928 6412 24968
rect 6452 24928 6461 24968
rect 12259 24928 12268 24968
rect 12308 24928 12556 24968
rect 12596 24928 12605 24968
rect 16483 24928 16492 24968
rect 16532 24928 19852 24968
rect 19892 24928 19901 24968
rect 20039 24928 20048 24968
rect 20088 24928 20130 24968
rect 20170 24928 20212 24968
rect 20252 24928 20294 24968
rect 20334 24928 20376 24968
rect 20416 24928 20425 24968
rect 20812 24928 21504 24968
rect 0 24908 80 24928
rect 6403 24927 6461 24928
rect 16483 24927 16541 24928
rect 21424 24908 21504 24928
rect 16579 24884 16637 24885
rect 5443 24844 5452 24884
rect 5492 24844 16588 24884
rect 16628 24844 16637 24884
rect 18499 24844 18508 24884
rect 18548 24844 18836 24884
rect 16579 24843 16637 24844
rect 2851 24800 2909 24801
rect 7843 24800 7901 24801
rect 17347 24800 17405 24801
rect 2755 24760 2764 24800
rect 2804 24760 2860 24800
rect 2900 24760 2909 24800
rect 3139 24760 3148 24800
rect 3188 24760 3436 24800
rect 3476 24760 3485 24800
rect 7843 24760 7852 24800
rect 7892 24760 8236 24800
rect 8276 24760 8285 24800
rect 17251 24760 17260 24800
rect 17300 24760 17356 24800
rect 17396 24760 17405 24800
rect 2851 24759 2909 24760
rect 7843 24759 7901 24760
rect 17347 24759 17405 24760
rect 9667 24676 9676 24716
rect 9716 24676 9964 24716
rect 10004 24676 10013 24716
rect 2947 24632 3005 24633
rect 3523 24632 3581 24633
rect 10147 24632 10205 24633
rect 11011 24632 11069 24633
rect 18796 24632 18836 24844
rect 21424 24632 21504 24652
rect 1219 24592 1228 24632
rect 1268 24592 1516 24632
rect 1556 24592 1900 24632
rect 1940 24592 1949 24632
rect 2862 24592 2956 24632
rect 2996 24592 3532 24632
rect 3572 24592 3581 24632
rect 6691 24592 6700 24632
rect 6740 24592 7180 24632
rect 7220 24592 7229 24632
rect 7843 24592 7852 24632
rect 7892 24592 8236 24632
rect 8276 24592 10156 24632
rect 10196 24592 10205 24632
rect 10926 24592 11020 24632
rect 11060 24592 11069 24632
rect 15139 24592 15148 24632
rect 15188 24592 15197 24632
rect 17539 24592 17548 24632
rect 17588 24592 18412 24632
rect 18452 24592 18461 24632
rect 18787 24592 18796 24632
rect 18836 24592 18845 24632
rect 20515 24592 20524 24632
rect 20564 24592 21504 24632
rect 2947 24591 3005 24592
rect 3523 24591 3581 24592
rect 10147 24591 10205 24592
rect 11011 24591 11069 24592
rect 13795 24548 13853 24549
rect 15148 24548 15188 24592
rect 21424 24572 21504 24592
rect 10147 24508 10156 24548
rect 10196 24508 10540 24548
rect 10580 24508 10732 24548
rect 10772 24508 10781 24548
rect 13795 24508 13804 24548
rect 13844 24508 14764 24548
rect 14804 24508 17452 24548
rect 17492 24508 17501 24548
rect 18211 24508 18220 24548
rect 18260 24508 18988 24548
rect 19028 24508 19037 24548
rect 13795 24507 13853 24508
rect 0 24464 80 24484
rect 5635 24464 5693 24465
rect 17059 24464 17117 24465
rect 0 24424 2540 24464
rect 0 24404 80 24424
rect 2500 24296 2540 24424
rect 5635 24424 5644 24464
rect 5684 24424 10444 24464
rect 10484 24424 11308 24464
rect 11348 24424 11357 24464
rect 16291 24424 16300 24464
rect 16340 24424 16492 24464
rect 16532 24424 16541 24464
rect 16974 24424 17068 24464
rect 17108 24424 17356 24464
rect 17396 24424 17405 24464
rect 5635 24423 5693 24424
rect 17059 24423 17117 24424
rect 2659 24340 2668 24380
rect 2708 24340 2956 24380
rect 2996 24340 3005 24380
rect 7843 24340 7852 24380
rect 7892 24340 9580 24380
rect 9620 24340 9629 24380
rect 19171 24340 19180 24380
rect 19220 24340 20180 24380
rect 10627 24296 10685 24297
rect 20140 24296 20180 24340
rect 21424 24296 21504 24316
rect 2500 24256 10636 24296
rect 10676 24256 10685 24296
rect 14371 24256 14380 24296
rect 14420 24256 15820 24296
rect 15860 24256 17548 24296
rect 17588 24256 17597 24296
rect 20140 24256 21504 24296
rect 10627 24255 10685 24256
rect 21424 24236 21504 24256
rect 3679 24172 3688 24212
rect 3728 24172 3770 24212
rect 3810 24172 3852 24212
rect 3892 24172 3934 24212
rect 3974 24172 4016 24212
rect 4056 24172 4065 24212
rect 18799 24172 18808 24212
rect 18848 24172 18890 24212
rect 18930 24172 18972 24212
rect 19012 24172 19054 24212
rect 19094 24172 19136 24212
rect 19176 24172 19185 24212
rect 4867 24004 4876 24044
rect 4916 24004 5740 24044
rect 5780 24004 5789 24044
rect 15235 24004 15244 24044
rect 15284 24004 15628 24044
rect 15668 24004 15677 24044
rect 0 23961 80 23980
rect 0 23960 125 23961
rect 11299 23960 11357 23961
rect 17635 23960 17693 23961
rect 19843 23960 19901 23961
rect 21424 23960 21504 23980
rect 0 23920 76 23960
rect 116 23920 125 23960
rect 1603 23920 1612 23960
rect 1652 23920 2380 23960
rect 2420 23920 11308 23960
rect 11348 23920 11357 23960
rect 15523 23920 15532 23960
rect 15572 23920 17164 23960
rect 17204 23920 17213 23960
rect 17635 23920 17644 23960
rect 17684 23920 17778 23960
rect 18115 23920 18124 23960
rect 18164 23920 18316 23960
rect 18356 23920 18365 23960
rect 19843 23920 19852 23960
rect 19892 23920 21504 23960
rect 0 23919 125 23920
rect 11299 23919 11357 23920
rect 17635 23919 17693 23920
rect 19843 23919 19901 23920
rect 0 23900 80 23919
rect 21424 23900 21504 23920
rect 18307 23876 18365 23877
rect 1228 23836 1420 23876
rect 1460 23836 1469 23876
rect 2947 23836 2956 23876
rect 2996 23836 3340 23876
rect 3380 23836 3389 23876
rect 4003 23836 4012 23876
rect 4052 23836 8908 23876
rect 8948 23836 8957 23876
rect 10915 23836 10924 23876
rect 10964 23836 11308 23876
rect 11348 23836 11357 23876
rect 17923 23836 17932 23876
rect 17972 23836 18316 23876
rect 18356 23836 18365 23876
rect 1228 23792 1268 23836
rect 18307 23835 18365 23836
rect 5443 23792 5501 23793
rect 5731 23792 5789 23793
rect 8227 23792 8285 23793
rect 13891 23792 13949 23793
rect 1219 23752 1228 23792
rect 1268 23752 1277 23792
rect 2755 23752 2764 23792
rect 2804 23752 3052 23792
rect 3092 23752 3101 23792
rect 4483 23752 4492 23792
rect 4532 23752 5164 23792
rect 5204 23752 5452 23792
rect 5492 23752 5501 23792
rect 5635 23752 5644 23792
rect 5684 23752 5740 23792
rect 5780 23752 5836 23792
rect 5876 23752 5904 23792
rect 6499 23752 6508 23792
rect 6548 23752 6892 23792
rect 6932 23752 6941 23792
rect 8227 23752 8236 23792
rect 8276 23752 9004 23792
rect 9044 23752 9053 23792
rect 10723 23752 10732 23792
rect 10772 23752 10781 23792
rect 13806 23752 13900 23792
rect 13940 23752 13949 23792
rect 5443 23751 5501 23752
rect 5731 23751 5789 23752
rect 6892 23708 6932 23752
rect 8227 23751 8285 23752
rect 8611 23708 8669 23709
rect 10732 23708 10772 23752
rect 13891 23751 13949 23752
rect 17731 23792 17789 23793
rect 17731 23752 17740 23792
rect 17780 23752 18316 23792
rect 18356 23752 18365 23792
rect 18499 23752 18508 23792
rect 18548 23752 18892 23792
rect 18932 23752 18941 23792
rect 17731 23751 17789 23752
rect 4291 23668 4300 23708
rect 4340 23668 5068 23708
rect 5108 23668 6028 23708
rect 6068 23668 6077 23708
rect 6892 23668 8524 23708
rect 8564 23668 8620 23708
rect 8660 23668 8688 23708
rect 10435 23668 10444 23708
rect 10484 23668 10772 23708
rect 11011 23708 11069 23709
rect 11299 23708 11357 23709
rect 17923 23708 17981 23709
rect 18508 23708 18548 23752
rect 11011 23668 11020 23708
rect 11060 23668 11116 23708
rect 11156 23668 11165 23708
rect 11299 23668 11308 23708
rect 11348 23668 12076 23708
rect 12116 23668 12125 23708
rect 14851 23668 14860 23708
rect 14900 23668 17932 23708
rect 17972 23668 18548 23708
rect 19660 23668 20044 23708
rect 20084 23668 20093 23708
rect 8611 23667 8669 23668
rect 11011 23667 11069 23668
rect 11299 23667 11357 23668
rect 5539 23624 5597 23625
rect 8323 23624 8381 23625
rect 11788 23624 11828 23668
rect 17923 23667 17981 23668
rect 19660 23624 19700 23668
rect 21424 23624 21504 23644
rect 1795 23584 1804 23624
rect 1844 23584 2284 23624
rect 2324 23584 2333 23624
rect 3139 23584 3148 23624
rect 3188 23584 3532 23624
rect 3572 23584 3581 23624
rect 4099 23584 4108 23624
rect 4148 23584 4588 23624
rect 4628 23584 4972 23624
rect 5012 23584 5021 23624
rect 5443 23584 5452 23624
rect 5492 23584 5548 23624
rect 5588 23584 5597 23624
rect 7075 23584 7084 23624
rect 7124 23584 7564 23624
rect 7604 23584 8140 23624
rect 8180 23584 8189 23624
rect 8323 23584 8332 23624
rect 8372 23584 8466 23624
rect 8707 23584 8716 23624
rect 8756 23584 9292 23624
rect 9332 23584 9341 23624
rect 11779 23584 11788 23624
rect 11828 23584 11868 23624
rect 19651 23584 19660 23624
rect 19700 23584 19709 23624
rect 19939 23584 19948 23624
rect 19988 23584 21504 23624
rect 5539 23583 5597 23584
rect 8323 23583 8381 23584
rect 21424 23564 21504 23584
rect 4675 23540 4733 23541
rect 2467 23500 2476 23540
rect 2516 23500 4684 23540
rect 4724 23500 11360 23540
rect 16771 23500 16780 23540
rect 16820 23500 17780 23540
rect 4675 23499 4733 23500
rect 0 23456 80 23476
rect 5443 23456 5501 23457
rect 0 23416 3820 23456
rect 3860 23416 3869 23456
rect 4919 23416 4928 23456
rect 4968 23416 5010 23456
rect 5050 23416 5092 23456
rect 5132 23416 5174 23456
rect 5214 23416 5256 23456
rect 5296 23416 5305 23456
rect 5443 23416 5452 23456
rect 5492 23416 5644 23456
rect 5684 23416 5693 23456
rect 6019 23416 6028 23456
rect 6068 23416 6892 23456
rect 6932 23416 6941 23456
rect 9475 23416 9484 23456
rect 9524 23416 10732 23456
rect 10772 23416 10781 23456
rect 0 23396 80 23416
rect 5443 23415 5501 23416
rect 6787 23372 6845 23373
rect 3331 23332 3340 23372
rect 3380 23332 4396 23372
rect 4436 23332 6700 23372
rect 6740 23332 6796 23372
rect 6836 23332 6864 23372
rect 10339 23332 10348 23372
rect 10388 23332 10828 23372
rect 10868 23332 10877 23372
rect 6787 23331 6845 23332
rect 11320 23288 11360 23500
rect 17740 23456 17780 23500
rect 17731 23416 17740 23456
rect 17780 23416 17789 23456
rect 20039 23416 20048 23456
rect 20088 23416 20130 23456
rect 20170 23416 20212 23456
rect 20252 23416 20294 23456
rect 20334 23416 20376 23456
rect 20416 23416 20425 23456
rect 21424 23288 21504 23308
rect 3244 23248 4492 23288
rect 4532 23248 4541 23288
rect 4771 23248 4780 23288
rect 4820 23248 4829 23288
rect 6115 23248 6124 23288
rect 6164 23248 6173 23288
rect 8611 23248 8620 23288
rect 8660 23248 9772 23288
rect 9812 23248 9821 23288
rect 11320 23248 11404 23288
rect 11444 23248 11453 23288
rect 19267 23248 19276 23288
rect 19316 23248 19564 23288
rect 19604 23248 19613 23288
rect 20035 23248 20044 23288
rect 20084 23248 21504 23288
rect 3244 23204 3284 23248
rect 2851 23164 2860 23204
rect 2900 23164 3244 23204
rect 3284 23164 3293 23204
rect 3523 23164 3532 23204
rect 3572 23164 3724 23204
rect 3764 23164 3773 23204
rect 163 23120 221 23121
rect 4780 23120 4820 23248
rect 6124 23120 6164 23248
rect 21424 23228 21504 23248
rect 6307 23164 6316 23204
rect 6356 23164 6604 23204
rect 6644 23164 6988 23204
rect 7028 23164 7037 23204
rect 8323 23164 8332 23204
rect 8372 23164 9196 23204
rect 9236 23164 9245 23204
rect 10243 23164 10252 23204
rect 10292 23164 11980 23204
rect 12020 23164 13612 23204
rect 13652 23164 14764 23204
rect 14804 23164 14813 23204
rect 8707 23120 8765 23121
rect 163 23080 172 23120
rect 212 23080 1420 23120
rect 1460 23080 1469 23120
rect 4780 23080 5356 23120
rect 5396 23080 5405 23120
rect 5548 23080 7660 23120
rect 7700 23080 7709 23120
rect 8707 23080 8716 23120
rect 8756 23080 8812 23120
rect 8852 23080 8861 23120
rect 9283 23080 9292 23120
rect 9332 23080 9676 23120
rect 9716 23080 9725 23120
rect 11587 23080 11596 23120
rect 11636 23080 18316 23120
rect 18356 23080 18365 23120
rect 163 23079 221 23080
rect 4099 23036 4157 23037
rect 3715 22996 3724 23036
rect 3764 22996 4108 23036
rect 4148 22996 4157 23036
rect 4099 22995 4157 22996
rect 0 22952 80 22972
rect 5548 22952 5588 23080
rect 8707 23079 8765 23080
rect 6307 23036 6365 23037
rect 7075 23036 7133 23037
rect 5923 22996 5932 23036
rect 5972 22996 6316 23036
rect 6356 22996 7084 23036
rect 7124 22996 7133 23036
rect 8131 22996 8140 23036
rect 8180 22996 9484 23036
rect 9524 22996 9533 23036
rect 15523 22996 15532 23036
rect 15572 22996 19948 23036
rect 19988 22996 19997 23036
rect 6307 22995 6365 22996
rect 7075 22995 7133 22996
rect 21424 22952 21504 22972
rect 0 22912 3628 22952
rect 3668 22912 3677 22952
rect 4483 22912 4492 22952
rect 4532 22912 4780 22952
rect 4820 22912 5164 22952
rect 5204 22912 5213 22952
rect 5539 22912 5548 22952
rect 5588 22912 5597 22952
rect 6307 22912 6316 22952
rect 6356 22912 7468 22952
rect 7508 22912 7517 22952
rect 9571 22912 9580 22952
rect 9620 22912 10060 22952
rect 10100 22912 10109 22952
rect 19843 22912 19852 22952
rect 19892 22912 21504 22952
rect 0 22892 80 22912
rect 21424 22892 21504 22912
rect 7171 22868 7229 22869
rect 4099 22828 4108 22868
rect 4148 22828 6028 22868
rect 6068 22828 6077 22868
rect 7086 22828 7180 22868
rect 7220 22828 7229 22868
rect 15523 22828 15532 22868
rect 15572 22828 16396 22868
rect 16436 22828 16445 22868
rect 5539 22784 5597 22785
rect 6028 22784 6068 22828
rect 7171 22827 7229 22828
rect 8323 22784 8381 22785
rect 5539 22744 5548 22784
rect 5588 22744 5644 22784
rect 5684 22744 5693 22784
rect 6028 22744 8332 22784
rect 8372 22744 8524 22784
rect 8564 22744 8573 22784
rect 5539 22743 5597 22744
rect 8323 22743 8381 22744
rect 3679 22660 3688 22700
rect 3728 22660 3770 22700
rect 3810 22660 3852 22700
rect 3892 22660 3934 22700
rect 3974 22660 4016 22700
rect 4056 22660 4065 22700
rect 6883 22660 6892 22700
rect 6932 22660 7084 22700
rect 7124 22660 7133 22700
rect 7948 22660 8428 22700
rect 8468 22660 8477 22700
rect 12931 22660 12940 22700
rect 12980 22660 13228 22700
rect 13268 22660 13277 22700
rect 15811 22660 15820 22700
rect 15860 22660 16876 22700
rect 16916 22660 16925 22700
rect 18799 22660 18808 22700
rect 18848 22660 18890 22700
rect 18930 22660 18972 22700
rect 19012 22660 19054 22700
rect 19094 22660 19136 22700
rect 19176 22660 19185 22700
rect 7948 22616 7988 22660
rect 21424 22616 21504 22636
rect 5635 22576 5644 22616
rect 5684 22576 7756 22616
rect 7796 22576 7805 22616
rect 7939 22576 7948 22616
rect 7988 22576 7997 22616
rect 12451 22576 12460 22616
rect 12500 22576 19756 22616
rect 19796 22576 19805 22616
rect 21283 22576 21292 22616
rect 21332 22576 21504 22616
rect 21424 22556 21504 22576
rect 8419 22492 8428 22532
rect 8468 22492 10156 22532
rect 10196 22492 10205 22532
rect 12643 22492 12652 22532
rect 12692 22492 13132 22532
rect 13172 22492 13516 22532
rect 13556 22492 13565 22532
rect 16483 22492 16492 22532
rect 16532 22492 17452 22532
rect 17492 22492 18412 22532
rect 18452 22492 19564 22532
rect 19604 22492 19613 22532
rect 20131 22492 20140 22532
rect 20180 22492 20908 22532
rect 20948 22492 20957 22532
rect 0 22448 80 22468
rect 0 22408 8140 22448
rect 8180 22408 8189 22448
rect 19651 22408 19660 22448
rect 19700 22408 21332 22448
rect 0 22388 80 22408
rect 10915 22364 10973 22365
rect 13795 22364 13853 22365
rect 6211 22324 6220 22364
rect 6260 22324 7756 22364
rect 7796 22324 7805 22364
rect 9187 22324 9196 22364
rect 9236 22324 10540 22364
rect 10580 22324 10924 22364
rect 10964 22324 10973 22364
rect 12835 22324 12844 22364
rect 12884 22324 13804 22364
rect 13844 22324 13853 22364
rect 14659 22324 14668 22364
rect 14708 22324 19508 22364
rect 10915 22323 10973 22324
rect 13795 22323 13853 22324
rect 11011 22280 11069 22281
rect 2755 22240 2764 22280
rect 2804 22240 4300 22280
rect 4340 22240 4349 22280
rect 4963 22240 4972 22280
rect 5012 22240 5452 22280
rect 5492 22240 5501 22280
rect 7267 22240 7276 22280
rect 7316 22240 7660 22280
rect 7700 22240 7709 22280
rect 9283 22240 9292 22280
rect 9332 22240 9484 22280
rect 9524 22240 10252 22280
rect 10292 22240 10301 22280
rect 10435 22240 10444 22280
rect 10484 22240 11020 22280
rect 11060 22240 11069 22280
rect 11011 22239 11069 22240
rect 13027 22280 13085 22281
rect 14371 22280 14429 22281
rect 13027 22240 13036 22280
rect 13076 22240 13132 22280
rect 13172 22240 14380 22280
rect 14420 22240 14764 22280
rect 14804 22240 16108 22280
rect 16148 22240 16157 22280
rect 16963 22240 16972 22280
rect 17012 22240 17452 22280
rect 17492 22240 17501 22280
rect 13027 22239 13085 22240
rect 14371 22239 14429 22240
rect 6499 22196 6557 22197
rect 2851 22156 2860 22196
rect 2900 22156 5356 22196
rect 5396 22156 5405 22196
rect 6211 22156 6220 22196
rect 6260 22156 6508 22196
rect 6548 22156 6557 22196
rect 6499 22155 6557 22156
rect 7651 22196 7709 22197
rect 7651 22156 7660 22196
rect 7700 22156 11360 22196
rect 11683 22156 11692 22196
rect 11732 22156 19372 22196
rect 19412 22156 19421 22196
rect 7651 22155 7709 22156
rect 2851 22112 2909 22113
rect 11320 22112 11360 22156
rect 2832 22072 2860 22112
rect 2900 22072 2956 22112
rect 2996 22072 10004 22112
rect 11320 22072 12652 22112
rect 12692 22072 12701 22112
rect 12835 22072 12844 22112
rect 12884 22072 13324 22112
rect 13364 22072 13373 22112
rect 2851 22071 2909 22072
rect 7651 22028 7709 22029
rect 9676 22028 9716 22072
rect 1507 21988 1516 22028
rect 1556 21988 7660 22028
rect 7700 21988 7709 22028
rect 9667 21988 9676 22028
rect 9716 21988 9756 22028
rect 7651 21987 7709 21988
rect 0 21944 80 21964
rect 9964 21944 10004 22072
rect 19468 22028 19508 22324
rect 21292 22280 21332 22408
rect 21424 22280 21504 22300
rect 21292 22240 21504 22280
rect 21424 22220 21504 22240
rect 19555 22072 19564 22112
rect 19604 22072 21332 22112
rect 20611 22028 20669 22029
rect 19468 21988 20620 22028
rect 20660 21988 20669 22028
rect 20611 21987 20669 21988
rect 21292 21944 21332 22072
rect 21424 21944 21504 21964
rect 0 21904 1804 21944
rect 1844 21904 1853 21944
rect 4919 21904 4928 21944
rect 4968 21904 5010 21944
rect 5050 21904 5092 21944
rect 5132 21904 5174 21944
rect 5214 21904 5256 21944
rect 5296 21904 5305 21944
rect 8611 21904 8620 21944
rect 8660 21904 9196 21944
rect 9236 21904 9245 21944
rect 9379 21904 9388 21944
rect 9428 21904 9868 21944
rect 9908 21904 9917 21944
rect 9964 21904 12556 21944
rect 12596 21904 14860 21944
rect 14900 21904 14909 21944
rect 20039 21904 20048 21944
rect 20088 21904 20130 21944
rect 20170 21904 20212 21944
rect 20252 21904 20294 21944
rect 20334 21904 20376 21944
rect 20416 21904 20425 21944
rect 21292 21904 21504 21944
rect 0 21884 80 21904
rect 21424 21884 21504 21904
rect 6892 21820 9292 21860
rect 9332 21820 9341 21860
rect 11299 21820 11308 21860
rect 11348 21820 11500 21860
rect 11540 21820 11549 21860
rect 12451 21820 12460 21860
rect 12500 21820 12940 21860
rect 12980 21820 13324 21860
rect 13364 21820 13373 21860
rect 6892 21776 6932 21820
rect 5251 21736 5260 21776
rect 5300 21736 5740 21776
rect 5780 21736 6892 21776
rect 6932 21736 6941 21776
rect 7075 21736 7084 21776
rect 7124 21736 7468 21776
rect 7508 21736 7517 21776
rect 9187 21736 9196 21776
rect 9236 21736 18988 21776
rect 19028 21736 19037 21776
rect 2179 21652 2188 21692
rect 2228 21652 5644 21692
rect 5684 21652 5693 21692
rect 5740 21652 10348 21692
rect 10388 21652 13420 21692
rect 13460 21652 13469 21692
rect 18691 21652 18700 21692
rect 18740 21652 19468 21692
rect 19508 21652 19517 21692
rect 2659 21608 2717 21609
rect 5740 21608 5780 21652
rect 7939 21608 7997 21609
rect 13987 21608 14045 21609
rect 17443 21608 17501 21609
rect 21424 21608 21504 21628
rect 2659 21568 2668 21608
rect 2708 21568 3628 21608
rect 3668 21568 3677 21608
rect 4003 21568 4012 21608
rect 4052 21568 5684 21608
rect 5731 21568 5740 21608
rect 5780 21568 5789 21608
rect 7854 21568 7948 21608
rect 7988 21568 7997 21608
rect 8515 21568 8524 21608
rect 8564 21568 9772 21608
rect 9812 21568 9821 21608
rect 11107 21568 11116 21608
rect 11156 21568 11980 21608
rect 12020 21568 12029 21608
rect 13891 21568 13900 21608
rect 13940 21568 13996 21608
rect 14036 21568 14045 21608
rect 14371 21568 14380 21608
rect 14420 21568 14956 21608
rect 14996 21568 15005 21608
rect 17358 21568 17452 21608
rect 17492 21568 17501 21608
rect 20899 21568 20908 21608
rect 20948 21568 21504 21608
rect 2659 21567 2717 21568
rect 5644 21524 5684 21568
rect 7939 21567 7997 21568
rect 6691 21524 6749 21525
rect 8515 21524 8573 21525
rect 2500 21484 4684 21524
rect 4724 21484 4733 21524
rect 5644 21484 6700 21524
rect 6740 21484 8524 21524
rect 8564 21484 8573 21524
rect 9772 21524 9812 21568
rect 13987 21567 14045 21568
rect 17443 21567 17501 21568
rect 21424 21548 21504 21568
rect 9772 21484 11020 21524
rect 11060 21484 11069 21524
rect 14563 21484 14572 21524
rect 14612 21484 19372 21524
rect 19412 21484 19421 21524
rect 0 21440 80 21460
rect 2500 21440 2540 21484
rect 6691 21483 6749 21484
rect 8515 21483 8573 21484
rect 0 21400 2540 21440
rect 7555 21400 7564 21440
rect 7604 21400 8332 21440
rect 8372 21400 8381 21440
rect 16099 21400 16108 21440
rect 16148 21400 16300 21440
rect 16340 21400 16349 21440
rect 17539 21400 17548 21440
rect 17588 21400 18508 21440
rect 18548 21400 18796 21440
rect 18836 21400 18845 21440
rect 19555 21400 19564 21440
rect 19604 21400 21100 21440
rect 21140 21400 21149 21440
rect 0 21380 80 21400
rect 5443 21316 5452 21356
rect 5492 21316 6124 21356
rect 6164 21316 6173 21356
rect 8035 21316 8044 21356
rect 8084 21316 8620 21356
rect 8660 21316 8669 21356
rect 13891 21316 13900 21356
rect 13940 21316 14476 21356
rect 14516 21316 14525 21356
rect 19075 21316 19084 21356
rect 19124 21316 20180 21356
rect 20140 21272 20180 21316
rect 21424 21272 21504 21292
rect 15331 21232 15340 21272
rect 15380 21232 17548 21272
rect 17588 21232 17597 21272
rect 20140 21232 21504 21272
rect 21424 21212 21504 21232
rect 3679 21148 3688 21188
rect 3728 21148 3770 21188
rect 3810 21148 3852 21188
rect 3892 21148 3934 21188
rect 3974 21148 4016 21188
rect 4056 21148 4065 21188
rect 18799 21148 18808 21188
rect 18848 21148 18890 21188
rect 18930 21148 18972 21188
rect 19012 21148 19054 21188
rect 19094 21148 19136 21188
rect 19176 21148 19185 21188
rect 7747 21104 7805 21105
rect 1027 21064 1036 21104
rect 1076 21064 7756 21104
rect 7796 21064 7805 21104
rect 7747 21063 7805 21064
rect 17827 21020 17885 21021
rect 18115 21020 18173 21021
rect 4291 20980 4300 21020
rect 4340 20980 5548 21020
rect 5588 20980 5597 21020
rect 8995 20980 9004 21020
rect 9044 20980 9484 21020
rect 9524 20980 9533 21020
rect 17827 20980 17836 21020
rect 17876 20980 18124 21020
rect 18164 20980 18173 21020
rect 17827 20979 17885 20980
rect 18115 20979 18173 20980
rect 0 20936 80 20956
rect 163 20936 221 20937
rect 6307 20936 6365 20937
rect 21424 20936 21504 20956
rect 0 20896 172 20936
rect 212 20896 221 20936
rect 4099 20896 4108 20936
rect 4148 20896 6316 20936
rect 6356 20896 6365 20936
rect 10147 20896 10156 20936
rect 10196 20896 14284 20936
rect 14324 20896 14333 20936
rect 15907 20896 15916 20936
rect 15956 20896 18028 20936
rect 18068 20896 18412 20936
rect 18452 20896 18604 20936
rect 18644 20896 18653 20936
rect 19267 20896 19276 20936
rect 19316 20896 21504 20936
rect 0 20876 80 20896
rect 163 20895 221 20896
rect 6307 20895 6365 20896
rect 21424 20876 21504 20896
rect 4675 20852 4733 20853
rect 12451 20852 12509 20853
rect 4590 20812 4684 20852
rect 4724 20812 4733 20852
rect 6787 20812 6796 20852
rect 6836 20812 7180 20852
rect 7220 20812 7229 20852
rect 8131 20812 8140 20852
rect 8180 20812 12460 20852
rect 12500 20812 12509 20852
rect 4675 20811 4733 20812
rect 12451 20811 12509 20812
rect 12556 20812 13228 20852
rect 13268 20812 13708 20852
rect 13748 20812 13757 20852
rect 16099 20812 16108 20852
rect 16148 20812 16396 20852
rect 16436 20812 16445 20852
rect 16579 20812 16588 20852
rect 16628 20812 19852 20852
rect 19892 20812 19901 20852
rect 12556 20769 12596 20812
rect 4099 20768 4157 20769
rect 5923 20768 5981 20769
rect 4099 20728 4108 20768
rect 4148 20728 5068 20768
rect 5108 20728 5932 20768
rect 5972 20728 5981 20768
rect 4099 20727 4157 20728
rect 5923 20727 5981 20728
rect 6403 20768 6461 20769
rect 6691 20768 6749 20769
rect 6403 20728 6412 20768
rect 6452 20728 6700 20768
rect 6740 20728 6749 20768
rect 6403 20727 6461 20728
rect 6691 20727 6749 20728
rect 7843 20768 7901 20769
rect 12547 20768 12605 20769
rect 12739 20768 12797 20769
rect 14371 20768 14429 20769
rect 17635 20768 17693 20769
rect 7843 20728 7852 20768
rect 7892 20728 8044 20768
rect 8084 20728 8093 20768
rect 12547 20728 12556 20768
rect 12596 20728 12605 20768
rect 12654 20728 12748 20768
rect 12788 20728 12797 20768
rect 14286 20728 14380 20768
rect 14420 20728 14429 20768
rect 7843 20727 7901 20728
rect 12547 20727 12605 20728
rect 12739 20727 12797 20728
rect 14371 20727 14429 20728
rect 17620 20728 17644 20768
rect 17684 20728 17778 20768
rect 18019 20728 18028 20768
rect 18068 20728 18508 20768
rect 18548 20728 18557 20768
rect 17620 20727 17693 20728
rect 4291 20684 4349 20685
rect 14275 20684 14333 20685
rect 17155 20684 17213 20685
rect 3043 20644 3052 20684
rect 3092 20644 3148 20684
rect 3188 20644 3628 20684
rect 3668 20644 3677 20684
rect 4291 20644 4300 20684
rect 4340 20644 5932 20684
rect 5972 20644 6604 20684
rect 6644 20644 6653 20684
rect 8131 20644 8140 20684
rect 8180 20644 8716 20684
rect 8756 20644 8765 20684
rect 12451 20644 12460 20684
rect 12500 20644 12940 20684
rect 12980 20644 12989 20684
rect 14190 20644 14284 20684
rect 14324 20644 14333 20684
rect 17070 20644 17164 20684
rect 17204 20644 17213 20684
rect 4291 20643 4349 20644
rect 14275 20643 14333 20644
rect 17155 20643 17213 20644
rect 10243 20600 10301 20601
rect 17620 20600 17660 20727
rect 21424 20600 21504 20620
rect 10243 20560 10252 20600
rect 10292 20560 17660 20600
rect 19267 20560 19276 20600
rect 19316 20560 19852 20600
rect 19892 20560 19901 20600
rect 20803 20560 20812 20600
rect 20852 20560 21504 20600
rect 10243 20559 10301 20560
rect 21424 20540 21504 20560
rect 8035 20476 8044 20516
rect 8084 20476 8236 20516
rect 8276 20476 8285 20516
rect 15235 20476 15244 20516
rect 15284 20476 15820 20516
rect 15860 20476 15869 20516
rect 0 20432 80 20452
rect 547 20432 605 20433
rect 0 20392 556 20432
rect 596 20392 605 20432
rect 4919 20392 4928 20432
rect 4968 20392 5010 20432
rect 5050 20392 5092 20432
rect 5132 20392 5174 20432
rect 5214 20392 5256 20432
rect 5296 20392 5305 20432
rect 15427 20392 15436 20432
rect 15476 20392 17068 20432
rect 17108 20392 17117 20432
rect 20039 20392 20048 20432
rect 20088 20392 20130 20432
rect 20170 20392 20212 20432
rect 20252 20392 20294 20432
rect 20334 20392 20376 20432
rect 20416 20392 20425 20432
rect 0 20372 80 20392
rect 547 20391 605 20392
rect 4675 20308 4684 20348
rect 4724 20308 7372 20348
rect 7412 20308 7421 20348
rect 3427 20264 3485 20265
rect 16396 20264 16436 20392
rect 17635 20308 17644 20348
rect 17684 20308 18028 20348
rect 18068 20308 18077 20348
rect 19651 20308 19660 20348
rect 19700 20308 20180 20348
rect 20140 20264 20180 20308
rect 21424 20264 21504 20284
rect 3427 20224 3436 20264
rect 3476 20224 3532 20264
rect 3572 20224 3581 20264
rect 16300 20224 16436 20264
rect 17251 20224 17260 20264
rect 17300 20224 17548 20264
rect 17588 20224 17597 20264
rect 20140 20224 21504 20264
rect 3427 20223 3485 20224
rect 2947 20180 3005 20181
rect 2947 20140 2956 20180
rect 2996 20140 6740 20180
rect 7620 20140 7660 20180
rect 7700 20140 7709 20180
rect 12364 20140 12844 20180
rect 12884 20140 12893 20180
rect 15588 20140 15628 20180
rect 15668 20140 15677 20180
rect 2947 20139 3005 20140
rect 5347 20096 5405 20097
rect 3331 20056 3340 20096
rect 3380 20056 4396 20096
rect 4436 20056 4445 20096
rect 5262 20056 5356 20096
rect 5396 20056 5405 20096
rect 5347 20055 5405 20056
rect 6700 20012 6740 20140
rect 7660 20096 7700 20140
rect 8611 20096 8669 20097
rect 12364 20096 12404 20140
rect 15628 20096 15668 20140
rect 16300 20096 16340 20224
rect 21424 20204 21504 20224
rect 19651 20096 19709 20097
rect 6787 20056 6796 20096
rect 6836 20056 7700 20096
rect 8227 20056 8236 20096
rect 8276 20056 8620 20096
rect 8660 20056 8669 20096
rect 8899 20056 8908 20096
rect 8948 20056 10732 20096
rect 10772 20056 10781 20096
rect 12163 20056 12172 20096
rect 12212 20056 12404 20096
rect 12739 20056 12748 20096
rect 12788 20056 12940 20096
rect 12980 20056 12989 20096
rect 15628 20056 15764 20096
rect 15907 20056 15916 20096
rect 15956 20056 16340 20096
rect 17731 20056 17740 20096
rect 17780 20056 18220 20096
rect 18260 20056 18269 20096
rect 19459 20056 19468 20096
rect 19508 20056 19660 20096
rect 19700 20056 19709 20096
rect 8611 20055 8669 20056
rect 3235 19972 3244 20012
rect 3284 19972 4108 20012
rect 4148 19972 4588 20012
rect 4628 19972 4637 20012
rect 6700 19972 7756 20012
rect 7796 19972 9292 20012
rect 9332 19972 9341 20012
rect 12643 19972 12652 20012
rect 12692 19972 13420 20012
rect 13460 19972 13469 20012
rect 0 19928 80 19948
rect 11875 19928 11933 19929
rect 15724 19928 15764 20056
rect 19651 20055 19709 20056
rect 16579 20012 16637 20013
rect 15811 19972 15820 20012
rect 15860 19972 16588 20012
rect 16628 19972 16637 20012
rect 16579 19971 16637 19972
rect 21424 19928 21504 19948
rect 0 19888 2540 19928
rect 2947 19888 2956 19928
rect 2996 19888 3916 19928
rect 3956 19888 4492 19928
rect 4532 19888 5260 19928
rect 5300 19888 5309 19928
rect 8419 19888 8428 19928
rect 8468 19888 8716 19928
rect 8756 19888 8765 19928
rect 10435 19888 10444 19928
rect 10484 19888 11692 19928
rect 11732 19888 11741 19928
rect 11875 19888 11884 19928
rect 11924 19888 14956 19928
rect 14996 19888 15005 19928
rect 15724 19888 16204 19928
rect 16244 19888 16253 19928
rect 20035 19888 20044 19928
rect 20084 19888 21504 19928
rect 0 19868 80 19888
rect 2500 19844 2540 19888
rect 11875 19887 11933 19888
rect 21424 19868 21504 19888
rect 3139 19844 3197 19845
rect 7171 19844 7229 19845
rect 13987 19844 14045 19845
rect 2500 19804 3148 19844
rect 3188 19804 3197 19844
rect 3811 19804 3820 19844
rect 3860 19804 7180 19844
rect 7220 19804 7229 19844
rect 3139 19803 3197 19804
rect 7171 19803 7229 19804
rect 7276 19804 9196 19844
rect 9236 19804 12364 19844
rect 12404 19804 12413 19844
rect 13987 19804 13996 19844
rect 14036 19804 14996 19844
rect 15043 19804 15052 19844
rect 15092 19804 15724 19844
rect 15764 19804 15773 19844
rect 3427 19760 3485 19761
rect 7276 19760 7316 19804
rect 13987 19803 14045 19804
rect 14956 19760 14996 19804
rect 3235 19720 3244 19760
rect 3284 19720 3436 19760
rect 3476 19720 6988 19760
rect 7028 19720 7037 19760
rect 7267 19720 7276 19760
rect 7316 19720 7325 19760
rect 10147 19720 10156 19760
rect 10196 19720 14476 19760
rect 14516 19720 14525 19760
rect 14956 19720 16780 19760
rect 16820 19720 17068 19760
rect 17108 19720 17117 19760
rect 3427 19719 3485 19720
rect 13411 19676 13469 19677
rect 3679 19636 3688 19676
rect 3728 19636 3770 19676
rect 3810 19636 3852 19676
rect 3892 19636 3934 19676
rect 3974 19636 4016 19676
rect 4056 19636 4065 19676
rect 5836 19636 8908 19676
rect 8948 19636 8957 19676
rect 10435 19636 10444 19676
rect 10484 19636 11020 19676
rect 11060 19636 11069 19676
rect 13411 19636 13420 19676
rect 13460 19636 15244 19676
rect 15284 19636 15532 19676
rect 15572 19636 15581 19676
rect 18799 19636 18808 19676
rect 18848 19636 18890 19676
rect 18930 19636 18972 19676
rect 19012 19636 19054 19676
rect 19094 19636 19136 19676
rect 19176 19636 19185 19676
rect 5836 19592 5876 19636
rect 13411 19635 13469 19636
rect 2083 19552 2092 19592
rect 2132 19552 3340 19592
rect 3380 19552 5876 19592
rect 7171 19592 7229 19593
rect 21424 19592 21504 19612
rect 7171 19552 7180 19592
rect 7220 19552 16588 19592
rect 16628 19552 16637 19592
rect 19555 19552 19564 19592
rect 19604 19552 21504 19592
rect 7171 19551 7229 19552
rect 21424 19532 21504 19552
rect 2659 19508 2717 19509
rect 2574 19468 2668 19508
rect 2708 19468 2717 19508
rect 6979 19468 6988 19508
rect 7028 19468 10444 19508
rect 10484 19468 10493 19508
rect 11683 19468 11692 19508
rect 11732 19468 18988 19508
rect 19028 19468 19037 19508
rect 2659 19467 2717 19468
rect 0 19424 80 19444
rect 13411 19424 13469 19425
rect 0 19384 556 19424
rect 596 19384 605 19424
rect 1315 19384 1324 19424
rect 1364 19384 1900 19424
rect 1940 19384 13420 19424
rect 13460 19384 13469 19424
rect 0 19364 80 19384
rect 13411 19383 13469 19384
rect 13891 19424 13949 19425
rect 14275 19424 14333 19425
rect 13891 19384 13900 19424
rect 13940 19384 14284 19424
rect 14324 19384 17548 19424
rect 17588 19384 17597 19424
rect 13891 19383 13949 19384
rect 14275 19383 14333 19384
rect 3811 19300 3820 19340
rect 3860 19300 4396 19340
rect 4436 19300 4445 19340
rect 7843 19300 7852 19340
rect 7892 19300 19372 19340
rect 19412 19300 19421 19340
rect 12835 19256 12893 19257
rect 17923 19256 17981 19257
rect 21424 19256 21504 19276
rect 2083 19216 2092 19256
rect 2132 19216 2476 19256
rect 2516 19216 2764 19256
rect 2804 19216 2813 19256
rect 3907 19216 3916 19256
rect 3956 19216 4492 19256
rect 4532 19216 4541 19256
rect 5347 19216 5356 19256
rect 5396 19216 6412 19256
rect 6452 19216 8620 19256
rect 8660 19216 9484 19256
rect 9524 19216 10156 19256
rect 10196 19216 10205 19256
rect 11107 19216 11116 19256
rect 11156 19216 12844 19256
rect 12884 19216 12893 19256
rect 12835 19215 12893 19216
rect 12940 19247 13172 19256
rect 12940 19216 13132 19247
rect 12940 19172 12980 19216
rect 13123 19207 13132 19216
rect 13172 19207 13181 19247
rect 13315 19216 13324 19256
rect 13364 19216 13373 19256
rect 13507 19216 13516 19256
rect 13556 19216 13900 19256
rect 13940 19216 13949 19256
rect 14371 19216 14380 19256
rect 14420 19216 14956 19256
rect 14996 19216 15005 19256
rect 16483 19216 16492 19256
rect 16532 19216 17164 19256
rect 17204 19216 17213 19256
rect 17923 19216 17932 19256
rect 17972 19216 18028 19256
rect 18068 19216 18796 19256
rect 18836 19216 18845 19256
rect 20611 19216 20620 19256
rect 20660 19216 21504 19256
rect 12451 19132 12460 19172
rect 12500 19132 12980 19172
rect 7843 19088 7901 19089
rect 8803 19088 8861 19089
rect 13324 19088 13364 19216
rect 17923 19215 17981 19216
rect 21424 19196 21504 19216
rect 13795 19132 13804 19172
rect 13844 19132 14668 19172
rect 14708 19132 15572 19172
rect 18691 19132 18700 19172
rect 18740 19132 19756 19172
rect 19796 19132 19805 19172
rect 7843 19048 7852 19088
rect 7892 19048 8524 19088
rect 8564 19048 8573 19088
rect 8803 19048 8812 19088
rect 8852 19048 12940 19088
rect 12980 19048 12989 19088
rect 13219 19048 13228 19088
rect 13268 19048 13364 19088
rect 14083 19048 14092 19088
rect 14132 19048 15436 19088
rect 15476 19048 15485 19088
rect 7843 19047 7901 19048
rect 8803 19047 8861 19048
rect 15532 19004 15572 19132
rect 16579 19048 16588 19088
rect 16628 19048 17068 19088
rect 17108 19048 17117 19088
rect 19939 19048 19948 19088
rect 19988 19048 21332 19088
rect 13699 18964 13708 19004
rect 13748 18964 14668 19004
rect 14708 18964 14717 19004
rect 15139 18964 15148 19004
rect 15188 18964 15572 19004
rect 15715 19004 15773 19005
rect 15715 18964 15724 19004
rect 15764 18964 17740 19004
rect 17780 18964 17789 19004
rect 15715 18963 15773 18964
rect 0 18920 80 18940
rect 1219 18920 1277 18921
rect 6211 18920 6269 18921
rect 21292 18920 21332 19048
rect 21424 18920 21504 18940
rect 0 18880 1228 18920
rect 1268 18880 1277 18920
rect 0 18860 80 18880
rect 1219 18879 1277 18880
rect 2284 18880 3244 18920
rect 3284 18880 3293 18920
rect 4919 18880 4928 18920
rect 4968 18880 5010 18920
rect 5050 18880 5092 18920
rect 5132 18880 5174 18920
rect 5214 18880 5256 18920
rect 5296 18880 5305 18920
rect 6211 18880 6220 18920
rect 6260 18880 8812 18920
rect 8852 18880 9100 18920
rect 9140 18880 9149 18920
rect 13027 18880 13036 18920
rect 13076 18880 15820 18920
rect 15860 18880 15869 18920
rect 16291 18880 16300 18920
rect 16340 18880 17452 18920
rect 17492 18880 18316 18920
rect 18356 18880 18365 18920
rect 20039 18880 20048 18920
rect 20088 18880 20130 18920
rect 20170 18880 20212 18920
rect 20252 18880 20294 18920
rect 20334 18880 20376 18920
rect 20416 18880 20425 18920
rect 21292 18880 21504 18920
rect 1891 18712 1900 18752
rect 1940 18712 2188 18752
rect 2228 18712 2237 18752
rect 2284 18668 2324 18880
rect 6211 18879 6269 18880
rect 21424 18860 21504 18880
rect 19267 18836 19325 18837
rect 4099 18796 4108 18836
rect 4148 18796 10828 18836
rect 10868 18796 11212 18836
rect 11252 18796 11261 18836
rect 13891 18796 13900 18836
rect 13940 18796 14572 18836
rect 14612 18796 14621 18836
rect 15043 18796 15052 18836
rect 15092 18796 16012 18836
rect 16052 18796 16061 18836
rect 19267 18796 19276 18836
rect 19316 18796 21292 18836
rect 21332 18796 21341 18836
rect 4195 18752 4253 18753
rect 5164 18752 5204 18796
rect 19267 18795 19325 18796
rect 11971 18752 12029 18753
rect 17059 18752 17117 18753
rect 4110 18712 4204 18752
rect 4244 18712 4253 18752
rect 5155 18712 5164 18752
rect 5204 18712 5213 18752
rect 11971 18712 11980 18752
rect 12020 18712 13324 18752
rect 13364 18712 13373 18752
rect 14755 18712 14764 18752
rect 14804 18712 15628 18752
rect 15668 18712 15677 18752
rect 15811 18712 15820 18752
rect 15860 18712 17068 18752
rect 17108 18712 17117 18752
rect 4195 18711 4253 18712
rect 11971 18711 12029 18712
rect 17059 18711 17117 18712
rect 2188 18628 2324 18668
rect 3235 18668 3293 18669
rect 17155 18668 17213 18669
rect 3235 18628 3244 18668
rect 3284 18628 3340 18668
rect 3380 18628 3389 18668
rect 11299 18628 11308 18668
rect 11348 18628 11360 18668
rect 13507 18628 13516 18668
rect 13556 18628 17164 18668
rect 17204 18628 17213 18668
rect 17443 18628 17452 18668
rect 17492 18628 17740 18668
rect 17780 18628 17789 18668
rect 2188 18584 2228 18628
rect 3235 18627 3293 18628
rect 11320 18584 11360 18628
rect 17155 18627 17213 18628
rect 17539 18584 17597 18585
rect 18595 18584 18653 18585
rect 21424 18584 21504 18604
rect 2179 18544 2188 18584
rect 2228 18544 2237 18584
rect 2563 18544 2572 18584
rect 2612 18544 3244 18584
rect 3284 18544 3293 18584
rect 8227 18544 8236 18584
rect 8276 18544 8428 18584
rect 8468 18544 8477 18584
rect 9283 18544 9292 18584
rect 9332 18544 9676 18584
rect 9716 18544 9725 18584
rect 11320 18544 11596 18584
rect 11636 18544 11645 18584
rect 11779 18544 11788 18584
rect 11828 18544 16012 18584
rect 16052 18544 16061 18584
rect 17539 18544 17548 18584
rect 17588 18544 17836 18584
rect 17876 18544 17885 18584
rect 18595 18544 18604 18584
rect 18644 18544 18796 18584
rect 18836 18544 18845 18584
rect 19843 18544 19852 18584
rect 19892 18544 21504 18584
rect 17539 18543 17597 18544
rect 18595 18543 18653 18544
rect 21424 18524 21504 18544
rect 18307 18500 18365 18501
rect 259 18460 268 18500
rect 308 18460 5548 18500
rect 5588 18460 5597 18500
rect 7747 18460 7756 18500
rect 7796 18460 14860 18500
rect 14900 18460 14909 18500
rect 18222 18460 18316 18500
rect 18356 18460 18365 18500
rect 18307 18459 18365 18460
rect 0 18416 80 18436
rect 14755 18416 14813 18417
rect 0 18376 12460 18416
rect 12500 18376 12509 18416
rect 14755 18376 14764 18416
rect 14804 18376 16972 18416
rect 17012 18376 17021 18416
rect 0 18356 80 18376
rect 14755 18375 14813 18376
rect 6019 18332 6077 18333
rect 17347 18332 17405 18333
rect 643 18292 652 18332
rect 692 18292 6028 18332
rect 6068 18292 6077 18332
rect 9667 18292 9676 18332
rect 9716 18292 10732 18332
rect 10772 18292 10781 18332
rect 13987 18292 13996 18332
rect 14036 18292 14380 18332
rect 14420 18292 14429 18332
rect 14947 18292 14956 18332
rect 14996 18292 15724 18332
rect 15764 18292 15773 18332
rect 17251 18292 17260 18332
rect 17300 18292 17356 18332
rect 17396 18292 17405 18332
rect 19171 18292 19180 18332
rect 19220 18292 20180 18332
rect 6019 18291 6077 18292
rect 17347 18291 17405 18292
rect 16099 18248 16157 18249
rect 3139 18208 3148 18248
rect 3188 18208 3532 18248
rect 3572 18208 5932 18248
rect 5972 18208 5981 18248
rect 7459 18208 7468 18248
rect 7508 18208 9868 18248
rect 9908 18208 9917 18248
rect 11779 18208 11788 18248
rect 11828 18208 15628 18248
rect 15668 18208 15677 18248
rect 16003 18208 16012 18248
rect 16052 18208 16108 18248
rect 16148 18208 16157 18248
rect 20140 18248 20180 18292
rect 21424 18248 21504 18268
rect 20140 18208 21504 18248
rect 16099 18207 16157 18208
rect 21424 18188 21504 18208
rect 9187 18164 9245 18165
rect 3679 18124 3688 18164
rect 3728 18124 3770 18164
rect 3810 18124 3852 18164
rect 3892 18124 3934 18164
rect 3974 18124 4016 18164
rect 4056 18124 4065 18164
rect 9102 18124 9196 18164
rect 9236 18124 9245 18164
rect 11203 18124 11212 18164
rect 11252 18124 18316 18164
rect 18356 18124 18365 18164
rect 18799 18124 18808 18164
rect 18848 18124 18890 18164
rect 18930 18124 18972 18164
rect 19012 18124 19054 18164
rect 19094 18124 19136 18164
rect 19176 18124 19185 18164
rect 9187 18123 9245 18124
rect 7171 18040 7180 18080
rect 7220 18040 20044 18080
rect 20084 18040 20093 18080
rect 13795 17996 13853 17997
rect 18595 17996 18653 17997
rect 8227 17956 8236 17996
rect 8276 17956 9580 17996
rect 9620 17956 9629 17996
rect 9676 17956 13804 17996
rect 13844 17956 14572 17996
rect 14612 17956 14621 17996
rect 15235 17956 15244 17996
rect 15284 17956 16012 17996
rect 16052 17956 16061 17996
rect 16195 17956 16204 17996
rect 16244 17956 16684 17996
rect 16724 17956 16733 17996
rect 18595 17956 18604 17996
rect 18644 17956 18796 17996
rect 18836 17956 18845 17996
rect 0 17912 80 17932
rect 8227 17912 8285 17913
rect 9676 17912 9716 17956
rect 13795 17955 13853 17956
rect 18595 17955 18653 17956
rect 19267 17912 19325 17913
rect 21424 17912 21504 17932
rect 0 17872 76 17912
rect 116 17872 125 17912
rect 5251 17872 5260 17912
rect 5300 17872 6028 17912
rect 6068 17872 8236 17912
rect 8276 17872 8285 17912
rect 8707 17872 8716 17912
rect 8756 17872 9196 17912
rect 9236 17872 9245 17912
rect 9667 17872 9676 17912
rect 9716 17872 9725 17912
rect 15244 17872 16780 17912
rect 16820 17872 16829 17912
rect 18499 17872 18508 17912
rect 18548 17872 18836 17912
rect 19075 17872 19084 17912
rect 19124 17872 19276 17912
rect 19316 17872 19325 17912
rect 20227 17872 20236 17912
rect 20276 17872 21504 17912
rect 0 17852 80 17872
rect 8227 17871 8285 17872
rect 4099 17828 4157 17829
rect 8131 17828 8189 17829
rect 14755 17828 14813 17829
rect 15244 17828 15284 17872
rect 18796 17828 18836 17872
rect 19267 17871 19325 17872
rect 21424 17852 21504 17872
rect 19651 17828 19709 17829
rect 4099 17788 4108 17828
rect 4148 17788 7276 17828
rect 7316 17788 8140 17828
rect 8180 17788 8189 17828
rect 4099 17787 4157 17788
rect 8131 17787 8189 17788
rect 9292 17788 10388 17828
rect 10435 17788 10444 17828
rect 10484 17788 10924 17828
rect 10964 17788 10973 17828
rect 14659 17788 14668 17828
rect 14708 17788 14764 17828
rect 14804 17788 14813 17828
rect 15235 17788 15244 17828
rect 15284 17788 15293 17828
rect 15715 17788 15724 17828
rect 15764 17788 16204 17828
rect 16244 17788 16253 17828
rect 18211 17788 18220 17828
rect 18260 17788 18740 17828
rect 18796 17788 19660 17828
rect 19700 17788 19709 17828
rect 9292 17744 9332 17788
rect 10243 17744 10301 17745
rect 6499 17704 6508 17744
rect 6548 17704 6988 17744
rect 7028 17704 7037 17744
rect 9283 17704 9292 17744
rect 9332 17704 9341 17744
rect 10158 17704 10252 17744
rect 10292 17704 10301 17744
rect 10348 17744 10388 17788
rect 14755 17787 14813 17788
rect 12259 17744 12317 17745
rect 16771 17744 16829 17745
rect 10348 17704 12268 17744
rect 12308 17704 12317 17744
rect 13795 17704 13804 17744
rect 13844 17704 16012 17744
rect 16052 17704 16061 17744
rect 16771 17704 16780 17744
rect 16820 17704 17164 17744
rect 17204 17704 18508 17744
rect 18548 17704 18557 17744
rect 10243 17703 10301 17704
rect 12259 17703 12317 17704
rect 16771 17703 16829 17704
rect 7939 17660 7997 17661
rect 451 17620 460 17660
rect 500 17620 7756 17660
rect 7796 17620 7805 17660
rect 7939 17620 7948 17660
rect 7988 17620 8082 17660
rect 9091 17620 9100 17660
rect 9140 17620 9772 17660
rect 9812 17620 9821 17660
rect 7939 17619 7997 17620
rect 18700 17576 18740 17788
rect 19651 17787 19709 17788
rect 19459 17704 19468 17744
rect 19508 17704 20524 17744
rect 20564 17704 20573 17744
rect 19651 17660 19709 17661
rect 19566 17620 19660 17660
rect 19700 17620 19709 17660
rect 19939 17620 19948 17660
rect 19988 17620 20180 17660
rect 19651 17619 19709 17620
rect 19459 17576 19517 17577
rect 2275 17536 2284 17576
rect 2324 17536 8044 17576
rect 8084 17536 8093 17576
rect 10915 17536 10924 17576
rect 10964 17536 18028 17576
rect 18068 17536 18077 17576
rect 18700 17536 19468 17576
rect 19508 17536 19517 17576
rect 20140 17576 20180 17620
rect 21424 17576 21504 17596
rect 20140 17536 21504 17576
rect 19459 17535 19517 17536
rect 21424 17516 21504 17536
rect 14659 17492 14717 17493
rect 1411 17452 1420 17492
rect 1460 17452 2572 17492
rect 2612 17452 9484 17492
rect 9524 17452 9533 17492
rect 9955 17452 9964 17492
rect 10004 17452 14668 17492
rect 14708 17452 15052 17492
rect 15092 17452 15101 17492
rect 14659 17451 14717 17452
rect 0 17408 80 17428
rect 4195 17408 4253 17409
rect 0 17368 2860 17408
rect 2900 17368 2909 17408
rect 3043 17368 3052 17408
rect 3092 17368 4204 17408
rect 4244 17368 4253 17408
rect 4919 17368 4928 17408
rect 4968 17368 5010 17408
rect 5050 17368 5092 17408
rect 5132 17368 5174 17408
rect 5214 17368 5256 17408
rect 5296 17368 5305 17408
rect 8899 17368 8908 17408
rect 8948 17368 19948 17408
rect 19988 17368 19997 17408
rect 20039 17368 20048 17408
rect 20088 17368 20130 17408
rect 20170 17368 20212 17408
rect 20252 17368 20294 17408
rect 20334 17368 20376 17408
rect 20416 17368 20425 17408
rect 0 17348 80 17368
rect 4195 17367 4253 17368
rect 17827 17324 17885 17325
rect 14947 17284 14956 17324
rect 14996 17284 15148 17324
rect 15188 17284 15197 17324
rect 17635 17284 17644 17324
rect 17684 17284 17836 17324
rect 17876 17284 17885 17324
rect 17827 17283 17885 17284
rect 21424 17240 21504 17260
rect 3043 17200 3052 17240
rect 3092 17200 3340 17240
rect 3380 17200 3389 17240
rect 11395 17200 11404 17240
rect 11444 17200 11692 17240
rect 11732 17200 11741 17240
rect 13900 17200 14764 17240
rect 14804 17200 14813 17240
rect 19267 17200 19276 17240
rect 19316 17200 19852 17240
rect 19892 17200 19901 17240
rect 21091 17200 21100 17240
rect 21140 17200 21504 17240
rect 13900 17156 13940 17200
rect 21424 17180 21504 17200
rect 14563 17156 14621 17157
rect 18403 17156 18461 17157
rect 1315 17116 1324 17156
rect 1364 17116 2284 17156
rect 2324 17116 2333 17156
rect 3523 17116 3532 17156
rect 3572 17116 8524 17156
rect 8564 17116 8573 17156
rect 9091 17116 9100 17156
rect 9140 17116 11212 17156
rect 11252 17116 13132 17156
rect 13172 17116 13900 17156
rect 13940 17116 13949 17156
rect 14563 17116 14572 17156
rect 14612 17116 15148 17156
rect 15188 17116 15197 17156
rect 18307 17116 18316 17156
rect 18356 17116 18412 17156
rect 18452 17116 18461 17156
rect 14563 17115 14621 17116
rect 18403 17115 18461 17116
rect 2467 17032 2476 17072
rect 2516 17032 3820 17072
rect 3860 17032 4780 17072
rect 4820 17032 4829 17072
rect 8035 17032 8044 17072
rect 8084 17032 9196 17072
rect 9236 17032 9964 17072
rect 10004 17032 10013 17072
rect 13699 17032 13708 17072
rect 13748 17032 14188 17072
rect 14228 17032 15340 17072
rect 15380 17032 15389 17072
rect 16675 17032 16684 17072
rect 16724 17032 17164 17072
rect 17204 17032 17213 17072
rect 18211 16988 18269 16989
rect 2851 16948 2860 16988
rect 2900 16948 3340 16988
rect 3380 16948 3389 16988
rect 6787 16948 6796 16988
rect 6836 16948 7372 16988
rect 7412 16948 7421 16988
rect 18211 16948 18220 16988
rect 18260 16948 18316 16988
rect 18356 16948 18365 16988
rect 18211 16947 18269 16948
rect 0 16904 80 16924
rect 11779 16904 11837 16905
rect 21424 16904 21504 16924
rect 0 16864 11788 16904
rect 11828 16864 11837 16904
rect 20227 16864 20236 16904
rect 20276 16864 21504 16904
rect 0 16844 80 16864
rect 11779 16863 11837 16864
rect 21424 16844 21504 16864
rect 18595 16820 18653 16821
rect 3043 16780 3052 16820
rect 3092 16780 4780 16820
rect 4820 16780 4829 16820
rect 8515 16780 8524 16820
rect 8564 16780 13708 16820
rect 13748 16780 13757 16820
rect 18595 16780 18604 16820
rect 18644 16780 18796 16820
rect 18836 16780 18845 16820
rect 18595 16779 18653 16780
rect 9475 16696 9484 16736
rect 9524 16696 11980 16736
rect 12020 16696 15916 16736
rect 15956 16696 15965 16736
rect 10915 16652 10973 16653
rect 16579 16652 16637 16653
rect 18403 16652 18461 16653
rect 1699 16612 1708 16652
rect 1748 16612 3532 16652
rect 3572 16612 3581 16652
rect 3679 16612 3688 16652
rect 3728 16612 3770 16652
rect 3810 16612 3852 16652
rect 3892 16612 3934 16652
rect 3974 16612 4016 16652
rect 4056 16612 4065 16652
rect 9859 16612 9868 16652
rect 9908 16612 10924 16652
rect 10964 16612 10973 16652
rect 12259 16612 12268 16652
rect 12308 16612 14284 16652
rect 14324 16612 14668 16652
rect 14708 16612 14717 16652
rect 16483 16612 16492 16652
rect 16532 16612 16588 16652
rect 16628 16612 16637 16652
rect 16867 16612 16876 16652
rect 16916 16612 17548 16652
rect 17588 16612 17597 16652
rect 18211 16612 18220 16652
rect 18260 16612 18412 16652
rect 18452 16612 18461 16652
rect 18799 16612 18808 16652
rect 18848 16612 18890 16652
rect 18930 16612 18972 16652
rect 19012 16612 19054 16652
rect 19094 16612 19136 16652
rect 19176 16612 19185 16652
rect 10915 16611 10973 16612
rect 16579 16611 16637 16612
rect 18403 16611 18461 16612
rect 19267 16568 19325 16569
rect 21424 16568 21504 16588
rect 172 16528 19276 16568
rect 19316 16528 19325 16568
rect 20899 16528 20908 16568
rect 20948 16528 21504 16568
rect 0 16400 80 16420
rect 172 16400 212 16528
rect 19267 16527 19325 16528
rect 21424 16508 21504 16528
rect 4195 16484 4253 16485
rect 4675 16484 4733 16485
rect 3331 16444 3340 16484
rect 3380 16444 3628 16484
rect 3668 16444 3677 16484
rect 3811 16444 3820 16484
rect 3860 16444 4204 16484
rect 4244 16444 4684 16484
rect 4724 16444 4733 16484
rect 15619 16444 15628 16484
rect 15668 16444 17740 16484
rect 17780 16444 17789 16484
rect 4195 16443 4253 16444
rect 4675 16443 4733 16444
rect 0 16360 212 16400
rect 931 16400 989 16401
rect 3427 16400 3485 16401
rect 13219 16400 13277 16401
rect 17059 16400 17117 16401
rect 931 16360 940 16400
rect 980 16360 1132 16400
rect 1172 16360 1181 16400
rect 3342 16360 3436 16400
rect 3476 16360 3485 16400
rect 4483 16360 4492 16400
rect 4532 16360 5260 16400
rect 5300 16360 6700 16400
rect 6740 16360 7377 16400
rect 7417 16360 7426 16400
rect 8035 16360 8044 16400
rect 8084 16360 9868 16400
rect 9908 16360 11020 16400
rect 11060 16360 11069 16400
rect 13219 16360 13228 16400
rect 13268 16360 16300 16400
rect 16340 16360 16492 16400
rect 16532 16360 16541 16400
rect 16588 16360 16684 16400
rect 16724 16360 16733 16400
rect 16974 16360 17068 16400
rect 17108 16360 17117 16400
rect 0 16340 80 16360
rect 931 16359 989 16360
rect 3427 16359 3485 16360
rect 13219 16359 13277 16360
rect 9475 16316 9533 16317
rect 3907 16276 3916 16316
rect 3956 16276 5452 16316
rect 5492 16276 8524 16316
rect 8564 16276 8573 16316
rect 9390 16276 9484 16316
rect 9524 16276 9533 16316
rect 12163 16276 12172 16316
rect 12212 16276 14956 16316
rect 14996 16276 16204 16316
rect 16244 16276 16253 16316
rect 9475 16275 9533 16276
rect 4195 16232 4253 16233
rect 2755 16192 2764 16232
rect 2804 16192 3340 16232
rect 3380 16192 3389 16232
rect 4195 16192 4204 16232
rect 4244 16192 5164 16232
rect 5204 16192 5213 16232
rect 5539 16192 5548 16232
rect 5588 16192 7180 16232
rect 7220 16192 7229 16232
rect 7843 16192 7852 16232
rect 7892 16192 13036 16232
rect 13076 16192 13085 16232
rect 15523 16192 15532 16232
rect 15572 16192 15916 16232
rect 15956 16192 16492 16232
rect 16532 16192 16541 16232
rect 4195 16191 4253 16192
rect 5059 16148 5117 16149
rect 4974 16108 5068 16148
rect 5108 16108 5117 16148
rect 5059 16107 5117 16108
rect 5731 16148 5789 16149
rect 5731 16108 5740 16148
rect 5780 16108 6220 16148
rect 6260 16108 6269 16148
rect 5731 16107 5789 16108
rect 16588 16064 16628 16360
rect 17059 16359 17117 16360
rect 17347 16276 17356 16316
rect 17396 16276 17740 16316
rect 17780 16276 17789 16316
rect 21424 16232 21504 16252
rect 16675 16192 16684 16232
rect 16724 16192 16876 16232
rect 16916 16192 17836 16232
rect 17876 16192 17885 16232
rect 18307 16192 18316 16232
rect 18356 16192 21504 16232
rect 21424 16172 21504 16192
rect 19651 16108 19660 16148
rect 19700 16108 20180 16148
rect 20140 16064 20180 16108
rect 2851 16024 2860 16064
rect 2900 16024 3052 16064
rect 3092 16024 3101 16064
rect 4387 16024 4396 16064
rect 4436 16024 6700 16064
rect 6740 16024 7084 16064
rect 7124 16024 7133 16064
rect 8515 16024 8524 16064
rect 8564 16024 10444 16064
rect 10484 16024 10493 16064
rect 16579 16024 16588 16064
rect 16628 16024 16637 16064
rect 19363 16024 19372 16064
rect 19412 16024 19852 16064
rect 19892 16024 19901 16064
rect 20131 16024 20140 16064
rect 20180 16024 20189 16064
rect 5731 15980 5789 15981
rect 2500 15940 5740 15980
rect 5780 15940 5789 15980
rect 6499 15940 6508 15980
rect 6548 15940 12076 15980
rect 12116 15940 12125 15980
rect 16195 15940 16204 15980
rect 16244 15940 20852 15980
rect 0 15896 80 15916
rect 2500 15896 2540 15940
rect 5731 15939 5789 15940
rect 18595 15896 18653 15897
rect 20812 15896 20852 15940
rect 21424 15896 21504 15916
rect 0 15856 2540 15896
rect 4919 15856 4928 15896
rect 4968 15856 5010 15896
rect 5050 15856 5092 15896
rect 5132 15856 5174 15896
rect 5214 15856 5256 15896
rect 5296 15856 5305 15896
rect 11395 15856 11404 15896
rect 11444 15856 11453 15896
rect 11875 15856 11884 15896
rect 11924 15856 18604 15896
rect 18644 15856 18653 15896
rect 20039 15856 20048 15896
rect 20088 15856 20130 15896
rect 20170 15856 20212 15896
rect 20252 15856 20294 15896
rect 20334 15856 20376 15896
rect 20416 15856 20425 15896
rect 20812 15856 21504 15896
rect 0 15836 80 15856
rect 11299 15812 11357 15813
rect 11404 15812 11444 15856
rect 18595 15855 18653 15856
rect 21424 15836 21504 15856
rect 4291 15772 4300 15812
rect 4340 15772 4588 15812
rect 4628 15772 6988 15812
rect 7028 15772 7037 15812
rect 11280 15772 11308 15812
rect 11348 15772 11444 15812
rect 11299 15771 11357 15772
rect 7939 15728 7997 15729
rect 4195 15688 4204 15728
rect 4244 15688 6892 15728
rect 6932 15688 6941 15728
rect 7854 15688 7948 15728
rect 7988 15688 7997 15728
rect 8419 15688 8428 15728
rect 8468 15688 10540 15728
rect 10580 15688 10589 15728
rect 11107 15688 11116 15728
rect 11156 15688 12364 15728
rect 12404 15688 12413 15728
rect 12643 15688 12652 15728
rect 12692 15688 12940 15728
rect 12980 15688 12989 15728
rect 17443 15688 17452 15728
rect 17492 15688 17932 15728
rect 17972 15688 17981 15728
rect 19075 15688 19084 15728
rect 19124 15688 19852 15728
rect 19892 15688 19901 15728
rect 7939 15687 7997 15688
rect 20707 15644 20765 15645
rect 6211 15604 6220 15644
rect 6260 15604 11212 15644
rect 11252 15604 11261 15644
rect 11587 15604 11596 15644
rect 11636 15604 14284 15644
rect 14324 15604 14476 15644
rect 14516 15604 14525 15644
rect 15724 15604 16628 15644
rect 16675 15604 16684 15644
rect 16724 15604 18988 15644
rect 19028 15604 19037 15644
rect 19564 15604 20716 15644
rect 20756 15604 20765 15644
rect 4099 15560 4157 15561
rect 15724 15560 15764 15604
rect 16588 15560 16628 15604
rect 19564 15560 19604 15604
rect 20707 15603 20765 15604
rect 21424 15560 21504 15580
rect 1315 15520 1324 15560
rect 1364 15520 1900 15560
rect 1940 15520 1949 15560
rect 3043 15520 3052 15560
rect 3092 15520 3820 15560
rect 3860 15520 3869 15560
rect 4014 15520 4108 15560
rect 4148 15520 4157 15560
rect 4771 15520 4780 15560
rect 4820 15520 6508 15560
rect 6548 15520 6557 15560
rect 7459 15520 7468 15560
rect 7508 15520 9100 15560
rect 9140 15520 9149 15560
rect 10915 15520 10924 15560
rect 10964 15520 10973 15560
rect 11395 15520 11404 15560
rect 11444 15520 12556 15560
rect 12596 15520 12605 15560
rect 12739 15520 12748 15560
rect 12788 15520 13036 15560
rect 13076 15520 13085 15560
rect 13987 15520 13996 15560
rect 14036 15520 15724 15560
rect 15764 15520 15773 15560
rect 15907 15520 15916 15560
rect 15956 15520 16204 15560
rect 16244 15520 16253 15560
rect 16579 15520 16588 15560
rect 16628 15520 16637 15560
rect 17251 15520 17260 15560
rect 17300 15520 19564 15560
rect 19604 15520 19613 15560
rect 19660 15520 21504 15560
rect 4099 15519 4157 15520
rect 10924 15476 10964 15520
rect 2467 15436 2476 15476
rect 2516 15436 2525 15476
rect 3427 15436 3436 15476
rect 3476 15436 5740 15476
rect 5780 15436 5789 15476
rect 10924 15436 16300 15476
rect 16340 15436 16349 15476
rect 16771 15436 16780 15476
rect 16820 15436 19084 15476
rect 19124 15436 19133 15476
rect 0 15392 80 15412
rect 2476 15392 2516 15436
rect 4291 15392 4349 15393
rect 0 15352 1172 15392
rect 2275 15352 2284 15392
rect 2324 15352 2516 15392
rect 3139 15352 3148 15392
rect 3188 15352 4300 15392
rect 4340 15352 4349 15392
rect 4483 15352 4492 15392
rect 4532 15352 4876 15392
rect 4916 15352 4925 15392
rect 8611 15352 8620 15392
rect 8660 15352 11360 15392
rect 12547 15352 12556 15392
rect 12596 15352 13420 15392
rect 13460 15352 18220 15392
rect 18260 15352 18269 15392
rect 0 15332 80 15352
rect 1132 15308 1172 15352
rect 4291 15351 4349 15352
rect 9379 15308 9437 15309
rect 11320 15308 11360 15352
rect 19660 15308 19700 15520
rect 21424 15500 21504 15520
rect 19843 15436 19852 15476
rect 19892 15436 20180 15476
rect 20140 15392 20180 15436
rect 20140 15352 21388 15392
rect 21428 15352 21437 15392
rect 1132 15268 2860 15308
rect 2900 15268 2909 15308
rect 3619 15268 3628 15308
rect 3668 15268 4108 15308
rect 4148 15268 4157 15308
rect 9379 15268 9388 15308
rect 9428 15268 10924 15308
rect 10964 15268 10973 15308
rect 11320 15268 19700 15308
rect 9379 15267 9437 15268
rect 20803 15224 20861 15225
rect 21424 15224 21504 15244
rect 10819 15184 10828 15224
rect 10868 15184 11980 15224
rect 12020 15184 12029 15224
rect 12556 15184 16684 15224
rect 16724 15184 16733 15224
rect 19555 15184 19564 15224
rect 19604 15184 20044 15224
rect 20084 15184 20093 15224
rect 20803 15184 20812 15224
rect 20852 15184 21504 15224
rect 12556 15141 12596 15184
rect 20803 15183 20861 15184
rect 21424 15164 21504 15184
rect 3235 15140 3293 15141
rect 8035 15140 8093 15141
rect 11011 15140 11069 15141
rect 12547 15140 12605 15141
rect 13891 15140 13949 15141
rect 16291 15140 16349 15141
rect 2947 15100 2956 15140
rect 2996 15100 3244 15140
rect 3284 15100 3293 15140
rect 3679 15100 3688 15140
rect 3728 15100 3770 15140
rect 3810 15100 3852 15140
rect 3892 15100 3934 15140
rect 3974 15100 4016 15140
rect 4056 15100 4065 15140
rect 8035 15100 8044 15140
rect 8084 15100 8908 15140
rect 8948 15100 8957 15140
rect 10723 15100 10732 15140
rect 10772 15100 11020 15140
rect 11060 15100 11069 15140
rect 11299 15100 11308 15140
rect 11348 15100 12556 15140
rect 12596 15100 12605 15140
rect 13027 15100 13036 15140
rect 13076 15100 13612 15140
rect 13652 15100 13661 15140
rect 13891 15100 13900 15140
rect 13940 15100 13996 15140
rect 14036 15100 14045 15140
rect 16206 15100 16300 15140
rect 16340 15100 18604 15140
rect 18644 15100 18653 15140
rect 18799 15100 18808 15140
rect 18848 15100 18890 15140
rect 18930 15100 18972 15140
rect 19012 15100 19054 15140
rect 19094 15100 19136 15140
rect 19176 15100 19185 15140
rect 3235 15099 3293 15100
rect 8035 15099 8093 15100
rect 11011 15099 11069 15100
rect 12547 15099 12605 15100
rect 13891 15099 13949 15100
rect 16291 15099 16349 15100
rect 1315 15016 1324 15056
rect 1364 15016 2380 15056
rect 2420 15016 6796 15056
rect 6836 15016 6845 15056
rect 12364 15016 15340 15056
rect 15380 15016 17836 15056
rect 17876 15016 17885 15056
rect 11299 14972 11357 14973
rect 9283 14932 9292 14972
rect 9332 14932 9676 14972
rect 9716 14932 9725 14972
rect 11299 14932 11308 14972
rect 11348 14932 11357 14972
rect 11299 14931 11357 14932
rect 0 14888 80 14908
rect 11308 14888 11348 14931
rect 0 14848 2540 14888
rect 3235 14848 3244 14888
rect 3284 14848 3293 14888
rect 5635 14848 5644 14888
rect 5684 14848 6892 14888
rect 6932 14848 7468 14888
rect 7508 14848 7517 14888
rect 9187 14848 9196 14888
rect 9236 14848 10772 14888
rect 11308 14848 11404 14888
rect 11444 14848 11453 14888
rect 0 14828 80 14848
rect 2500 14720 2540 14848
rect 3244 14804 3284 14848
rect 10732 14804 10772 14848
rect 12364 14804 12404 15016
rect 12451 14932 12460 14972
rect 12500 14932 13804 14972
rect 13844 14932 13853 14972
rect 14371 14932 14380 14972
rect 14420 14932 15724 14972
rect 15764 14932 16204 14972
rect 16244 14932 16253 14972
rect 18499 14932 18508 14972
rect 18548 14932 19084 14972
rect 19124 14932 19372 14972
rect 19412 14932 20140 14972
rect 20180 14932 20189 14972
rect 17635 14888 17693 14889
rect 21424 14888 21504 14908
rect 12931 14848 12940 14888
rect 12980 14848 14860 14888
rect 14900 14848 14909 14888
rect 17635 14848 17644 14888
rect 17684 14848 21504 14888
rect 17635 14847 17693 14848
rect 21424 14828 21504 14848
rect 16483 14804 16541 14805
rect 18403 14804 18461 14805
rect 3244 14764 4108 14804
rect 4148 14764 4157 14804
rect 6403 14764 6412 14804
rect 6452 14764 8620 14804
rect 8660 14764 8669 14804
rect 9091 14764 9100 14804
rect 9140 14764 10252 14804
rect 10292 14764 10636 14804
rect 10676 14764 10685 14804
rect 10732 14764 12404 14804
rect 13420 14764 14764 14804
rect 14804 14764 14813 14804
rect 16483 14764 16492 14804
rect 16532 14764 18412 14804
rect 18452 14764 18461 14804
rect 13420 14720 13460 14764
rect 16483 14763 16541 14764
rect 18403 14763 18461 14764
rect 19459 14720 19517 14721
rect 2500 14680 11360 14720
rect 12451 14680 12460 14720
rect 12500 14680 12748 14720
rect 12788 14680 13228 14720
rect 13268 14680 13277 14720
rect 13411 14680 13420 14720
rect 13460 14680 13469 14720
rect 13603 14680 13612 14720
rect 13652 14680 14949 14720
rect 14989 14680 14998 14720
rect 15043 14680 15052 14720
rect 15092 14680 15101 14720
rect 15235 14680 15244 14720
rect 15284 14680 15293 14720
rect 19374 14680 19468 14720
rect 19508 14680 19517 14720
rect 11320 14636 11360 14680
rect 15052 14636 15092 14680
rect 3139 14596 3148 14636
rect 3188 14596 3820 14636
rect 3860 14596 3869 14636
rect 5731 14596 5740 14636
rect 5780 14596 8140 14636
rect 8180 14596 8189 14636
rect 11320 14596 13804 14636
rect 13844 14596 13853 14636
rect 14083 14596 14092 14636
rect 14132 14596 15092 14636
rect 15244 14552 15284 14680
rect 19459 14679 19517 14680
rect 16675 14636 16733 14637
rect 16675 14596 16684 14636
rect 16724 14596 18604 14636
rect 18644 14596 18653 14636
rect 16675 14595 16733 14596
rect 21424 14552 21504 14572
rect 2659 14512 2668 14552
rect 2708 14512 3532 14552
rect 3572 14512 3581 14552
rect 4387 14512 4396 14552
rect 4436 14512 10732 14552
rect 10772 14512 10781 14552
rect 12643 14512 12652 14552
rect 12692 14512 15628 14552
rect 15668 14512 15677 14552
rect 16675 14512 16684 14552
rect 16724 14512 16972 14552
rect 17012 14512 20236 14552
rect 20276 14512 20285 14552
rect 21100 14512 21504 14552
rect 21100 14468 21140 14512
rect 21424 14492 21504 14512
rect 1804 14428 13036 14468
rect 13076 14428 13085 14468
rect 14659 14428 14668 14468
rect 14708 14428 14860 14468
rect 14900 14428 14909 14468
rect 17731 14428 17740 14468
rect 17780 14428 18412 14468
rect 18452 14428 18461 14468
rect 18595 14428 18604 14468
rect 18644 14428 21140 14468
rect 0 14384 80 14404
rect 1804 14384 1844 14428
rect 3427 14384 3485 14385
rect 0 14344 1844 14384
rect 2755 14344 2764 14384
rect 2804 14344 3244 14384
rect 3284 14344 3293 14384
rect 3427 14344 3436 14384
rect 3476 14344 3532 14384
rect 3572 14344 3581 14384
rect 4919 14344 4928 14384
rect 4968 14344 5010 14384
rect 5050 14344 5092 14384
rect 5132 14344 5174 14384
rect 5214 14344 5256 14384
rect 5296 14344 5305 14384
rect 11320 14344 18700 14384
rect 18740 14344 18749 14384
rect 20039 14344 20048 14384
rect 20088 14344 20130 14384
rect 20170 14344 20212 14384
rect 20252 14344 20294 14384
rect 20334 14344 20376 14384
rect 20416 14344 20425 14384
rect 0 14324 80 14344
rect 3427 14343 3485 14344
rect 6499 14300 6557 14301
rect 11320 14300 11360 14344
rect 13891 14300 13949 14301
rect 14947 14300 15005 14301
rect 6019 14260 6028 14300
rect 6068 14260 6508 14300
rect 6548 14260 11360 14300
rect 12259 14260 12268 14300
rect 12308 14260 13900 14300
rect 13940 14260 14092 14300
rect 14132 14260 14141 14300
rect 14275 14260 14284 14300
rect 14324 14260 14764 14300
rect 14804 14260 14813 14300
rect 14947 14260 14956 14300
rect 14996 14260 20180 14300
rect 6499 14259 6557 14260
rect 13891 14259 13949 14260
rect 14947 14259 15005 14260
rect 7267 14216 7325 14217
rect 2947 14176 2956 14216
rect 2996 14176 3340 14216
rect 3380 14176 3389 14216
rect 3907 14176 3916 14216
rect 3956 14176 4588 14216
rect 4628 14176 7276 14216
rect 7316 14176 7325 14216
rect 7267 14175 7325 14176
rect 8803 14216 8861 14217
rect 14659 14216 14717 14217
rect 20140 14216 20180 14260
rect 21424 14216 21504 14236
rect 8803 14176 8812 14216
rect 8852 14176 8946 14216
rect 12931 14176 12940 14216
rect 12980 14176 14188 14216
rect 14228 14176 14237 14216
rect 14659 14176 14668 14216
rect 14708 14176 14956 14216
rect 14996 14176 15005 14216
rect 18403 14176 18412 14216
rect 18452 14176 19948 14216
rect 19988 14176 19997 14216
rect 20140 14176 21504 14216
rect 8803 14175 8861 14176
rect 14659 14175 14717 14176
rect 21424 14156 21504 14176
rect 7075 14132 7133 14133
rect 11683 14132 11741 14133
rect 1603 14092 1612 14132
rect 1652 14092 2092 14132
rect 2132 14092 2141 14132
rect 4675 14092 4684 14132
rect 4724 14092 6508 14132
rect 6548 14092 7084 14132
rect 7124 14092 7133 14132
rect 7075 14091 7133 14092
rect 7180 14092 9100 14132
rect 9140 14092 9149 14132
rect 9283 14092 9292 14132
rect 9332 14092 9772 14132
rect 9812 14092 9821 14132
rect 11683 14092 11692 14132
rect 11732 14092 17644 14132
rect 17684 14092 17693 14132
rect 19555 14092 19564 14132
rect 19604 14092 20140 14132
rect 20180 14092 20189 14132
rect 3043 14048 3101 14049
rect 355 14008 364 14048
rect 404 14008 3052 14048
rect 3092 14008 3101 14048
rect 3043 14007 3101 14008
rect 5923 14048 5981 14049
rect 7180 14048 7220 14092
rect 11683 14091 11741 14092
rect 5923 14008 5932 14048
rect 5972 14008 6028 14048
rect 6068 14008 6077 14048
rect 6979 14008 6988 14048
rect 7028 14008 7220 14048
rect 7555 14008 7564 14048
rect 7604 14008 9580 14048
rect 9620 14008 9629 14048
rect 13219 14008 13228 14048
rect 13268 14008 14476 14048
rect 14516 14008 14525 14048
rect 14659 14008 14668 14048
rect 14708 14008 17260 14048
rect 17300 14008 17309 14048
rect 18883 14008 18892 14048
rect 18932 14008 19948 14048
rect 19988 14008 19997 14048
rect 5923 14007 5981 14008
rect 2851 13964 2909 13965
rect 8515 13964 8573 13965
rect 16675 13964 16733 13965
rect 1507 13924 1516 13964
rect 1556 13924 2860 13964
rect 2900 13924 2909 13964
rect 4099 13924 4108 13964
rect 4148 13924 4188 13964
rect 8515 13924 8524 13964
rect 8564 13924 11020 13964
rect 11060 13924 11069 13964
rect 11203 13924 11212 13964
rect 11252 13924 14764 13964
rect 14804 13924 16684 13964
rect 16724 13924 16733 13964
rect 17155 13924 17164 13964
rect 17204 13924 20180 13964
rect 2851 13923 2909 13924
rect 0 13880 80 13900
rect 4108 13880 4148 13924
rect 8515 13923 8573 13924
rect 16675 13923 16733 13924
rect 12163 13880 12221 13881
rect 14755 13880 14813 13881
rect 15619 13880 15677 13881
rect 20140 13880 20180 13924
rect 21424 13880 21504 13900
rect 0 13840 172 13880
rect 212 13840 221 13880
rect 1699 13840 1708 13880
rect 1748 13840 2092 13880
rect 2132 13840 2141 13880
rect 2851 13840 2860 13880
rect 2900 13840 4396 13880
rect 4436 13840 4445 13880
rect 5539 13840 5548 13880
rect 5588 13840 5836 13880
rect 5876 13840 5885 13880
rect 6211 13840 6220 13880
rect 6260 13840 11360 13880
rect 12078 13840 12172 13880
rect 12212 13840 12221 13880
rect 12355 13840 12364 13880
rect 12404 13840 14764 13880
rect 14804 13840 14813 13880
rect 14947 13840 14956 13880
rect 14996 13840 15628 13880
rect 15668 13840 15677 13880
rect 15811 13840 15820 13880
rect 15860 13840 17068 13880
rect 17108 13840 17117 13880
rect 20140 13840 21504 13880
rect 0 13820 80 13840
rect 11320 13796 11360 13840
rect 12163 13839 12221 13840
rect 14755 13839 14813 13840
rect 15619 13839 15677 13840
rect 21424 13820 21504 13840
rect 15715 13796 15773 13797
rect 3235 13756 3244 13796
rect 3284 13756 6604 13796
rect 6644 13756 6653 13796
rect 7747 13756 7756 13796
rect 7796 13756 8716 13796
rect 8756 13756 8765 13796
rect 11320 13756 12844 13796
rect 12884 13756 15724 13796
rect 15764 13756 15773 13796
rect 15715 13755 15773 13756
rect 3043 13712 3101 13713
rect 9187 13712 9245 13713
rect 3043 13672 3052 13712
rect 3092 13672 3340 13712
rect 3380 13672 3389 13712
rect 7555 13672 7564 13712
rect 7604 13672 8044 13712
rect 8084 13672 8093 13712
rect 8899 13672 8908 13712
rect 8948 13672 9196 13712
rect 9236 13672 9484 13712
rect 9524 13672 9533 13712
rect 14179 13672 14188 13712
rect 14228 13672 14476 13712
rect 14516 13672 14525 13712
rect 3043 13671 3101 13672
rect 9187 13671 9245 13672
rect 6499 13628 6557 13629
rect 8611 13628 8669 13629
rect 3679 13588 3688 13628
rect 3728 13588 3770 13628
rect 3810 13588 3852 13628
rect 3892 13588 3934 13628
rect 3974 13588 4016 13628
rect 4056 13588 4065 13628
rect 6499 13588 6508 13628
rect 6548 13588 6604 13628
rect 6644 13588 6653 13628
rect 8526 13588 8620 13628
rect 8660 13588 8669 13628
rect 15427 13588 15436 13628
rect 15476 13588 16972 13628
rect 17012 13588 17021 13628
rect 18799 13588 18808 13628
rect 18848 13588 18890 13628
rect 18930 13588 18972 13628
rect 19012 13588 19054 13628
rect 19094 13588 19136 13628
rect 19176 13588 19185 13628
rect 6499 13587 6557 13588
rect 8611 13587 8669 13588
rect 10531 13544 10589 13545
rect 17827 13544 17885 13545
rect 21424 13544 21504 13564
rect 2500 13504 7604 13544
rect 8515 13504 8524 13544
rect 8564 13504 8716 13544
rect 8756 13504 8765 13544
rect 10051 13504 10060 13544
rect 10100 13504 10540 13544
rect 10580 13504 10589 13544
rect 11683 13504 11692 13544
rect 11732 13504 11980 13544
rect 12020 13504 15148 13544
rect 15188 13504 15197 13544
rect 15244 13504 17836 13544
rect 17876 13504 17885 13544
rect 20611 13504 20620 13544
rect 20660 13504 21504 13544
rect 739 13460 797 13461
rect 2500 13460 2540 13504
rect 7564 13460 7604 13504
rect 10531 13503 10589 13504
rect 739 13420 748 13460
rect 788 13420 2540 13460
rect 7075 13420 7084 13460
rect 7124 13420 7468 13460
rect 7508 13420 7517 13460
rect 7564 13420 10676 13460
rect 10723 13420 10732 13460
rect 10772 13420 12460 13460
rect 12500 13420 12748 13460
rect 12788 13420 12797 13460
rect 739 13419 797 13420
rect 0 13376 80 13396
rect 10636 13376 10676 13420
rect 11299 13376 11357 13377
rect 15244 13376 15284 13504
rect 17827 13503 17885 13504
rect 21424 13484 21504 13504
rect 15523 13420 15532 13460
rect 15572 13420 16108 13460
rect 16148 13420 16157 13460
rect 0 13336 10444 13376
rect 10484 13336 10493 13376
rect 10636 13336 11308 13376
rect 11348 13336 11357 13376
rect 11683 13336 11692 13376
rect 11732 13336 15284 13376
rect 15907 13336 15916 13376
rect 15956 13336 16972 13376
rect 17012 13336 17021 13376
rect 0 13316 80 13336
rect 11299 13335 11357 13336
rect 1411 13292 1469 13293
rect 1411 13252 1420 13292
rect 1460 13252 6508 13292
rect 6548 13252 6557 13292
rect 10339 13252 10348 13292
rect 10388 13252 10397 13292
rect 16579 13252 16588 13292
rect 16628 13252 17356 13292
rect 17396 13252 17405 13292
rect 18211 13252 18220 13292
rect 18260 13252 20180 13292
rect 1411 13251 1469 13252
rect 9475 13208 9533 13209
rect 3715 13168 3724 13208
rect 3764 13168 4108 13208
rect 4148 13168 4157 13208
rect 5635 13168 5644 13208
rect 5684 13168 9484 13208
rect 9524 13168 9580 13208
rect 9620 13168 9629 13208
rect 9475 13167 9533 13168
rect 931 13084 940 13124
rect 980 13084 2572 13124
rect 2612 13084 2621 13124
rect 6316 13084 10060 13124
rect 10100 13084 10109 13124
rect 6316 12956 6356 13084
rect 7555 13040 7613 13041
rect 10348 13040 10388 13252
rect 20140 13208 20180 13252
rect 21424 13208 21504 13228
rect 11107 13168 11116 13208
rect 11156 13168 11360 13208
rect 14755 13168 14764 13208
rect 14804 13168 15052 13208
rect 15092 13168 15244 13208
rect 15284 13168 16780 13208
rect 16820 13168 16829 13208
rect 18595 13168 18604 13208
rect 18644 13168 19564 13208
rect 19604 13168 19613 13208
rect 20140 13168 21504 13208
rect 11320 13124 11360 13168
rect 21424 13148 21504 13168
rect 16483 13124 16541 13125
rect 11320 13084 12556 13124
rect 12596 13084 13132 13124
rect 13172 13084 13181 13124
rect 13699 13084 13708 13124
rect 13748 13084 15532 13124
rect 15572 13084 15581 13124
rect 16398 13084 16492 13124
rect 16532 13084 16541 13124
rect 16483 13083 16541 13084
rect 7267 13000 7276 13040
rect 7316 13000 7564 13040
rect 7604 13000 7613 13040
rect 8323 13000 8332 13040
rect 8372 13000 8524 13040
rect 8564 13000 8573 13040
rect 10348 13000 10732 13040
rect 10772 13000 10781 13040
rect 17827 13000 17836 13040
rect 17876 13000 18124 13040
rect 18164 13000 18173 13040
rect 7555 12999 7613 13000
rect 364 12916 6356 12956
rect 15043 12916 15052 12956
rect 15092 12916 15724 12956
rect 15764 12916 15773 12956
rect 0 12872 80 12892
rect 364 12872 404 12916
rect 12163 12872 12221 12873
rect 21424 12872 21504 12892
rect 0 12832 404 12872
rect 4919 12832 4928 12872
rect 4968 12832 5010 12872
rect 5050 12832 5092 12872
rect 5132 12832 5174 12872
rect 5214 12832 5256 12872
rect 5296 12832 5305 12872
rect 5443 12832 5452 12872
rect 5492 12832 6220 12872
rect 6260 12832 6269 12872
rect 12078 12832 12172 12872
rect 12212 12832 12221 12872
rect 17059 12832 17068 12872
rect 17108 12832 17356 12872
rect 17396 12832 17405 12872
rect 20039 12832 20048 12872
rect 20088 12832 20130 12872
rect 20170 12832 20212 12872
rect 20252 12832 20294 12872
rect 20334 12832 20376 12872
rect 20416 12832 20425 12872
rect 20812 12832 21504 12872
rect 0 12812 80 12832
rect 12163 12831 12221 12832
rect 20812 12788 20852 12832
rect 21424 12812 21504 12832
rect 11107 12748 11116 12788
rect 11156 12748 20852 12788
rect 18499 12704 18557 12705
rect 10147 12664 10156 12704
rect 10196 12664 12076 12704
rect 12116 12664 12125 12704
rect 13795 12664 13804 12704
rect 13844 12664 18508 12704
rect 18548 12664 18557 12704
rect 18499 12663 18557 12664
rect 3139 12620 3197 12621
rect 12163 12620 12221 12621
rect 13123 12620 13181 12621
rect 2275 12580 2284 12620
rect 2324 12580 2764 12620
rect 2804 12580 2813 12620
rect 3139 12580 3148 12620
rect 3188 12580 7660 12620
rect 7700 12580 7709 12620
rect 7843 12580 7852 12620
rect 7892 12580 11360 12620
rect 3139 12579 3197 12580
rect 3427 12536 3485 12537
rect 11320 12536 11360 12580
rect 12163 12580 12172 12620
rect 12212 12580 12844 12620
rect 12884 12580 12893 12620
rect 13038 12580 13132 12620
rect 13172 12580 13181 12620
rect 12163 12579 12221 12580
rect 13123 12579 13181 12580
rect 14659 12620 14717 12621
rect 18307 12620 18365 12621
rect 14659 12580 14668 12620
rect 14708 12580 18316 12620
rect 18356 12580 18365 12620
rect 14659 12579 14717 12580
rect 18307 12579 18365 12580
rect 16483 12536 16541 12537
rect 21424 12536 21504 12556
rect 2284 12496 2476 12536
rect 2516 12496 2525 12536
rect 3427 12496 3436 12536
rect 3476 12496 3532 12536
rect 3572 12496 3581 12536
rect 3907 12496 3916 12536
rect 3956 12496 5932 12536
rect 5972 12496 5981 12536
rect 6115 12496 6124 12536
rect 6164 12496 6412 12536
rect 6452 12496 6461 12536
rect 7459 12496 7468 12536
rect 7508 12496 7948 12536
rect 7988 12496 7997 12536
rect 8803 12496 8812 12536
rect 8852 12496 9292 12536
rect 9332 12496 9341 12536
rect 9571 12496 9580 12536
rect 9620 12496 10060 12536
rect 10100 12496 10109 12536
rect 11320 12496 12268 12536
rect 12308 12496 12317 12536
rect 13027 12496 13036 12536
rect 13076 12496 13324 12536
rect 13364 12496 13516 12536
rect 13556 12496 13565 12536
rect 15619 12496 15628 12536
rect 15668 12496 16492 12536
rect 16532 12496 17452 12536
rect 17492 12496 17501 12536
rect 18211 12496 18220 12536
rect 18260 12496 19564 12536
rect 19604 12496 19613 12536
rect 20140 12496 21504 12536
rect 0 12368 80 12388
rect 1219 12368 1277 12369
rect 2284 12368 2324 12496
rect 3427 12495 3485 12496
rect 6412 12368 6452 12496
rect 16483 12495 16541 12496
rect 8035 12452 8093 12453
rect 8035 12412 8044 12452
rect 8084 12412 13420 12452
rect 13460 12412 13469 12452
rect 13603 12412 13612 12452
rect 13652 12412 13804 12452
rect 13844 12412 13853 12452
rect 16099 12412 16108 12452
rect 16148 12412 17356 12452
rect 17396 12412 17405 12452
rect 18979 12412 18988 12452
rect 19028 12412 19660 12452
rect 19700 12412 19948 12452
rect 19988 12412 19997 12452
rect 8035 12411 8093 12412
rect 20140 12368 20180 12496
rect 21424 12476 21504 12496
rect 0 12328 1228 12368
rect 1268 12328 1277 12368
rect 2275 12328 2284 12368
rect 2324 12328 2333 12368
rect 6412 12328 9004 12368
rect 9044 12328 9053 12368
rect 11320 12328 20180 12368
rect 0 12308 80 12328
rect 1219 12327 1277 12328
rect 11320 12284 11360 12328
rect 3811 12244 3820 12284
rect 3860 12244 3869 12284
rect 5155 12244 5164 12284
rect 5204 12244 6124 12284
rect 6164 12244 6700 12284
rect 6740 12244 6892 12284
rect 6932 12244 6941 12284
rect 6988 12244 11360 12284
rect 11587 12244 11596 12284
rect 11636 12244 18412 12284
rect 18452 12244 18461 12284
rect 3820 12200 3860 12244
rect 6988 12200 7028 12244
rect 3820 12160 4492 12200
rect 4532 12160 7028 12200
rect 8611 12200 8669 12201
rect 15715 12200 15773 12201
rect 16099 12200 16157 12201
rect 8611 12160 8620 12200
rect 8660 12160 8716 12200
rect 8756 12160 8765 12200
rect 9283 12160 9292 12200
rect 9332 12160 15668 12200
rect 8611 12159 8669 12160
rect 3235 12116 3293 12117
rect 7939 12116 7997 12117
rect 15628 12116 15668 12160
rect 15715 12160 15724 12200
rect 15764 12160 15820 12200
rect 15860 12160 15869 12200
rect 16003 12160 16012 12200
rect 16052 12160 16108 12200
rect 16148 12160 16157 12200
rect 15715 12159 15773 12160
rect 16099 12159 16157 12160
rect 17731 12200 17789 12201
rect 21424 12200 21504 12220
rect 17731 12160 17740 12200
rect 17780 12160 17932 12200
rect 17972 12160 17981 12200
rect 18691 12160 18700 12200
rect 18740 12160 21504 12200
rect 17731 12159 17789 12160
rect 21424 12140 21504 12160
rect 17827 12116 17885 12117
rect 3150 12076 3244 12116
rect 3284 12076 3293 12116
rect 3679 12076 3688 12116
rect 3728 12076 3770 12116
rect 3810 12076 3852 12116
rect 3892 12076 3934 12116
rect 3974 12076 4016 12116
rect 4056 12076 4065 12116
rect 5260 12076 7948 12116
rect 7988 12076 7997 12116
rect 8611 12076 8620 12116
rect 8660 12076 10060 12116
rect 10100 12076 10109 12116
rect 11491 12076 11500 12116
rect 11540 12076 11788 12116
rect 11828 12076 15052 12116
rect 15092 12076 15101 12116
rect 15628 12076 17836 12116
rect 17876 12076 17885 12116
rect 18799 12076 18808 12116
rect 18848 12076 18890 12116
rect 18930 12076 18972 12116
rect 19012 12076 19054 12116
rect 19094 12076 19136 12116
rect 19176 12076 19185 12116
rect 3235 12075 3293 12076
rect 5260 11948 5300 12076
rect 7939 12075 7997 12076
rect 17827 12075 17885 12076
rect 17836 12032 17876 12075
rect 5443 11992 5452 12032
rect 5492 11992 10828 12032
rect 10868 11992 11596 12032
rect 11636 11992 11645 12032
rect 12547 11992 12556 12032
rect 12596 11992 13036 12032
rect 13076 11992 13085 12032
rect 13219 11992 13228 12032
rect 13268 11992 13612 12032
rect 13652 11992 13661 12032
rect 14083 11992 14092 12032
rect 14132 11992 14860 12032
rect 14900 11992 16780 12032
rect 16820 11992 16829 12032
rect 17836 11992 19660 12032
rect 19700 11992 19709 12032
rect 1228 11908 5300 11948
rect 5731 11948 5789 11949
rect 5731 11908 5740 11948
rect 5780 11908 9196 11948
rect 9236 11908 9245 11948
rect 9475 11908 9484 11948
rect 9524 11908 16876 11948
rect 16916 11908 16925 11948
rect 0 11864 80 11884
rect 1228 11864 1268 11908
rect 5731 11907 5789 11908
rect 7459 11864 7517 11865
rect 0 11824 1268 11864
rect 1315 11824 1324 11864
rect 1364 11824 5836 11864
rect 5876 11824 7468 11864
rect 7508 11824 7517 11864
rect 0 11804 80 11824
rect 7459 11823 7517 11824
rect 9484 11780 9524 11908
rect 21424 11864 21504 11884
rect 9571 11824 9580 11864
rect 9620 11824 10444 11864
rect 10484 11824 10493 11864
rect 11875 11824 11884 11864
rect 11924 11824 11933 11864
rect 13987 11824 13996 11864
rect 14036 11824 14045 11864
rect 14563 11824 14572 11864
rect 14612 11824 14860 11864
rect 14900 11824 14909 11864
rect 15523 11824 15532 11864
rect 15572 11824 18700 11864
rect 18740 11824 18749 11864
rect 20140 11824 21504 11864
rect 5923 11740 5932 11780
rect 5972 11740 9524 11780
rect 2467 11656 2476 11696
rect 2516 11656 8564 11696
rect 9187 11656 9196 11696
rect 9236 11656 9428 11696
rect 9859 11656 9868 11696
rect 9908 11656 10060 11696
rect 10100 11656 10109 11696
rect 4099 11612 4157 11613
rect 2500 11572 4108 11612
rect 4148 11572 4157 11612
rect 8524 11612 8564 11656
rect 9388 11612 9428 11656
rect 8524 11572 9292 11612
rect 9332 11572 9341 11612
rect 9388 11572 9772 11612
rect 9812 11572 9821 11612
rect 2500 11528 2540 11572
rect 4099 11571 4157 11572
rect 5635 11528 5693 11529
rect 1411 11488 1420 11528
rect 1460 11488 2540 11528
rect 2668 11488 5644 11528
rect 5684 11488 5693 11528
rect 7075 11488 7084 11528
rect 7124 11488 11788 11528
rect 11828 11488 11837 11528
rect 2668 11444 2708 11488
rect 5635 11487 5693 11488
rect 8323 11444 8381 11445
rect 11884 11444 11924 11824
rect 13996 11780 14036 11824
rect 20140 11780 20180 11824
rect 21424 11804 21504 11824
rect 12739 11740 12748 11780
rect 12788 11740 14036 11780
rect 15715 11740 15724 11780
rect 15764 11740 20180 11780
rect 17827 11696 17885 11697
rect 18499 11696 18557 11697
rect 13315 11656 13324 11696
rect 13364 11656 14476 11696
rect 14516 11656 14525 11696
rect 15139 11656 15148 11696
rect 15188 11656 16300 11696
rect 16340 11656 16780 11696
rect 16820 11656 16829 11696
rect 17827 11656 17836 11696
rect 17876 11656 18124 11696
rect 18164 11656 18173 11696
rect 18499 11656 18508 11696
rect 18548 11656 19084 11696
rect 19124 11656 19133 11696
rect 19267 11656 19276 11696
rect 19316 11656 19756 11696
rect 19796 11656 19805 11696
rect 20035 11656 20044 11696
rect 20084 11656 20093 11696
rect 17827 11655 17885 11656
rect 18499 11655 18557 11656
rect 12067 11612 12125 11613
rect 12835 11612 12893 11613
rect 13123 11612 13181 11613
rect 20044 11612 20084 11656
rect 12067 11572 12076 11612
rect 12116 11572 12210 11612
rect 12835 11572 12844 11612
rect 12884 11572 13132 11612
rect 13172 11572 13420 11612
rect 13460 11572 14284 11612
rect 14324 11572 14333 11612
rect 17731 11572 17740 11612
rect 17780 11572 17789 11612
rect 18307 11572 18316 11612
rect 18356 11572 18700 11612
rect 18740 11572 20084 11612
rect 12067 11571 12125 11572
rect 12835 11571 12893 11572
rect 13123 11571 13181 11572
rect 16579 11528 16637 11529
rect 12835 11488 12844 11528
rect 12884 11488 13612 11528
rect 13652 11488 13661 11528
rect 13891 11488 13900 11528
rect 13940 11488 14380 11528
rect 14420 11488 14429 11528
rect 16579 11488 16588 11528
rect 16628 11488 16876 11528
rect 16916 11488 16925 11528
rect 16579 11487 16637 11488
rect 2500 11404 2708 11444
rect 8238 11404 8332 11444
rect 8372 11404 8381 11444
rect 0 11360 80 11380
rect 2500 11360 2540 11404
rect 8323 11403 8381 11404
rect 11788 11404 11924 11444
rect 11980 11404 12748 11444
rect 12788 11404 13460 11444
rect 13507 11404 13516 11444
rect 13556 11404 14092 11444
rect 14132 11404 14141 11444
rect 14467 11404 14476 11444
rect 14516 11404 14956 11444
rect 14996 11404 15005 11444
rect 4579 11360 4637 11361
rect 9187 11360 9245 11361
rect 0 11320 2540 11360
rect 4494 11320 4588 11360
rect 4628 11320 4637 11360
rect 4919 11320 4928 11360
rect 4968 11320 5010 11360
rect 5050 11320 5092 11360
rect 5132 11320 5174 11360
rect 5214 11320 5256 11360
rect 5296 11320 5305 11360
rect 9102 11320 9196 11360
rect 9236 11320 9245 11360
rect 0 11300 80 11320
rect 4579 11319 4637 11320
rect 9187 11319 9245 11320
rect 547 11236 556 11276
rect 596 11236 2540 11276
rect 2659 11236 2668 11276
rect 2708 11236 4300 11276
rect 4340 11236 4349 11276
rect 8419 11236 8428 11276
rect 8468 11236 9484 11276
rect 9524 11236 9533 11276
rect 2500 11192 2540 11236
rect 8803 11192 8861 11193
rect 11788 11192 11828 11404
rect 11980 11360 12020 11404
rect 13420 11360 13460 11404
rect 11875 11320 11884 11360
rect 11924 11320 12020 11360
rect 13380 11320 13420 11360
rect 13460 11320 13469 11360
rect 17740 11276 17780 11572
rect 21424 11528 21504 11548
rect 20140 11488 21504 11528
rect 18499 11444 18557 11445
rect 20140 11444 20180 11488
rect 21424 11468 21504 11488
rect 18499 11404 18508 11444
rect 18548 11404 20180 11444
rect 18499 11403 18557 11404
rect 20039 11320 20048 11360
rect 20088 11320 20130 11360
rect 20170 11320 20212 11360
rect 20252 11320 20294 11360
rect 20334 11320 20376 11360
rect 20416 11320 20425 11360
rect 15715 11236 15724 11276
rect 15764 11236 17780 11276
rect 12067 11192 12125 11193
rect 17923 11192 17981 11193
rect 21424 11192 21504 11212
rect 2500 11152 3052 11192
rect 3092 11152 3101 11192
rect 3715 11152 3724 11192
rect 3764 11152 4972 11192
rect 5012 11152 5021 11192
rect 7267 11152 7276 11192
rect 7316 11152 8236 11192
rect 8276 11152 8285 11192
rect 8803 11152 8812 11192
rect 8852 11152 9004 11192
rect 9044 11152 9053 11192
rect 11788 11152 11884 11192
rect 11924 11152 11933 11192
rect 12067 11152 12076 11192
rect 12116 11152 12364 11192
rect 12404 11152 12413 11192
rect 12739 11152 12748 11192
rect 12788 11152 14572 11192
rect 14612 11152 14621 11192
rect 17731 11152 17740 11192
rect 17780 11152 17932 11192
rect 17972 11152 17981 11192
rect 19459 11152 19468 11192
rect 19508 11152 20044 11192
rect 20084 11152 20093 11192
rect 21283 11152 21292 11192
rect 21332 11152 21504 11192
rect 8803 11151 8861 11152
rect 12067 11151 12125 11152
rect 17923 11151 17981 11152
rect 21424 11132 21504 11152
rect 8323 11108 8381 11109
rect 17731 11108 17789 11109
rect 1603 11068 1612 11108
rect 1652 11068 8332 11108
rect 8372 11068 11788 11108
rect 11828 11068 12172 11108
rect 12212 11068 17356 11108
rect 17396 11068 17405 11108
rect 17731 11068 17740 11108
rect 17780 11068 18028 11108
rect 18068 11068 19948 11108
rect 19988 11068 19997 11108
rect 7084 11024 7124 11068
rect 8323 11067 8381 11068
rect 17731 11067 17789 11068
rect 9379 11024 9437 11025
rect 1219 10984 1228 11024
rect 1268 10984 2188 11024
rect 2228 10984 2237 11024
rect 4483 10984 4492 11024
rect 4532 10984 4876 11024
rect 4916 10984 4925 11024
rect 5155 10984 5164 11024
rect 5204 10984 6316 11024
rect 6356 10984 6365 11024
rect 7075 10984 7084 11024
rect 7124 10984 7133 11024
rect 7939 10984 7948 11024
rect 7988 10984 8332 11024
rect 8372 10984 8716 11024
rect 8756 10984 8765 11024
rect 8899 10984 8908 11024
rect 8948 10984 9388 11024
rect 9428 10984 9437 11024
rect 11587 10984 11596 11024
rect 11636 10984 13132 11024
rect 13172 10984 13181 11024
rect 17827 10984 17836 11024
rect 17876 10984 19852 11024
rect 19892 10984 19901 11024
rect 9379 10983 9437 10984
rect 17443 10940 17501 10941
rect 1315 10900 1324 10940
rect 1364 10900 1900 10940
rect 1940 10900 1949 10940
rect 2500 10900 17452 10940
rect 17492 10900 17501 10940
rect 17923 10900 17932 10940
rect 17972 10900 18796 10940
rect 18836 10900 18845 10940
rect 0 10856 80 10876
rect 2500 10856 2540 10900
rect 17443 10899 17501 10900
rect 12451 10856 12509 10857
rect 12835 10856 12893 10857
rect 21424 10856 21504 10876
rect 0 10816 2540 10856
rect 3715 10816 3724 10856
rect 3764 10816 3773 10856
rect 4387 10816 4396 10856
rect 4436 10816 5068 10856
rect 5108 10816 5117 10856
rect 12366 10816 12460 10856
rect 12500 10816 12509 10856
rect 12750 10816 12844 10856
rect 12884 10816 12893 10856
rect 18019 10816 18028 10856
rect 18068 10816 18508 10856
rect 18548 10816 18557 10856
rect 20140 10816 21504 10856
rect 0 10796 80 10816
rect 3235 10772 3293 10773
rect 2563 10732 2572 10772
rect 2612 10732 3244 10772
rect 3284 10732 3293 10772
rect 3235 10731 3293 10732
rect 3724 10688 3764 10816
rect 12451 10815 12509 10816
rect 12835 10815 12893 10816
rect 4771 10772 4829 10773
rect 18211 10772 18269 10773
rect 3811 10732 3820 10772
rect 3860 10732 4492 10772
rect 4532 10732 4541 10772
rect 4675 10732 4684 10772
rect 4724 10732 4780 10772
rect 4820 10732 7084 10772
rect 7124 10732 7133 10772
rect 8899 10732 8908 10772
rect 8948 10732 9388 10772
rect 9428 10732 9437 10772
rect 13219 10732 13228 10772
rect 13268 10732 18220 10772
rect 18260 10732 18269 10772
rect 4771 10731 4829 10732
rect 18211 10731 18269 10732
rect 11299 10688 11357 10689
rect 19747 10688 19805 10689
rect 3532 10648 3764 10688
rect 6892 10648 10924 10688
rect 10964 10648 10973 10688
rect 11299 10648 11308 10688
rect 11348 10648 14572 10688
rect 14612 10648 14621 10688
rect 15139 10648 15148 10688
rect 15188 10648 16012 10688
rect 16052 10648 16061 10688
rect 16675 10648 16684 10688
rect 16724 10648 19756 10688
rect 19796 10648 19805 10688
rect 3532 10604 3572 10648
rect 2659 10564 2668 10604
rect 2708 10564 3572 10604
rect 3679 10564 3688 10604
rect 3728 10564 3770 10604
rect 3810 10564 3852 10604
rect 3892 10564 3934 10604
rect 3974 10564 4016 10604
rect 4056 10564 4065 10604
rect 3043 10396 3052 10436
rect 3092 10396 4396 10436
rect 4436 10396 4445 10436
rect 0 10352 80 10372
rect 6892 10352 6932 10648
rect 11299 10647 11357 10648
rect 19747 10647 19805 10648
rect 10147 10564 10156 10604
rect 10196 10564 11308 10604
rect 11348 10564 11357 10604
rect 12931 10564 12940 10604
rect 12980 10564 13708 10604
rect 13748 10564 13757 10604
rect 14083 10564 14092 10604
rect 14132 10564 15724 10604
rect 15764 10564 15773 10604
rect 16300 10564 17932 10604
rect 17972 10564 18508 10604
rect 18548 10564 18557 10604
rect 18799 10564 18808 10604
rect 18848 10564 18890 10604
rect 18930 10564 18972 10604
rect 19012 10564 19054 10604
rect 19094 10564 19136 10604
rect 19176 10564 19185 10604
rect 9475 10520 9533 10521
rect 8995 10480 9004 10520
rect 9044 10480 9196 10520
rect 9236 10480 9484 10520
rect 9524 10480 9533 10520
rect 9475 10479 9533 10480
rect 10627 10520 10685 10521
rect 16300 10520 16340 10564
rect 20140 10520 20180 10816
rect 21424 10796 21504 10816
rect 10627 10480 10636 10520
rect 10676 10480 11404 10520
rect 11444 10480 13228 10520
rect 13268 10480 13277 10520
rect 13507 10480 13516 10520
rect 13556 10480 14188 10520
rect 14228 10480 14237 10520
rect 15427 10480 15436 10520
rect 15476 10480 16340 10520
rect 18211 10480 18220 10520
rect 18260 10480 20180 10520
rect 20707 10520 20765 10521
rect 21424 10520 21504 10540
rect 20707 10480 20716 10520
rect 20756 10480 21504 10520
rect 10627 10479 10685 10480
rect 20707 10479 20765 10480
rect 21424 10460 21504 10480
rect 9091 10436 9149 10437
rect 8227 10396 8236 10436
rect 8276 10396 8812 10436
rect 8852 10396 8861 10436
rect 9091 10396 9100 10436
rect 9140 10396 9292 10436
rect 9332 10396 9484 10436
rect 9524 10396 9533 10436
rect 9955 10396 9964 10436
rect 10004 10396 10636 10436
rect 10676 10396 10685 10436
rect 10732 10396 20180 10436
rect 9091 10395 9149 10396
rect 0 10312 6932 10352
rect 7555 10312 7564 10352
rect 7604 10312 8044 10352
rect 8084 10312 8093 10352
rect 0 10292 80 10312
rect 9379 10268 9437 10269
rect 10732 10268 10772 10396
rect 18115 10352 18173 10353
rect 10915 10312 10924 10352
rect 10964 10312 18124 10352
rect 18164 10312 18173 10352
rect 18115 10311 18173 10312
rect 18403 10352 18461 10353
rect 18403 10312 18412 10352
rect 18452 10312 19084 10352
rect 19124 10312 19133 10352
rect 18403 10311 18461 10312
rect 1603 10228 1612 10268
rect 1652 10228 2476 10268
rect 2516 10228 2525 10268
rect 7747 10228 7756 10268
rect 7796 10228 8140 10268
rect 8180 10228 8524 10268
rect 8564 10228 8573 10268
rect 9283 10228 9292 10268
rect 9332 10228 9388 10268
rect 9428 10228 9437 10268
rect 9379 10227 9437 10228
rect 9772 10228 10772 10268
rect 11299 10228 11308 10268
rect 11348 10228 15148 10268
rect 15188 10228 15197 10268
rect 15715 10228 15724 10268
rect 15764 10228 16012 10268
rect 16052 10228 16061 10268
rect 17347 10228 17356 10268
rect 17396 10228 17588 10268
rect 18115 10228 18124 10268
rect 18164 10228 18412 10268
rect 18452 10228 18461 10268
rect 4099 10184 4157 10185
rect 9772 10184 9812 10228
rect 10051 10184 10109 10185
rect 17155 10184 17213 10185
rect 17548 10184 17588 10228
rect 20140 10184 20180 10396
rect 21424 10184 21504 10204
rect 1219 10144 1228 10184
rect 1268 10144 2092 10184
rect 2132 10144 2284 10184
rect 2324 10144 2333 10184
rect 4014 10144 4108 10184
rect 4148 10144 4157 10184
rect 7555 10144 7564 10184
rect 7604 10144 7948 10184
rect 7988 10144 7997 10184
rect 8419 10144 8428 10184
rect 8468 10144 9772 10184
rect 9812 10144 9821 10184
rect 10051 10144 10060 10184
rect 10100 10144 11404 10184
rect 11444 10144 11453 10184
rect 13123 10144 13132 10184
rect 13172 10144 17164 10184
rect 17204 10144 17452 10184
rect 17492 10144 17501 10184
rect 17548 10144 18700 10184
rect 18740 10144 18749 10184
rect 20140 10144 21504 10184
rect 4099 10143 4157 10144
rect 10051 10143 10109 10144
rect 17155 10143 17213 10144
rect 21424 10124 21504 10144
rect 2851 10060 2860 10100
rect 2900 10060 3436 10100
rect 3476 10060 3485 10100
rect 8707 10060 8716 10100
rect 8756 10060 9196 10100
rect 9236 10060 9245 10100
rect 10156 10060 10348 10100
rect 10388 10060 10924 10100
rect 10964 10060 10973 10100
rect 11491 10060 11500 10100
rect 11540 10060 12652 10100
rect 12692 10060 13612 10100
rect 13652 10060 13661 10100
rect 14659 10060 14668 10100
rect 14708 10060 14949 10100
rect 14989 10060 14998 10100
rect 15043 10060 15052 10100
rect 15092 10060 18124 10100
rect 18164 10060 18173 10100
rect 18883 10060 18892 10100
rect 18932 10060 19564 10100
rect 19604 10060 19948 10100
rect 19988 10060 19997 10100
rect 3043 10016 3101 10017
rect 10156 10016 10196 10060
rect 3043 9976 3052 10016
rect 3092 9976 3532 10016
rect 3572 9976 8840 10016
rect 9475 9976 9484 10016
rect 9524 9976 10196 10016
rect 11320 9976 21332 10016
rect 3043 9975 3101 9976
rect 6691 9932 6749 9933
rect 2500 9892 6700 9932
rect 6740 9892 6749 9932
rect 8800 9932 8840 9976
rect 11320 9932 11360 9976
rect 8800 9892 11360 9932
rect 15523 9892 15532 9932
rect 15572 9892 16012 9932
rect 16052 9892 16061 9932
rect 16483 9892 16492 9932
rect 16532 9892 17740 9932
rect 17780 9892 17789 9932
rect 0 9848 80 9868
rect 2500 9848 2540 9892
rect 6691 9891 6749 9892
rect 9091 9848 9149 9849
rect 12739 9848 12797 9849
rect 21292 9848 21332 9976
rect 21424 9848 21504 9868
rect 0 9808 2540 9848
rect 4919 9808 4928 9848
rect 4968 9808 5010 9848
rect 5050 9808 5092 9848
rect 5132 9808 5174 9848
rect 5214 9808 5256 9848
rect 5296 9808 5305 9848
rect 5347 9808 5356 9848
rect 5396 9808 6988 9848
rect 7028 9808 7037 9848
rect 8995 9808 9004 9848
rect 9044 9808 9100 9848
rect 9140 9808 9149 9848
rect 0 9788 80 9808
rect 9091 9807 9149 9808
rect 11320 9808 12748 9848
rect 12788 9808 12797 9848
rect 15715 9808 15724 9848
rect 15764 9808 15916 9848
rect 15956 9808 15965 9848
rect 20039 9808 20048 9848
rect 20088 9808 20130 9848
rect 20170 9808 20212 9848
rect 20252 9808 20294 9848
rect 20334 9808 20376 9848
rect 20416 9808 20425 9848
rect 21292 9808 21504 9848
rect 11320 9764 11360 9808
rect 12739 9807 12797 9808
rect 21424 9788 21504 9808
rect 1603 9724 1612 9764
rect 1652 9724 11360 9764
rect 14467 9724 14476 9764
rect 14516 9724 16396 9764
rect 16436 9724 16445 9764
rect 835 9680 893 9681
rect 9187 9680 9245 9681
rect 835 9640 844 9680
rect 884 9640 5740 9680
rect 5780 9640 5789 9680
rect 8899 9640 8908 9680
rect 8948 9640 9196 9680
rect 9236 9640 9245 9680
rect 835 9639 893 9640
rect 9187 9639 9245 9640
rect 9475 9680 9533 9681
rect 9475 9640 9484 9680
rect 9524 9640 12556 9680
rect 12596 9640 12605 9680
rect 13027 9640 13036 9680
rect 13076 9640 13804 9680
rect 13844 9640 13853 9680
rect 17731 9640 17740 9680
rect 17780 9640 20236 9680
rect 20276 9640 20285 9680
rect 9475 9639 9533 9640
rect 7651 9596 7709 9597
rect 2179 9556 2188 9596
rect 2228 9556 5356 9596
rect 5396 9556 5405 9596
rect 5539 9556 5548 9596
rect 5588 9556 7468 9596
rect 7508 9556 7517 9596
rect 7651 9556 7660 9596
rect 7700 9556 7756 9596
rect 7796 9556 7805 9596
rect 8035 9556 8044 9596
rect 8084 9556 8428 9596
rect 8468 9556 8477 9596
rect 9187 9556 9196 9596
rect 9236 9556 9868 9596
rect 9908 9556 9917 9596
rect 12643 9556 12652 9596
rect 12692 9556 12940 9596
rect 12980 9556 12989 9596
rect 17635 9556 17644 9596
rect 17684 9556 18028 9596
rect 18068 9556 18077 9596
rect 7651 9555 7709 9556
rect 17731 9512 17789 9513
rect 21424 9512 21504 9532
rect 2947 9472 2956 9512
rect 2996 9472 3340 9512
rect 3380 9472 3389 9512
rect 3523 9472 3532 9512
rect 3572 9472 4588 9512
rect 4628 9472 4637 9512
rect 6979 9472 6988 9512
rect 7028 9472 10348 9512
rect 10388 9472 11116 9512
rect 11156 9472 11165 9512
rect 17155 9472 17164 9512
rect 17204 9472 17548 9512
rect 17588 9472 17740 9512
rect 17780 9472 17789 9512
rect 19075 9472 19084 9512
rect 19124 9472 19852 9512
rect 19892 9472 21504 9512
rect 17731 9471 17789 9472
rect 21424 9452 21504 9472
rect 3619 9428 3677 9429
rect 4195 9428 4253 9429
rect 10531 9428 10589 9429
rect 13219 9428 13277 9429
rect 14659 9428 14717 9429
rect 2467 9388 2476 9428
rect 2516 9388 2764 9428
rect 2804 9388 2813 9428
rect 3427 9388 3436 9428
rect 3476 9388 3628 9428
rect 3668 9388 3677 9428
rect 4099 9388 4108 9428
rect 4148 9388 4204 9428
rect 4244 9388 4684 9428
rect 4724 9388 4733 9428
rect 7468 9388 10540 9428
rect 10580 9388 10589 9428
rect 12739 9388 12748 9428
rect 12788 9388 13228 9428
rect 13268 9388 13277 9428
rect 14083 9388 14092 9428
rect 14132 9388 14668 9428
rect 14708 9388 14717 9428
rect 3619 9387 3677 9388
rect 4195 9387 4253 9388
rect 0 9344 80 9364
rect 7468 9344 7508 9388
rect 10531 9387 10589 9388
rect 13219 9387 13277 9388
rect 14659 9387 14717 9388
rect 18403 9428 18461 9429
rect 18403 9388 18412 9428
rect 18452 9388 18508 9428
rect 18548 9388 18557 9428
rect 18403 9387 18461 9388
rect 10915 9344 10973 9345
rect 11779 9344 11837 9345
rect 17635 9344 17693 9345
rect 0 9304 7508 9344
rect 7555 9304 7564 9344
rect 7604 9304 8716 9344
rect 8756 9304 8765 9344
rect 10051 9304 10060 9344
rect 10100 9304 10252 9344
rect 10292 9304 10540 9344
rect 10580 9304 10589 9344
rect 10915 9304 10924 9344
rect 10964 9304 11116 9344
rect 11156 9304 11165 9344
rect 11779 9304 11788 9344
rect 11828 9304 14860 9344
rect 14900 9304 14909 9344
rect 17059 9304 17068 9344
rect 17108 9304 17452 9344
rect 17492 9304 17501 9344
rect 17550 9304 17644 9344
rect 17684 9304 17693 9344
rect 0 9284 80 9304
rect 10915 9303 10973 9304
rect 11779 9303 11837 9304
rect 17635 9303 17693 9304
rect 3139 9260 3197 9261
rect 9571 9260 9629 9261
rect 10147 9260 10205 9261
rect 3054 9220 3148 9260
rect 3188 9220 3197 9260
rect 6883 9220 6892 9260
rect 6932 9220 9100 9260
rect 9140 9220 9292 9260
rect 9332 9220 9341 9260
rect 9571 9220 9580 9260
rect 9620 9220 10156 9260
rect 10196 9220 10205 9260
rect 3139 9219 3197 9220
rect 9571 9219 9629 9220
rect 10147 9219 10205 9220
rect 10531 9260 10589 9261
rect 18595 9260 18653 9261
rect 10531 9220 10540 9260
rect 10580 9220 10636 9260
rect 10676 9220 10685 9260
rect 14947 9220 14956 9260
rect 14996 9220 15628 9260
rect 15668 9220 15677 9260
rect 17731 9220 17740 9260
rect 17780 9220 18604 9260
rect 18644 9220 18653 9260
rect 10531 9219 10589 9220
rect 18595 9219 18653 9220
rect 4579 9176 4637 9177
rect 21424 9176 21504 9196
rect 4483 9136 4492 9176
rect 4532 9136 4588 9176
rect 4628 9136 4637 9176
rect 5347 9136 5356 9176
rect 5396 9136 5932 9176
rect 5972 9136 12460 9176
rect 12500 9136 12509 9176
rect 13699 9136 13708 9176
rect 13748 9136 21504 9176
rect 4579 9135 4637 9136
rect 21424 9116 21504 9136
rect 7555 9092 7613 9093
rect 11875 9092 11933 9093
rect 3679 9052 3688 9092
rect 3728 9052 3770 9092
rect 3810 9052 3852 9092
rect 3892 9052 3934 9092
rect 3974 9052 4016 9092
rect 4056 9052 4065 9092
rect 6595 9052 6604 9092
rect 6644 9052 7180 9092
rect 7220 9052 7229 9092
rect 7459 9052 7468 9092
rect 7508 9052 7564 9092
rect 7604 9052 7613 9092
rect 8515 9052 8524 9092
rect 8564 9052 11884 9092
rect 11924 9052 11933 9092
rect 18799 9052 18808 9092
rect 18848 9052 18890 9092
rect 18930 9052 18972 9092
rect 19012 9052 19054 9092
rect 19094 9052 19136 9092
rect 19176 9052 19185 9092
rect 7555 9051 7613 9052
rect 11875 9051 11933 9052
rect 14275 9008 14333 9009
rect 1420 8968 14284 9008
rect 14324 8968 14333 9008
rect 14947 8968 14956 9008
rect 14996 8968 15340 9008
rect 15380 8968 15389 9008
rect 17251 8968 17260 9008
rect 17300 8968 18604 9008
rect 18644 8968 20044 9008
rect 20084 8968 20093 9008
rect 0 8840 80 8860
rect 1420 8840 1460 8968
rect 14275 8967 14333 8968
rect 2659 8884 2668 8924
rect 2708 8884 3532 8924
rect 3572 8884 3581 8924
rect 3811 8884 3820 8924
rect 3860 8884 11360 8924
rect 16963 8884 16972 8924
rect 17012 8884 19564 8924
rect 19604 8884 19613 8924
rect 8803 8840 8861 8841
rect 0 8800 1460 8840
rect 1795 8800 1804 8840
rect 1844 8800 3052 8840
rect 3092 8800 3101 8840
rect 8044 8800 8812 8840
rect 8852 8800 8861 8840
rect 11320 8840 11360 8884
rect 21424 8840 21504 8860
rect 11320 8800 21504 8840
rect 0 8780 80 8800
rect 4195 8756 4253 8757
rect 8044 8756 8084 8800
rect 8803 8799 8861 8800
rect 21424 8780 21504 8800
rect 4110 8716 4204 8756
rect 4244 8716 4253 8756
rect 6403 8716 6412 8756
rect 6452 8716 8044 8756
rect 8084 8716 8093 8756
rect 8227 8716 8236 8756
rect 8276 8716 9676 8756
rect 9716 8716 10540 8756
rect 10580 8716 10589 8756
rect 11779 8716 11788 8756
rect 11828 8716 19948 8756
rect 19988 8716 19997 8756
rect 4195 8715 4253 8716
rect 10051 8672 10109 8673
rect 4099 8632 4108 8672
rect 4148 8632 4492 8672
rect 4532 8632 4541 8672
rect 5347 8632 5356 8672
rect 5396 8632 10060 8672
rect 10100 8632 10109 8672
rect 10051 8631 10109 8632
rect 12259 8672 12317 8673
rect 12259 8632 12268 8672
rect 12308 8632 14764 8672
rect 14804 8632 14813 8672
rect 14947 8632 14956 8672
rect 14996 8632 15340 8672
rect 15380 8632 15389 8672
rect 17443 8632 17452 8672
rect 17492 8632 17932 8672
rect 17972 8632 19084 8672
rect 19124 8632 19133 8672
rect 12259 8631 12317 8632
rect 18307 8588 18365 8589
rect 3043 8548 3052 8588
rect 3092 8548 3340 8588
rect 3380 8548 3389 8588
rect 4003 8548 4012 8588
rect 4052 8548 6220 8588
rect 6260 8548 9292 8588
rect 9332 8548 9341 8588
rect 14179 8548 14188 8588
rect 14228 8548 14476 8588
rect 14516 8548 14525 8588
rect 15139 8548 15148 8588
rect 15188 8548 17836 8588
rect 17876 8548 17885 8588
rect 18222 8548 18316 8588
rect 18356 8548 18365 8588
rect 18307 8547 18365 8548
rect 16963 8504 17021 8505
rect 21424 8504 21504 8524
rect 2947 8464 2956 8504
rect 2996 8464 4204 8504
rect 4244 8464 4253 8504
rect 4867 8464 4876 8504
rect 4916 8464 5452 8504
rect 5492 8464 5501 8504
rect 10147 8464 10156 8504
rect 10196 8464 10444 8504
rect 10484 8464 10493 8504
rect 15043 8464 15052 8504
rect 15092 8464 15729 8504
rect 15769 8464 15778 8504
rect 16963 8464 16972 8504
rect 17012 8464 21504 8504
rect 16963 8463 17021 8464
rect 21424 8444 21504 8464
rect 7651 8380 7660 8420
rect 7700 8380 7852 8420
rect 7892 8380 10252 8420
rect 10292 8380 10301 8420
rect 13987 8380 13996 8420
rect 14036 8380 14188 8420
rect 14228 8380 15436 8420
rect 15476 8380 15485 8420
rect 0 8336 80 8356
rect 18115 8336 18173 8337
rect 0 8296 4628 8336
rect 4919 8296 4928 8336
rect 4968 8296 5010 8336
rect 5050 8296 5092 8336
rect 5132 8296 5174 8336
rect 5214 8296 5256 8336
rect 5296 8296 5305 8336
rect 11203 8296 11212 8336
rect 11252 8296 16204 8336
rect 16244 8296 16253 8336
rect 18030 8296 18124 8336
rect 18164 8296 18173 8336
rect 20039 8296 20048 8336
rect 20088 8296 20130 8336
rect 20170 8296 20212 8336
rect 20252 8296 20294 8336
rect 20334 8296 20376 8336
rect 20416 8296 20425 8336
rect 0 8276 80 8296
rect 3427 8128 3436 8168
rect 3476 8128 4396 8168
rect 4436 8128 4445 8168
rect 2947 8084 3005 8085
rect 268 8044 2956 8084
rect 2996 8044 3005 8084
rect 0 7832 80 7852
rect 268 7832 308 8044
rect 2947 8043 3005 8044
rect 1987 7960 1996 8000
rect 2036 7960 2045 8000
rect 2179 7960 2188 8000
rect 2228 7960 2668 8000
rect 2708 7960 2717 8000
rect 1996 7916 2036 7960
rect 4588 7916 4628 8296
rect 18115 8295 18173 8296
rect 18019 8212 18028 8252
rect 18068 8212 18077 8252
rect 6499 8168 6557 8169
rect 6414 8128 6508 8168
rect 6548 8128 6557 8168
rect 15523 8128 15532 8168
rect 15572 8128 16204 8168
rect 16244 8128 16253 8168
rect 6499 8127 6557 8128
rect 5539 8044 5548 8084
rect 5588 8044 8140 8084
rect 8180 8044 8189 8084
rect 18028 8000 18068 8212
rect 21424 8168 21504 8188
rect 19267 8128 19276 8168
rect 19316 8128 21504 8168
rect 21424 8108 21504 8128
rect 19075 8044 19084 8084
rect 19124 8044 19564 8084
rect 19604 8044 19613 8084
rect 4675 7960 4684 8000
rect 4724 7960 8332 8000
rect 8372 7960 8381 8000
rect 9667 7960 9676 8000
rect 9716 7960 11212 8000
rect 11252 7960 11261 8000
rect 11320 7960 11692 8000
rect 11732 7960 13900 8000
rect 13940 7960 13949 8000
rect 15523 7960 15532 8000
rect 15572 7960 15916 8000
rect 15956 7960 15965 8000
rect 17635 7960 17644 8000
rect 17684 7960 18508 8000
rect 18548 7960 18557 8000
rect 19363 7960 19372 8000
rect 19412 7960 20524 8000
rect 20564 7960 20573 8000
rect 8332 7916 8372 7960
rect 11320 7916 11360 7960
rect 1996 7876 2860 7916
rect 2900 7876 4204 7916
rect 4244 7876 4253 7916
rect 4588 7876 5780 7916
rect 8332 7876 11360 7916
rect 3427 7832 3485 7833
rect 0 7792 308 7832
rect 1315 7792 1324 7832
rect 1364 7792 1996 7832
rect 2036 7792 2045 7832
rect 3427 7792 3436 7832
rect 3476 7792 3724 7832
rect 3764 7792 3773 7832
rect 0 7772 80 7792
rect 3427 7791 3485 7792
rect 2755 7708 2764 7748
rect 2804 7708 4108 7748
rect 4148 7708 5644 7748
rect 5684 7708 5693 7748
rect 5740 7664 5780 7876
rect 7459 7832 7517 7833
rect 16195 7832 16253 7833
rect 21424 7832 21504 7852
rect 6115 7792 6124 7832
rect 6164 7792 6412 7832
rect 6452 7792 6461 7832
rect 7459 7792 7468 7832
rect 7508 7792 10732 7832
rect 10772 7792 10781 7832
rect 11395 7792 11404 7832
rect 11444 7792 12460 7832
rect 12500 7792 12940 7832
rect 12980 7792 13900 7832
rect 13940 7792 14284 7832
rect 14324 7792 14333 7832
rect 16195 7792 16204 7832
rect 16244 7792 16876 7832
rect 16916 7792 16925 7832
rect 21379 7792 21388 7832
rect 21428 7792 21504 7832
rect 7459 7791 7517 7792
rect 16195 7791 16253 7792
rect 21424 7772 21504 7792
rect 10435 7748 10493 7749
rect 16771 7748 16829 7749
rect 6499 7708 6508 7748
rect 6548 7708 7468 7748
rect 7508 7708 7517 7748
rect 10051 7708 10060 7748
rect 10100 7708 10444 7748
rect 10484 7708 10636 7748
rect 10676 7708 10685 7748
rect 11299 7708 11308 7748
rect 11348 7708 16780 7748
rect 16820 7708 16829 7748
rect 10435 7707 10493 7708
rect 16771 7707 16829 7708
rect 16963 7748 17021 7749
rect 19075 7748 19133 7749
rect 16963 7708 16972 7748
rect 17012 7708 17106 7748
rect 18990 7708 19084 7748
rect 19124 7708 19133 7748
rect 16963 7707 17021 7708
rect 19075 7707 19133 7708
rect 17059 7664 17117 7665
rect 3427 7624 3436 7664
rect 3476 7624 4916 7664
rect 5740 7624 14092 7664
rect 14132 7624 14141 7664
rect 15715 7624 15724 7664
rect 15764 7624 15916 7664
rect 15956 7624 15965 7664
rect 16291 7624 16300 7664
rect 16340 7624 17068 7664
rect 17108 7624 17117 7664
rect 4771 7580 4829 7581
rect 2563 7540 2572 7580
rect 2612 7540 2652 7580
rect 3679 7540 3688 7580
rect 3728 7540 3770 7580
rect 3810 7540 3852 7580
rect 3892 7540 3934 7580
rect 3974 7540 4016 7580
rect 4056 7540 4065 7580
rect 4686 7540 4780 7580
rect 4820 7540 4829 7580
rect 4876 7580 4916 7624
rect 17059 7623 17117 7624
rect 4876 7540 6508 7580
rect 6548 7540 6557 7580
rect 6883 7540 6892 7580
rect 6932 7540 8236 7580
rect 8276 7540 8285 7580
rect 8611 7540 8620 7580
rect 8660 7540 9196 7580
rect 9236 7540 9245 7580
rect 10723 7540 10732 7580
rect 10772 7540 11308 7580
rect 11348 7540 16684 7580
rect 16724 7540 16733 7580
rect 18799 7540 18808 7580
rect 18848 7540 18890 7580
rect 18930 7540 18972 7580
rect 19012 7540 19054 7580
rect 19094 7540 19136 7580
rect 19176 7540 19185 7580
rect 2572 7496 2612 7540
rect 4771 7539 4829 7540
rect 21424 7496 21504 7516
rect 2083 7456 2092 7496
rect 2132 7456 4396 7496
rect 4436 7456 4445 7496
rect 6403 7456 6412 7496
rect 6452 7456 7756 7496
rect 7796 7456 9964 7496
rect 10004 7456 10013 7496
rect 12547 7456 12556 7496
rect 12596 7456 21504 7496
rect 21424 7436 21504 7456
rect 1315 7412 1373 7413
rect 1315 7372 1324 7412
rect 1364 7372 2572 7412
rect 2612 7372 2621 7412
rect 4579 7372 4588 7412
rect 4628 7372 9388 7412
rect 9428 7372 9437 7412
rect 11203 7372 11212 7412
rect 11252 7372 11404 7412
rect 11444 7372 11453 7412
rect 13987 7372 13996 7412
rect 14036 7372 18316 7412
rect 18356 7372 18365 7412
rect 1315 7371 1373 7372
rect 0 7328 80 7348
rect 4588 7328 4628 7372
rect 0 7288 652 7328
rect 692 7288 701 7328
rect 2500 7288 4628 7328
rect 14083 7288 14092 7328
rect 14132 7288 14476 7328
rect 14516 7288 14525 7328
rect 0 7268 80 7288
rect 2500 7244 2540 7288
rect 1315 7204 1324 7244
rect 1364 7204 2540 7244
rect 4291 7204 4300 7244
rect 4340 7204 7180 7244
rect 7220 7204 7229 7244
rect 9955 7204 9964 7244
rect 10004 7204 14324 7244
rect 14284 7160 14324 7204
rect 16387 7160 16445 7161
rect 21424 7160 21504 7180
rect 2467 7120 2476 7160
rect 2516 7120 3052 7160
rect 3092 7120 3101 7160
rect 3427 7120 3436 7160
rect 3476 7120 8332 7160
rect 8372 7120 8524 7160
rect 8564 7120 8573 7160
rect 12163 7120 12172 7160
rect 12212 7120 13420 7160
rect 13460 7120 13940 7160
rect 14275 7120 14284 7160
rect 14324 7120 14333 7160
rect 16387 7120 16396 7160
rect 16436 7120 21504 7160
rect 3331 7076 3389 7077
rect 3715 7076 3773 7077
rect 1315 7036 1324 7076
rect 1364 7036 3340 7076
rect 3380 7036 3724 7076
rect 3764 7036 3773 7076
rect 5923 7036 5932 7076
rect 5972 7036 7660 7076
rect 7700 7036 12460 7076
rect 12500 7036 12509 7076
rect 3331 7035 3389 7036
rect 3715 7035 3773 7036
rect 13411 6992 13469 6993
rect 1795 6952 1804 6992
rect 1844 6952 4780 6992
rect 4820 6952 4829 6992
rect 9763 6952 9772 6992
rect 9812 6952 10252 6992
rect 10292 6952 10301 6992
rect 13326 6952 13420 6992
rect 13460 6952 13469 6992
rect 13900 6992 13940 7120
rect 16387 7119 16445 7120
rect 21424 7100 21504 7120
rect 13987 7036 13996 7076
rect 14036 7036 16396 7076
rect 16436 7036 16445 7076
rect 17155 6992 17213 6993
rect 13900 6952 17164 6992
rect 17204 6952 20620 6992
rect 20660 6952 20669 6992
rect 13411 6951 13469 6952
rect 17155 6951 17213 6952
rect 2659 6908 2717 6909
rect 10243 6908 10301 6909
rect 2659 6868 2668 6908
rect 2708 6868 10252 6908
rect 10292 6868 10301 6908
rect 2659 6867 2717 6868
rect 10243 6867 10301 6868
rect 13219 6908 13277 6909
rect 13219 6868 13228 6908
rect 13268 6868 13612 6908
rect 13652 6868 13661 6908
rect 13219 6867 13277 6868
rect 0 6824 80 6844
rect 11395 6824 11453 6825
rect 21424 6824 21504 6844
rect 0 6784 2540 6824
rect 4919 6784 4928 6824
rect 4968 6784 5010 6824
rect 5050 6784 5092 6824
rect 5132 6784 5174 6824
rect 5214 6784 5256 6824
rect 5296 6784 5305 6824
rect 6211 6784 6220 6824
rect 6260 6784 8140 6824
rect 8180 6784 11404 6824
rect 11444 6784 11453 6824
rect 13795 6784 13804 6824
rect 13844 6784 18932 6824
rect 20039 6784 20048 6824
rect 20088 6784 20130 6824
rect 20170 6784 20212 6824
rect 20252 6784 20294 6824
rect 20334 6784 20376 6824
rect 20416 6784 20425 6824
rect 20812 6784 21504 6824
rect 0 6764 80 6784
rect 2500 6740 2540 6784
rect 11395 6783 11453 6784
rect 17443 6740 17501 6741
rect 2500 6700 15820 6740
rect 15860 6700 15869 6740
rect 17443 6700 17452 6740
rect 17492 6700 18412 6740
rect 18452 6700 18461 6740
rect 17443 6699 17501 6700
rect 3715 6656 3773 6657
rect 18892 6656 18932 6784
rect 20812 6740 20852 6784
rect 21424 6764 21504 6784
rect 18979 6700 18988 6740
rect 19028 6700 20852 6740
rect 2659 6616 2668 6656
rect 2708 6616 3532 6656
rect 3572 6616 3581 6656
rect 3715 6616 3724 6656
rect 3764 6616 7124 6656
rect 7171 6616 7180 6656
rect 7220 6616 11404 6656
rect 11444 6616 11453 6656
rect 11779 6616 11788 6656
rect 11828 6616 18796 6656
rect 18836 6616 18845 6656
rect 18892 6616 20180 6656
rect 3715 6615 3773 6616
rect 7084 6572 7124 6616
rect 1507 6532 1516 6572
rect 1556 6532 3436 6572
rect 3476 6532 3485 6572
rect 7084 6532 11116 6572
rect 11156 6532 11165 6572
rect 12259 6532 12268 6572
rect 12308 6532 18892 6572
rect 18932 6532 18941 6572
rect 5635 6488 5693 6489
rect 20140 6488 20180 6616
rect 21424 6488 21504 6508
rect 2371 6448 2380 6488
rect 2420 6448 3148 6488
rect 3188 6448 3197 6488
rect 5550 6448 5644 6488
rect 5684 6448 5693 6488
rect 5923 6448 5932 6488
rect 5972 6448 9772 6488
rect 9812 6448 9821 6488
rect 13411 6448 13420 6488
rect 13460 6448 13804 6488
rect 13844 6448 13853 6488
rect 15907 6448 15916 6488
rect 15956 6448 17068 6488
rect 17108 6448 17117 6488
rect 17827 6448 17836 6488
rect 17876 6448 19852 6488
rect 19892 6448 19901 6488
rect 20140 6448 21504 6488
rect 5635 6447 5693 6448
rect 21424 6428 21504 6448
rect 3052 6364 5260 6404
rect 5300 6364 5309 6404
rect 17923 6364 17932 6404
rect 17972 6364 18700 6404
rect 18740 6364 18988 6404
rect 19028 6364 19037 6404
rect 0 6320 80 6340
rect 3052 6320 3092 6364
rect 0 6280 500 6320
rect 2563 6280 2572 6320
rect 2612 6280 3052 6320
rect 3092 6280 3101 6320
rect 3235 6280 3244 6320
rect 3284 6280 4588 6320
rect 4628 6280 4637 6320
rect 6595 6280 6604 6320
rect 6644 6280 7084 6320
rect 7124 6280 7133 6320
rect 15619 6280 15628 6320
rect 15668 6280 16876 6320
rect 16916 6280 16925 6320
rect 18019 6280 18028 6320
rect 18068 6280 20236 6320
rect 20276 6280 20285 6320
rect 0 6260 80 6280
rect 460 6236 500 6280
rect 2659 6236 2717 6237
rect 17923 6236 17981 6237
rect 460 6196 2668 6236
rect 2708 6196 2717 6236
rect 4099 6196 4108 6236
rect 4148 6196 4300 6236
rect 4340 6196 4349 6236
rect 4675 6196 4684 6236
rect 4724 6196 5452 6236
rect 5492 6196 6316 6236
rect 6356 6196 6365 6236
rect 6979 6196 6988 6236
rect 7028 6196 15148 6236
rect 15188 6196 15197 6236
rect 15427 6196 15436 6236
rect 15476 6196 16204 6236
rect 16244 6196 16253 6236
rect 16579 6196 16588 6236
rect 16628 6196 17068 6236
rect 17108 6196 17117 6236
rect 17731 6196 17740 6236
rect 17780 6196 17932 6236
rect 17972 6196 17981 6236
rect 18883 6196 18892 6236
rect 18932 6196 19660 6236
rect 19700 6196 19709 6236
rect 2659 6195 2717 6196
rect 17923 6195 17981 6196
rect 18499 6152 18557 6153
rect 21424 6152 21504 6172
rect 1612 6112 5836 6152
rect 5876 6112 5885 6152
rect 6883 6112 6892 6152
rect 6932 6112 9580 6152
rect 9620 6112 9629 6152
rect 13324 6112 18508 6152
rect 18548 6112 18557 6152
rect 67 6028 76 6068
rect 116 6028 1516 6068
rect 1556 6028 1565 6068
rect 0 5816 80 5836
rect 1612 5816 1652 6112
rect 12259 6068 12317 6069
rect 3679 6028 3688 6068
rect 3728 6028 3770 6068
rect 3810 6028 3852 6068
rect 3892 6028 3934 6068
rect 3974 6028 4016 6068
rect 4056 6028 4065 6068
rect 6892 6028 12268 6068
rect 12308 6028 12317 6068
rect 6892 5984 6932 6028
rect 12259 6027 12317 6028
rect 13324 5984 13364 6112
rect 18499 6111 18557 6112
rect 20140 6112 21504 6152
rect 18307 6068 18365 6069
rect 15139 6028 15148 6068
rect 15188 6028 18316 6068
rect 18356 6028 18365 6068
rect 18799 6028 18808 6068
rect 18848 6028 18890 6068
rect 18930 6028 18972 6068
rect 19012 6028 19054 6068
rect 19094 6028 19136 6068
rect 19176 6028 19185 6068
rect 18307 6027 18365 6028
rect 17635 5984 17693 5985
rect 18403 5984 18461 5985
rect 2083 5944 2092 5984
rect 2132 5944 6932 5984
rect 9187 5944 9196 5984
rect 9236 5944 13364 5984
rect 13411 5944 13420 5984
rect 13460 5944 13612 5984
rect 13652 5944 16396 5984
rect 16436 5944 17644 5984
rect 17684 5944 17693 5984
rect 18019 5944 18028 5984
rect 18068 5944 18412 5984
rect 18452 5944 18461 5984
rect 17635 5943 17693 5944
rect 18403 5943 18461 5944
rect 20140 5900 20180 6112
rect 21424 6092 21504 6112
rect 3331 5860 3340 5900
rect 3380 5860 3724 5900
rect 3764 5860 6892 5900
rect 6932 5860 6941 5900
rect 7075 5860 7084 5900
rect 7124 5860 9332 5900
rect 9571 5860 9580 5900
rect 9620 5860 20180 5900
rect 4771 5816 4829 5817
rect 9292 5816 9332 5860
rect 15619 5816 15677 5817
rect 21424 5816 21504 5836
rect 0 5776 1652 5816
rect 3139 5776 3148 5816
rect 3188 5776 4780 5816
rect 4820 5776 9196 5816
rect 9236 5776 9245 5816
rect 9292 5776 13228 5816
rect 13268 5776 13277 5816
rect 15534 5776 15628 5816
rect 15668 5776 15677 5816
rect 17635 5776 17644 5816
rect 17684 5776 18412 5816
rect 18452 5776 18461 5816
rect 20140 5776 21504 5816
rect 0 5756 80 5776
rect 4771 5775 4829 5776
rect 15619 5775 15677 5776
rect 3427 5732 3485 5733
rect 4675 5732 4733 5733
rect 3427 5692 3436 5732
rect 3476 5692 3628 5732
rect 3668 5692 3677 5732
rect 4675 5692 4684 5732
rect 4724 5692 9292 5732
rect 9332 5692 9341 5732
rect 13027 5692 13036 5732
rect 13076 5692 13420 5732
rect 13460 5692 13469 5732
rect 14947 5692 14956 5732
rect 14996 5692 16300 5732
rect 16340 5692 16349 5732
rect 16675 5692 16684 5732
rect 16724 5692 17356 5732
rect 17396 5692 17972 5732
rect 3427 5691 3485 5692
rect 4675 5691 4733 5692
rect 2755 5608 2764 5648
rect 2804 5608 4780 5648
rect 4820 5608 4829 5648
rect 5155 5608 5164 5648
rect 5204 5608 6988 5648
rect 7028 5608 7037 5648
rect 8227 5608 8236 5648
rect 8276 5608 8524 5648
rect 8564 5608 8573 5648
rect 15619 5608 15628 5648
rect 15668 5608 16972 5648
rect 17012 5608 17021 5648
rect 17251 5608 17260 5648
rect 17300 5608 17644 5648
rect 17684 5608 17693 5648
rect 17932 5564 17972 5692
rect 20140 5564 20180 5776
rect 21424 5756 21504 5776
rect 4099 5524 4108 5564
rect 4148 5524 7468 5564
rect 7508 5524 7517 5564
rect 13699 5524 13708 5564
rect 13748 5524 16300 5564
rect 16340 5524 16349 5564
rect 17923 5524 17932 5564
rect 17972 5524 17981 5564
rect 18412 5524 20180 5564
rect 1891 5440 1900 5480
rect 1940 5440 2476 5480
rect 2516 5440 2525 5480
rect 3139 5440 3148 5480
rect 3188 5440 8908 5480
rect 8948 5440 8957 5480
rect 13219 5440 13228 5480
rect 13268 5440 18316 5480
rect 18356 5440 18365 5480
rect 7075 5396 7133 5397
rect 18412 5396 18452 5524
rect 21424 5480 21504 5500
rect 19651 5440 19660 5480
rect 19700 5440 21504 5480
rect 21424 5420 21504 5440
rect 4387 5356 4396 5396
rect 4436 5356 4684 5396
rect 4724 5356 5932 5396
rect 5972 5356 5981 5396
rect 6307 5356 6316 5396
rect 6356 5356 6796 5396
rect 6836 5356 6845 5396
rect 7075 5356 7084 5396
rect 7124 5356 18452 5396
rect 7075 5355 7133 5356
rect 0 5312 80 5332
rect 0 5272 2540 5312
rect 4919 5272 4928 5312
rect 4968 5272 5010 5312
rect 5050 5272 5092 5312
rect 5132 5272 5174 5312
rect 5214 5272 5256 5312
rect 5296 5272 5305 5312
rect 6595 5272 6604 5312
rect 6644 5272 7180 5312
rect 7220 5272 7229 5312
rect 8803 5272 8812 5312
rect 8852 5272 9292 5312
rect 9332 5272 9341 5312
rect 15235 5272 15244 5312
rect 15284 5272 15628 5312
rect 15668 5272 16684 5312
rect 16724 5272 16733 5312
rect 20039 5272 20048 5312
rect 20088 5272 20130 5312
rect 20170 5272 20212 5312
rect 20252 5272 20294 5312
rect 20334 5272 20376 5312
rect 20416 5272 20425 5312
rect 0 5252 80 5272
rect 2500 5228 2540 5272
rect 2500 5188 7756 5228
rect 7796 5188 7805 5228
rect 8812 5144 8852 5272
rect 12643 5228 12701 5229
rect 12643 5188 12652 5228
rect 12692 5188 15532 5228
rect 15572 5188 15581 5228
rect 16483 5188 16492 5228
rect 16532 5188 16780 5228
rect 16820 5188 16829 5228
rect 12643 5187 12701 5188
rect 12547 5144 12605 5145
rect 21424 5144 21504 5164
rect 4291 5104 4300 5144
rect 4340 5104 8852 5144
rect 12355 5104 12364 5144
rect 12404 5104 12556 5144
rect 12596 5104 21504 5144
rect 12547 5103 12605 5104
rect 21424 5084 21504 5104
rect 4675 5060 4733 5061
rect 16579 5060 16637 5061
rect 2275 5020 2284 5060
rect 2324 5020 3340 5060
rect 3380 5020 3389 5060
rect 4195 5020 4204 5060
rect 4244 5020 4284 5060
rect 4675 5020 4684 5060
rect 4724 5020 4780 5060
rect 4820 5020 4829 5060
rect 12451 5020 12460 5060
rect 12500 5020 12652 5060
rect 12692 5020 14572 5060
rect 14612 5020 15188 5060
rect 4204 4976 4244 5020
rect 4675 5019 4733 5020
rect 6787 4976 6845 4977
rect 7171 4976 7229 4977
rect 2846 4936 2855 4976
rect 2895 4936 2904 4976
rect 2947 4936 2956 4976
rect 2996 4936 4492 4976
rect 4532 4936 4541 4976
rect 6787 4936 6796 4976
rect 6836 4936 7180 4976
rect 7220 4936 7229 4976
rect 8995 4936 9004 4976
rect 9044 4936 11404 4976
rect 11444 4936 11453 4976
rect 2860 4893 2900 4936
rect 6787 4935 6845 4936
rect 7171 4935 7229 4936
rect 2851 4892 2909 4893
rect 12460 4892 12500 5020
rect 13507 4976 13565 4977
rect 13795 4976 13853 4977
rect 15148 4976 15188 5020
rect 16579 5020 16588 5060
rect 16628 5020 17644 5060
rect 17684 5020 17693 5060
rect 16579 5019 16637 5020
rect 17443 4976 17501 4977
rect 17731 4976 17789 4977
rect 13507 4936 13516 4976
rect 13556 4936 13804 4976
rect 13844 4936 15052 4976
rect 15092 4936 15101 4976
rect 15148 4936 15436 4976
rect 15476 4936 16300 4976
rect 16340 4936 16349 4976
rect 17059 4936 17068 4976
rect 17108 4936 17452 4976
rect 17492 4936 17501 4976
rect 17646 4936 17740 4976
rect 17780 4936 17789 4976
rect 17923 4936 17932 4976
rect 17972 4936 19084 4976
rect 19124 4936 19133 4976
rect 19459 4936 19468 4976
rect 19508 4936 20236 4976
rect 20276 4936 20285 4976
rect 13507 4935 13565 4936
rect 13795 4935 13853 4936
rect 17068 4892 17108 4936
rect 17443 4935 17501 4936
rect 17731 4935 17789 4936
rect 18019 4892 18077 4893
rect 2851 4852 2860 4892
rect 2900 4852 2909 4892
rect 4387 4852 4396 4892
rect 4436 4852 7372 4892
rect 7412 4852 7421 4892
rect 7651 4852 7660 4892
rect 7700 4852 8660 4892
rect 11011 4852 11020 4892
rect 11060 4852 12500 4892
rect 13027 4852 13036 4892
rect 13076 4852 13228 4892
rect 13268 4852 17108 4892
rect 17155 4852 17164 4892
rect 17204 4852 18028 4892
rect 18068 4852 18077 4892
rect 2851 4851 2909 4852
rect 0 4808 80 4828
rect 1219 4808 1277 4809
rect 8620 4808 8660 4852
rect 18019 4851 18077 4852
rect 21424 4808 21504 4828
rect 0 4768 1228 4808
rect 1268 4768 1277 4808
rect 2179 4768 2188 4808
rect 2228 4768 2668 4808
rect 2708 4768 2717 4808
rect 2851 4768 2860 4808
rect 2900 4768 3148 4808
rect 3188 4768 3197 4808
rect 4099 4768 4108 4808
rect 4148 4768 6508 4808
rect 6548 4768 8524 4808
rect 8564 4768 8573 4808
rect 8620 4768 9100 4808
rect 9140 4768 21504 4808
rect 0 4748 80 4768
rect 1219 4767 1277 4768
rect 21424 4748 21504 4768
rect 5539 4724 5597 4725
rect 1315 4684 1324 4724
rect 1364 4684 5548 4724
rect 5588 4684 5597 4724
rect 6691 4684 6700 4724
rect 6740 4684 7084 4724
rect 7124 4684 7133 4724
rect 7363 4684 7372 4724
rect 7412 4684 10252 4724
rect 10292 4684 10301 4724
rect 11971 4684 11980 4724
rect 12020 4684 13228 4724
rect 13268 4684 13277 4724
rect 14947 4684 14956 4724
rect 14996 4684 17932 4724
rect 17972 4684 17981 4724
rect 18595 4684 18604 4724
rect 18644 4684 19948 4724
rect 19988 4684 19997 4724
rect 5539 4683 5597 4684
rect 1987 4600 1996 4640
rect 2036 4600 5260 4640
rect 5300 4600 5309 4640
rect 16195 4600 16204 4640
rect 16244 4600 17356 4640
rect 17396 4600 18412 4640
rect 18452 4600 18461 4640
rect 19363 4556 19421 4557
rect 3679 4516 3688 4556
rect 3728 4516 3770 4556
rect 3810 4516 3852 4556
rect 3892 4516 3934 4556
rect 3974 4516 4016 4556
rect 4056 4516 4065 4556
rect 18799 4516 18808 4556
rect 18848 4516 18890 4556
rect 18930 4516 18972 4556
rect 19012 4516 19054 4556
rect 19094 4516 19136 4556
rect 19176 4516 19185 4556
rect 19363 4516 19372 4556
rect 19412 4516 19506 4556
rect 19363 4515 19421 4516
rect 2851 4472 2909 4473
rect 7459 4472 7517 4473
rect 11587 4472 11645 4473
rect 2851 4432 2860 4472
rect 2900 4432 7316 4472
rect 2851 4431 2909 4432
rect 7276 4388 7316 4432
rect 7459 4432 7468 4472
rect 7508 4432 7602 4472
rect 7939 4432 7948 4472
rect 7988 4432 11596 4472
rect 11636 4432 11645 4472
rect 7459 4431 7517 4432
rect 11587 4431 11645 4432
rect 17635 4472 17693 4473
rect 21424 4472 21504 4492
rect 17635 4432 17644 4472
rect 17684 4432 21504 4472
rect 17635 4431 17693 4432
rect 21424 4412 21504 4432
rect 19363 4388 19421 4389
rect 2500 4348 7220 4388
rect 7276 4348 14668 4388
rect 14708 4348 14717 4388
rect 15907 4348 15916 4388
rect 15956 4348 16300 4388
rect 16340 4348 16349 4388
rect 18787 4348 18796 4388
rect 18836 4348 19372 4388
rect 19412 4348 19421 4388
rect 0 4304 80 4324
rect 2500 4304 2540 4348
rect 0 4264 364 4304
rect 404 4264 413 4304
rect 1315 4264 1324 4304
rect 1364 4264 2540 4304
rect 0 4244 80 4264
rect 2860 3968 2900 4348
rect 4483 4304 4541 4305
rect 3523 4264 3532 4304
rect 3572 4264 4492 4304
rect 4532 4264 4972 4304
rect 5012 4264 5452 4304
rect 5492 4264 5501 4304
rect 5548 4264 6508 4304
rect 6548 4264 6557 4304
rect 4483 4263 4541 4264
rect 5548 4220 5588 4264
rect 5923 4220 5981 4221
rect 3235 4180 3244 4220
rect 3284 4180 4108 4220
rect 4148 4180 4157 4220
rect 4579 4180 4588 4220
rect 4628 4180 5588 4220
rect 5827 4180 5836 4220
rect 5876 4180 5932 4220
rect 5972 4180 5981 4220
rect 7180 4220 7220 4348
rect 19363 4347 19421 4348
rect 16675 4304 16733 4305
rect 7267 4264 7276 4304
rect 7316 4264 8660 4304
rect 9859 4264 9868 4304
rect 9908 4264 10060 4304
rect 10100 4264 10252 4304
rect 10292 4264 10301 4304
rect 16590 4264 16684 4304
rect 16724 4264 16733 4304
rect 8620 4220 8660 4264
rect 16675 4263 16733 4264
rect 7180 4180 8084 4220
rect 8611 4180 8620 4220
rect 8660 4180 8669 4220
rect 8716 4180 10636 4220
rect 10676 4180 10685 4220
rect 19075 4180 19084 4220
rect 19124 4180 19660 4220
rect 19700 4180 19709 4220
rect 5923 4179 5981 4180
rect 5731 4136 5789 4137
rect 8044 4136 8084 4180
rect 8716 4136 8756 4180
rect 21424 4141 21504 4156
rect 16579 4136 16637 4137
rect 16963 4136 17021 4137
rect 3139 4096 3148 4136
rect 3188 4096 4492 4136
rect 4532 4096 4541 4136
rect 4588 4096 5740 4136
rect 5780 4096 5789 4136
rect 6403 4096 6412 4136
rect 6452 4096 7948 4136
rect 7988 4096 7997 4136
rect 8044 4096 8756 4136
rect 8899 4096 8908 4136
rect 8948 4096 11980 4136
rect 12020 4096 12268 4136
rect 12308 4096 12317 4136
rect 15139 4096 15148 4136
rect 15188 4096 15916 4136
rect 15956 4096 16588 4136
rect 16628 4096 16684 4136
rect 16724 4096 16733 4136
rect 16878 4096 16972 4136
rect 17012 4096 17021 4136
rect 2659 3928 2668 3968
rect 2708 3928 2717 3968
rect 2851 3928 2860 3968
rect 2900 3928 2909 3968
rect 2668 3884 2708 3928
rect 2668 3844 2956 3884
rect 2996 3844 3005 3884
rect 0 3800 80 3820
rect 4588 3800 4628 4096
rect 5731 4095 5789 4096
rect 16579 4095 16637 4096
rect 16963 4095 17021 4096
rect 17155 4136 17213 4137
rect 17155 4096 17164 4136
rect 17204 4096 17260 4136
rect 17300 4096 17309 4136
rect 17731 4096 17740 4136
rect 17780 4096 18124 4136
rect 18164 4096 19564 4136
rect 19604 4096 19613 4136
rect 21292 4101 21504 4141
rect 17155 4095 17213 4096
rect 17260 4052 17300 4096
rect 4771 4012 4780 4052
rect 4820 4012 5356 4052
rect 5396 4012 5405 4052
rect 7075 4012 7084 4052
rect 7124 4012 12460 4052
rect 12500 4012 12509 4052
rect 17260 4012 19468 4052
rect 19508 4012 19517 4052
rect 21292 3968 21332 4101
rect 21388 4096 21504 4101
rect 21424 4076 21504 4096
rect 5232 3928 5260 3968
rect 5300 3928 9004 3968
rect 9044 3928 9053 3968
rect 9571 3928 9580 3968
rect 9620 3928 13132 3968
rect 13172 3928 13181 3968
rect 13699 3928 13708 3968
rect 13748 3928 18028 3968
rect 18068 3928 21332 3968
rect 5356 3884 5396 3928
rect 5347 3844 5356 3884
rect 5396 3844 5405 3884
rect 7564 3844 7660 3884
rect 7700 3844 7709 3884
rect 8515 3844 8524 3884
rect 8564 3844 10060 3884
rect 10100 3844 10109 3884
rect 10627 3844 10636 3884
rect 10676 3844 12844 3884
rect 12884 3844 12893 3884
rect 13411 3844 13420 3884
rect 13460 3844 20852 3884
rect 7564 3800 7604 3844
rect 0 3760 4628 3800
rect 4919 3760 4928 3800
rect 4968 3760 5010 3800
rect 5050 3760 5092 3800
rect 5132 3760 5174 3800
rect 5214 3760 5256 3800
rect 5296 3760 5305 3800
rect 6115 3760 6124 3800
rect 6164 3760 7604 3800
rect 7651 3800 7709 3801
rect 16579 3800 16637 3801
rect 18307 3800 18365 3801
rect 20812 3800 20852 3844
rect 21424 3800 21504 3820
rect 7651 3760 7660 3800
rect 7700 3760 8812 3800
rect 8852 3760 8861 3800
rect 10339 3760 10348 3800
rect 10388 3760 11020 3800
rect 11060 3760 11069 3800
rect 15427 3760 15436 3800
rect 15476 3760 15724 3800
rect 15764 3760 15773 3800
rect 16579 3760 16588 3800
rect 16628 3760 18316 3800
rect 18356 3760 18365 3800
rect 20039 3760 20048 3800
rect 20088 3760 20130 3800
rect 20170 3760 20212 3800
rect 20252 3760 20294 3800
rect 20334 3760 20376 3800
rect 20416 3760 20425 3800
rect 20812 3760 21504 3800
rect 0 3740 80 3760
rect 7651 3759 7709 3760
rect 16579 3759 16637 3760
rect 18307 3759 18365 3760
rect 21424 3740 21504 3760
rect 6883 3716 6941 3717
rect 1987 3676 1996 3716
rect 2036 3676 6892 3716
rect 6932 3676 6941 3716
rect 6883 3675 6941 3676
rect 7267 3716 7325 3717
rect 7267 3676 7276 3716
rect 7316 3676 15340 3716
rect 15380 3676 15389 3716
rect 16195 3676 16204 3716
rect 16244 3676 16876 3716
rect 16916 3676 16925 3716
rect 17059 3676 17068 3716
rect 17108 3676 17356 3716
rect 17396 3676 17405 3716
rect 7267 3675 7325 3676
rect 8515 3632 8573 3633
rect 13315 3632 13373 3633
rect 3139 3592 3148 3632
rect 3188 3592 4684 3632
rect 4724 3592 4733 3632
rect 5059 3592 5068 3632
rect 5108 3592 7660 3632
rect 7700 3592 7709 3632
rect 8419 3592 8428 3632
rect 8468 3592 8524 3632
rect 8564 3592 8573 3632
rect 9955 3592 9964 3632
rect 10004 3592 10444 3632
rect 10484 3592 10493 3632
rect 13315 3592 13324 3632
rect 13364 3592 18028 3632
rect 18068 3592 18077 3632
rect 8515 3591 8573 3592
rect 13315 3591 13373 3592
rect 67 3548 125 3549
rect 7267 3548 7325 3549
rect 7555 3548 7613 3549
rect 8995 3548 9053 3549
rect 67 3508 76 3548
rect 116 3508 4588 3548
rect 4628 3508 4637 3548
rect 6499 3508 6508 3548
rect 6548 3508 7276 3548
rect 7316 3508 7325 3548
rect 7470 3508 7564 3548
rect 7604 3508 7613 3548
rect 7843 3508 7852 3548
rect 7892 3508 8140 3548
rect 8180 3508 8189 3548
rect 8910 3508 9004 3548
rect 9044 3508 9053 3548
rect 9283 3508 9292 3548
rect 9332 3508 10924 3548
rect 10964 3508 10973 3548
rect 11107 3508 11116 3548
rect 11156 3508 18412 3548
rect 18452 3508 18461 3548
rect 67 3507 125 3508
rect 7267 3507 7325 3508
rect 7555 3507 7613 3508
rect 8995 3507 9053 3508
rect 4195 3464 4253 3465
rect 7075 3464 7133 3465
rect 18211 3464 18269 3465
rect 21424 3464 21504 3484
rect 3619 3424 3628 3464
rect 3668 3424 4204 3464
rect 4244 3424 6220 3464
rect 6260 3424 6269 3464
rect 7075 3424 7084 3464
rect 7124 3424 7180 3464
rect 7220 3424 7229 3464
rect 8035 3424 8044 3464
rect 8084 3424 11404 3464
rect 11444 3424 12364 3464
rect 12404 3424 12413 3464
rect 12835 3424 12844 3464
rect 12884 3424 14188 3464
rect 14228 3424 14237 3464
rect 16963 3424 16972 3464
rect 17012 3424 17644 3464
rect 17684 3424 17693 3464
rect 18115 3424 18124 3464
rect 18164 3424 18220 3464
rect 18260 3424 18269 3464
rect 4195 3423 4253 3424
rect 7075 3423 7133 3424
rect 18211 3423 18269 3424
rect 20140 3424 21504 3464
rect 3907 3380 3965 3381
rect 17635 3380 17693 3381
rect 3715 3340 3724 3380
rect 3764 3340 3916 3380
rect 3956 3340 3965 3380
rect 8419 3340 8428 3380
rect 8468 3340 8716 3380
rect 8756 3340 9484 3380
rect 9524 3340 9533 3380
rect 11320 3340 17644 3380
rect 17684 3340 17693 3380
rect 3907 3339 3965 3340
rect 0 3296 80 3316
rect 0 3256 268 3296
rect 308 3256 317 3296
rect 4867 3256 4876 3296
rect 4916 3256 6988 3296
rect 7028 3256 7037 3296
rect 7747 3256 7756 3296
rect 7796 3256 8812 3296
rect 8852 3256 8861 3296
rect 0 3236 80 3256
rect 11320 3212 11360 3340
rect 17635 3339 17693 3340
rect 18019 3296 18077 3297
rect 1411 3172 1420 3212
rect 1460 3172 2188 3212
rect 2228 3172 2237 3212
rect 6211 3172 6220 3212
rect 6260 3172 11360 3212
rect 11884 3256 15956 3296
rect 16291 3256 16300 3296
rect 16340 3256 16780 3296
rect 16820 3256 16829 3296
rect 17347 3256 17356 3296
rect 17396 3256 18028 3296
rect 18068 3256 19660 3296
rect 19700 3256 19709 3296
rect 1603 3088 1612 3128
rect 1652 3088 2284 3128
rect 2324 3088 2333 3128
rect 8611 3088 8620 3128
rect 8660 3088 9100 3128
rect 9140 3088 9149 3128
rect 3679 3004 3688 3044
rect 3728 3004 3770 3044
rect 3810 3004 3852 3044
rect 3892 3004 3934 3044
rect 3974 3004 4016 3044
rect 4056 3004 4065 3044
rect 7267 3004 7276 3044
rect 7316 3004 9868 3044
rect 9908 3004 9917 3044
rect 11884 2960 11924 3256
rect 15916 3212 15956 3256
rect 18019 3255 18077 3256
rect 20140 3212 20180 3424
rect 21424 3404 21504 3424
rect 15427 3172 15436 3212
rect 15476 3172 15820 3212
rect 15860 3172 15869 3212
rect 15916 3172 20180 3212
rect 17923 3128 17981 3129
rect 20803 3128 20861 3129
rect 21424 3128 21504 3148
rect 16492 3088 17932 3128
rect 17972 3088 19276 3128
rect 19316 3088 19325 3128
rect 20803 3088 20812 3128
rect 20852 3088 21504 3128
rect 16492 3044 16532 3088
rect 17923 3087 17981 3088
rect 20803 3087 20861 3088
rect 21424 3068 21504 3088
rect 11971 3004 11980 3044
rect 12020 3004 16532 3044
rect 16579 3004 16588 3044
rect 16628 3004 18220 3044
rect 18260 3004 18269 3044
rect 18799 3004 18808 3044
rect 18848 3004 18890 3044
rect 18930 3004 18972 3044
rect 19012 3004 19054 3044
rect 19094 3004 19136 3044
rect 19176 3004 19185 3044
rect 6499 2920 6508 2960
rect 6548 2920 7084 2960
rect 7124 2920 8332 2960
rect 8372 2920 8381 2960
rect 8428 2920 11924 2960
rect 16483 2920 16492 2960
rect 16532 2920 18124 2960
rect 18164 2920 18173 2960
rect 8428 2876 8468 2920
rect 2659 2836 2668 2876
rect 2708 2836 3436 2876
rect 3476 2836 3485 2876
rect 4963 2836 4972 2876
rect 5012 2836 5260 2876
rect 5300 2836 5309 2876
rect 6883 2836 6892 2876
rect 6932 2836 8140 2876
rect 8180 2836 8189 2876
rect 8419 2836 8428 2876
rect 8468 2836 8477 2876
rect 9187 2836 9196 2876
rect 9236 2836 10156 2876
rect 10196 2836 18316 2876
rect 18356 2836 18365 2876
rect 18595 2836 18604 2876
rect 18644 2836 20180 2876
rect 0 2792 80 2812
rect 5260 2792 5300 2836
rect 16291 2792 16349 2793
rect 20140 2792 20180 2836
rect 21424 2792 21504 2812
rect 0 2752 460 2792
rect 500 2752 509 2792
rect 5260 2752 6796 2792
rect 6836 2752 6845 2792
rect 8035 2752 8044 2792
rect 8084 2752 11500 2792
rect 11540 2752 14324 2792
rect 15331 2752 15340 2792
rect 15380 2752 15820 2792
rect 15860 2752 15869 2792
rect 15916 2752 16300 2792
rect 16340 2752 16349 2792
rect 16483 2752 16492 2792
rect 16532 2752 17452 2792
rect 17492 2752 17501 2792
rect 20140 2752 21504 2792
rect 0 2732 80 2752
rect 6691 2708 6749 2709
rect 3907 2668 3916 2708
rect 3956 2668 6700 2708
rect 6740 2668 6749 2708
rect 6691 2667 6749 2668
rect 7459 2708 7517 2709
rect 14179 2708 14237 2709
rect 7459 2668 7468 2708
rect 7508 2668 7948 2708
rect 7988 2668 8428 2708
rect 8468 2668 8477 2708
rect 14094 2668 14188 2708
rect 14228 2668 14237 2708
rect 14284 2708 14324 2752
rect 15916 2708 15956 2752
rect 16291 2751 16349 2752
rect 21424 2732 21504 2752
rect 14284 2668 15956 2708
rect 17443 2708 17501 2709
rect 17443 2668 17452 2708
rect 17492 2668 17501 2708
rect 18499 2668 18508 2708
rect 18548 2668 19180 2708
rect 19220 2668 19564 2708
rect 19604 2668 19613 2708
rect 7459 2667 7517 2668
rect 14179 2667 14237 2668
rect 17443 2667 17501 2668
rect 16291 2624 16349 2625
rect 17155 2624 17213 2625
rect 17452 2624 17492 2667
rect 1603 2584 1612 2624
rect 1652 2584 5836 2624
rect 5876 2584 5885 2624
rect 6796 2584 7180 2624
rect 7220 2584 7229 2624
rect 8707 2584 8716 2624
rect 8756 2584 9100 2624
rect 9140 2584 9676 2624
rect 9716 2584 10100 2624
rect 11011 2584 11020 2624
rect 11060 2584 13036 2624
rect 13076 2584 13085 2624
rect 14851 2584 14860 2624
rect 14900 2584 14909 2624
rect 15715 2584 15724 2624
rect 15764 2584 16012 2624
rect 16052 2584 16061 2624
rect 16108 2584 16300 2624
rect 16340 2584 16349 2624
rect 16675 2584 16684 2624
rect 16724 2584 16972 2624
rect 17012 2584 17021 2624
rect 17155 2584 17164 2624
rect 17204 2584 17260 2624
rect 17300 2584 17492 2624
rect 18595 2584 18604 2624
rect 18644 2584 18653 2624
rect 19363 2584 19372 2624
rect 19412 2584 19756 2624
rect 19796 2584 19805 2624
rect 1699 2500 1708 2540
rect 1748 2500 2540 2540
rect 2500 2456 2540 2500
rect 6796 2456 6836 2584
rect 10060 2540 10100 2584
rect 7236 2500 7276 2540
rect 7316 2500 7325 2540
rect 7524 2500 7564 2540
rect 7604 2500 7613 2540
rect 10051 2500 10060 2540
rect 10100 2500 10109 2540
rect 11203 2500 11212 2540
rect 11252 2500 11540 2540
rect 12612 2500 12652 2540
rect 12692 2500 12701 2540
rect 7276 2456 7316 2500
rect 2500 2416 6836 2456
rect 6892 2416 7316 2456
rect 7564 2456 7604 2500
rect 11500 2456 11540 2500
rect 12652 2456 12692 2500
rect 14860 2456 14900 2584
rect 7564 2416 8908 2456
rect 8948 2416 8957 2456
rect 11320 2416 11444 2456
rect 11500 2416 12692 2456
rect 14851 2416 14860 2456
rect 14900 2416 14909 2456
rect 6892 2372 6932 2416
rect 7651 2372 7709 2373
rect 6883 2332 6892 2372
rect 6932 2332 6941 2372
rect 7555 2332 7564 2372
rect 7604 2332 7660 2372
rect 7700 2332 7709 2372
rect 7651 2331 7709 2332
rect 7843 2372 7901 2373
rect 8611 2372 8669 2373
rect 11320 2372 11360 2416
rect 7843 2332 7852 2372
rect 7892 2332 8620 2372
rect 8660 2332 11360 2372
rect 11404 2372 11444 2416
rect 11404 2332 15244 2372
rect 15284 2332 15293 2372
rect 7843 2331 7901 2332
rect 8611 2331 8669 2332
rect 13891 2288 13949 2289
rect 16108 2288 16148 2584
rect 16291 2583 16349 2584
rect 17155 2583 17213 2584
rect 16579 2540 16637 2541
rect 16494 2500 16588 2540
rect 16628 2500 16637 2540
rect 16579 2499 16637 2500
rect 16675 2456 16733 2457
rect 16483 2416 16492 2456
rect 16532 2416 16684 2456
rect 16724 2416 16733 2456
rect 18604 2456 18644 2584
rect 19812 2500 19852 2540
rect 19892 2500 19901 2540
rect 19852 2456 19892 2500
rect 21424 2456 21504 2476
rect 18604 2416 19892 2456
rect 20140 2416 21504 2456
rect 16675 2415 16733 2416
rect 16195 2372 16253 2373
rect 20140 2372 20180 2416
rect 21424 2396 21504 2416
rect 16195 2332 16204 2372
rect 16244 2332 16588 2372
rect 16628 2332 16637 2372
rect 18508 2332 20180 2372
rect 16195 2331 16253 2332
rect 18508 2288 18548 2332
rect 4919 2248 4928 2288
rect 4968 2248 5010 2288
rect 5050 2248 5092 2288
rect 5132 2248 5174 2288
rect 5214 2248 5256 2288
rect 5296 2248 5305 2288
rect 7267 2248 7276 2288
rect 7316 2248 7660 2288
rect 7700 2248 7709 2288
rect 8035 2248 8044 2288
rect 8084 2248 8716 2288
rect 8756 2248 8765 2288
rect 10147 2248 10156 2288
rect 10196 2248 12748 2288
rect 12788 2248 12797 2288
rect 13891 2248 13900 2288
rect 13940 2248 15724 2288
rect 15764 2248 15773 2288
rect 16108 2248 18548 2288
rect 20039 2248 20048 2288
rect 20088 2248 20130 2288
rect 20170 2248 20212 2288
rect 20252 2248 20294 2288
rect 20334 2248 20376 2288
rect 20416 2248 20425 2288
rect 13891 2247 13949 2248
rect 8515 2204 8573 2205
rect 6691 2164 6700 2204
rect 6740 2164 7180 2204
rect 7220 2164 7229 2204
rect 7276 2164 8524 2204
rect 8564 2164 8573 2204
rect 13411 2164 13420 2204
rect 13460 2164 13804 2204
rect 13844 2164 13853 2204
rect 14083 2164 14092 2204
rect 14132 2164 14956 2204
rect 14996 2164 15005 2204
rect 16963 2164 16972 2204
rect 17012 2164 17260 2204
rect 17300 2164 17309 2204
rect 18019 2164 18028 2204
rect 18068 2164 18508 2204
rect 18548 2164 18557 2204
rect 7276 2120 7316 2164
rect 8515 2163 8573 2164
rect 4771 2080 4780 2120
rect 4820 2080 7316 2120
rect 7555 2120 7613 2121
rect 21424 2120 21504 2140
rect 7555 2080 7564 2120
rect 7604 2080 21504 2120
rect 7555 2079 7613 2080
rect 21424 2060 21504 2080
rect 18115 2036 18173 2037
rect 5635 1996 5644 2036
rect 5684 1996 9676 2036
rect 9716 1996 9725 2036
rect 13804 1996 18124 2036
rect 18164 1996 19948 2036
rect 19988 1996 19997 2036
rect 5539 1952 5597 1953
rect 1315 1912 1324 1952
rect 1364 1912 4780 1952
rect 4820 1912 4829 1952
rect 4963 1912 4972 1952
rect 5012 1912 5548 1952
rect 5588 1912 5597 1952
rect 6307 1912 6316 1952
rect 6356 1912 6988 1952
rect 7028 1912 7037 1952
rect 7171 1912 7180 1952
rect 7220 1912 8236 1952
rect 8276 1912 8285 1952
rect 8428 1912 9004 1952
rect 9044 1912 9484 1952
rect 9524 1912 9772 1952
rect 9812 1912 9821 1952
rect 10156 1912 12596 1952
rect 5539 1911 5597 1912
rect 2275 1868 2333 1869
rect 8428 1868 8468 1912
rect 8611 1868 8669 1869
rect 10156 1868 10196 1912
rect 10339 1868 10397 1869
rect 10819 1868 10877 1869
rect 11107 1868 11165 1869
rect 2275 1828 2284 1868
rect 2324 1828 2956 1868
rect 2996 1828 3005 1868
rect 6403 1828 6412 1868
rect 6452 1828 7852 1868
rect 7892 1828 8428 1868
rect 8468 1828 8477 1868
rect 8611 1828 8620 1868
rect 8660 1828 10196 1868
rect 10254 1828 10348 1868
rect 10388 1828 10397 1868
rect 10723 1828 10732 1868
rect 10772 1828 10828 1868
rect 10868 1828 10877 1868
rect 11022 1828 11116 1868
rect 11156 1828 11165 1868
rect 2275 1827 2333 1828
rect 8611 1827 8669 1828
rect 10339 1827 10397 1828
rect 10819 1827 10877 1828
rect 11107 1827 11165 1828
rect 7459 1784 7517 1785
rect 8515 1784 8573 1785
rect 3523 1744 3532 1784
rect 3572 1744 4108 1784
rect 4148 1744 5356 1784
rect 5396 1744 6220 1784
rect 6260 1744 7468 1784
rect 7508 1744 7517 1784
rect 7651 1744 7660 1784
rect 7700 1744 8044 1784
rect 8084 1744 8093 1784
rect 8515 1744 8524 1784
rect 8564 1744 11500 1784
rect 11540 1744 11549 1784
rect 7459 1743 7517 1744
rect 8515 1743 8573 1744
rect 12556 1700 12596 1912
rect 13804 1868 13844 1996
rect 18115 1995 18173 1996
rect 14371 1912 14380 1952
rect 14420 1912 14956 1952
rect 14996 1912 15005 1952
rect 16387 1912 16396 1952
rect 16436 1912 17164 1952
rect 17204 1912 17213 1952
rect 18115 1912 18124 1952
rect 18164 1912 18173 1952
rect 18124 1868 18164 1912
rect 12643 1828 12652 1868
rect 12692 1828 13804 1868
rect 13844 1828 13853 1868
rect 16771 1828 16780 1868
rect 16820 1828 18164 1868
rect 20899 1784 20957 1785
rect 21424 1784 21504 1804
rect 12739 1744 12748 1784
rect 12788 1744 14188 1784
rect 14228 1744 16492 1784
rect 16532 1744 17260 1784
rect 17300 1744 17309 1784
rect 20899 1744 20908 1784
rect 20948 1744 21504 1784
rect 20899 1743 20957 1744
rect 21424 1724 21504 1744
rect 13219 1700 13277 1701
rect 1795 1660 1804 1700
rect 1844 1660 2540 1700
rect 3139 1660 3148 1700
rect 3188 1660 8908 1700
rect 8948 1660 8957 1700
rect 11299 1660 11308 1700
rect 11348 1660 12364 1700
rect 12404 1660 12413 1700
rect 12556 1660 13228 1700
rect 13268 1660 16012 1700
rect 16052 1660 16061 1700
rect 2500 1616 2540 1660
rect 13219 1659 13277 1660
rect 15043 1616 15101 1617
rect 2500 1576 3340 1616
rect 3380 1576 5012 1616
rect 6595 1576 6604 1616
rect 6644 1576 14860 1616
rect 14900 1576 14909 1616
rect 15043 1576 15052 1616
rect 15092 1576 19276 1616
rect 19316 1576 19325 1616
rect 4972 1532 5012 1576
rect 15043 1575 15101 1576
rect 1795 1492 1804 1532
rect 1844 1492 2092 1532
rect 2132 1492 2141 1532
rect 3679 1492 3688 1532
rect 3728 1492 3770 1532
rect 3810 1492 3852 1532
rect 3892 1492 3934 1532
rect 3974 1492 4016 1532
rect 4056 1492 4065 1532
rect 4963 1492 4972 1532
rect 5012 1492 7660 1532
rect 7700 1492 7709 1532
rect 8419 1492 8428 1532
rect 8468 1492 14572 1532
rect 14612 1492 14621 1532
rect 15820 1492 17932 1532
rect 17972 1492 17981 1532
rect 18799 1492 18808 1532
rect 18848 1492 18890 1532
rect 18930 1492 18972 1532
rect 19012 1492 19054 1532
rect 19094 1492 19136 1532
rect 19176 1492 19185 1532
rect 13699 1448 13757 1449
rect 15820 1448 15860 1492
rect 21424 1448 21504 1468
rect 4867 1408 4876 1448
rect 4916 1408 5932 1448
rect 5972 1408 5981 1448
rect 6499 1408 6508 1448
rect 6548 1408 6892 1448
rect 6932 1408 6941 1448
rect 7939 1408 7948 1448
rect 7988 1408 8716 1448
rect 8756 1408 8765 1448
rect 9379 1408 9388 1448
rect 9428 1408 11116 1448
rect 11156 1408 11165 1448
rect 13699 1408 13708 1448
rect 13748 1408 15860 1448
rect 16195 1408 16204 1448
rect 16244 1408 19468 1448
rect 19508 1408 19517 1448
rect 19939 1408 19948 1448
rect 19988 1408 21504 1448
rect 13699 1407 13757 1408
rect 21424 1388 21504 1408
rect 6019 1324 6028 1364
rect 6068 1324 8140 1364
rect 8180 1324 8189 1364
rect 10915 1324 10924 1364
rect 10964 1324 12172 1364
rect 12212 1324 12221 1364
rect 13987 1324 13996 1364
rect 14036 1324 16684 1364
rect 16724 1324 16733 1364
rect 16963 1324 16972 1364
rect 17012 1324 17260 1364
rect 17300 1324 17309 1364
rect 3331 1280 3389 1281
rect 3246 1240 3340 1280
rect 3380 1240 3389 1280
rect 3331 1239 3389 1240
rect 3523 1280 3581 1281
rect 5443 1280 5501 1281
rect 6595 1280 6653 1281
rect 7747 1280 7805 1281
rect 9283 1280 9341 1281
rect 14083 1280 14141 1281
rect 16771 1280 16829 1281
rect 17539 1280 17597 1281
rect 18691 1280 18749 1281
rect 19459 1280 19517 1281
rect 3523 1240 3532 1280
rect 3572 1240 3724 1280
rect 3764 1240 5300 1280
rect 5358 1240 5452 1280
rect 5492 1240 5501 1280
rect 6115 1240 6124 1280
rect 6164 1240 6604 1280
rect 6644 1240 6653 1280
rect 6787 1240 6796 1280
rect 6836 1240 7084 1280
rect 7124 1240 7133 1280
rect 7662 1240 7756 1280
rect 7796 1240 7805 1280
rect 3523 1239 3581 1240
rect 643 1196 701 1197
rect 5260 1196 5300 1240
rect 5443 1239 5501 1240
rect 6595 1239 6653 1240
rect 7747 1239 7805 1240
rect 7852 1240 8180 1280
rect 8323 1240 8332 1280
rect 8372 1240 9292 1280
rect 9332 1240 9341 1280
rect 10531 1240 10540 1280
rect 10580 1240 11692 1280
rect 11732 1240 11741 1280
rect 12547 1240 12556 1280
rect 12596 1240 14092 1280
rect 14132 1240 14141 1280
rect 16686 1240 16780 1280
rect 16820 1240 16829 1280
rect 17454 1240 17548 1280
rect 17588 1240 17597 1280
rect 18606 1240 18700 1280
rect 18740 1240 18749 1280
rect 19374 1240 19468 1280
rect 19508 1240 19517 1280
rect 7171 1196 7229 1197
rect 7852 1196 7892 1240
rect 8035 1196 8093 1197
rect 643 1156 652 1196
rect 692 1156 3916 1196
rect 3956 1156 3965 1196
rect 5260 1156 5644 1196
rect 5684 1156 5693 1196
rect 6883 1156 6892 1196
rect 6932 1156 6941 1196
rect 7171 1156 7180 1196
rect 7220 1156 7892 1196
rect 7950 1156 8044 1196
rect 8084 1156 8093 1196
rect 8140 1196 8180 1240
rect 9283 1239 9341 1240
rect 14083 1239 14141 1240
rect 16771 1239 16829 1240
rect 17539 1239 17597 1240
rect 18691 1239 18749 1240
rect 19459 1239 19517 1240
rect 9571 1196 9629 1197
rect 10051 1196 10109 1197
rect 8140 1156 9100 1196
rect 9140 1156 9149 1196
rect 9571 1156 9580 1196
rect 9620 1156 9868 1196
rect 9908 1156 9917 1196
rect 10051 1156 10060 1196
rect 10100 1156 10348 1196
rect 10388 1156 10397 1196
rect 10627 1156 10636 1196
rect 10676 1156 14860 1196
rect 14900 1156 14909 1196
rect 15523 1156 15532 1196
rect 15572 1156 16396 1196
rect 16436 1156 16445 1196
rect 16492 1156 20180 1196
rect 643 1155 701 1156
rect 4771 1112 4829 1113
rect 6892 1112 6932 1156
rect 7171 1155 7229 1156
rect 8035 1155 8093 1156
rect 9571 1155 9629 1156
rect 10051 1155 10109 1156
rect 14467 1112 14525 1113
rect 16492 1112 16532 1156
rect 20140 1112 20180 1156
rect 21424 1112 21504 1132
rect 4195 1072 4204 1112
rect 4244 1072 4780 1112
rect 4820 1072 4829 1112
rect 5059 1072 5068 1112
rect 5108 1072 6508 1112
rect 6548 1072 6557 1112
rect 6604 1072 7372 1112
rect 7412 1072 7421 1112
rect 7468 1072 11360 1112
rect 12739 1072 12748 1112
rect 12788 1072 14476 1112
rect 14516 1072 14525 1112
rect 4771 1071 4829 1072
rect 1123 1028 1181 1029
rect 6604 1028 6644 1072
rect 7468 1028 7508 1072
rect 10819 1028 10877 1029
rect 11203 1028 11261 1029
rect 1123 988 1132 1028
rect 1172 988 3532 1028
rect 3572 988 3581 1028
rect 4483 988 4492 1028
rect 4532 988 5740 1028
rect 5780 988 5789 1028
rect 5836 988 6644 1028
rect 7075 988 7084 1028
rect 7124 988 7412 1028
rect 7456 988 7465 1028
rect 7505 988 7514 1028
rect 7756 988 8716 1028
rect 8756 988 8765 1028
rect 9091 988 9100 1028
rect 9140 988 10828 1028
rect 10868 988 10877 1028
rect 11118 988 11212 1028
rect 11252 988 11261 1028
rect 11320 1028 11360 1072
rect 14467 1071 14525 1072
rect 14572 1072 16532 1112
rect 17155 1072 17164 1112
rect 17204 1072 17644 1112
rect 17684 1072 17693 1112
rect 20140 1072 21504 1112
rect 13507 1028 13565 1029
rect 11320 988 12652 1028
rect 12692 988 12701 1028
rect 13422 988 13516 1028
rect 13556 988 13565 1028
rect 1123 987 1181 988
rect 2755 944 2813 945
rect 4099 944 4157 945
rect 4771 944 4829 945
rect 5836 944 5876 988
rect 7372 944 7412 988
rect 7756 944 7796 988
rect 10819 987 10877 988
rect 11203 987 11261 988
rect 13507 987 13565 988
rect 7939 944 7997 945
rect 14572 944 14612 1072
rect 21424 1052 21504 1072
rect 17827 1028 17885 1029
rect 16387 988 16396 1028
rect 16436 988 17836 1028
rect 17876 988 19372 1028
rect 19412 988 19660 1028
rect 19700 988 19709 1028
rect 17827 987 17885 988
rect 15907 944 15965 945
rect 18115 944 18173 945
rect 19267 944 19325 945
rect 2670 904 2764 944
rect 2804 904 2813 944
rect 4014 904 4108 944
rect 4148 904 4157 944
rect 4579 904 4588 944
rect 4628 904 4637 944
rect 4771 904 4780 944
rect 4820 904 5356 944
rect 5396 904 5876 944
rect 6595 904 6604 944
rect 6644 904 7180 944
rect 7220 904 7229 944
rect 7372 904 7796 944
rect 7854 904 7948 944
rect 7988 904 7997 944
rect 8611 904 8620 944
rect 8660 904 9484 944
rect 9524 904 9533 944
rect 10243 904 10252 944
rect 10292 904 10732 944
rect 10772 904 10781 944
rect 11395 904 11404 944
rect 11444 904 11980 944
rect 12020 904 12029 944
rect 13315 904 13324 944
rect 13364 904 14612 944
rect 14851 904 14860 944
rect 14900 904 15340 944
rect 15380 904 15389 944
rect 15907 904 15916 944
rect 15956 904 17740 944
rect 17780 904 17789 944
rect 18030 904 18124 944
rect 18164 904 18173 944
rect 18883 904 18892 944
rect 18932 904 19276 944
rect 19316 904 19325 944
rect 2755 903 2813 904
rect 4099 903 4157 904
rect 4588 860 4628 904
rect 4771 903 4829 904
rect 7939 903 7997 904
rect 15907 903 15965 904
rect 18115 903 18173 904
rect 19267 903 19325 904
rect 14275 860 14333 861
rect 16867 860 16925 861
rect 17923 860 17981 861
rect 4588 820 9100 860
rect 9140 820 9149 860
rect 10819 820 10828 860
rect 10868 820 13420 860
rect 13460 820 13469 860
rect 14190 820 14284 860
rect 14324 820 14333 860
rect 14467 820 14476 860
rect 14516 820 16876 860
rect 16916 820 16925 860
rect 17443 820 17452 860
rect 17492 820 17932 860
rect 17972 820 17981 860
rect 14275 819 14333 820
rect 16867 819 16925 820
rect 17923 819 17981 820
rect 2563 776 2621 777
rect 6979 776 7037 777
rect 13699 776 13757 777
rect 21424 776 21504 796
rect 2563 736 2572 776
rect 2612 736 2706 776
rect 4919 736 4928 776
rect 4968 736 5010 776
rect 5050 736 5092 776
rect 5132 736 5174 776
rect 5214 736 5256 776
rect 5296 736 5305 776
rect 6979 736 6988 776
rect 7028 736 8524 776
rect 8564 736 8573 776
rect 9283 736 9292 776
rect 9332 736 11360 776
rect 13614 736 13708 776
rect 13748 736 13757 776
rect 16099 736 16108 776
rect 16148 736 17164 776
rect 17204 736 17213 776
rect 20039 736 20048 776
rect 20088 736 20130 776
rect 20170 736 20212 776
rect 20252 736 20294 776
rect 20334 736 20376 776
rect 20416 736 20425 776
rect 21292 736 21504 776
rect 2563 735 2621 736
rect 6979 735 7037 736
rect 5923 692 5981 693
rect 2659 652 2668 692
rect 2708 652 5780 692
rect 5827 652 5836 692
rect 5876 652 5932 692
rect 5972 652 5981 692
rect 1027 608 1085 609
rect 4675 608 4733 609
rect 5347 608 5405 609
rect 1027 568 1036 608
rect 1076 568 4300 608
rect 4340 568 4349 608
rect 4675 568 4684 608
rect 4724 568 4876 608
rect 4916 568 4925 608
rect 5251 568 5260 608
rect 5300 568 5356 608
rect 5396 568 5405 608
rect 5740 608 5780 652
rect 5923 651 5981 652
rect 6499 692 6557 693
rect 11320 692 11360 736
rect 13699 735 13757 736
rect 6499 652 6508 692
rect 6548 652 7564 692
rect 7604 652 7613 692
rect 7843 652 7852 692
rect 7892 652 10444 692
rect 10484 652 10493 692
rect 11320 652 20180 692
rect 6499 651 6557 652
rect 7939 608 7997 609
rect 8131 608 8189 609
rect 15427 608 15485 609
rect 5740 568 7948 608
rect 7988 568 7997 608
rect 8046 568 8140 608
rect 8180 568 8189 608
rect 9859 568 9868 608
rect 9908 568 11596 608
rect 11636 568 11645 608
rect 13315 568 13324 608
rect 13364 568 15436 608
rect 15476 568 15485 608
rect 1027 567 1085 568
rect 4675 567 4733 568
rect 5347 567 5405 568
rect 7939 567 7997 568
rect 8131 567 8189 568
rect 15427 567 15485 568
rect 17059 608 17117 609
rect 20140 608 20180 652
rect 21292 608 21332 736
rect 21424 716 21504 736
rect 17059 568 17068 608
rect 17108 568 18508 608
rect 18548 568 18557 608
rect 20140 568 21332 608
rect 17059 567 17117 568
rect 2467 524 2525 525
rect 7363 524 7421 525
rect 14851 524 14909 525
rect 2467 484 2476 524
rect 2516 484 5068 524
rect 5108 484 5117 524
rect 5635 484 5644 524
rect 5684 484 6548 524
rect 7278 484 7372 524
rect 7412 484 7421 524
rect 8227 484 8236 524
rect 8276 484 9292 524
rect 9332 484 9341 524
rect 10531 484 10540 524
rect 10580 484 11404 524
rect 11444 484 11453 524
rect 13123 484 13132 524
rect 13172 484 14860 524
rect 14900 484 14909 524
rect 16675 484 16684 524
rect 16724 484 17356 524
rect 17396 484 17405 524
rect 2467 483 2525 484
rect 6403 440 6461 441
rect 6318 400 6412 440
rect 6452 400 6461 440
rect 6508 440 6548 484
rect 7363 483 7421 484
rect 14851 483 14909 484
rect 15235 440 15293 441
rect 21424 440 21504 460
rect 6508 400 7316 440
rect 10147 400 10156 440
rect 10196 400 11596 440
rect 11636 400 11645 440
rect 12931 400 12940 440
rect 12980 400 15244 440
rect 15284 400 15293 440
rect 6403 399 6461 400
rect 2371 356 2429 357
rect 6883 356 6941 357
rect 2371 316 2380 356
rect 2420 316 6836 356
rect 2371 315 2429 316
rect 2179 272 2237 273
rect 6796 272 6836 316
rect 6883 316 6892 356
rect 6932 316 7180 356
rect 7220 316 7229 356
rect 6883 315 6941 316
rect 7276 272 7316 400
rect 15235 399 15293 400
rect 20140 400 21504 440
rect 14083 356 14141 357
rect 20140 356 20180 400
rect 21424 380 21504 400
rect 8995 316 9004 356
rect 9044 316 11020 356
rect 11060 316 11069 356
rect 13998 316 14092 356
rect 14132 316 14141 356
rect 14083 315 14141 316
rect 15820 316 20180 356
rect 12163 272 12221 273
rect 15715 272 15773 273
rect 1891 232 1900 272
rect 1940 232 2036 272
rect 1996 104 2036 232
rect 2179 232 2188 272
rect 2228 232 6604 272
rect 6644 232 6653 272
rect 6796 232 6988 272
rect 7028 232 7037 272
rect 7276 232 12172 272
rect 12212 232 12221 272
rect 13891 232 13900 272
rect 13940 232 15724 272
rect 15764 232 15773 272
rect 2179 231 2237 232
rect 12163 231 12221 232
rect 15715 231 15773 232
rect 13603 188 13661 189
rect 7276 148 13612 188
rect 13652 148 13661 188
rect 7276 104 7316 148
rect 13603 147 13661 148
rect 1987 64 1996 104
rect 2036 64 2045 104
rect 6211 64 6220 104
rect 6260 64 7316 104
rect 7939 104 7997 105
rect 10819 104 10877 105
rect 15820 104 15860 316
rect 17251 272 17309 273
rect 17251 232 17260 272
rect 17300 232 19084 272
rect 19124 232 19133 272
rect 17251 231 17309 232
rect 7939 64 7948 104
rect 7988 64 10636 104
rect 10676 64 10685 104
rect 10819 64 10828 104
rect 10868 64 15860 104
rect 17155 104 17213 105
rect 21424 104 21504 124
rect 17155 64 17164 104
rect 17204 64 21504 104
rect 7939 63 7997 64
rect 10819 63 10877 64
rect 17155 63 17213 64
rect 21424 44 21504 64
<< via3 >>
rect 20620 42736 20660 42776
rect 4108 42568 4148 42608
rect 11788 42568 11828 42608
rect 14668 42568 14708 42608
rect 1900 42232 1940 42272
rect 18700 42148 18740 42188
rect 1516 42064 1556 42104
rect 4928 41560 4968 41600
rect 5010 41560 5050 41600
rect 5092 41560 5132 41600
rect 5174 41560 5214 41600
rect 5256 41560 5296 41600
rect 9868 41560 9908 41600
rect 10060 41560 10100 41600
rect 11404 41560 11444 41600
rect 11596 41560 11636 41600
rect 17932 41560 17972 41600
rect 18508 41560 18548 41600
rect 20048 41560 20088 41600
rect 20130 41560 20170 41600
rect 20212 41560 20252 41600
rect 20294 41560 20334 41600
rect 20376 41560 20416 41600
rect 20812 41392 20852 41432
rect 1804 41224 1844 41264
rect 2764 41224 2804 41264
rect 16684 41224 16724 41264
rect 8044 41140 8084 41180
rect 19756 41140 19796 41180
rect 13324 40972 13364 41012
rect 19852 41056 19892 41096
rect 15628 40972 15668 41012
rect 16012 40972 16052 41012
rect 3052 40804 3092 40844
rect 3688 40804 3728 40844
rect 3770 40804 3810 40844
rect 3852 40804 3892 40844
rect 3934 40804 3974 40844
rect 4016 40804 4056 40844
rect 4204 40804 4244 40844
rect 17644 40804 17684 40844
rect 18808 40804 18848 40844
rect 18890 40804 18930 40844
rect 18972 40804 19012 40844
rect 19054 40804 19094 40844
rect 19136 40804 19176 40844
rect 10924 40636 10964 40676
rect 3340 40552 3380 40592
rect 14092 40552 14132 40592
rect 14476 40552 14516 40592
rect 14860 40552 14900 40592
rect 5836 40384 5876 40424
rect 10828 40384 10868 40424
rect 15148 40552 15188 40592
rect 15820 40552 15860 40592
rect 16396 40552 16436 40592
rect 18892 40468 18932 40508
rect 19660 40468 19700 40508
rect 9772 40300 9812 40340
rect 14956 40300 14996 40340
rect 15244 40300 15284 40340
rect 3052 40216 3092 40256
rect 10252 40216 10292 40256
rect 15628 40300 15668 40340
rect 17356 40300 17396 40340
rect 19852 40300 19892 40340
rect 18700 40216 18740 40256
rect 3148 40048 3188 40088
rect 4928 40048 4968 40088
rect 5010 40048 5050 40088
rect 5092 40048 5132 40088
rect 5174 40048 5214 40088
rect 5256 40048 5296 40088
rect 17932 40048 17972 40088
rect 20048 40048 20088 40088
rect 20130 40048 20170 40088
rect 20212 40048 20252 40088
rect 20294 40048 20334 40088
rect 20376 40048 20416 40088
rect 17164 39796 17204 39836
rect 1612 39712 1652 39752
rect 20812 39712 20852 39752
rect 10924 39628 10964 39668
rect 11116 39628 11156 39668
rect 2476 39544 2516 39584
rect 12364 39544 12404 39584
rect 17260 39544 17300 39584
rect 16876 39460 16916 39500
rect 3688 39292 3728 39332
rect 3770 39292 3810 39332
rect 3852 39292 3892 39332
rect 3934 39292 3974 39332
rect 4016 39292 4056 39332
rect 12940 39292 12980 39332
rect 18808 39292 18848 39332
rect 18890 39292 18930 39332
rect 18972 39292 19012 39332
rect 19054 39292 19094 39332
rect 19136 39292 19176 39332
rect 8908 39208 8948 39248
rect 11788 39124 11828 39164
rect 13516 39124 13556 39164
rect 1420 38956 1460 38996
rect 17644 38956 17684 38996
rect 1708 38872 1748 38912
rect 14188 38872 14228 38912
rect 16684 38872 16724 38912
rect 11212 38788 11252 38828
rect 18220 38704 18260 38744
rect 18988 38704 19028 38744
rect 2092 38620 2132 38660
rect 4928 38536 4968 38576
rect 5010 38536 5050 38576
rect 5092 38536 5132 38576
rect 5174 38536 5214 38576
rect 5256 38536 5296 38576
rect 8620 38536 8660 38576
rect 20048 38536 20088 38576
rect 20130 38536 20170 38576
rect 20212 38536 20252 38576
rect 20294 38536 20334 38576
rect 20376 38536 20416 38576
rect 12652 38368 12692 38408
rect 12844 38368 12884 38408
rect 20140 38284 20180 38324
rect 9580 38200 9620 38240
rect 10348 38200 10388 38240
rect 12652 38200 12692 38240
rect 14188 38200 14228 38240
rect 7372 38116 7412 38156
rect 8428 38116 8468 38156
rect 1804 38032 1844 38072
rect 4204 37948 4244 37988
rect 2572 37864 2612 37904
rect 11212 37864 11252 37904
rect 17356 37864 17396 37904
rect 1804 37780 1844 37820
rect 3688 37780 3728 37820
rect 3770 37780 3810 37820
rect 3852 37780 3892 37820
rect 3934 37780 3974 37820
rect 4016 37780 4056 37820
rect 2476 37696 2516 37736
rect 18808 37780 18848 37820
rect 18890 37780 18930 37820
rect 18972 37780 19012 37820
rect 19054 37780 19094 37820
rect 19136 37780 19176 37820
rect 8332 37696 8372 37736
rect 15724 37696 15764 37736
rect 2476 37528 2516 37568
rect 2764 37444 2804 37484
rect 652 37360 692 37400
rect 2380 37360 2420 37400
rect 2572 37360 2612 37400
rect 4204 37360 4244 37400
rect 7564 37360 7604 37400
rect 18124 37360 18164 37400
rect 1228 37276 1268 37316
rect 8332 37276 8372 37316
rect 19660 37276 19700 37316
rect 1996 37192 2036 37232
rect 6892 37192 6932 37232
rect 9196 37108 9236 37148
rect 9388 37108 9428 37148
rect 16300 37108 16340 37148
rect 172 37024 212 37064
rect 4928 37024 4968 37064
rect 5010 37024 5050 37064
rect 5092 37024 5132 37064
rect 5174 37024 5214 37064
rect 5256 37024 5296 37064
rect 20048 37024 20088 37064
rect 20130 37024 20170 37064
rect 20212 37024 20252 37064
rect 20294 37024 20334 37064
rect 20376 37024 20416 37064
rect 2284 36772 2324 36812
rect 2476 36856 2516 36896
rect 3532 36856 3572 36896
rect 14668 36856 14708 36896
rect 21004 36772 21044 36812
rect 5836 36688 5876 36728
rect 12652 36688 12692 36728
rect 11980 36604 12020 36644
rect 6700 36520 6740 36560
rect 18508 36520 18548 36560
rect 21196 36520 21236 36560
rect 940 36436 980 36476
rect 3688 36268 3728 36308
rect 3770 36268 3810 36308
rect 3852 36268 3892 36308
rect 3934 36268 3974 36308
rect 4016 36268 4056 36308
rect 18808 36268 18848 36308
rect 18890 36268 18930 36308
rect 18972 36268 19012 36308
rect 19054 36268 19094 36308
rect 19136 36268 19176 36308
rect 4108 36100 4148 36140
rect 3532 36016 3572 36056
rect 8812 35932 8852 35972
rect 16300 35932 16340 35972
rect 19948 35932 19988 35972
rect 6604 35848 6644 35888
rect 9676 35848 9716 35888
rect 18220 35764 18260 35804
rect 2188 35680 2228 35720
rect 4492 35680 4532 35720
rect 9004 35680 9044 35720
rect 4928 35512 4968 35552
rect 5010 35512 5050 35552
rect 5092 35512 5132 35552
rect 5174 35512 5214 35552
rect 5256 35512 5296 35552
rect 16492 35512 16532 35552
rect 20048 35512 20088 35552
rect 20130 35512 20170 35552
rect 20212 35512 20252 35552
rect 20294 35512 20334 35552
rect 20376 35512 20416 35552
rect 7468 35428 7508 35468
rect 9580 35428 9620 35468
rect 14764 35428 14804 35468
rect 20620 35428 20660 35468
rect 16108 35344 16148 35384
rect 8716 35260 8756 35300
rect 9292 35260 9332 35300
rect 2572 35176 2612 35216
rect 2764 35176 2804 35216
rect 12652 35176 12692 35216
rect 17644 35176 17684 35216
rect 19948 35176 19988 35216
rect 748 35092 788 35132
rect 12844 35092 12884 35132
rect 15916 35092 15956 35132
rect 8716 35008 8756 35048
rect 17068 35008 17108 35048
rect 1132 34840 1172 34880
rect 13036 34840 13076 34880
rect 14668 34840 14708 34880
rect 16108 34840 16148 34880
rect 3688 34756 3728 34796
rect 3770 34756 3810 34796
rect 3852 34756 3892 34796
rect 3934 34756 3974 34796
rect 4016 34756 4056 34796
rect 18808 34756 18848 34796
rect 18890 34756 18930 34796
rect 18972 34756 19012 34796
rect 19054 34756 19094 34796
rect 19136 34756 19176 34796
rect 3148 34672 3188 34712
rect 9388 34672 9428 34712
rect 13804 34672 13844 34712
rect 2668 34588 2708 34628
rect 2092 34504 2132 34544
rect 6604 34420 6644 34460
rect 1132 34336 1172 34376
rect 8140 34336 8180 34376
rect 16780 34336 16820 34376
rect 13804 34252 13844 34292
rect 18508 34168 18548 34208
rect 19564 34168 19604 34208
rect 4928 34000 4968 34040
rect 5010 34000 5050 34040
rect 5092 34000 5132 34040
rect 5174 34000 5214 34040
rect 5256 34000 5296 34040
rect 10444 34000 10484 34040
rect 15436 34000 15476 34040
rect 20048 34000 20088 34040
rect 20130 34000 20170 34040
rect 20212 34000 20252 34040
rect 20294 34000 20334 34040
rect 20376 34000 20416 34040
rect 1036 33916 1076 33956
rect 2476 33916 2516 33956
rect 5452 33664 5492 33704
rect 8236 33664 8276 33704
rect 10444 33664 10484 33704
rect 844 33580 884 33620
rect 4684 33580 4724 33620
rect 18604 33580 18644 33620
rect 2860 33496 2900 33536
rect 2476 33412 2516 33452
rect 9292 33412 9332 33452
rect 18412 33412 18452 33452
rect 20812 33412 20852 33452
rect 12652 33328 12692 33368
rect 3688 33244 3728 33284
rect 3770 33244 3810 33284
rect 3852 33244 3892 33284
rect 3934 33244 3974 33284
rect 4016 33244 4056 33284
rect 6220 33244 6260 33284
rect 7180 33244 7220 33284
rect 9292 33244 9332 33284
rect 1516 33160 1556 33200
rect 1900 33160 1940 33200
rect 5836 33160 5876 33200
rect 18808 33244 18848 33284
rect 18890 33244 18930 33284
rect 18972 33244 19012 33284
rect 19054 33244 19094 33284
rect 19136 33244 19176 33284
rect 19852 33160 19892 33200
rect 14572 33076 14612 33116
rect 16972 33076 17012 33116
rect 19660 33076 19700 33116
rect 17452 32992 17492 33032
rect 1324 32908 1364 32948
rect 2572 32908 2612 32948
rect 3724 32908 3764 32948
rect 1804 32824 1844 32864
rect 4204 32824 4244 32864
rect 10156 32824 10196 32864
rect 12652 32824 12692 32864
rect 4300 32740 4340 32780
rect 7084 32740 7124 32780
rect 19948 32740 19988 32780
rect 6220 32656 6260 32696
rect 8620 32572 8660 32612
rect 4928 32488 4968 32528
rect 5010 32488 5050 32528
rect 5092 32488 5132 32528
rect 5174 32488 5214 32528
rect 5256 32488 5296 32528
rect 20048 32488 20088 32528
rect 20130 32488 20170 32528
rect 20212 32488 20252 32528
rect 20294 32488 20334 32528
rect 20376 32488 20416 32528
rect 16972 32320 17012 32360
rect 17452 32320 17492 32360
rect 19564 32320 19604 32360
rect 2476 32236 2516 32276
rect 4684 32152 4724 32192
rect 8620 32152 8660 32192
rect 12268 32068 12308 32108
rect 13612 32068 13652 32108
rect 3688 31732 3728 31772
rect 3770 31732 3810 31772
rect 3852 31732 3892 31772
rect 3934 31732 3974 31772
rect 4016 31732 4056 31772
rect 18808 31732 18848 31772
rect 18890 31732 18930 31772
rect 18972 31732 19012 31772
rect 19054 31732 19094 31772
rect 19136 31732 19176 31772
rect 7756 31648 7796 31688
rect 7084 31564 7124 31604
rect 2380 31480 2420 31520
rect 2668 31312 2708 31352
rect 6988 31312 7028 31352
rect 10636 31564 10676 31604
rect 19852 31480 19892 31520
rect 20524 31480 20564 31520
rect 16492 31396 16532 31436
rect 19852 31312 19892 31352
rect 18604 31144 18644 31184
rect 19276 31144 19316 31184
rect 4928 30976 4968 31016
rect 5010 30976 5050 31016
rect 5092 30976 5132 31016
rect 5174 30976 5214 31016
rect 5256 30976 5296 31016
rect 20048 30976 20088 31016
rect 20130 30976 20170 31016
rect 20212 30976 20252 31016
rect 20294 30976 20334 31016
rect 20376 30976 20416 31016
rect 21196 30976 21236 31016
rect 4780 30808 4820 30848
rect 7468 30808 7508 30848
rect 16684 30808 16724 30848
rect 17068 30808 17108 30848
rect 7276 30640 7316 30680
rect 15724 30640 15764 30680
rect 16780 30640 16820 30680
rect 18604 30640 18644 30680
rect 19948 30640 19988 30680
rect 1132 30472 1172 30512
rect 14572 30472 14612 30512
rect 19660 30304 19700 30344
rect 1708 30220 1748 30260
rect 3688 30220 3728 30260
rect 3770 30220 3810 30260
rect 3852 30220 3892 30260
rect 3934 30220 3974 30260
rect 4016 30220 4056 30260
rect 14764 30220 14804 30260
rect 18808 30220 18848 30260
rect 18890 30220 18930 30260
rect 18972 30220 19012 30260
rect 19054 30220 19094 30260
rect 19136 30220 19176 30260
rect 19948 30220 19988 30260
rect 7084 29884 7124 29924
rect 17740 29884 17780 29924
rect 2668 29800 2708 29840
rect 17548 29800 17588 29840
rect 17836 29800 17876 29840
rect 7180 29716 7220 29756
rect 15436 29716 15476 29756
rect 1708 29464 1748 29504
rect 4928 29464 4968 29504
rect 5010 29464 5050 29504
rect 5092 29464 5132 29504
rect 5174 29464 5214 29504
rect 5256 29464 5296 29504
rect 20048 29464 20088 29504
rect 20130 29464 20170 29504
rect 20212 29464 20252 29504
rect 20294 29464 20334 29504
rect 20376 29464 20416 29504
rect 12844 29296 12884 29336
rect 18316 29296 18356 29336
rect 20812 29296 20852 29336
rect 5452 29212 5492 29252
rect 2284 29044 2324 29084
rect 21004 28960 21044 29000
rect 18316 28876 18356 28916
rect 3688 28708 3728 28748
rect 3770 28708 3810 28748
rect 3852 28708 3892 28748
rect 3934 28708 3974 28748
rect 4016 28708 4056 28748
rect 6700 28708 6740 28748
rect 11500 28708 11540 28748
rect 18808 28708 18848 28748
rect 18890 28708 18930 28748
rect 18972 28708 19012 28748
rect 19054 28708 19094 28748
rect 19136 28708 19176 28748
rect 18412 28624 18452 28664
rect 7468 28456 7508 28496
rect 7756 28372 7796 28412
rect 15436 28456 15476 28496
rect 19276 28372 19316 28412
rect 17836 28288 17876 28328
rect 18028 28288 18068 28328
rect 18508 28288 18548 28328
rect 18124 28204 18164 28244
rect 18316 28204 18356 28244
rect 4928 27952 4968 27992
rect 5010 27952 5050 27992
rect 5092 27952 5132 27992
rect 5174 27952 5214 27992
rect 5256 27952 5296 27992
rect 20048 27952 20088 27992
rect 20130 27952 20170 27992
rect 20212 27952 20252 27992
rect 20294 27952 20334 27992
rect 20376 27952 20416 27992
rect 16684 27868 16724 27908
rect 6220 27784 6260 27824
rect 3148 27700 3188 27740
rect 7180 27700 7220 27740
rect 11020 27700 11060 27740
rect 19948 27700 19988 27740
rect 14572 27616 14612 27656
rect 3052 27532 3092 27572
rect 5356 27448 5396 27488
rect 17740 27448 17780 27488
rect 10156 27364 10196 27404
rect 3688 27196 3728 27236
rect 3770 27196 3810 27236
rect 3852 27196 3892 27236
rect 3934 27196 3974 27236
rect 4016 27196 4056 27236
rect 18808 27196 18848 27236
rect 18890 27196 18930 27236
rect 18972 27196 19012 27236
rect 19054 27196 19094 27236
rect 19136 27196 19176 27236
rect 13900 27028 13940 27068
rect 17644 26860 17684 26900
rect 10156 26776 10196 26816
rect 18220 26692 18260 26732
rect 6220 26524 6260 26564
rect 18604 26524 18644 26564
rect 4928 26440 4968 26480
rect 5010 26440 5050 26480
rect 5092 26440 5132 26480
rect 5174 26440 5214 26480
rect 5256 26440 5296 26480
rect 14668 26440 14708 26480
rect 20048 26440 20088 26480
rect 20130 26440 20170 26480
rect 20212 26440 20252 26480
rect 20294 26440 20334 26480
rect 20376 26440 20416 26480
rect 14572 26272 14612 26312
rect 14764 26272 14804 26312
rect 3244 26188 3284 26228
rect 4108 26188 4148 26228
rect 6700 26104 6740 26144
rect 13804 26104 13844 26144
rect 4300 26020 4340 26060
rect 5356 26020 5396 26060
rect 11884 26020 11924 26060
rect 17740 26020 17780 26060
rect 1612 25936 1652 25976
rect 3688 25684 3728 25724
rect 3770 25684 3810 25724
rect 3852 25684 3892 25724
rect 3934 25684 3974 25724
rect 4016 25684 4056 25724
rect 16492 25684 16532 25724
rect 18808 25684 18848 25724
rect 18890 25684 18930 25724
rect 18972 25684 19012 25724
rect 19054 25684 19094 25724
rect 19136 25684 19176 25724
rect 6220 25264 6260 25304
rect 6508 25264 6548 25304
rect 7948 25264 7988 25304
rect 16588 25264 16628 25304
rect 6028 25180 6068 25220
rect 14284 25180 14324 25220
rect 4928 24928 4968 24968
rect 5010 24928 5050 24968
rect 5092 24928 5132 24968
rect 5174 24928 5214 24968
rect 5256 24928 5296 24968
rect 6412 24928 6452 24968
rect 16492 24928 16532 24968
rect 20048 24928 20088 24968
rect 20130 24928 20170 24968
rect 20212 24928 20252 24968
rect 20294 24928 20334 24968
rect 20376 24928 20416 24968
rect 16588 24844 16628 24884
rect 2860 24760 2900 24800
rect 7852 24760 7892 24800
rect 17356 24760 17396 24800
rect 2956 24592 2996 24632
rect 3532 24592 3572 24632
rect 10156 24592 10196 24632
rect 11020 24592 11060 24632
rect 13804 24508 13844 24548
rect 5644 24424 5684 24464
rect 17068 24424 17108 24464
rect 10636 24256 10676 24296
rect 3688 24172 3728 24212
rect 3770 24172 3810 24212
rect 3852 24172 3892 24212
rect 3934 24172 3974 24212
rect 4016 24172 4056 24212
rect 18808 24172 18848 24212
rect 18890 24172 18930 24212
rect 18972 24172 19012 24212
rect 19054 24172 19094 24212
rect 19136 24172 19176 24212
rect 76 23920 116 23960
rect 11308 23920 11348 23960
rect 17644 23920 17684 23960
rect 19852 23920 19892 23960
rect 18316 23836 18356 23876
rect 5452 23752 5492 23792
rect 5740 23752 5780 23792
rect 8236 23752 8276 23792
rect 13900 23752 13940 23792
rect 17740 23752 17780 23792
rect 8620 23668 8660 23708
rect 11020 23668 11060 23708
rect 11308 23668 11348 23708
rect 17932 23668 17972 23708
rect 5548 23584 5588 23624
rect 8332 23584 8372 23624
rect 4684 23500 4724 23540
rect 4928 23416 4968 23456
rect 5010 23416 5050 23456
rect 5092 23416 5132 23456
rect 5174 23416 5214 23456
rect 5256 23416 5296 23456
rect 5452 23416 5492 23456
rect 6796 23332 6836 23372
rect 20048 23416 20088 23456
rect 20130 23416 20170 23456
rect 20212 23416 20252 23456
rect 20294 23416 20334 23456
rect 20376 23416 20416 23456
rect 172 23080 212 23120
rect 8716 23080 8756 23120
rect 4108 22996 4148 23036
rect 6316 22996 6356 23036
rect 7084 22996 7124 23036
rect 7180 22828 7220 22868
rect 5548 22744 5588 22784
rect 8332 22744 8372 22784
rect 3688 22660 3728 22700
rect 3770 22660 3810 22700
rect 3852 22660 3892 22700
rect 3934 22660 3974 22700
rect 4016 22660 4056 22700
rect 18808 22660 18848 22700
rect 18890 22660 18930 22700
rect 18972 22660 19012 22700
rect 19054 22660 19094 22700
rect 19136 22660 19176 22700
rect 10924 22324 10964 22364
rect 13804 22324 13844 22364
rect 11020 22240 11060 22280
rect 13036 22240 13076 22280
rect 14380 22240 14420 22280
rect 6508 22156 6548 22196
rect 7660 22156 7700 22196
rect 2860 22072 2900 22112
rect 7660 21988 7700 22028
rect 20620 21988 20660 22028
rect 4928 21904 4968 21944
rect 5010 21904 5050 21944
rect 5092 21904 5132 21944
rect 5174 21904 5214 21944
rect 5256 21904 5296 21944
rect 20048 21904 20088 21944
rect 20130 21904 20170 21944
rect 20212 21904 20252 21944
rect 20294 21904 20334 21944
rect 20376 21904 20416 21944
rect 2668 21568 2708 21608
rect 7948 21568 7988 21608
rect 13996 21568 14036 21608
rect 17452 21568 17492 21608
rect 6700 21484 6740 21524
rect 8524 21484 8564 21524
rect 3688 21148 3728 21188
rect 3770 21148 3810 21188
rect 3852 21148 3892 21188
rect 3934 21148 3974 21188
rect 4016 21148 4056 21188
rect 18808 21148 18848 21188
rect 18890 21148 18930 21188
rect 18972 21148 19012 21188
rect 19054 21148 19094 21188
rect 19136 21148 19176 21188
rect 7756 21064 7796 21104
rect 17836 20980 17876 21020
rect 18124 20980 18164 21020
rect 172 20896 212 20936
rect 6316 20896 6356 20936
rect 4684 20812 4724 20852
rect 12460 20812 12500 20852
rect 4108 20728 4148 20768
rect 5932 20728 5972 20768
rect 6412 20728 6452 20768
rect 6700 20728 6740 20768
rect 7852 20728 7892 20768
rect 12556 20728 12596 20768
rect 12748 20728 12788 20768
rect 14380 20728 14420 20768
rect 17644 20728 17684 20768
rect 4300 20644 4340 20684
rect 14284 20644 14324 20684
rect 17164 20644 17204 20684
rect 10252 20560 10292 20600
rect 556 20392 596 20432
rect 4928 20392 4968 20432
rect 5010 20392 5050 20432
rect 5092 20392 5132 20432
rect 5174 20392 5214 20432
rect 5256 20392 5296 20432
rect 20048 20392 20088 20432
rect 20130 20392 20170 20432
rect 20212 20392 20252 20432
rect 20294 20392 20334 20432
rect 20376 20392 20416 20432
rect 3436 20224 3476 20264
rect 2956 20140 2996 20180
rect 5356 20056 5396 20096
rect 8620 20056 8660 20096
rect 19660 20056 19700 20096
rect 16588 19972 16628 20012
rect 11884 19888 11924 19928
rect 3148 19804 3188 19844
rect 7180 19804 7220 19844
rect 13996 19804 14036 19844
rect 3436 19720 3476 19760
rect 3688 19636 3728 19676
rect 3770 19636 3810 19676
rect 3852 19636 3892 19676
rect 3934 19636 3974 19676
rect 4016 19636 4056 19676
rect 13420 19636 13460 19676
rect 18808 19636 18848 19676
rect 18890 19636 18930 19676
rect 18972 19636 19012 19676
rect 19054 19636 19094 19676
rect 19136 19636 19176 19676
rect 7180 19552 7220 19592
rect 2668 19468 2708 19508
rect 13420 19384 13460 19424
rect 13900 19384 13940 19424
rect 14284 19384 14324 19424
rect 12844 19216 12884 19256
rect 17932 19216 17972 19256
rect 7852 19048 7892 19088
rect 8812 19048 8852 19088
rect 15724 18964 15764 19004
rect 1228 18880 1268 18920
rect 4928 18880 4968 18920
rect 5010 18880 5050 18920
rect 5092 18880 5132 18920
rect 5174 18880 5214 18920
rect 5256 18880 5296 18920
rect 6220 18880 6260 18920
rect 20048 18880 20088 18920
rect 20130 18880 20170 18920
rect 20212 18880 20252 18920
rect 20294 18880 20334 18920
rect 20376 18880 20416 18920
rect 19276 18796 19316 18836
rect 4204 18712 4244 18752
rect 11980 18712 12020 18752
rect 17068 18712 17108 18752
rect 3244 18628 3284 18668
rect 17164 18628 17204 18668
rect 17548 18544 17588 18584
rect 18604 18544 18644 18584
rect 18316 18460 18356 18500
rect 14764 18376 14804 18416
rect 6028 18292 6068 18332
rect 17356 18292 17396 18332
rect 16108 18208 16148 18248
rect 3688 18124 3728 18164
rect 3770 18124 3810 18164
rect 3852 18124 3892 18164
rect 3934 18124 3974 18164
rect 4016 18124 4056 18164
rect 9196 18124 9236 18164
rect 18808 18124 18848 18164
rect 18890 18124 18930 18164
rect 18972 18124 19012 18164
rect 19054 18124 19094 18164
rect 19136 18124 19176 18164
rect 13804 17956 13844 17996
rect 18604 17956 18644 17996
rect 8236 17872 8276 17912
rect 19276 17872 19316 17912
rect 4108 17788 4148 17828
rect 8140 17788 8180 17828
rect 14764 17788 14804 17828
rect 19660 17788 19700 17828
rect 10252 17704 10292 17744
rect 12268 17704 12308 17744
rect 16780 17704 16820 17744
rect 7948 17620 7988 17660
rect 19660 17620 19700 17660
rect 19468 17536 19508 17576
rect 14668 17452 14708 17492
rect 4204 17368 4244 17408
rect 4928 17368 4968 17408
rect 5010 17368 5050 17408
rect 5092 17368 5132 17408
rect 5174 17368 5214 17408
rect 5256 17368 5296 17408
rect 20048 17368 20088 17408
rect 20130 17368 20170 17408
rect 20212 17368 20252 17408
rect 20294 17368 20334 17408
rect 20376 17368 20416 17408
rect 17836 17284 17876 17324
rect 14572 17116 14612 17156
rect 18412 17116 18452 17156
rect 18220 16948 18260 16988
rect 11788 16864 11828 16904
rect 18604 16780 18644 16820
rect 3688 16612 3728 16652
rect 3770 16612 3810 16652
rect 3852 16612 3892 16652
rect 3934 16612 3974 16652
rect 4016 16612 4056 16652
rect 10924 16612 10964 16652
rect 16588 16612 16628 16652
rect 18412 16612 18452 16652
rect 18808 16612 18848 16652
rect 18890 16612 18930 16652
rect 18972 16612 19012 16652
rect 19054 16612 19094 16652
rect 19136 16612 19176 16652
rect 19276 16528 19316 16568
rect 4204 16444 4244 16484
rect 4684 16444 4724 16484
rect 940 16360 980 16400
rect 3436 16360 3476 16400
rect 13228 16360 13268 16400
rect 17068 16360 17108 16400
rect 9484 16276 9524 16316
rect 4204 16192 4244 16232
rect 5068 16108 5108 16148
rect 5740 16108 5780 16148
rect 5740 15940 5780 15980
rect 4928 15856 4968 15896
rect 5010 15856 5050 15896
rect 5092 15856 5132 15896
rect 5174 15856 5214 15896
rect 5256 15856 5296 15896
rect 18604 15856 18644 15896
rect 20048 15856 20088 15896
rect 20130 15856 20170 15896
rect 20212 15856 20252 15896
rect 20294 15856 20334 15896
rect 20376 15856 20416 15896
rect 11308 15772 11348 15812
rect 7948 15688 7988 15728
rect 20716 15604 20756 15644
rect 4108 15520 4148 15560
rect 4300 15352 4340 15392
rect 9388 15268 9428 15308
rect 20812 15184 20852 15224
rect 3244 15100 3284 15140
rect 3688 15100 3728 15140
rect 3770 15100 3810 15140
rect 3852 15100 3892 15140
rect 3934 15100 3974 15140
rect 4016 15100 4056 15140
rect 8044 15100 8084 15140
rect 11020 15100 11060 15140
rect 12556 15100 12596 15140
rect 13900 15100 13940 15140
rect 16300 15100 16340 15140
rect 18808 15100 18848 15140
rect 18890 15100 18930 15140
rect 18972 15100 19012 15140
rect 19054 15100 19094 15140
rect 19136 15100 19176 15140
rect 11308 14932 11348 14972
rect 17644 14848 17684 14888
rect 16492 14764 16532 14804
rect 18412 14764 18452 14804
rect 19468 14680 19508 14720
rect 16684 14596 16724 14636
rect 3436 14344 3476 14384
rect 4928 14344 4968 14384
rect 5010 14344 5050 14384
rect 5092 14344 5132 14384
rect 5174 14344 5214 14384
rect 5256 14344 5296 14384
rect 20048 14344 20088 14384
rect 20130 14344 20170 14384
rect 20212 14344 20252 14384
rect 20294 14344 20334 14384
rect 20376 14344 20416 14384
rect 6508 14260 6548 14300
rect 13900 14260 13940 14300
rect 14956 14260 14996 14300
rect 7276 14176 7316 14216
rect 8812 14176 8852 14216
rect 14668 14176 14708 14216
rect 7084 14092 7124 14132
rect 11692 14092 11732 14132
rect 3052 14008 3092 14048
rect 5932 14008 5972 14048
rect 2860 13924 2900 13964
rect 8524 13924 8564 13964
rect 16684 13924 16724 13964
rect 12172 13840 12212 13880
rect 14764 13840 14804 13880
rect 15628 13840 15668 13880
rect 15724 13756 15764 13796
rect 3052 13672 3092 13712
rect 9196 13672 9236 13712
rect 3688 13588 3728 13628
rect 3770 13588 3810 13628
rect 3852 13588 3892 13628
rect 3934 13588 3974 13628
rect 4016 13588 4056 13628
rect 6508 13588 6548 13628
rect 8620 13588 8660 13628
rect 18808 13588 18848 13628
rect 18890 13588 18930 13628
rect 18972 13588 19012 13628
rect 19054 13588 19094 13628
rect 19136 13588 19176 13628
rect 10540 13504 10580 13544
rect 17836 13504 17876 13544
rect 748 13420 788 13460
rect 11308 13336 11348 13376
rect 1420 13252 1460 13292
rect 9484 13168 9524 13208
rect 16492 13084 16532 13124
rect 7564 13000 7604 13040
rect 4928 12832 4968 12872
rect 5010 12832 5050 12872
rect 5092 12832 5132 12872
rect 5174 12832 5214 12872
rect 5256 12832 5296 12872
rect 12172 12832 12212 12872
rect 20048 12832 20088 12872
rect 20130 12832 20170 12872
rect 20212 12832 20252 12872
rect 20294 12832 20334 12872
rect 20376 12832 20416 12872
rect 18508 12664 18548 12704
rect 3148 12580 3188 12620
rect 12172 12580 12212 12620
rect 13132 12580 13172 12620
rect 14668 12580 14708 12620
rect 18316 12580 18356 12620
rect 3436 12496 3476 12536
rect 16492 12496 16532 12536
rect 8044 12412 8084 12452
rect 1228 12328 1268 12368
rect 8620 12160 8660 12200
rect 15724 12160 15764 12200
rect 16108 12160 16148 12200
rect 17740 12160 17780 12200
rect 3244 12076 3284 12116
rect 3688 12076 3728 12116
rect 3770 12076 3810 12116
rect 3852 12076 3892 12116
rect 3934 12076 3974 12116
rect 4016 12076 4056 12116
rect 7948 12076 7988 12116
rect 17836 12076 17876 12116
rect 18808 12076 18848 12116
rect 18890 12076 18930 12116
rect 18972 12076 19012 12116
rect 19054 12076 19094 12116
rect 19136 12076 19176 12116
rect 5740 11908 5780 11948
rect 7468 11824 7508 11864
rect 4108 11572 4148 11612
rect 5644 11488 5684 11528
rect 17836 11656 17876 11696
rect 18508 11656 18548 11696
rect 12076 11572 12116 11612
rect 12844 11572 12884 11612
rect 13132 11572 13172 11612
rect 16588 11488 16628 11528
rect 8332 11404 8372 11444
rect 4588 11320 4628 11360
rect 4928 11320 4968 11360
rect 5010 11320 5050 11360
rect 5092 11320 5132 11360
rect 5174 11320 5214 11360
rect 5256 11320 5296 11360
rect 9196 11320 9236 11360
rect 18508 11404 18548 11444
rect 20048 11320 20088 11360
rect 20130 11320 20170 11360
rect 20212 11320 20252 11360
rect 20294 11320 20334 11360
rect 20376 11320 20416 11360
rect 8812 11152 8852 11192
rect 12076 11152 12116 11192
rect 17932 11152 17972 11192
rect 8332 11068 8372 11108
rect 17740 11068 17780 11108
rect 9388 10984 9428 11024
rect 17452 10900 17492 10940
rect 12460 10816 12500 10856
rect 12844 10816 12884 10856
rect 3244 10732 3284 10772
rect 4780 10732 4820 10772
rect 18220 10732 18260 10772
rect 11308 10648 11348 10688
rect 19756 10648 19796 10688
rect 3688 10564 3728 10604
rect 3770 10564 3810 10604
rect 3852 10564 3892 10604
rect 3934 10564 3974 10604
rect 4016 10564 4056 10604
rect 18808 10564 18848 10604
rect 18890 10564 18930 10604
rect 18972 10564 19012 10604
rect 19054 10564 19094 10604
rect 19136 10564 19176 10604
rect 9484 10480 9524 10520
rect 10636 10480 10676 10520
rect 20716 10480 20756 10520
rect 9100 10396 9140 10436
rect 18124 10312 18164 10352
rect 18412 10312 18452 10352
rect 9388 10228 9428 10268
rect 4108 10144 4148 10184
rect 10060 10144 10100 10184
rect 17164 10144 17204 10184
rect 3052 9976 3092 10016
rect 6700 9892 6740 9932
rect 4928 9808 4968 9848
rect 5010 9808 5050 9848
rect 5092 9808 5132 9848
rect 5174 9808 5214 9848
rect 5256 9808 5296 9848
rect 9100 9808 9140 9848
rect 12748 9808 12788 9848
rect 20048 9808 20088 9848
rect 20130 9808 20170 9848
rect 20212 9808 20252 9848
rect 20294 9808 20334 9848
rect 20376 9808 20416 9848
rect 844 9640 884 9680
rect 9196 9640 9236 9680
rect 9484 9640 9524 9680
rect 7660 9556 7700 9596
rect 17740 9472 17780 9512
rect 3628 9388 3668 9428
rect 4204 9388 4244 9428
rect 10540 9388 10580 9428
rect 13228 9388 13268 9428
rect 14668 9388 14708 9428
rect 18412 9388 18452 9428
rect 10924 9304 10964 9344
rect 11788 9304 11828 9344
rect 17644 9304 17684 9344
rect 3148 9220 3188 9260
rect 9580 9220 9620 9260
rect 10156 9220 10196 9260
rect 10540 9220 10580 9260
rect 18604 9220 18644 9260
rect 4588 9136 4628 9176
rect 3688 9052 3728 9092
rect 3770 9052 3810 9092
rect 3852 9052 3892 9092
rect 3934 9052 3974 9092
rect 4016 9052 4056 9092
rect 7564 9052 7604 9092
rect 11884 9052 11924 9092
rect 18808 9052 18848 9092
rect 18890 9052 18930 9092
rect 18972 9052 19012 9092
rect 19054 9052 19094 9092
rect 19136 9052 19176 9092
rect 14284 8968 14324 9008
rect 8812 8800 8852 8840
rect 4204 8716 4244 8756
rect 10060 8632 10100 8672
rect 12268 8632 12308 8672
rect 18316 8548 18356 8588
rect 16972 8464 17012 8504
rect 4928 8296 4968 8336
rect 5010 8296 5050 8336
rect 5092 8296 5132 8336
rect 5174 8296 5214 8336
rect 5256 8296 5296 8336
rect 18124 8296 18164 8336
rect 20048 8296 20088 8336
rect 20130 8296 20170 8336
rect 20212 8296 20252 8336
rect 20294 8296 20334 8336
rect 20376 8296 20416 8336
rect 2956 8044 2996 8084
rect 6508 8128 6548 8168
rect 3436 7792 3476 7832
rect 7468 7792 7508 7832
rect 16204 7792 16244 7832
rect 10444 7708 10484 7748
rect 16780 7708 16820 7748
rect 16972 7708 17012 7748
rect 19084 7708 19124 7748
rect 17068 7624 17108 7664
rect 3688 7540 3728 7580
rect 3770 7540 3810 7580
rect 3852 7540 3892 7580
rect 3934 7540 3974 7580
rect 4016 7540 4056 7580
rect 4780 7540 4820 7580
rect 18808 7540 18848 7580
rect 18890 7540 18930 7580
rect 18972 7540 19012 7580
rect 19054 7540 19094 7580
rect 19136 7540 19176 7580
rect 1324 7372 1364 7412
rect 16396 7120 16436 7160
rect 3340 7036 3380 7076
rect 3724 7036 3764 7076
rect 13420 6952 13460 6992
rect 17164 6952 17204 6992
rect 2668 6868 2708 6908
rect 10252 6868 10292 6908
rect 13228 6868 13268 6908
rect 4928 6784 4968 6824
rect 5010 6784 5050 6824
rect 5092 6784 5132 6824
rect 5174 6784 5214 6824
rect 5256 6784 5296 6824
rect 11404 6784 11444 6824
rect 20048 6784 20088 6824
rect 20130 6784 20170 6824
rect 20212 6784 20252 6824
rect 20294 6784 20334 6824
rect 20376 6784 20416 6824
rect 17452 6700 17492 6740
rect 3724 6616 3764 6656
rect 5644 6448 5684 6488
rect 2668 6196 2708 6236
rect 17932 6196 17972 6236
rect 18508 6112 18548 6152
rect 3688 6028 3728 6068
rect 3770 6028 3810 6068
rect 3852 6028 3892 6068
rect 3934 6028 3974 6068
rect 4016 6028 4056 6068
rect 12268 6028 12308 6068
rect 18316 6028 18356 6068
rect 18808 6028 18848 6068
rect 18890 6028 18930 6068
rect 18972 6028 19012 6068
rect 19054 6028 19094 6068
rect 19136 6028 19176 6068
rect 17644 5944 17684 5984
rect 18412 5944 18452 5984
rect 4780 5776 4820 5816
rect 15628 5776 15668 5816
rect 3436 5692 3476 5732
rect 4684 5692 4724 5732
rect 7084 5356 7124 5396
rect 4928 5272 4968 5312
rect 5010 5272 5050 5312
rect 5092 5272 5132 5312
rect 5174 5272 5214 5312
rect 5256 5272 5296 5312
rect 20048 5272 20088 5312
rect 20130 5272 20170 5312
rect 20212 5272 20252 5312
rect 20294 5272 20334 5312
rect 20376 5272 20416 5312
rect 12652 5188 12692 5228
rect 12556 5104 12596 5144
rect 4684 5020 4724 5060
rect 6796 4936 6836 4976
rect 7180 4936 7220 4976
rect 16588 5020 16628 5060
rect 13516 4936 13556 4976
rect 13804 4936 13844 4976
rect 17452 4936 17492 4976
rect 17740 4936 17780 4976
rect 2860 4852 2900 4892
rect 18028 4852 18068 4892
rect 1228 4768 1268 4808
rect 5548 4684 5588 4724
rect 3688 4516 3728 4556
rect 3770 4516 3810 4556
rect 3852 4516 3892 4556
rect 3934 4516 3974 4556
rect 4016 4516 4056 4556
rect 18808 4516 18848 4556
rect 18890 4516 18930 4556
rect 18972 4516 19012 4556
rect 19054 4516 19094 4556
rect 19136 4516 19176 4556
rect 19372 4516 19412 4556
rect 2860 4432 2900 4472
rect 7468 4432 7508 4472
rect 11596 4432 11636 4472
rect 17644 4432 17684 4472
rect 19372 4348 19412 4388
rect 4492 4264 4532 4304
rect 5932 4180 5972 4220
rect 16684 4264 16724 4304
rect 5740 4096 5780 4136
rect 16588 4096 16628 4136
rect 16972 4096 17012 4136
rect 17164 4096 17204 4136
rect 4928 3760 4968 3800
rect 5010 3760 5050 3800
rect 5092 3760 5132 3800
rect 5174 3760 5214 3800
rect 5256 3760 5296 3800
rect 7660 3760 7700 3800
rect 16588 3760 16628 3800
rect 18316 3760 18356 3800
rect 20048 3760 20088 3800
rect 20130 3760 20170 3800
rect 20212 3760 20252 3800
rect 20294 3760 20334 3800
rect 20376 3760 20416 3800
rect 6892 3676 6932 3716
rect 7276 3676 7316 3716
rect 8524 3592 8564 3632
rect 13324 3592 13364 3632
rect 76 3508 116 3548
rect 7276 3508 7316 3548
rect 7564 3508 7604 3548
rect 9004 3508 9044 3548
rect 4204 3424 4244 3464
rect 7084 3424 7124 3464
rect 18220 3424 18260 3464
rect 3916 3340 3956 3380
rect 17644 3340 17684 3380
rect 18028 3256 18068 3296
rect 3688 3004 3728 3044
rect 3770 3004 3810 3044
rect 3852 3004 3892 3044
rect 3934 3004 3974 3044
rect 4016 3004 4056 3044
rect 17932 3088 17972 3128
rect 20812 3088 20852 3128
rect 18808 3004 18848 3044
rect 18890 3004 18930 3044
rect 18972 3004 19012 3044
rect 19054 3004 19094 3044
rect 19136 3004 19176 3044
rect 16300 2752 16340 2792
rect 6700 2668 6740 2708
rect 7468 2668 7508 2708
rect 14188 2668 14228 2708
rect 17452 2668 17492 2708
rect 16300 2584 16340 2624
rect 17164 2584 17204 2624
rect 7660 2332 7700 2372
rect 7852 2332 7892 2372
rect 8620 2332 8660 2372
rect 16588 2500 16628 2540
rect 16684 2416 16724 2456
rect 16204 2332 16244 2372
rect 4928 2248 4968 2288
rect 5010 2248 5050 2288
rect 5092 2248 5132 2288
rect 5174 2248 5214 2288
rect 5256 2248 5296 2288
rect 13900 2248 13940 2288
rect 20048 2248 20088 2288
rect 20130 2248 20170 2288
rect 20212 2248 20252 2288
rect 20294 2248 20334 2288
rect 20376 2248 20416 2288
rect 8524 2164 8564 2204
rect 7564 2080 7604 2120
rect 18124 1996 18164 2036
rect 5548 1912 5588 1952
rect 2284 1828 2324 1868
rect 8620 1828 8660 1868
rect 10348 1828 10388 1868
rect 10828 1828 10868 1868
rect 11116 1828 11156 1868
rect 7468 1744 7508 1784
rect 8524 1744 8564 1784
rect 20908 1744 20948 1784
rect 13228 1660 13268 1700
rect 15052 1576 15092 1616
rect 3688 1492 3728 1532
rect 3770 1492 3810 1532
rect 3852 1492 3892 1532
rect 3934 1492 3974 1532
rect 4016 1492 4056 1532
rect 18808 1492 18848 1532
rect 18890 1492 18930 1532
rect 18972 1492 19012 1532
rect 19054 1492 19094 1532
rect 19136 1492 19176 1532
rect 13708 1408 13748 1448
rect 3340 1240 3380 1280
rect 3532 1240 3572 1280
rect 5452 1240 5492 1280
rect 6604 1240 6644 1280
rect 7756 1240 7796 1280
rect 9292 1240 9332 1280
rect 14092 1240 14132 1280
rect 16780 1240 16820 1280
rect 17548 1240 17588 1280
rect 18700 1240 18740 1280
rect 19468 1240 19508 1280
rect 652 1156 692 1196
rect 7180 1156 7220 1196
rect 8044 1156 8084 1196
rect 9580 1156 9620 1196
rect 10060 1156 10100 1196
rect 4780 1072 4820 1112
rect 14476 1072 14516 1112
rect 1132 988 1172 1028
rect 10828 988 10868 1028
rect 11212 988 11252 1028
rect 13516 988 13556 1028
rect 17836 988 17876 1028
rect 2764 904 2804 944
rect 4108 904 4148 944
rect 4780 904 4820 944
rect 7948 904 7988 944
rect 15916 904 15956 944
rect 18124 904 18164 944
rect 19276 904 19316 944
rect 14284 820 14324 860
rect 16876 820 16916 860
rect 17932 820 17972 860
rect 2572 736 2612 776
rect 4928 736 4968 776
rect 5010 736 5050 776
rect 5092 736 5132 776
rect 5174 736 5214 776
rect 5256 736 5296 776
rect 6988 736 7028 776
rect 13708 736 13748 776
rect 20048 736 20088 776
rect 20130 736 20170 776
rect 20212 736 20252 776
rect 20294 736 20334 776
rect 20376 736 20416 776
rect 5932 652 5972 692
rect 1036 568 1076 608
rect 4684 568 4724 608
rect 5356 568 5396 608
rect 6508 652 6548 692
rect 7948 568 7988 608
rect 8140 568 8180 608
rect 15436 568 15476 608
rect 17068 568 17108 608
rect 2476 484 2516 524
rect 7372 484 7412 524
rect 14860 484 14900 524
rect 6412 400 6452 440
rect 15244 400 15284 440
rect 2380 316 2420 356
rect 6892 316 6932 356
rect 14092 316 14132 356
rect 2188 232 2228 272
rect 12172 232 12212 272
rect 15724 232 15764 272
rect 13612 148 13652 188
rect 17260 232 17300 272
rect 7948 64 7988 104
rect 10828 64 10868 104
rect 17164 64 17204 104
<< metal4 >>
rect 20620 42776 20660 42785
rect 4108 42608 4148 42617
rect 1900 42272 1940 42281
rect 1516 42104 1556 42113
rect 1420 38996 1460 39005
rect 652 37400 692 37409
rect 172 37064 212 37073
rect 76 23960 116 23969
rect 76 3548 116 23920
rect 172 23120 212 37024
rect 172 23071 212 23080
rect 172 20936 212 20945
rect 172 7757 212 20896
rect 556 20432 596 20441
rect 459 20012 501 20021
rect 459 19972 460 20012
rect 500 19972 501 20012
rect 459 19963 501 19972
rect 460 16157 500 19963
rect 556 16325 596 20392
rect 555 16316 597 16325
rect 555 16276 556 16316
rect 596 16276 597 16316
rect 555 16267 597 16276
rect 459 16148 501 16157
rect 459 16108 460 16148
rect 500 16108 501 16148
rect 459 16099 501 16108
rect 171 7748 213 7757
rect 171 7708 172 7748
rect 212 7708 213 7748
rect 171 7699 213 7708
rect 76 3499 116 3508
rect 652 1196 692 37360
rect 1228 37316 1268 37325
rect 940 36476 980 36485
rect 748 35132 788 35141
rect 748 20021 788 35092
rect 844 33620 884 33629
rect 747 20012 789 20021
rect 747 19972 748 20012
rect 788 19972 789 20012
rect 747 19963 789 19972
rect 844 19508 884 33580
rect 748 19468 884 19508
rect 748 13460 788 19468
rect 940 19424 980 36436
rect 1132 34880 1172 34889
rect 1132 34376 1172 34840
rect 748 13411 788 13420
rect 844 19384 980 19424
rect 1036 33956 1076 33965
rect 844 9680 884 19384
rect 844 9631 884 9640
rect 940 16400 980 16409
rect 940 7001 980 16360
rect 939 6992 981 7001
rect 939 6952 940 6992
rect 980 6952 981 6992
rect 939 6943 981 6952
rect 652 1147 692 1156
rect 1036 608 1076 33916
rect 1132 30512 1172 34336
rect 1132 30463 1172 30472
rect 1228 20180 1268 37276
rect 1132 20140 1268 20180
rect 1324 32948 1364 32957
rect 1132 1028 1172 20140
rect 1227 19088 1269 19097
rect 1227 19048 1228 19088
rect 1268 19048 1269 19088
rect 1227 19039 1269 19048
rect 1228 18920 1268 19039
rect 1228 18871 1268 18880
rect 1227 12368 1269 12377
rect 1227 12328 1228 12368
rect 1268 12328 1269 12368
rect 1227 12319 1269 12328
rect 1228 12234 1268 12319
rect 1324 7412 1364 32908
rect 1420 13292 1460 38956
rect 1516 33200 1556 42064
rect 1804 41264 1844 41273
rect 1516 33151 1556 33160
rect 1612 39752 1652 39761
rect 1612 25976 1652 39712
rect 1708 38912 1748 38921
rect 1708 30260 1748 38872
rect 1804 38072 1844 41224
rect 1804 37820 1844 38032
rect 1804 32864 1844 37780
rect 1900 33200 1940 42232
rect 2764 41264 2804 41273
rect 2476 39584 2516 39593
rect 2092 38660 2132 38669
rect 1900 33151 1940 33160
rect 1996 37232 2036 37241
rect 1804 32815 1844 32824
rect 1708 29504 1748 30220
rect 1708 29455 1748 29464
rect 1612 25927 1652 25936
rect 1420 13243 1460 13252
rect 1324 7363 1364 7372
rect 1227 4808 1269 4817
rect 1227 4768 1228 4808
rect 1268 4768 1269 4808
rect 1227 4759 1269 4768
rect 1228 4674 1268 4759
rect 1132 979 1172 988
rect 1036 559 1076 568
rect 1996 449 2036 37192
rect 2092 34544 2132 38620
rect 2476 37736 2516 39544
rect 2571 38072 2613 38081
rect 2571 38032 2572 38072
rect 2612 38032 2613 38072
rect 2571 38023 2613 38032
rect 2572 37904 2612 38023
rect 2572 37855 2612 37864
rect 2764 37820 2804 41224
rect 3052 40844 3092 40853
rect 3052 40256 3092 40804
rect 3688 40844 4056 40853
rect 3728 40804 3770 40844
rect 3810 40804 3852 40844
rect 3892 40804 3934 40844
rect 3974 40804 4016 40844
rect 3688 40795 4056 40804
rect 3052 40207 3092 40216
rect 3340 40592 3380 40601
rect 3148 40088 3188 40097
rect 2955 38072 2997 38081
rect 2955 38032 2956 38072
rect 2996 38032 2997 38072
rect 2955 38023 2997 38032
rect 2764 37780 2900 37820
rect 2476 37687 2516 37696
rect 2476 37568 2516 37577
rect 2380 37528 2476 37568
rect 2380 37400 2420 37528
rect 2476 37519 2516 37528
rect 2764 37484 2804 37493
rect 2380 37351 2420 37360
rect 2572 37400 2612 37409
rect 2476 36896 2516 36905
rect 2284 36856 2476 36896
rect 2284 36812 2324 36856
rect 2476 36847 2516 36856
rect 2284 36763 2324 36772
rect 2092 34495 2132 34504
rect 2188 35720 2228 35729
rect 1995 440 2037 449
rect 1995 400 1996 440
rect 2036 400 2037 440
rect 1995 391 2037 400
rect 2188 272 2228 35680
rect 2572 35216 2612 37360
rect 2572 35167 2612 35176
rect 2764 35216 2804 37444
rect 2668 34628 2708 34637
rect 2476 33956 2516 33965
rect 2476 33452 2516 33916
rect 2476 33403 2516 33412
rect 2572 32948 2612 32957
rect 2476 32276 2516 32285
rect 2380 31520 2420 31529
rect 2284 29084 2324 29093
rect 2284 1868 2324 29044
rect 2284 1819 2324 1828
rect 2380 356 2420 31480
rect 2476 524 2516 32236
rect 2572 776 2612 32908
rect 2668 31352 2708 34588
rect 2668 29840 2708 31312
rect 2668 29791 2708 29800
rect 2668 21608 2708 21617
rect 2668 19508 2708 21568
rect 2668 19459 2708 19468
rect 2668 6908 2708 6917
rect 2668 6236 2708 6868
rect 2668 6187 2708 6196
rect 2764 944 2804 35176
rect 2860 33536 2900 37780
rect 2860 33487 2900 33496
rect 2860 24800 2900 24809
rect 2860 22112 2900 24760
rect 2956 24632 2996 38023
rect 3148 34712 3188 40048
rect 3340 38249 3380 40552
rect 3688 39332 4056 39341
rect 3728 39292 3770 39332
rect 3810 39292 3852 39332
rect 3892 39292 3934 39332
rect 3974 39292 4016 39332
rect 3688 39283 4056 39292
rect 3339 38240 3381 38249
rect 3339 38200 3340 38240
rect 3380 38200 3381 38240
rect 3339 38191 3381 38200
rect 3148 27740 3188 34672
rect 3148 27691 3188 27700
rect 2956 24583 2996 24592
rect 3052 27572 3092 27581
rect 2860 22063 2900 22072
rect 2956 20180 2996 20189
rect 2860 13964 2900 13973
rect 2860 4892 2900 13924
rect 2956 8084 2996 20140
rect 3052 14048 3092 27532
rect 3244 26228 3284 26237
rect 3052 13999 3092 14008
rect 3148 19844 3188 19853
rect 3052 13712 3092 13721
rect 3052 10016 3092 13672
rect 3148 12620 3188 19804
rect 3244 18668 3284 26188
rect 3244 18619 3284 18628
rect 3148 12571 3188 12580
rect 3244 15140 3284 15149
rect 3244 12452 3284 15100
rect 3052 9967 3092 9976
rect 3148 12412 3284 12452
rect 3148 9260 3188 12412
rect 3244 12116 3284 12125
rect 3244 10772 3284 12076
rect 3244 10723 3284 10732
rect 3148 9211 3188 9220
rect 3340 8252 3380 38191
rect 3688 37820 4056 37829
rect 3728 37780 3770 37820
rect 3810 37780 3852 37820
rect 3892 37780 3934 37820
rect 3974 37780 4016 37820
rect 3688 37771 4056 37780
rect 3532 36896 3572 36905
rect 3532 36056 3572 36856
rect 3688 36308 4056 36317
rect 3728 36268 3770 36308
rect 3810 36268 3852 36308
rect 3892 36268 3934 36308
rect 3974 36268 4016 36308
rect 3688 36259 4056 36268
rect 4108 36140 4148 42568
rect 11788 42608 11828 42617
rect 4928 41600 5296 41609
rect 4968 41560 5010 41600
rect 5050 41560 5092 41600
rect 5132 41560 5174 41600
rect 5214 41560 5256 41600
rect 4928 41551 5296 41560
rect 9868 41600 9908 41609
rect 8044 41180 8084 41189
rect 4204 40844 4244 40853
rect 4204 37988 4244 40804
rect 5836 40424 5876 40433
rect 4928 40088 5296 40097
rect 4968 40048 5010 40088
rect 5050 40048 5092 40088
rect 5132 40048 5174 40088
rect 5214 40048 5256 40088
rect 4928 40039 5296 40048
rect 4928 38576 5296 38585
rect 4968 38536 5010 38576
rect 5050 38536 5092 38576
rect 5132 38536 5174 38576
rect 5214 38536 5256 38576
rect 4928 38527 5296 38536
rect 4204 37939 4244 37948
rect 4108 36091 4148 36100
rect 4204 37400 4244 37409
rect 3532 36007 3572 36016
rect 4204 35300 4244 37360
rect 4928 37064 5296 37073
rect 4968 37024 5010 37064
rect 5050 37024 5092 37064
rect 5132 37024 5174 37064
rect 5214 37024 5256 37064
rect 4928 37015 5296 37024
rect 5836 36728 5876 40384
rect 7372 38156 7412 38165
rect 5836 36679 5876 36688
rect 6892 37232 6932 37241
rect 6700 36560 6740 36569
rect 6604 35888 6644 35897
rect 4492 35720 4532 35729
rect 4204 35260 4340 35300
rect 3688 34796 4056 34805
rect 3728 34756 3770 34796
rect 3810 34756 3852 34796
rect 3892 34756 3934 34796
rect 3974 34756 4016 34796
rect 3688 34747 4056 34756
rect 3688 33284 4056 33293
rect 3728 33244 3770 33284
rect 3810 33244 3852 33284
rect 3892 33244 3934 33284
rect 3974 33244 4016 33284
rect 3688 33235 4056 33244
rect 3723 32948 3765 32957
rect 3723 32908 3724 32948
rect 3764 32908 3765 32948
rect 3723 32899 3765 32908
rect 3724 32814 3764 32899
rect 4204 32864 4244 32873
rect 3688 31772 4056 31781
rect 3728 31732 3770 31772
rect 3810 31732 3852 31772
rect 3892 31732 3934 31772
rect 3974 31732 4016 31772
rect 3688 31723 4056 31732
rect 3688 30260 4056 30269
rect 3728 30220 3770 30260
rect 3810 30220 3852 30260
rect 3892 30220 3934 30260
rect 3974 30220 4016 30260
rect 3688 30211 4056 30220
rect 3688 28748 4056 28757
rect 3728 28708 3770 28748
rect 3810 28708 3852 28748
rect 3892 28708 3934 28748
rect 3974 28708 4016 28748
rect 3688 28699 4056 28708
rect 3688 27236 4056 27245
rect 3728 27196 3770 27236
rect 3810 27196 3852 27236
rect 3892 27196 3934 27236
rect 3974 27196 4016 27236
rect 3688 27187 4056 27196
rect 4108 26228 4148 26237
rect 3688 25724 4056 25733
rect 3728 25684 3770 25724
rect 3810 25684 3852 25724
rect 3892 25684 3934 25724
rect 3974 25684 4016 25724
rect 3688 25675 4056 25684
rect 3532 24632 3572 24641
rect 3436 20264 3476 20273
rect 3436 19760 3476 20224
rect 3436 19711 3476 19720
rect 3436 16400 3476 16409
rect 3436 14384 3476 16360
rect 3436 14335 3476 14344
rect 2956 8035 2996 8044
rect 3148 8212 3380 8252
rect 3436 12536 3476 12545
rect 2860 4472 2900 4852
rect 2860 4423 2900 4432
rect 3148 2540 3188 8212
rect 3436 8084 3476 12496
rect 3340 8044 3476 8084
rect 3340 7076 3380 8044
rect 3340 7027 3380 7036
rect 3436 7832 3476 7841
rect 3436 5732 3476 7792
rect 3436 5683 3476 5692
rect 3148 2500 3380 2540
rect 3340 1280 3380 2500
rect 3340 1231 3380 1240
rect 3532 1280 3572 24592
rect 3688 24212 4056 24221
rect 3728 24172 3770 24212
rect 3810 24172 3852 24212
rect 3892 24172 3934 24212
rect 3974 24172 4016 24212
rect 3688 24163 4056 24172
rect 4108 23036 4148 26188
rect 3688 22700 4056 22709
rect 3728 22660 3770 22700
rect 3810 22660 3852 22700
rect 3892 22660 3934 22700
rect 3974 22660 4016 22700
rect 3688 22651 4056 22660
rect 3688 21188 4056 21197
rect 3728 21148 3770 21188
rect 3810 21148 3852 21188
rect 3892 21148 3934 21188
rect 3974 21148 4016 21188
rect 3688 21139 4056 21148
rect 4108 20768 4148 22996
rect 4108 20719 4148 20728
rect 3688 19676 4056 19685
rect 3728 19636 3770 19676
rect 3810 19636 3852 19676
rect 3892 19636 3934 19676
rect 3974 19636 4016 19676
rect 3688 19627 4056 19636
rect 4204 18752 4244 32824
rect 4300 32780 4340 35260
rect 4300 32731 4340 32740
rect 4300 26060 4340 26069
rect 4300 20684 4340 26020
rect 4300 20635 4340 20644
rect 4204 18703 4244 18712
rect 3688 18164 4056 18173
rect 3728 18124 3770 18164
rect 3810 18124 3852 18164
rect 3892 18124 3934 18164
rect 3974 18124 4016 18164
rect 3688 18115 4056 18124
rect 4108 17828 4148 17837
rect 3688 16652 4056 16661
rect 3728 16612 3770 16652
rect 3810 16612 3852 16652
rect 3892 16612 3934 16652
rect 3974 16612 4016 16652
rect 3688 16603 4056 16612
rect 4108 15560 4148 17788
rect 4204 17408 4244 17417
rect 4204 16484 4244 17368
rect 4204 16435 4244 16444
rect 3688 15140 4056 15149
rect 3728 15100 3770 15140
rect 3810 15100 3852 15140
rect 3892 15100 3934 15140
rect 3974 15100 4016 15140
rect 3688 15091 4056 15100
rect 3688 13628 4056 13637
rect 3728 13588 3770 13628
rect 3810 13588 3852 13628
rect 3892 13588 3934 13628
rect 3974 13588 4016 13628
rect 3688 13579 4056 13588
rect 3688 12116 4056 12125
rect 3728 12076 3770 12116
rect 3810 12076 3852 12116
rect 3892 12076 3934 12116
rect 3974 12076 4016 12116
rect 3688 12067 4056 12076
rect 4108 11612 4148 15520
rect 4108 11563 4148 11572
rect 4204 16232 4244 16241
rect 3688 10604 4056 10613
rect 3728 10564 3770 10604
rect 3810 10564 3852 10604
rect 3892 10564 3934 10604
rect 3974 10564 4016 10604
rect 3688 10555 4056 10564
rect 4107 10184 4149 10193
rect 4107 10144 4108 10184
rect 4148 10144 4149 10184
rect 4107 10135 4149 10144
rect 4108 10050 4148 10135
rect 3627 9428 3669 9437
rect 3627 9388 3628 9428
rect 3668 9388 3669 9428
rect 3627 9379 3669 9388
rect 4204 9428 4244 16192
rect 4300 15392 4340 15401
rect 4300 9437 4340 15352
rect 4204 9379 4244 9388
rect 4299 9428 4341 9437
rect 4299 9388 4300 9428
rect 4340 9388 4341 9428
rect 4299 9379 4341 9388
rect 3628 9294 3668 9379
rect 3688 9092 4056 9101
rect 3728 9052 3770 9092
rect 3810 9052 3852 9092
rect 3892 9052 3934 9092
rect 3974 9052 4016 9092
rect 3688 9043 4056 9052
rect 4204 8756 4244 8765
rect 3688 7580 4056 7589
rect 3728 7540 3770 7580
rect 3810 7540 3852 7580
rect 3892 7540 3934 7580
rect 3974 7540 4016 7580
rect 3688 7531 4056 7540
rect 3724 7076 3764 7085
rect 3724 6656 3764 7036
rect 3724 6607 3764 6616
rect 3688 6068 4056 6077
rect 3728 6028 3770 6068
rect 3810 6028 3852 6068
rect 3892 6028 3934 6068
rect 3974 6028 4016 6068
rect 3688 6019 4056 6028
rect 3688 4556 4056 4565
rect 3728 4516 3770 4556
rect 3810 4516 3852 4556
rect 3892 4516 3934 4556
rect 3974 4516 4016 4556
rect 3688 4507 4056 4516
rect 4204 3464 4244 8716
rect 4492 4304 4532 35680
rect 4928 35552 5296 35561
rect 4968 35512 5010 35552
rect 5050 35512 5092 35552
rect 5132 35512 5174 35552
rect 5214 35512 5256 35552
rect 4928 35503 5296 35512
rect 6604 34460 6644 35848
rect 4928 34040 5296 34049
rect 4968 34000 5010 34040
rect 5050 34000 5092 34040
rect 5132 34000 5174 34040
rect 5214 34000 5256 34040
rect 4928 33991 5296 34000
rect 5452 33704 5492 33713
rect 4684 33620 4724 33629
rect 4684 32192 4724 33580
rect 4928 32528 5296 32537
rect 4968 32488 5010 32528
rect 5050 32488 5092 32528
rect 5132 32488 5174 32528
rect 5214 32488 5256 32528
rect 4928 32479 5296 32488
rect 4684 23540 4724 32152
rect 4928 31016 5296 31025
rect 4968 30976 5010 31016
rect 5050 30976 5092 31016
rect 5132 30976 5174 31016
rect 5214 30976 5256 31016
rect 4928 30967 5296 30976
rect 4684 23491 4724 23500
rect 4780 30848 4820 30857
rect 4684 20852 4724 20861
rect 4684 19517 4724 20812
rect 4683 19508 4725 19517
rect 4683 19468 4684 19508
rect 4724 19468 4725 19508
rect 4683 19459 4725 19468
rect 4684 16484 4724 16493
rect 4684 14561 4724 16444
rect 4780 15317 4820 30808
rect 4928 29504 5296 29513
rect 4968 29464 5010 29504
rect 5050 29464 5092 29504
rect 5132 29464 5174 29504
rect 5214 29464 5256 29504
rect 4928 29455 5296 29464
rect 5452 29252 5492 33664
rect 6220 33284 6260 33293
rect 5452 29000 5492 29212
rect 5356 28960 5492 29000
rect 5836 33200 5876 33209
rect 4928 27992 5296 28001
rect 4968 27952 5010 27992
rect 5050 27952 5092 27992
rect 5132 27952 5174 27992
rect 5214 27952 5256 27992
rect 4928 27943 5296 27952
rect 5356 27488 5396 28960
rect 4928 26480 5296 26489
rect 4968 26440 5010 26480
rect 5050 26440 5092 26480
rect 5132 26440 5174 26480
rect 5214 26440 5256 26480
rect 4928 26431 5296 26440
rect 5356 26060 5396 27448
rect 4928 24968 5296 24977
rect 4968 24928 5010 24968
rect 5050 24928 5092 24968
rect 5132 24928 5174 24968
rect 5214 24928 5256 24968
rect 4928 24919 5296 24928
rect 4928 23456 5296 23465
rect 4968 23416 5010 23456
rect 5050 23416 5092 23456
rect 5132 23416 5174 23456
rect 5214 23416 5256 23456
rect 4928 23407 5296 23416
rect 4928 21944 5296 21953
rect 4968 21904 5010 21944
rect 5050 21904 5092 21944
rect 5132 21904 5174 21944
rect 5214 21904 5256 21944
rect 4928 21895 5296 21904
rect 4928 20432 5296 20441
rect 4968 20392 5010 20432
rect 5050 20392 5092 20432
rect 5132 20392 5174 20432
rect 5214 20392 5256 20432
rect 4928 20383 5296 20392
rect 5356 20096 5396 26020
rect 5644 24464 5684 24473
rect 5452 23792 5492 23801
rect 5452 23456 5492 23752
rect 5452 23407 5492 23416
rect 5548 23624 5588 23633
rect 5548 22784 5588 23584
rect 5548 22735 5588 22744
rect 4928 18920 5296 18929
rect 4968 18880 5010 18920
rect 5050 18880 5092 18920
rect 5132 18880 5174 18920
rect 5214 18880 5256 18920
rect 4928 18871 5296 18880
rect 4928 17408 5296 17417
rect 4968 17368 5010 17408
rect 5050 17368 5092 17408
rect 5132 17368 5174 17408
rect 5214 17368 5256 17408
rect 4928 17359 5296 17368
rect 5067 16148 5109 16157
rect 5067 16108 5068 16148
rect 5108 16108 5109 16148
rect 5067 16099 5109 16108
rect 5068 16014 5108 16099
rect 4928 15896 5296 15905
rect 4968 15856 5010 15896
rect 5050 15856 5092 15896
rect 5132 15856 5174 15896
rect 5214 15856 5256 15896
rect 4928 15847 5296 15856
rect 4779 15308 4821 15317
rect 4779 15268 4780 15308
rect 4820 15268 4821 15308
rect 4779 15259 4821 15268
rect 4683 14552 4725 14561
rect 4683 14512 4684 14552
rect 4724 14512 4725 14552
rect 4683 14503 4725 14512
rect 4588 11360 4628 11369
rect 4588 10193 4628 11320
rect 4587 10184 4629 10193
rect 4587 10144 4588 10184
rect 4628 10144 4629 10184
rect 4587 10135 4629 10144
rect 4492 4255 4532 4264
rect 4588 9176 4628 9185
rect 4204 3415 4244 3424
rect 3916 3380 3956 3391
rect 3916 3305 3956 3340
rect 4588 3305 4628 9136
rect 4684 5732 4724 14503
rect 4780 10772 4820 15259
rect 4928 14384 5296 14393
rect 4968 14344 5010 14384
rect 5050 14344 5092 14384
rect 5132 14344 5174 14384
rect 5214 14344 5256 14384
rect 4928 14335 5296 14344
rect 4928 12872 5296 12881
rect 4968 12832 5010 12872
rect 5050 12832 5092 12872
rect 5132 12832 5174 12872
rect 5214 12832 5256 12872
rect 4928 12823 5296 12832
rect 4928 11360 5296 11369
rect 4968 11320 5010 11360
rect 5050 11320 5092 11360
rect 5132 11320 5174 11360
rect 5214 11320 5256 11360
rect 5356 11360 5396 20056
rect 5644 11528 5684 24424
rect 5740 23792 5780 23801
rect 5740 16148 5780 23752
rect 5740 16099 5780 16108
rect 5740 15980 5780 15989
rect 5740 11948 5780 15940
rect 5740 11899 5780 11908
rect 5739 11780 5781 11789
rect 5739 11740 5740 11780
rect 5780 11740 5781 11780
rect 5739 11731 5781 11740
rect 5644 11479 5684 11488
rect 5356 11320 5588 11360
rect 4928 11311 5296 11320
rect 4780 10723 4820 10732
rect 4928 9848 5296 9857
rect 4968 9808 5010 9848
rect 5050 9808 5092 9848
rect 5132 9808 5174 9848
rect 5214 9808 5256 9848
rect 4928 9799 5296 9808
rect 4928 8336 5296 8345
rect 4968 8296 5010 8336
rect 5050 8296 5092 8336
rect 5132 8296 5174 8336
rect 5214 8296 5256 8336
rect 4928 8287 5296 8296
rect 4780 7580 4820 7589
rect 4780 5816 4820 7540
rect 4928 6824 5296 6833
rect 4968 6784 5010 6824
rect 5050 6784 5092 6824
rect 5132 6784 5174 6824
rect 5214 6784 5256 6824
rect 4928 6775 5296 6784
rect 5451 6152 5493 6161
rect 5451 6112 5452 6152
rect 5492 6112 5493 6152
rect 5451 6103 5493 6112
rect 5355 5984 5397 5993
rect 5355 5944 5356 5984
rect 5396 5944 5397 5984
rect 5355 5935 5397 5944
rect 4780 5767 4820 5776
rect 4684 5060 4724 5692
rect 4928 5312 5296 5321
rect 4968 5272 5010 5312
rect 5050 5272 5092 5312
rect 5132 5272 5174 5312
rect 5214 5272 5256 5312
rect 4928 5263 5296 5272
rect 4684 5011 4724 5020
rect 4928 3800 5296 3809
rect 4968 3760 5010 3800
rect 5050 3760 5092 3800
rect 5132 3760 5174 3800
rect 5214 3760 5256 3800
rect 4928 3751 5296 3760
rect 3915 3296 3957 3305
rect 3915 3256 3916 3296
rect 3956 3256 3957 3296
rect 3915 3247 3957 3256
rect 4587 3296 4629 3305
rect 4587 3256 4588 3296
rect 4628 3256 4629 3296
rect 4587 3247 4629 3256
rect 3688 3044 4056 3053
rect 3728 3004 3770 3044
rect 3810 3004 3852 3044
rect 3892 3004 3934 3044
rect 3974 3004 4016 3044
rect 3688 2995 4056 3004
rect 4928 2288 5296 2297
rect 4968 2248 5010 2288
rect 5050 2248 5092 2288
rect 5132 2248 5174 2288
rect 5214 2248 5256 2288
rect 4928 2239 5296 2248
rect 3688 1532 4056 1541
rect 3728 1492 3770 1532
rect 3810 1492 3852 1532
rect 3892 1492 3934 1532
rect 3974 1492 4016 1532
rect 3688 1483 4056 1492
rect 4107 1364 4149 1373
rect 4107 1324 4108 1364
rect 4148 1324 4149 1364
rect 4107 1315 4149 1324
rect 3532 1231 3572 1240
rect 2764 895 2804 904
rect 4108 944 4148 1315
rect 4683 1280 4725 1289
rect 4683 1240 4684 1280
rect 4724 1240 4725 1280
rect 4683 1231 4725 1240
rect 4108 895 4148 904
rect 2572 727 2612 736
rect 4684 608 4724 1231
rect 4780 1112 4820 1121
rect 4780 944 4820 1072
rect 4780 895 4820 904
rect 4928 776 5296 785
rect 4968 736 5010 776
rect 5050 736 5092 776
rect 5132 736 5174 776
rect 5214 736 5256 776
rect 4928 727 5296 736
rect 4684 559 4724 568
rect 5356 608 5396 5935
rect 5452 1280 5492 6103
rect 5548 4724 5588 11320
rect 5643 6488 5685 6497
rect 5643 6448 5644 6488
rect 5684 6448 5685 6488
rect 5643 6439 5685 6448
rect 5644 6354 5684 6439
rect 5548 2297 5588 4684
rect 5740 4136 5780 11731
rect 5740 4087 5780 4096
rect 5836 2540 5876 33160
rect 6220 32696 6260 33244
rect 6220 32647 6260 32656
rect 6220 27824 6260 27833
rect 6220 26564 6260 27784
rect 6220 26515 6260 26524
rect 6220 25304 6260 25313
rect 6028 25220 6068 25229
rect 5932 20768 5972 20777
rect 5932 14048 5972 20728
rect 6028 18332 6068 25180
rect 6028 18283 6068 18292
rect 6220 18920 6260 25264
rect 6508 25304 6548 25313
rect 6412 24968 6452 24977
rect 6316 23036 6356 23045
rect 6316 20936 6356 22996
rect 6316 20887 6356 20896
rect 6412 20768 6452 24928
rect 6508 22196 6548 25264
rect 6508 22147 6548 22156
rect 6412 20719 6452 20728
rect 5932 11360 5972 14008
rect 6220 11789 6260 18880
rect 6508 14300 6548 14309
rect 6508 13628 6548 14260
rect 6508 13579 6548 13588
rect 6219 11780 6261 11789
rect 6219 11740 6220 11780
rect 6260 11740 6261 11780
rect 6219 11731 6261 11740
rect 5932 11320 6068 11360
rect 5931 4220 5973 4229
rect 5931 4180 5932 4220
rect 5972 4180 5973 4220
rect 5931 4171 5973 4180
rect 5932 4086 5972 4171
rect 6028 3221 6068 11320
rect 6508 8168 6548 8177
rect 6027 3212 6069 3221
rect 6027 3172 6028 3212
rect 6068 3172 6069 3212
rect 6027 3163 6069 3172
rect 5836 2500 5972 2540
rect 5547 2288 5589 2297
rect 5547 2248 5548 2288
rect 5588 2248 5589 2288
rect 5547 2239 5589 2248
rect 5548 1952 5588 2239
rect 5548 1903 5588 1912
rect 5452 1231 5492 1240
rect 5932 692 5972 2500
rect 5932 643 5972 652
rect 6508 692 6548 8128
rect 6604 1280 6644 34420
rect 6700 28748 6740 36520
rect 6700 28699 6740 28708
rect 6700 26144 6740 26153
rect 6700 21524 6740 26104
rect 6700 21475 6740 21484
rect 6796 23372 6836 23381
rect 6700 20768 6740 20777
rect 6700 9932 6740 20728
rect 6700 9883 6740 9892
rect 6796 4976 6836 23332
rect 6796 4927 6836 4936
rect 6892 3884 6932 37192
rect 7180 33284 7220 33293
rect 7084 32780 7124 32789
rect 7084 31604 7124 32740
rect 6796 3844 6932 3884
rect 6988 31352 7028 31361
rect 6700 2708 6740 2717
rect 6700 2381 6740 2668
rect 6796 2540 6836 3844
rect 6891 3716 6933 3725
rect 6891 3676 6892 3716
rect 6932 3676 6933 3716
rect 6891 3667 6933 3676
rect 6892 3582 6932 3667
rect 6796 2500 6932 2540
rect 6699 2372 6741 2381
rect 6699 2332 6700 2372
rect 6740 2332 6741 2372
rect 6699 2323 6741 2332
rect 6604 1231 6644 1240
rect 6508 643 6548 652
rect 5356 559 5396 568
rect 2476 475 2516 484
rect 6411 440 6453 449
rect 6411 400 6412 440
rect 6452 400 6453 440
rect 6411 391 6453 400
rect 2380 307 2420 316
rect 6412 306 6452 391
rect 6892 356 6932 2500
rect 6988 776 7028 31312
rect 7084 29924 7124 31564
rect 7084 29875 7124 29884
rect 7180 29756 7220 33244
rect 7180 29707 7220 29716
rect 7276 30680 7316 30689
rect 7180 27740 7220 27749
rect 7083 23036 7125 23045
rect 7083 22996 7084 23036
rect 7124 22996 7125 23036
rect 7083 22987 7125 22996
rect 7084 22902 7124 22987
rect 7180 22868 7220 27700
rect 7180 19844 7220 22828
rect 7180 19592 7220 19804
rect 7180 19543 7220 19552
rect 7276 14216 7316 30640
rect 7276 14167 7316 14176
rect 7084 14132 7124 14141
rect 7084 5396 7124 14092
rect 7084 3464 7124 5356
rect 7084 3415 7124 3424
rect 7180 4976 7220 4985
rect 7180 1196 7220 4936
rect 7276 3716 7316 3725
rect 7276 3548 7316 3676
rect 7276 3499 7316 3508
rect 7180 1147 7220 1156
rect 6988 727 7028 736
rect 7372 524 7412 38116
rect 7564 37400 7604 37409
rect 7468 35468 7508 35477
rect 7468 30848 7508 35428
rect 7468 28496 7508 30808
rect 7468 28447 7508 28456
rect 7564 13040 7604 37360
rect 7756 31688 7796 31697
rect 7756 28412 7796 31648
rect 7756 28363 7796 28372
rect 7948 25304 7988 25313
rect 7852 24800 7892 24809
rect 7564 12991 7604 13000
rect 7660 22196 7700 22205
rect 7660 22028 7700 22156
rect 7468 11864 7508 11873
rect 7468 7832 7508 11824
rect 7660 9596 7700 21988
rect 7660 9547 7700 9556
rect 7756 21104 7796 21113
rect 7563 9428 7605 9437
rect 7563 9388 7564 9428
rect 7604 9388 7605 9428
rect 7563 9379 7605 9388
rect 7564 9092 7604 9379
rect 7564 9043 7604 9052
rect 7468 7783 7508 7792
rect 7468 4472 7508 4481
rect 7468 2708 7508 4432
rect 7660 3800 7700 3809
rect 7468 2659 7508 2668
rect 7564 3548 7604 3557
rect 7564 2120 7604 3508
rect 7660 2372 7700 3760
rect 7660 2323 7700 2332
rect 7564 2071 7604 2080
rect 7467 1868 7509 1877
rect 7467 1828 7468 1868
rect 7508 1828 7509 1868
rect 7467 1819 7509 1828
rect 7468 1784 7508 1819
rect 7468 1733 7508 1744
rect 7756 1280 7796 21064
rect 7852 20768 7892 24760
rect 7852 19088 7892 20728
rect 7852 19039 7892 19048
rect 7948 21608 7988 25264
rect 7948 17660 7988 21568
rect 7948 17611 7988 17620
rect 7948 15728 7988 15737
rect 7948 12116 7988 15688
rect 8044 15140 8084 41140
rect 9772 40340 9812 40349
rect 8908 39248 8948 39257
rect 8620 38576 8660 38585
rect 8428 38156 8468 38165
rect 8332 37736 8372 37745
rect 8332 37316 8372 37696
rect 8332 37267 8372 37276
rect 8140 34376 8180 34385
rect 8140 17828 8180 34336
rect 8236 33704 8276 33713
rect 8236 23792 8276 33664
rect 8236 17912 8276 23752
rect 8332 23624 8372 23633
rect 8332 22784 8372 23584
rect 8332 22735 8372 22744
rect 8236 17863 8276 17872
rect 8140 17779 8180 17788
rect 8044 15091 8084 15100
rect 7948 12067 7988 12076
rect 8044 12452 8084 12461
rect 7851 2372 7893 2381
rect 7851 2332 7852 2372
rect 7892 2332 7893 2372
rect 7851 2323 7893 2332
rect 7852 2238 7892 2323
rect 7756 1231 7796 1240
rect 8044 1196 8084 12412
rect 8332 11444 8372 11453
rect 8332 11108 8372 11404
rect 8332 11059 8372 11068
rect 8428 1289 8468 38116
rect 8620 32612 8660 38536
rect 8812 35972 8852 35981
rect 8716 35300 8756 35309
rect 8716 35048 8756 35260
rect 8716 34999 8756 35008
rect 8620 32192 8660 32572
rect 8620 32143 8660 32152
rect 8620 23708 8660 23717
rect 8524 21524 8564 21533
rect 8524 13964 8564 21484
rect 8620 20096 8660 23668
rect 8620 20047 8660 20056
rect 8716 23120 8756 23129
rect 8524 11360 8564 13924
rect 8620 13628 8660 13637
rect 8620 12200 8660 13588
rect 8620 12151 8660 12160
rect 8524 11320 8660 11360
rect 8524 3632 8564 3641
rect 8524 2204 8564 3592
rect 8620 2372 8660 11320
rect 8716 3809 8756 23080
rect 8812 19088 8852 35932
rect 8812 19039 8852 19048
rect 8812 14216 8852 14225
rect 8812 11192 8852 14176
rect 8812 11143 8852 11152
rect 8811 9344 8853 9353
rect 8811 9304 8812 9344
rect 8852 9304 8853 9344
rect 8811 9295 8853 9304
rect 8812 8840 8852 9295
rect 8812 8791 8852 8800
rect 8908 6161 8948 39208
rect 9579 38240 9621 38249
rect 9579 38200 9580 38240
rect 9620 38200 9621 38240
rect 9579 38191 9621 38200
rect 9580 38106 9620 38191
rect 9196 37148 9236 37157
rect 9388 37148 9428 37157
rect 9236 37108 9388 37148
rect 9196 37099 9236 37108
rect 9388 37099 9428 37108
rect 9676 35888 9716 35897
rect 9004 35720 9044 35729
rect 8907 6152 8949 6161
rect 8907 6112 8908 6152
rect 8948 6112 8949 6152
rect 8907 6103 8949 6112
rect 8715 3800 8757 3809
rect 8715 3760 8716 3800
rect 8756 3760 8757 3800
rect 8715 3751 8757 3760
rect 9004 3548 9044 35680
rect 9580 35468 9620 35477
rect 9292 35300 9332 35309
rect 9292 33452 9332 35260
rect 9292 33403 9332 33412
rect 9388 34712 9428 34721
rect 9292 33284 9332 33293
rect 9196 18164 9236 18173
rect 9196 13712 9236 18124
rect 9196 13663 9236 13672
rect 9196 11360 9236 11369
rect 9100 10436 9140 10445
rect 9100 9848 9140 10396
rect 9100 9799 9140 9808
rect 9196 9680 9236 11320
rect 9196 9631 9236 9640
rect 9004 3499 9044 3508
rect 8620 2323 8660 2332
rect 8524 1784 8564 2164
rect 8619 1868 8661 1877
rect 8619 1828 8620 1868
rect 8660 1828 8661 1868
rect 8619 1819 8661 1828
rect 8524 1735 8564 1744
rect 8620 1734 8660 1819
rect 8427 1280 8469 1289
rect 8427 1240 8428 1280
rect 8468 1240 8469 1280
rect 8427 1231 8469 1240
rect 9292 1280 9332 33244
rect 9388 15308 9428 34672
rect 9580 32957 9620 35428
rect 9579 32948 9621 32957
rect 9579 32908 9580 32948
rect 9620 32908 9621 32948
rect 9579 32899 9621 32908
rect 9388 15259 9428 15268
rect 9484 16316 9524 16325
rect 9484 13208 9524 16276
rect 9484 13159 9524 13168
rect 9388 11024 9428 11033
rect 9388 10268 9428 10984
rect 9388 10219 9428 10228
rect 9484 10520 9524 10529
rect 9484 9680 9524 10480
rect 9484 9631 9524 9640
rect 9580 9260 9620 9269
rect 9580 4229 9620 9220
rect 9579 4220 9621 4229
rect 9579 4180 9580 4220
rect 9620 4180 9621 4220
rect 9579 4171 9621 4180
rect 9292 1231 9332 1240
rect 8044 1147 8084 1156
rect 9580 1196 9620 4171
rect 9676 1373 9716 35848
rect 9772 5993 9812 40300
rect 9868 6497 9908 41560
rect 10060 41600 10100 41609
rect 10060 10352 10100 41560
rect 11404 41600 11444 41609
rect 10924 40676 10964 40685
rect 10828 40424 10868 40433
rect 10252 40256 10292 40265
rect 10252 38081 10292 40216
rect 10348 38240 10388 38249
rect 10251 38072 10293 38081
rect 10251 38032 10252 38072
rect 10292 38032 10293 38072
rect 10251 38023 10293 38032
rect 10156 32864 10196 32873
rect 10156 27404 10196 32824
rect 10156 26816 10196 27364
rect 10156 26767 10196 26776
rect 10156 24632 10196 24641
rect 10156 10529 10196 24592
rect 10252 20600 10292 20609
rect 10252 17744 10292 20560
rect 10155 10520 10197 10529
rect 10155 10480 10156 10520
rect 10196 10480 10197 10520
rect 10155 10471 10197 10480
rect 10060 10312 10196 10352
rect 10060 10184 10100 10193
rect 10060 8672 10100 10144
rect 10156 9260 10196 10312
rect 10156 9211 10196 9220
rect 10060 8623 10100 8632
rect 10252 6908 10292 17704
rect 10252 6859 10292 6868
rect 9867 6488 9909 6497
rect 9867 6448 9868 6488
rect 9908 6448 9909 6488
rect 9867 6439 9909 6448
rect 9771 5984 9813 5993
rect 9771 5944 9772 5984
rect 9812 5944 9813 5984
rect 9771 5935 9813 5944
rect 9868 2540 9908 6439
rect 9868 2500 10100 2540
rect 9675 1364 9717 1373
rect 9675 1324 9676 1364
rect 9716 1324 9717 1364
rect 9675 1315 9717 1324
rect 9580 1147 9620 1156
rect 10060 1196 10100 2500
rect 10348 1868 10388 38200
rect 10444 34040 10484 34049
rect 10444 33704 10484 34000
rect 10444 33655 10484 33664
rect 10636 31604 10676 31613
rect 10636 24296 10676 31564
rect 10540 13544 10580 13553
rect 10443 10520 10485 10529
rect 10443 10480 10444 10520
rect 10484 10480 10485 10520
rect 10443 10471 10485 10480
rect 10444 7748 10484 10471
rect 10540 9428 10580 13504
rect 10636 10520 10676 24256
rect 10636 10471 10676 10480
rect 10540 9260 10580 9388
rect 10540 9211 10580 9220
rect 10444 7699 10484 7708
rect 10348 1819 10388 1828
rect 10828 1868 10868 40384
rect 10924 39668 10964 40636
rect 10924 39619 10964 39628
rect 11116 39668 11156 39677
rect 11020 27740 11060 27749
rect 11020 24632 11060 27700
rect 10924 24592 11020 24632
rect 10924 22364 10964 24592
rect 11020 24583 11060 24592
rect 10924 22315 10964 22324
rect 11020 23708 11060 23717
rect 11020 22280 11060 23668
rect 11020 22231 11060 22240
rect 10924 16652 10964 16661
rect 10924 9353 10964 16612
rect 11019 15476 11061 15485
rect 11019 15436 11020 15476
rect 11060 15436 11061 15476
rect 11019 15427 11061 15436
rect 11020 15140 11060 15427
rect 11020 15091 11060 15100
rect 10923 9344 10965 9353
rect 10923 9304 10924 9344
rect 10964 9304 10965 9344
rect 10923 9295 10965 9304
rect 10924 9210 10964 9295
rect 10828 1819 10868 1828
rect 11116 1868 11156 39628
rect 11116 1819 11156 1828
rect 11212 38828 11252 38837
rect 11212 37904 11252 38788
rect 10060 1147 10100 1156
rect 10828 1028 10868 1037
rect 7947 944 7989 953
rect 7947 904 7948 944
rect 7988 904 7989 944
rect 7947 895 7989 904
rect 7948 810 7988 895
rect 7372 475 7412 484
rect 7948 608 7988 617
rect 6892 307 6932 316
rect 2188 223 2228 232
rect 7948 104 7988 568
rect 8139 608 8181 617
rect 8139 568 8140 608
rect 8180 568 8181 608
rect 8139 559 8181 568
rect 8140 474 8180 559
rect 7948 55 7988 64
rect 10828 104 10868 988
rect 11212 1028 11252 37864
rect 11308 23960 11348 23969
rect 11308 23708 11348 23920
rect 11308 23659 11348 23668
rect 11308 15812 11348 15821
rect 11308 14972 11348 15772
rect 11308 14923 11348 14932
rect 11308 13376 11348 13385
rect 11308 10688 11348 13336
rect 11308 10639 11348 10648
rect 11404 6824 11444 41560
rect 11596 41600 11636 41609
rect 11404 6775 11444 6784
rect 11500 28748 11540 28757
rect 11212 979 11252 988
rect 11500 953 11540 28708
rect 11596 4472 11636 41560
rect 11788 39164 11828 42568
rect 14668 42608 14708 42617
rect 13324 41012 13364 41021
rect 11788 39115 11828 39124
rect 12364 39584 12404 39593
rect 11980 36644 12020 36653
rect 11884 26060 11924 26069
rect 11884 19928 11924 26020
rect 11788 16904 11828 16913
rect 11691 15476 11733 15485
rect 11691 15436 11692 15476
rect 11732 15436 11733 15476
rect 11691 15427 11733 15436
rect 11692 14132 11732 15427
rect 11692 14083 11732 14092
rect 11788 9344 11828 16864
rect 11788 9295 11828 9304
rect 11884 9092 11924 19888
rect 11980 18752 12020 36604
rect 11980 18703 12020 18712
rect 12268 32108 12308 32117
rect 12268 17744 12308 32068
rect 12172 13880 12212 13889
rect 12172 12872 12212 13840
rect 12172 12823 12212 12832
rect 12172 12620 12212 12629
rect 12076 11612 12116 11621
rect 12076 11192 12116 11572
rect 12076 11143 12116 11152
rect 11884 9043 11924 9052
rect 11596 4423 11636 4432
rect 11499 944 11541 953
rect 11499 904 11500 944
rect 11540 904 11541 944
rect 11499 895 11541 904
rect 12172 272 12212 12580
rect 12268 8672 12308 17704
rect 12268 6068 12308 8632
rect 12268 6019 12308 6028
rect 12364 1457 12404 39544
rect 12940 39332 12980 39341
rect 12652 38408 12692 38417
rect 12652 38240 12692 38368
rect 12843 38408 12885 38417
rect 12843 38368 12844 38408
rect 12884 38368 12885 38408
rect 12843 38359 12885 38368
rect 12844 38274 12884 38359
rect 12652 38191 12692 38200
rect 12652 36728 12692 36737
rect 12652 35216 12692 36688
rect 12652 33368 12692 35176
rect 12652 33319 12692 33328
rect 12844 35132 12884 35141
rect 12652 32864 12692 32873
rect 12460 20852 12500 20861
rect 12460 10856 12500 20812
rect 12556 20768 12596 20777
rect 12556 15485 12596 20728
rect 12555 15476 12597 15485
rect 12555 15436 12556 15476
rect 12596 15436 12597 15476
rect 12555 15427 12597 15436
rect 12460 10807 12500 10816
rect 12556 15140 12596 15149
rect 12556 5144 12596 15100
rect 12652 5228 12692 32824
rect 12844 29336 12884 35092
rect 12748 20768 12788 20777
rect 12748 9848 12788 20728
rect 12844 19256 12884 29296
rect 12844 19207 12884 19216
rect 12844 11612 12884 11621
rect 12844 10856 12884 11572
rect 12844 10807 12884 10816
rect 12748 9799 12788 9808
rect 12652 5179 12692 5188
rect 12556 5095 12596 5104
rect 12363 1448 12405 1457
rect 12363 1408 12364 1448
rect 12404 1408 12405 1448
rect 12363 1399 12405 1408
rect 12940 617 12980 39292
rect 13036 34880 13076 34889
rect 13036 22280 13076 34840
rect 13036 22231 13076 22240
rect 13228 16400 13268 16409
rect 13132 12620 13172 12629
rect 13132 11612 13172 12580
rect 13132 11563 13172 11572
rect 13228 9428 13268 16360
rect 13228 9379 13268 9388
rect 13228 6908 13268 6917
rect 13228 1700 13268 6868
rect 13324 3632 13364 40972
rect 14092 40592 14132 40601
rect 13516 39164 13556 39173
rect 13420 19676 13460 19685
rect 13420 19424 13460 19636
rect 13420 11360 13460 19384
rect 13516 12629 13556 39124
rect 13707 38660 13749 38669
rect 13707 38620 13708 38660
rect 13748 38620 13749 38660
rect 13707 38611 13749 38620
rect 13612 32108 13652 32117
rect 13515 12620 13557 12629
rect 13515 12580 13516 12620
rect 13556 12580 13557 12620
rect 13515 12571 13557 12580
rect 13420 11320 13556 11360
rect 13419 6992 13461 7001
rect 13419 6952 13420 6992
rect 13460 6952 13461 6992
rect 13419 6943 13461 6952
rect 13420 6858 13460 6943
rect 13516 4976 13556 11320
rect 13516 4927 13556 4936
rect 13324 3583 13364 3592
rect 13228 1651 13268 1660
rect 13515 1028 13557 1037
rect 13515 988 13516 1028
rect 13556 988 13557 1028
rect 13515 979 13557 988
rect 13516 894 13556 979
rect 12939 608 12981 617
rect 12939 568 12940 608
rect 12980 568 12981 608
rect 12939 559 12981 568
rect 12172 223 12212 232
rect 13612 188 13652 32068
rect 13708 1448 13748 38611
rect 13804 34712 13844 34721
rect 13804 34292 13844 34672
rect 13804 34243 13844 34252
rect 13900 27068 13940 27077
rect 13804 26144 13844 26153
rect 13804 24548 13844 26104
rect 13804 24499 13844 24508
rect 13900 23792 13940 27028
rect 13804 22364 13844 22373
rect 13804 17996 13844 22324
rect 13900 19424 13940 23752
rect 13900 19375 13940 19384
rect 13996 21608 14036 21617
rect 13996 19844 14036 21568
rect 13804 17947 13844 17956
rect 13900 15140 13940 15149
rect 13900 14300 13940 15100
rect 13900 14251 13940 14260
rect 13804 4976 13844 4985
rect 13804 3725 13844 4936
rect 13996 4817 14036 19804
rect 13995 4808 14037 4817
rect 13995 4768 13996 4808
rect 14036 4768 14037 4808
rect 13995 4759 14037 4768
rect 13803 3716 13845 3725
rect 13803 3676 13804 3716
rect 13844 3676 13845 3716
rect 13803 3667 13845 3676
rect 13899 2288 13941 2297
rect 13899 2248 13900 2288
rect 13940 2248 13941 2288
rect 13899 2239 13941 2248
rect 13900 2154 13940 2239
rect 13708 1399 13748 1408
rect 14092 1280 14132 40552
rect 14476 40592 14516 40601
rect 14188 38912 14228 38921
rect 14188 38240 14228 38872
rect 14188 38191 14228 38200
rect 14284 25220 14324 25229
rect 14284 20684 14324 25180
rect 14380 22280 14420 22289
rect 14380 20768 14420 22240
rect 14380 20719 14420 20728
rect 14284 20635 14324 20644
rect 14284 19424 14324 19433
rect 14284 9008 14324 19384
rect 14284 8959 14324 8968
rect 14187 3800 14229 3809
rect 14187 3760 14188 3800
rect 14228 3760 14229 3800
rect 14187 3751 14229 3760
rect 14188 2708 14228 3751
rect 14188 2659 14228 2668
rect 14092 1231 14132 1240
rect 14476 1112 14516 40552
rect 14668 36896 14708 42568
rect 18700 42188 18740 42197
rect 17932 41600 17972 41609
rect 16684 41264 16724 41273
rect 15628 41012 15668 41021
rect 15532 40972 15628 41012
rect 14668 36847 14708 36856
rect 14860 40592 14900 40601
rect 14764 35468 14804 35477
rect 14668 34880 14708 34889
rect 14572 33116 14612 33125
rect 14572 30512 14612 33076
rect 14572 27656 14612 30472
rect 14572 27607 14612 27616
rect 14668 26480 14708 34840
rect 14764 30260 14804 35428
rect 14764 30211 14804 30220
rect 14668 26431 14708 26440
rect 14572 26312 14612 26321
rect 14572 17156 14612 26272
rect 14764 26312 14804 26321
rect 14764 18416 14804 26272
rect 14764 17828 14804 18376
rect 14764 17779 14804 17788
rect 14572 17107 14612 17116
rect 14668 17492 14708 17501
rect 14668 14216 14708 17452
rect 14763 16652 14805 16661
rect 14763 16612 14764 16652
rect 14804 16612 14805 16652
rect 14763 16603 14805 16612
rect 14668 14167 14708 14176
rect 14764 13880 14804 16603
rect 14764 13831 14804 13840
rect 14668 12620 14708 12629
rect 14668 9428 14708 12580
rect 14668 9379 14708 9388
rect 14476 1063 14516 1072
rect 14283 860 14325 869
rect 14283 820 14284 860
rect 14324 820 14325 860
rect 14283 811 14325 820
rect 13707 776 13749 785
rect 13707 736 13708 776
rect 13748 736 13749 776
rect 13707 727 13749 736
rect 13708 642 13748 727
rect 14284 726 14324 811
rect 14860 524 14900 40552
rect 15148 40592 15188 40601
rect 14956 40340 14996 40349
rect 14956 16661 14996 40300
rect 15051 38744 15093 38753
rect 15051 38704 15052 38744
rect 15092 38704 15093 38744
rect 15051 38695 15093 38704
rect 14955 16652 14997 16661
rect 14955 16612 14956 16652
rect 14996 16612 14997 16652
rect 14955 16603 14997 16612
rect 14955 14552 14997 14561
rect 14955 14512 14956 14552
rect 14996 14512 14997 14552
rect 14955 14503 14997 14512
rect 14956 14300 14996 14503
rect 14956 14251 14996 14260
rect 15052 1616 15092 38695
rect 15052 1567 15092 1576
rect 15148 1037 15188 40552
rect 15244 40340 15284 40349
rect 15147 1028 15189 1037
rect 15147 988 15148 1028
rect 15188 988 15189 1028
rect 15147 979 15189 988
rect 14860 475 14900 484
rect 15244 440 15284 40300
rect 15436 34040 15476 34049
rect 15436 29756 15476 34000
rect 15436 28496 15476 29716
rect 15436 28447 15476 28456
rect 15532 2540 15572 40972
rect 15628 40963 15668 40972
rect 16012 41012 16052 41021
rect 15820 40592 15860 40601
rect 15628 40340 15668 40349
rect 15628 13880 15668 40300
rect 15724 37736 15764 37745
rect 15724 30680 15764 37696
rect 15724 30631 15764 30640
rect 15628 13831 15668 13840
rect 15724 19004 15764 19013
rect 15724 13796 15764 18964
rect 15724 12200 15764 13756
rect 15724 12151 15764 12160
rect 15627 5816 15669 5825
rect 15627 5776 15628 5816
rect 15668 5776 15669 5816
rect 15627 5767 15669 5776
rect 15628 5682 15668 5767
rect 15820 2540 15860 40552
rect 15436 2500 15572 2540
rect 15724 2500 15860 2540
rect 15916 35132 15956 35141
rect 15436 608 15476 2500
rect 15436 559 15476 568
rect 15244 391 15284 400
rect 14091 356 14133 365
rect 14091 316 14092 356
rect 14132 316 14133 356
rect 14091 307 14133 316
rect 14092 222 14132 307
rect 15724 272 15764 2500
rect 15916 944 15956 35092
rect 15916 895 15956 904
rect 16012 785 16052 40972
rect 16396 40592 16436 40601
rect 16300 37148 16340 37157
rect 16300 35972 16340 37108
rect 16300 35923 16340 35932
rect 16108 35384 16148 35393
rect 16108 34880 16148 35344
rect 16108 34831 16148 34840
rect 16108 18248 16148 18257
rect 16108 12200 16148 18208
rect 16108 12151 16148 12160
rect 16300 15140 16340 15149
rect 16204 7832 16244 7841
rect 16204 2372 16244 7792
rect 16300 2792 16340 15100
rect 16396 11360 16436 40552
rect 16684 38912 16724 41224
rect 17644 40844 17684 40853
rect 17356 40340 17396 40349
rect 17163 39836 17205 39845
rect 17163 39796 17164 39836
rect 17204 39796 17205 39836
rect 17163 39787 17205 39796
rect 17164 39702 17204 39787
rect 17260 39584 17300 39593
rect 16684 38863 16724 38872
rect 16876 39500 16916 39509
rect 16492 35552 16532 35561
rect 16492 31436 16532 35512
rect 16492 29000 16532 31396
rect 16780 34376 16820 34385
rect 16684 30848 16724 30857
rect 16492 28960 16628 29000
rect 16492 25724 16532 25733
rect 16492 24968 16532 25684
rect 16492 24919 16532 24928
rect 16588 25304 16628 28960
rect 16684 27908 16724 30808
rect 16780 30680 16820 34336
rect 16780 30631 16820 30640
rect 16684 27859 16724 27868
rect 16588 24884 16628 25264
rect 16588 20012 16628 24844
rect 16588 19963 16628 19972
rect 16491 19088 16533 19097
rect 16491 19048 16492 19088
rect 16532 19048 16533 19088
rect 16491 19039 16533 19048
rect 16492 14804 16532 19039
rect 16780 17744 16820 17753
rect 16492 14755 16532 14764
rect 16588 16652 16628 16661
rect 16492 13124 16532 13133
rect 16492 12536 16532 13084
rect 16492 12487 16532 12496
rect 16588 11528 16628 16612
rect 16684 14636 16724 14645
rect 16684 13964 16724 14596
rect 16684 13915 16724 13924
rect 16588 11479 16628 11488
rect 16396 11320 16532 11360
rect 16395 10184 16437 10193
rect 16395 10144 16396 10184
rect 16436 10144 16437 10184
rect 16395 10135 16437 10144
rect 16396 7160 16436 10135
rect 16396 7111 16436 7120
rect 16300 2624 16340 2752
rect 16300 2575 16340 2584
rect 16204 2323 16244 2332
rect 16011 776 16053 785
rect 16011 736 16012 776
rect 16052 736 16053 776
rect 16011 727 16053 736
rect 16492 365 16532 11320
rect 16780 7748 16820 17704
rect 16588 5060 16628 5069
rect 16588 4136 16628 5020
rect 16588 4087 16628 4096
rect 16684 4304 16724 4313
rect 16588 3800 16628 3809
rect 16588 2540 16628 3760
rect 16588 2491 16628 2500
rect 16684 2456 16724 4264
rect 16684 2407 16724 2416
rect 16780 1280 16820 7708
rect 16780 1231 16820 1240
rect 16876 860 16916 39460
rect 17068 35048 17108 35057
rect 16972 33116 17012 33125
rect 16972 32360 17012 33076
rect 16972 32311 17012 32320
rect 17068 30848 17108 35008
rect 17068 30799 17108 30808
rect 17068 24464 17108 24473
rect 16971 19508 17013 19517
rect 16971 19468 16972 19508
rect 17012 19468 17013 19508
rect 16971 19459 17013 19468
rect 16972 8504 17012 19459
rect 17068 18752 17108 24424
rect 17068 18703 17108 18712
rect 17164 20684 17204 20693
rect 17164 18668 17204 20644
rect 17067 16400 17109 16409
rect 17067 16360 17068 16400
rect 17108 16360 17109 16400
rect 17067 16351 17109 16360
rect 17068 16266 17108 16351
rect 17164 10184 17204 18628
rect 17164 10135 17204 10144
rect 16972 8455 17012 8464
rect 16972 7748 17012 7757
rect 16972 4136 17012 7708
rect 16972 4087 17012 4096
rect 17068 7664 17108 7673
rect 16876 811 16916 820
rect 17068 608 17108 7624
rect 17164 6992 17204 7001
rect 17164 4136 17204 6952
rect 17164 4087 17204 4096
rect 17068 559 17108 568
rect 17164 2624 17204 2633
rect 16491 356 16533 365
rect 16491 316 16492 356
rect 16532 316 16533 356
rect 16491 307 16533 316
rect 15724 223 15764 232
rect 13612 139 13652 148
rect 10828 55 10868 64
rect 17164 104 17204 2584
rect 17260 272 17300 39544
rect 17356 37904 17396 40300
rect 17644 38996 17684 40804
rect 17932 40088 17972 41560
rect 17932 40039 17972 40048
rect 18508 41600 18548 41609
rect 17644 38947 17684 38956
rect 18219 38744 18261 38753
rect 18219 38704 18220 38744
rect 18260 38704 18261 38744
rect 18219 38695 18261 38704
rect 18220 38610 18260 38695
rect 17356 37855 17396 37864
rect 18124 37400 18164 37409
rect 17644 35216 17684 35225
rect 17452 33032 17492 33041
rect 17452 32360 17492 32992
rect 17452 32311 17492 32320
rect 17548 29840 17588 29849
rect 17356 24800 17396 24809
rect 17356 18332 17396 24760
rect 17356 18283 17396 18292
rect 17452 21608 17492 21617
rect 17355 12620 17397 12629
rect 17355 12580 17356 12620
rect 17396 12580 17397 12620
rect 17355 12571 17397 12580
rect 17356 2540 17396 12571
rect 17452 10940 17492 21568
rect 17548 18584 17588 29800
rect 17644 26900 17684 35176
rect 17740 29924 17780 29933
rect 17740 27488 17780 29884
rect 17740 27439 17780 27448
rect 17836 29840 17876 29849
rect 17836 28328 17876 29800
rect 17644 26851 17684 26860
rect 17740 26060 17780 26069
rect 17644 23960 17684 23969
rect 17644 20768 17684 23920
rect 17644 20719 17684 20728
rect 17740 23792 17780 26020
rect 17548 18535 17588 18544
rect 17452 10891 17492 10900
rect 17644 14888 17684 14897
rect 17644 9344 17684 14848
rect 17740 12377 17780 23752
rect 17836 21020 17876 28288
rect 18028 28328 18068 28337
rect 17836 20971 17876 20980
rect 17932 23708 17972 23717
rect 17932 19256 17972 23668
rect 17932 19207 17972 19216
rect 17836 17324 17876 17333
rect 17836 13544 17876 17284
rect 17876 13504 17972 13544
rect 17836 13495 17876 13504
rect 17739 12368 17781 12377
rect 17739 12328 17740 12368
rect 17780 12328 17781 12368
rect 17739 12319 17781 12328
rect 17740 12200 17780 12209
rect 17740 11108 17780 12160
rect 17740 11059 17780 11068
rect 17836 12116 17876 12125
rect 17836 11696 17876 12076
rect 17452 6740 17492 6749
rect 17452 4976 17492 6700
rect 17644 5984 17684 9304
rect 17644 5935 17684 5944
rect 17740 9512 17780 9521
rect 17452 2708 17492 4936
rect 17740 4976 17780 9472
rect 17740 4927 17780 4936
rect 17644 4472 17684 4481
rect 17644 3380 17684 4432
rect 17644 3331 17684 3340
rect 17452 2659 17492 2668
rect 17356 2500 17588 2540
rect 17548 1280 17588 2500
rect 17548 1231 17588 1240
rect 17836 1028 17876 11656
rect 17932 11192 17972 13504
rect 17932 11143 17972 11152
rect 17836 979 17876 988
rect 17932 6236 17972 6245
rect 17932 3128 17972 6196
rect 18028 4892 18068 28288
rect 18124 28244 18164 37360
rect 18508 36560 18548 41560
rect 18700 40256 18740 42148
rect 20048 41600 20416 41609
rect 20088 41560 20130 41600
rect 20170 41560 20212 41600
rect 20252 41560 20294 41600
rect 20334 41560 20376 41600
rect 20048 41551 20416 41560
rect 19756 41180 19796 41189
rect 18808 40844 19176 40853
rect 18848 40804 18890 40844
rect 18930 40804 18972 40844
rect 19012 40804 19054 40844
rect 19094 40804 19136 40844
rect 18808 40795 19176 40804
rect 18891 40508 18933 40517
rect 18891 40468 18892 40508
rect 18932 40468 18933 40508
rect 18891 40459 18933 40468
rect 19660 40508 19700 40517
rect 18892 40374 18932 40459
rect 18700 40207 18740 40216
rect 18808 39332 19176 39341
rect 18848 39292 18890 39332
rect 18930 39292 18972 39332
rect 19012 39292 19054 39332
rect 19094 39292 19136 39332
rect 18808 39283 19176 39292
rect 18988 38744 19028 38755
rect 18988 38669 19028 38704
rect 18987 38660 19029 38669
rect 18987 38620 18988 38660
rect 19028 38620 19029 38660
rect 18987 38611 19029 38620
rect 18699 38408 18741 38417
rect 18699 38368 18700 38408
rect 18740 38368 18741 38408
rect 18699 38359 18741 38368
rect 18508 36511 18548 36520
rect 18124 28195 18164 28204
rect 18220 35804 18260 35813
rect 18220 26732 18260 35764
rect 18508 34208 18548 34217
rect 18412 33452 18452 33461
rect 18316 29336 18356 29345
rect 18316 28916 18356 29296
rect 18316 28867 18356 28876
rect 18412 28664 18452 33412
rect 18412 28615 18452 28624
rect 18508 28328 18548 34168
rect 18604 33620 18644 33629
rect 18604 31184 18644 33580
rect 18604 31135 18644 31144
rect 18508 28279 18548 28288
rect 18604 30680 18644 30689
rect 18220 26683 18260 26692
rect 18316 28244 18356 28253
rect 18316 23876 18356 28204
rect 18604 26564 18644 30640
rect 18604 26515 18644 26524
rect 18124 21020 18164 21029
rect 18124 10352 18164 20980
rect 18316 18500 18356 23836
rect 18124 10303 18164 10312
rect 18220 16988 18260 16997
rect 18220 10772 18260 16948
rect 18316 12620 18356 18460
rect 18604 18584 18644 18593
rect 18604 17996 18644 18544
rect 18604 17947 18644 17956
rect 18412 17156 18452 17165
rect 18412 16652 18452 17116
rect 18412 16603 18452 16612
rect 18604 16820 18644 16829
rect 18604 15896 18644 16780
rect 18316 12571 18356 12580
rect 18412 14804 18452 14813
rect 18028 3296 18068 4852
rect 18028 3247 18068 3256
rect 18124 8336 18164 8345
rect 17932 860 17972 3088
rect 18124 2036 18164 8296
rect 18220 3464 18260 10732
rect 18412 10352 18452 14764
rect 18508 12704 18548 12713
rect 18508 11696 18548 12664
rect 18508 11647 18548 11656
rect 18412 10303 18452 10312
rect 18508 11444 18548 11453
rect 18412 9428 18452 9437
rect 18316 8588 18356 8597
rect 18316 6068 18356 8548
rect 18316 3800 18356 6028
rect 18412 5984 18452 9388
rect 18508 6152 18548 11404
rect 18604 9260 18644 15856
rect 18604 9211 18644 9220
rect 18508 6103 18548 6112
rect 18412 5935 18452 5944
rect 18316 3751 18356 3760
rect 18220 3415 18260 3424
rect 18124 1987 18164 1996
rect 18123 1448 18165 1457
rect 18123 1408 18124 1448
rect 18164 1408 18165 1448
rect 18123 1399 18165 1408
rect 18124 944 18164 1399
rect 18700 1280 18740 38359
rect 18808 37820 19176 37829
rect 18848 37780 18890 37820
rect 18930 37780 18972 37820
rect 19012 37780 19054 37820
rect 19094 37780 19136 37820
rect 18808 37771 19176 37780
rect 19660 37316 19700 40468
rect 19660 37267 19700 37276
rect 18808 36308 19176 36317
rect 18848 36268 18890 36308
rect 18930 36268 18972 36308
rect 19012 36268 19054 36308
rect 19094 36268 19136 36308
rect 18808 36259 19176 36268
rect 18808 34796 19176 34805
rect 18848 34756 18890 34796
rect 18930 34756 18972 34796
rect 19012 34756 19054 34796
rect 19094 34756 19136 34796
rect 18808 34747 19176 34756
rect 19564 34208 19604 34217
rect 18808 33284 19176 33293
rect 18848 33244 18890 33284
rect 18930 33244 18972 33284
rect 19012 33244 19054 33284
rect 19094 33244 19136 33284
rect 18808 33235 19176 33244
rect 19564 32360 19604 34168
rect 19564 32311 19604 32320
rect 19660 33116 19700 33125
rect 18808 31772 19176 31781
rect 18848 31732 18890 31772
rect 18930 31732 18972 31772
rect 19012 31732 19054 31772
rect 19094 31732 19136 31772
rect 18808 31723 19176 31732
rect 19276 31184 19316 31193
rect 18808 30260 19176 30269
rect 18848 30220 18890 30260
rect 18930 30220 18972 30260
rect 19012 30220 19054 30260
rect 19094 30220 19136 30260
rect 18808 30211 19176 30220
rect 18808 28748 19176 28757
rect 18848 28708 18890 28748
rect 18930 28708 18972 28748
rect 19012 28708 19054 28748
rect 19094 28708 19136 28748
rect 18808 28699 19176 28708
rect 19276 28412 19316 31144
rect 19660 30344 19700 33076
rect 19660 30295 19700 30304
rect 19276 28363 19316 28372
rect 18808 27236 19176 27245
rect 18848 27196 18890 27236
rect 18930 27196 18972 27236
rect 19012 27196 19054 27236
rect 19094 27196 19136 27236
rect 18808 27187 19176 27196
rect 18808 25724 19176 25733
rect 18848 25684 18890 25724
rect 18930 25684 18972 25724
rect 19012 25684 19054 25724
rect 19094 25684 19136 25724
rect 18808 25675 19176 25684
rect 18808 24212 19176 24221
rect 18848 24172 18890 24212
rect 18930 24172 18972 24212
rect 19012 24172 19054 24212
rect 19094 24172 19136 24212
rect 18808 24163 19176 24172
rect 19275 23036 19317 23045
rect 19275 22996 19276 23036
rect 19316 22996 19317 23036
rect 19275 22987 19317 22996
rect 18808 22700 19176 22709
rect 18848 22660 18890 22700
rect 18930 22660 18972 22700
rect 19012 22660 19054 22700
rect 19094 22660 19136 22700
rect 18808 22651 19176 22660
rect 18808 21188 19176 21197
rect 18848 21148 18890 21188
rect 18930 21148 18972 21188
rect 19012 21148 19054 21188
rect 19094 21148 19136 21188
rect 18808 21139 19176 21148
rect 18808 19676 19176 19685
rect 18848 19636 18890 19676
rect 18930 19636 18972 19676
rect 19012 19636 19054 19676
rect 19094 19636 19136 19676
rect 18808 19627 19176 19636
rect 19276 18836 19316 22987
rect 19276 18787 19316 18796
rect 19660 20096 19700 20105
rect 18808 18164 19176 18173
rect 18848 18124 18890 18164
rect 18930 18124 18972 18164
rect 19012 18124 19054 18164
rect 19094 18124 19136 18164
rect 18808 18115 19176 18124
rect 19276 17912 19316 17921
rect 18808 16652 19176 16661
rect 18848 16612 18890 16652
rect 18930 16612 18972 16652
rect 19012 16612 19054 16652
rect 19094 16612 19136 16652
rect 18808 16603 19176 16612
rect 19276 16568 19316 17872
rect 19660 17828 19700 20056
rect 19660 17660 19700 17788
rect 19660 17611 19700 17620
rect 19276 16519 19316 16528
rect 19468 17576 19508 17585
rect 18808 15140 19176 15149
rect 18848 15100 18890 15140
rect 18930 15100 18972 15140
rect 19012 15100 19054 15140
rect 19094 15100 19136 15140
rect 18808 15091 19176 15100
rect 19468 14720 19508 17536
rect 19468 14671 19508 14680
rect 18808 13628 19176 13637
rect 18848 13588 18890 13628
rect 18930 13588 18972 13628
rect 19012 13588 19054 13628
rect 19094 13588 19136 13628
rect 18808 13579 19176 13588
rect 18808 12116 19176 12125
rect 18848 12076 18890 12116
rect 18930 12076 18972 12116
rect 19012 12076 19054 12116
rect 19094 12076 19136 12116
rect 18808 12067 19176 12076
rect 19756 10688 19796 41140
rect 19852 41096 19892 41105
rect 19852 40340 19892 41056
rect 19852 40291 19892 40300
rect 20048 40088 20416 40097
rect 20088 40048 20130 40088
rect 20170 40048 20212 40088
rect 20252 40048 20294 40088
rect 20334 40048 20376 40088
rect 20048 40039 20416 40048
rect 20048 38576 20416 38585
rect 20088 38536 20130 38576
rect 20170 38536 20212 38576
rect 20252 38536 20294 38576
rect 20334 38536 20376 38576
rect 20048 38527 20416 38536
rect 20139 38324 20181 38333
rect 20139 38284 20140 38324
rect 20180 38284 20181 38324
rect 20139 38275 20181 38284
rect 20140 38190 20180 38275
rect 20048 37064 20416 37073
rect 20088 37024 20130 37064
rect 20170 37024 20212 37064
rect 20252 37024 20294 37064
rect 20334 37024 20376 37064
rect 20048 37015 20416 37024
rect 19948 35972 19988 35981
rect 19948 35216 19988 35932
rect 20048 35552 20416 35561
rect 20088 35512 20130 35552
rect 20170 35512 20212 35552
rect 20252 35512 20294 35552
rect 20334 35512 20376 35552
rect 20048 35503 20416 35512
rect 20620 35468 20660 42736
rect 20812 41432 20852 41441
rect 20812 39752 20852 41392
rect 20812 39703 20852 39712
rect 20620 35419 20660 35428
rect 21004 36812 21044 36821
rect 19948 35167 19988 35176
rect 20048 34040 20416 34049
rect 20088 34000 20130 34040
rect 20170 34000 20212 34040
rect 20252 34000 20294 34040
rect 20334 34000 20376 34040
rect 20048 33991 20416 34000
rect 20812 33452 20852 33461
rect 19852 33200 19892 33209
rect 19852 31520 19892 33160
rect 19852 31471 19892 31480
rect 19948 32780 19988 32789
rect 19852 31352 19892 31361
rect 19852 23960 19892 31312
rect 19948 30680 19988 32740
rect 20048 32528 20416 32537
rect 20088 32488 20130 32528
rect 20170 32488 20212 32528
rect 20252 32488 20294 32528
rect 20334 32488 20376 32528
rect 20048 32479 20416 32488
rect 20524 31520 20564 31529
rect 20048 31016 20416 31025
rect 20088 30976 20130 31016
rect 20170 30976 20212 31016
rect 20252 30976 20294 31016
rect 20334 30976 20376 31016
rect 20048 30967 20416 30976
rect 19948 30631 19988 30640
rect 19948 30260 19988 30269
rect 19948 27740 19988 30220
rect 20048 29504 20416 29513
rect 20088 29464 20130 29504
rect 20170 29464 20212 29504
rect 20252 29464 20294 29504
rect 20334 29464 20376 29504
rect 20048 29455 20416 29464
rect 20048 27992 20416 28001
rect 20088 27952 20130 27992
rect 20170 27952 20212 27992
rect 20252 27952 20294 27992
rect 20334 27952 20376 27992
rect 20048 27943 20416 27952
rect 19948 27691 19988 27700
rect 20048 26480 20416 26489
rect 20088 26440 20130 26480
rect 20170 26440 20212 26480
rect 20252 26440 20294 26480
rect 20334 26440 20376 26480
rect 20048 26431 20416 26440
rect 20048 24968 20416 24977
rect 20088 24928 20130 24968
rect 20170 24928 20212 24968
rect 20252 24928 20294 24968
rect 20334 24928 20376 24968
rect 20048 24919 20416 24928
rect 19852 23911 19892 23920
rect 20048 23456 20416 23465
rect 20088 23416 20130 23456
rect 20170 23416 20212 23456
rect 20252 23416 20294 23456
rect 20334 23416 20376 23456
rect 20048 23407 20416 23416
rect 20048 21944 20416 21953
rect 20088 21904 20130 21944
rect 20170 21904 20212 21944
rect 20252 21904 20294 21944
rect 20334 21904 20376 21944
rect 20048 21895 20416 21904
rect 20048 20432 20416 20441
rect 20088 20392 20130 20432
rect 20170 20392 20212 20432
rect 20252 20392 20294 20432
rect 20334 20392 20376 20432
rect 20048 20383 20416 20392
rect 20048 18920 20416 18929
rect 20088 18880 20130 18920
rect 20170 18880 20212 18920
rect 20252 18880 20294 18920
rect 20334 18880 20376 18920
rect 20048 18871 20416 18880
rect 20048 17408 20416 17417
rect 20088 17368 20130 17408
rect 20170 17368 20212 17408
rect 20252 17368 20294 17408
rect 20334 17368 20376 17408
rect 20048 17359 20416 17368
rect 20048 15896 20416 15905
rect 20088 15856 20130 15896
rect 20170 15856 20212 15896
rect 20252 15856 20294 15896
rect 20334 15856 20376 15896
rect 20048 15847 20416 15856
rect 20048 14384 20416 14393
rect 20088 14344 20130 14384
rect 20170 14344 20212 14384
rect 20252 14344 20294 14384
rect 20334 14344 20376 14384
rect 20048 14335 20416 14344
rect 20048 12872 20416 12881
rect 20088 12832 20130 12872
rect 20170 12832 20212 12872
rect 20252 12832 20294 12872
rect 20334 12832 20376 12872
rect 20048 12823 20416 12832
rect 20048 11360 20416 11369
rect 20088 11320 20130 11360
rect 20170 11320 20212 11360
rect 20252 11320 20294 11360
rect 20334 11320 20376 11360
rect 20048 11311 20416 11320
rect 19756 10639 19796 10648
rect 18808 10604 19176 10613
rect 18848 10564 18890 10604
rect 18930 10564 18972 10604
rect 19012 10564 19054 10604
rect 19094 10564 19136 10604
rect 18808 10555 19176 10564
rect 20048 9848 20416 9857
rect 20088 9808 20130 9848
rect 20170 9808 20212 9848
rect 20252 9808 20294 9848
rect 20334 9808 20376 9848
rect 20048 9799 20416 9808
rect 18808 9092 19176 9101
rect 18848 9052 18890 9092
rect 18930 9052 18972 9092
rect 19012 9052 19054 9092
rect 19094 9052 19136 9092
rect 18808 9043 19176 9052
rect 20048 8336 20416 8345
rect 20088 8296 20130 8336
rect 20170 8296 20212 8336
rect 20252 8296 20294 8336
rect 20334 8296 20376 8336
rect 20048 8287 20416 8296
rect 19084 7757 19124 7842
rect 19083 7748 19125 7757
rect 19083 7708 19084 7748
rect 19124 7708 19125 7748
rect 19083 7699 19125 7708
rect 18808 7580 19176 7589
rect 18848 7540 18890 7580
rect 18930 7540 18972 7580
rect 19012 7540 19054 7580
rect 19094 7540 19136 7580
rect 18808 7531 19176 7540
rect 19467 7076 19509 7085
rect 19467 7036 19468 7076
rect 19508 7036 19509 7076
rect 19467 7027 19509 7036
rect 19275 6992 19317 7001
rect 19275 6952 19276 6992
rect 19316 6952 19317 6992
rect 19275 6943 19317 6952
rect 18808 6068 19176 6077
rect 18848 6028 18890 6068
rect 18930 6028 18972 6068
rect 19012 6028 19054 6068
rect 19094 6028 19136 6068
rect 18808 6019 19176 6028
rect 18808 4556 19176 4565
rect 18848 4516 18890 4556
rect 18930 4516 18972 4556
rect 19012 4516 19054 4556
rect 19094 4516 19136 4556
rect 18808 4507 19176 4516
rect 18808 3044 19176 3053
rect 18848 3004 18890 3044
rect 18930 3004 18972 3044
rect 19012 3004 19054 3044
rect 19094 3004 19136 3044
rect 18808 2995 19176 3004
rect 18808 1532 19176 1541
rect 18848 1492 18890 1532
rect 18930 1492 18972 1532
rect 19012 1492 19054 1532
rect 19094 1492 19136 1532
rect 18808 1483 19176 1492
rect 18700 1231 18740 1240
rect 18124 895 18164 904
rect 19276 944 19316 6943
rect 19372 4556 19412 4565
rect 19372 4388 19412 4516
rect 19372 4339 19412 4348
rect 19468 1280 19508 7027
rect 20524 7001 20564 31480
rect 20812 29336 20852 33412
rect 20812 29287 20852 29296
rect 21004 29000 21044 36772
rect 21196 36560 21236 36569
rect 21196 31016 21236 36520
rect 21196 30967 21236 30976
rect 21004 28951 21044 28960
rect 20620 22028 20660 22037
rect 20620 7085 20660 21988
rect 20716 15644 20756 15653
rect 20716 10520 20756 15604
rect 20811 15308 20853 15317
rect 20811 15268 20812 15308
rect 20852 15268 20853 15308
rect 20811 15259 20853 15268
rect 20812 15224 20852 15259
rect 20812 15173 20852 15184
rect 20716 10471 20756 10480
rect 20619 7076 20661 7085
rect 20619 7036 20620 7076
rect 20660 7036 20661 7076
rect 20619 7027 20661 7036
rect 20523 6992 20565 7001
rect 20523 6952 20524 6992
rect 20564 6952 20565 6992
rect 20523 6943 20565 6952
rect 20048 6824 20416 6833
rect 20088 6784 20130 6824
rect 20170 6784 20212 6824
rect 20252 6784 20294 6824
rect 20334 6784 20376 6824
rect 20048 6775 20416 6784
rect 20048 5312 20416 5321
rect 20088 5272 20130 5312
rect 20170 5272 20212 5312
rect 20252 5272 20294 5312
rect 20334 5272 20376 5312
rect 20048 5263 20416 5272
rect 20048 3800 20416 3809
rect 20088 3760 20130 3800
rect 20170 3760 20212 3800
rect 20252 3760 20294 3800
rect 20334 3760 20376 3800
rect 20048 3751 20416 3760
rect 20907 3296 20949 3305
rect 20907 3256 20908 3296
rect 20948 3256 20949 3296
rect 20907 3247 20949 3256
rect 20811 3212 20853 3221
rect 20811 3172 20812 3212
rect 20852 3172 20853 3212
rect 20811 3163 20853 3172
rect 20812 3128 20852 3163
rect 20812 3077 20852 3088
rect 20048 2288 20416 2297
rect 20088 2248 20130 2288
rect 20170 2248 20212 2288
rect 20252 2248 20294 2288
rect 20334 2248 20376 2288
rect 20048 2239 20416 2248
rect 20908 1784 20948 3247
rect 20908 1735 20948 1744
rect 19468 1231 19508 1240
rect 19276 895 19316 904
rect 17932 811 17972 820
rect 20048 776 20416 785
rect 20088 736 20130 776
rect 20170 736 20212 776
rect 20252 736 20294 776
rect 20334 736 20376 776
rect 20048 727 20416 736
rect 17260 223 17300 232
rect 17164 55 17204 64
<< via4 >>
rect 460 19972 500 20012
rect 556 16276 596 16316
rect 460 16108 500 16148
rect 172 7708 212 7748
rect 748 19972 788 20012
rect 940 6952 980 6992
rect 1228 19048 1268 19088
rect 1228 12328 1268 12368
rect 1228 4768 1268 4808
rect 2572 38032 2612 38072
rect 3688 40804 3728 40844
rect 3770 40804 3810 40844
rect 3852 40804 3892 40844
rect 3934 40804 3974 40844
rect 4016 40804 4056 40844
rect 2956 38032 2996 38072
rect 1996 400 2036 440
rect 3688 39292 3728 39332
rect 3770 39292 3810 39332
rect 3852 39292 3892 39332
rect 3934 39292 3974 39332
rect 4016 39292 4056 39332
rect 3340 38200 3380 38240
rect 3688 37780 3728 37820
rect 3770 37780 3810 37820
rect 3852 37780 3892 37820
rect 3934 37780 3974 37820
rect 4016 37780 4056 37820
rect 3688 36268 3728 36308
rect 3770 36268 3810 36308
rect 3852 36268 3892 36308
rect 3934 36268 3974 36308
rect 4016 36268 4056 36308
rect 4928 41560 4968 41600
rect 5010 41560 5050 41600
rect 5092 41560 5132 41600
rect 5174 41560 5214 41600
rect 5256 41560 5296 41600
rect 4928 40048 4968 40088
rect 5010 40048 5050 40088
rect 5092 40048 5132 40088
rect 5174 40048 5214 40088
rect 5256 40048 5296 40088
rect 4928 38536 4968 38576
rect 5010 38536 5050 38576
rect 5092 38536 5132 38576
rect 5174 38536 5214 38576
rect 5256 38536 5296 38576
rect 4928 37024 4968 37064
rect 5010 37024 5050 37064
rect 5092 37024 5132 37064
rect 5174 37024 5214 37064
rect 5256 37024 5296 37064
rect 3688 34756 3728 34796
rect 3770 34756 3810 34796
rect 3852 34756 3892 34796
rect 3934 34756 3974 34796
rect 4016 34756 4056 34796
rect 3688 33244 3728 33284
rect 3770 33244 3810 33284
rect 3852 33244 3892 33284
rect 3934 33244 3974 33284
rect 4016 33244 4056 33284
rect 3724 32908 3764 32948
rect 3688 31732 3728 31772
rect 3770 31732 3810 31772
rect 3852 31732 3892 31772
rect 3934 31732 3974 31772
rect 4016 31732 4056 31772
rect 3688 30220 3728 30260
rect 3770 30220 3810 30260
rect 3852 30220 3892 30260
rect 3934 30220 3974 30260
rect 4016 30220 4056 30260
rect 3688 28708 3728 28748
rect 3770 28708 3810 28748
rect 3852 28708 3892 28748
rect 3934 28708 3974 28748
rect 4016 28708 4056 28748
rect 3688 27196 3728 27236
rect 3770 27196 3810 27236
rect 3852 27196 3892 27236
rect 3934 27196 3974 27236
rect 4016 27196 4056 27236
rect 3688 25684 3728 25724
rect 3770 25684 3810 25724
rect 3852 25684 3892 25724
rect 3934 25684 3974 25724
rect 4016 25684 4056 25724
rect 3688 24172 3728 24212
rect 3770 24172 3810 24212
rect 3852 24172 3892 24212
rect 3934 24172 3974 24212
rect 4016 24172 4056 24212
rect 3688 22660 3728 22700
rect 3770 22660 3810 22700
rect 3852 22660 3892 22700
rect 3934 22660 3974 22700
rect 4016 22660 4056 22700
rect 3688 21148 3728 21188
rect 3770 21148 3810 21188
rect 3852 21148 3892 21188
rect 3934 21148 3974 21188
rect 4016 21148 4056 21188
rect 3688 19636 3728 19676
rect 3770 19636 3810 19676
rect 3852 19636 3892 19676
rect 3934 19636 3974 19676
rect 4016 19636 4056 19676
rect 3688 18124 3728 18164
rect 3770 18124 3810 18164
rect 3852 18124 3892 18164
rect 3934 18124 3974 18164
rect 4016 18124 4056 18164
rect 3688 16612 3728 16652
rect 3770 16612 3810 16652
rect 3852 16612 3892 16652
rect 3934 16612 3974 16652
rect 4016 16612 4056 16652
rect 3688 15100 3728 15140
rect 3770 15100 3810 15140
rect 3852 15100 3892 15140
rect 3934 15100 3974 15140
rect 4016 15100 4056 15140
rect 3688 13588 3728 13628
rect 3770 13588 3810 13628
rect 3852 13588 3892 13628
rect 3934 13588 3974 13628
rect 4016 13588 4056 13628
rect 3688 12076 3728 12116
rect 3770 12076 3810 12116
rect 3852 12076 3892 12116
rect 3934 12076 3974 12116
rect 4016 12076 4056 12116
rect 3688 10564 3728 10604
rect 3770 10564 3810 10604
rect 3852 10564 3892 10604
rect 3934 10564 3974 10604
rect 4016 10564 4056 10604
rect 4108 10144 4148 10184
rect 3628 9388 3668 9428
rect 4300 9388 4340 9428
rect 3688 9052 3728 9092
rect 3770 9052 3810 9092
rect 3852 9052 3892 9092
rect 3934 9052 3974 9092
rect 4016 9052 4056 9092
rect 3688 7540 3728 7580
rect 3770 7540 3810 7580
rect 3852 7540 3892 7580
rect 3934 7540 3974 7580
rect 4016 7540 4056 7580
rect 3688 6028 3728 6068
rect 3770 6028 3810 6068
rect 3852 6028 3892 6068
rect 3934 6028 3974 6068
rect 4016 6028 4056 6068
rect 3688 4516 3728 4556
rect 3770 4516 3810 4556
rect 3852 4516 3892 4556
rect 3934 4516 3974 4556
rect 4016 4516 4056 4556
rect 4928 35512 4968 35552
rect 5010 35512 5050 35552
rect 5092 35512 5132 35552
rect 5174 35512 5214 35552
rect 5256 35512 5296 35552
rect 4928 34000 4968 34040
rect 5010 34000 5050 34040
rect 5092 34000 5132 34040
rect 5174 34000 5214 34040
rect 5256 34000 5296 34040
rect 4928 32488 4968 32528
rect 5010 32488 5050 32528
rect 5092 32488 5132 32528
rect 5174 32488 5214 32528
rect 5256 32488 5296 32528
rect 4928 30976 4968 31016
rect 5010 30976 5050 31016
rect 5092 30976 5132 31016
rect 5174 30976 5214 31016
rect 5256 30976 5296 31016
rect 4684 19468 4724 19508
rect 4928 29464 4968 29504
rect 5010 29464 5050 29504
rect 5092 29464 5132 29504
rect 5174 29464 5214 29504
rect 5256 29464 5296 29504
rect 4928 27952 4968 27992
rect 5010 27952 5050 27992
rect 5092 27952 5132 27992
rect 5174 27952 5214 27992
rect 5256 27952 5296 27992
rect 4928 26440 4968 26480
rect 5010 26440 5050 26480
rect 5092 26440 5132 26480
rect 5174 26440 5214 26480
rect 5256 26440 5296 26480
rect 4928 24928 4968 24968
rect 5010 24928 5050 24968
rect 5092 24928 5132 24968
rect 5174 24928 5214 24968
rect 5256 24928 5296 24968
rect 4928 23416 4968 23456
rect 5010 23416 5050 23456
rect 5092 23416 5132 23456
rect 5174 23416 5214 23456
rect 5256 23416 5296 23456
rect 4928 21904 4968 21944
rect 5010 21904 5050 21944
rect 5092 21904 5132 21944
rect 5174 21904 5214 21944
rect 5256 21904 5296 21944
rect 4928 20392 4968 20432
rect 5010 20392 5050 20432
rect 5092 20392 5132 20432
rect 5174 20392 5214 20432
rect 5256 20392 5296 20432
rect 4928 18880 4968 18920
rect 5010 18880 5050 18920
rect 5092 18880 5132 18920
rect 5174 18880 5214 18920
rect 5256 18880 5296 18920
rect 4928 17368 4968 17408
rect 5010 17368 5050 17408
rect 5092 17368 5132 17408
rect 5174 17368 5214 17408
rect 5256 17368 5296 17408
rect 5068 16108 5108 16148
rect 4928 15856 4968 15896
rect 5010 15856 5050 15896
rect 5092 15856 5132 15896
rect 5174 15856 5214 15896
rect 5256 15856 5296 15896
rect 4780 15268 4820 15308
rect 4684 14512 4724 14552
rect 4588 10144 4628 10184
rect 4928 14344 4968 14384
rect 5010 14344 5050 14384
rect 5092 14344 5132 14384
rect 5174 14344 5214 14384
rect 5256 14344 5296 14384
rect 4928 12832 4968 12872
rect 5010 12832 5050 12872
rect 5092 12832 5132 12872
rect 5174 12832 5214 12872
rect 5256 12832 5296 12872
rect 4928 11320 4968 11360
rect 5010 11320 5050 11360
rect 5092 11320 5132 11360
rect 5174 11320 5214 11360
rect 5256 11320 5296 11360
rect 5740 11740 5780 11780
rect 4928 9808 4968 9848
rect 5010 9808 5050 9848
rect 5092 9808 5132 9848
rect 5174 9808 5214 9848
rect 5256 9808 5296 9848
rect 4928 8296 4968 8336
rect 5010 8296 5050 8336
rect 5092 8296 5132 8336
rect 5174 8296 5214 8336
rect 5256 8296 5296 8336
rect 4928 6784 4968 6824
rect 5010 6784 5050 6824
rect 5092 6784 5132 6824
rect 5174 6784 5214 6824
rect 5256 6784 5296 6824
rect 5452 6112 5492 6152
rect 5356 5944 5396 5984
rect 4928 5272 4968 5312
rect 5010 5272 5050 5312
rect 5092 5272 5132 5312
rect 5174 5272 5214 5312
rect 5256 5272 5296 5312
rect 4928 3760 4968 3800
rect 5010 3760 5050 3800
rect 5092 3760 5132 3800
rect 5174 3760 5214 3800
rect 5256 3760 5296 3800
rect 3916 3256 3956 3296
rect 4588 3256 4628 3296
rect 3688 3004 3728 3044
rect 3770 3004 3810 3044
rect 3852 3004 3892 3044
rect 3934 3004 3974 3044
rect 4016 3004 4056 3044
rect 4928 2248 4968 2288
rect 5010 2248 5050 2288
rect 5092 2248 5132 2288
rect 5174 2248 5214 2288
rect 5256 2248 5296 2288
rect 3688 1492 3728 1532
rect 3770 1492 3810 1532
rect 3852 1492 3892 1532
rect 3934 1492 3974 1532
rect 4016 1492 4056 1532
rect 4108 1324 4148 1364
rect 4684 1240 4724 1280
rect 4928 736 4968 776
rect 5010 736 5050 776
rect 5092 736 5132 776
rect 5174 736 5214 776
rect 5256 736 5296 776
rect 5644 6448 5684 6488
rect 6220 11740 6260 11780
rect 5932 4180 5972 4220
rect 6028 3172 6068 3212
rect 5548 2248 5588 2288
rect 6892 3676 6932 3716
rect 6700 2332 6740 2372
rect 6412 400 6452 440
rect 7084 22996 7124 23036
rect 7564 9388 7604 9428
rect 7468 1828 7508 1868
rect 7852 2332 7892 2372
rect 8812 9304 8852 9344
rect 9580 38200 9620 38240
rect 8908 6112 8948 6152
rect 8716 3760 8756 3800
rect 8620 1828 8660 1868
rect 8428 1240 8468 1280
rect 9580 32908 9620 32948
rect 9580 4180 9620 4220
rect 10252 38032 10292 38072
rect 10156 10480 10196 10520
rect 9868 6448 9908 6488
rect 9772 5944 9812 5984
rect 9676 1324 9716 1364
rect 10444 10480 10484 10520
rect 11020 15436 11060 15476
rect 10924 9304 10964 9344
rect 7948 904 7988 944
rect 8140 568 8180 608
rect 11692 15436 11732 15476
rect 11500 904 11540 944
rect 12844 38368 12884 38408
rect 12556 15436 12596 15476
rect 12364 1408 12404 1448
rect 13708 38620 13748 38660
rect 13516 12580 13556 12620
rect 13420 6952 13460 6992
rect 13516 988 13556 1028
rect 12940 568 12980 608
rect 13996 4768 14036 4808
rect 13804 3676 13844 3716
rect 13900 2248 13940 2288
rect 14188 3760 14228 3800
rect 14764 16612 14804 16652
rect 14284 820 14324 860
rect 13708 736 13748 776
rect 15052 38704 15092 38744
rect 14956 16612 14996 16652
rect 14956 14512 14996 14552
rect 15148 988 15188 1028
rect 15628 5776 15668 5816
rect 14092 316 14132 356
rect 17164 39796 17204 39836
rect 16492 19048 16532 19088
rect 16396 10144 16436 10184
rect 16012 736 16052 776
rect 16972 19468 17012 19508
rect 17068 16360 17108 16400
rect 16492 316 16532 356
rect 18220 38704 18260 38744
rect 17356 12580 17396 12620
rect 17740 12328 17780 12368
rect 20048 41560 20088 41600
rect 20130 41560 20170 41600
rect 20212 41560 20252 41600
rect 20294 41560 20334 41600
rect 20376 41560 20416 41600
rect 18808 40804 18848 40844
rect 18890 40804 18930 40844
rect 18972 40804 19012 40844
rect 19054 40804 19094 40844
rect 19136 40804 19176 40844
rect 18892 40468 18932 40508
rect 18808 39292 18848 39332
rect 18890 39292 18930 39332
rect 18972 39292 19012 39332
rect 19054 39292 19094 39332
rect 19136 39292 19176 39332
rect 18988 38620 19028 38660
rect 18700 38368 18740 38408
rect 18124 1408 18164 1448
rect 18808 37780 18848 37820
rect 18890 37780 18930 37820
rect 18972 37780 19012 37820
rect 19054 37780 19094 37820
rect 19136 37780 19176 37820
rect 18808 36268 18848 36308
rect 18890 36268 18930 36308
rect 18972 36268 19012 36308
rect 19054 36268 19094 36308
rect 19136 36268 19176 36308
rect 18808 34756 18848 34796
rect 18890 34756 18930 34796
rect 18972 34756 19012 34796
rect 19054 34756 19094 34796
rect 19136 34756 19176 34796
rect 18808 33244 18848 33284
rect 18890 33244 18930 33284
rect 18972 33244 19012 33284
rect 19054 33244 19094 33284
rect 19136 33244 19176 33284
rect 18808 31732 18848 31772
rect 18890 31732 18930 31772
rect 18972 31732 19012 31772
rect 19054 31732 19094 31772
rect 19136 31732 19176 31772
rect 18808 30220 18848 30260
rect 18890 30220 18930 30260
rect 18972 30220 19012 30260
rect 19054 30220 19094 30260
rect 19136 30220 19176 30260
rect 18808 28708 18848 28748
rect 18890 28708 18930 28748
rect 18972 28708 19012 28748
rect 19054 28708 19094 28748
rect 19136 28708 19176 28748
rect 18808 27196 18848 27236
rect 18890 27196 18930 27236
rect 18972 27196 19012 27236
rect 19054 27196 19094 27236
rect 19136 27196 19176 27236
rect 18808 25684 18848 25724
rect 18890 25684 18930 25724
rect 18972 25684 19012 25724
rect 19054 25684 19094 25724
rect 19136 25684 19176 25724
rect 18808 24172 18848 24212
rect 18890 24172 18930 24212
rect 18972 24172 19012 24212
rect 19054 24172 19094 24212
rect 19136 24172 19176 24212
rect 19276 22996 19316 23036
rect 18808 22660 18848 22700
rect 18890 22660 18930 22700
rect 18972 22660 19012 22700
rect 19054 22660 19094 22700
rect 19136 22660 19176 22700
rect 18808 21148 18848 21188
rect 18890 21148 18930 21188
rect 18972 21148 19012 21188
rect 19054 21148 19094 21188
rect 19136 21148 19176 21188
rect 18808 19636 18848 19676
rect 18890 19636 18930 19676
rect 18972 19636 19012 19676
rect 19054 19636 19094 19676
rect 19136 19636 19176 19676
rect 18808 18124 18848 18164
rect 18890 18124 18930 18164
rect 18972 18124 19012 18164
rect 19054 18124 19094 18164
rect 19136 18124 19176 18164
rect 18808 16612 18848 16652
rect 18890 16612 18930 16652
rect 18972 16612 19012 16652
rect 19054 16612 19094 16652
rect 19136 16612 19176 16652
rect 18808 15100 18848 15140
rect 18890 15100 18930 15140
rect 18972 15100 19012 15140
rect 19054 15100 19094 15140
rect 19136 15100 19176 15140
rect 18808 13588 18848 13628
rect 18890 13588 18930 13628
rect 18972 13588 19012 13628
rect 19054 13588 19094 13628
rect 19136 13588 19176 13628
rect 18808 12076 18848 12116
rect 18890 12076 18930 12116
rect 18972 12076 19012 12116
rect 19054 12076 19094 12116
rect 19136 12076 19176 12116
rect 20048 40048 20088 40088
rect 20130 40048 20170 40088
rect 20212 40048 20252 40088
rect 20294 40048 20334 40088
rect 20376 40048 20416 40088
rect 20048 38536 20088 38576
rect 20130 38536 20170 38576
rect 20212 38536 20252 38576
rect 20294 38536 20334 38576
rect 20376 38536 20416 38576
rect 20140 38284 20180 38324
rect 20048 37024 20088 37064
rect 20130 37024 20170 37064
rect 20212 37024 20252 37064
rect 20294 37024 20334 37064
rect 20376 37024 20416 37064
rect 20048 35512 20088 35552
rect 20130 35512 20170 35552
rect 20212 35512 20252 35552
rect 20294 35512 20334 35552
rect 20376 35512 20416 35552
rect 20048 34000 20088 34040
rect 20130 34000 20170 34040
rect 20212 34000 20252 34040
rect 20294 34000 20334 34040
rect 20376 34000 20416 34040
rect 20048 32488 20088 32528
rect 20130 32488 20170 32528
rect 20212 32488 20252 32528
rect 20294 32488 20334 32528
rect 20376 32488 20416 32528
rect 20048 30976 20088 31016
rect 20130 30976 20170 31016
rect 20212 30976 20252 31016
rect 20294 30976 20334 31016
rect 20376 30976 20416 31016
rect 20048 29464 20088 29504
rect 20130 29464 20170 29504
rect 20212 29464 20252 29504
rect 20294 29464 20334 29504
rect 20376 29464 20416 29504
rect 20048 27952 20088 27992
rect 20130 27952 20170 27992
rect 20212 27952 20252 27992
rect 20294 27952 20334 27992
rect 20376 27952 20416 27992
rect 20048 26440 20088 26480
rect 20130 26440 20170 26480
rect 20212 26440 20252 26480
rect 20294 26440 20334 26480
rect 20376 26440 20416 26480
rect 20048 24928 20088 24968
rect 20130 24928 20170 24968
rect 20212 24928 20252 24968
rect 20294 24928 20334 24968
rect 20376 24928 20416 24968
rect 20048 23416 20088 23456
rect 20130 23416 20170 23456
rect 20212 23416 20252 23456
rect 20294 23416 20334 23456
rect 20376 23416 20416 23456
rect 20048 21904 20088 21944
rect 20130 21904 20170 21944
rect 20212 21904 20252 21944
rect 20294 21904 20334 21944
rect 20376 21904 20416 21944
rect 20048 20392 20088 20432
rect 20130 20392 20170 20432
rect 20212 20392 20252 20432
rect 20294 20392 20334 20432
rect 20376 20392 20416 20432
rect 20048 18880 20088 18920
rect 20130 18880 20170 18920
rect 20212 18880 20252 18920
rect 20294 18880 20334 18920
rect 20376 18880 20416 18920
rect 20048 17368 20088 17408
rect 20130 17368 20170 17408
rect 20212 17368 20252 17408
rect 20294 17368 20334 17408
rect 20376 17368 20416 17408
rect 20048 15856 20088 15896
rect 20130 15856 20170 15896
rect 20212 15856 20252 15896
rect 20294 15856 20334 15896
rect 20376 15856 20416 15896
rect 20048 14344 20088 14384
rect 20130 14344 20170 14384
rect 20212 14344 20252 14384
rect 20294 14344 20334 14384
rect 20376 14344 20416 14384
rect 20048 12832 20088 12872
rect 20130 12832 20170 12872
rect 20212 12832 20252 12872
rect 20294 12832 20334 12872
rect 20376 12832 20416 12872
rect 20048 11320 20088 11360
rect 20130 11320 20170 11360
rect 20212 11320 20252 11360
rect 20294 11320 20334 11360
rect 20376 11320 20416 11360
rect 18808 10564 18848 10604
rect 18890 10564 18930 10604
rect 18972 10564 19012 10604
rect 19054 10564 19094 10604
rect 19136 10564 19176 10604
rect 20048 9808 20088 9848
rect 20130 9808 20170 9848
rect 20212 9808 20252 9848
rect 20294 9808 20334 9848
rect 20376 9808 20416 9848
rect 18808 9052 18848 9092
rect 18890 9052 18930 9092
rect 18972 9052 19012 9092
rect 19054 9052 19094 9092
rect 19136 9052 19176 9092
rect 20048 8296 20088 8336
rect 20130 8296 20170 8336
rect 20212 8296 20252 8336
rect 20294 8296 20334 8336
rect 20376 8296 20416 8336
rect 19084 7708 19124 7748
rect 18808 7540 18848 7580
rect 18890 7540 18930 7580
rect 18972 7540 19012 7580
rect 19054 7540 19094 7580
rect 19136 7540 19176 7580
rect 19468 7036 19508 7076
rect 19276 6952 19316 6992
rect 18808 6028 18848 6068
rect 18890 6028 18930 6068
rect 18972 6028 19012 6068
rect 19054 6028 19094 6068
rect 19136 6028 19176 6068
rect 18808 4516 18848 4556
rect 18890 4516 18930 4556
rect 18972 4516 19012 4556
rect 19054 4516 19094 4556
rect 19136 4516 19176 4556
rect 18808 3004 18848 3044
rect 18890 3004 18930 3044
rect 18972 3004 19012 3044
rect 19054 3004 19094 3044
rect 19136 3004 19176 3044
rect 18808 1492 18848 1532
rect 18890 1492 18930 1532
rect 18972 1492 19012 1532
rect 19054 1492 19094 1532
rect 19136 1492 19176 1532
rect 20812 15268 20852 15308
rect 20620 7036 20660 7076
rect 20524 6952 20564 6992
rect 20048 6784 20088 6824
rect 20130 6784 20170 6824
rect 20212 6784 20252 6824
rect 20294 6784 20334 6824
rect 20376 6784 20416 6824
rect 20048 5272 20088 5312
rect 20130 5272 20170 5312
rect 20212 5272 20252 5312
rect 20294 5272 20334 5312
rect 20376 5272 20416 5312
rect 20048 3760 20088 3800
rect 20130 3760 20170 3800
rect 20212 3760 20252 3800
rect 20294 3760 20334 3800
rect 20376 3760 20416 3800
rect 20908 3256 20948 3296
rect 20812 3172 20852 3212
rect 20048 2248 20088 2288
rect 20130 2248 20170 2288
rect 20212 2248 20252 2288
rect 20294 2248 20334 2288
rect 20376 2248 20416 2288
rect 20048 736 20088 776
rect 20130 736 20170 776
rect 20212 736 20252 776
rect 20294 736 20334 776
rect 20376 736 20416 776
<< metal5 >>
rect 4919 41623 5305 41642
rect 4919 41600 4985 41623
rect 5071 41600 5153 41623
rect 5239 41600 5305 41623
rect 4919 41560 4928 41600
rect 4968 41560 4985 41600
rect 5071 41560 5092 41600
rect 5132 41560 5153 41600
rect 5239 41560 5256 41600
rect 5296 41560 5305 41600
rect 4919 41537 4985 41560
rect 5071 41537 5153 41560
rect 5239 41537 5305 41560
rect 4919 41518 5305 41537
rect 20039 41623 20425 41642
rect 20039 41600 20105 41623
rect 20191 41600 20273 41623
rect 20359 41600 20425 41623
rect 20039 41560 20048 41600
rect 20088 41560 20105 41600
rect 20191 41560 20212 41600
rect 20252 41560 20273 41600
rect 20359 41560 20376 41600
rect 20416 41560 20425 41600
rect 20039 41537 20105 41560
rect 20191 41537 20273 41560
rect 20359 41537 20425 41560
rect 20039 41518 20425 41537
rect 3679 40867 4065 40886
rect 3679 40844 3745 40867
rect 3831 40844 3913 40867
rect 3999 40844 4065 40867
rect 3679 40804 3688 40844
rect 3728 40804 3745 40844
rect 3831 40804 3852 40844
rect 3892 40804 3913 40844
rect 3999 40804 4016 40844
rect 4056 40804 4065 40844
rect 3679 40781 3745 40804
rect 3831 40781 3913 40804
rect 3999 40781 4065 40804
rect 3679 40762 4065 40781
rect 18799 40867 19185 40886
rect 18799 40844 18865 40867
rect 18951 40844 19033 40867
rect 19119 40844 19185 40867
rect 18799 40804 18808 40844
rect 18848 40804 18865 40844
rect 18951 40804 18972 40844
rect 19012 40804 19033 40844
rect 19119 40804 19136 40844
rect 19176 40804 19185 40844
rect 18799 40781 18865 40804
rect 18951 40781 19033 40804
rect 19119 40781 19185 40804
rect 18799 40762 19185 40781
rect 12122 40531 12246 40550
rect 12122 40445 12141 40531
rect 12227 40508 12246 40531
rect 12227 40468 18892 40508
rect 18932 40468 18941 40508
rect 12227 40445 12246 40468
rect 12122 40426 12246 40445
rect 4919 40111 5305 40130
rect 4919 40088 4985 40111
rect 5071 40088 5153 40111
rect 5239 40088 5305 40111
rect 4919 40048 4928 40088
rect 4968 40048 4985 40088
rect 5071 40048 5092 40088
rect 5132 40048 5153 40088
rect 5239 40048 5256 40088
rect 5296 40048 5305 40088
rect 4919 40025 4985 40048
rect 5071 40025 5153 40048
rect 5239 40025 5305 40048
rect 4919 40006 5305 40025
rect 20039 40111 20425 40130
rect 20039 40088 20105 40111
rect 20191 40088 20273 40111
rect 20359 40088 20425 40111
rect 20039 40048 20048 40088
rect 20088 40048 20105 40088
rect 20191 40048 20212 40088
rect 20252 40048 20273 40088
rect 20359 40048 20376 40088
rect 20416 40048 20425 40088
rect 20039 40025 20105 40048
rect 20191 40025 20273 40048
rect 20359 40025 20425 40048
rect 20039 40006 20425 40025
rect 17138 39859 17262 39878
rect 17138 39773 17157 39859
rect 17243 39773 17262 39859
rect 17138 39754 17262 39773
rect 3679 39355 4065 39374
rect 3679 39332 3745 39355
rect 3831 39332 3913 39355
rect 3999 39332 4065 39355
rect 3679 39292 3688 39332
rect 3728 39292 3745 39332
rect 3831 39292 3852 39332
rect 3892 39292 3913 39332
rect 3999 39292 4016 39332
rect 4056 39292 4065 39332
rect 3679 39269 3745 39292
rect 3831 39269 3913 39292
rect 3999 39269 4065 39292
rect 3679 39250 4065 39269
rect 18799 39355 19185 39374
rect 18799 39332 18865 39355
rect 18951 39332 19033 39355
rect 19119 39332 19185 39355
rect 18799 39292 18808 39332
rect 18848 39292 18865 39332
rect 18951 39292 18972 39332
rect 19012 39292 19033 39332
rect 19119 39292 19136 39332
rect 19176 39292 19185 39332
rect 18799 39269 18865 39292
rect 18951 39269 19033 39292
rect 19119 39269 19185 39292
rect 18799 39250 19185 39269
rect 15043 38704 15052 38744
rect 15092 38704 18220 38744
rect 18260 38704 18269 38744
rect 13699 38620 13708 38660
rect 13748 38620 18988 38660
rect 19028 38620 19037 38660
rect 4919 38599 5305 38618
rect 4919 38576 4985 38599
rect 5071 38576 5153 38599
rect 5239 38576 5305 38599
rect 4919 38536 4928 38576
rect 4968 38536 4985 38576
rect 5071 38536 5092 38576
rect 5132 38536 5153 38576
rect 5239 38536 5256 38576
rect 5296 38536 5305 38576
rect 4919 38513 4985 38536
rect 5071 38513 5153 38536
rect 5239 38513 5305 38536
rect 4919 38494 5305 38513
rect 20039 38599 20425 38618
rect 20039 38576 20105 38599
rect 20191 38576 20273 38599
rect 20359 38576 20425 38599
rect 20039 38536 20048 38576
rect 20088 38536 20105 38576
rect 20191 38536 20212 38576
rect 20252 38536 20273 38576
rect 20359 38536 20376 38576
rect 20416 38536 20425 38576
rect 20039 38513 20105 38536
rect 20191 38513 20273 38536
rect 20359 38513 20425 38536
rect 20039 38494 20425 38513
rect 12835 38368 12844 38408
rect 12884 38368 18700 38408
rect 18740 38368 19044 38408
rect 19004 38324 19044 38368
rect 19004 38284 20140 38324
rect 20180 38284 20189 38324
rect 3331 38200 3340 38240
rect 3380 38200 9580 38240
rect 9620 38200 9629 38240
rect 2563 38032 2572 38072
rect 2612 38032 2956 38072
rect 2996 38032 10252 38072
rect 10292 38032 10301 38072
rect 3679 37843 4065 37862
rect 3679 37820 3745 37843
rect 3831 37820 3913 37843
rect 3999 37820 4065 37843
rect 3679 37780 3688 37820
rect 3728 37780 3745 37820
rect 3831 37780 3852 37820
rect 3892 37780 3913 37820
rect 3999 37780 4016 37820
rect 4056 37780 4065 37820
rect 3679 37757 3745 37780
rect 3831 37757 3913 37780
rect 3999 37757 4065 37780
rect 3679 37738 4065 37757
rect 18799 37843 19185 37862
rect 18799 37820 18865 37843
rect 18951 37820 19033 37843
rect 19119 37820 19185 37843
rect 18799 37780 18808 37820
rect 18848 37780 18865 37820
rect 18951 37780 18972 37820
rect 19012 37780 19033 37820
rect 19119 37780 19136 37820
rect 19176 37780 19185 37820
rect 18799 37757 18865 37780
rect 18951 37757 19033 37780
rect 19119 37757 19185 37780
rect 18799 37738 19185 37757
rect 4919 37087 5305 37106
rect 4919 37064 4985 37087
rect 5071 37064 5153 37087
rect 5239 37064 5305 37087
rect 4919 37024 4928 37064
rect 4968 37024 4985 37064
rect 5071 37024 5092 37064
rect 5132 37024 5153 37064
rect 5239 37024 5256 37064
rect 5296 37024 5305 37064
rect 4919 37001 4985 37024
rect 5071 37001 5153 37024
rect 5239 37001 5305 37024
rect 4919 36982 5305 37001
rect 20039 37087 20425 37106
rect 20039 37064 20105 37087
rect 20191 37064 20273 37087
rect 20359 37064 20425 37087
rect 20039 37024 20048 37064
rect 20088 37024 20105 37064
rect 20191 37024 20212 37064
rect 20252 37024 20273 37064
rect 20359 37024 20376 37064
rect 20416 37024 20425 37064
rect 20039 37001 20105 37024
rect 20191 37001 20273 37024
rect 20359 37001 20425 37024
rect 20039 36982 20425 37001
rect 3679 36331 4065 36350
rect 3679 36308 3745 36331
rect 3831 36308 3913 36331
rect 3999 36308 4065 36331
rect 3679 36268 3688 36308
rect 3728 36268 3745 36308
rect 3831 36268 3852 36308
rect 3892 36268 3913 36308
rect 3999 36268 4016 36308
rect 4056 36268 4065 36308
rect 3679 36245 3745 36268
rect 3831 36245 3913 36268
rect 3999 36245 4065 36268
rect 3679 36226 4065 36245
rect 18799 36331 19185 36350
rect 18799 36308 18865 36331
rect 18951 36308 19033 36331
rect 19119 36308 19185 36331
rect 18799 36268 18808 36308
rect 18848 36268 18865 36308
rect 18951 36268 18972 36308
rect 19012 36268 19033 36308
rect 19119 36268 19136 36308
rect 19176 36268 19185 36308
rect 18799 36245 18865 36268
rect 18951 36245 19033 36268
rect 19119 36245 19185 36268
rect 18799 36226 19185 36245
rect 4919 35575 5305 35594
rect 4919 35552 4985 35575
rect 5071 35552 5153 35575
rect 5239 35552 5305 35575
rect 4919 35512 4928 35552
rect 4968 35512 4985 35552
rect 5071 35512 5092 35552
rect 5132 35512 5153 35552
rect 5239 35512 5256 35552
rect 5296 35512 5305 35552
rect 4919 35489 4985 35512
rect 5071 35489 5153 35512
rect 5239 35489 5305 35512
rect 4919 35470 5305 35489
rect 20039 35575 20425 35594
rect 20039 35552 20105 35575
rect 20191 35552 20273 35575
rect 20359 35552 20425 35575
rect 20039 35512 20048 35552
rect 20088 35512 20105 35552
rect 20191 35512 20212 35552
rect 20252 35512 20273 35552
rect 20359 35512 20376 35552
rect 20416 35512 20425 35552
rect 20039 35489 20105 35512
rect 20191 35489 20273 35512
rect 20359 35489 20425 35512
rect 20039 35470 20425 35489
rect 3679 34819 4065 34838
rect 3679 34796 3745 34819
rect 3831 34796 3913 34819
rect 3999 34796 4065 34819
rect 3679 34756 3688 34796
rect 3728 34756 3745 34796
rect 3831 34756 3852 34796
rect 3892 34756 3913 34796
rect 3999 34756 4016 34796
rect 4056 34756 4065 34796
rect 3679 34733 3745 34756
rect 3831 34733 3913 34756
rect 3999 34733 4065 34756
rect 3679 34714 4065 34733
rect 18799 34819 19185 34838
rect 18799 34796 18865 34819
rect 18951 34796 19033 34819
rect 19119 34796 19185 34819
rect 18799 34756 18808 34796
rect 18848 34756 18865 34796
rect 18951 34756 18972 34796
rect 19012 34756 19033 34796
rect 19119 34756 19136 34796
rect 19176 34756 19185 34796
rect 18799 34733 18865 34756
rect 18951 34733 19033 34756
rect 19119 34733 19185 34756
rect 18799 34714 19185 34733
rect 4919 34063 5305 34082
rect 4919 34040 4985 34063
rect 5071 34040 5153 34063
rect 5239 34040 5305 34063
rect 4919 34000 4928 34040
rect 4968 34000 4985 34040
rect 5071 34000 5092 34040
rect 5132 34000 5153 34040
rect 5239 34000 5256 34040
rect 5296 34000 5305 34040
rect 4919 33977 4985 34000
rect 5071 33977 5153 34000
rect 5239 33977 5305 34000
rect 4919 33958 5305 33977
rect 20039 34063 20425 34082
rect 20039 34040 20105 34063
rect 20191 34040 20273 34063
rect 20359 34040 20425 34063
rect 20039 34000 20048 34040
rect 20088 34000 20105 34040
rect 20191 34000 20212 34040
rect 20252 34000 20273 34040
rect 20359 34000 20376 34040
rect 20416 34000 20425 34040
rect 20039 33977 20105 34000
rect 20191 33977 20273 34000
rect 20359 33977 20425 34000
rect 20039 33958 20425 33977
rect 3679 33307 4065 33326
rect 3679 33284 3745 33307
rect 3831 33284 3913 33307
rect 3999 33284 4065 33307
rect 3679 33244 3688 33284
rect 3728 33244 3745 33284
rect 3831 33244 3852 33284
rect 3892 33244 3913 33284
rect 3999 33244 4016 33284
rect 4056 33244 4065 33284
rect 3679 33221 3745 33244
rect 3831 33221 3913 33244
rect 3999 33221 4065 33244
rect 3679 33202 4065 33221
rect 18799 33307 19185 33326
rect 18799 33284 18865 33307
rect 18951 33284 19033 33307
rect 19119 33284 19185 33307
rect 18799 33244 18808 33284
rect 18848 33244 18865 33284
rect 18951 33244 18972 33284
rect 19012 33244 19033 33284
rect 19119 33244 19136 33284
rect 19176 33244 19185 33284
rect 18799 33221 18865 33244
rect 18951 33221 19033 33244
rect 19119 33221 19185 33244
rect 18799 33202 19185 33221
rect 3715 32908 3724 32948
rect 3764 32908 9580 32948
rect 9620 32908 9629 32948
rect 4919 32551 5305 32570
rect 4919 32528 4985 32551
rect 5071 32528 5153 32551
rect 5239 32528 5305 32551
rect 4919 32488 4928 32528
rect 4968 32488 4985 32528
rect 5071 32488 5092 32528
rect 5132 32488 5153 32528
rect 5239 32488 5256 32528
rect 5296 32488 5305 32528
rect 4919 32465 4985 32488
rect 5071 32465 5153 32488
rect 5239 32465 5305 32488
rect 4919 32446 5305 32465
rect 20039 32551 20425 32570
rect 20039 32528 20105 32551
rect 20191 32528 20273 32551
rect 20359 32528 20425 32551
rect 20039 32488 20048 32528
rect 20088 32488 20105 32528
rect 20191 32488 20212 32528
rect 20252 32488 20273 32528
rect 20359 32488 20376 32528
rect 20416 32488 20425 32528
rect 20039 32465 20105 32488
rect 20191 32465 20273 32488
rect 20359 32465 20425 32488
rect 20039 32446 20425 32465
rect 3679 31795 4065 31814
rect 3679 31772 3745 31795
rect 3831 31772 3913 31795
rect 3999 31772 4065 31795
rect 3679 31732 3688 31772
rect 3728 31732 3745 31772
rect 3831 31732 3852 31772
rect 3892 31732 3913 31772
rect 3999 31732 4016 31772
rect 4056 31732 4065 31772
rect 3679 31709 3745 31732
rect 3831 31709 3913 31732
rect 3999 31709 4065 31732
rect 3679 31690 4065 31709
rect 18799 31795 19185 31814
rect 18799 31772 18865 31795
rect 18951 31772 19033 31795
rect 19119 31772 19185 31795
rect 18799 31732 18808 31772
rect 18848 31732 18865 31772
rect 18951 31732 18972 31772
rect 19012 31732 19033 31772
rect 19119 31732 19136 31772
rect 19176 31732 19185 31772
rect 18799 31709 18865 31732
rect 18951 31709 19033 31732
rect 19119 31709 19185 31732
rect 18799 31690 19185 31709
rect 4919 31039 5305 31058
rect 4919 31016 4985 31039
rect 5071 31016 5153 31039
rect 5239 31016 5305 31039
rect 4919 30976 4928 31016
rect 4968 30976 4985 31016
rect 5071 30976 5092 31016
rect 5132 30976 5153 31016
rect 5239 30976 5256 31016
rect 5296 30976 5305 31016
rect 4919 30953 4985 30976
rect 5071 30953 5153 30976
rect 5239 30953 5305 30976
rect 4919 30934 5305 30953
rect 20039 31039 20425 31058
rect 20039 31016 20105 31039
rect 20191 31016 20273 31039
rect 20359 31016 20425 31039
rect 20039 30976 20048 31016
rect 20088 30976 20105 31016
rect 20191 30976 20212 31016
rect 20252 30976 20273 31016
rect 20359 30976 20376 31016
rect 20416 30976 20425 31016
rect 20039 30953 20105 30976
rect 20191 30953 20273 30976
rect 20359 30953 20425 30976
rect 20039 30934 20425 30953
rect 3679 30283 4065 30302
rect 3679 30260 3745 30283
rect 3831 30260 3913 30283
rect 3999 30260 4065 30283
rect 3679 30220 3688 30260
rect 3728 30220 3745 30260
rect 3831 30220 3852 30260
rect 3892 30220 3913 30260
rect 3999 30220 4016 30260
rect 4056 30220 4065 30260
rect 3679 30197 3745 30220
rect 3831 30197 3913 30220
rect 3999 30197 4065 30220
rect 3679 30178 4065 30197
rect 18799 30283 19185 30302
rect 18799 30260 18865 30283
rect 18951 30260 19033 30283
rect 19119 30260 19185 30283
rect 18799 30220 18808 30260
rect 18848 30220 18865 30260
rect 18951 30220 18972 30260
rect 19012 30220 19033 30260
rect 19119 30220 19136 30260
rect 19176 30220 19185 30260
rect 18799 30197 18865 30220
rect 18951 30197 19033 30220
rect 19119 30197 19185 30220
rect 18799 30178 19185 30197
rect 4919 29527 5305 29546
rect 4919 29504 4985 29527
rect 5071 29504 5153 29527
rect 5239 29504 5305 29527
rect 4919 29464 4928 29504
rect 4968 29464 4985 29504
rect 5071 29464 5092 29504
rect 5132 29464 5153 29504
rect 5239 29464 5256 29504
rect 5296 29464 5305 29504
rect 4919 29441 4985 29464
rect 5071 29441 5153 29464
rect 5239 29441 5305 29464
rect 4919 29422 5305 29441
rect 20039 29527 20425 29546
rect 20039 29504 20105 29527
rect 20191 29504 20273 29527
rect 20359 29504 20425 29527
rect 20039 29464 20048 29504
rect 20088 29464 20105 29504
rect 20191 29464 20212 29504
rect 20252 29464 20273 29504
rect 20359 29464 20376 29504
rect 20416 29464 20425 29504
rect 20039 29441 20105 29464
rect 20191 29441 20273 29464
rect 20359 29441 20425 29464
rect 20039 29422 20425 29441
rect 3679 28771 4065 28790
rect 3679 28748 3745 28771
rect 3831 28748 3913 28771
rect 3999 28748 4065 28771
rect 3679 28708 3688 28748
rect 3728 28708 3745 28748
rect 3831 28708 3852 28748
rect 3892 28708 3913 28748
rect 3999 28708 4016 28748
rect 4056 28708 4065 28748
rect 3679 28685 3745 28708
rect 3831 28685 3913 28708
rect 3999 28685 4065 28708
rect 3679 28666 4065 28685
rect 18799 28771 19185 28790
rect 18799 28748 18865 28771
rect 18951 28748 19033 28771
rect 19119 28748 19185 28771
rect 18799 28708 18808 28748
rect 18848 28708 18865 28748
rect 18951 28708 18972 28748
rect 19012 28708 19033 28748
rect 19119 28708 19136 28748
rect 19176 28708 19185 28748
rect 18799 28685 18865 28708
rect 18951 28685 19033 28708
rect 19119 28685 19185 28708
rect 18799 28666 19185 28685
rect 4919 28015 5305 28034
rect 4919 27992 4985 28015
rect 5071 27992 5153 28015
rect 5239 27992 5305 28015
rect 4919 27952 4928 27992
rect 4968 27952 4985 27992
rect 5071 27952 5092 27992
rect 5132 27952 5153 27992
rect 5239 27952 5256 27992
rect 5296 27952 5305 27992
rect 4919 27929 4985 27952
rect 5071 27929 5153 27952
rect 5239 27929 5305 27952
rect 4919 27910 5305 27929
rect 20039 28015 20425 28034
rect 20039 27992 20105 28015
rect 20191 27992 20273 28015
rect 20359 27992 20425 28015
rect 20039 27952 20048 27992
rect 20088 27952 20105 27992
rect 20191 27952 20212 27992
rect 20252 27952 20273 27992
rect 20359 27952 20376 27992
rect 20416 27952 20425 27992
rect 20039 27929 20105 27952
rect 20191 27929 20273 27952
rect 20359 27929 20425 27952
rect 20039 27910 20425 27929
rect 3679 27259 4065 27278
rect 3679 27236 3745 27259
rect 3831 27236 3913 27259
rect 3999 27236 4065 27259
rect 3679 27196 3688 27236
rect 3728 27196 3745 27236
rect 3831 27196 3852 27236
rect 3892 27196 3913 27236
rect 3999 27196 4016 27236
rect 4056 27196 4065 27236
rect 3679 27173 3745 27196
rect 3831 27173 3913 27196
rect 3999 27173 4065 27196
rect 3679 27154 4065 27173
rect 18799 27259 19185 27278
rect 18799 27236 18865 27259
rect 18951 27236 19033 27259
rect 19119 27236 19185 27259
rect 18799 27196 18808 27236
rect 18848 27196 18865 27236
rect 18951 27196 18972 27236
rect 19012 27196 19033 27236
rect 19119 27196 19136 27236
rect 19176 27196 19185 27236
rect 18799 27173 18865 27196
rect 18951 27173 19033 27196
rect 19119 27173 19185 27196
rect 18799 27154 19185 27173
rect 4919 26503 5305 26522
rect 4919 26480 4985 26503
rect 5071 26480 5153 26503
rect 5239 26480 5305 26503
rect 4919 26440 4928 26480
rect 4968 26440 4985 26480
rect 5071 26440 5092 26480
rect 5132 26440 5153 26480
rect 5239 26440 5256 26480
rect 5296 26440 5305 26480
rect 4919 26417 4985 26440
rect 5071 26417 5153 26440
rect 5239 26417 5305 26440
rect 4919 26398 5305 26417
rect 20039 26503 20425 26522
rect 20039 26480 20105 26503
rect 20191 26480 20273 26503
rect 20359 26480 20425 26503
rect 20039 26440 20048 26480
rect 20088 26440 20105 26480
rect 20191 26440 20212 26480
rect 20252 26440 20273 26480
rect 20359 26440 20376 26480
rect 20416 26440 20425 26480
rect 20039 26417 20105 26440
rect 20191 26417 20273 26440
rect 20359 26417 20425 26440
rect 20039 26398 20425 26417
rect 3679 25747 4065 25766
rect 3679 25724 3745 25747
rect 3831 25724 3913 25747
rect 3999 25724 4065 25747
rect 3679 25684 3688 25724
rect 3728 25684 3745 25724
rect 3831 25684 3852 25724
rect 3892 25684 3913 25724
rect 3999 25684 4016 25724
rect 4056 25684 4065 25724
rect 3679 25661 3745 25684
rect 3831 25661 3913 25684
rect 3999 25661 4065 25684
rect 3679 25642 4065 25661
rect 18799 25747 19185 25766
rect 18799 25724 18865 25747
rect 18951 25724 19033 25747
rect 19119 25724 19185 25747
rect 18799 25684 18808 25724
rect 18848 25684 18865 25724
rect 18951 25684 18972 25724
rect 19012 25684 19033 25724
rect 19119 25684 19136 25724
rect 19176 25684 19185 25724
rect 18799 25661 18865 25684
rect 18951 25661 19033 25684
rect 19119 25661 19185 25684
rect 18799 25642 19185 25661
rect 4919 24991 5305 25010
rect 4919 24968 4985 24991
rect 5071 24968 5153 24991
rect 5239 24968 5305 24991
rect 4919 24928 4928 24968
rect 4968 24928 4985 24968
rect 5071 24928 5092 24968
rect 5132 24928 5153 24968
rect 5239 24928 5256 24968
rect 5296 24928 5305 24968
rect 4919 24905 4985 24928
rect 5071 24905 5153 24928
rect 5239 24905 5305 24928
rect 4919 24886 5305 24905
rect 20039 24991 20425 25010
rect 20039 24968 20105 24991
rect 20191 24968 20273 24991
rect 20359 24968 20425 24991
rect 20039 24928 20048 24968
rect 20088 24928 20105 24968
rect 20191 24928 20212 24968
rect 20252 24928 20273 24968
rect 20359 24928 20376 24968
rect 20416 24928 20425 24968
rect 20039 24905 20105 24928
rect 20191 24905 20273 24928
rect 20359 24905 20425 24928
rect 20039 24886 20425 24905
rect 3679 24235 4065 24254
rect 3679 24212 3745 24235
rect 3831 24212 3913 24235
rect 3999 24212 4065 24235
rect 3679 24172 3688 24212
rect 3728 24172 3745 24212
rect 3831 24172 3852 24212
rect 3892 24172 3913 24212
rect 3999 24172 4016 24212
rect 4056 24172 4065 24212
rect 3679 24149 3745 24172
rect 3831 24149 3913 24172
rect 3999 24149 4065 24172
rect 3679 24130 4065 24149
rect 18799 24235 19185 24254
rect 18799 24212 18865 24235
rect 18951 24212 19033 24235
rect 19119 24212 19185 24235
rect 18799 24172 18808 24212
rect 18848 24172 18865 24212
rect 18951 24172 18972 24212
rect 19012 24172 19033 24212
rect 19119 24172 19136 24212
rect 19176 24172 19185 24212
rect 18799 24149 18865 24172
rect 18951 24149 19033 24172
rect 19119 24149 19185 24172
rect 18799 24130 19185 24149
rect 4919 23479 5305 23498
rect 4919 23456 4985 23479
rect 5071 23456 5153 23479
rect 5239 23456 5305 23479
rect 4919 23416 4928 23456
rect 4968 23416 4985 23456
rect 5071 23416 5092 23456
rect 5132 23416 5153 23456
rect 5239 23416 5256 23456
rect 5296 23416 5305 23456
rect 4919 23393 4985 23416
rect 5071 23393 5153 23416
rect 5239 23393 5305 23416
rect 4919 23374 5305 23393
rect 20039 23479 20425 23498
rect 20039 23456 20105 23479
rect 20191 23456 20273 23479
rect 20359 23456 20425 23479
rect 20039 23416 20048 23456
rect 20088 23416 20105 23456
rect 20191 23416 20212 23456
rect 20252 23416 20273 23456
rect 20359 23416 20376 23456
rect 20416 23416 20425 23456
rect 20039 23393 20105 23416
rect 20191 23393 20273 23416
rect 20359 23393 20425 23416
rect 20039 23374 20425 23393
rect 7075 22996 7084 23036
rect 7124 22996 19276 23036
rect 19316 22996 19325 23036
rect 3679 22723 4065 22742
rect 3679 22700 3745 22723
rect 3831 22700 3913 22723
rect 3999 22700 4065 22723
rect 3679 22660 3688 22700
rect 3728 22660 3745 22700
rect 3831 22660 3852 22700
rect 3892 22660 3913 22700
rect 3999 22660 4016 22700
rect 4056 22660 4065 22700
rect 3679 22637 3745 22660
rect 3831 22637 3913 22660
rect 3999 22637 4065 22660
rect 3679 22618 4065 22637
rect 18799 22723 19185 22742
rect 18799 22700 18865 22723
rect 18951 22700 19033 22723
rect 19119 22700 19185 22723
rect 18799 22660 18808 22700
rect 18848 22660 18865 22700
rect 18951 22660 18972 22700
rect 19012 22660 19033 22700
rect 19119 22660 19136 22700
rect 19176 22660 19185 22700
rect 18799 22637 18865 22660
rect 18951 22637 19033 22660
rect 19119 22637 19185 22660
rect 18799 22618 19185 22637
rect 4919 21967 5305 21986
rect 4919 21944 4985 21967
rect 5071 21944 5153 21967
rect 5239 21944 5305 21967
rect 4919 21904 4928 21944
rect 4968 21904 4985 21944
rect 5071 21904 5092 21944
rect 5132 21904 5153 21944
rect 5239 21904 5256 21944
rect 5296 21904 5305 21944
rect 4919 21881 4985 21904
rect 5071 21881 5153 21904
rect 5239 21881 5305 21904
rect 4919 21862 5305 21881
rect 20039 21967 20425 21986
rect 20039 21944 20105 21967
rect 20191 21944 20273 21967
rect 20359 21944 20425 21967
rect 20039 21904 20048 21944
rect 20088 21904 20105 21944
rect 20191 21904 20212 21944
rect 20252 21904 20273 21944
rect 20359 21904 20376 21944
rect 20416 21904 20425 21944
rect 20039 21881 20105 21904
rect 20191 21881 20273 21904
rect 20359 21881 20425 21904
rect 20039 21862 20425 21881
rect 3679 21211 4065 21230
rect 3679 21188 3745 21211
rect 3831 21188 3913 21211
rect 3999 21188 4065 21211
rect 3679 21148 3688 21188
rect 3728 21148 3745 21188
rect 3831 21148 3852 21188
rect 3892 21148 3913 21188
rect 3999 21148 4016 21188
rect 4056 21148 4065 21188
rect 3679 21125 3745 21148
rect 3831 21125 3913 21148
rect 3999 21125 4065 21148
rect 3679 21106 4065 21125
rect 18799 21211 19185 21230
rect 18799 21188 18865 21211
rect 18951 21188 19033 21211
rect 19119 21188 19185 21211
rect 18799 21148 18808 21188
rect 18848 21148 18865 21188
rect 18951 21148 18972 21188
rect 19012 21148 19033 21188
rect 19119 21148 19136 21188
rect 19176 21148 19185 21188
rect 18799 21125 18865 21148
rect 18951 21125 19033 21148
rect 19119 21125 19185 21148
rect 18799 21106 19185 21125
rect 4919 20455 5305 20474
rect 4919 20432 4985 20455
rect 5071 20432 5153 20455
rect 5239 20432 5305 20455
rect 4919 20392 4928 20432
rect 4968 20392 4985 20432
rect 5071 20392 5092 20432
rect 5132 20392 5153 20432
rect 5239 20392 5256 20432
rect 5296 20392 5305 20432
rect 4919 20369 4985 20392
rect 5071 20369 5153 20392
rect 5239 20369 5305 20392
rect 4919 20350 5305 20369
rect 20039 20455 20425 20474
rect 20039 20432 20105 20455
rect 20191 20432 20273 20455
rect 20359 20432 20425 20455
rect 20039 20392 20048 20432
rect 20088 20392 20105 20432
rect 20191 20392 20212 20432
rect 20252 20392 20273 20432
rect 20359 20392 20376 20432
rect 20416 20392 20425 20432
rect 20039 20369 20105 20392
rect 20191 20369 20273 20392
rect 20359 20369 20425 20392
rect 20039 20350 20425 20369
rect 451 19972 460 20012
rect 500 19972 748 20012
rect 788 19972 797 20012
rect 3679 19699 4065 19718
rect 3679 19676 3745 19699
rect 3831 19676 3913 19699
rect 3999 19676 4065 19699
rect 3679 19636 3688 19676
rect 3728 19636 3745 19676
rect 3831 19636 3852 19676
rect 3892 19636 3913 19676
rect 3999 19636 4016 19676
rect 4056 19636 4065 19676
rect 3679 19613 3745 19636
rect 3831 19613 3913 19636
rect 3999 19613 4065 19636
rect 3679 19594 4065 19613
rect 18799 19699 19185 19718
rect 18799 19676 18865 19699
rect 18951 19676 19033 19699
rect 19119 19676 19185 19699
rect 18799 19636 18808 19676
rect 18848 19636 18865 19676
rect 18951 19636 18972 19676
rect 19012 19636 19033 19676
rect 19119 19636 19136 19676
rect 19176 19636 19185 19676
rect 18799 19613 18865 19636
rect 18951 19613 19033 19636
rect 19119 19613 19185 19636
rect 18799 19594 19185 19613
rect 4675 19468 4684 19508
rect 4724 19468 16972 19508
rect 17012 19468 17021 19508
rect 1219 19048 1228 19088
rect 1268 19048 16492 19088
rect 16532 19048 16541 19088
rect 4919 18943 5305 18962
rect 4919 18920 4985 18943
rect 5071 18920 5153 18943
rect 5239 18920 5305 18943
rect 4919 18880 4928 18920
rect 4968 18880 4985 18920
rect 5071 18880 5092 18920
rect 5132 18880 5153 18920
rect 5239 18880 5256 18920
rect 5296 18880 5305 18920
rect 4919 18857 4985 18880
rect 5071 18857 5153 18880
rect 5239 18857 5305 18880
rect 4919 18838 5305 18857
rect 20039 18943 20425 18962
rect 20039 18920 20105 18943
rect 20191 18920 20273 18943
rect 20359 18920 20425 18943
rect 20039 18880 20048 18920
rect 20088 18880 20105 18920
rect 20191 18880 20212 18920
rect 20252 18880 20273 18920
rect 20359 18880 20376 18920
rect 20416 18880 20425 18920
rect 20039 18857 20105 18880
rect 20191 18857 20273 18880
rect 20359 18857 20425 18880
rect 20039 18838 20425 18857
rect 3679 18187 4065 18206
rect 3679 18164 3745 18187
rect 3831 18164 3913 18187
rect 3999 18164 4065 18187
rect 3679 18124 3688 18164
rect 3728 18124 3745 18164
rect 3831 18124 3852 18164
rect 3892 18124 3913 18164
rect 3999 18124 4016 18164
rect 4056 18124 4065 18164
rect 3679 18101 3745 18124
rect 3831 18101 3913 18124
rect 3999 18101 4065 18124
rect 3679 18082 4065 18101
rect 18799 18187 19185 18206
rect 18799 18164 18865 18187
rect 18951 18164 19033 18187
rect 19119 18164 19185 18187
rect 18799 18124 18808 18164
rect 18848 18124 18865 18164
rect 18951 18124 18972 18164
rect 19012 18124 19033 18164
rect 19119 18124 19136 18164
rect 19176 18124 19185 18164
rect 18799 18101 18865 18124
rect 18951 18101 19033 18124
rect 19119 18101 19185 18124
rect 18799 18082 19185 18101
rect 4919 17431 5305 17450
rect 4919 17408 4985 17431
rect 5071 17408 5153 17431
rect 5239 17408 5305 17431
rect 4919 17368 4928 17408
rect 4968 17368 4985 17408
rect 5071 17368 5092 17408
rect 5132 17368 5153 17408
rect 5239 17368 5256 17408
rect 5296 17368 5305 17408
rect 4919 17345 4985 17368
rect 5071 17345 5153 17368
rect 5239 17345 5305 17368
rect 4919 17326 5305 17345
rect 20039 17431 20425 17450
rect 20039 17408 20105 17431
rect 20191 17408 20273 17431
rect 20359 17408 20425 17431
rect 20039 17368 20048 17408
rect 20088 17368 20105 17408
rect 20191 17368 20212 17408
rect 20252 17368 20273 17408
rect 20359 17368 20376 17408
rect 20416 17368 20425 17408
rect 20039 17345 20105 17368
rect 20191 17345 20273 17368
rect 20359 17345 20425 17368
rect 20039 17326 20425 17345
rect 3679 16675 4065 16694
rect 3679 16652 3745 16675
rect 3831 16652 3913 16675
rect 3999 16652 4065 16675
rect 18799 16675 19185 16694
rect 18799 16652 18865 16675
rect 18951 16652 19033 16675
rect 19119 16652 19185 16675
rect 3679 16612 3688 16652
rect 3728 16612 3745 16652
rect 3831 16612 3852 16652
rect 3892 16612 3913 16652
rect 3999 16612 4016 16652
rect 4056 16612 4065 16652
rect 14755 16612 14764 16652
rect 14804 16612 14956 16652
rect 14996 16612 15005 16652
rect 18799 16612 18808 16652
rect 18848 16612 18865 16652
rect 18951 16612 18972 16652
rect 19012 16612 19033 16652
rect 19119 16612 19136 16652
rect 19176 16612 19185 16652
rect 3679 16589 3745 16612
rect 3831 16589 3913 16612
rect 3999 16589 4065 16612
rect 3679 16570 4065 16589
rect 18799 16589 18865 16612
rect 18951 16589 19033 16612
rect 19119 16589 19185 16612
rect 18799 16570 19185 16589
rect 2500 16360 17068 16400
rect 17108 16360 17117 16400
rect 2500 16316 2540 16360
rect 547 16276 556 16316
rect 596 16276 2540 16316
rect 451 16108 460 16148
rect 500 16108 5068 16148
rect 5108 16108 5117 16148
rect 4919 15919 5305 15938
rect 4919 15896 4985 15919
rect 5071 15896 5153 15919
rect 5239 15896 5305 15919
rect 4919 15856 4928 15896
rect 4968 15856 4985 15896
rect 5071 15856 5092 15896
rect 5132 15856 5153 15896
rect 5239 15856 5256 15896
rect 5296 15856 5305 15896
rect 4919 15833 4985 15856
rect 5071 15833 5153 15856
rect 5239 15833 5305 15856
rect 4919 15814 5305 15833
rect 20039 15919 20425 15938
rect 20039 15896 20105 15919
rect 20191 15896 20273 15919
rect 20359 15896 20425 15919
rect 20039 15856 20048 15896
rect 20088 15856 20105 15896
rect 20191 15856 20212 15896
rect 20252 15856 20273 15896
rect 20359 15856 20376 15896
rect 20416 15856 20425 15896
rect 20039 15833 20105 15856
rect 20191 15833 20273 15856
rect 20359 15833 20425 15856
rect 20039 15814 20425 15833
rect 11011 15436 11020 15476
rect 11060 15436 11692 15476
rect 11732 15436 12556 15476
rect 12596 15436 12605 15476
rect 4771 15268 4780 15308
rect 4820 15268 20812 15308
rect 20852 15268 20861 15308
rect 3679 15163 4065 15182
rect 3679 15140 3745 15163
rect 3831 15140 3913 15163
rect 3999 15140 4065 15163
rect 3679 15100 3688 15140
rect 3728 15100 3745 15140
rect 3831 15100 3852 15140
rect 3892 15100 3913 15140
rect 3999 15100 4016 15140
rect 4056 15100 4065 15140
rect 3679 15077 3745 15100
rect 3831 15077 3913 15100
rect 3999 15077 4065 15100
rect 3679 15058 4065 15077
rect 18799 15163 19185 15182
rect 18799 15140 18865 15163
rect 18951 15140 19033 15163
rect 19119 15140 19185 15163
rect 18799 15100 18808 15140
rect 18848 15100 18865 15140
rect 18951 15100 18972 15140
rect 19012 15100 19033 15140
rect 19119 15100 19136 15140
rect 19176 15100 19185 15140
rect 18799 15077 18865 15100
rect 18951 15077 19033 15100
rect 19119 15077 19185 15100
rect 18799 15058 19185 15077
rect 4675 14512 4684 14552
rect 4724 14512 14956 14552
rect 14996 14512 15005 14552
rect 4919 14407 5305 14426
rect 4919 14384 4985 14407
rect 5071 14384 5153 14407
rect 5239 14384 5305 14407
rect 4919 14344 4928 14384
rect 4968 14344 4985 14384
rect 5071 14344 5092 14384
rect 5132 14344 5153 14384
rect 5239 14344 5256 14384
rect 5296 14344 5305 14384
rect 4919 14321 4985 14344
rect 5071 14321 5153 14344
rect 5239 14321 5305 14344
rect 4919 14302 5305 14321
rect 20039 14407 20425 14426
rect 20039 14384 20105 14407
rect 20191 14384 20273 14407
rect 20359 14384 20425 14407
rect 20039 14344 20048 14384
rect 20088 14344 20105 14384
rect 20191 14344 20212 14384
rect 20252 14344 20273 14384
rect 20359 14344 20376 14384
rect 20416 14344 20425 14384
rect 20039 14321 20105 14344
rect 20191 14321 20273 14344
rect 20359 14321 20425 14344
rect 20039 14302 20425 14321
rect 3679 13651 4065 13670
rect 3679 13628 3745 13651
rect 3831 13628 3913 13651
rect 3999 13628 4065 13651
rect 3679 13588 3688 13628
rect 3728 13588 3745 13628
rect 3831 13588 3852 13628
rect 3892 13588 3913 13628
rect 3999 13588 4016 13628
rect 4056 13588 4065 13628
rect 3679 13565 3745 13588
rect 3831 13565 3913 13588
rect 3999 13565 4065 13588
rect 3679 13546 4065 13565
rect 18799 13651 19185 13670
rect 18799 13628 18865 13651
rect 18951 13628 19033 13651
rect 19119 13628 19185 13651
rect 18799 13588 18808 13628
rect 18848 13588 18865 13628
rect 18951 13588 18972 13628
rect 19012 13588 19033 13628
rect 19119 13588 19136 13628
rect 19176 13588 19185 13628
rect 18799 13565 18865 13588
rect 18951 13565 19033 13588
rect 19119 13565 19185 13588
rect 18799 13546 19185 13565
rect 4919 12895 5305 12914
rect 4919 12872 4985 12895
rect 5071 12872 5153 12895
rect 5239 12872 5305 12895
rect 4919 12832 4928 12872
rect 4968 12832 4985 12872
rect 5071 12832 5092 12872
rect 5132 12832 5153 12872
rect 5239 12832 5256 12872
rect 5296 12832 5305 12872
rect 4919 12809 4985 12832
rect 5071 12809 5153 12832
rect 5239 12809 5305 12832
rect 4919 12790 5305 12809
rect 20039 12895 20425 12914
rect 20039 12872 20105 12895
rect 20191 12872 20273 12895
rect 20359 12872 20425 12895
rect 20039 12832 20048 12872
rect 20088 12832 20105 12872
rect 20191 12832 20212 12872
rect 20252 12832 20273 12872
rect 20359 12832 20376 12872
rect 20416 12832 20425 12872
rect 20039 12809 20105 12832
rect 20191 12809 20273 12832
rect 20359 12809 20425 12832
rect 20039 12790 20425 12809
rect 13507 12580 13516 12620
rect 13556 12580 17356 12620
rect 17396 12580 17405 12620
rect 1219 12328 1228 12368
rect 1268 12328 17740 12368
rect 17780 12328 17789 12368
rect 3679 12139 4065 12158
rect 3679 12116 3745 12139
rect 3831 12116 3913 12139
rect 3999 12116 4065 12139
rect 3679 12076 3688 12116
rect 3728 12076 3745 12116
rect 3831 12076 3852 12116
rect 3892 12076 3913 12116
rect 3999 12076 4016 12116
rect 4056 12076 4065 12116
rect 3679 12053 3745 12076
rect 3831 12053 3913 12076
rect 3999 12053 4065 12076
rect 3679 12034 4065 12053
rect 18799 12139 19185 12158
rect 18799 12116 18865 12139
rect 18951 12116 19033 12139
rect 19119 12116 19185 12139
rect 18799 12076 18808 12116
rect 18848 12076 18865 12116
rect 18951 12076 18972 12116
rect 19012 12076 19033 12116
rect 19119 12076 19136 12116
rect 19176 12076 19185 12116
rect 18799 12053 18865 12076
rect 18951 12053 19033 12076
rect 19119 12053 19185 12076
rect 18799 12034 19185 12053
rect 5731 11740 5740 11780
rect 5780 11740 6220 11780
rect 6260 11740 6269 11780
rect 4919 11383 5305 11402
rect 4919 11360 4985 11383
rect 5071 11360 5153 11383
rect 5239 11360 5305 11383
rect 4919 11320 4928 11360
rect 4968 11320 4985 11360
rect 5071 11320 5092 11360
rect 5132 11320 5153 11360
rect 5239 11320 5256 11360
rect 5296 11320 5305 11360
rect 4919 11297 4985 11320
rect 5071 11297 5153 11320
rect 5239 11297 5305 11320
rect 4919 11278 5305 11297
rect 20039 11383 20425 11402
rect 20039 11360 20105 11383
rect 20191 11360 20273 11383
rect 20359 11360 20425 11383
rect 20039 11320 20048 11360
rect 20088 11320 20105 11360
rect 20191 11320 20212 11360
rect 20252 11320 20273 11360
rect 20359 11320 20376 11360
rect 20416 11320 20425 11360
rect 20039 11297 20105 11320
rect 20191 11297 20273 11320
rect 20359 11297 20425 11320
rect 20039 11278 20425 11297
rect 3679 10627 4065 10646
rect 3679 10604 3745 10627
rect 3831 10604 3913 10627
rect 3999 10604 4065 10627
rect 3679 10564 3688 10604
rect 3728 10564 3745 10604
rect 3831 10564 3852 10604
rect 3892 10564 3913 10604
rect 3999 10564 4016 10604
rect 4056 10564 4065 10604
rect 3679 10541 3745 10564
rect 3831 10541 3913 10564
rect 3999 10541 4065 10564
rect 3679 10522 4065 10541
rect 18799 10627 19185 10646
rect 18799 10604 18865 10627
rect 18951 10604 19033 10627
rect 19119 10604 19185 10627
rect 18799 10564 18808 10604
rect 18848 10564 18865 10604
rect 18951 10564 18972 10604
rect 19012 10564 19033 10604
rect 19119 10564 19136 10604
rect 19176 10564 19185 10604
rect 18799 10541 18865 10564
rect 18951 10541 19033 10564
rect 19119 10541 19185 10564
rect 18799 10522 19185 10541
rect 10147 10480 10156 10520
rect 10196 10480 10444 10520
rect 10484 10480 10493 10520
rect 4099 10144 4108 10184
rect 4148 10144 4588 10184
rect 4628 10144 16396 10184
rect 16436 10144 16445 10184
rect 4919 9871 5305 9890
rect 4919 9848 4985 9871
rect 5071 9848 5153 9871
rect 5239 9848 5305 9871
rect 4919 9808 4928 9848
rect 4968 9808 4985 9848
rect 5071 9808 5092 9848
rect 5132 9808 5153 9848
rect 5239 9808 5256 9848
rect 5296 9808 5305 9848
rect 4919 9785 4985 9808
rect 5071 9785 5153 9808
rect 5239 9785 5305 9808
rect 4919 9766 5305 9785
rect 20039 9871 20425 9890
rect 20039 9848 20105 9871
rect 20191 9848 20273 9871
rect 20359 9848 20425 9871
rect 20039 9808 20048 9848
rect 20088 9808 20105 9848
rect 20191 9808 20212 9848
rect 20252 9808 20273 9848
rect 20359 9808 20376 9848
rect 20416 9808 20425 9848
rect 20039 9785 20105 9808
rect 20191 9785 20273 9808
rect 20359 9785 20425 9808
rect 20039 9766 20425 9785
rect 3619 9388 3628 9428
rect 3668 9388 4300 9428
rect 4340 9388 7564 9428
rect 7604 9388 7613 9428
rect 8803 9304 8812 9344
rect 8852 9304 10924 9344
rect 10964 9304 10973 9344
rect 3679 9115 4065 9134
rect 3679 9092 3745 9115
rect 3831 9092 3913 9115
rect 3999 9092 4065 9115
rect 3679 9052 3688 9092
rect 3728 9052 3745 9092
rect 3831 9052 3852 9092
rect 3892 9052 3913 9092
rect 3999 9052 4016 9092
rect 4056 9052 4065 9092
rect 3679 9029 3745 9052
rect 3831 9029 3913 9052
rect 3999 9029 4065 9052
rect 3679 9010 4065 9029
rect 18799 9115 19185 9134
rect 18799 9092 18865 9115
rect 18951 9092 19033 9115
rect 19119 9092 19185 9115
rect 18799 9052 18808 9092
rect 18848 9052 18865 9092
rect 18951 9052 18972 9092
rect 19012 9052 19033 9092
rect 19119 9052 19136 9092
rect 19176 9052 19185 9092
rect 18799 9029 18865 9052
rect 18951 9029 19033 9052
rect 19119 9029 19185 9052
rect 18799 9010 19185 9029
rect 4919 8359 5305 8378
rect 4919 8336 4985 8359
rect 5071 8336 5153 8359
rect 5239 8336 5305 8359
rect 4919 8296 4928 8336
rect 4968 8296 4985 8336
rect 5071 8296 5092 8336
rect 5132 8296 5153 8336
rect 5239 8296 5256 8336
rect 5296 8296 5305 8336
rect 4919 8273 4985 8296
rect 5071 8273 5153 8296
rect 5239 8273 5305 8296
rect 4919 8254 5305 8273
rect 20039 8359 20425 8378
rect 20039 8336 20105 8359
rect 20191 8336 20273 8359
rect 20359 8336 20425 8359
rect 20039 8296 20048 8336
rect 20088 8296 20105 8336
rect 20191 8296 20212 8336
rect 20252 8296 20273 8336
rect 20359 8296 20376 8336
rect 20416 8296 20425 8336
rect 20039 8273 20105 8296
rect 20191 8273 20273 8296
rect 20359 8273 20425 8296
rect 20039 8254 20425 8273
rect 163 7708 172 7748
rect 212 7708 19084 7748
rect 19124 7708 19133 7748
rect 3679 7603 4065 7622
rect 3679 7580 3745 7603
rect 3831 7580 3913 7603
rect 3999 7580 4065 7603
rect 3679 7540 3688 7580
rect 3728 7540 3745 7580
rect 3831 7540 3852 7580
rect 3892 7540 3913 7580
rect 3999 7540 4016 7580
rect 4056 7540 4065 7580
rect 3679 7517 3745 7540
rect 3831 7517 3913 7540
rect 3999 7517 4065 7540
rect 3679 7498 4065 7517
rect 18799 7603 19185 7622
rect 18799 7580 18865 7603
rect 18951 7580 19033 7603
rect 19119 7580 19185 7603
rect 18799 7540 18808 7580
rect 18848 7540 18865 7580
rect 18951 7540 18972 7580
rect 19012 7540 19033 7580
rect 19119 7540 19136 7580
rect 19176 7540 19185 7580
rect 18799 7517 18865 7540
rect 18951 7517 19033 7540
rect 19119 7517 19185 7540
rect 18799 7498 19185 7517
rect 19459 7036 19468 7076
rect 19508 7036 20620 7076
rect 20660 7036 20669 7076
rect 931 6952 940 6992
rect 980 6952 13420 6992
rect 13460 6952 13469 6992
rect 19267 6952 19276 6992
rect 19316 6952 20524 6992
rect 20564 6952 20573 6992
rect 4919 6847 5305 6866
rect 4919 6824 4985 6847
rect 5071 6824 5153 6847
rect 5239 6824 5305 6847
rect 4919 6784 4928 6824
rect 4968 6784 4985 6824
rect 5071 6784 5092 6824
rect 5132 6784 5153 6824
rect 5239 6784 5256 6824
rect 5296 6784 5305 6824
rect 4919 6761 4985 6784
rect 5071 6761 5153 6784
rect 5239 6761 5305 6784
rect 4919 6742 5305 6761
rect 20039 6847 20425 6866
rect 20039 6824 20105 6847
rect 20191 6824 20273 6847
rect 20359 6824 20425 6847
rect 20039 6784 20048 6824
rect 20088 6784 20105 6824
rect 20191 6784 20212 6824
rect 20252 6784 20273 6824
rect 20359 6784 20376 6824
rect 20416 6784 20425 6824
rect 20039 6761 20105 6784
rect 20191 6761 20273 6784
rect 20359 6761 20425 6784
rect 20039 6742 20425 6761
rect 5635 6448 5644 6488
rect 5684 6448 9868 6488
rect 9908 6448 9917 6488
rect 5443 6112 5452 6152
rect 5492 6112 8908 6152
rect 8948 6112 8957 6152
rect 3679 6091 4065 6110
rect 3679 6068 3745 6091
rect 3831 6068 3913 6091
rect 3999 6068 4065 6091
rect 3679 6028 3688 6068
rect 3728 6028 3745 6068
rect 3831 6028 3852 6068
rect 3892 6028 3913 6068
rect 3999 6028 4016 6068
rect 4056 6028 4065 6068
rect 3679 6005 3745 6028
rect 3831 6005 3913 6028
rect 3999 6005 4065 6028
rect 3679 5986 4065 6005
rect 18799 6091 19185 6110
rect 18799 6068 18865 6091
rect 18951 6068 19033 6091
rect 19119 6068 19185 6091
rect 18799 6028 18808 6068
rect 18848 6028 18865 6068
rect 18951 6028 18972 6068
rect 19012 6028 19033 6068
rect 19119 6028 19136 6068
rect 19176 6028 19185 6068
rect 18799 6005 18865 6028
rect 18951 6005 19033 6028
rect 19119 6005 19185 6028
rect 18799 5986 19185 6005
rect 5347 5944 5356 5984
rect 5396 5944 9772 5984
rect 9812 5944 9821 5984
rect 12122 5839 12246 5858
rect 12122 5753 12141 5839
rect 12227 5816 12246 5839
rect 12227 5776 15628 5816
rect 15668 5776 15677 5816
rect 12227 5753 12246 5776
rect 12122 5734 12246 5753
rect 4919 5335 5305 5354
rect 4919 5312 4985 5335
rect 5071 5312 5153 5335
rect 5239 5312 5305 5335
rect 4919 5272 4928 5312
rect 4968 5272 4985 5312
rect 5071 5272 5092 5312
rect 5132 5272 5153 5312
rect 5239 5272 5256 5312
rect 5296 5272 5305 5312
rect 4919 5249 4985 5272
rect 5071 5249 5153 5272
rect 5239 5249 5305 5272
rect 4919 5230 5305 5249
rect 20039 5335 20425 5354
rect 20039 5312 20105 5335
rect 20191 5312 20273 5335
rect 20359 5312 20425 5335
rect 20039 5272 20048 5312
rect 20088 5272 20105 5312
rect 20191 5272 20212 5312
rect 20252 5272 20273 5312
rect 20359 5272 20376 5312
rect 20416 5272 20425 5312
rect 20039 5249 20105 5272
rect 20191 5249 20273 5272
rect 20359 5249 20425 5272
rect 20039 5230 20425 5249
rect 1219 4768 1228 4808
rect 1268 4768 13996 4808
rect 14036 4768 14045 4808
rect 3679 4579 4065 4598
rect 3679 4556 3745 4579
rect 3831 4556 3913 4579
rect 3999 4556 4065 4579
rect 3679 4516 3688 4556
rect 3728 4516 3745 4556
rect 3831 4516 3852 4556
rect 3892 4516 3913 4556
rect 3999 4516 4016 4556
rect 4056 4516 4065 4556
rect 3679 4493 3745 4516
rect 3831 4493 3913 4516
rect 3999 4493 4065 4516
rect 3679 4474 4065 4493
rect 18799 4579 19185 4598
rect 18799 4556 18865 4579
rect 18951 4556 19033 4579
rect 19119 4556 19185 4579
rect 18799 4516 18808 4556
rect 18848 4516 18865 4556
rect 18951 4516 18972 4556
rect 19012 4516 19033 4556
rect 19119 4516 19136 4556
rect 19176 4516 19185 4556
rect 18799 4493 18865 4516
rect 18951 4493 19033 4516
rect 19119 4493 19185 4516
rect 18799 4474 19185 4493
rect 5923 4180 5932 4220
rect 5972 4180 9580 4220
rect 9620 4180 9629 4220
rect 4919 3823 5305 3842
rect 4919 3800 4985 3823
rect 5071 3800 5153 3823
rect 5239 3800 5305 3823
rect 20039 3823 20425 3842
rect 20039 3800 20105 3823
rect 20191 3800 20273 3823
rect 20359 3800 20425 3823
rect 4919 3760 4928 3800
rect 4968 3760 4985 3800
rect 5071 3760 5092 3800
rect 5132 3760 5153 3800
rect 5239 3760 5256 3800
rect 5296 3760 5305 3800
rect 8707 3760 8716 3800
rect 8756 3760 14188 3800
rect 14228 3760 14237 3800
rect 20039 3760 20048 3800
rect 20088 3760 20105 3800
rect 20191 3760 20212 3800
rect 20252 3760 20273 3800
rect 20359 3760 20376 3800
rect 20416 3760 20425 3800
rect 4919 3737 4985 3760
rect 5071 3737 5153 3760
rect 5239 3737 5305 3760
rect 4919 3718 5305 3737
rect 20039 3737 20105 3760
rect 20191 3737 20273 3760
rect 20359 3737 20425 3760
rect 20039 3718 20425 3737
rect 6883 3676 6892 3716
rect 6932 3676 13804 3716
rect 13844 3676 13853 3716
rect 3907 3256 3916 3296
rect 3956 3256 4588 3296
rect 4628 3256 20908 3296
rect 20948 3256 20957 3296
rect 6019 3172 6028 3212
rect 6068 3172 20812 3212
rect 20852 3172 20861 3212
rect 3679 3067 4065 3086
rect 3679 3044 3745 3067
rect 3831 3044 3913 3067
rect 3999 3044 4065 3067
rect 3679 3004 3688 3044
rect 3728 3004 3745 3044
rect 3831 3004 3852 3044
rect 3892 3004 3913 3044
rect 3999 3004 4016 3044
rect 4056 3004 4065 3044
rect 3679 2981 3745 3004
rect 3831 2981 3913 3004
rect 3999 2981 4065 3004
rect 3679 2962 4065 2981
rect 18799 3067 19185 3086
rect 18799 3044 18865 3067
rect 18951 3044 19033 3067
rect 19119 3044 19185 3067
rect 18799 3004 18808 3044
rect 18848 3004 18865 3044
rect 18951 3004 18972 3044
rect 19012 3004 19033 3044
rect 19119 3004 19136 3044
rect 19176 3004 19185 3044
rect 18799 2981 18865 3004
rect 18951 2981 19033 3004
rect 19119 2981 19185 3004
rect 18799 2962 19185 2981
rect 6691 2332 6700 2372
rect 6740 2332 7852 2372
rect 7892 2332 7901 2372
rect 4919 2311 5305 2330
rect 4919 2288 4985 2311
rect 5071 2288 5153 2311
rect 5239 2288 5305 2311
rect 20039 2311 20425 2330
rect 20039 2288 20105 2311
rect 20191 2288 20273 2311
rect 20359 2288 20425 2311
rect 4919 2248 4928 2288
rect 4968 2248 4985 2288
rect 5071 2248 5092 2288
rect 5132 2248 5153 2288
rect 5239 2248 5256 2288
rect 5296 2248 5305 2288
rect 5539 2248 5548 2288
rect 5588 2248 13900 2288
rect 13940 2248 13949 2288
rect 20039 2248 20048 2288
rect 20088 2248 20105 2288
rect 20191 2248 20212 2288
rect 20252 2248 20273 2288
rect 20359 2248 20376 2288
rect 20416 2248 20425 2288
rect 4919 2225 4985 2248
rect 5071 2225 5153 2248
rect 5239 2225 5305 2248
rect 4919 2206 5305 2225
rect 20039 2225 20105 2248
rect 20191 2225 20273 2248
rect 20359 2225 20425 2248
rect 20039 2206 20425 2225
rect 7459 1828 7468 1868
rect 7508 1828 8620 1868
rect 8660 1828 8669 1868
rect 3679 1555 4065 1574
rect 3679 1532 3745 1555
rect 3831 1532 3913 1555
rect 3999 1532 4065 1555
rect 3679 1492 3688 1532
rect 3728 1492 3745 1532
rect 3831 1492 3852 1532
rect 3892 1492 3913 1532
rect 3999 1492 4016 1532
rect 4056 1492 4065 1532
rect 3679 1469 3745 1492
rect 3831 1469 3913 1492
rect 3999 1469 4065 1492
rect 3679 1450 4065 1469
rect 18799 1555 19185 1574
rect 18799 1532 18865 1555
rect 18951 1532 19033 1555
rect 19119 1532 19185 1555
rect 18799 1492 18808 1532
rect 18848 1492 18865 1532
rect 18951 1492 18972 1532
rect 19012 1492 19033 1532
rect 19119 1492 19136 1532
rect 19176 1492 19185 1532
rect 18799 1469 18865 1492
rect 18951 1469 19033 1492
rect 19119 1469 19185 1492
rect 18799 1450 19185 1469
rect 12355 1408 12364 1448
rect 12404 1408 18124 1448
rect 18164 1408 18173 1448
rect 4099 1324 4108 1364
rect 4148 1324 9676 1364
rect 9716 1324 9725 1364
rect 4675 1240 4684 1280
rect 4724 1240 8428 1280
rect 8468 1240 8477 1280
rect 13507 988 13516 1028
rect 13556 988 15148 1028
rect 15188 988 15197 1028
rect 7939 904 7948 944
rect 7988 904 11500 944
rect 11540 904 11549 944
rect 17138 883 17262 902
rect 17138 860 17157 883
rect 14275 820 14284 860
rect 14324 820 17157 860
rect 4919 799 5305 818
rect 4919 776 4985 799
rect 5071 776 5153 799
rect 5239 776 5305 799
rect 17138 797 17157 820
rect 17243 797 17262 883
rect 17138 778 17262 797
rect 20039 799 20425 818
rect 20039 776 20105 799
rect 20191 776 20273 799
rect 20359 776 20425 799
rect 4919 736 4928 776
rect 4968 736 4985 776
rect 5071 736 5092 776
rect 5132 736 5153 776
rect 5239 736 5256 776
rect 5296 736 5305 776
rect 13699 736 13708 776
rect 13748 736 16012 776
rect 16052 736 16061 776
rect 20039 736 20048 776
rect 20088 736 20105 776
rect 20191 736 20212 776
rect 20252 736 20273 776
rect 20359 736 20376 776
rect 20416 736 20425 776
rect 4919 713 4985 736
rect 5071 713 5153 736
rect 5239 713 5305 736
rect 4919 694 5305 713
rect 20039 713 20105 736
rect 20191 713 20273 736
rect 20359 713 20425 736
rect 20039 694 20425 713
rect 8131 568 8140 608
rect 8180 568 12940 608
rect 12980 568 12989 608
rect 1987 400 1996 440
rect 2036 400 6412 440
rect 6452 400 6461 440
rect 14083 316 14092 356
rect 14132 316 16492 356
rect 16532 316 16541 356
<< via5 >>
rect 4985 41600 5071 41623
rect 5153 41600 5239 41623
rect 4985 41560 5010 41600
rect 5010 41560 5050 41600
rect 5050 41560 5071 41600
rect 5153 41560 5174 41600
rect 5174 41560 5214 41600
rect 5214 41560 5239 41600
rect 4985 41537 5071 41560
rect 5153 41537 5239 41560
rect 20105 41600 20191 41623
rect 20273 41600 20359 41623
rect 20105 41560 20130 41600
rect 20130 41560 20170 41600
rect 20170 41560 20191 41600
rect 20273 41560 20294 41600
rect 20294 41560 20334 41600
rect 20334 41560 20359 41600
rect 20105 41537 20191 41560
rect 20273 41537 20359 41560
rect 3745 40844 3831 40867
rect 3913 40844 3999 40867
rect 3745 40804 3770 40844
rect 3770 40804 3810 40844
rect 3810 40804 3831 40844
rect 3913 40804 3934 40844
rect 3934 40804 3974 40844
rect 3974 40804 3999 40844
rect 3745 40781 3831 40804
rect 3913 40781 3999 40804
rect 18865 40844 18951 40867
rect 19033 40844 19119 40867
rect 18865 40804 18890 40844
rect 18890 40804 18930 40844
rect 18930 40804 18951 40844
rect 19033 40804 19054 40844
rect 19054 40804 19094 40844
rect 19094 40804 19119 40844
rect 18865 40781 18951 40804
rect 19033 40781 19119 40804
rect 12141 40445 12227 40531
rect 4985 40088 5071 40111
rect 5153 40088 5239 40111
rect 4985 40048 5010 40088
rect 5010 40048 5050 40088
rect 5050 40048 5071 40088
rect 5153 40048 5174 40088
rect 5174 40048 5214 40088
rect 5214 40048 5239 40088
rect 4985 40025 5071 40048
rect 5153 40025 5239 40048
rect 20105 40088 20191 40111
rect 20273 40088 20359 40111
rect 20105 40048 20130 40088
rect 20130 40048 20170 40088
rect 20170 40048 20191 40088
rect 20273 40048 20294 40088
rect 20294 40048 20334 40088
rect 20334 40048 20359 40088
rect 20105 40025 20191 40048
rect 20273 40025 20359 40048
rect 17157 39836 17243 39859
rect 17157 39796 17164 39836
rect 17164 39796 17204 39836
rect 17204 39796 17243 39836
rect 17157 39773 17243 39796
rect 3745 39332 3831 39355
rect 3913 39332 3999 39355
rect 3745 39292 3770 39332
rect 3770 39292 3810 39332
rect 3810 39292 3831 39332
rect 3913 39292 3934 39332
rect 3934 39292 3974 39332
rect 3974 39292 3999 39332
rect 3745 39269 3831 39292
rect 3913 39269 3999 39292
rect 18865 39332 18951 39355
rect 19033 39332 19119 39355
rect 18865 39292 18890 39332
rect 18890 39292 18930 39332
rect 18930 39292 18951 39332
rect 19033 39292 19054 39332
rect 19054 39292 19094 39332
rect 19094 39292 19119 39332
rect 18865 39269 18951 39292
rect 19033 39269 19119 39292
rect 4985 38576 5071 38599
rect 5153 38576 5239 38599
rect 4985 38536 5010 38576
rect 5010 38536 5050 38576
rect 5050 38536 5071 38576
rect 5153 38536 5174 38576
rect 5174 38536 5214 38576
rect 5214 38536 5239 38576
rect 4985 38513 5071 38536
rect 5153 38513 5239 38536
rect 20105 38576 20191 38599
rect 20273 38576 20359 38599
rect 20105 38536 20130 38576
rect 20130 38536 20170 38576
rect 20170 38536 20191 38576
rect 20273 38536 20294 38576
rect 20294 38536 20334 38576
rect 20334 38536 20359 38576
rect 20105 38513 20191 38536
rect 20273 38513 20359 38536
rect 3745 37820 3831 37843
rect 3913 37820 3999 37843
rect 3745 37780 3770 37820
rect 3770 37780 3810 37820
rect 3810 37780 3831 37820
rect 3913 37780 3934 37820
rect 3934 37780 3974 37820
rect 3974 37780 3999 37820
rect 3745 37757 3831 37780
rect 3913 37757 3999 37780
rect 18865 37820 18951 37843
rect 19033 37820 19119 37843
rect 18865 37780 18890 37820
rect 18890 37780 18930 37820
rect 18930 37780 18951 37820
rect 19033 37780 19054 37820
rect 19054 37780 19094 37820
rect 19094 37780 19119 37820
rect 18865 37757 18951 37780
rect 19033 37757 19119 37780
rect 4985 37064 5071 37087
rect 5153 37064 5239 37087
rect 4985 37024 5010 37064
rect 5010 37024 5050 37064
rect 5050 37024 5071 37064
rect 5153 37024 5174 37064
rect 5174 37024 5214 37064
rect 5214 37024 5239 37064
rect 4985 37001 5071 37024
rect 5153 37001 5239 37024
rect 20105 37064 20191 37087
rect 20273 37064 20359 37087
rect 20105 37024 20130 37064
rect 20130 37024 20170 37064
rect 20170 37024 20191 37064
rect 20273 37024 20294 37064
rect 20294 37024 20334 37064
rect 20334 37024 20359 37064
rect 20105 37001 20191 37024
rect 20273 37001 20359 37024
rect 3745 36308 3831 36331
rect 3913 36308 3999 36331
rect 3745 36268 3770 36308
rect 3770 36268 3810 36308
rect 3810 36268 3831 36308
rect 3913 36268 3934 36308
rect 3934 36268 3974 36308
rect 3974 36268 3999 36308
rect 3745 36245 3831 36268
rect 3913 36245 3999 36268
rect 18865 36308 18951 36331
rect 19033 36308 19119 36331
rect 18865 36268 18890 36308
rect 18890 36268 18930 36308
rect 18930 36268 18951 36308
rect 19033 36268 19054 36308
rect 19054 36268 19094 36308
rect 19094 36268 19119 36308
rect 18865 36245 18951 36268
rect 19033 36245 19119 36268
rect 4985 35552 5071 35575
rect 5153 35552 5239 35575
rect 4985 35512 5010 35552
rect 5010 35512 5050 35552
rect 5050 35512 5071 35552
rect 5153 35512 5174 35552
rect 5174 35512 5214 35552
rect 5214 35512 5239 35552
rect 4985 35489 5071 35512
rect 5153 35489 5239 35512
rect 20105 35552 20191 35575
rect 20273 35552 20359 35575
rect 20105 35512 20130 35552
rect 20130 35512 20170 35552
rect 20170 35512 20191 35552
rect 20273 35512 20294 35552
rect 20294 35512 20334 35552
rect 20334 35512 20359 35552
rect 20105 35489 20191 35512
rect 20273 35489 20359 35512
rect 3745 34796 3831 34819
rect 3913 34796 3999 34819
rect 3745 34756 3770 34796
rect 3770 34756 3810 34796
rect 3810 34756 3831 34796
rect 3913 34756 3934 34796
rect 3934 34756 3974 34796
rect 3974 34756 3999 34796
rect 3745 34733 3831 34756
rect 3913 34733 3999 34756
rect 18865 34796 18951 34819
rect 19033 34796 19119 34819
rect 18865 34756 18890 34796
rect 18890 34756 18930 34796
rect 18930 34756 18951 34796
rect 19033 34756 19054 34796
rect 19054 34756 19094 34796
rect 19094 34756 19119 34796
rect 18865 34733 18951 34756
rect 19033 34733 19119 34756
rect 4985 34040 5071 34063
rect 5153 34040 5239 34063
rect 4985 34000 5010 34040
rect 5010 34000 5050 34040
rect 5050 34000 5071 34040
rect 5153 34000 5174 34040
rect 5174 34000 5214 34040
rect 5214 34000 5239 34040
rect 4985 33977 5071 34000
rect 5153 33977 5239 34000
rect 20105 34040 20191 34063
rect 20273 34040 20359 34063
rect 20105 34000 20130 34040
rect 20130 34000 20170 34040
rect 20170 34000 20191 34040
rect 20273 34000 20294 34040
rect 20294 34000 20334 34040
rect 20334 34000 20359 34040
rect 20105 33977 20191 34000
rect 20273 33977 20359 34000
rect 3745 33284 3831 33307
rect 3913 33284 3999 33307
rect 3745 33244 3770 33284
rect 3770 33244 3810 33284
rect 3810 33244 3831 33284
rect 3913 33244 3934 33284
rect 3934 33244 3974 33284
rect 3974 33244 3999 33284
rect 3745 33221 3831 33244
rect 3913 33221 3999 33244
rect 18865 33284 18951 33307
rect 19033 33284 19119 33307
rect 18865 33244 18890 33284
rect 18890 33244 18930 33284
rect 18930 33244 18951 33284
rect 19033 33244 19054 33284
rect 19054 33244 19094 33284
rect 19094 33244 19119 33284
rect 18865 33221 18951 33244
rect 19033 33221 19119 33244
rect 4985 32528 5071 32551
rect 5153 32528 5239 32551
rect 4985 32488 5010 32528
rect 5010 32488 5050 32528
rect 5050 32488 5071 32528
rect 5153 32488 5174 32528
rect 5174 32488 5214 32528
rect 5214 32488 5239 32528
rect 4985 32465 5071 32488
rect 5153 32465 5239 32488
rect 20105 32528 20191 32551
rect 20273 32528 20359 32551
rect 20105 32488 20130 32528
rect 20130 32488 20170 32528
rect 20170 32488 20191 32528
rect 20273 32488 20294 32528
rect 20294 32488 20334 32528
rect 20334 32488 20359 32528
rect 20105 32465 20191 32488
rect 20273 32465 20359 32488
rect 3745 31772 3831 31795
rect 3913 31772 3999 31795
rect 3745 31732 3770 31772
rect 3770 31732 3810 31772
rect 3810 31732 3831 31772
rect 3913 31732 3934 31772
rect 3934 31732 3974 31772
rect 3974 31732 3999 31772
rect 3745 31709 3831 31732
rect 3913 31709 3999 31732
rect 18865 31772 18951 31795
rect 19033 31772 19119 31795
rect 18865 31732 18890 31772
rect 18890 31732 18930 31772
rect 18930 31732 18951 31772
rect 19033 31732 19054 31772
rect 19054 31732 19094 31772
rect 19094 31732 19119 31772
rect 18865 31709 18951 31732
rect 19033 31709 19119 31732
rect 4985 31016 5071 31039
rect 5153 31016 5239 31039
rect 4985 30976 5010 31016
rect 5010 30976 5050 31016
rect 5050 30976 5071 31016
rect 5153 30976 5174 31016
rect 5174 30976 5214 31016
rect 5214 30976 5239 31016
rect 4985 30953 5071 30976
rect 5153 30953 5239 30976
rect 20105 31016 20191 31039
rect 20273 31016 20359 31039
rect 20105 30976 20130 31016
rect 20130 30976 20170 31016
rect 20170 30976 20191 31016
rect 20273 30976 20294 31016
rect 20294 30976 20334 31016
rect 20334 30976 20359 31016
rect 20105 30953 20191 30976
rect 20273 30953 20359 30976
rect 3745 30260 3831 30283
rect 3913 30260 3999 30283
rect 3745 30220 3770 30260
rect 3770 30220 3810 30260
rect 3810 30220 3831 30260
rect 3913 30220 3934 30260
rect 3934 30220 3974 30260
rect 3974 30220 3999 30260
rect 3745 30197 3831 30220
rect 3913 30197 3999 30220
rect 18865 30260 18951 30283
rect 19033 30260 19119 30283
rect 18865 30220 18890 30260
rect 18890 30220 18930 30260
rect 18930 30220 18951 30260
rect 19033 30220 19054 30260
rect 19054 30220 19094 30260
rect 19094 30220 19119 30260
rect 18865 30197 18951 30220
rect 19033 30197 19119 30220
rect 4985 29504 5071 29527
rect 5153 29504 5239 29527
rect 4985 29464 5010 29504
rect 5010 29464 5050 29504
rect 5050 29464 5071 29504
rect 5153 29464 5174 29504
rect 5174 29464 5214 29504
rect 5214 29464 5239 29504
rect 4985 29441 5071 29464
rect 5153 29441 5239 29464
rect 20105 29504 20191 29527
rect 20273 29504 20359 29527
rect 20105 29464 20130 29504
rect 20130 29464 20170 29504
rect 20170 29464 20191 29504
rect 20273 29464 20294 29504
rect 20294 29464 20334 29504
rect 20334 29464 20359 29504
rect 20105 29441 20191 29464
rect 20273 29441 20359 29464
rect 3745 28748 3831 28771
rect 3913 28748 3999 28771
rect 3745 28708 3770 28748
rect 3770 28708 3810 28748
rect 3810 28708 3831 28748
rect 3913 28708 3934 28748
rect 3934 28708 3974 28748
rect 3974 28708 3999 28748
rect 3745 28685 3831 28708
rect 3913 28685 3999 28708
rect 18865 28748 18951 28771
rect 19033 28748 19119 28771
rect 18865 28708 18890 28748
rect 18890 28708 18930 28748
rect 18930 28708 18951 28748
rect 19033 28708 19054 28748
rect 19054 28708 19094 28748
rect 19094 28708 19119 28748
rect 18865 28685 18951 28708
rect 19033 28685 19119 28708
rect 4985 27992 5071 28015
rect 5153 27992 5239 28015
rect 4985 27952 5010 27992
rect 5010 27952 5050 27992
rect 5050 27952 5071 27992
rect 5153 27952 5174 27992
rect 5174 27952 5214 27992
rect 5214 27952 5239 27992
rect 4985 27929 5071 27952
rect 5153 27929 5239 27952
rect 20105 27992 20191 28015
rect 20273 27992 20359 28015
rect 20105 27952 20130 27992
rect 20130 27952 20170 27992
rect 20170 27952 20191 27992
rect 20273 27952 20294 27992
rect 20294 27952 20334 27992
rect 20334 27952 20359 27992
rect 20105 27929 20191 27952
rect 20273 27929 20359 27952
rect 3745 27236 3831 27259
rect 3913 27236 3999 27259
rect 3745 27196 3770 27236
rect 3770 27196 3810 27236
rect 3810 27196 3831 27236
rect 3913 27196 3934 27236
rect 3934 27196 3974 27236
rect 3974 27196 3999 27236
rect 3745 27173 3831 27196
rect 3913 27173 3999 27196
rect 18865 27236 18951 27259
rect 19033 27236 19119 27259
rect 18865 27196 18890 27236
rect 18890 27196 18930 27236
rect 18930 27196 18951 27236
rect 19033 27196 19054 27236
rect 19054 27196 19094 27236
rect 19094 27196 19119 27236
rect 18865 27173 18951 27196
rect 19033 27173 19119 27196
rect 4985 26480 5071 26503
rect 5153 26480 5239 26503
rect 4985 26440 5010 26480
rect 5010 26440 5050 26480
rect 5050 26440 5071 26480
rect 5153 26440 5174 26480
rect 5174 26440 5214 26480
rect 5214 26440 5239 26480
rect 4985 26417 5071 26440
rect 5153 26417 5239 26440
rect 20105 26480 20191 26503
rect 20273 26480 20359 26503
rect 20105 26440 20130 26480
rect 20130 26440 20170 26480
rect 20170 26440 20191 26480
rect 20273 26440 20294 26480
rect 20294 26440 20334 26480
rect 20334 26440 20359 26480
rect 20105 26417 20191 26440
rect 20273 26417 20359 26440
rect 3745 25724 3831 25747
rect 3913 25724 3999 25747
rect 3745 25684 3770 25724
rect 3770 25684 3810 25724
rect 3810 25684 3831 25724
rect 3913 25684 3934 25724
rect 3934 25684 3974 25724
rect 3974 25684 3999 25724
rect 3745 25661 3831 25684
rect 3913 25661 3999 25684
rect 18865 25724 18951 25747
rect 19033 25724 19119 25747
rect 18865 25684 18890 25724
rect 18890 25684 18930 25724
rect 18930 25684 18951 25724
rect 19033 25684 19054 25724
rect 19054 25684 19094 25724
rect 19094 25684 19119 25724
rect 18865 25661 18951 25684
rect 19033 25661 19119 25684
rect 4985 24968 5071 24991
rect 5153 24968 5239 24991
rect 4985 24928 5010 24968
rect 5010 24928 5050 24968
rect 5050 24928 5071 24968
rect 5153 24928 5174 24968
rect 5174 24928 5214 24968
rect 5214 24928 5239 24968
rect 4985 24905 5071 24928
rect 5153 24905 5239 24928
rect 20105 24968 20191 24991
rect 20273 24968 20359 24991
rect 20105 24928 20130 24968
rect 20130 24928 20170 24968
rect 20170 24928 20191 24968
rect 20273 24928 20294 24968
rect 20294 24928 20334 24968
rect 20334 24928 20359 24968
rect 20105 24905 20191 24928
rect 20273 24905 20359 24928
rect 3745 24212 3831 24235
rect 3913 24212 3999 24235
rect 3745 24172 3770 24212
rect 3770 24172 3810 24212
rect 3810 24172 3831 24212
rect 3913 24172 3934 24212
rect 3934 24172 3974 24212
rect 3974 24172 3999 24212
rect 3745 24149 3831 24172
rect 3913 24149 3999 24172
rect 18865 24212 18951 24235
rect 19033 24212 19119 24235
rect 18865 24172 18890 24212
rect 18890 24172 18930 24212
rect 18930 24172 18951 24212
rect 19033 24172 19054 24212
rect 19054 24172 19094 24212
rect 19094 24172 19119 24212
rect 18865 24149 18951 24172
rect 19033 24149 19119 24172
rect 4985 23456 5071 23479
rect 5153 23456 5239 23479
rect 4985 23416 5010 23456
rect 5010 23416 5050 23456
rect 5050 23416 5071 23456
rect 5153 23416 5174 23456
rect 5174 23416 5214 23456
rect 5214 23416 5239 23456
rect 4985 23393 5071 23416
rect 5153 23393 5239 23416
rect 20105 23456 20191 23479
rect 20273 23456 20359 23479
rect 20105 23416 20130 23456
rect 20130 23416 20170 23456
rect 20170 23416 20191 23456
rect 20273 23416 20294 23456
rect 20294 23416 20334 23456
rect 20334 23416 20359 23456
rect 20105 23393 20191 23416
rect 20273 23393 20359 23416
rect 3745 22700 3831 22723
rect 3913 22700 3999 22723
rect 3745 22660 3770 22700
rect 3770 22660 3810 22700
rect 3810 22660 3831 22700
rect 3913 22660 3934 22700
rect 3934 22660 3974 22700
rect 3974 22660 3999 22700
rect 3745 22637 3831 22660
rect 3913 22637 3999 22660
rect 18865 22700 18951 22723
rect 19033 22700 19119 22723
rect 18865 22660 18890 22700
rect 18890 22660 18930 22700
rect 18930 22660 18951 22700
rect 19033 22660 19054 22700
rect 19054 22660 19094 22700
rect 19094 22660 19119 22700
rect 18865 22637 18951 22660
rect 19033 22637 19119 22660
rect 4985 21944 5071 21967
rect 5153 21944 5239 21967
rect 4985 21904 5010 21944
rect 5010 21904 5050 21944
rect 5050 21904 5071 21944
rect 5153 21904 5174 21944
rect 5174 21904 5214 21944
rect 5214 21904 5239 21944
rect 4985 21881 5071 21904
rect 5153 21881 5239 21904
rect 20105 21944 20191 21967
rect 20273 21944 20359 21967
rect 20105 21904 20130 21944
rect 20130 21904 20170 21944
rect 20170 21904 20191 21944
rect 20273 21904 20294 21944
rect 20294 21904 20334 21944
rect 20334 21904 20359 21944
rect 20105 21881 20191 21904
rect 20273 21881 20359 21904
rect 3745 21188 3831 21211
rect 3913 21188 3999 21211
rect 3745 21148 3770 21188
rect 3770 21148 3810 21188
rect 3810 21148 3831 21188
rect 3913 21148 3934 21188
rect 3934 21148 3974 21188
rect 3974 21148 3999 21188
rect 3745 21125 3831 21148
rect 3913 21125 3999 21148
rect 18865 21188 18951 21211
rect 19033 21188 19119 21211
rect 18865 21148 18890 21188
rect 18890 21148 18930 21188
rect 18930 21148 18951 21188
rect 19033 21148 19054 21188
rect 19054 21148 19094 21188
rect 19094 21148 19119 21188
rect 18865 21125 18951 21148
rect 19033 21125 19119 21148
rect 4985 20432 5071 20455
rect 5153 20432 5239 20455
rect 4985 20392 5010 20432
rect 5010 20392 5050 20432
rect 5050 20392 5071 20432
rect 5153 20392 5174 20432
rect 5174 20392 5214 20432
rect 5214 20392 5239 20432
rect 4985 20369 5071 20392
rect 5153 20369 5239 20392
rect 20105 20432 20191 20455
rect 20273 20432 20359 20455
rect 20105 20392 20130 20432
rect 20130 20392 20170 20432
rect 20170 20392 20191 20432
rect 20273 20392 20294 20432
rect 20294 20392 20334 20432
rect 20334 20392 20359 20432
rect 20105 20369 20191 20392
rect 20273 20369 20359 20392
rect 3745 19676 3831 19699
rect 3913 19676 3999 19699
rect 3745 19636 3770 19676
rect 3770 19636 3810 19676
rect 3810 19636 3831 19676
rect 3913 19636 3934 19676
rect 3934 19636 3974 19676
rect 3974 19636 3999 19676
rect 3745 19613 3831 19636
rect 3913 19613 3999 19636
rect 18865 19676 18951 19699
rect 19033 19676 19119 19699
rect 18865 19636 18890 19676
rect 18890 19636 18930 19676
rect 18930 19636 18951 19676
rect 19033 19636 19054 19676
rect 19054 19636 19094 19676
rect 19094 19636 19119 19676
rect 18865 19613 18951 19636
rect 19033 19613 19119 19636
rect 4985 18920 5071 18943
rect 5153 18920 5239 18943
rect 4985 18880 5010 18920
rect 5010 18880 5050 18920
rect 5050 18880 5071 18920
rect 5153 18880 5174 18920
rect 5174 18880 5214 18920
rect 5214 18880 5239 18920
rect 4985 18857 5071 18880
rect 5153 18857 5239 18880
rect 20105 18920 20191 18943
rect 20273 18920 20359 18943
rect 20105 18880 20130 18920
rect 20130 18880 20170 18920
rect 20170 18880 20191 18920
rect 20273 18880 20294 18920
rect 20294 18880 20334 18920
rect 20334 18880 20359 18920
rect 20105 18857 20191 18880
rect 20273 18857 20359 18880
rect 3745 18164 3831 18187
rect 3913 18164 3999 18187
rect 3745 18124 3770 18164
rect 3770 18124 3810 18164
rect 3810 18124 3831 18164
rect 3913 18124 3934 18164
rect 3934 18124 3974 18164
rect 3974 18124 3999 18164
rect 3745 18101 3831 18124
rect 3913 18101 3999 18124
rect 18865 18164 18951 18187
rect 19033 18164 19119 18187
rect 18865 18124 18890 18164
rect 18890 18124 18930 18164
rect 18930 18124 18951 18164
rect 19033 18124 19054 18164
rect 19054 18124 19094 18164
rect 19094 18124 19119 18164
rect 18865 18101 18951 18124
rect 19033 18101 19119 18124
rect 4985 17408 5071 17431
rect 5153 17408 5239 17431
rect 4985 17368 5010 17408
rect 5010 17368 5050 17408
rect 5050 17368 5071 17408
rect 5153 17368 5174 17408
rect 5174 17368 5214 17408
rect 5214 17368 5239 17408
rect 4985 17345 5071 17368
rect 5153 17345 5239 17368
rect 20105 17408 20191 17431
rect 20273 17408 20359 17431
rect 20105 17368 20130 17408
rect 20130 17368 20170 17408
rect 20170 17368 20191 17408
rect 20273 17368 20294 17408
rect 20294 17368 20334 17408
rect 20334 17368 20359 17408
rect 20105 17345 20191 17368
rect 20273 17345 20359 17368
rect 3745 16652 3831 16675
rect 3913 16652 3999 16675
rect 18865 16652 18951 16675
rect 19033 16652 19119 16675
rect 3745 16612 3770 16652
rect 3770 16612 3810 16652
rect 3810 16612 3831 16652
rect 3913 16612 3934 16652
rect 3934 16612 3974 16652
rect 3974 16612 3999 16652
rect 18865 16612 18890 16652
rect 18890 16612 18930 16652
rect 18930 16612 18951 16652
rect 19033 16612 19054 16652
rect 19054 16612 19094 16652
rect 19094 16612 19119 16652
rect 3745 16589 3831 16612
rect 3913 16589 3999 16612
rect 18865 16589 18951 16612
rect 19033 16589 19119 16612
rect 4985 15896 5071 15919
rect 5153 15896 5239 15919
rect 4985 15856 5010 15896
rect 5010 15856 5050 15896
rect 5050 15856 5071 15896
rect 5153 15856 5174 15896
rect 5174 15856 5214 15896
rect 5214 15856 5239 15896
rect 4985 15833 5071 15856
rect 5153 15833 5239 15856
rect 20105 15896 20191 15919
rect 20273 15896 20359 15919
rect 20105 15856 20130 15896
rect 20130 15856 20170 15896
rect 20170 15856 20191 15896
rect 20273 15856 20294 15896
rect 20294 15856 20334 15896
rect 20334 15856 20359 15896
rect 20105 15833 20191 15856
rect 20273 15833 20359 15856
rect 3745 15140 3831 15163
rect 3913 15140 3999 15163
rect 3745 15100 3770 15140
rect 3770 15100 3810 15140
rect 3810 15100 3831 15140
rect 3913 15100 3934 15140
rect 3934 15100 3974 15140
rect 3974 15100 3999 15140
rect 3745 15077 3831 15100
rect 3913 15077 3999 15100
rect 18865 15140 18951 15163
rect 19033 15140 19119 15163
rect 18865 15100 18890 15140
rect 18890 15100 18930 15140
rect 18930 15100 18951 15140
rect 19033 15100 19054 15140
rect 19054 15100 19094 15140
rect 19094 15100 19119 15140
rect 18865 15077 18951 15100
rect 19033 15077 19119 15100
rect 4985 14384 5071 14407
rect 5153 14384 5239 14407
rect 4985 14344 5010 14384
rect 5010 14344 5050 14384
rect 5050 14344 5071 14384
rect 5153 14344 5174 14384
rect 5174 14344 5214 14384
rect 5214 14344 5239 14384
rect 4985 14321 5071 14344
rect 5153 14321 5239 14344
rect 20105 14384 20191 14407
rect 20273 14384 20359 14407
rect 20105 14344 20130 14384
rect 20130 14344 20170 14384
rect 20170 14344 20191 14384
rect 20273 14344 20294 14384
rect 20294 14344 20334 14384
rect 20334 14344 20359 14384
rect 20105 14321 20191 14344
rect 20273 14321 20359 14344
rect 3745 13628 3831 13651
rect 3913 13628 3999 13651
rect 3745 13588 3770 13628
rect 3770 13588 3810 13628
rect 3810 13588 3831 13628
rect 3913 13588 3934 13628
rect 3934 13588 3974 13628
rect 3974 13588 3999 13628
rect 3745 13565 3831 13588
rect 3913 13565 3999 13588
rect 18865 13628 18951 13651
rect 19033 13628 19119 13651
rect 18865 13588 18890 13628
rect 18890 13588 18930 13628
rect 18930 13588 18951 13628
rect 19033 13588 19054 13628
rect 19054 13588 19094 13628
rect 19094 13588 19119 13628
rect 18865 13565 18951 13588
rect 19033 13565 19119 13588
rect 4985 12872 5071 12895
rect 5153 12872 5239 12895
rect 4985 12832 5010 12872
rect 5010 12832 5050 12872
rect 5050 12832 5071 12872
rect 5153 12832 5174 12872
rect 5174 12832 5214 12872
rect 5214 12832 5239 12872
rect 4985 12809 5071 12832
rect 5153 12809 5239 12832
rect 20105 12872 20191 12895
rect 20273 12872 20359 12895
rect 20105 12832 20130 12872
rect 20130 12832 20170 12872
rect 20170 12832 20191 12872
rect 20273 12832 20294 12872
rect 20294 12832 20334 12872
rect 20334 12832 20359 12872
rect 20105 12809 20191 12832
rect 20273 12809 20359 12832
rect 3745 12116 3831 12139
rect 3913 12116 3999 12139
rect 3745 12076 3770 12116
rect 3770 12076 3810 12116
rect 3810 12076 3831 12116
rect 3913 12076 3934 12116
rect 3934 12076 3974 12116
rect 3974 12076 3999 12116
rect 3745 12053 3831 12076
rect 3913 12053 3999 12076
rect 18865 12116 18951 12139
rect 19033 12116 19119 12139
rect 18865 12076 18890 12116
rect 18890 12076 18930 12116
rect 18930 12076 18951 12116
rect 19033 12076 19054 12116
rect 19054 12076 19094 12116
rect 19094 12076 19119 12116
rect 18865 12053 18951 12076
rect 19033 12053 19119 12076
rect 4985 11360 5071 11383
rect 5153 11360 5239 11383
rect 4985 11320 5010 11360
rect 5010 11320 5050 11360
rect 5050 11320 5071 11360
rect 5153 11320 5174 11360
rect 5174 11320 5214 11360
rect 5214 11320 5239 11360
rect 4985 11297 5071 11320
rect 5153 11297 5239 11320
rect 20105 11360 20191 11383
rect 20273 11360 20359 11383
rect 20105 11320 20130 11360
rect 20130 11320 20170 11360
rect 20170 11320 20191 11360
rect 20273 11320 20294 11360
rect 20294 11320 20334 11360
rect 20334 11320 20359 11360
rect 20105 11297 20191 11320
rect 20273 11297 20359 11320
rect 3745 10604 3831 10627
rect 3913 10604 3999 10627
rect 3745 10564 3770 10604
rect 3770 10564 3810 10604
rect 3810 10564 3831 10604
rect 3913 10564 3934 10604
rect 3934 10564 3974 10604
rect 3974 10564 3999 10604
rect 3745 10541 3831 10564
rect 3913 10541 3999 10564
rect 18865 10604 18951 10627
rect 19033 10604 19119 10627
rect 18865 10564 18890 10604
rect 18890 10564 18930 10604
rect 18930 10564 18951 10604
rect 19033 10564 19054 10604
rect 19054 10564 19094 10604
rect 19094 10564 19119 10604
rect 18865 10541 18951 10564
rect 19033 10541 19119 10564
rect 4985 9848 5071 9871
rect 5153 9848 5239 9871
rect 4985 9808 5010 9848
rect 5010 9808 5050 9848
rect 5050 9808 5071 9848
rect 5153 9808 5174 9848
rect 5174 9808 5214 9848
rect 5214 9808 5239 9848
rect 4985 9785 5071 9808
rect 5153 9785 5239 9808
rect 20105 9848 20191 9871
rect 20273 9848 20359 9871
rect 20105 9808 20130 9848
rect 20130 9808 20170 9848
rect 20170 9808 20191 9848
rect 20273 9808 20294 9848
rect 20294 9808 20334 9848
rect 20334 9808 20359 9848
rect 20105 9785 20191 9808
rect 20273 9785 20359 9808
rect 3745 9092 3831 9115
rect 3913 9092 3999 9115
rect 3745 9052 3770 9092
rect 3770 9052 3810 9092
rect 3810 9052 3831 9092
rect 3913 9052 3934 9092
rect 3934 9052 3974 9092
rect 3974 9052 3999 9092
rect 3745 9029 3831 9052
rect 3913 9029 3999 9052
rect 18865 9092 18951 9115
rect 19033 9092 19119 9115
rect 18865 9052 18890 9092
rect 18890 9052 18930 9092
rect 18930 9052 18951 9092
rect 19033 9052 19054 9092
rect 19054 9052 19094 9092
rect 19094 9052 19119 9092
rect 18865 9029 18951 9052
rect 19033 9029 19119 9052
rect 4985 8336 5071 8359
rect 5153 8336 5239 8359
rect 4985 8296 5010 8336
rect 5010 8296 5050 8336
rect 5050 8296 5071 8336
rect 5153 8296 5174 8336
rect 5174 8296 5214 8336
rect 5214 8296 5239 8336
rect 4985 8273 5071 8296
rect 5153 8273 5239 8296
rect 20105 8336 20191 8359
rect 20273 8336 20359 8359
rect 20105 8296 20130 8336
rect 20130 8296 20170 8336
rect 20170 8296 20191 8336
rect 20273 8296 20294 8336
rect 20294 8296 20334 8336
rect 20334 8296 20359 8336
rect 20105 8273 20191 8296
rect 20273 8273 20359 8296
rect 3745 7580 3831 7603
rect 3913 7580 3999 7603
rect 3745 7540 3770 7580
rect 3770 7540 3810 7580
rect 3810 7540 3831 7580
rect 3913 7540 3934 7580
rect 3934 7540 3974 7580
rect 3974 7540 3999 7580
rect 3745 7517 3831 7540
rect 3913 7517 3999 7540
rect 18865 7580 18951 7603
rect 19033 7580 19119 7603
rect 18865 7540 18890 7580
rect 18890 7540 18930 7580
rect 18930 7540 18951 7580
rect 19033 7540 19054 7580
rect 19054 7540 19094 7580
rect 19094 7540 19119 7580
rect 18865 7517 18951 7540
rect 19033 7517 19119 7540
rect 4985 6824 5071 6847
rect 5153 6824 5239 6847
rect 4985 6784 5010 6824
rect 5010 6784 5050 6824
rect 5050 6784 5071 6824
rect 5153 6784 5174 6824
rect 5174 6784 5214 6824
rect 5214 6784 5239 6824
rect 4985 6761 5071 6784
rect 5153 6761 5239 6784
rect 20105 6824 20191 6847
rect 20273 6824 20359 6847
rect 20105 6784 20130 6824
rect 20130 6784 20170 6824
rect 20170 6784 20191 6824
rect 20273 6784 20294 6824
rect 20294 6784 20334 6824
rect 20334 6784 20359 6824
rect 20105 6761 20191 6784
rect 20273 6761 20359 6784
rect 3745 6068 3831 6091
rect 3913 6068 3999 6091
rect 3745 6028 3770 6068
rect 3770 6028 3810 6068
rect 3810 6028 3831 6068
rect 3913 6028 3934 6068
rect 3934 6028 3974 6068
rect 3974 6028 3999 6068
rect 3745 6005 3831 6028
rect 3913 6005 3999 6028
rect 18865 6068 18951 6091
rect 19033 6068 19119 6091
rect 18865 6028 18890 6068
rect 18890 6028 18930 6068
rect 18930 6028 18951 6068
rect 19033 6028 19054 6068
rect 19054 6028 19094 6068
rect 19094 6028 19119 6068
rect 18865 6005 18951 6028
rect 19033 6005 19119 6028
rect 12141 5753 12227 5839
rect 4985 5312 5071 5335
rect 5153 5312 5239 5335
rect 4985 5272 5010 5312
rect 5010 5272 5050 5312
rect 5050 5272 5071 5312
rect 5153 5272 5174 5312
rect 5174 5272 5214 5312
rect 5214 5272 5239 5312
rect 4985 5249 5071 5272
rect 5153 5249 5239 5272
rect 20105 5312 20191 5335
rect 20273 5312 20359 5335
rect 20105 5272 20130 5312
rect 20130 5272 20170 5312
rect 20170 5272 20191 5312
rect 20273 5272 20294 5312
rect 20294 5272 20334 5312
rect 20334 5272 20359 5312
rect 20105 5249 20191 5272
rect 20273 5249 20359 5272
rect 3745 4556 3831 4579
rect 3913 4556 3999 4579
rect 3745 4516 3770 4556
rect 3770 4516 3810 4556
rect 3810 4516 3831 4556
rect 3913 4516 3934 4556
rect 3934 4516 3974 4556
rect 3974 4516 3999 4556
rect 3745 4493 3831 4516
rect 3913 4493 3999 4516
rect 18865 4556 18951 4579
rect 19033 4556 19119 4579
rect 18865 4516 18890 4556
rect 18890 4516 18930 4556
rect 18930 4516 18951 4556
rect 19033 4516 19054 4556
rect 19054 4516 19094 4556
rect 19094 4516 19119 4556
rect 18865 4493 18951 4516
rect 19033 4493 19119 4516
rect 4985 3800 5071 3823
rect 5153 3800 5239 3823
rect 20105 3800 20191 3823
rect 20273 3800 20359 3823
rect 4985 3760 5010 3800
rect 5010 3760 5050 3800
rect 5050 3760 5071 3800
rect 5153 3760 5174 3800
rect 5174 3760 5214 3800
rect 5214 3760 5239 3800
rect 20105 3760 20130 3800
rect 20130 3760 20170 3800
rect 20170 3760 20191 3800
rect 20273 3760 20294 3800
rect 20294 3760 20334 3800
rect 20334 3760 20359 3800
rect 4985 3737 5071 3760
rect 5153 3737 5239 3760
rect 20105 3737 20191 3760
rect 20273 3737 20359 3760
rect 3745 3044 3831 3067
rect 3913 3044 3999 3067
rect 3745 3004 3770 3044
rect 3770 3004 3810 3044
rect 3810 3004 3831 3044
rect 3913 3004 3934 3044
rect 3934 3004 3974 3044
rect 3974 3004 3999 3044
rect 3745 2981 3831 3004
rect 3913 2981 3999 3004
rect 18865 3044 18951 3067
rect 19033 3044 19119 3067
rect 18865 3004 18890 3044
rect 18890 3004 18930 3044
rect 18930 3004 18951 3044
rect 19033 3004 19054 3044
rect 19054 3004 19094 3044
rect 19094 3004 19119 3044
rect 18865 2981 18951 3004
rect 19033 2981 19119 3004
rect 4985 2288 5071 2311
rect 5153 2288 5239 2311
rect 20105 2288 20191 2311
rect 20273 2288 20359 2311
rect 4985 2248 5010 2288
rect 5010 2248 5050 2288
rect 5050 2248 5071 2288
rect 5153 2248 5174 2288
rect 5174 2248 5214 2288
rect 5214 2248 5239 2288
rect 20105 2248 20130 2288
rect 20130 2248 20170 2288
rect 20170 2248 20191 2288
rect 20273 2248 20294 2288
rect 20294 2248 20334 2288
rect 20334 2248 20359 2288
rect 4985 2225 5071 2248
rect 5153 2225 5239 2248
rect 20105 2225 20191 2248
rect 20273 2225 20359 2248
rect 3745 1532 3831 1555
rect 3913 1532 3999 1555
rect 3745 1492 3770 1532
rect 3770 1492 3810 1532
rect 3810 1492 3831 1532
rect 3913 1492 3934 1532
rect 3934 1492 3974 1532
rect 3974 1492 3999 1532
rect 3745 1469 3831 1492
rect 3913 1469 3999 1492
rect 18865 1532 18951 1555
rect 19033 1532 19119 1555
rect 18865 1492 18890 1532
rect 18890 1492 18930 1532
rect 18930 1492 18951 1532
rect 19033 1492 19054 1532
rect 19054 1492 19094 1532
rect 19094 1492 19119 1532
rect 18865 1469 18951 1492
rect 19033 1469 19119 1492
rect 4985 776 5071 799
rect 5153 776 5239 799
rect 17157 797 17243 883
rect 20105 776 20191 799
rect 20273 776 20359 799
rect 4985 736 5010 776
rect 5010 736 5050 776
rect 5050 736 5071 776
rect 5153 736 5174 776
rect 5174 736 5214 776
rect 5214 736 5239 776
rect 20105 736 20130 776
rect 20130 736 20170 776
rect 20170 736 20191 776
rect 20273 736 20294 776
rect 20294 736 20334 776
rect 20334 736 20359 776
rect 4985 713 5071 736
rect 5153 713 5239 736
rect 20105 713 20191 736
rect 20273 713 20359 736
<< metal6 >>
rect 3652 40867 4092 43008
rect 3652 40781 3745 40867
rect 3831 40781 3913 40867
rect 3999 40781 4092 40867
rect 3652 39355 4092 40781
rect 3652 39269 3745 39355
rect 3831 39269 3913 39355
rect 3999 39269 4092 39355
rect 3652 37843 4092 39269
rect 3652 37757 3745 37843
rect 3831 37757 3913 37843
rect 3999 37757 4092 37843
rect 3652 36331 4092 37757
rect 3652 36245 3745 36331
rect 3831 36245 3913 36331
rect 3999 36245 4092 36331
rect 3652 34819 4092 36245
rect 3652 34733 3745 34819
rect 3831 34733 3913 34819
rect 3999 34733 4092 34819
rect 3652 33307 4092 34733
rect 3652 33221 3745 33307
rect 3831 33221 3913 33307
rect 3999 33221 4092 33307
rect 3652 31795 4092 33221
rect 3652 31709 3745 31795
rect 3831 31709 3913 31795
rect 3999 31709 4092 31795
rect 3652 30283 4092 31709
rect 3652 30197 3745 30283
rect 3831 30197 3913 30283
rect 3999 30197 4092 30283
rect 3652 28771 4092 30197
rect 3652 28685 3745 28771
rect 3831 28685 3913 28771
rect 3999 28685 4092 28771
rect 3652 27259 4092 28685
rect 3652 27173 3745 27259
rect 3831 27173 3913 27259
rect 3999 27173 4092 27259
rect 3652 25747 4092 27173
rect 3652 25661 3745 25747
rect 3831 25661 3913 25747
rect 3999 25661 4092 25747
rect 3652 24235 4092 25661
rect 3652 24149 3745 24235
rect 3831 24149 3913 24235
rect 3999 24149 4092 24235
rect 3652 22723 4092 24149
rect 3652 22637 3745 22723
rect 3831 22637 3913 22723
rect 3999 22637 4092 22723
rect 3652 21211 4092 22637
rect 3652 21125 3745 21211
rect 3831 21125 3913 21211
rect 3999 21125 4092 21211
rect 3652 19699 4092 21125
rect 3652 19613 3745 19699
rect 3831 19613 3913 19699
rect 3999 19613 4092 19699
rect 3652 18187 4092 19613
rect 3652 18101 3745 18187
rect 3831 18101 3913 18187
rect 3999 18101 4092 18187
rect 3652 16675 4092 18101
rect 3652 16589 3745 16675
rect 3831 16589 3913 16675
rect 3999 16589 4092 16675
rect 3652 15163 4092 16589
rect 3652 15077 3745 15163
rect 3831 15077 3913 15163
rect 3999 15077 4092 15163
rect 3652 13651 4092 15077
rect 3652 13565 3745 13651
rect 3831 13565 3913 13651
rect 3999 13565 4092 13651
rect 3652 12139 4092 13565
rect 3652 12053 3745 12139
rect 3831 12053 3913 12139
rect 3999 12053 4092 12139
rect 3652 10627 4092 12053
rect 3652 10541 3745 10627
rect 3831 10541 3913 10627
rect 3999 10541 4092 10627
rect 3652 9115 4092 10541
rect 3652 9029 3745 9115
rect 3831 9029 3913 9115
rect 3999 9029 4092 9115
rect 3652 7603 4092 9029
rect 3652 7517 3745 7603
rect 3831 7517 3913 7603
rect 3999 7517 4092 7603
rect 3652 6091 4092 7517
rect 3652 6005 3745 6091
rect 3831 6005 3913 6091
rect 3999 6005 4092 6091
rect 3652 4579 4092 6005
rect 3652 4493 3745 4579
rect 3831 4493 3913 4579
rect 3999 4493 4092 4579
rect 3652 3067 4092 4493
rect 3652 2981 3745 3067
rect 3831 2981 3913 3067
rect 3999 2981 4092 3067
rect 3652 1555 4092 2981
rect 3652 1469 3745 1555
rect 3831 1469 3913 1555
rect 3999 1469 4092 1555
rect 3652 0 4092 1469
rect 4892 41623 5332 43008
rect 4892 41537 4985 41623
rect 5071 41537 5153 41623
rect 5239 41537 5332 41623
rect 4892 40111 5332 41537
rect 18772 40867 19212 43008
rect 18772 40781 18865 40867
rect 18951 40781 19033 40867
rect 19119 40781 19212 40867
rect 4892 40025 4985 40111
rect 5071 40025 5153 40111
rect 5239 40025 5332 40111
rect 4892 38599 5332 40025
rect 4892 38513 4985 38599
rect 5071 38513 5153 38599
rect 5239 38513 5332 38599
rect 4892 37087 5332 38513
rect 4892 37001 4985 37087
rect 5071 37001 5153 37087
rect 5239 37001 5332 37087
rect 4892 35575 5332 37001
rect 4892 35489 4985 35575
rect 5071 35489 5153 35575
rect 5239 35489 5332 35575
rect 4892 34063 5332 35489
rect 4892 33977 4985 34063
rect 5071 33977 5153 34063
rect 5239 33977 5332 34063
rect 4892 32551 5332 33977
rect 4892 32465 4985 32551
rect 5071 32465 5153 32551
rect 5239 32465 5332 32551
rect 4892 31039 5332 32465
rect 4892 30953 4985 31039
rect 5071 30953 5153 31039
rect 5239 30953 5332 31039
rect 4892 29527 5332 30953
rect 4892 29441 4985 29527
rect 5071 29441 5153 29527
rect 5239 29441 5332 29527
rect 4892 28015 5332 29441
rect 4892 27929 4985 28015
rect 5071 27929 5153 28015
rect 5239 27929 5332 28015
rect 4892 26503 5332 27929
rect 4892 26417 4985 26503
rect 5071 26417 5153 26503
rect 5239 26417 5332 26503
rect 4892 24991 5332 26417
rect 4892 24905 4985 24991
rect 5071 24905 5153 24991
rect 5239 24905 5332 24991
rect 4892 23479 5332 24905
rect 4892 23393 4985 23479
rect 5071 23393 5153 23479
rect 5239 23393 5332 23479
rect 4892 21967 5332 23393
rect 4892 21881 4985 21967
rect 5071 21881 5153 21967
rect 5239 21881 5332 21967
rect 4892 20455 5332 21881
rect 4892 20369 4985 20455
rect 5071 20369 5153 20455
rect 5239 20369 5332 20455
rect 4892 18943 5332 20369
rect 4892 18857 4985 18943
rect 5071 18857 5153 18943
rect 5239 18857 5332 18943
rect 4892 17431 5332 18857
rect 4892 17345 4985 17431
rect 5071 17345 5153 17431
rect 5239 17345 5332 17431
rect 4892 15919 5332 17345
rect 4892 15833 4985 15919
rect 5071 15833 5153 15919
rect 5239 15833 5332 15919
rect 4892 14407 5332 15833
rect 4892 14321 4985 14407
rect 5071 14321 5153 14407
rect 5239 14321 5332 14407
rect 4892 12895 5332 14321
rect 4892 12809 4985 12895
rect 5071 12809 5153 12895
rect 5239 12809 5332 12895
rect 4892 11383 5332 12809
rect 4892 11297 4985 11383
rect 5071 11297 5153 11383
rect 5239 11297 5332 11383
rect 4892 9871 5332 11297
rect 4892 9785 4985 9871
rect 5071 9785 5153 9871
rect 5239 9785 5332 9871
rect 4892 8359 5332 9785
rect 4892 8273 4985 8359
rect 5071 8273 5153 8359
rect 5239 8273 5332 8359
rect 4892 6847 5332 8273
rect 4892 6761 4985 6847
rect 5071 6761 5153 6847
rect 5239 6761 5332 6847
rect 4892 5335 5332 6761
rect 12020 40531 12348 40652
rect 12020 40445 12141 40531
rect 12227 40445 12348 40531
rect 12020 5839 12348 40445
rect 12020 5753 12141 5839
rect 12227 5753 12348 5839
rect 12020 5632 12348 5753
rect 17036 39859 17364 39980
rect 17036 39773 17157 39859
rect 17243 39773 17364 39859
rect 4892 5249 4985 5335
rect 5071 5249 5153 5335
rect 5239 5249 5332 5335
rect 4892 3823 5332 5249
rect 4892 3737 4985 3823
rect 5071 3737 5153 3823
rect 5239 3737 5332 3823
rect 4892 2311 5332 3737
rect 4892 2225 4985 2311
rect 5071 2225 5153 2311
rect 5239 2225 5332 2311
rect 4892 799 5332 2225
rect 4892 713 4985 799
rect 5071 713 5153 799
rect 5239 713 5332 799
rect 4892 0 5332 713
rect 17036 883 17364 39773
rect 17036 797 17157 883
rect 17243 797 17364 883
rect 17036 676 17364 797
rect 18772 39355 19212 40781
rect 18772 39269 18865 39355
rect 18951 39269 19033 39355
rect 19119 39269 19212 39355
rect 18772 37843 19212 39269
rect 18772 37757 18865 37843
rect 18951 37757 19033 37843
rect 19119 37757 19212 37843
rect 18772 36331 19212 37757
rect 18772 36245 18865 36331
rect 18951 36245 19033 36331
rect 19119 36245 19212 36331
rect 18772 34819 19212 36245
rect 18772 34733 18865 34819
rect 18951 34733 19033 34819
rect 19119 34733 19212 34819
rect 18772 33307 19212 34733
rect 18772 33221 18865 33307
rect 18951 33221 19033 33307
rect 19119 33221 19212 33307
rect 18772 31795 19212 33221
rect 18772 31709 18865 31795
rect 18951 31709 19033 31795
rect 19119 31709 19212 31795
rect 18772 30283 19212 31709
rect 18772 30197 18865 30283
rect 18951 30197 19033 30283
rect 19119 30197 19212 30283
rect 18772 28771 19212 30197
rect 18772 28685 18865 28771
rect 18951 28685 19033 28771
rect 19119 28685 19212 28771
rect 18772 27259 19212 28685
rect 18772 27173 18865 27259
rect 18951 27173 19033 27259
rect 19119 27173 19212 27259
rect 18772 25747 19212 27173
rect 18772 25661 18865 25747
rect 18951 25661 19033 25747
rect 19119 25661 19212 25747
rect 18772 24235 19212 25661
rect 18772 24149 18865 24235
rect 18951 24149 19033 24235
rect 19119 24149 19212 24235
rect 18772 22723 19212 24149
rect 18772 22637 18865 22723
rect 18951 22637 19033 22723
rect 19119 22637 19212 22723
rect 18772 21211 19212 22637
rect 18772 21125 18865 21211
rect 18951 21125 19033 21211
rect 19119 21125 19212 21211
rect 18772 19699 19212 21125
rect 18772 19613 18865 19699
rect 18951 19613 19033 19699
rect 19119 19613 19212 19699
rect 18772 18187 19212 19613
rect 18772 18101 18865 18187
rect 18951 18101 19033 18187
rect 19119 18101 19212 18187
rect 18772 16675 19212 18101
rect 18772 16589 18865 16675
rect 18951 16589 19033 16675
rect 19119 16589 19212 16675
rect 18772 15163 19212 16589
rect 18772 15077 18865 15163
rect 18951 15077 19033 15163
rect 19119 15077 19212 15163
rect 18772 13651 19212 15077
rect 18772 13565 18865 13651
rect 18951 13565 19033 13651
rect 19119 13565 19212 13651
rect 18772 12139 19212 13565
rect 18772 12053 18865 12139
rect 18951 12053 19033 12139
rect 19119 12053 19212 12139
rect 18772 10627 19212 12053
rect 18772 10541 18865 10627
rect 18951 10541 19033 10627
rect 19119 10541 19212 10627
rect 18772 9115 19212 10541
rect 18772 9029 18865 9115
rect 18951 9029 19033 9115
rect 19119 9029 19212 9115
rect 18772 7603 19212 9029
rect 18772 7517 18865 7603
rect 18951 7517 19033 7603
rect 19119 7517 19212 7603
rect 18772 6091 19212 7517
rect 18772 6005 18865 6091
rect 18951 6005 19033 6091
rect 19119 6005 19212 6091
rect 18772 4579 19212 6005
rect 18772 4493 18865 4579
rect 18951 4493 19033 4579
rect 19119 4493 19212 4579
rect 18772 3067 19212 4493
rect 18772 2981 18865 3067
rect 18951 2981 19033 3067
rect 19119 2981 19212 3067
rect 18772 1555 19212 2981
rect 18772 1469 18865 1555
rect 18951 1469 19033 1555
rect 19119 1469 19212 1555
rect 18772 0 19212 1469
rect 20012 41623 20452 43008
rect 20012 41537 20105 41623
rect 20191 41537 20273 41623
rect 20359 41537 20452 41623
rect 20012 40111 20452 41537
rect 20012 40025 20105 40111
rect 20191 40025 20273 40111
rect 20359 40025 20452 40111
rect 20012 38599 20452 40025
rect 20012 38513 20105 38599
rect 20191 38513 20273 38599
rect 20359 38513 20452 38599
rect 20012 37087 20452 38513
rect 20012 37001 20105 37087
rect 20191 37001 20273 37087
rect 20359 37001 20452 37087
rect 20012 35575 20452 37001
rect 20012 35489 20105 35575
rect 20191 35489 20273 35575
rect 20359 35489 20452 35575
rect 20012 34063 20452 35489
rect 20012 33977 20105 34063
rect 20191 33977 20273 34063
rect 20359 33977 20452 34063
rect 20012 32551 20452 33977
rect 20012 32465 20105 32551
rect 20191 32465 20273 32551
rect 20359 32465 20452 32551
rect 20012 31039 20452 32465
rect 20012 30953 20105 31039
rect 20191 30953 20273 31039
rect 20359 30953 20452 31039
rect 20012 29527 20452 30953
rect 20012 29441 20105 29527
rect 20191 29441 20273 29527
rect 20359 29441 20452 29527
rect 20012 28015 20452 29441
rect 20012 27929 20105 28015
rect 20191 27929 20273 28015
rect 20359 27929 20452 28015
rect 20012 26503 20452 27929
rect 20012 26417 20105 26503
rect 20191 26417 20273 26503
rect 20359 26417 20452 26503
rect 20012 24991 20452 26417
rect 20012 24905 20105 24991
rect 20191 24905 20273 24991
rect 20359 24905 20452 24991
rect 20012 23479 20452 24905
rect 20012 23393 20105 23479
rect 20191 23393 20273 23479
rect 20359 23393 20452 23479
rect 20012 21967 20452 23393
rect 20012 21881 20105 21967
rect 20191 21881 20273 21967
rect 20359 21881 20452 21967
rect 20012 20455 20452 21881
rect 20012 20369 20105 20455
rect 20191 20369 20273 20455
rect 20359 20369 20452 20455
rect 20012 18943 20452 20369
rect 20012 18857 20105 18943
rect 20191 18857 20273 18943
rect 20359 18857 20452 18943
rect 20012 17431 20452 18857
rect 20012 17345 20105 17431
rect 20191 17345 20273 17431
rect 20359 17345 20452 17431
rect 20012 15919 20452 17345
rect 20012 15833 20105 15919
rect 20191 15833 20273 15919
rect 20359 15833 20452 15919
rect 20012 14407 20452 15833
rect 20012 14321 20105 14407
rect 20191 14321 20273 14407
rect 20359 14321 20452 14407
rect 20012 12895 20452 14321
rect 20012 12809 20105 12895
rect 20191 12809 20273 12895
rect 20359 12809 20452 12895
rect 20012 11383 20452 12809
rect 20012 11297 20105 11383
rect 20191 11297 20273 11383
rect 20359 11297 20452 11383
rect 20012 9871 20452 11297
rect 20012 9785 20105 9871
rect 20191 9785 20273 9871
rect 20359 9785 20452 9871
rect 20012 8359 20452 9785
rect 20012 8273 20105 8359
rect 20191 8273 20273 8359
rect 20359 8273 20452 8359
rect 20012 6847 20452 8273
rect 20012 6761 20105 6847
rect 20191 6761 20273 6847
rect 20359 6761 20452 6847
rect 20012 5335 20452 6761
rect 20012 5249 20105 5335
rect 20191 5249 20273 5335
rect 20359 5249 20452 5335
rect 20012 3823 20452 5249
rect 20012 3737 20105 3823
rect 20191 3737 20273 3823
rect 20359 3737 20452 3823
rect 20012 2311 20452 3737
rect 20012 2225 20105 2311
rect 20191 2225 20273 2311
rect 20359 2225 20452 2311
rect 20012 799 20452 2225
rect 20012 713 20105 799
rect 20191 713 20273 799
rect 20359 713 20452 799
rect 20012 0 20452 713
use sg13g2_inv_1  _209_
timestamp 1676382929
transform 1 0 7008 0 -1 6804
box -48 -56 336 834
use sg13g2_inv_1  _210_
timestamp 1676382929
transform -1 0 6432 0 1 756
box -48 -56 336 834
use sg13g2_inv_1  _211_
timestamp 1676382929
transform 1 0 12384 0 -1 21924
box -48 -56 336 834
use sg13g2_inv_1  _212_
timestamp 1676382929
transform -1 0 7584 0 -1 18900
box -48 -56 336 834
use sg13g2_inv_1  _213_
timestamp 1676382929
transform 1 0 2976 0 1 30996
box -48 -56 336 834
use sg13g2_inv_1  _214_
timestamp 1676382929
transform 1 0 14784 0 -1 9828
box -48 -56 336 834
use sg13g2_inv_1  _215_
timestamp 1676382929
transform 1 0 7296 0 -1 30996
box -48 -56 336 834
use sg13g2_inv_1  _216_
timestamp 1676382929
transform 1 0 18432 0 -1 8316
box -48 -56 336 834
use sg13g2_inv_1  _217_
timestamp 1676382929
transform 1 0 19968 0 1 11340
box -48 -56 336 834
use sg13g2_inv_1  _218_
timestamp 1676382929
transform -1 0 14880 0 1 12852
box -48 -56 336 834
use sg13g2_inv_1  _219_
timestamp 1676382929
transform -1 0 15744 0 -1 12852
box -48 -56 336 834
use sg13g2_inv_1  _220_
timestamp 1676382929
transform 1 0 17568 0 1 756
box -48 -56 336 834
use sg13g2_inv_1  _221_
timestamp 1676382929
transform -1 0 18240 0 -1 2268
box -48 -56 336 834
use sg13g2_inv_1  _222_
timestamp 1676382929
transform 1 0 13632 0 1 17388
box -48 -56 336 834
use sg13g2_inv_1  _223_
timestamp 1676382929
transform -1 0 14016 0 1 18900
box -48 -56 336 834
use sg13g2_inv_1  _224_
timestamp 1676382929
transform -1 0 6144 0 1 34020
box -48 -56 336 834
use sg13g2_inv_1  _225_
timestamp 1676382929
transform 1 0 7680 0 1 32508
box -48 -56 336 834
use sg13g2_inv_1  _226_
timestamp 1676382929
transform -1 0 4320 0 1 30996
box -48 -56 336 834
use sg13g2_inv_1  _227_
timestamp 1676382929
transform -1 0 16800 0 1 3780
box -48 -56 336 834
use sg13g2_inv_1  _228_
timestamp 1676382929
transform -1 0 16512 0 1 3780
box -48 -56 336 834
use sg13g2_mux2_1  _229_
timestamp 1677247768
transform -1 0 6720 0 1 2268
box -48 -56 1008 834
use sg13g2_nand2_1  _230_
timestamp 1676557249
transform 1 0 1536 0 1 2268
box -48 -56 432 834
use sg13g2_mux2_1  _231_
timestamp 1677247768
transform -1 0 8544 0 1 2268
box -48 -56 1008 834
use sg13g2_a21oi_1  _232_
timestamp 1683973020
transform 1 0 6912 0 -1 2268
box -48 -56 528 834
use sg13g2_mux2_1  _233_
timestamp 1677247768
transform 1 0 5184 0 1 756
box -48 -56 1008 834
use sg13g2_nand2b_1  _234_
timestamp 1676567195
transform -1 0 7584 0 1 756
box -48 -56 528 834
use sg13g2_o21ai_1  _235_
timestamp 1685175443
transform 1 0 4704 0 1 756
box -48 -56 538 834
use sg13g2_nand2b_1  _236_
timestamp 1676567195
transform 1 0 6432 0 1 756
box -48 -56 528 834
use sg13g2_a21oi_1  _237_
timestamp 1683973020
transform -1 0 8544 0 -1 2268
box -48 -56 528 834
use sg13g2_a221oi_1  _238_
timestamp 1685197497
transform 1 0 6720 0 1 2268
box -48 -56 816 834
use sg13g2_nor2_1  _239_
timestamp 1676627187
transform -1 0 9792 0 1 2268
box -48 -56 432 834
use sg13g2_nor2b_1  _240_
timestamp 1685181386
transform -1 0 10176 0 -1 2268
box -54 -56 528 834
use sg13g2_nor2b_1  _241_
timestamp 1685181386
transform -1 0 9120 0 1 2268
box -54 -56 528 834
use sg13g2_a22oi_1  _242_
timestamp 1685173987
transform 1 0 7968 0 -1 3780
box -48 -56 624 834
use sg13g2_a21oi_1  _243_
timestamp 1683973020
transform 1 0 6912 0 -1 3780
box -48 -56 528 834
use sg13g2_o21ai_1  _244_
timestamp 1685175443
transform 1 0 7584 0 -1 2268
box -48 -56 538 834
use sg13g2_a22oi_1  _245_
timestamp 1685173987
transform 1 0 8544 0 -1 3780
box -48 -56 624 834
use sg13g2_and2_1  _246_
timestamp 1676901763
transform 1 0 8544 0 -1 2268
box -48 -56 528 834
use sg13g2_a22oi_1  _247_
timestamp 1685173987
transform -1 0 7968 0 -1 3780
box -48 -56 624 834
use sg13g2_a21o_1  _248_
timestamp 1677175127
transform 1 0 4512 0 -1 3780
box -48 -56 720 834
use sg13g2_mux4_1  _249_
timestamp 1677257233
transform 1 0 10848 0 -1 40068
box -48 -56 2064 834
use sg13g2_inv_1  _250_
timestamp 1676382929
transform -1 0 17856 0 -1 12852
box -48 -56 336 834
use sg13g2_mux4_1  _251_
timestamp 1677257233
transform 1 0 12288 0 -1 34020
box -48 -56 2064 834
use sg13g2_nor2b_1  _252_
timestamp 1685181386
transform -1 0 13824 0 -1 11340
box -54 -56 528 834
use sg13g2_a21oi_1  _253_
timestamp 1683973020
transform 1 0 13728 0 1 11340
box -48 -56 528 834
use sg13g2_nand3b_1  _254_
timestamp 1676573470
transform 1 0 12768 0 -1 12852
box -48 -56 720 834
use sg13g2_o21ai_1  _255_
timestamp 1685175443
transform 1 0 14208 0 1 11340
box -48 -56 538 834
use sg13g2_mux4_1  _256_
timestamp 1677257233
transform 1 0 11712 0 1 11340
box -48 -56 2064 834
use sg13g2_mux2_1  _257_
timestamp 1677247768
transform -1 0 13344 0 -1 11340
box -48 -56 1008 834
use sg13g2_mux4_1  _258_
timestamp 1677257233
transform 1 0 9984 0 1 40068
box -48 -56 2064 834
use sg13g2_mux4_1  _259_
timestamp 1677257233
transform 1 0 7776 0 1 34020
box -48 -56 2064 834
use sg13g2_nor2b_1  _260_
timestamp 1685181386
transform -1 0 4896 0 1 8316
box -54 -56 528 834
use sg13g2_a21oi_1  _261_
timestamp 1683973020
transform -1 0 4416 0 1 8316
box -48 -56 528 834
use sg13g2_nand3b_1  _262_
timestamp 1676573470
transform 1 0 1824 0 -1 8316
box -48 -56 720 834
use sg13g2_o21ai_1  _263_
timestamp 1685175443
transform 1 0 2880 0 -1 6804
box -48 -56 538 834
use sg13g2_mux4_1  _264_
timestamp 1677257233
transform 1 0 2496 0 -1 8316
box -48 -56 2064 834
use sg13g2_mux2_1  _265_
timestamp 1677247768
transform -1 0 3936 0 1 8316
box -48 -56 1008 834
use sg13g2_mux4_1  _266_
timestamp 1677257233
transform 1 0 1728 0 -1 34020
box -48 -56 2064 834
use sg13g2_mux4_1  _267_
timestamp 1677257233
transform 1 0 4608 0 -1 38556
box -48 -56 2064 834
use sg13g2_mux4_1  _268_
timestamp 1677257233
transform 1 0 3072 0 -1 23436
box -48 -56 2064 834
use sg13g2_nand3b_1  _269_
timestamp 1676573470
transform 1 0 4320 0 1 23436
box -48 -56 720 834
use sg13g2_nor2b_1  _270_
timestamp 1685181386
transform -1 0 6048 0 -1 23436
box -54 -56 528 834
use sg13g2_a21oi_1  _271_
timestamp 1683973020
transform -1 0 5472 0 1 23436
box -48 -56 528 834
use sg13g2_o21ai_1  _272_
timestamp 1685175443
transform 1 0 5088 0 -1 23436
box -48 -56 538 834
use sg13g2_mux2_1  _273_
timestamp 1677247768
transform -1 0 5568 0 1 21924
box -48 -56 1008 834
use sg13g2_mux4_1  _274_
timestamp 1677257233
transform 1 0 12288 0 -1 32508
box -48 -56 2064 834
use sg13g2_mux4_1  _275_
timestamp 1677257233
transform 1 0 9792 0 -1 38556
box -48 -56 2064 834
use sg13g2_inv_1  _276_
timestamp 1676382929
transform -1 0 17568 0 1 756
box -48 -56 336 834
use sg13g2_nor2b_1  _277_
timestamp 1685181386
transform 1 0 17952 0 -1 8316
box -54 -56 528 834
use sg13g2_a21oi_1  _278_
timestamp 1683973020
transform -1 0 18720 0 -1 5292
box -48 -56 528 834
use sg13g2_nand3b_1  _279_
timestamp 1676573470
transform 1 0 17472 0 -1 6804
box -48 -56 720 834
use sg13g2_o21ai_1  _280_
timestamp 1685175443
transform 1 0 19872 0 1 5292
box -48 -56 538 834
use sg13g2_mux4_1  _281_
timestamp 1677257233
transform 1 0 18144 0 -1 6804
box -48 -56 2064 834
use sg13g2_mux2_1  _282_
timestamp 1677247768
transform -1 0 19968 0 -1 8316
box -48 -56 1008 834
use sg13g2_mux4_1  _283_
timestamp 1677257233
transform 1 0 13152 0 1 34020
box -48 -56 2064 834
use sg13g2_mux4_1  _284_
timestamp 1677257233
transform 1 0 5184 0 1 3780
box -48 -56 2064 834
use sg13g2_nand3b_1  _285_
timestamp 1676573470
transform 1 0 16320 0 1 15876
box -48 -56 720 834
use sg13g2_nor2b_1  _286_
timestamp 1685181386
transform -1 0 16320 0 1 15876
box -54 -56 528 834
use sg13g2_a21oi_1  _287_
timestamp 1683973020
transform -1 0 15840 0 1 15876
box -48 -56 528 834
use sg13g2_o21ai_1  _288_
timestamp 1685175443
transform -1 0 17952 0 -1 17388
box -48 -56 538 834
use sg13g2_mux4_1  _289_
timestamp 1677257233
transform 1 0 16032 0 -1 15876
box -48 -56 2064 834
use sg13g2_mux2_1  _290_
timestamp 1677247768
transform -1 0 17952 0 1 15876
box -48 -56 1008 834
use sg13g2_mux4_1  _291_
timestamp 1677257233
transform 1 0 7680 0 1 38556
box -48 -56 2064 834
use sg13g2_mux4_1  _292_
timestamp 1677257233
transform 1 0 4992 0 -1 6804
box -48 -56 2064 834
use sg13g2_mux4_1  _293_
timestamp 1677257233
transform -1 0 9696 0 -1 11340
box -48 -56 2064 834
use sg13g2_nand3b_1  _294_
timestamp 1676573470
transform -1 0 8544 0 1 9828
box -48 -56 720 834
use sg13g2_nor2b_1  _295_
timestamp 1685181386
transform -1 0 9120 0 1 11340
box -54 -56 528 834
use sg13g2_a21oi_1  _296_
timestamp 1683973020
transform -1 0 8832 0 -1 14364
box -48 -56 528 834
use sg13g2_o21ai_1  _297_
timestamp 1685175443
transform -1 0 7872 0 1 9828
box -48 -56 538 834
use sg13g2_mux2_1  _298_
timestamp 1677247768
transform -1 0 8544 0 -1 12852
box -48 -56 1008 834
use sg13g2_mux4_1  _299_
timestamp 1677257233
transform 1 0 2304 0 1 37044
box -48 -56 2064 834
use sg13g2_mux4_1  _300_
timestamp 1677257233
transform 1 0 3744 0 -1 35532
box -48 -56 2064 834
use sg13g2_nor2b_1  _301_
timestamp 1685181386
transform -1 0 4800 0 -1 11340
box -54 -56 528 834
use sg13g2_a21oi_1  _302_
timestamp 1683973020
transform 1 0 4800 0 -1 11340
box -48 -56 528 834
use sg13g2_nand3b_1  _303_
timestamp 1676573470
transform 1 0 3168 0 -1 9828
box -48 -56 720 834
use sg13g2_o21ai_1  _304_
timestamp 1685175443
transform -1 0 3936 0 1 11340
box -48 -56 538 834
use sg13g2_mux4_1  _305_
timestamp 1677257233
transform -1 0 4800 0 1 9828
box -48 -56 2064 834
use sg13g2_mux2_1  _306_
timestamp 1677247768
transform -1 0 3936 0 -1 11340
box -48 -56 1008 834
use sg13g2_mux4_1  _307_
timestamp 1677257233
transform 1 0 9312 0 1 35532
box -48 -56 2064 834
use sg13g2_inv_1  _308_
timestamp 1676382929
transform 1 0 16320 0 1 6804
box -48 -56 336 834
use sg13g2_mux4_1  _309_
timestamp 1677257233
transform 1 0 14784 0 1 38556
box -48 -56 2064 834
use sg13g2_inv_1  _310_
timestamp 1676382929
transform -1 0 17856 0 -1 5292
box -48 -56 336 834
use sg13g2_nand3_1  _311_
timestamp 1683988354
transform -1 0 20352 0 -1 9828
box -48 -56 528 834
use sg13g2_or2_1  _312_
timestamp 1684236171
transform -1 0 17856 0 -1 9828
box -48 -56 528 834
use sg13g2_o21ai_1  _313_
timestamp 1685175443
transform -1 0 17376 0 -1 9828
box -48 -56 538 834
use sg13g2_o21ai_1  _314_
timestamp 1685175443
transform 1 0 19392 0 1 8316
box -48 -56 538 834
use sg13g2_mux4_1  _315_
timestamp 1677257233
transform 1 0 17856 0 -1 9828
box -48 -56 2064 834
use sg13g2_mux2_1  _316_
timestamp 1677247768
transform -1 0 19968 0 1 9828
box -48 -56 1008 834
use sg13g2_mux4_1  _317_
timestamp 1677257233
transform 1 0 12288 0 -1 37044
box -48 -56 2064 834
use sg13g2_mux4_1  _318_
timestamp 1677257233
transform 1 0 12480 0 1 12852
box -48 -56 2064 834
use sg13g2_nand3b_1  _319_
timestamp 1676573470
transform 1 0 13056 0 1 14364
box -48 -56 720 834
use sg13g2_nor2b_1  _320_
timestamp 1685181386
transform -1 0 14880 0 -1 14364
box -54 -56 528 834
use sg13g2_a21oi_1  _321_
timestamp 1683973020
transform -1 0 13056 0 1 14364
box -48 -56 528 834
use sg13g2_o21ai_1  _322_
timestamp 1685175443
transform 1 0 14688 0 1 14364
box -48 -56 538 834
use sg13g2_mux2_1  _323_
timestamp 1677247768
transform -1 0 14688 0 1 14364
box -48 -56 1008 834
use sg13g2_mux4_1  _324_
timestamp 1677257233
transform 1 0 5664 0 1 38556
box -48 -56 2064 834
use sg13g2_mux4_1  _325_
timestamp 1677257233
transform -1 0 4416 0 1 5292
box -48 -56 2064 834
use sg13g2_nand3b_1  _326_
timestamp 1676573470
transform 1 0 4416 0 1 5292
box -48 -56 720 834
use sg13g2_nor2b_1  _327_
timestamp 1685181386
transform -1 0 4896 0 -1 5292
box -54 -56 528 834
use sg13g2_a21oi_1  _328_
timestamp 1683973020
transform -1 0 3264 0 1 3780
box -48 -56 528 834
use sg13g2_o21ai_1  _329_
timestamp 1685175443
transform 1 0 4416 0 1 6804
box -48 -56 538 834
use sg13g2_mux2_1  _330_
timestamp 1677247768
transform -1 0 2400 0 1 5292
box -48 -56 1008 834
use sg13g2_mux4_1  _331_
timestamp 1677257233
transform 1 0 2304 0 -1 38556
box -48 -56 2064 834
use sg13g2_nor2b_1  _332_
timestamp 1685181386
transform -1 0 3648 0 -1 20412
box -54 -56 528 834
use sg13g2_a21oi_1  _333_
timestamp 1683973020
transform 1 0 4320 0 -1 20412
box -48 -56 528 834
use sg13g2_nand3b_1  _334_
timestamp 1676573470
transform -1 0 4320 0 -1 20412
box -48 -56 720 834
use sg13g2_o21ai_1  _335_
timestamp 1685175443
transform -1 0 4032 0 1 18900
box -48 -56 538 834
use sg13g2_mux4_1  _336_
timestamp 1677257233
transform -1 0 5376 0 1 20412
box -48 -56 2064 834
use sg13g2_mux2_1  _337_
timestamp 1677247768
transform -1 0 3840 0 -1 21924
box -48 -56 1008 834
use sg13g2_mux4_1  _338_
timestamp 1677257233
transform 1 0 15168 0 -1 38556
box -48 -56 2064 834
use sg13g2_nor2b_1  _339_
timestamp 1685181386
transform 1 0 19680 0 -1 3780
box -54 -56 528 834
use sg13g2_a21oi_1  _340_
timestamp 1683973020
transform -1 0 20064 0 1 2268
box -48 -56 528 834
use sg13g2_nand3b_1  _341_
timestamp 1676573470
transform -1 0 19584 0 1 2268
box -48 -56 720 834
use sg13g2_o21ai_1  _342_
timestamp 1685175443
transform 1 0 18432 0 1 2268
box -48 -56 538 834
use sg13g2_mux4_1  _343_
timestamp 1677257233
transform 1 0 18336 0 1 3780
box -48 -56 2064 834
use sg13g2_mux2_1  _344_
timestamp 1677247768
transform -1 0 19968 0 -1 5292
box -48 -56 1008 834
use sg13g2_mux4_1  _345_
timestamp 1677257233
transform 1 0 12960 0 1 35532
box -48 -56 2064 834
use sg13g2_mux4_1  _346_
timestamp 1677257233
transform 1 0 18336 0 -1 15876
box -48 -56 2064 834
use sg13g2_nand3b_1  _347_
timestamp 1676573470
transform 1 0 19200 0 1 14364
box -48 -56 720 834
use sg13g2_nor2b_1  _348_
timestamp 1685181386
transform 1 0 18144 0 -1 14364
box -54 -56 528 834
use sg13g2_a21oi_1  _349_
timestamp 1683973020
transform 1 0 19872 0 1 14364
box -48 -56 528 834
use sg13g2_o21ai_1  _350_
timestamp 1685175443
transform -1 0 20256 0 1 15876
box -48 -56 538 834
use sg13g2_mux2_1  _351_
timestamp 1677247768
transform -1 0 19968 0 1 17388
box -48 -56 1008 834
use sg13g2_mux4_1  _352_
timestamp 1677257233
transform 1 0 7488 0 1 37044
box -48 -56 2064 834
use sg13g2_mux4_1  _353_
timestamp 1677257233
transform 1 0 8544 0 1 9828
box -48 -56 2064 834
use sg13g2_nand3b_1  _354_
timestamp 1676573470
transform -1 0 10272 0 -1 9828
box -48 -56 720 834
use sg13g2_nor2b_1  _355_
timestamp 1685181386
transform 1 0 10272 0 -1 9828
box -54 -56 528 834
use sg13g2_a21oi_1  _356_
timestamp 1683973020
transform 1 0 10560 0 1 9828
box -48 -56 528 834
use sg13g2_o21ai_1  _357_
timestamp 1685175443
transform -1 0 10176 0 -1 11340
box -48 -56 538 834
use sg13g2_mux2_1  _358_
timestamp 1677247768
transform -1 0 10080 0 1 11340
box -48 -56 1008 834
use sg13g2_mux4_1  _359_
timestamp 1677257233
transform 1 0 1728 0 -1 35532
box -48 -56 2064 834
use sg13g2_nor2b_1  _360_
timestamp 1685181386
transform 1 0 2976 0 -1 17388
box -54 -56 528 834
use sg13g2_a21oi_1  _361_
timestamp 1683973020
transform 1 0 3552 0 -1 15876
box -48 -56 528 834
use sg13g2_nand3b_1  _362_
timestamp 1676573470
transform 1 0 2880 0 -1 15876
box -48 -56 720 834
use sg13g2_o21ai_1  _363_
timestamp 1685175443
transform -1 0 4224 0 1 14364
box -48 -56 538 834
use sg13g2_mux4_1  _364_
timestamp 1677257233
transform -1 0 4608 0 -1 14364
box -48 -56 2064 834
use sg13g2_mux2_1  _365_
timestamp 1677247768
transform -1 0 3744 0 1 14364
box -48 -56 1008 834
use sg13g2_mux4_1  _366_
timestamp 1677257233
transform 1 0 15168 0 -1 37044
box -48 -56 2064 834
use sg13g2_nand3_1  _367_
timestamp 1683988354
transform 1 0 17664 0 -1 11340
box -48 -56 528 834
use sg13g2_or2_1  _368_
timestamp 1684236171
transform -1 0 18912 0 1 11340
box -48 -56 528 834
use sg13g2_o21ai_1  _369_
timestamp 1685175443
transform 1 0 17856 0 -1 12852
box -48 -56 538 834
use sg13g2_o21ai_1  _370_
timestamp 1685175443
transform -1 0 19872 0 1 12852
box -48 -56 538 834
use sg13g2_mux4_1  _371_
timestamp 1677257233
transform 1 0 18144 0 -1 11340
box -48 -56 2064 834
use sg13g2_mux2_1  _372_
timestamp 1677247768
transform -1 0 19968 0 1 11340
box -48 -56 1008 834
use sg13g2_o21ai_1  _373_
timestamp 1685175443
transform 1 0 16512 0 -1 14364
box -48 -56 538 834
use sg13g2_a21o_1  _374_
timestamp 1677175127
transform 1 0 16896 0 1 12852
box -48 -56 720 834
use sg13g2_mux2_1  _375_
timestamp 1677247768
transform 1 0 16224 0 -1 12852
box -48 -56 1008 834
use sg13g2_a21oi_1  _376_
timestamp 1683973020
transform 1 0 16992 0 -1 14364
box -48 -56 528 834
use sg13g2_mux4_1  _377_
timestamp 1677257233
transform 1 0 14880 0 1 12852
box -48 -56 2064 834
use sg13g2_nor2_1  _378_
timestamp 1676627187
transform -1 0 17568 0 -1 12852
box -48 -56 432 834
use sg13g2_a21oi_1  _379_
timestamp 1683973020
transform -1 0 16224 0 -1 12852
box -48 -56 528 834
use sg13g2_mux4_1  _380_
timestamp 1677257233
transform 1 0 8544 0 1 5292
box -48 -56 2064 834
use sg13g2_mux4_1  _381_
timestamp 1677257233
transform 1 0 8544 0 -1 6804
box -48 -56 2064 834
use sg13g2_mux2_1  _382_
timestamp 1677247768
transform 1 0 9792 0 1 2268
box -48 -56 1008 834
use sg13g2_mux4_1  _383_
timestamp 1677257233
transform 1 0 6432 0 -1 23436
box -48 -56 2064 834
use sg13g2_nand2b_1  _384_
timestamp 1676567195
transform -1 0 9408 0 -1 23436
box -48 -56 528 834
use sg13g2_mux2_1  _385_
timestamp 1677247768
transform 1 0 7008 0 -1 24948
box -48 -56 1008 834
use sg13g2_nand2b_1  _386_
timestamp 1676567195
transform 1 0 6912 0 1 21924
box -48 -56 528 834
use sg13g2_nand2_1  _387_
timestamp 1676557249
transform 1 0 6048 0 -1 23436
box -48 -56 432 834
use sg13g2_and3_1  _388_
timestamp 1676971669
transform 1 0 7392 0 1 21924
box -48 -56 720 834
use sg13g2_o21ai_1  _389_
timestamp 1685175443
transform 1 0 9408 0 -1 23436
box -48 -56 538 834
use sg13g2_o21ai_1  _390_
timestamp 1685175443
transform 1 0 8448 0 -1 23436
box -48 -56 538 834
use sg13g2_o21ai_1  _391_
timestamp 1685175443
transform -1 0 16800 0 1 2268
box -48 -56 538 834
use sg13g2_a21o_1  _392_
timestamp 1677175127
transform 1 0 16800 0 -1 2268
box -48 -56 720 834
use sg13g2_mux2_1  _393_
timestamp 1677247768
transform 1 0 16800 0 1 3780
box -48 -56 1008 834
use sg13g2_a21oi_1  _394_
timestamp 1683973020
transform -1 0 17952 0 -1 2268
box -48 -56 528 834
use sg13g2_o21ai_1  _395_
timestamp 1685175443
transform -1 0 17856 0 -1 3780
box -48 -56 538 834
use sg13g2_a21o_1  _396_
timestamp 1677175127
transform 1 0 16704 0 -1 3780
box -48 -56 720 834
use sg13g2_mux2_1  _397_
timestamp 1677247768
transform 1 0 16800 0 1 2268
box -48 -56 1008 834
use sg13g2_a21oi_1  _398_
timestamp 1683973020
transform -1 0 18240 0 1 2268
box -48 -56 528 834
use sg13g2_a22oi_1  _399_
timestamp 1685173987
transform 1 0 16128 0 -1 3780
box -48 -56 624 834
use sg13g2_mux4_1  _400_
timestamp 1677257233
transform -1 0 15936 0 1 17388
box -48 -56 2064 834
use sg13g2_nand2b_1  _401_
timestamp 1676567195
transform 1 0 15072 0 -1 20412
box -48 -56 528 834
use sg13g2_a21oi_1  _402_
timestamp 1683973020
transform 1 0 15264 0 -1 17388
box -48 -56 528 834
use sg13g2_nand2b_1  _403_
timestamp 1676567195
transform -1 0 14496 0 1 18900
box -48 -56 528 834
use sg13g2_a21oi_1  _404_
timestamp 1683973020
transform 1 0 15936 0 1 17388
box -48 -56 528 834
use sg13g2_a221oi_1  _405_
timestamp 1685197497
transform 1 0 15072 0 -1 18900
box -48 -56 816 834
use sg13g2_a21o_1  _406_
timestamp 1677175127
transform -1 0 15168 0 1 18900
box -48 -56 720 834
use sg13g2_mux4_1  _407_
timestamp 1677257233
transform 1 0 7872 0 1 14364
box -48 -56 2064 834
use sg13g2_mux4_1  _408_
timestamp 1677257233
transform 1 0 7776 0 -1 15876
box -48 -56 2064 834
use sg13g2_mux2_1  _409_
timestamp 1677247768
transform -1 0 9792 0 -1 14364
box -48 -56 1008 834
use sg13g2_nor2_1  _410_
timestamp 1676627187
transform 1 0 6912 0 -1 30996
box -48 -56 432 834
use sg13g2_o21ai_1  _411_
timestamp 1685175443
transform 1 0 6240 0 -1 30996
box -48 -56 538 834
use sg13g2_or2_1  _412_
timestamp 1684236171
transform 1 0 7488 0 -1 32508
box -48 -56 528 834
use sg13g2_mux2_1  _413_
timestamp 1677247768
transform 1 0 6336 0 -1 32508
box -48 -56 1008 834
use sg13g2_a21oi_1  _414_
timestamp 1683973020
transform -1 0 7200 0 1 32508
box -48 -56 528 834
use sg13g2_a21oi_1  _415_
timestamp 1683973020
transform 1 0 7200 0 1 32508
box -48 -56 528 834
use sg13g2_o21ai_1  _416_
timestamp 1685175443
transform 1 0 7968 0 -1 32508
box -48 -56 538 834
use sg13g2_mux2_1  _417_
timestamp 1677247768
transform -1 0 6720 0 1 32508
box -48 -56 1008 834
use sg13g2_a21oi_1  _418_
timestamp 1683973020
transform -1 0 3744 0 1 34020
box -48 -56 528 834
use sg13g2_a22oi_1  _419_
timestamp 1685173987
transform -1 0 7968 0 -1 34020
box -48 -56 624 834
use sg13g2_o21ai_1  _420_
timestamp 1685175443
transform -1 0 15360 0 1 5292
box -48 -56 538 834
use sg13g2_a21o_1  _421_
timestamp 1677175127
transform 1 0 16128 0 -1 6804
box -48 -56 720 834
use sg13g2_mux2_1  _422_
timestamp 1677247768
transform -1 0 16896 0 1 5292
box -48 -56 1008 834
use sg13g2_a21oi_1  _423_
timestamp 1683973020
transform 1 0 15648 0 -1 6804
box -48 -56 528 834
use sg13g2_mux2_1  _424_
timestamp 1677247768
transform 1 0 16608 0 -1 5292
box -48 -56 1008 834
use sg13g2_o21ai_1  _425_
timestamp 1685175443
transform -1 0 18048 0 1 5292
box -48 -56 538 834
use sg13g2_a21o_1  _426_
timestamp 1677175127
transform 1 0 16896 0 1 5292
box -48 -56 720 834
use sg13g2_a21oi_1  _427_
timestamp 1683973020
transform 1 0 16800 0 -1 6804
box -48 -56 528 834
use sg13g2_a22oi_1  _428_
timestamp 1685173987
transform 1 0 15360 0 1 5292
box -48 -56 624 834
use sg13g2_o21ai_1  _429_
timestamp 1685175443
transform 1 0 2784 0 1 23436
box -48 -56 538 834
use sg13g2_nand2b_1  _430_
timestamp 1676567195
transform 1 0 2784 0 -1 24948
box -48 -56 528 834
use sg13g2_o21ai_1  _431_
timestamp 1685175443
transform 1 0 3264 0 1 23436
box -48 -56 538 834
use sg13g2_mux4_1  _432_
timestamp 1677257233
transform 1 0 17568 0 1 37044
box -48 -56 2064 834
use sg13g2_mux4_1  _433_
timestamp 1677257233
transform 1 0 7584 0 1 30996
box -48 -56 2064 834
use sg13g2_mux4_1  _434_
timestamp 1677257233
transform 1 0 9888 0 1 30996
box -48 -56 2064 834
use sg13g2_mux4_1  _435_
timestamp 1677257233
transform 1 0 17376 0 -1 35532
box -48 -56 2064 834
use sg13g2_mux4_1  _436_
timestamp 1677257233
transform 1 0 17568 0 -1 30996
box -48 -56 2064 834
use sg13g2_mux4_1  _437_
timestamp 1677257233
transform 1 0 6720 0 1 29484
box -48 -56 2064 834
use sg13g2_mux4_1  _438_
timestamp 1677257233
transform 1 0 10272 0 1 29484
box -48 -56 2064 834
use sg13g2_mux4_1  _439_
timestamp 1677257233
transform 1 0 16992 0 1 32508
box -48 -56 2064 834
use sg13g2_mux4_1  _440_
timestamp 1677257233
transform 1 0 14592 0 -1 32508
box -48 -56 2064 834
use sg13g2_mux4_1  _441_
timestamp 1677257233
transform 1 0 6336 0 1 35532
box -48 -56 2064 834
use sg13g2_mux4_1  _442_
timestamp 1677257233
transform 1 0 9792 0 -1 34020
box -48 -56 2064 834
use sg13g2_mux4_1  _443_
timestamp 1677257233
transform 1 0 15840 0 -1 34020
box -48 -56 2064 834
use sg13g2_mux4_1  _444_
timestamp 1677257233
transform 1 0 16992 0 1 29484
box -48 -56 2064 834
use sg13g2_mux4_1  _445_
timestamp 1677257233
transform 1 0 5376 0 -1 27972
box -48 -56 2064 834
use sg13g2_mux4_1  _446_
timestamp 1677257233
transform 1 0 9984 0 1 27972
box -48 -56 2064 834
use sg13g2_mux4_1  _447_
timestamp 1677257233
transform 1 0 14592 0 -1 27972
box -48 -56 2064 834
use sg13g2_mux4_1  _448_
timestamp 1677257233
transform 1 0 17376 0 1 27972
box -48 -56 2064 834
use sg13g2_mux4_1  _449_
timestamp 1677257233
transform 1 0 7392 0 -1 27972
box -48 -56 2064 834
use sg13g2_mux4_1  _450_
timestamp 1677257233
transform 1 0 10272 0 -1 27972
box -48 -56 2064 834
use sg13g2_mux4_1  _451_
timestamp 1677257233
transform 1 0 16416 0 1 26460
box -48 -56 2064 834
use sg13g2_mux4_1  _452_
timestamp 1677257233
transform 1 0 17280 0 -1 26460
box -48 -56 2064 834
use sg13g2_mux4_1  _453_
timestamp 1677257233
transform 1 0 6912 0 1 24948
box -48 -56 2064 834
use sg13g2_mux4_1  _454_
timestamp 1677257233
transform 1 0 9792 0 -1 24948
box -48 -56 2064 834
use sg13g2_mux4_1  _455_
timestamp 1677257233
transform 1 0 16320 0 -1 24948
box -48 -56 2064 834
use sg13g2_mux4_1  _456_
timestamp 1677257233
transform 1 0 13728 0 1 29484
box -48 -56 2064 834
use sg13g2_mux4_1  _457_
timestamp 1677257233
transform 1 0 3552 0 1 24948
box -48 -56 2064 834
use sg13g2_mux4_1  _458_
timestamp 1677257233
transform 1 0 10560 0 1 23436
box -48 -56 2064 834
use sg13g2_mux4_1  _459_
timestamp 1677257233
transform 1 0 13536 0 1 24948
box -48 -56 2064 834
use sg13g2_mux4_1  _460_
timestamp 1677257233
transform 1 0 13152 0 1 27972
box -48 -56 2064 834
use sg13g2_mux4_1  _461_
timestamp 1677257233
transform 1 0 3168 0 -1 26460
box -48 -56 2064 834
use sg13g2_mux4_1  _462_
timestamp 1677257233
transform 1 0 9792 0 1 21924
box -48 -56 2064 834
use sg13g2_mux4_1  _463_
timestamp 1677257233
transform 1 0 13632 0 1 23436
box -48 -56 2064 834
use sg13g2_mux4_1  _464_
timestamp 1677257233
transform 1 0 17664 0 1 23436
box -48 -56 2064 834
use sg13g2_mux4_1  _465_
timestamp 1677257233
transform 1 0 7296 0 -1 21924
box -48 -56 2064 834
use sg13g2_mux4_1  _466_
timestamp 1677257233
transform 1 0 10656 0 1 24948
box -48 -56 2064 834
use sg13g2_mux4_1  _467_
timestamp 1677257233
transform 1 0 16800 0 -1 21924
box -48 -56 2064 834
use sg13g2_mux4_1  _468_
timestamp 1677257233
transform 1 0 17376 0 1 20412
box -48 -56 2064 834
use sg13g2_mux4_1  _469_
timestamp 1677257233
transform 1 0 5952 0 1 20412
box -48 -56 2064 834
use sg13g2_mux4_1  _470_
timestamp 1677257233
transform 1 0 9888 0 1 8316
box -48 -56 2064 834
use sg13g2_mux4_1  _471_
timestamp 1677257233
transform 1 0 16800 0 1 18900
box -48 -56 2064 834
use sg13g2_mux4_1  _472_
timestamp 1677257233
transform 1 0 17568 0 -1 18900
box -48 -56 2064 834
use sg13g2_mux4_1  _473_
timestamp 1677257233
transform 1 0 8544 0 -1 20412
box -48 -56 2064 834
use sg13g2_mux4_1  _474_
timestamp 1677257233
transform 1 0 5280 0 -1 18900
box -48 -56 2064 834
use sg13g2_mux4_1  _475_
timestamp 1677257233
transform 1 0 14688 0 1 20412
box -48 -56 2064 834
use sg13g2_mux4_1  _476_
timestamp 1677257233
transform 1 0 12672 0 -1 21924
box -48 -56 2064 834
use sg13g2_mux4_1  _477_
timestamp 1677257233
transform 1 0 7008 0 1 17388
box -48 -56 2064 834
use sg13g2_mux4_1  _478_
timestamp 1677257233
transform 1 0 2304 0 -1 27972
box -48 -56 2064 834
use sg13g2_mux4_1  _479_
timestamp 1677257233
transform 1 0 9024 0 1 17388
box -48 -56 2064 834
use sg13g2_mux4_1  _480_
timestamp 1677257233
transform 1 0 13056 0 -1 2268
box -48 -56 2064 834
use sg13g2_mux4_1  _481_
timestamp 1677257233
transform -1 0 4416 0 -1 3780
box -48 -56 2064 834
use sg13g2_mux4_1  _482_
timestamp 1677257233
transform 1 0 6912 0 -1 5292
box -48 -56 2064 834
use sg13g2_mux4_1  _483_
timestamp 1677257233
transform 1 0 10752 0 1 2268
box -48 -56 2064 834
use sg13g2_mux4_1  _484_
timestamp 1677257233
transform 1 0 11232 0 1 3780
box -48 -56 2064 834
use sg13g2_mux4_1  _485_
timestamp 1677257233
transform 1 0 5760 0 -1 14364
box -48 -56 2064 834
use sg13g2_mux4_1  _486_
timestamp 1677257233
transform 1 0 6240 0 -1 8316
box -48 -56 2064 834
use sg13g2_mux4_1  _487_
timestamp 1677257233
transform 1 0 12768 0 -1 6804
box -48 -56 2064 834
use sg13g2_nor3_1  _488_
timestamp 1676639442
transform 1 0 12576 0 1 20412
box -48 -56 528 834
use sg13g2_nand2b_1  _489_
timestamp 1676567195
transform 1 0 13152 0 1 18900
box -48 -56 528 834
use sg13g2_a221oi_1  _490_
timestamp 1685197497
transform -1 0 13056 0 -1 20412
box -48 -56 816 834
use sg13g2_mux4_1  _491_
timestamp 1677257233
transform 1 0 11520 0 -1 17388
box -48 -56 2064 834
use sg13g2_nor3_1  _492_
timestamp 1676639442
transform 1 0 4032 0 -1 15876
box -48 -56 528 834
use sg13g2_nand2b_1  _493_
timestamp 1676567195
transform 1 0 5184 0 -1 17388
box -48 -56 528 834
use sg13g2_a221oi_1  _494_
timestamp 1685197497
transform 1 0 6816 0 1 15876
box -48 -56 816 834
use sg13g2_mux4_1  _495_
timestamp 1677257233
transform 1 0 5472 0 -1 12852
box -48 -56 2064 834
use sg13g2_nor3_1  _496_
timestamp 1676639442
transform 1 0 2112 0 -1 30996
box -48 -56 528 834
use sg13g2_nand2b_1  _497_
timestamp 1676567195
transform 1 0 3552 0 1 29484
box -48 -56 528 834
use sg13g2_a221oi_1  _498_
timestamp 1685197497
transform 1 0 2784 0 1 29484
box -48 -56 816 834
use sg13g2_mux4_1  _499_
timestamp 1677257233
transform 1 0 4224 0 -1 30996
box -48 -56 2064 834
use sg13g2_nor3_1  _500_
timestamp 1676639442
transform 1 0 14688 0 1 8316
box -48 -56 528 834
use sg13g2_nand2b_1  _501_
timestamp 1676567195
transform 1 0 15840 0 1 6804
box -48 -56 528 834
use sg13g2_a221oi_1  _502_
timestamp 1685197497
transform 1 0 15168 0 1 8316
box -48 -56 816 834
use sg13g2_mux4_1  _503_
timestamp 1677257233
transform 1 0 12960 0 -1 5292
box -48 -56 2064 834
use sg13g2_mux4_1  _504_
timestamp 1677257233
transform 1 0 14784 0 1 9828
box -48 -56 2064 834
use sg13g2_mux4_1  _505_
timestamp 1677257233
transform -1 0 4512 0 1 12852
box -48 -56 2064 834
use sg13g2_mux4_1  _506_
timestamp 1677257233
transform -1 0 7680 0 -1 9828
box -48 -56 2064 834
use sg13g2_mux4_1  _507_
timestamp 1677257233
transform 1 0 10656 0 -1 15876
box -48 -56 2064 834
use sg13g2_mux4_1  _508_
timestamp 1677257233
transform 1 0 11520 0 1 6804
box -48 -56 2064 834
use sg13g2_mux4_1  _509_
timestamp 1677257233
transform 1 0 3456 0 1 27972
box -48 -56 2064 834
use sg13g2_mux4_1  _510_
timestamp 1677257233
transform 1 0 2304 0 -1 18900
box -48 -56 2064 834
use sg13g2_mux4_1  _511_
timestamp 1677257233
transform 1 0 10464 0 1 12852
box -48 -56 2064 834
use sg13g2_mux4_1  _512_
timestamp 1677257233
transform 1 0 11424 0 -1 18900
box -48 -56 2064 834
use sg13g2_mux4_1  _513_
timestamp 1677257233
transform 1 0 3168 0 1 15876
box -48 -56 2064 834
use sg13g2_mux4_1  _514_
timestamp 1677257233
transform -1 0 4704 0 -1 32508
box -48 -56 2064 834
use sg13g2_mux4_1  _515_
timestamp 1677257233
transform 1 0 12768 0 -1 9828
box -48 -56 2064 834
use sg13g2_dlhq_1  _516_
timestamp 1678805552
transform 1 0 11136 0 -1 9828
box -50 -56 1692 834
use sg13g2_dlhq_1  _517_
timestamp 1678805552
transform 1 0 12960 0 1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _518_
timestamp 1678805552
transform 1 0 1152 0 1 34020
box -50 -56 1692 834
use sg13g2_dlhq_1  _519_
timestamp 1678805552
transform -1 0 3840 0 1 32508
box -50 -56 1692 834
use sg13g2_dlhq_1  _520_
timestamp 1678805552
transform 1 0 1152 0 -1 15876
box -50 -56 1692 834
use sg13g2_dlhq_1  _521_
timestamp 1678805552
transform 1 0 3456 0 -1 17388
box -50 -56 1692 834
use sg13g2_dlhq_1  _522_
timestamp 1678805552
transform 1 0 9792 0 -1 18900
box -50 -56 1692 834
use sg13g2_dlhq_1  _523_
timestamp 1678805552
transform 1 0 11520 0 1 18900
box -50 -56 1692 834
use sg13g2_dlhq_1  _524_
timestamp 1678805552
transform 1 0 8832 0 1 12852
box -50 -56 1692 834
use sg13g2_dlhq_1  _525_
timestamp 1678805552
transform 1 0 10752 0 -1 12852
box -50 -56 1692 834
use sg13g2_dlhq_1  _526_
timestamp 1678805552
transform 1 0 1152 0 -1 17388
box -50 -56 1692 834
use sg13g2_dlhq_1  _527_
timestamp 1678805552
transform 1 0 2496 0 1 17388
box -50 -56 1692 834
use sg13g2_dlhq_1  _528_
timestamp 1678805552
transform 1 0 3744 0 -1 29484
box -50 -56 1692 834
use sg13g2_dlhq_1  _529_
timestamp 1678805552
transform 1 0 1440 0 -1 29484
box -50 -56 1692 834
use sg13g2_dlhq_1  _530_
timestamp 1678805552
transform 1 0 11616 0 -1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _531_
timestamp 1678805552
transform 1 0 9888 0 1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _532_
timestamp 1678805552
transform 1 0 9408 0 1 15876
box -50 -56 1692 834
use sg13g2_dlhq_1  _533_
timestamp 1678805552
transform 1 0 10656 0 1 14364
box -50 -56 1692 834
use sg13g2_dlhq_1  _534_
timestamp 1678805552
transform -1 0 7296 0 1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _535_
timestamp 1678805552
transform 1 0 4032 0 -1 9828
box -50 -56 1692 834
use sg13g2_dlhq_1  _536_
timestamp 1678805552
transform -1 0 3840 0 -1 12852
box -50 -56 1692 834
use sg13g2_dlhq_1  _537_
timestamp 1678805552
transform 1 0 1152 0 -1 11340
box -50 -56 1692 834
use sg13g2_dlhq_1  _538_
timestamp 1678805552
transform 1 0 13152 0 1 9828
box -50 -56 1692 834
use sg13g2_dlhq_1  _539_
timestamp 1678805552
transform 1 0 15072 0 -1 9828
box -50 -56 1692 834
use sg13g2_dlhq_1  _540_
timestamp 1678805552
transform 1 0 14688 0 1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _541_
timestamp 1678805552
transform 1 0 14976 0 -1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _542_
timestamp 1678805552
transform 1 0 14112 0 -1 3780
box -50 -56 1692 834
use sg13g2_dlhq_1  _543_
timestamp 1678805552
transform 1 0 4128 0 1 34020
box -50 -56 1692 834
use sg13g2_dlhq_1  _544_
timestamp 1678805552
transform 1 0 4128 0 -1 34020
box -50 -56 1692 834
use sg13g2_dlhq_1  _545_
timestamp 1678805552
transform 1 0 3936 0 1 32508
box -50 -56 1692 834
use sg13g2_dlhq_1  _546_
timestamp 1678805552
transform 1 0 6144 0 1 14364
box -50 -56 1692 834
use sg13g2_dlhq_1  _547_
timestamp 1678805552
transform 1 0 7776 0 1 15876
box -50 -56 1692 834
use sg13g2_dlhq_1  _548_
timestamp 1678805552
transform 1 0 6144 0 -1 15876
box -50 -56 1692 834
use sg13g2_dlhq_1  _549_
timestamp 1678805552
transform 1 0 13440 0 -1 18900
box -50 -56 1692 834
use sg13g2_dlhq_1  _550_
timestamp 1678805552
transform -1 0 15264 0 -1 17388
box -50 -56 1692 834
use sg13g2_dlhq_1  _551_
timestamp 1678805552
transform -1 0 15072 0 -1 20412
box -50 -56 1692 834
use sg13g2_dlhq_1  _552_
timestamp 1678805552
transform 1 0 11328 0 -1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _553_
timestamp 1678805552
transform 1 0 13248 0 1 3780
box -50 -56 1692 834
use sg13g2_dlhq_1  _554_
timestamp 1678805552
transform 1 0 2592 0 -1 30996
box -50 -56 1692 834
use sg13g2_dlhq_1  _555_
timestamp 1678805552
transform 1 0 4320 0 1 30996
box -50 -56 1692 834
use sg13g2_dlhq_1  _556_
timestamp 1678805552
transform 1 0 3840 0 -1 12852
box -50 -56 1692 834
use sg13g2_dlhq_1  _557_
timestamp 1678805552
transform 1 0 5376 0 1 11340
box -50 -56 1692 834
use sg13g2_dlhq_1  _558_
timestamp 1678805552
transform 1 0 9888 0 -1 17388
box -50 -56 1692 834
use sg13g2_dlhq_1  _559_
timestamp 1678805552
transform 1 0 11808 0 1 15876
box -50 -56 1692 834
use sg13g2_dlhq_1  _560_
timestamp 1678805552
transform 1 0 11136 0 -1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _561_
timestamp 1678805552
transform 1 0 13152 0 1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _562_
timestamp 1678805552
transform 1 0 4608 0 -1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _563_
timestamp 1678805552
transform 1 0 6336 0 1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _564_
timestamp 1678805552
transform 1 0 5568 0 1 12852
box -50 -56 1692 834
use sg13g2_dlhq_1  _565_
timestamp 1678805552
transform 1 0 4320 0 1 14364
box -50 -56 1692 834
use sg13g2_dlhq_1  _566_
timestamp 1678805552
transform 1 0 11328 0 1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _567_
timestamp 1678805552
transform 1 0 9696 0 -1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _568_
timestamp 1678805552
transform 1 0 11136 0 -1 3780
box -50 -56 1692 834
use sg13g2_dlhq_1  _569_
timestamp 1678805552
transform 1 0 9120 0 -1 3780
box -50 -56 1692 834
use sg13g2_dlhq_1  _570_
timestamp 1678805552
transform 1 0 5184 0 -1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _571_
timestamp 1678805552
transform 1 0 7200 0 1 3780
box -50 -56 1692 834
use sg13g2_dlhq_1  _572_
timestamp 1678805552
transform 1 0 2784 0 -1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _573_
timestamp 1678805552
transform 1 0 1920 0 1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _574_
timestamp 1678805552
transform 1 0 13152 0 1 756
box -50 -56 1692 834
use sg13g2_dlhq_1  _575_
timestamp 1678805552
transform 1 0 11424 0 -1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _576_
timestamp 1678805552
transform 1 0 15648 0 1 756
box -50 -56 1692 834
use sg13g2_dlhq_1  _577_
timestamp 1678805552
transform 1 0 15168 0 -1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _578_
timestamp 1678805552
transform 1 0 15456 0 -1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _579_
timestamp 1678805552
transform 1 0 5184 0 -1 24948
box -50 -56 1692 834
use sg13g2_dlhq_1  _580_
timestamp 1678805552
transform 1 0 5568 0 1 23436
box -50 -56 1692 834
use sg13g2_dlhq_1  _581_
timestamp 1678805552
transform 1 0 7200 0 1 23436
box -50 -56 1692 834
use sg13g2_dlhq_1  _582_
timestamp 1678805552
transform 1 0 6912 0 1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _583_
timestamp 1678805552
transform 1 0 8256 0 1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _584_
timestamp 1678805552
transform 1 0 8928 0 1 3780
box -50 -56 1692 834
use sg13g2_dlhq_1  _585_
timestamp 1678805552
transform 1 0 13728 0 -1 12852
box -50 -56 1692 834
use sg13g2_dlhq_1  _586_
timestamp 1678805552
transform 1 0 14880 0 -1 14364
box -50 -56 1692 834
use sg13g2_dlhq_1  _587_
timestamp 1678805552
transform 1 0 14976 0 1 11340
box -50 -56 1692 834
use sg13g2_dlhq_1  _588_
timestamp 1678805552
transform 1 0 7200 0 1 18900
box -50 -56 1692 834
use sg13g2_dlhq_1  _589_
timestamp 1678805552
transform 1 0 8160 0 -1 18900
box -50 -56 1692 834
use sg13g2_dlhq_1  _590_
timestamp 1678805552
transform 1 0 1152 0 1 26460
box -50 -56 1692 834
use sg13g2_dlhq_1  _591_
timestamp 1678805552
transform 1 0 1824 0 1 27972
box -50 -56 1692 834
use sg13g2_dlhq_1  _592_
timestamp 1678805552
transform 1 0 5664 0 -1 17388
box -50 -56 1692 834
use sg13g2_dlhq_1  _593_
timestamp 1678805552
transform 1 0 7392 0 -1 17388
box -50 -56 1692 834
use sg13g2_dlhq_1  _594_
timestamp 1678805552
transform 1 0 11808 0 1 21924
box -50 -56 1692 834
use sg13g2_dlhq_1  _595_
timestamp 1678805552
transform 1 0 13440 0 1 21924
box -50 -56 1692 834
use sg13g2_dlhq_1  _596_
timestamp 1678805552
transform 1 0 14784 0 -1 21924
box -50 -56 1692 834
use sg13g2_dlhq_1  _597_
timestamp 1678805552
transform 1 0 13056 0 1 20412
box -50 -56 1692 834
use sg13g2_dlhq_1  _598_
timestamp 1678805552
transform 1 0 5184 0 1 17388
box -50 -56 1692 834
use sg13g2_dlhq_1  _599_
timestamp 1678805552
transform 1 0 4032 0 1 18900
box -50 -56 1692 834
use sg13g2_dlhq_1  _600_
timestamp 1678805552
transform 1 0 8832 0 1 18900
box -50 -56 1692 834
use sg13g2_dlhq_1  _601_
timestamp 1678805552
transform 1 0 6912 0 -1 20412
box -50 -56 1692 834
use sg13g2_dlhq_1  _602_
timestamp 1678805552
transform 1 0 18336 0 -1 17388
box -50 -56 1692 834
use sg13g2_dlhq_1  _603_
timestamp 1678805552
transform 1 0 15936 0 -1 18900
box -50 -56 1692 834
use sg13g2_dlhq_1  _604_
timestamp 1678805552
transform 1 0 17184 0 1 17388
box -50 -56 1692 834
use sg13g2_dlhq_1  _605_
timestamp 1678805552
transform 1 0 15168 0 1 18900
box -50 -56 1692 834
use sg13g2_dlhq_1  _606_
timestamp 1678805552
transform 1 0 9984 0 -1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _607_
timestamp 1678805552
transform 1 0 8352 0 -1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _608_
timestamp 1678805552
transform 1 0 5280 0 -1 20412
box -50 -56 1692 834
use sg13g2_dlhq_1  _609_
timestamp 1678805552
transform 1 0 3936 0 -1 21924
box -50 -56 1692 834
use sg13g2_dlhq_1  _610_
timestamp 1678805552
transform 1 0 18144 0 -1 20412
box -50 -56 1692 834
use sg13g2_dlhq_1  _611_
timestamp 1678805552
transform 1 0 15744 0 -1 20412
box -50 -56 1692 834
use sg13g2_dlhq_1  _612_
timestamp 1678805552
transform 1 0 15168 0 1 21924
box -50 -56 1692 834
use sg13g2_dlhq_1  _613_
timestamp 1678805552
transform 1 0 17088 0 1 21924
box -50 -56 1692 834
use sg13g2_dlhq_1  _614_
timestamp 1678805552
transform 1 0 9120 0 -1 26460
box -50 -56 1692 834
use sg13g2_dlhq_1  _615_
timestamp 1678805552
transform 1 0 10752 0 -1 26460
box -50 -56 1692 834
use sg13g2_dlhq_1  _616_
timestamp 1678805552
transform 1 0 5568 0 -1 21924
box -50 -56 1692 834
use sg13g2_dlhq_1  _617_
timestamp 1678805552
transform 1 0 7968 0 1 20412
box -50 -56 1692 834
use sg13g2_dlhq_1  _618_
timestamp 1678805552
transform 1 0 16032 0 1 23436
box -50 -56 1692 834
use sg13g2_dlhq_1  _619_
timestamp 1678805552
transform 1 0 18240 0 -1 23436
box -50 -56 1692 834
use sg13g2_dlhq_1  _620_
timestamp 1678805552
transform 1 0 12288 0 -1 23436
box -50 -56 1692 834
use sg13g2_dlhq_1  _621_
timestamp 1678805552
transform 1 0 13824 0 -1 24948
box -50 -56 1692 834
use sg13g2_dlhq_1  _622_
timestamp 1678805552
transform 1 0 8160 0 1 21924
box -50 -56 1692 834
use sg13g2_dlhq_1  _623_
timestamp 1678805552
transform 1 0 9792 0 -1 21924
box -50 -56 1692 834
use sg13g2_dlhq_1  _624_
timestamp 1678805552
transform 1 0 1632 0 1 24948
box -50 -56 1692 834
use sg13g2_dlhq_1  _625_
timestamp 1678805552
transform 1 0 2784 0 1 26460
box -50 -56 1692 834
use sg13g2_dlhq_1  _626_
timestamp 1678805552
transform 1 0 11904 0 -1 29484
box -50 -56 1692 834
use sg13g2_dlhq_1  _627_
timestamp 1678805552
transform 1 0 13536 0 -1 29484
box -50 -56 1692 834
use sg13g2_dlhq_1  _628_
timestamp 1678805552
transform 1 0 12384 0 -1 26460
box -50 -56 1692 834
use sg13g2_dlhq_1  _629_
timestamp 1678805552
transform 1 0 13536 0 1 26460
box -50 -56 1692 834
use sg13g2_dlhq_1  _630_
timestamp 1678805552
transform 1 0 8928 0 1 23436
box -50 -56 1692 834
use sg13g2_dlhq_1  _631_
timestamp 1678805552
transform 1 0 10656 0 -1 23436
box -50 -56 1692 834
use sg13g2_dlhq_1  _632_
timestamp 1678805552
transform 1 0 1536 0 -1 26460
box -50 -56 1692 834
use sg13g2_dlhq_1  _633_
timestamp 1678805552
transform 1 0 3552 0 -1 24948
box -50 -56 1692 834
use sg13g2_dlhq_1  _634_
timestamp 1678805552
transform 1 0 12384 0 -1 30996
box -50 -56 1692 834
use sg13g2_dlhq_1  _635_
timestamp 1678805552
transform 1 0 14016 0 -1 30996
box -50 -56 1692 834
use sg13g2_dlhq_1  _636_
timestamp 1678805552
transform 1 0 14784 0 -1 26460
box -50 -56 1692 834
use sg13g2_dlhq_1  _637_
timestamp 1678805552
transform 1 0 16320 0 1 24948
box -50 -56 1692 834
use sg13g2_dlhq_1  _638_
timestamp 1678805552
transform 1 0 8160 0 -1 24948
box -50 -56 1692 834
use sg13g2_dlhq_1  _639_
timestamp 1678805552
transform 1 0 9024 0 1 24948
box -50 -56 1692 834
use sg13g2_dlhq_1  _640_
timestamp 1678805552
transform 1 0 5376 0 -1 26460
box -50 -56 1692 834
use sg13g2_dlhq_1  _641_
timestamp 1678805552
transform 1 0 7008 0 -1 26460
box -50 -56 1692 834
use sg13g2_dlhq_1  _642_
timestamp 1678805552
transform 1 0 16608 0 -1 27972
box -50 -56 1692 834
use sg13g2_dlhq_1  _643_
timestamp 1678805552
transform 1 0 17952 0 1 24948
box -50 -56 1692 834
use sg13g2_dlhq_1  _644_
timestamp 1678805552
transform -1 0 20064 0 1 26460
box -50 -56 1692 834
use sg13g2_dlhq_1  _645_
timestamp 1678805552
transform 1 0 15168 0 1 27972
box -50 -56 1692 834
use sg13g2_dlhq_1  _646_
timestamp 1678805552
transform 1 0 10752 0 1 26460
box -50 -56 1692 834
use sg13g2_dlhq_1  _647_
timestamp 1678805552
transform 1 0 8832 0 1 26460
box -50 -56 1692 834
use sg13g2_dlhq_1  _648_
timestamp 1678805552
transform 1 0 7680 0 1 27972
box -50 -56 1692 834
use sg13g2_dlhq_1  _649_
timestamp 1678805552
transform 1 0 5856 0 1 27972
box -50 -56 1692 834
use sg13g2_dlhq_1  _650_
timestamp 1678805552
transform 1 0 18240 0 -1 27972
box -50 -56 1692 834
use sg13g2_dlhq_1  _651_
timestamp 1678805552
transform -1 0 18432 0 -1 29484
box -50 -56 1692 834
use sg13g2_dlhq_1  _652_
timestamp 1678805552
transform 1 0 15168 0 -1 29484
box -50 -56 1692 834
use sg13g2_dlhq_1  _653_
timestamp 1678805552
transform 1 0 12960 0 -1 27972
box -50 -56 1692 834
use sg13g2_dlhq_1  _654_
timestamp 1678805552
transform 1 0 10272 0 -1 29484
box -50 -56 1692 834
use sg13g2_dlhq_1  _655_
timestamp 1678805552
transform 1 0 8640 0 -1 29484
box -50 -56 1692 834
use sg13g2_dlhq_1  _656_
timestamp 1678805552
transform 1 0 6048 0 1 26460
box -50 -56 1692 834
use sg13g2_dlhq_1  _657_
timestamp 1678805552
transform 1 0 4416 0 1 26460
box -50 -56 1692 834
use sg13g2_dlhq_1  _658_
timestamp 1678805552
transform 1 0 18432 0 -1 29484
box -50 -56 1692 834
use sg13g2_dlhq_1  _659_
timestamp 1678805552
transform 1 0 15648 0 -1 30996
box -50 -56 1692 834
use sg13g2_dlhq_1  _660_
timestamp 1678805552
transform 1 0 15168 0 1 34020
box -50 -56 1692 834
use sg13g2_dlhq_1  _661_
timestamp 1678805552
transform 1 0 16800 0 1 34020
box -50 -56 1692 834
use sg13g2_dlhq_1  _662_
timestamp 1678805552
transform 1 0 8160 0 -1 34020
box -50 -56 1692 834
use sg13g2_dlhq_1  _663_
timestamp 1678805552
transform 1 0 9312 0 -1 35532
box -50 -56 1692 834
use sg13g2_dlhq_1  _664_
timestamp 1678805552
transform 1 0 4896 0 -1 37044
box -50 -56 1692 834
use sg13g2_dlhq_1  _665_
timestamp 1678805552
transform 1 0 6048 0 -1 35532
box -50 -56 1692 834
use sg13g2_dlhq_1  _666_
timestamp 1678805552
transform 1 0 13248 0 1 32508
box -50 -56 1692 834
use sg13g2_dlhq_1  _667_
timestamp 1678805552
transform 1 0 14784 0 1 30996
box -50 -56 1692 834
use sg13g2_dlhq_1  _668_
timestamp 1678805552
transform 1 0 17376 0 -1 32508
box -50 -56 1692 834
use sg13g2_dlhq_1  _669_
timestamp 1678805552
transform 1 0 15360 0 1 32508
box -50 -56 1692 834
use sg13g2_dlhq_1  _670_
timestamp 1678805552
transform 1 0 10752 0 -1 30996
box -50 -56 1692 834
use sg13g2_dlhq_1  _671_
timestamp 1678805552
transform 1 0 8832 0 -1 30996
box -50 -56 1692 834
use sg13g2_dlhq_1  _672_
timestamp 1678805552
transform 1 0 6912 0 -1 29484
box -50 -56 1692 834
use sg13g2_dlhq_1  _673_
timestamp 1678805552
transform 1 0 5088 0 1 29484
box -50 -56 1692 834
use sg13g2_dlhq_1  _674_
timestamp 1678805552
transform 1 0 18336 0 1 30996
box -50 -56 1692 834
use sg13g2_dlhq_1  _675_
timestamp 1678805552
transform 1 0 16416 0 1 30996
box -50 -56 1692 834
use sg13g2_dlhq_1  _676_
timestamp 1678805552
transform 1 0 18240 0 1 35532
box -50 -56 1692 834
use sg13g2_dlhq_1  _677_
timestamp 1678805552
transform -1 0 18816 0 -1 37044
box -50 -56 1692 834
use sg13g2_dlhq_1  _678_
timestamp 1678805552
transform 1 0 10080 0 1 32508
box -50 -56 1692 834
use sg13g2_dlhq_1  _679_
timestamp 1678805552
transform 1 0 8544 0 -1 32508
box -50 -56 1692 834
use sg13g2_dlhq_1  _680_
timestamp 1678805552
transform 1 0 7968 0 1 32508
box -50 -56 1692 834
use sg13g2_dlhq_1  _681_
timestamp 1678805552
transform 1 0 5952 0 1 30996
box -50 -56 1692 834
use sg13g2_dlhq_1  _682_
timestamp 1678805552
transform 1 0 16608 0 -1 41580
box -50 -56 1692 834
use sg13g2_dlhq_1  _683_
timestamp 1678805552
transform -1 0 18816 0 -1 38556
box -50 -56 1692 834
use sg13g2_dlhq_1  _684_
timestamp 1678805552
transform 1 0 16800 0 1 11340
box -50 -56 1692 834
use sg13g2_dlhq_1  _685_
timestamp 1678805552
transform 1 0 18336 0 -1 12852
box -50 -56 1692 834
use sg13g2_dlhq_1  _686_
timestamp 1678805552
transform 1 0 17760 0 1 12852
box -50 -56 1692 834
use sg13g2_dlhq_1  _687_
timestamp 1678805552
transform 1 0 1344 0 1 15876
box -50 -56 1692 834
use sg13g2_dlhq_1  _688_
timestamp 1678805552
transform 1 0 1152 0 1 11340
box -50 -56 1692 834
use sg13g2_dlhq_1  _689_
timestamp 1678805552
transform 1 0 1152 0 1 14364
box -50 -56 1692 834
use sg13g2_dlhq_1  _690_
timestamp 1678805552
transform 1 0 8256 0 1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _691_
timestamp 1678805552
transform 1 0 7680 0 -1 9828
box -50 -56 1692 834
use sg13g2_dlhq_1  _692_
timestamp 1678805552
transform -1 0 10176 0 -1 12852
box -50 -56 1692 834
use sg13g2_dlhq_1  _693_
timestamp 1678805552
transform 1 0 17568 0 1 14364
box -50 -56 1692 834
use sg13g2_dlhq_1  _694_
timestamp 1678805552
transform 1 0 18624 0 -1 14364
box -50 -56 1692 834
use sg13g2_dlhq_1  _695_
timestamp 1678805552
transform 1 0 18144 0 1 15876
box -50 -56 1692 834
use sg13g2_dlhq_1  _696_
timestamp 1678805552
transform 1 0 18336 0 -1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _697_
timestamp 1678805552
transform 1 0 18048 0 1 756
box -50 -56 1692 834
use sg13g2_dlhq_1  _698_
timestamp 1678805552
transform 1 0 18048 0 -1 3780
box -50 -56 1692 834
use sg13g2_dlhq_1  _699_
timestamp 1678805552
transform 1 0 1536 0 1 20412
box -50 -56 1692 834
use sg13g2_dlhq_1  _700_
timestamp 1678805552
transform 1 0 1440 0 -1 20412
box -50 -56 1692 834
use sg13g2_dlhq_1  _701_
timestamp 1678805552
transform 1 0 1152 0 1 18900
box -50 -56 1692 834
use sg13g2_dlhq_1  _702_
timestamp 1678805552
transform 1 0 1152 0 1 3780
box -50 -56 1692 834
use sg13g2_dlhq_1  _703_
timestamp 1678805552
transform 1 0 1248 0 -1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _704_
timestamp 1678805552
transform 1 0 1152 0 -1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _705_
timestamp 1678805552
transform 1 0 10944 0 -1 14364
box -50 -56 1692 834
use sg13g2_dlhq_1  _706_
timestamp 1678805552
transform 1 0 12768 0 -1 14364
box -50 -56 1692 834
use sg13g2_dlhq_1  _707_
timestamp 1678805552
transform 1 0 12672 0 -1 15876
box -50 -56 1692 834
use sg13g2_dlhq_1  _708_
timestamp 1678805552
transform 1 0 16128 0 1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _709_
timestamp 1678805552
transform 1 0 17376 0 1 9828
box -50 -56 1692 834
use sg13g2_dlhq_1  _710_
timestamp 1678805552
transform 1 0 17760 0 1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _711_
timestamp 1678805552
transform 1 0 1440 0 -1 9828
box -50 -56 1692 834
use sg13g2_dlhq_1  _712_
timestamp 1678805552
transform 1 0 1152 0 1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _713_
timestamp 1678805552
transform 1 0 1152 0 1 9828
box -50 -56 1692 834
use sg13g2_dlhq_1  _714_
timestamp 1678805552
transform 1 0 7200 0 1 12852
box -50 -56 1692 834
use sg13g2_dlhq_1  _715_
timestamp 1678805552
transform 1 0 7008 0 1 11340
box -50 -56 1692 834
use sg13g2_dlhq_1  _716_
timestamp 1678805552
transform 1 0 5760 0 -1 11340
box -50 -56 1692 834
use sg13g2_dlhq_1  _717_
timestamp 1678805552
transform 1 0 14400 0 -1 15876
box -50 -56 1692 834
use sg13g2_dlhq_1  _718_
timestamp 1678805552
transform 1 0 15264 0 1 14364
box -50 -56 1692 834
use sg13g2_dlhq_1  _719_
timestamp 1678805552
transform 1 0 15840 0 -1 17388
box -50 -56 1692 834
use sg13g2_dlhq_1  _720_
timestamp 1678805552
transform 1 0 16608 0 1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _721_
timestamp 1678805552
transform 1 0 18240 0 1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _722_
timestamp 1678805552
transform 1 0 18240 0 1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _723_
timestamp 1678805552
transform 1 0 1344 0 -1 23436
box -50 -56 1692 834
use sg13g2_dlhq_1  _724_
timestamp 1678805552
transform 1 0 2976 0 1 21924
box -50 -56 1692 834
use sg13g2_dlhq_1  _725_
timestamp 1678805552
transform 1 0 1344 0 1 21924
box -50 -56 1692 834
use sg13g2_dlhq_1  _726_
timestamp 1678805552
transform -1 0 4416 0 1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _727_
timestamp 1678805552
transform 1 0 1152 0 1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _728_
timestamp 1678805552
transform 1 0 1152 0 -1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _729_
timestamp 1678805552
transform 1 0 10464 0 -1 11340
box -50 -56 1692 834
use sg13g2_dlhq_1  _730_
timestamp 1678805552
transform 1 0 11328 0 1 9828
box -50 -56 1692 834
use sg13g2_dlhq_1  _731_
timestamp 1678805552
transform 1 0 10080 0 1 11340
box -50 -56 1692 834
use sg13g2_dlhq_1  _732_
timestamp 1678805552
transform 1 0 1152 0 1 23436
box -50 -56 1692 834
use sg13g2_dlhq_1  _733_
timestamp 1678805552
transform 1 0 1152 0 -1 24948
box -50 -56 1692 834
use sg13g2_dlhq_1  _734_
timestamp 1678805552
transform 1 0 2688 0 1 756
box -50 -56 1692 834
use sg13g2_dlhq_1  _735_
timestamp 1678805552
transform -1 0 4896 0 -1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _736_
timestamp 1678805552
transform 1 0 4896 0 -1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _737_
timestamp 1678805552
transform 1 0 3744 0 1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _738_
timestamp 1678805552
transform -1 0 16608 0 1 35532
box -50 -56 1692 834
use sg13g2_dlhq_1  _739_
timestamp 1678805552
transform -1 0 18240 0 1 35532
box -50 -56 1692 834
use sg13g2_dlhq_1  _740_
timestamp 1678805552
transform -1 0 6336 0 -1 32508
box -50 -56 1692 834
use sg13g2_dlhq_1  _741_
timestamp 1678805552
transform -1 0 7392 0 -1 34020
box -50 -56 1692 834
use sg13g2_dlhq_1  _742_
timestamp 1678805552
transform 1 0 5568 0 1 37044
box -50 -56 1692 834
use sg13g2_dlhq_1  _743_
timestamp 1678805552
transform 1 0 7776 0 -1 38556
box -50 -56 1692 834
use sg13g2_dlhq_1  _744_
timestamp 1678805552
transform 1 0 11424 0 1 37044
box -50 -56 1692 834
use sg13g2_dlhq_1  _745_
timestamp 1678805552
transform 1 0 13248 0 1 37044
box -50 -56 1692 834
use sg13g2_dlhq_1  _746_
timestamp 1678805552
transform 1 0 13536 0 -1 38556
box -50 -56 1692 834
use sg13g2_dlhq_1  _747_
timestamp 1678805552
transform 1 0 15552 0 1 37044
box -50 -56 1692 834
use sg13g2_dlhq_1  _748_
timestamp 1678805552
transform -1 0 7680 0 -1 41580
box -50 -56 1692 834
use sg13g2_dlhq_1  _749_
timestamp 1678805552
transform -1 0 15168 0 -1 41580
box -50 -56 1692 834
use sg13g2_dlhq_1  _750_
timestamp 1678805552
transform 1 0 2016 0 1 40068
box -50 -56 1692 834
use sg13g2_dlhq_1  _751_
timestamp 1678805552
transform 1 0 4320 0 -1 40068
box -50 -56 1692 834
use sg13g2_dlhq_1  _752_
timestamp 1678805552
transform 1 0 10656 0 -1 37044
box -50 -56 1692 834
use sg13g2_dlhq_1  _753_
timestamp 1678805552
transform 1 0 12480 0 1 38556
box -50 -56 1692 834
use sg13g2_dlhq_1  _754_
timestamp 1678805552
transform 1 0 13248 0 -1 40068
box -50 -56 1692 834
use sg13g2_dlhq_1  _755_
timestamp 1678805552
transform 1 0 15168 0 -1 40068
box -50 -56 1692 834
use sg13g2_dlhq_1  _756_
timestamp 1678805552
transform -1 0 13536 0 -1 41580
box -50 -56 1692 834
use sg13g2_dlhq_1  _757_
timestamp 1678805552
transform 1 0 1728 0 -1 41580
box -50 -56 1692 834
use sg13g2_dlhq_1  _758_
timestamp 1678805552
transform 1 0 6336 0 1 40068
box -50 -56 1692 834
use sg13g2_dlhq_1  _759_
timestamp 1678805552
transform 1 0 6912 0 -1 40068
box -50 -56 1692 834
use sg13g2_dlhq_1  _760_
timestamp 1678805552
transform 1 0 10944 0 -1 35532
box -50 -56 1692 834
use sg13g2_dlhq_1  _761_
timestamp 1678805552
transform -1 0 15840 0 -1 35532
box -50 -56 1692 834
use sg13g2_dlhq_1  _762_
timestamp 1678805552
transform 1 0 10656 0 -1 32508
box -50 -56 1692 834
use sg13g2_dlhq_1  _763_
timestamp 1678805552
transform 1 0 12480 0 1 30996
box -50 -56 1692 834
use sg13g2_dlhq_1  _764_
timestamp 1678805552
transform -1 0 11136 0 1 37044
box -50 -56 1692 834
use sg13g2_dlhq_1  _765_
timestamp 1678805552
transform 1 0 1632 0 -1 40068
box -50 -56 1692 834
use sg13g2_dlhq_1  _766_
timestamp 1678805552
transform 1 0 6144 0 1 34020
box -50 -56 1692 834
use sg13g2_dlhq_1  _767_
timestamp 1678805552
transform 1 0 7680 0 -1 35532
box -50 -56 1692 834
use sg13g2_dlhq_1  _768_
timestamp 1678805552
transform 1 0 10944 0 1 34020
box -50 -56 1692 834
use sg13g2_dlhq_1  _769_
timestamp 1678805552
transform 1 0 12576 0 -1 35532
box -50 -56 1692 834
use sg13g2_dlhq_1  _770_
timestamp 1678805552
transform 1 0 7392 0 -1 37044
box -50 -56 1692 834
use sg13g2_dlhq_1  _771_
timestamp 1678805552
transform 1 0 9024 0 -1 37044
box -50 -56 1692 834
use sg13g2_dlhq_1  _772_
timestamp 1678805552
transform 1 0 1632 0 1 38556
box -50 -56 1692 834
use sg13g2_dlhq_1  _773_
timestamp 1678805552
transform -1 0 6336 0 1 35532
box -50 -56 1692 834
use sg13g2_dlhq_1  _774_
timestamp 1678805552
transform 1 0 5088 0 1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _775_
timestamp 1678805552
transform 1 0 3360 0 -1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _776_
timestamp 1678805552
transform 1 0 5184 0 -1 3780
box -50 -56 1692 834
use sg13g2_dlhq_1  _777_
timestamp 1678805552
transform 1 0 3264 0 1 3780
box -50 -56 1692 834
use sg13g2_dlhq_1  _778_
timestamp 1678805552
transform 1 0 8544 0 -1 40068
box -50 -56 1692 834
use sg13g2_dlhq_1  _779_
timestamp 1678805552
transform 1 0 10176 0 1 38556
box -50 -56 1692 834
use sg13g2_dlhq_1  _780_
timestamp 1678805552
transform 1 0 3360 0 -1 41580
box -50 -56 1692 834
use sg13g2_dlhq_1  _781_
timestamp 1678805552
transform 1 0 4032 0 1 40068
box -50 -56 1692 834
use sg13g2_dlhq_1  _782_
timestamp 1678805552
transform 1 0 8640 0 -1 41580
box -50 -56 1692 834
use sg13g2_dlhq_1  _783_
timestamp 1678805552
transform 1 0 10272 0 -1 41580
box -50 -56 1692 834
use sg13g2_dlhq_1  _784_
timestamp 1678805552
transform 1 0 8064 0 1 40068
box -50 -56 1692 834
use sg13g2_dlhq_1  _785_
timestamp 1678805552
transform -1 0 13632 0 1 40068
box -50 -56 1692 834
use sg13g2_dlhq_1  _786_
timestamp 1678805552
transform 1 0 13824 0 -1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _787_
timestamp 1678805552
transform 1 0 14208 0 1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _788_
timestamp 1678805552
transform 1 0 1152 0 1 30996
box -50 -56 1692 834
use sg13g2_dlhq_1  _789_
timestamp 1678805552
transform 1 0 1152 0 1 29484
box -50 -56 1692 834
use sg13g2_dlhq_1  _790_
timestamp 1678805552
transform -1 0 6144 0 -1 15876
box -50 -56 1692 834
use sg13g2_dlhq_1  _791_
timestamp 1678805552
transform 1 0 5184 0 1 15876
box -50 -56 1692 834
use sg13g2_dlhq_1  _792_
timestamp 1678805552
transform 1 0 10656 0 -1 20412
box -50 -56 1692 834
use sg13g2_dlhq_1  _793_
timestamp 1678805552
transform 1 0 10944 0 1 20412
box -50 -56 1692 834
use sg13g2_buf_1  _794_
timestamp 1676381911
transform -1 0 4128 0 1 23436
box -48 -56 432 834
use sg13g2_buf_1  _795_
timestamp 1676381911
transform 1 0 17952 0 -1 17388
box -48 -56 432 834
use sg13g2_buf_1  _796_
timestamp 1676381911
transform 1 0 19584 0 -1 30996
box -48 -56 432 834
use sg13g2_buf_1  _797_
timestamp 1676381911
transform 1 0 19968 0 -1 17388
box -48 -56 432 834
use sg13g2_buf_1  _798_
timestamp 1676381911
transform 1 0 19296 0 -1 21924
box -48 -56 432 834
use sg13g2_buf_1  _799_
timestamp 1676381911
transform 1 0 19776 0 1 20412
box -48 -56 432 834
use sg13g2_buf_1  _800_
timestamp 1676381911
transform 1 0 19968 0 -1 18900
box -48 -56 432 834
use sg13g2_buf_1  _801_
timestamp 1676381911
transform 1 0 18912 0 1 18900
box -48 -56 432 834
use sg13g2_buf_1  _802_
timestamp 1676381911
transform 1 0 19584 0 -1 18900
box -48 -56 432 834
use sg13g2_buf_1  _803_
timestamp 1676381911
transform 1 0 19680 0 1 18900
box -48 -56 432 834
use sg13g2_buf_1  _804_
timestamp 1676381911
transform 1 0 19872 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  _805_
timestamp 1676381911
transform 1 0 19296 0 1 18900
box -48 -56 432 834
use sg13g2_buf_1  _806_
timestamp 1676381911
transform 1 0 19776 0 -1 20412
box -48 -56 432 834
use sg13g2_buf_1  _807_
timestamp 1676381911
transform 1 0 19392 0 1 20412
box -48 -56 432 834
use sg13g2_buf_1  _808_
timestamp 1676381911
transform 1 0 19584 0 1 24948
box -48 -56 432 834
use sg13g2_buf_1  _809_
timestamp 1676381911
transform 1 0 18912 0 -1 21924
box -48 -56 432 834
use sg13g2_buf_1  _810_
timestamp 1676381911
transform 1 0 18912 0 1 21924
box -48 -56 432 834
use sg13g2_buf_1  _811_
timestamp 1676381911
transform 1 0 19872 0 -1 23436
box -48 -56 432 834
use sg13g2_buf_1  _812_
timestamp 1676381911
transform 1 0 19296 0 1 21924
box -48 -56 432 834
use sg13g2_buf_1  _813_
timestamp 1676381911
transform 1 0 19680 0 -1 26460
box -48 -56 432 834
use sg13g2_buf_1  _814_
timestamp 1676381911
transform 1 0 19968 0 -1 30996
box -48 -56 432 834
use sg13g2_buf_1  _815_
timestamp 1676381911
transform 1 0 18528 0 1 34020
box -48 -56 432 834
use sg13g2_buf_1  _816_
timestamp 1676381911
transform 1 0 18144 0 -1 34020
box -48 -56 432 834
use sg13g2_buf_1  _817_
timestamp 1676381911
transform 1 0 18912 0 -1 37044
box -48 -56 432 834
use sg13g2_buf_1  _818_
timestamp 1676381911
transform 1 0 19680 0 -1 34020
box -48 -56 432 834
use sg13g2_buf_1  _819_
timestamp 1676381911
transform 1 0 18528 0 -1 34020
box -48 -56 432 834
use sg13g2_buf_1  _820_
timestamp 1676381911
transform 1 0 16032 0 1 29484
box -48 -56 432 834
use sg13g2_buf_1  _821_
timestamp 1676381911
transform 1 0 19296 0 1 32508
box -48 -56 432 834
use sg13g2_buf_1  _822_
timestamp 1676381911
transform 1 0 19680 0 1 32508
box -48 -56 432 834
use sg13g2_buf_1  _823_
timestamp 1676381911
transform 1 0 19680 0 -1 37044
box -48 -56 432 834
use sg13g2_buf_1  _824_
timestamp 1676381911
transform 1 0 19296 0 -1 34020
box -48 -56 432 834
use sg13g2_buf_1  _825_
timestamp 1676381911
transform 1 0 18912 0 -1 34020
box -48 -56 432 834
use sg13g2_buf_1  _826_
timestamp 1676381911
transform 1 0 19584 0 1 38556
box -48 -56 432 834
use sg13g2_buf_1  _827_
timestamp 1676381911
transform 1 0 19296 0 -1 24948
box -48 -56 432 834
use sg13g2_buf_1  _828_
timestamp 1676381911
transform 1 0 19680 0 1 21924
box -48 -56 432 834
use sg13g2_buf_1  _829_
timestamp 1676381911
transform 1 0 19680 0 -1 24948
box -48 -56 432 834
use sg13g2_buf_1  _830_
timestamp 1676381911
transform 1 0 19680 0 -1 32508
box -48 -56 432 834
use sg13g2_buf_1  _831_
timestamp 1676381911
transform 1 0 18912 0 -1 24948
box -48 -56 432 834
use sg13g2_buf_1  _832_
timestamp 1676381911
transform 1 0 19968 0 1 24948
box -48 -56 432 834
use sg13g2_buf_1  _833_
timestamp 1676381911
transform 1 0 19296 0 -1 26460
box -48 -56 432 834
use sg13g2_buf_1  _834_
timestamp 1676381911
transform 1 0 18528 0 -1 24948
box -48 -56 432 834
use sg13g2_buf_1  _835_
timestamp 1676381911
transform 1 0 19872 0 -1 27972
box -48 -56 432 834
use sg13g2_buf_1  _836_
timestamp 1676381911
transform 1 0 19392 0 1 27972
box -48 -56 432 834
use sg13g2_buf_1  _837_
timestamp 1676381911
transform 1 0 19776 0 1 27972
box -48 -56 432 834
use sg13g2_buf_1  _838_
timestamp 1676381911
transform 1 0 16992 0 1 27972
box -48 -56 432 834
use sg13g2_buf_1  _839_
timestamp 1676381911
transform 1 0 19296 0 1 29484
box -48 -56 432 834
use sg13g2_buf_1  _840_
timestamp 1676381911
transform 1 0 19968 0 1 30996
box -48 -56 432 834
use sg13g2_buf_1  _841_
timestamp 1676381911
transform 1 0 19680 0 1 29484
box -48 -56 432 834
use sg13g2_buf_1  _842_
timestamp 1676381911
transform 1 0 19296 0 -1 32508
box -48 -56 432 834
use sg13g2_buf_1  _843_
timestamp 1676381911
transform 1 0 19296 0 1 34020
box -48 -56 432 834
use sg13g2_buf_1  _844_
timestamp 1676381911
transform 1 0 16992 0 -1 32508
box -48 -56 432 834
use sg13g2_buf_1  _845_
timestamp 1676381911
transform 1 0 19680 0 1 34020
box -48 -56 432 834
use sg13g2_buf_1  _846_
timestamp 1676381911
transform 1 0 18912 0 1 34020
box -48 -56 432 834
use sg13g2_buf_1  _847_
timestamp 1676381911
transform 1 0 19392 0 -1 35532
box -48 -56 432 834
use sg13g2_buf_1  _848_
timestamp 1676381911
transform 1 0 19776 0 -1 35532
box -48 -56 432 834
use sg13g2_buf_1  _849_
timestamp 1676381911
transform 1 0 19872 0 1 35532
box -48 -56 432 834
use sg13g2_buf_1  _850_
timestamp 1676381911
transform 1 0 19296 0 -1 37044
box -48 -56 432 834
use sg13g2_buf_1  _851_
timestamp 1676381911
transform 1 0 16992 0 -1 35532
box -48 -56 432 834
use sg13g2_buf_1  _852_
timestamp 1676381911
transform 1 0 19584 0 1 37044
box -48 -56 432 834
use sg13g2_buf_1  _853_
timestamp 1676381911
transform 1 0 19968 0 1 37044
box -48 -56 432 834
use sg13g2_buf_1  _854_
timestamp 1676381911
transform 1 0 19296 0 -1 38556
box -48 -56 432 834
use sg13g2_buf_1  _855_
timestamp 1676381911
transform 1 0 19680 0 -1 38556
box -48 -56 432 834
use sg13g2_buf_1  _856_
timestamp 1676381911
transform 1 0 18912 0 -1 38556
box -48 -56 432 834
use sg13g2_buf_1  _857_
timestamp 1676381911
transform 1 0 11328 0 1 35532
box -48 -56 432 834
use sg13g2_buf_1  _858_
timestamp 1676381911
transform 1 0 17184 0 1 37044
box -48 -56 432 834
use sg13g2_buf_1  _859_
timestamp 1676381911
transform 1 0 19968 0 1 38556
box -48 -56 432 834
use sg13g2_buf_1  _860_
timestamp 1676381911
transform 1 0 19200 0 1 38556
box -48 -56 432 834
use sg13g2_buf_1  _861_
timestamp 1676381911
transform 1 0 12384 0 -1 38556
box -48 -56 432 834
use sg13g2_buf_1  _862_
timestamp 1676381911
transform 1 0 19680 0 -1 40068
box -48 -56 432 834
use sg13g2_buf_1  _863_
timestamp 1676381911
transform 1 0 16608 0 -1 32508
box -48 -56 432 834
use sg13g2_buf_1  _864_
timestamp 1676381911
transform 1 0 19296 0 -1 40068
box -48 -56 432 834
use sg13g2_buf_1  _865_
timestamp 1676381911
transform 1 0 12000 0 1 38556
box -48 -56 432 834
use sg13g2_buf_1  _866_
timestamp 1676381911
transform 1 0 14784 0 -1 37044
box -48 -56 432 834
use sg13g2_buf_1  _867_
timestamp 1676381911
transform 1 0 16224 0 -1 35532
box -48 -56 432 834
use sg13g2_buf_1  _868_
timestamp 1676381911
transform 1 0 19680 0 -1 41580
box -48 -56 432 834
use sg13g2_buf_1  _869_
timestamp 1676381911
transform 1 0 16800 0 1 38556
box -48 -56 432 834
use sg13g2_buf_1  _870_
timestamp 1676381911
transform 1 0 12000 0 -1 38556
box -48 -56 432 834
use sg13g2_buf_1  _871_
timestamp 1676381911
transform 1 0 15168 0 1 37044
box -48 -56 432 834
use sg13g2_buf_1  _872_
timestamp 1676381911
transform 1 0 17184 0 1 38556
box -48 -56 432 834
use sg13g2_buf_1  _873_
timestamp 1676381911
transform 1 0 12864 0 -1 40068
box -48 -56 432 834
use sg13g2_buf_1  _874_
timestamp 1676381911
transform 1 0 16608 0 -1 35532
box -48 -56 432 834
use sg13g2_buf_1  _875_
timestamp 1676381911
transform -1 0 18912 0 -1 41580
box -48 -56 432 834
use sg13g2_buf_1  _876_
timestamp 1676381911
transform -1 0 19296 0 -1 41580
box -48 -56 432 834
use sg13g2_buf_1  _877_
timestamp 1676381911
transform 1 0 15648 0 1 23436
box -48 -56 432 834
use sg13g2_buf_1  _878_
timestamp 1676381911
transform -1 0 17952 0 1 38556
box -48 -56 432 834
use sg13g2_buf_1  _879_
timestamp 1676381911
transform -1 0 18816 0 1 38556
box -48 -56 432 834
use sg13g2_buf_1  _880_
timestamp 1676381911
transform 1 0 16416 0 1 29484
box -48 -56 432 834
use sg13g2_buf_1  _881_
timestamp 1676381911
transform 1 0 13152 0 -1 38556
box -48 -56 432 834
use sg13g2_buf_1  _882_
timestamp 1676381911
transform -1 0 19392 0 1 40068
box -48 -56 432 834
use sg13g2_buf_1  _883_
timestamp 1676381911
transform 1 0 14400 0 -1 37044
box -48 -56 432 834
use sg13g2_buf_1  _884_
timestamp 1676381911
transform -1 0 18912 0 -1 40068
box -48 -56 432 834
use sg13g2_buf_1  _885_
timestamp 1676381911
transform 1 0 15840 0 -1 35532
box -48 -56 432 834
use sg13g2_buf_1  _886_
timestamp 1676381911
transform -1 0 19296 0 -1 40068
box -48 -56 432 834
use sg13g2_buf_1  _887_
timestamp 1676381911
transform -1 0 20160 0 1 40068
box -48 -56 432 834
use sg13g2_buf_1  _888_
timestamp 1676381911
transform -1 0 18624 0 1 40068
box -48 -56 432 834
use sg13g2_buf_1  _889_
timestamp 1676381911
transform 1 0 15456 0 -1 34020
box -48 -56 432 834
use sg13g2_buf_1  _890_
timestamp 1676381911
transform 1 0 12768 0 -1 38556
box -48 -56 432 834
use sg13g2_buf_1  _891_
timestamp 1676381911
transform -1 0 19776 0 1 40068
box -48 -56 432 834
use sg13g2_buf_1  _892_
timestamp 1676381911
transform 1 0 17184 0 1 40068
box -48 -56 432 834
use sg13g2_buf_1  _893_
timestamp 1676381911
transform 1 0 18144 0 -1 40068
box -48 -56 432 834
use sg13g2_buf_1  _894_
timestamp 1676381911
transform 1 0 14400 0 1 38556
box -48 -56 432 834
use sg13g2_buf_1  _895_
timestamp 1676381911
transform 1 0 1344 0 -1 34020
box -48 -56 432 834
use sg13g2_buf_1  _896_
timestamp 1676381911
transform 1 0 1248 0 1 35532
box -48 -56 432 834
use sg13g2_buf_1  _897_
timestamp 1676381911
transform 1 0 1344 0 -1 35532
box -48 -56 432 834
use sg13g2_buf_1  _898_
timestamp 1676381911
transform 1 0 1248 0 -1 37044
box -48 -56 432 834
use sg13g2_buf_1  _899_
timestamp 1676381911
transform -1 0 14016 0 1 40068
box -48 -56 432 834
use sg13g2_buf_1  _900_
timestamp 1676381911
transform -1 0 3264 0 1 34020
box -48 -56 432 834
use sg13g2_buf_1  _901_
timestamp 1676381911
transform 1 0 1152 0 -1 38556
box -48 -56 432 834
use sg13g2_buf_1  _902_
timestamp 1676381911
transform 1 0 1152 0 1 37044
box -48 -56 432 834
use sg13g2_buf_1  _903_
timestamp 1676381911
transform -1 0 3744 0 1 35532
box -48 -56 432 834
use sg13g2_buf_1  _904_
timestamp 1676381911
transform 1 0 1632 0 -1 37044
box -48 -56 432 834
use sg13g2_buf_1  _905_
timestamp 1676381911
transform 1 0 1152 0 -1 40068
box -48 -56 432 834
use sg13g2_buf_1  _906_
timestamp 1676381911
transform -1 0 19680 0 -1 41580
box -48 -56 432 834
use sg13g2_buf_1  _907_
timestamp 1676381911
transform 1 0 1632 0 1 32508
box -48 -56 432 834
use sg13g2_buf_1  _908_
timestamp 1676381911
transform 1 0 1536 0 1 37044
box -48 -56 432 834
use sg13g2_buf_1  _909_
timestamp 1676381911
transform 1 0 1248 0 1 32508
box -48 -56 432 834
use sg13g2_buf_1  _910_
timestamp 1676381911
transform 1 0 4416 0 -1 37044
box -48 -56 432 834
use sg13g2_buf_1  _911_
timestamp 1676381911
transform 1 0 1440 0 1 40068
box -48 -56 432 834
use sg13g2_buf_1  _912_
timestamp 1676381911
transform 1 0 4416 0 1 37044
box -48 -56 432 834
use sg13g2_buf_1  _913_
timestamp 1676381911
transform 1 0 1536 0 -1 38556
box -48 -56 432 834
use sg13g2_buf_1  _914_
timestamp 1676381911
transform 1 0 4800 0 1 37044
box -48 -56 432 834
use sg13g2_buf_1  _915_
timestamp 1676381911
transform 1 0 1920 0 -1 38556
box -48 -56 432 834
use sg13g2_buf_1  _916_
timestamp 1676381911
transform 1 0 2112 0 -1 37044
box -48 -56 432 834
use sg13g2_buf_1  _917_
timestamp 1676381911
transform 1 0 5184 0 1 37044
box -48 -56 432 834
use sg13g2_buf_1  _918_
timestamp 1676381911
transform 1 0 3744 0 1 35532
box -48 -56 432 834
use sg13g2_buf_1  _919_
timestamp 1676381911
transform -1 0 7584 0 -1 38556
box -48 -56 432 834
use sg13g2_buf_1  _920_
timestamp 1676381911
transform -1 0 7200 0 -1 38556
box -48 -56 432 834
use sg13g2_buf_1  _921_
timestamp 1676381911
transform 1 0 1248 0 1 38556
box -48 -56 432 834
use sg13g2_buf_1  _922_
timestamp 1676381911
transform 1 0 3264 0 -1 40068
box -48 -56 432 834
use sg13g2_buf_1  _923_
timestamp 1676381911
transform 1 0 6816 0 -1 37044
box -48 -56 432 834
use sg13g2_buf_1  _924_
timestamp 1676381911
transform 1 0 3648 0 1 40068
box -48 -56 432 834
use sg13g2_buf_1  _925_
timestamp 1676381911
transform -1 0 10560 0 -1 40068
box -48 -56 432 834
use sg13g2_buf_1  _926_
timestamp 1676381911
transform 1 0 5952 0 1 40068
box -48 -56 432 834
use sg13g2_buf_1  _927_
timestamp 1676381911
transform -1 0 19008 0 1 40068
box -48 -56 432 834
use sg13g2_buf_1  _928_
timestamp 1676381911
transform 1 0 4128 0 1 38556
box -48 -56 432 834
use sg13g2_buf_1  _929_
timestamp 1676381911
transform 1 0 7968 0 -1 41580
box -48 -56 432 834
use sg13g2_buf_1  _930_
timestamp 1676381911
transform -1 0 15936 0 1 40068
box -48 -56 432 834
use sg13g2_buf_1  _931_
timestamp 1676381911
transform 1 0 6528 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _932_
timestamp 1676381911
transform 1 0 2880 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _933_
timestamp 1676381911
transform 1 0 4320 0 1 756
box -48 -56 432 834
use sg13g2_buf_1  _934_
timestamp 1676381911
transform 1 0 7968 0 1 756
box -48 -56 432 834
use sg13g2_buf_1  _935_
timestamp 1676381911
transform 1 0 8352 0 1 756
box -48 -56 432 834
use sg13g2_buf_1  _936_
timestamp 1676381911
transform 1 0 5376 0 1 2268
box -48 -56 432 834
use sg13g2_buf_1  _937_
timestamp 1676381911
transform -1 0 11904 0 1 756
box -48 -56 432 834
use sg13g2_buf_1  _938_
timestamp 1676381911
transform 1 0 9504 0 1 756
box -48 -56 432 834
use sg13g2_buf_1  _939_
timestamp 1676381911
transform -1 0 11040 0 1 756
box -48 -56 432 834
use sg13g2_buf_1  _940_
timestamp 1676381911
transform 1 0 7584 0 1 756
box -48 -56 432 834
use sg13g2_buf_1  _941_
timestamp 1676381911
transform 1 0 2304 0 1 756
box -48 -56 432 834
use sg13g2_buf_1  _942_
timestamp 1676381911
transform -1 0 14112 0 1 2268
box -48 -56 432 834
use sg13g2_buf_1  _943_
timestamp 1676381911
transform 1 0 8736 0 1 756
box -48 -56 432 834
use sg13g2_buf_1  _944_
timestamp 1676381911
transform 1 0 9120 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _945_
timestamp 1676381911
transform 1 0 10272 0 1 756
box -48 -56 432 834
use sg13g2_buf_1  _946_
timestamp 1676381911
transform 1 0 9888 0 1 756
box -48 -56 432 834
use sg13g2_buf_1  _947_
timestamp 1676381911
transform 1 0 10272 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _948_
timestamp 1676381911
transform 1 0 11136 0 1 756
box -48 -56 432 834
use sg13g2_buf_1  _949_
timestamp 1676381911
transform 1 0 10656 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _950_
timestamp 1676381911
transform 1 0 11040 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _951_
timestamp 1676381911
transform -1 0 14400 0 1 40068
box -48 -56 432 834
use sg13g2_buf_1  _952_
timestamp 1676381911
transform -1 0 14784 0 1 40068
box -48 -56 432 834
use sg13g2_buf_1  _953_
timestamp 1676381911
transform -1 0 15552 0 -1 41580
box -48 -56 432 834
use sg13g2_buf_1  _954_
timestamp 1676381911
transform -1 0 15168 0 1 40068
box -48 -56 432 834
use sg13g2_buf_1  _955_
timestamp 1676381911
transform -1 0 15936 0 -1 41580
box -48 -56 432 834
use sg13g2_buf_1  _956_
timestamp 1676381911
transform -1 0 15552 0 1 40068
box -48 -56 432 834
use sg13g2_buf_1  _957_
timestamp 1676381911
transform -1 0 16320 0 -1 41580
box -48 -56 432 834
use sg13g2_buf_1  _958_
timestamp 1676381911
transform -1 0 16320 0 1 40068
box -48 -56 432 834
use sg13g2_buf_1  _959_
timestamp 1676381911
transform -1 0 16704 0 1 40068
box -48 -56 432 834
use sg13g2_buf_1  _960_
timestamp 1676381911
transform -1 0 17088 0 1 40068
box -48 -56 432 834
use sg13g2_buf_1  _961_
timestamp 1676381911
transform -1 0 17184 0 -1 40068
box -48 -56 432 834
use sg13g2_buf_1  _962_
timestamp 1676381911
transform -1 0 17952 0 1 40068
box -48 -56 432 834
use sg13g2_buf_1  _963_
timestamp 1676381911
transform -1 0 15648 0 1 756
box -48 -56 432 834
use sg13g2_buf_1  _964_
timestamp 1676381911
transform 1 0 14112 0 1 2268
box -48 -56 432 834
use sg13g2_buf_1  _965_
timestamp 1676381911
transform 1 0 14784 0 1 756
box -48 -56 432 834
use sg13g2_buf_1  _966_
timestamp 1676381911
transform -1 0 16128 0 -1 3780
box -48 -56 432 834
use sg13g2_buf_1  _967_
timestamp 1676381911
transform -1 0 17856 0 -1 40068
box -48 -56 432 834
use sg13g2_antennanp  ANTENNA_1
timestamp 1679999689
transform 1 0 20064 0 -1 40068
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_2
timestamp 1679999689
transform 1 0 20064 0 -1 38556
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_3
timestamp 1679999689
transform -1 0 18240 0 1 40068
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_4
timestamp 1679999689
transform -1 0 18144 0 -1 40068
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_5
timestamp 1679999689
transform 1 0 9696 0 1 40068
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_6
timestamp 1679999689
transform -1 0 10848 0 -1 40068
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_7
timestamp 1679999689
transform 1 0 4416 0 1 35532
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_8
timestamp 1679999689
transform 1 0 4896 0 1 3780
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_9
timestamp 1679999689
transform -1 0 4416 0 -1 37044
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_10
timestamp 1679999689
transform -1 0 1440 0 1 40068
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_11
timestamp 1679999689
transform 1 0 9504 0 -1 38556
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_12
timestamp 1679999689
transform -1 0 1440 0 -1 41580
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_13
timestamp 1679999689
transform 1 0 7200 0 1 37044
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_14
timestamp 1679999689
transform 1 0 18912 0 1 38556
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_15
timestamp 1679999689
transform 1 0 18240 0 -1 41580
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_16
timestamp 1679999689
transform 1 0 17184 0 -1 40068
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_17
timestamp 1679999689
transform 1 0 18144 0 1 38556
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_18
timestamp 1679999689
transform -1 0 6816 0 -1 37044
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_19
timestamp 1679999689
transform 1 0 3648 0 -1 40068
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_20
timestamp 1679999689
transform 1 0 5952 0 -1 40068
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_21
timestamp 1679999689
transform 1 0 1920 0 1 37044
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_22
timestamp 1679999689
transform 1 0 2112 0 1 35532
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_23
timestamp 1679999689
transform -1 0 4032 0 -1 37044
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_24
timestamp 1679999689
transform -1 0 4032 0 1 34020
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_25
timestamp 1679999689
transform -1 0 9408 0 1 756
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_26
timestamp 1679999689
transform -1 0 4032 0 -1 34020
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_27
timestamp 1679999689
transform 1 0 9120 0 1 2268
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_28
timestamp 1679999689
transform -1 0 15456 0 -1 34020
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_29
timestamp 1679999689
transform 1 0 3264 0 1 38556
box -48 -56 336 834
use sg13g2_buf_8  clkbuf_0_UserCLK
timestamp 1676451365
transform -1 0 12960 0 1 32508
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_1_0__f_UserCLK
timestamp 1676451365
transform -1 0 9984 0 1 29484
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_1_1__f_UserCLK
timestamp 1676451365
transform 1 0 11712 0 1 35532
box -48 -56 1296 834
use sg13g2_decap_8  FILLER_0_0
timestamp 1679581782
transform 1 0 1152 0 1 756
box -48 -56 720 834
use sg13g2_decap_4  FILLER_0_7
timestamp 1679577901
transform 1 0 1824 0 1 756
box -48 -56 432 834
use sg13g2_fill_1  FILLER_0_11
timestamp 1677579658
transform 1 0 2208 0 1 756
box -48 -56 144 834
use sg13g2_fill_2  FILLER_0_60
timestamp 1677580104
transform 1 0 6912 0 1 756
box -48 -56 240 834
use sg13g2_fill_1  FILLER_0_86
timestamp 1677579658
transform 1 0 9408 0 1 756
box -48 -56 144 834
use sg13g2_fill_1  FILLER_0_103
timestamp 1677579658
transform 1 0 11040 0 1 756
box -48 -56 144 834
use sg13g2_decap_8  FILLER_0_112
timestamp 1679581782
transform 1 0 11904 0 1 756
box -48 -56 720 834
use sg13g2_decap_4  FILLER_0_119
timestamp 1679577901
transform 1 0 12576 0 1 756
box -48 -56 432 834
use sg13g2_fill_2  FILLER_0_123
timestamp 1677580104
transform 1 0 12960 0 1 756
box -48 -56 240 834
use sg13g2_fill_1  FILLER_0_146
timestamp 1677579658
transform 1 0 15168 0 1 756
box -48 -56 144 834
use sg13g2_fill_2  FILLER_0_174
timestamp 1677580104
transform 1 0 17856 0 1 756
box -48 -56 240 834
use sg13g2_decap_8  FILLER_0_193
timestamp 1679581782
transform 1 0 19680 0 1 756
box -48 -56 720 834
use sg13g2_fill_1  FILLER_1_0
timestamp 1677579658
transform 1 0 1152 0 -1 2268
box -48 -56 144 834
use sg13g2_fill_2  FILLER_1_65
timestamp 1677580104
transform 1 0 7392 0 -1 2268
box -48 -56 240 834
use sg13g2_fill_1  FILLER_1_82
timestamp 1677579658
transform 1 0 9024 0 -1 2268
box -48 -56 144 834
use sg13g2_fill_2  FILLER_1_87
timestamp 1677580104
transform 1 0 9504 0 -1 2268
box -48 -56 240 834
use sg13g2_fill_1  FILLER_1_94
timestamp 1677579658
transform 1 0 10176 0 -1 2268
box -48 -56 144 834
use sg13g2_fill_1  FILLER_1_145
timestamp 1677579658
transform 1 0 15072 0 -1 2268
box -48 -56 144 834
use sg13g2_fill_1  FILLER_1_178
timestamp 1677579658
transform 1 0 18240 0 -1 2268
box -48 -56 144 834
use sg13g2_decap_4  FILLER_1_196
timestamp 1679577901
transform 1 0 19968 0 -1 2268
box -48 -56 432 834
use sg13g2_decap_4  FILLER_2_0
timestamp 1679577901
transform 1 0 1152 0 1 2268
box -48 -56 432 834
use sg13g2_fill_2  FILLER_2_25
timestamp 1677580104
transform 1 0 3552 0 1 2268
box -48 -56 240 834
use sg13g2_fill_1  FILLER_2_66
timestamp 1677579658
transform 1 0 7488 0 1 2268
box -48 -56 144 834
use sg13g2_fill_1  FILLER_2_77
timestamp 1677579658
transform 1 0 8544 0 1 2268
box -48 -56 144 834
use sg13g2_decap_8  FILLER_2_121
timestamp 1679581782
transform 1 0 12768 0 1 2268
box -48 -56 720 834
use sg13g2_fill_2  FILLER_2_128
timestamp 1677580104
transform 1 0 13440 0 1 2268
box -48 -56 240 834
use sg13g2_fill_1  FILLER_2_130
timestamp 1677579658
transform 1 0 13632 0 1 2268
box -48 -56 144 834
use sg13g2_fill_2  FILLER_2_139
timestamp 1677580104
transform 1 0 14496 0 1 2268
box -48 -56 240 834
use sg13g2_fill_2  FILLER_2_178
timestamp 1677580104
transform 1 0 18240 0 1 2268
box -48 -56 240 834
use sg13g2_fill_2  FILLER_2_197
timestamp 1677580104
transform 1 0 20064 0 1 2268
box -48 -56 240 834
use sg13g2_fill_1  FILLER_2_199
timestamp 1677579658
transform 1 0 20256 0 1 2268
box -48 -56 144 834
use sg13g2_decap_8  FILLER_3_0
timestamp 1679581782
transform 1 0 1152 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_4  FILLER_3_7
timestamp 1679577901
transform 1 0 1824 0 -1 3780
box -48 -56 432 834
use sg13g2_fill_2  FILLER_3_11
timestamp 1677580104
transform 1 0 2208 0 -1 3780
box -48 -56 240 834
use sg13g2_fill_1  FILLER_3_34
timestamp 1677579658
transform 1 0 4416 0 -1 3780
box -48 -56 144 834
use sg13g2_fill_1  FILLER_3_59
timestamp 1677579658
transform 1 0 6816 0 -1 3780
box -48 -56 144 834
use sg13g2_decap_4  FILLER_3_100
timestamp 1679577901
transform 1 0 10752 0 -1 3780
box -48 -56 432 834
use sg13g2_decap_8  FILLER_3_121
timestamp 1679581782
transform 1 0 12768 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_128
timestamp 1679581782
transform 1 0 13440 0 -1 3780
box -48 -56 720 834
use sg13g2_fill_2  FILLER_3_174
timestamp 1677580104
transform 1 0 17856 0 -1 3780
box -48 -56 240 834
use sg13g2_fill_2  FILLER_3_198
timestamp 1677580104
transform 1 0 20160 0 -1 3780
box -48 -56 240 834
use sg13g2_fill_1  FILLER_4_80
timestamp 1677579658
transform 1 0 8832 0 1 3780
box -48 -56 144 834
use sg13g2_decap_8  FILLER_4_98
timestamp 1679581782
transform 1 0 10560 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_143
timestamp 1679581782
transform 1 0 14880 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_150
timestamp 1679581782
transform 1 0 15552 0 1 3780
box -48 -56 720 834
use sg13g2_decap_4  FILLER_4_173
timestamp 1679577901
transform 1 0 17760 0 1 3780
box -48 -56 432 834
use sg13g2_fill_2  FILLER_4_177
timestamp 1677580104
transform 1 0 18144 0 1 3780
box -48 -56 240 834
use sg13g2_fill_2  FILLER_5_39
timestamp 1677580104
transform 1 0 4896 0 -1 5292
box -48 -56 240 834
use sg13g2_fill_1  FILLER_5_41
timestamp 1677579658
transform 1 0 5088 0 -1 5292
box -48 -56 144 834
use sg13g2_fill_1  FILLER_5_59
timestamp 1677579658
transform 1 0 6816 0 -1 5292
box -48 -56 144 834
use sg13g2_decap_8  FILLER_5_81
timestamp 1679581782
transform 1 0 8928 0 -1 5292
box -48 -56 720 834
use sg13g2_fill_1  FILLER_5_88
timestamp 1677579658
transform 1 0 9600 0 -1 5292
box -48 -56 144 834
use sg13g2_decap_4  FILLER_5_174
timestamp 1679577901
transform 1 0 17856 0 -1 5292
box -48 -56 432 834
use sg13g2_fill_2  FILLER_5_183
timestamp 1677580104
transform 1 0 18720 0 -1 5292
box -48 -56 240 834
use sg13g2_fill_1  FILLER_5_185
timestamp 1677579658
transform 1 0 18912 0 -1 5292
box -48 -56 144 834
use sg13g2_decap_4  FILLER_5_196
timestamp 1679577901
transform 1 0 19968 0 -1 5292
box -48 -56 432 834
use sg13g2_fill_2  FILLER_6_0
timestamp 1677580104
transform 1 0 1152 0 1 5292
box -48 -56 240 834
use sg13g2_fill_1  FILLER_6_2
timestamp 1677579658
transform 1 0 1344 0 1 5292
box -48 -56 144 834
use sg13g2_fill_2  FILLER_6_58
timestamp 1677580104
transform 1 0 6720 0 1 5292
box -48 -56 240 834
use sg13g2_decap_8  FILLER_6_98
timestamp 1679581782
transform 1 0 10560 0 1 5292
box -48 -56 720 834
use sg13g2_fill_1  FILLER_6_105
timestamp 1677579658
transform 1 0 11232 0 1 5292
box -48 -56 144 834
use sg13g2_fill_2  FILLER_6_123
timestamp 1677580104
transform 1 0 12960 0 1 5292
box -48 -56 240 834
use sg13g2_fill_1  FILLER_6_142
timestamp 1677579658
transform 1 0 14784 0 1 5292
box -48 -56 144 834
use sg13g2_fill_2  FILLER_6_176
timestamp 1677580104
transform 1 0 18048 0 1 5292
box -48 -56 240 834
use sg13g2_fill_1  FILLER_7_17
timestamp 1677579658
transform 1 0 2784 0 -1 6804
box -48 -56 144 834
use sg13g2_decap_8  FILLER_7_64
timestamp 1679581782
transform 1 0 7296 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_4  FILLER_7_71
timestamp 1679577901
transform 1 0 7968 0 -1 6804
box -48 -56 432 834
use sg13g2_fill_2  FILLER_7_75
timestamp 1677580104
transform 1 0 8352 0 -1 6804
box -48 -56 240 834
use sg13g2_decap_4  FILLER_7_98
timestamp 1679577901
transform 1 0 10560 0 -1 6804
box -48 -56 432 834
use sg13g2_fill_2  FILLER_7_102
timestamp 1677580104
transform 1 0 10944 0 -1 6804
box -48 -56 240 834
use sg13g2_decap_8  FILLER_7_142
timestamp 1679581782
transform 1 0 14784 0 -1 6804
box -48 -56 720 834
use sg13g2_fill_2  FILLER_7_149
timestamp 1677580104
transform 1 0 15456 0 -1 6804
box -48 -56 240 834
use sg13g2_fill_2  FILLER_7_168
timestamp 1677580104
transform 1 0 17280 0 -1 6804
box -48 -56 240 834
use sg13g2_fill_2  FILLER_7_198
timestamp 1677580104
transform 1 0 20160 0 -1 6804
box -48 -56 240 834
use sg13g2_decap_8  FILLER_8_39
timestamp 1679581782
transform 1 0 4896 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_46
timestamp 1679581782
transform 1 0 5568 0 1 6804
box -48 -56 720 834
use sg13g2_fill_1  FILLER_8_53
timestamp 1677579658
transform 1 0 6240 0 1 6804
box -48 -56 144 834
use sg13g2_fill_2  FILLER_8_71
timestamp 1677580104
transform 1 0 7968 0 1 6804
box -48 -56 240 834
use sg13g2_fill_1  FILLER_8_73
timestamp 1677579658
transform 1 0 8160 0 1 6804
box -48 -56 144 834
use sg13g2_decap_8  FILLER_8_129
timestamp 1679581782
transform 1 0 13536 0 1 6804
box -48 -56 720 834
use sg13g2_decap_4  FILLER_8_195
timestamp 1679577901
transform 1 0 19872 0 1 6804
box -48 -56 432 834
use sg13g2_fill_1  FILLER_8_199
timestamp 1677579658
transform 1 0 20256 0 1 6804
box -48 -56 144 834
use sg13g2_decap_8  FILLER_9_0
timestamp 1679581782
transform 1 0 1152 0 -1 8316
box -48 -56 720 834
use sg13g2_fill_1  FILLER_9_35
timestamp 1677579658
transform 1 0 4512 0 -1 8316
box -48 -56 144 834
use sg13g2_fill_1  FILLER_9_74
timestamp 1677579658
transform 1 0 8256 0 -1 8316
box -48 -56 144 834
use sg13g2_decap_4  FILLER_9_126
timestamp 1679577901
transform 1 0 13248 0 -1 8316
box -48 -56 432 834
use sg13g2_fill_2  FILLER_9_130
timestamp 1677580104
transform 1 0 13632 0 -1 8316
box -48 -56 240 834
use sg13g2_decap_8  FILLER_9_166
timestamp 1679581782
transform 1 0 17088 0 -1 8316
box -48 -56 720 834
use sg13g2_fill_2  FILLER_9_173
timestamp 1677580104
transform 1 0 17760 0 -1 8316
box -48 -56 240 834
use sg13g2_fill_2  FILLER_9_183
timestamp 1677580104
transform 1 0 18720 0 -1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_9_185
timestamp 1677579658
transform 1 0 18912 0 -1 8316
box -48 -56 144 834
use sg13g2_decap_4  FILLER_9_196
timestamp 1679577901
transform 1 0 19968 0 -1 8316
box -48 -56 432 834
use sg13g2_fill_2  FILLER_10_17
timestamp 1677580104
transform 1 0 2784 0 1 8316
box -48 -56 240 834
use sg13g2_decap_8  FILLER_10_39
timestamp 1679581782
transform 1 0 4896 0 1 8316
box -48 -56 720 834
use sg13g2_fill_1  FILLER_10_46
timestamp 1677579658
transform 1 0 5568 0 1 8316
box -48 -56 144 834
use sg13g2_decap_8  FILLER_10_64
timestamp 1679581782
transform 1 0 7296 0 1 8316
box -48 -56 720 834
use sg13g2_fill_2  FILLER_10_71
timestamp 1677580104
transform 1 0 7968 0 1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_10_73
timestamp 1677579658
transform 1 0 8160 0 1 8316
box -48 -56 144 834
use sg13g2_decap_8  FILLER_10_112
timestamp 1679581782
transform 1 0 11904 0 1 8316
box -48 -56 720 834
use sg13g2_decap_4  FILLER_10_119
timestamp 1679577901
transform 1 0 12576 0 1 8316
box -48 -56 432 834
use sg13g2_fill_1  FILLER_10_140
timestamp 1677579658
transform 1 0 14592 0 1 8316
box -48 -56 144 834
use sg13g2_fill_2  FILLER_10_154
timestamp 1677580104
transform 1 0 15936 0 1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_10_199
timestamp 1677579658
transform 1 0 20256 0 1 8316
box -48 -56 144 834
use sg13g2_fill_2  FILLER_11_0
timestamp 1677580104
transform 1 0 1152 0 -1 9828
box -48 -56 240 834
use sg13g2_fill_1  FILLER_11_2
timestamp 1677579658
transform 1 0 1344 0 -1 9828
box -48 -56 144 834
use sg13g2_fill_1  FILLER_11_20
timestamp 1677579658
transform 1 0 3072 0 -1 9828
box -48 -56 144 834
use sg13g2_fill_2  FILLER_11_28
timestamp 1677580104
transform 1 0 3840 0 -1 9828
box -48 -56 240 834
use sg13g2_fill_2  FILLER_11_85
timestamp 1677580104
transform 1 0 9312 0 -1 9828
box -48 -56 240 834
use sg13g2_fill_1  FILLER_11_87
timestamp 1677579658
transform 1 0 9504 0 -1 9828
box -48 -56 144 834
use sg13g2_decap_4  FILLER_11_100
timestamp 1679577901
transform 1 0 10752 0 -1 9828
box -48 -56 432 834
use sg13g2_fill_2  FILLER_11_162
timestamp 1677580104
transform 1 0 16704 0 -1 9828
box -48 -56 240 834
use sg13g2_decap_8  FILLER_12_38
timestamp 1679581782
transform 1 0 4800 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_45
timestamp 1679581782
transform 1 0 5472 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_52
timestamp 1679581782
transform 1 0 6144 0 1 9828
box -48 -56 720 834
use sg13g2_decap_4  FILLER_12_59
timestamp 1679577901
transform 1 0 6816 0 1 9828
box -48 -56 432 834
use sg13g2_fill_2  FILLER_12_63
timestamp 1677580104
transform 1 0 7200 0 1 9828
box -48 -56 240 834
use sg13g2_fill_2  FILLER_12_103
timestamp 1677580104
transform 1 0 11040 0 1 9828
box -48 -56 240 834
use sg13g2_fill_1  FILLER_12_105
timestamp 1677579658
transform 1 0 11232 0 1 9828
box -48 -56 144 834
use sg13g2_fill_2  FILLER_12_123
timestamp 1677580104
transform 1 0 12960 0 1 9828
box -48 -56 240 834
use sg13g2_decap_4  FILLER_12_163
timestamp 1679577901
transform 1 0 16800 0 1 9828
box -48 -56 432 834
use sg13g2_fill_2  FILLER_12_167
timestamp 1677580104
transform 1 0 17184 0 1 9828
box -48 -56 240 834
use sg13g2_decap_4  FILLER_12_196
timestamp 1679577901
transform 1 0 19968 0 1 9828
box -48 -56 432 834
use sg13g2_fill_2  FILLER_13_17
timestamp 1677580104
transform 1 0 2784 0 -1 11340
box -48 -56 240 834
use sg13g2_decap_4  FILLER_13_29
timestamp 1679577901
transform 1 0 3936 0 -1 11340
box -48 -56 432 834
use sg13g2_decap_4  FILLER_13_43
timestamp 1679577901
transform 1 0 5280 0 -1 11340
box -48 -56 432 834
use sg13g2_fill_1  FILLER_13_47
timestamp 1677579658
transform 1 0 5664 0 -1 11340
box -48 -56 144 834
use sg13g2_fill_2  FILLER_13_65
timestamp 1677580104
transform 1 0 7392 0 -1 11340
box -48 -56 240 834
use sg13g2_fill_1  FILLER_13_67
timestamp 1677579658
transform 1 0 7584 0 -1 11340
box -48 -56 144 834
use sg13g2_fill_2  FILLER_13_94
timestamp 1677580104
transform 1 0 10176 0 -1 11340
box -48 -56 240 834
use sg13g2_fill_1  FILLER_13_96
timestamp 1677579658
transform 1 0 10368 0 -1 11340
box -48 -56 144 834
use sg13g2_fill_2  FILLER_13_114
timestamp 1677580104
transform 1 0 12096 0 -1 11340
box -48 -56 240 834
use sg13g2_fill_1  FILLER_13_116
timestamp 1677579658
transform 1 0 12288 0 -1 11340
box -48 -56 144 834
use sg13g2_decap_8  FILLER_13_132
timestamp 1679581782
transform 1 0 13824 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_139
timestamp 1679581782
transform 1 0 14496 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_146
timestamp 1679581782
transform 1 0 15168 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_153
timestamp 1679581782
transform 1 0 15840 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_160
timestamp 1679581782
transform 1 0 16512 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_4  FILLER_13_167
timestamp 1679577901
transform 1 0 17184 0 -1 11340
box -48 -56 432 834
use sg13g2_fill_1  FILLER_13_171
timestamp 1677579658
transform 1 0 17568 0 -1 11340
box -48 -56 144 834
use sg13g2_fill_2  FILLER_13_198
timestamp 1677580104
transform 1 0 20160 0 -1 11340
box -48 -56 240 834
use sg13g2_decap_8  FILLER_14_17
timestamp 1679581782
transform 1 0 2784 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_29
timestamp 1679581782
transform 1 0 3936 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_36
timestamp 1679581782
transform 1 0 4608 0 1 11340
box -48 -56 720 834
use sg13g2_fill_1  FILLER_14_43
timestamp 1677579658
transform 1 0 5280 0 1 11340
box -48 -56 144 834
use sg13g2_fill_2  FILLER_14_141
timestamp 1677580104
transform 1 0 14688 0 1 11340
box -48 -56 240 834
use sg13g2_fill_1  FILLER_14_143
timestamp 1677579658
transform 1 0 14880 0 1 11340
box -48 -56 144 834
use sg13g2_fill_2  FILLER_14_161
timestamp 1677580104
transform 1 0 16608 0 1 11340
box -48 -56 240 834
use sg13g2_fill_1  FILLER_14_185
timestamp 1677579658
transform 1 0 18912 0 1 11340
box -48 -56 144 834
use sg13g2_fill_1  FILLER_14_199
timestamp 1677579658
transform 1 0 20256 0 1 11340
box -48 -56 144 834
use sg13g2_decap_8  FILLER_15_0
timestamp 1679581782
transform 1 0 1152 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_4  FILLER_15_7
timestamp 1679577901
transform 1 0 1824 0 -1 12852
box -48 -56 432 834
use sg13g2_fill_1  FILLER_15_66
timestamp 1677579658
transform 1 0 7488 0 -1 12852
box -48 -56 144 834
use sg13g2_decap_4  FILLER_15_94
timestamp 1679577901
transform 1 0 10176 0 -1 12852
box -48 -56 432 834
use sg13g2_fill_2  FILLER_15_98
timestamp 1677580104
transform 1 0 10560 0 -1 12852
box -48 -56 240 834
use sg13g2_decap_4  FILLER_15_117
timestamp 1679577901
transform 1 0 12384 0 -1 12852
box -48 -56 432 834
use sg13g2_fill_2  FILLER_15_128
timestamp 1677580104
transform 1 0 13440 0 -1 12852
box -48 -56 240 834
use sg13g2_fill_1  FILLER_15_130
timestamp 1677579658
transform 1 0 13632 0 -1 12852
box -48 -56 144 834
use sg13g2_fill_1  FILLER_15_148
timestamp 1677579658
transform 1 0 15360 0 -1 12852
box -48 -56 144 834
use sg13g2_decap_4  FILLER_15_196
timestamp 1679577901
transform 1 0 19968 0 -1 12852
box -48 -56 432 834
use sg13g2_decap_8  FILLER_16_0
timestamp 1679581782
transform 1 0 1152 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_7
timestamp 1679581782
transform 1 0 1824 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_35
timestamp 1679581782
transform 1 0 4512 0 1 12852
box -48 -56 720 834
use sg13g2_decap_4  FILLER_16_42
timestamp 1679577901
transform 1 0 5184 0 1 12852
box -48 -56 432 834
use sg13g2_fill_1  FILLER_16_139
timestamp 1677579658
transform 1 0 14496 0 1 12852
box -48 -56 144 834
use sg13g2_fill_2  FILLER_16_171
timestamp 1677580104
transform 1 0 17568 0 1 12852
box -48 -56 240 834
use sg13g2_decap_4  FILLER_16_195
timestamp 1679577901
transform 1 0 19872 0 1 12852
box -48 -56 432 834
use sg13g2_fill_1  FILLER_16_199
timestamp 1677579658
transform 1 0 20256 0 1 12852
box -48 -56 144 834
use sg13g2_decap_8  FILLER_17_0
timestamp 1679581782
transform 1 0 1152 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_7
timestamp 1679581782
transform 1 0 1824 0 -1 14364
box -48 -56 720 834
use sg13g2_fill_1  FILLER_17_14
timestamp 1677579658
transform 1 0 2496 0 -1 14364
box -48 -56 144 834
use sg13g2_decap_8  FILLER_17_36
timestamp 1679581782
transform 1 0 4608 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_4  FILLER_17_43
timestamp 1679577901
transform 1 0 5280 0 -1 14364
box -48 -56 432 834
use sg13g2_fill_1  FILLER_17_47
timestamp 1677579658
transform 1 0 5664 0 -1 14364
box -48 -56 144 834
use sg13g2_decap_4  FILLER_17_69
timestamp 1679577901
transform 1 0 7776 0 -1 14364
box -48 -56 432 834
use sg13g2_fill_2  FILLER_17_73
timestamp 1677580104
transform 1 0 8160 0 -1 14364
box -48 -56 240 834
use sg13g2_decap_8  FILLER_17_90
timestamp 1679581782
transform 1 0 9792 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_4  FILLER_17_97
timestamp 1679577901
transform 1 0 10464 0 -1 14364
box -48 -56 432 834
use sg13g2_fill_1  FILLER_17_101
timestamp 1677579658
transform 1 0 10848 0 -1 14364
box -48 -56 144 834
use sg13g2_fill_2  FILLER_17_119
timestamp 1677580104
transform 1 0 12576 0 -1 14364
box -48 -56 240 834
use sg13g2_decap_8  FILLER_17_170
timestamp 1679581782
transform 1 0 17472 0 -1 14364
box -48 -56 720 834
use sg13g2_fill_1  FILLER_17_199
timestamp 1677579658
transform 1 0 20256 0 -1 14364
box -48 -56 144 834
use sg13g2_fill_1  FILLER_18_32
timestamp 1677579658
transform 1 0 4224 0 1 14364
box -48 -56 144 834
use sg13g2_fill_2  FILLER_18_50
timestamp 1677580104
transform 1 0 5952 0 1 14364
box -48 -56 240 834
use sg13g2_fill_1  FILLER_18_69
timestamp 1677579658
transform 1 0 7776 0 1 14364
box -48 -56 144 834
use sg13g2_decap_8  FILLER_18_91
timestamp 1679581782
transform 1 0 9888 0 1 14364
box -48 -56 720 834
use sg13g2_fill_1  FILLER_18_98
timestamp 1677579658
transform 1 0 10560 0 1 14364
box -48 -56 144 834
use sg13g2_fill_2  FILLER_18_116
timestamp 1677580104
transform 1 0 12288 0 1 14364
box -48 -56 240 834
use sg13g2_fill_1  FILLER_18_118
timestamp 1677579658
transform 1 0 12480 0 1 14364
box -48 -56 144 834
use sg13g2_fill_1  FILLER_18_146
timestamp 1677579658
transform 1 0 15168 0 1 14364
box -48 -56 144 834
use sg13g2_decap_8  FILLER_18_164
timestamp 1679581782
transform 1 0 16896 0 1 14364
box -48 -56 720 834
use sg13g2_fill_1  FILLER_19_17
timestamp 1677579658
transform 1 0 2784 0 -1 15876
box -48 -56 144 834
use sg13g2_decap_8  FILLER_19_90
timestamp 1679581782
transform 1 0 9792 0 -1 15876
box -48 -56 720 834
use sg13g2_fill_2  FILLER_19_97
timestamp 1677580104
transform 1 0 10464 0 -1 15876
box -48 -56 240 834
use sg13g2_fill_1  FILLER_19_137
timestamp 1677579658
transform 1 0 14304 0 -1 15876
box -48 -56 144 834
use sg13g2_fill_2  FILLER_19_176
timestamp 1677580104
transform 1 0 18048 0 -1 15876
box -48 -56 240 834
use sg13g2_fill_1  FILLER_19_178
timestamp 1677579658
transform 1 0 18240 0 -1 15876
box -48 -56 144 834
use sg13g2_fill_2  FILLER_20_0
timestamp 1677580104
transform 1 0 1152 0 1 15876
box -48 -56 240 834
use sg13g2_fill_2  FILLER_20_19
timestamp 1677580104
transform 1 0 2976 0 1 15876
box -48 -56 240 834
use sg13g2_fill_2  FILLER_20_67
timestamp 1677580104
transform 1 0 7584 0 1 15876
box -48 -56 240 834
use sg13g2_decap_8  FILLER_20_103
timestamp 1679581782
transform 1 0 11040 0 1 15876
box -48 -56 720 834
use sg13g2_fill_1  FILLER_20_110
timestamp 1677579658
transform 1 0 11712 0 1 15876
box -48 -56 144 834
use sg13g2_decap_8  FILLER_20_128
timestamp 1679581782
transform 1 0 13440 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_135
timestamp 1679581782
transform 1 0 14112 0 1 15876
box -48 -56 720 834
use sg13g2_decap_4  FILLER_20_142
timestamp 1679577901
transform 1 0 14784 0 1 15876
box -48 -56 432 834
use sg13g2_fill_2  FILLER_20_146
timestamp 1677580104
transform 1 0 15168 0 1 15876
box -48 -56 240 834
use sg13g2_fill_2  FILLER_20_175
timestamp 1677580104
transform 1 0 17952 0 1 15876
box -48 -56 240 834
use sg13g2_fill_1  FILLER_20_199
timestamp 1677579658
transform 1 0 20256 0 1 15876
box -48 -56 144 834
use sg13g2_fill_2  FILLER_21_17
timestamp 1677580104
transform 1 0 2784 0 -1 17388
box -48 -56 240 834
use sg13g2_fill_1  FILLER_21_41
timestamp 1677579658
transform 1 0 5088 0 -1 17388
box -48 -56 144 834
use sg13g2_fill_1  FILLER_21_64
timestamp 1677579658
transform 1 0 7296 0 -1 17388
box -48 -56 144 834
use sg13g2_decap_8  FILLER_21_82
timestamp 1679581782
transform 1 0 9024 0 -1 17388
box -48 -56 720 834
use sg13g2_fill_2  FILLER_21_89
timestamp 1677580104
transform 1 0 9696 0 -1 17388
box -48 -56 240 834
use sg13g2_fill_1  FILLER_21_129
timestamp 1677579658
transform 1 0 13536 0 -1 17388
box -48 -56 144 834
use sg13g2_fill_1  FILLER_21_152
timestamp 1677579658
transform 1 0 15744 0 -1 17388
box -48 -56 144 834
use sg13g2_decap_8  FILLER_22_0
timestamp 1679581782
transform 1 0 1152 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_7
timestamp 1679581782
transform 1 0 1824 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_31
timestamp 1679581782
transform 1 0 4128 0 1 17388
box -48 -56 720 834
use sg13g2_decap_4  FILLER_22_38
timestamp 1679577901
transform 1 0 4800 0 1 17388
box -48 -56 432 834
use sg13g2_fill_2  FILLER_22_59
timestamp 1677580104
transform 1 0 6816 0 1 17388
box -48 -56 240 834
use sg13g2_decap_8  FILLER_22_103
timestamp 1679581782
transform 1 0 11040 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_110
timestamp 1679581782
transform 1 0 11712 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_117
timestamp 1679581782
transform 1 0 12384 0 1 17388
box -48 -56 720 834
use sg13g2_decap_4  FILLER_22_124
timestamp 1679577901
transform 1 0 13056 0 1 17388
box -48 -56 432 834
use sg13g2_fill_2  FILLER_22_128
timestamp 1677580104
transform 1 0 13440 0 1 17388
box -48 -56 240 834
use sg13g2_decap_8  FILLER_22_159
timestamp 1679581782
transform 1 0 16416 0 1 17388
box -48 -56 720 834
use sg13g2_fill_1  FILLER_22_166
timestamp 1677579658
transform 1 0 17088 0 1 17388
box -48 -56 144 834
use sg13g2_fill_2  FILLER_22_184
timestamp 1677580104
transform 1 0 18816 0 1 17388
box -48 -56 240 834
use sg13g2_decap_4  FILLER_22_196
timestamp 1679577901
transform 1 0 19968 0 1 17388
box -48 -56 432 834
use sg13g2_decap_8  FILLER_23_0
timestamp 1679581782
transform 1 0 1152 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_4  FILLER_23_7
timestamp 1679577901
transform 1 0 1824 0 -1 18900
box -48 -56 432 834
use sg13g2_fill_1  FILLER_23_11
timestamp 1677579658
transform 1 0 2208 0 -1 18900
box -48 -56 144 834
use sg13g2_decap_8  FILLER_23_33
timestamp 1679581782
transform 1 0 4320 0 -1 18900
box -48 -56 720 834
use sg13g2_fill_2  FILLER_23_40
timestamp 1677580104
transform 1 0 4992 0 -1 18900
box -48 -56 240 834
use sg13g2_fill_1  FILLER_23_42
timestamp 1677579658
transform 1 0 5184 0 -1 18900
box -48 -56 144 834
use sg13g2_decap_4  FILLER_23_67
timestamp 1679577901
transform 1 0 7584 0 -1 18900
box -48 -56 432 834
use sg13g2_fill_2  FILLER_23_71
timestamp 1677580104
transform 1 0 7968 0 -1 18900
box -48 -56 240 834
use sg13g2_fill_1  FILLER_23_153
timestamp 1677579658
transform 1 0 15840 0 -1 18900
box -48 -56 144 834
use sg13g2_decap_8  FILLER_24_17
timestamp 1679581782
transform 1 0 2784 0 1 18900
box -48 -56 720 834
use sg13g2_fill_1  FILLER_24_24
timestamp 1677579658
transform 1 0 3456 0 1 18900
box -48 -56 144 834
use sg13g2_decap_8  FILLER_24_47
timestamp 1679581782
transform 1 0 5664 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_54
timestamp 1679581782
transform 1 0 6336 0 1 18900
box -48 -56 720 834
use sg13g2_fill_2  FILLER_24_61
timestamp 1677580104
transform 1 0 7008 0 1 18900
box -48 -56 240 834
use sg13g2_decap_8  FILLER_24_97
timestamp 1679581782
transform 1 0 10464 0 1 18900
box -48 -56 720 834
use sg13g2_decap_4  FILLER_24_104
timestamp 1679577901
transform 1 0 11136 0 1 18900
box -48 -56 432 834
use sg13g2_fill_1  FILLER_24_130
timestamp 1677579658
transform 1 0 13632 0 1 18900
box -48 -56 144 834
use sg13g2_fill_1  FILLER_24_184
timestamp 1677579658
transform 1 0 18816 0 1 18900
box -48 -56 144 834
use sg13g2_fill_2  FILLER_24_197
timestamp 1677580104
transform 1 0 20064 0 1 18900
box -48 -56 240 834
use sg13g2_fill_1  FILLER_24_199
timestamp 1677579658
transform 1 0 20256 0 1 18900
box -48 -56 144 834
use sg13g2_fill_2  FILLER_25_0
timestamp 1677580104
transform 1 0 1152 0 -1 20412
box -48 -56 240 834
use sg13g2_fill_1  FILLER_25_2
timestamp 1677579658
transform 1 0 1344 0 -1 20412
box -48 -56 144 834
use sg13g2_fill_1  FILLER_25_20
timestamp 1677579658
transform 1 0 3072 0 -1 20412
box -48 -56 144 834
use sg13g2_decap_4  FILLER_25_38
timestamp 1679577901
transform 1 0 4800 0 -1 20412
box -48 -56 432 834
use sg13g2_fill_1  FILLER_25_42
timestamp 1677579658
transform 1 0 5184 0 -1 20412
box -48 -56 144 834
use sg13g2_fill_1  FILLER_25_98
timestamp 1677579658
transform 1 0 10560 0 -1 20412
box -48 -56 144 834
use sg13g2_decap_4  FILLER_25_124
timestamp 1679577901
transform 1 0 13056 0 -1 20412
box -48 -56 432 834
use sg13g2_fill_2  FILLER_25_150
timestamp 1677580104
transform 1 0 15552 0 -1 20412
box -48 -56 240 834
use sg13g2_decap_8  FILLER_25_169
timestamp 1679581782
transform 1 0 17376 0 -1 20412
box -48 -56 720 834
use sg13g2_fill_1  FILLER_25_176
timestamp 1677579658
transform 1 0 18048 0 -1 20412
box -48 -56 144 834
use sg13g2_fill_2  FILLER_25_198
timestamp 1677580104
transform 1 0 20160 0 -1 20412
box -48 -56 240 834
use sg13g2_decap_4  FILLER_26_0
timestamp 1679577901
transform 1 0 1152 0 1 20412
box -48 -56 432 834
use sg13g2_fill_2  FILLER_26_21
timestamp 1677580104
transform 1 0 3168 0 1 20412
box -48 -56 240 834
use sg13g2_decap_4  FILLER_26_44
timestamp 1679577901
transform 1 0 5376 0 1 20412
box -48 -56 432 834
use sg13g2_fill_2  FILLER_26_48
timestamp 1677580104
transform 1 0 5760 0 1 20412
box -48 -56 240 834
use sg13g2_decap_8  FILLER_26_88
timestamp 1679581782
transform 1 0 9600 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_95
timestamp 1679581782
transform 1 0 10272 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_162
timestamp 1679581782
transform 1 0 16704 0 1 20412
box -48 -56 720 834
use sg13g2_fill_2  FILLER_26_198
timestamp 1677580104
transform 1 0 20160 0 1 20412
box -48 -56 240 834
use sg13g2_decap_8  FILLER_27_0
timestamp 1679581782
transform 1 0 1152 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_7
timestamp 1679581782
transform 1 0 1824 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_4  FILLER_27_14
timestamp 1679577901
transform 1 0 2496 0 -1 21924
box -48 -56 432 834
use sg13g2_fill_1  FILLER_27_28
timestamp 1677579658
transform 1 0 3840 0 -1 21924
box -48 -56 144 834
use sg13g2_fill_1  FILLER_27_63
timestamp 1677579658
transform 1 0 7200 0 -1 21924
box -48 -56 144 834
use sg13g2_decap_4  FILLER_27_85
timestamp 1679577901
transform 1 0 9312 0 -1 21924
box -48 -56 432 834
use sg13g2_fill_1  FILLER_27_89
timestamp 1677579658
transform 1 0 9696 0 -1 21924
box -48 -56 144 834
use sg13g2_decap_8  FILLER_27_107
timestamp 1679581782
transform 1 0 11424 0 -1 21924
box -48 -56 720 834
use sg13g2_fill_2  FILLER_27_114
timestamp 1677580104
transform 1 0 12096 0 -1 21924
box -48 -56 240 834
use sg13g2_fill_1  FILLER_27_116
timestamp 1677579658
transform 1 0 12288 0 -1 21924
box -48 -56 144 834
use sg13g2_fill_1  FILLER_27_141
timestamp 1677579658
transform 1 0 14688 0 -1 21924
box -48 -56 144 834
use sg13g2_decap_4  FILLER_27_159
timestamp 1679577901
transform 1 0 16416 0 -1 21924
box -48 -56 432 834
use sg13g2_fill_1  FILLER_27_184
timestamp 1677579658
transform 1 0 18816 0 -1 21924
box -48 -56 144 834
use sg13g2_decap_8  FILLER_27_193
timestamp 1679581782
transform 1 0 19680 0 -1 21924
box -48 -56 720 834
use sg13g2_fill_2  FILLER_28_0
timestamp 1677580104
transform 1 0 1152 0 1 21924
box -48 -56 240 834
use sg13g2_decap_8  FILLER_28_46
timestamp 1679581782
transform 1 0 5568 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_53
timestamp 1679581782
transform 1 0 6240 0 1 21924
box -48 -56 720 834
use sg13g2_fill_1  FILLER_28_72
timestamp 1677579658
transform 1 0 8064 0 1 21924
box -48 -56 144 834
use sg13g2_fill_1  FILLER_28_145
timestamp 1677579658
transform 1 0 15072 0 1 21924
box -48 -56 144 834
use sg13g2_fill_2  FILLER_28_163
timestamp 1677580104
transform 1 0 16800 0 1 21924
box -48 -56 240 834
use sg13g2_fill_1  FILLER_28_165
timestamp 1677579658
transform 1 0 16992 0 1 21924
box -48 -56 144 834
use sg13g2_fill_2  FILLER_28_183
timestamp 1677580104
transform 1 0 18720 0 1 21924
box -48 -56 240 834
use sg13g2_fill_2  FILLER_28_197
timestamp 1677580104
transform 1 0 20064 0 1 21924
box -48 -56 240 834
use sg13g2_fill_1  FILLER_28_199
timestamp 1677579658
transform 1 0 20256 0 1 21924
box -48 -56 144 834
use sg13g2_fill_2  FILLER_29_0
timestamp 1677580104
transform 1 0 1152 0 -1 23436
box -48 -56 240 834
use sg13g2_fill_1  FILLER_29_19
timestamp 1677579658
transform 1 0 2976 0 -1 23436
box -48 -56 144 834
use sg13g2_decap_8  FILLER_29_91
timestamp 1679581782
transform 1 0 9888 0 -1 23436
box -48 -56 720 834
use sg13g2_fill_1  FILLER_29_98
timestamp 1677579658
transform 1 0 10560 0 -1 23436
box -48 -56 144 834
use sg13g2_decap_8  FILLER_29_133
timestamp 1679581782
transform 1 0 13920 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_140
timestamp 1679581782
transform 1 0 14592 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_147
timestamp 1679581782
transform 1 0 15264 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_154
timestamp 1679581782
transform 1 0 15936 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_161
timestamp 1679581782
transform 1 0 16608 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_168
timestamp 1679581782
transform 1 0 17280 0 -1 23436
box -48 -56 720 834
use sg13g2_fill_2  FILLER_29_175
timestamp 1677580104
transform 1 0 17952 0 -1 23436
box -48 -56 240 834
use sg13g2_fill_1  FILLER_29_177
timestamp 1677579658
transform 1 0 18144 0 -1 23436
box -48 -56 144 834
use sg13g2_fill_1  FILLER_29_199
timestamp 1677579658
transform 1 0 20256 0 -1 23436
box -48 -56 144 834
use sg13g2_fill_2  FILLER_30_31
timestamp 1677580104
transform 1 0 4128 0 1 23436
box -48 -56 240 834
use sg13g2_fill_1  FILLER_30_45
timestamp 1677579658
transform 1 0 5472 0 1 23436
box -48 -56 144 834
use sg13g2_fill_1  FILLER_30_80
timestamp 1677579658
transform 1 0 8832 0 1 23436
box -48 -56 144 834
use sg13g2_decap_8  FILLER_30_119
timestamp 1679581782
transform 1 0 12576 0 1 23436
box -48 -56 720 834
use sg13g2_decap_4  FILLER_30_126
timestamp 1679577901
transform 1 0 13248 0 1 23436
box -48 -56 432 834
use sg13g2_decap_8  FILLER_30_193
timestamp 1679581782
transform 1 0 19680 0 1 23436
box -48 -56 720 834
use sg13g2_fill_2  FILLER_31_22
timestamp 1677580104
transform 1 0 3264 0 -1 24948
box -48 -56 240 834
use sg13g2_fill_1  FILLER_31_24
timestamp 1677579658
transform 1 0 3456 0 -1 24948
box -48 -56 144 834
use sg13g2_fill_2  FILLER_31_59
timestamp 1677580104
transform 1 0 6816 0 -1 24948
box -48 -56 240 834
use sg13g2_fill_2  FILLER_31_71
timestamp 1677580104
transform 1 0 7968 0 -1 24948
box -48 -56 240 834
use sg13g2_decap_8  FILLER_31_111
timestamp 1679581782
transform 1 0 11808 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_118
timestamp 1679581782
transform 1 0 12480 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_125
timestamp 1679581782
transform 1 0 13152 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_149
timestamp 1679581782
transform 1 0 15456 0 -1 24948
box -48 -56 720 834
use sg13g2_fill_2  FILLER_31_156
timestamp 1677580104
transform 1 0 16128 0 -1 24948
box -48 -56 240 834
use sg13g2_fill_2  FILLER_31_179
timestamp 1677580104
transform 1 0 18336 0 -1 24948
box -48 -56 240 834
use sg13g2_fill_2  FILLER_31_197
timestamp 1677580104
transform 1 0 20064 0 -1 24948
box -48 -56 240 834
use sg13g2_fill_1  FILLER_31_199
timestamp 1677579658
transform 1 0 20256 0 -1 24948
box -48 -56 144 834
use sg13g2_decap_4  FILLER_32_0
timestamp 1679577901
transform 1 0 1152 0 1 24948
box -48 -56 432 834
use sg13g2_fill_1  FILLER_32_4
timestamp 1677579658
transform 1 0 1536 0 1 24948
box -48 -56 144 834
use sg13g2_fill_2  FILLER_32_22
timestamp 1677580104
transform 1 0 3264 0 1 24948
box -48 -56 240 834
use sg13g2_fill_1  FILLER_32_24
timestamp 1677579658
transform 1 0 3456 0 1 24948
box -48 -56 144 834
use sg13g2_decap_8  FILLER_32_46
timestamp 1679581782
transform 1 0 5568 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_53
timestamp 1679581782
transform 1 0 6240 0 1 24948
box -48 -56 720 834
use sg13g2_fill_1  FILLER_32_81
timestamp 1677579658
transform 1 0 8928 0 1 24948
box -48 -56 144 834
use sg13g2_decap_8  FILLER_32_120
timestamp 1679581782
transform 1 0 12672 0 1 24948
box -48 -56 720 834
use sg13g2_fill_2  FILLER_32_127
timestamp 1677580104
transform 1 0 13344 0 1 24948
box -48 -56 240 834
use sg13g2_decap_8  FILLER_32_150
timestamp 1679581782
transform 1 0 15552 0 1 24948
box -48 -56 720 834
use sg13g2_fill_1  FILLER_32_157
timestamp 1677579658
transform 1 0 16224 0 1 24948
box -48 -56 144 834
use sg13g2_decap_4  FILLER_33_0
timestamp 1679577901
transform 1 0 1152 0 -1 26460
box -48 -56 432 834
use sg13g2_fill_2  FILLER_33_42
timestamp 1677580104
transform 1 0 5184 0 -1 26460
box -48 -56 240 834
use sg13g2_decap_4  FILLER_33_78
timestamp 1679577901
transform 1 0 8640 0 -1 26460
box -48 -56 432 834
use sg13g2_fill_1  FILLER_33_82
timestamp 1677579658
transform 1 0 9024 0 -1 26460
box -48 -56 144 834
use sg13g2_decap_8  FILLER_33_134
timestamp 1679581782
transform 1 0 14016 0 -1 26460
box -48 -56 720 834
use sg13g2_fill_1  FILLER_33_141
timestamp 1677579658
transform 1 0 14688 0 -1 26460
box -48 -56 144 834
use sg13g2_decap_8  FILLER_33_159
timestamp 1679581782
transform 1 0 16416 0 -1 26460
box -48 -56 720 834
use sg13g2_fill_2  FILLER_33_166
timestamp 1677580104
transform 1 0 17088 0 -1 26460
box -48 -56 240 834
use sg13g2_fill_2  FILLER_33_197
timestamp 1677580104
transform 1 0 20064 0 -1 26460
box -48 -56 240 834
use sg13g2_fill_1  FILLER_33_199
timestamp 1677579658
transform 1 0 20256 0 -1 26460
box -48 -56 144 834
use sg13g2_decap_8  FILLER_34_68
timestamp 1679581782
transform 1 0 7680 0 1 26460
box -48 -56 720 834
use sg13g2_decap_4  FILLER_34_75
timestamp 1679577901
transform 1 0 8352 0 1 26460
box -48 -56 432 834
use sg13g2_fill_1  FILLER_34_79
timestamp 1677579658
transform 1 0 8736 0 1 26460
box -48 -56 144 834
use sg13g2_fill_2  FILLER_34_97
timestamp 1677580104
transform 1 0 10464 0 1 26460
box -48 -56 240 834
use sg13g2_fill_1  FILLER_34_99
timestamp 1677579658
transform 1 0 10656 0 1 26460
box -48 -56 144 834
use sg13g2_decap_8  FILLER_34_117
timestamp 1679581782
transform 1 0 12384 0 1 26460
box -48 -56 720 834
use sg13g2_decap_4  FILLER_34_124
timestamp 1679577901
transform 1 0 13056 0 1 26460
box -48 -56 432 834
use sg13g2_fill_1  FILLER_34_128
timestamp 1677579658
transform 1 0 13440 0 1 26460
box -48 -56 144 834
use sg13g2_decap_8  FILLER_34_146
timestamp 1679581782
transform 1 0 15168 0 1 26460
box -48 -56 720 834
use sg13g2_decap_4  FILLER_34_153
timestamp 1679577901
transform 1 0 15840 0 1 26460
box -48 -56 432 834
use sg13g2_fill_2  FILLER_34_157
timestamp 1677580104
transform 1 0 16224 0 1 26460
box -48 -56 240 834
use sg13g2_fill_2  FILLER_34_197
timestamp 1677580104
transform 1 0 20064 0 1 26460
box -48 -56 240 834
use sg13g2_fill_1  FILLER_34_199
timestamp 1677579658
transform 1 0 20256 0 1 26460
box -48 -56 144 834
use sg13g2_decap_8  FILLER_35_0
timestamp 1679581782
transform 1 0 1152 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_4  FILLER_35_7
timestamp 1679577901
transform 1 0 1824 0 -1 27972
box -48 -56 432 834
use sg13g2_fill_1  FILLER_35_11
timestamp 1677579658
transform 1 0 2208 0 -1 27972
box -48 -56 144 834
use sg13g2_decap_8  FILLER_35_33
timestamp 1679581782
transform 1 0 4320 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_4  FILLER_35_40
timestamp 1679577901
transform 1 0 4992 0 -1 27972
box -48 -56 432 834
use sg13g2_decap_8  FILLER_35_86
timestamp 1679581782
transform 1 0 9408 0 -1 27972
box -48 -56 720 834
use sg13g2_fill_2  FILLER_35_93
timestamp 1677580104
transform 1 0 10080 0 -1 27972
box -48 -56 240 834
use sg13g2_decap_8  FILLER_35_116
timestamp 1679581782
transform 1 0 12288 0 -1 27972
box -48 -56 720 834
use sg13g2_fill_1  FILLER_35_199
timestamp 1677579658
transform 1 0 20256 0 -1 27972
box -48 -56 144 834
use sg13g2_decap_8  FILLER_36_0
timestamp 1679581782
transform 1 0 1152 0 1 27972
box -48 -56 720 834
use sg13g2_decap_4  FILLER_36_45
timestamp 1679577901
transform 1 0 5472 0 1 27972
box -48 -56 432 834
use sg13g2_fill_2  FILLER_36_66
timestamp 1677580104
transform 1 0 7488 0 1 27972
box -48 -56 240 834
use sg13g2_decap_8  FILLER_36_85
timestamp 1679581782
transform 1 0 9312 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_113
timestamp 1679581782
transform 1 0 12000 0 1 27972
box -48 -56 720 834
use sg13g2_decap_4  FILLER_36_120
timestamp 1679577901
transform 1 0 12672 0 1 27972
box -48 -56 432 834
use sg13g2_fill_1  FILLER_36_124
timestamp 1677579658
transform 1 0 13056 0 1 27972
box -48 -56 144 834
use sg13g2_fill_2  FILLER_36_163
timestamp 1677580104
transform 1 0 16800 0 1 27972
box -48 -56 240 834
use sg13g2_fill_2  FILLER_36_198
timestamp 1677580104
transform 1 0 20160 0 1 27972
box -48 -56 240 834
use sg13g2_fill_2  FILLER_37_0
timestamp 1677580104
transform 1 0 1152 0 -1 29484
box -48 -56 240 834
use sg13g2_fill_1  FILLER_37_2
timestamp 1677579658
transform 1 0 1344 0 -1 29484
box -48 -56 144 834
use sg13g2_decap_8  FILLER_37_20
timestamp 1679581782
transform 1 0 3072 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_44
timestamp 1679581782
transform 1 0 5376 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_51
timestamp 1679581782
transform 1 0 6048 0 -1 29484
box -48 -56 720 834
use sg13g2_fill_2  FILLER_37_58
timestamp 1677580104
transform 1 0 6720 0 -1 29484
box -48 -56 240 834
use sg13g2_fill_1  FILLER_37_77
timestamp 1677579658
transform 1 0 8544 0 -1 29484
box -48 -56 144 834
use sg13g2_fill_2  FILLER_37_197
timestamp 1677580104
transform 1 0 20064 0 -1 29484
box -48 -56 240 834
use sg13g2_fill_1  FILLER_37_199
timestamp 1677579658
transform 1 0 20256 0 -1 29484
box -48 -56 144 834
use sg13g2_decap_8  FILLER_38_30
timestamp 1679581782
transform 1 0 4032 0 1 29484
box -48 -56 720 834
use sg13g2_decap_4  FILLER_38_37
timestamp 1679577901
transform 1 0 4704 0 1 29484
box -48 -56 432 834
use sg13g2_fill_2  FILLER_38_92
timestamp 1677580104
transform 1 0 9984 0 1 29484
box -48 -56 240 834
use sg13g2_fill_1  FILLER_38_94
timestamp 1677579658
transform 1 0 10176 0 1 29484
box -48 -56 144 834
use sg13g2_decap_8  FILLER_38_116
timestamp 1679581782
transform 1 0 12288 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_123
timestamp 1679581782
transform 1 0 12960 0 1 29484
box -48 -56 720 834
use sg13g2_fill_1  FILLER_38_130
timestamp 1677579658
transform 1 0 13632 0 1 29484
box -48 -56 144 834
use sg13g2_fill_2  FILLER_38_152
timestamp 1677580104
transform 1 0 15744 0 1 29484
box -48 -56 240 834
use sg13g2_fill_1  FILLER_38_154
timestamp 1677579658
transform 1 0 15936 0 1 29484
box -48 -56 144 834
use sg13g2_fill_2  FILLER_38_163
timestamp 1677580104
transform 1 0 16800 0 1 29484
box -48 -56 240 834
use sg13g2_fill_2  FILLER_38_186
timestamp 1677580104
transform 1 0 19008 0 1 29484
box -48 -56 240 834
use sg13g2_fill_1  FILLER_38_188
timestamp 1677579658
transform 1 0 19200 0 1 29484
box -48 -56 144 834
use sg13g2_fill_2  FILLER_38_197
timestamp 1677580104
transform 1 0 20064 0 1 29484
box -48 -56 240 834
use sg13g2_fill_1  FILLER_38_199
timestamp 1677579658
transform 1 0 20256 0 1 29484
box -48 -56 144 834
use sg13g2_decap_8  FILLER_39_0
timestamp 1679581782
transform 1 0 1152 0 -1 30996
box -48 -56 720 834
use sg13g2_fill_2  FILLER_39_7
timestamp 1677580104
transform 1 0 1824 0 -1 30996
box -48 -56 240 834
use sg13g2_fill_1  FILLER_39_9
timestamp 1677579658
transform 1 0 2016 0 -1 30996
box -48 -56 144 834
use sg13g2_fill_2  FILLER_39_58
timestamp 1677580104
transform 1 0 6720 0 -1 30996
box -48 -56 240 834
use sg13g2_decap_8  FILLER_39_67
timestamp 1679581782
transform 1 0 7584 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_4  FILLER_39_74
timestamp 1679577901
transform 1 0 8256 0 -1 30996
box -48 -56 432 834
use sg13g2_fill_2  FILLER_39_78
timestamp 1677580104
transform 1 0 8640 0 -1 30996
box -48 -56 240 834
use sg13g2_fill_2  FILLER_39_97
timestamp 1677580104
transform 1 0 10464 0 -1 30996
box -48 -56 240 834
use sg13g2_fill_1  FILLER_39_99
timestamp 1677579658
transform 1 0 10656 0 -1 30996
box -48 -56 144 834
use sg13g2_fill_2  FILLER_39_168
timestamp 1677580104
transform 1 0 17280 0 -1 30996
box -48 -56 240 834
use sg13g2_fill_1  FILLER_39_170
timestamp 1677579658
transform 1 0 17472 0 -1 30996
box -48 -56 144 834
use sg13g2_fill_2  FILLER_40_17
timestamp 1677580104
transform 1 0 2784 0 1 30996
box -48 -56 240 834
use sg13g2_decap_8  FILLER_40_22
timestamp 1679581782
transform 1 0 3264 0 1 30996
box -48 -56 720 834
use sg13g2_fill_1  FILLER_40_29
timestamp 1677579658
transform 1 0 3936 0 1 30996
box -48 -56 144 834
use sg13g2_fill_2  FILLER_40_88
timestamp 1677580104
transform 1 0 9600 0 1 30996
box -48 -56 240 834
use sg13g2_fill_1  FILLER_40_90
timestamp 1677579658
transform 1 0 9792 0 1 30996
box -48 -56 144 834
use sg13g2_decap_4  FILLER_40_112
timestamp 1679577901
transform 1 0 11904 0 1 30996
box -48 -56 432 834
use sg13g2_fill_2  FILLER_40_116
timestamp 1677580104
transform 1 0 12288 0 1 30996
box -48 -56 240 834
use sg13g2_decap_8  FILLER_40_135
timestamp 1679581782
transform 1 0 14112 0 1 30996
box -48 -56 720 834
use sg13g2_fill_2  FILLER_40_176
timestamp 1677580104
transform 1 0 18048 0 1 30996
box -48 -56 240 834
use sg13g2_fill_1  FILLER_40_178
timestamp 1677579658
transform 1 0 18240 0 1 30996
box -48 -56 144 834
use sg13g2_decap_8  FILLER_41_0
timestamp 1679581782
transform 1 0 1152 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_7
timestamp 1679581782
transform 1 0 1824 0 -1 32508
box -48 -56 720 834
use sg13g2_fill_2  FILLER_41_14
timestamp 1677580104
transform 1 0 2496 0 -1 32508
box -48 -56 240 834
use sg13g2_fill_2  FILLER_41_64
timestamp 1677580104
transform 1 0 7296 0 -1 32508
box -48 -56 240 834
use sg13g2_fill_1  FILLER_41_76
timestamp 1677579658
transform 1 0 8448 0 -1 32508
box -48 -56 144 834
use sg13g2_decap_4  FILLER_41_94
timestamp 1679577901
transform 1 0 10176 0 -1 32508
box -48 -56 432 834
use sg13g2_fill_1  FILLER_41_98
timestamp 1677579658
transform 1 0 10560 0 -1 32508
box -48 -56 144 834
use sg13g2_fill_2  FILLER_41_137
timestamp 1677580104
transform 1 0 14304 0 -1 32508
box -48 -56 240 834
use sg13g2_fill_1  FILLER_41_139
timestamp 1677579658
transform 1 0 14496 0 -1 32508
box -48 -56 144 834
use sg13g2_fill_2  FILLER_41_186
timestamp 1677580104
transform 1 0 19008 0 -1 32508
box -48 -56 240 834
use sg13g2_fill_1  FILLER_41_188
timestamp 1677579658
transform 1 0 19200 0 -1 32508
box -48 -56 144 834
use sg13g2_fill_2  FILLER_41_197
timestamp 1677580104
transform 1 0 20064 0 -1 32508
box -48 -56 240 834
use sg13g2_fill_1  FILLER_41_199
timestamp 1677579658
transform 1 0 20256 0 -1 32508
box -48 -56 144 834
use sg13g2_fill_1  FILLER_42_0
timestamp 1677579658
transform 1 0 1152 0 1 32508
box -48 -56 144 834
use sg13g2_fill_2  FILLER_42_9
timestamp 1677580104
transform 1 0 2016 0 1 32508
box -48 -56 240 834
use sg13g2_fill_1  FILLER_42_28
timestamp 1677579658
transform 1 0 3840 0 1 32508
box -48 -56 144 834
use sg13g2_fill_2  FILLER_42_46
timestamp 1677580104
transform 1 0 5568 0 1 32508
box -48 -56 240 834
use sg13g2_decap_4  FILLER_42_88
timestamp 1679577901
transform 1 0 9600 0 1 32508
box -48 -56 432 834
use sg13g2_fill_1  FILLER_42_92
timestamp 1677579658
transform 1 0 9984 0 1 32508
box -48 -56 144 834
use sg13g2_fill_2  FILLER_42_123
timestamp 1677580104
transform 1 0 12960 0 1 32508
box -48 -56 240 834
use sg13g2_fill_1  FILLER_42_125
timestamp 1677579658
transform 1 0 13152 0 1 32508
box -48 -56 144 834
use sg13g2_decap_4  FILLER_42_143
timestamp 1679577901
transform 1 0 14880 0 1 32508
box -48 -56 432 834
use sg13g2_fill_1  FILLER_42_147
timestamp 1677579658
transform 1 0 15264 0 1 32508
box -48 -56 144 834
use sg13g2_fill_2  FILLER_42_186
timestamp 1677580104
transform 1 0 19008 0 1 32508
box -48 -56 240 834
use sg13g2_fill_1  FILLER_42_188
timestamp 1677579658
transform 1 0 19200 0 1 32508
box -48 -56 144 834
use sg13g2_fill_2  FILLER_42_197
timestamp 1677580104
transform 1 0 20064 0 1 32508
box -48 -56 240 834
use sg13g2_fill_1  FILLER_42_199
timestamp 1677579658
transform 1 0 20256 0 1 32508
box -48 -56 144 834
use sg13g2_fill_2  FILLER_43_0
timestamp 1677580104
transform 1 0 1152 0 -1 34020
box -48 -56 240 834
use sg13g2_fill_1  FILLER_43_30
timestamp 1677579658
transform 1 0 4032 0 -1 34020
box -48 -56 144 834
use sg13g2_fill_2  FILLER_43_71
timestamp 1677580104
transform 1 0 7968 0 -1 34020
box -48 -56 240 834
use sg13g2_decap_4  FILLER_43_111
timestamp 1679577901
transform 1 0 11808 0 -1 34020
box -48 -56 432 834
use sg13g2_fill_1  FILLER_43_115
timestamp 1677579658
transform 1 0 12192 0 -1 34020
box -48 -56 144 834
use sg13g2_decap_8  FILLER_43_137
timestamp 1679581782
transform 1 0 14304 0 -1 34020
box -48 -56 720 834
use sg13g2_fill_2  FILLER_43_144
timestamp 1677580104
transform 1 0 14976 0 -1 34020
box -48 -56 240 834
use sg13g2_fill_2  FILLER_43_174
timestamp 1677580104
transform 1 0 17856 0 -1 34020
box -48 -56 240 834
use sg13g2_fill_1  FILLER_43_176
timestamp 1677579658
transform 1 0 18048 0 -1 34020
box -48 -56 144 834
use sg13g2_fill_2  FILLER_43_197
timestamp 1677580104
transform 1 0 20064 0 -1 34020
box -48 -56 240 834
use sg13g2_fill_1  FILLER_43_199
timestamp 1677579658
transform 1 0 20256 0 -1 34020
box -48 -56 144 834
use sg13g2_fill_1  FILLER_44_17
timestamp 1677579658
transform 1 0 2784 0 1 34020
box -48 -56 144 834
use sg13g2_fill_1  FILLER_44_30
timestamp 1677579658
transform 1 0 4032 0 1 34020
box -48 -56 144 834
use sg13g2_fill_1  FILLER_44_48
timestamp 1677579658
transform 1 0 5760 0 1 34020
box -48 -56 144 834
use sg13g2_decap_8  FILLER_44_90
timestamp 1679581782
transform 1 0 9792 0 1 34020
box -48 -56 720 834
use sg13g2_decap_4  FILLER_44_97
timestamp 1679577901
transform 1 0 10464 0 1 34020
box -48 -56 432 834
use sg13g2_fill_1  FILLER_44_101
timestamp 1677579658
transform 1 0 10848 0 1 34020
box -48 -56 144 834
use sg13g2_decap_4  FILLER_44_119
timestamp 1679577901
transform 1 0 12576 0 1 34020
box -48 -56 432 834
use sg13g2_fill_2  FILLER_44_123
timestamp 1677580104
transform 1 0 12960 0 1 34020
box -48 -56 240 834
use sg13g2_fill_1  FILLER_44_180
timestamp 1677579658
transform 1 0 18432 0 1 34020
box -48 -56 144 834
use sg13g2_fill_2  FILLER_44_197
timestamp 1677580104
transform 1 0 20064 0 1 34020
box -48 -56 240 834
use sg13g2_fill_1  FILLER_44_199
timestamp 1677579658
transform 1 0 20256 0 1 34020
box -48 -56 144 834
use sg13g2_fill_2  FILLER_45_0
timestamp 1677580104
transform 1 0 1152 0 -1 35532
box -48 -56 240 834
use sg13g2_fill_2  FILLER_45_48
timestamp 1677580104
transform 1 0 5760 0 -1 35532
box -48 -56 240 834
use sg13g2_fill_1  FILLER_45_50
timestamp 1677579658
transform 1 0 5952 0 -1 35532
box -48 -56 144 834
use sg13g2_fill_2  FILLER_45_198
timestamp 1677580104
transform 1 0 20160 0 -1 35532
box -48 -56 240 834
use sg13g2_fill_1  FILLER_46_0
timestamp 1677579658
transform 1 0 1152 0 1 35532
box -48 -56 144 834
use sg13g2_decap_4  FILLER_46_5
timestamp 1679577901
transform 1 0 1632 0 1 35532
box -48 -56 432 834
use sg13g2_fill_1  FILLER_46_9
timestamp 1677579658
transform 1 0 2016 0 1 35532
box -48 -56 144 834
use sg13g2_decap_8  FILLER_46_13
timestamp 1679581782
transform 1 0 2400 0 1 35532
box -48 -56 720 834
use sg13g2_fill_2  FILLER_46_20
timestamp 1677580104
transform 1 0 3072 0 1 35532
box -48 -56 240 834
use sg13g2_fill_1  FILLER_46_22
timestamp 1677579658
transform 1 0 3264 0 1 35532
box -48 -56 144 834
use sg13g2_fill_2  FILLER_46_31
timestamp 1677580104
transform 1 0 4128 0 1 35532
box -48 -56 240 834
use sg13g2_fill_1  FILLER_46_33
timestamp 1677579658
transform 1 0 4320 0 1 35532
box -48 -56 144 834
use sg13g2_decap_8  FILLER_46_75
timestamp 1679581782
transform 1 0 8352 0 1 35532
box -48 -56 720 834
use sg13g2_fill_2  FILLER_46_82
timestamp 1677580104
transform 1 0 9024 0 1 35532
box -48 -56 240 834
use sg13g2_fill_1  FILLER_46_84
timestamp 1677579658
transform 1 0 9216 0 1 35532
box -48 -56 144 834
use sg13g2_fill_1  FILLER_46_199
timestamp 1677579658
transform 1 0 20256 0 1 35532
box -48 -56 144 834
use sg13g2_fill_1  FILLER_47_0
timestamp 1677579658
transform 1 0 1152 0 -1 37044
box -48 -56 144 834
use sg13g2_fill_1  FILLER_47_9
timestamp 1677579658
transform 1 0 2016 0 -1 37044
box -48 -56 144 834
use sg13g2_decap_8  FILLER_47_14
timestamp 1679581782
transform 1 0 2496 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_4  FILLER_47_21
timestamp 1679577901
transform 1 0 3168 0 -1 37044
box -48 -56 432 834
use sg13g2_fill_2  FILLER_47_25
timestamp 1677580104
transform 1 0 3552 0 -1 37044
box -48 -56 240 834
use sg13g2_fill_1  FILLER_47_30
timestamp 1677579658
transform 1 0 4032 0 -1 37044
box -48 -56 144 834
use sg13g2_fill_1  FILLER_47_38
timestamp 1677579658
transform 1 0 4800 0 -1 37044
box -48 -56 144 834
use sg13g2_fill_2  FILLER_47_63
timestamp 1677580104
transform 1 0 7200 0 -1 37044
box -48 -56 240 834
use sg13g2_fill_1  FILLER_47_137
timestamp 1677579658
transform 1 0 14304 0 -1 37044
box -48 -56 144 834
use sg13g2_fill_1  FILLER_47_184
timestamp 1677579658
transform 1 0 18816 0 -1 37044
box -48 -56 144 834
use sg13g2_fill_2  FILLER_47_197
timestamp 1677580104
transform 1 0 20064 0 -1 37044
box -48 -56 240 834
use sg13g2_fill_1  FILLER_47_199
timestamp 1677579658
transform 1 0 20256 0 -1 37044
box -48 -56 144 834
use sg13g2_fill_1  FILLER_48_11
timestamp 1677579658
transform 1 0 2208 0 1 37044
box -48 -56 144 834
use sg13g2_fill_1  FILLER_48_33
timestamp 1677579658
transform 1 0 4320 0 1 37044
box -48 -56 144 834
use sg13g2_fill_2  FILLER_48_104
timestamp 1677580104
transform 1 0 11136 0 1 37044
box -48 -56 240 834
use sg13g2_fill_1  FILLER_48_106
timestamp 1677579658
transform 1 0 11328 0 1 37044
box -48 -56 144 834
use sg13g2_fill_2  FILLER_48_124
timestamp 1677580104
transform 1 0 13056 0 1 37044
box -48 -56 240 834
use sg13g2_fill_2  FILLER_48_143
timestamp 1677580104
transform 1 0 14880 0 1 37044
box -48 -56 240 834
use sg13g2_fill_1  FILLER_48_145
timestamp 1677579658
transform 1 0 15072 0 1 37044
box -48 -56 144 834
use sg13g2_fill_2  FILLER_49_33
timestamp 1677580104
transform 1 0 4320 0 -1 38556
box -48 -56 240 834
use sg13g2_fill_1  FILLER_49_35
timestamp 1677579658
transform 1 0 4512 0 -1 38556
box -48 -56 144 834
use sg13g2_fill_2  FILLER_49_57
timestamp 1677580104
transform 1 0 6624 0 -1 38556
box -48 -56 240 834
use sg13g2_fill_2  FILLER_49_67
timestamp 1677580104
transform 1 0 7584 0 -1 38556
box -48 -56 240 834
use sg13g2_fill_1  FILLER_49_86
timestamp 1677579658
transform 1 0 9408 0 -1 38556
box -48 -56 144 834
use sg13g2_fill_2  FILLER_49_111
timestamp 1677580104
transform 1 0 11808 0 -1 38556
box -48 -56 240 834
use sg13g2_fill_1  FILLER_49_184
timestamp 1677579658
transform 1 0 18816 0 -1 38556
box -48 -56 144 834
use sg13g2_fill_1  FILLER_50_0
timestamp 1677579658
transform 1 0 1152 0 1 38556
box -48 -56 144 834
use sg13g2_decap_4  FILLER_50_25
timestamp 1679577901
transform 1 0 3552 0 1 38556
box -48 -56 432 834
use sg13g2_fill_2  FILLER_50_29
timestamp 1677580104
transform 1 0 3936 0 1 38556
box -48 -56 240 834
use sg13g2_decap_8  FILLER_50_35
timestamp 1679581782
transform 1 0 4512 0 1 38556
box -48 -56 720 834
use sg13g2_decap_4  FILLER_50_42
timestamp 1679577901
transform 1 0 5184 0 1 38556
box -48 -56 432 834
use sg13g2_fill_1  FILLER_50_46
timestamp 1677579658
transform 1 0 5568 0 1 38556
box -48 -56 144 834
use sg13g2_decap_4  FILLER_50_89
timestamp 1679577901
transform 1 0 9696 0 1 38556
box -48 -56 432 834
use sg13g2_fill_1  FILLER_50_93
timestamp 1677579658
transform 1 0 10080 0 1 38556
box -48 -56 144 834
use sg13g2_fill_2  FILLER_50_111
timestamp 1677580104
transform 1 0 11808 0 1 38556
box -48 -56 240 834
use sg13g2_fill_1  FILLER_50_117
timestamp 1677579658
transform 1 0 12384 0 1 38556
box -48 -56 144 834
use sg13g2_fill_2  FILLER_50_135
timestamp 1677580104
transform 1 0 14112 0 1 38556
box -48 -56 240 834
use sg13g2_fill_1  FILLER_50_137
timestamp 1677579658
transform 1 0 14304 0 1 38556
box -48 -56 144 834
use sg13g2_fill_2  FILLER_50_175
timestamp 1677580104
transform 1 0 17952 0 1 38556
box -48 -56 240 834
use sg13g2_fill_1  FILLER_50_184
timestamp 1677579658
transform 1 0 18816 0 1 38556
box -48 -56 144 834
use sg13g2_fill_1  FILLER_51_4
timestamp 1677579658
transform 1 0 1536 0 -1 40068
box -48 -56 144 834
use sg13g2_decap_4  FILLER_51_29
timestamp 1679577901
transform 1 0 3936 0 -1 40068
box -48 -56 432 834
use sg13g2_decap_8  FILLER_51_53
timestamp 1679581782
transform 1 0 6240 0 -1 40068
box -48 -56 720 834
use sg13g2_fill_2  FILLER_51_143
timestamp 1677580104
transform 1 0 14880 0 -1 40068
box -48 -56 240 834
use sg13g2_fill_1  FILLER_51_145
timestamp 1677579658
transform 1 0 15072 0 -1 40068
box -48 -56 144 834
use sg13g2_fill_2  FILLER_52_7
timestamp 1677580104
transform 1 0 1824 0 1 40068
box -48 -56 240 834
use sg13g2_fill_2  FILLER_52_47
timestamp 1677580104
transform 1 0 5664 0 1 40068
box -48 -56 240 834
use sg13g2_fill_1  FILLER_52_49
timestamp 1677579658
transform 1 0 5856 0 1 40068
box -48 -56 144 834
use sg13g2_fill_1  FILLER_52_71
timestamp 1677579658
transform 1 0 7968 0 1 40068
box -48 -56 144 834
use sg13g2_fill_1  FILLER_52_166
timestamp 1677579658
transform 1 0 17088 0 1 40068
box -48 -56 144 834
use sg13g2_fill_2  FILLER_52_198
timestamp 1677580104
transform 1 0 20160 0 1 40068
box -48 -56 240 834
use sg13g2_fill_2  FILLER_53_3
timestamp 1677580104
transform 1 0 1440 0 -1 41580
box -48 -56 240 834
use sg13g2_fill_1  FILLER_53_5
timestamp 1677579658
transform 1 0 1632 0 -1 41580
box -48 -56 144 834
use sg13g2_decap_8  FILLER_53_40
timestamp 1679581782
transform 1 0 4992 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_4  FILLER_53_47
timestamp 1679577901
transform 1 0 5664 0 -1 41580
box -48 -56 432 834
use sg13g2_fill_2  FILLER_53_68
timestamp 1677580104
transform 1 0 7680 0 -1 41580
box -48 -56 240 834
use sg13g2_fill_1  FILLER_53_70
timestamp 1677579658
transform 1 0 7872 0 -1 41580
box -48 -56 144 834
use sg13g2_fill_2  FILLER_53_75
timestamp 1677580104
transform 1 0 8352 0 -1 41580
box -48 -56 240 834
use sg13g2_fill_1  FILLER_53_77
timestamp 1677579658
transform 1 0 8544 0 -1 41580
box -48 -56 144 834
use sg13g2_fill_2  FILLER_53_158
timestamp 1677580104
transform 1 0 16320 0 -1 41580
box -48 -56 240 834
use sg13g2_fill_1  FILLER_53_160
timestamp 1677579658
transform 1 0 16512 0 -1 41580
box -48 -56 144 834
use sg13g2_fill_2  FILLER_53_197
timestamp 1677580104
transform 1 0 20064 0 -1 41580
box -48 -56 240 834
use sg13g2_fill_1  FILLER_53_199
timestamp 1677579658
transform 1 0 20256 0 -1 41580
box -48 -56 144 834
<< labels >>
flabel metal3 s 0 23396 80 23476 0 FreeSans 320 0 0 0 CLK_TT_PROJECT
port 0 nsew signal output
flabel metal3 s 21424 16172 21504 16252 0 FreeSans 320 0 0 0 E1BEG[0]
port 1 nsew signal output
flabel metal3 s 21424 16508 21504 16588 0 FreeSans 320 0 0 0 E1BEG[1]
port 2 nsew signal output
flabel metal3 s 21424 16844 21504 16924 0 FreeSans 320 0 0 0 E1BEG[2]
port 3 nsew signal output
flabel metal3 s 21424 17180 21504 17260 0 FreeSans 320 0 0 0 E1BEG[3]
port 4 nsew signal output
flabel metal3 s 21424 17516 21504 17596 0 FreeSans 320 0 0 0 E2BEG[0]
port 5 nsew signal output
flabel metal3 s 21424 17852 21504 17932 0 FreeSans 320 0 0 0 E2BEG[1]
port 6 nsew signal output
flabel metal3 s 21424 18188 21504 18268 0 FreeSans 320 0 0 0 E2BEG[2]
port 7 nsew signal output
flabel metal3 s 21424 18524 21504 18604 0 FreeSans 320 0 0 0 E2BEG[3]
port 8 nsew signal output
flabel metal3 s 21424 18860 21504 18940 0 FreeSans 320 0 0 0 E2BEG[4]
port 9 nsew signal output
flabel metal3 s 21424 19196 21504 19276 0 FreeSans 320 0 0 0 E2BEG[5]
port 10 nsew signal output
flabel metal3 s 21424 19532 21504 19612 0 FreeSans 320 0 0 0 E2BEG[6]
port 11 nsew signal output
flabel metal3 s 21424 19868 21504 19948 0 FreeSans 320 0 0 0 E2BEG[7]
port 12 nsew signal output
flabel metal3 s 21424 20204 21504 20284 0 FreeSans 320 0 0 0 E2BEGb[0]
port 13 nsew signal output
flabel metal3 s 21424 20540 21504 20620 0 FreeSans 320 0 0 0 E2BEGb[1]
port 14 nsew signal output
flabel metal3 s 21424 20876 21504 20956 0 FreeSans 320 0 0 0 E2BEGb[2]
port 15 nsew signal output
flabel metal3 s 21424 21212 21504 21292 0 FreeSans 320 0 0 0 E2BEGb[3]
port 16 nsew signal output
flabel metal3 s 21424 21548 21504 21628 0 FreeSans 320 0 0 0 E2BEGb[4]
port 17 nsew signal output
flabel metal3 s 21424 21884 21504 21964 0 FreeSans 320 0 0 0 E2BEGb[5]
port 18 nsew signal output
flabel metal3 s 21424 22220 21504 22300 0 FreeSans 320 0 0 0 E2BEGb[6]
port 19 nsew signal output
flabel metal3 s 21424 22556 21504 22636 0 FreeSans 320 0 0 0 E2BEGb[7]
port 20 nsew signal output
flabel metal3 s 21424 28268 21504 28348 0 FreeSans 320 0 0 0 E6BEG[0]
port 21 nsew signal output
flabel metal3 s 21424 31628 21504 31708 0 FreeSans 320 0 0 0 E6BEG[10]
port 22 nsew signal output
flabel metal3 s 21424 31964 21504 32044 0 FreeSans 320 0 0 0 E6BEG[11]
port 23 nsew signal output
flabel metal3 s 21424 28604 21504 28684 0 FreeSans 320 0 0 0 E6BEG[1]
port 24 nsew signal output
flabel metal3 s 21424 28940 21504 29020 0 FreeSans 320 0 0 0 E6BEG[2]
port 25 nsew signal output
flabel metal3 s 21424 29276 21504 29356 0 FreeSans 320 0 0 0 E6BEG[3]
port 26 nsew signal output
flabel metal3 s 21424 29612 21504 29692 0 FreeSans 320 0 0 0 E6BEG[4]
port 27 nsew signal output
flabel metal3 s 21424 29948 21504 30028 0 FreeSans 320 0 0 0 E6BEG[5]
port 28 nsew signal output
flabel metal3 s 21424 30284 21504 30364 0 FreeSans 320 0 0 0 E6BEG[6]
port 29 nsew signal output
flabel metal3 s 21424 30620 21504 30700 0 FreeSans 320 0 0 0 E6BEG[7]
port 30 nsew signal output
flabel metal3 s 21424 30956 21504 31036 0 FreeSans 320 0 0 0 E6BEG[8]
port 31 nsew signal output
flabel metal3 s 21424 31292 21504 31372 0 FreeSans 320 0 0 0 E6BEG[9]
port 32 nsew signal output
flabel metal3 s 21424 22892 21504 22972 0 FreeSans 320 0 0 0 EE4BEG[0]
port 33 nsew signal output
flabel metal3 s 21424 26252 21504 26332 0 FreeSans 320 0 0 0 EE4BEG[10]
port 34 nsew signal output
flabel metal3 s 21424 26588 21504 26668 0 FreeSans 320 0 0 0 EE4BEG[11]
port 35 nsew signal output
flabel metal3 s 21424 26924 21504 27004 0 FreeSans 320 0 0 0 EE4BEG[12]
port 36 nsew signal output
flabel metal3 s 21424 27260 21504 27340 0 FreeSans 320 0 0 0 EE4BEG[13]
port 37 nsew signal output
flabel metal3 s 21424 27596 21504 27676 0 FreeSans 320 0 0 0 EE4BEG[14]
port 38 nsew signal output
flabel metal3 s 21424 27932 21504 28012 0 FreeSans 320 0 0 0 EE4BEG[15]
port 39 nsew signal output
flabel metal3 s 21424 23228 21504 23308 0 FreeSans 320 0 0 0 EE4BEG[1]
port 40 nsew signal output
flabel metal3 s 21424 23564 21504 23644 0 FreeSans 320 0 0 0 EE4BEG[2]
port 41 nsew signal output
flabel metal3 s 21424 23900 21504 23980 0 FreeSans 320 0 0 0 EE4BEG[3]
port 42 nsew signal output
flabel metal3 s 21424 24236 21504 24316 0 FreeSans 320 0 0 0 EE4BEG[4]
port 43 nsew signal output
flabel metal3 s 21424 24572 21504 24652 0 FreeSans 320 0 0 0 EE4BEG[5]
port 44 nsew signal output
flabel metal3 s 21424 24908 21504 24988 0 FreeSans 320 0 0 0 EE4BEG[6]
port 45 nsew signal output
flabel metal3 s 21424 25244 21504 25324 0 FreeSans 320 0 0 0 EE4BEG[7]
port 46 nsew signal output
flabel metal3 s 21424 25580 21504 25660 0 FreeSans 320 0 0 0 EE4BEG[8]
port 47 nsew signal output
flabel metal3 s 21424 25916 21504 25996 0 FreeSans 320 0 0 0 EE4BEG[9]
port 48 nsew signal output
flabel metal3 s 0 22892 80 22972 0 FreeSans 320 0 0 0 ENA_TT_PROJECT
port 49 nsew signal output
flabel metal3 s 0 24404 80 24484 0 FreeSans 320 0 0 0 FrameData[0]
port 50 nsew signal input
flabel metal3 s 0 29444 80 29524 0 FreeSans 320 0 0 0 FrameData[10]
port 51 nsew signal input
flabel metal3 s 0 29948 80 30028 0 FreeSans 320 0 0 0 FrameData[11]
port 52 nsew signal input
flabel metal3 s 0 30452 80 30532 0 FreeSans 320 0 0 0 FrameData[12]
port 53 nsew signal input
flabel metal3 s 0 30956 80 31036 0 FreeSans 320 0 0 0 FrameData[13]
port 54 nsew signal input
flabel metal3 s 0 31460 80 31540 0 FreeSans 320 0 0 0 FrameData[14]
port 55 nsew signal input
flabel metal3 s 0 31964 80 32044 0 FreeSans 320 0 0 0 FrameData[15]
port 56 nsew signal input
flabel metal3 s 0 32468 80 32548 0 FreeSans 320 0 0 0 FrameData[16]
port 57 nsew signal input
flabel metal3 s 0 32972 80 33052 0 FreeSans 320 0 0 0 FrameData[17]
port 58 nsew signal input
flabel metal3 s 0 33476 80 33556 0 FreeSans 320 0 0 0 FrameData[18]
port 59 nsew signal input
flabel metal3 s 0 33980 80 34060 0 FreeSans 320 0 0 0 FrameData[19]
port 60 nsew signal input
flabel metal3 s 0 24908 80 24988 0 FreeSans 320 0 0 0 FrameData[1]
port 61 nsew signal input
flabel metal3 s 0 34484 80 34564 0 FreeSans 320 0 0 0 FrameData[20]
port 62 nsew signal input
flabel metal3 s 0 34988 80 35068 0 FreeSans 320 0 0 0 FrameData[21]
port 63 nsew signal input
flabel metal3 s 0 35492 80 35572 0 FreeSans 320 0 0 0 FrameData[22]
port 64 nsew signal input
flabel metal3 s 0 35996 80 36076 0 FreeSans 320 0 0 0 FrameData[23]
port 65 nsew signal input
flabel metal3 s 0 36500 80 36580 0 FreeSans 320 0 0 0 FrameData[24]
port 66 nsew signal input
flabel metal3 s 0 37004 80 37084 0 FreeSans 320 0 0 0 FrameData[25]
port 67 nsew signal input
flabel metal3 s 0 37508 80 37588 0 FreeSans 320 0 0 0 FrameData[26]
port 68 nsew signal input
flabel metal3 s 0 38012 80 38092 0 FreeSans 320 0 0 0 FrameData[27]
port 69 nsew signal input
flabel metal3 s 0 38516 80 38596 0 FreeSans 320 0 0 0 FrameData[28]
port 70 nsew signal input
flabel metal3 s 0 39020 80 39100 0 FreeSans 320 0 0 0 FrameData[29]
port 71 nsew signal input
flabel metal3 s 0 25412 80 25492 0 FreeSans 320 0 0 0 FrameData[2]
port 72 nsew signal input
flabel metal3 s 0 39524 80 39604 0 FreeSans 320 0 0 0 FrameData[30]
port 73 nsew signal input
flabel metal3 s 0 40028 80 40108 0 FreeSans 320 0 0 0 FrameData[31]
port 74 nsew signal input
flabel metal3 s 0 25916 80 25996 0 FreeSans 320 0 0 0 FrameData[3]
port 75 nsew signal input
flabel metal3 s 0 26420 80 26500 0 FreeSans 320 0 0 0 FrameData[4]
port 76 nsew signal input
flabel metal3 s 0 26924 80 27004 0 FreeSans 320 0 0 0 FrameData[5]
port 77 nsew signal input
flabel metal3 s 0 27428 80 27508 0 FreeSans 320 0 0 0 FrameData[6]
port 78 nsew signal input
flabel metal3 s 0 27932 80 28012 0 FreeSans 320 0 0 0 FrameData[7]
port 79 nsew signal input
flabel metal3 s 0 28436 80 28516 0 FreeSans 320 0 0 0 FrameData[8]
port 80 nsew signal input
flabel metal3 s 0 28940 80 29020 0 FreeSans 320 0 0 0 FrameData[9]
port 81 nsew signal input
flabel metal3 s 21424 32300 21504 32380 0 FreeSans 320 0 0 0 FrameData_O[0]
port 82 nsew signal output
flabel metal3 s 21424 35660 21504 35740 0 FreeSans 320 0 0 0 FrameData_O[10]
port 83 nsew signal output
flabel metal3 s 21424 35996 21504 36076 0 FreeSans 320 0 0 0 FrameData_O[11]
port 84 nsew signal output
flabel metal3 s 21424 36332 21504 36412 0 FreeSans 320 0 0 0 FrameData_O[12]
port 85 nsew signal output
flabel metal3 s 21424 36668 21504 36748 0 FreeSans 320 0 0 0 FrameData_O[13]
port 86 nsew signal output
flabel metal3 s 21424 37004 21504 37084 0 FreeSans 320 0 0 0 FrameData_O[14]
port 87 nsew signal output
flabel metal3 s 21424 37340 21504 37420 0 FreeSans 320 0 0 0 FrameData_O[15]
port 88 nsew signal output
flabel metal3 s 21424 37676 21504 37756 0 FreeSans 320 0 0 0 FrameData_O[16]
port 89 nsew signal output
flabel metal3 s 21424 38012 21504 38092 0 FreeSans 320 0 0 0 FrameData_O[17]
port 90 nsew signal output
flabel metal3 s 21424 38348 21504 38428 0 FreeSans 320 0 0 0 FrameData_O[18]
port 91 nsew signal output
flabel metal3 s 21424 38684 21504 38764 0 FreeSans 320 0 0 0 FrameData_O[19]
port 92 nsew signal output
flabel metal3 s 21424 32636 21504 32716 0 FreeSans 320 0 0 0 FrameData_O[1]
port 93 nsew signal output
flabel metal3 s 21424 39020 21504 39100 0 FreeSans 320 0 0 0 FrameData_O[20]
port 94 nsew signal output
flabel metal3 s 21424 39356 21504 39436 0 FreeSans 320 0 0 0 FrameData_O[21]
port 95 nsew signal output
flabel metal3 s 21424 39692 21504 39772 0 FreeSans 320 0 0 0 FrameData_O[22]
port 96 nsew signal output
flabel metal3 s 21424 40028 21504 40108 0 FreeSans 320 0 0 0 FrameData_O[23]
port 97 nsew signal output
flabel metal3 s 21424 40364 21504 40444 0 FreeSans 320 0 0 0 FrameData_O[24]
port 98 nsew signal output
flabel metal3 s 21424 40700 21504 40780 0 FreeSans 320 0 0 0 FrameData_O[25]
port 99 nsew signal output
flabel metal3 s 21424 41036 21504 41116 0 FreeSans 320 0 0 0 FrameData_O[26]
port 100 nsew signal output
flabel metal3 s 21424 41372 21504 41452 0 FreeSans 320 0 0 0 FrameData_O[27]
port 101 nsew signal output
flabel metal3 s 21424 41708 21504 41788 0 FreeSans 320 0 0 0 FrameData_O[28]
port 102 nsew signal output
flabel metal3 s 21424 42044 21504 42124 0 FreeSans 320 0 0 0 FrameData_O[29]
port 103 nsew signal output
flabel metal3 s 21424 32972 21504 33052 0 FreeSans 320 0 0 0 FrameData_O[2]
port 104 nsew signal output
flabel metal3 s 21424 42380 21504 42460 0 FreeSans 320 0 0 0 FrameData_O[30]
port 105 nsew signal output
flabel metal3 s 21424 42716 21504 42796 0 FreeSans 320 0 0 0 FrameData_O[31]
port 106 nsew signal output
flabel metal3 s 21424 33308 21504 33388 0 FreeSans 320 0 0 0 FrameData_O[3]
port 107 nsew signal output
flabel metal3 s 21424 33644 21504 33724 0 FreeSans 320 0 0 0 FrameData_O[4]
port 108 nsew signal output
flabel metal3 s 21424 33980 21504 34060 0 FreeSans 320 0 0 0 FrameData_O[5]
port 109 nsew signal output
flabel metal3 s 21424 34316 21504 34396 0 FreeSans 320 0 0 0 FrameData_O[6]
port 110 nsew signal output
flabel metal3 s 21424 34652 21504 34732 0 FreeSans 320 0 0 0 FrameData_O[7]
port 111 nsew signal output
flabel metal3 s 21424 34988 21504 35068 0 FreeSans 320 0 0 0 FrameData_O[8]
port 112 nsew signal output
flabel metal3 s 21424 35324 21504 35404 0 FreeSans 320 0 0 0 FrameData_O[9]
port 113 nsew signal output
flabel metal2 s 15800 0 15880 80 0 FreeSans 320 0 0 0 FrameStrobe[0]
port 114 nsew signal input
flabel metal2 s 17720 0 17800 80 0 FreeSans 320 0 0 0 FrameStrobe[10]
port 115 nsew signal input
flabel metal2 s 17912 0 17992 80 0 FreeSans 320 0 0 0 FrameStrobe[11]
port 116 nsew signal input
flabel metal2 s 18104 0 18184 80 0 FreeSans 320 0 0 0 FrameStrobe[12]
port 117 nsew signal input
flabel metal2 s 18296 0 18376 80 0 FreeSans 320 0 0 0 FrameStrobe[13]
port 118 nsew signal input
flabel metal2 s 18488 0 18568 80 0 FreeSans 320 0 0 0 FrameStrobe[14]
port 119 nsew signal input
flabel metal2 s 18680 0 18760 80 0 FreeSans 320 0 0 0 FrameStrobe[15]
port 120 nsew signal input
flabel metal2 s 18872 0 18952 80 0 FreeSans 320 0 0 0 FrameStrobe[16]
port 121 nsew signal input
flabel metal2 s 19064 0 19144 80 0 FreeSans 320 0 0 0 FrameStrobe[17]
port 122 nsew signal input
flabel metal2 s 19256 0 19336 80 0 FreeSans 320 0 0 0 FrameStrobe[18]
port 123 nsew signal input
flabel metal2 s 19448 0 19528 80 0 FreeSans 320 0 0 0 FrameStrobe[19]
port 124 nsew signal input
flabel metal2 s 15992 0 16072 80 0 FreeSans 320 0 0 0 FrameStrobe[1]
port 125 nsew signal input
flabel metal2 s 16184 0 16264 80 0 FreeSans 320 0 0 0 FrameStrobe[2]
port 126 nsew signal input
flabel metal2 s 16376 0 16456 80 0 FreeSans 320 0 0 0 FrameStrobe[3]
port 127 nsew signal input
flabel metal2 s 16568 0 16648 80 0 FreeSans 320 0 0 0 FrameStrobe[4]
port 128 nsew signal input
flabel metal2 s 16760 0 16840 80 0 FreeSans 320 0 0 0 FrameStrobe[5]
port 129 nsew signal input
flabel metal2 s 16952 0 17032 80 0 FreeSans 320 0 0 0 FrameStrobe[6]
port 130 nsew signal input
flabel metal2 s 17144 0 17224 80 0 FreeSans 320 0 0 0 FrameStrobe[7]
port 131 nsew signal input
flabel metal2 s 17336 0 17416 80 0 FreeSans 320 0 0 0 FrameStrobe[8]
port 132 nsew signal input
flabel metal2 s 17528 0 17608 80 0 FreeSans 320 0 0 0 FrameStrobe[9]
port 133 nsew signal input
flabel metal2 s 15800 42928 15880 43008 0 FreeSans 320 0 0 0 FrameStrobe_O[0]
port 134 nsew signal output
flabel metal2 s 17720 42928 17800 43008 0 FreeSans 320 0 0 0 FrameStrobe_O[10]
port 135 nsew signal output
flabel metal2 s 17912 42928 17992 43008 0 FreeSans 320 0 0 0 FrameStrobe_O[11]
port 136 nsew signal output
flabel metal2 s 18104 42928 18184 43008 0 FreeSans 320 0 0 0 FrameStrobe_O[12]
port 137 nsew signal output
flabel metal2 s 18296 42928 18376 43008 0 FreeSans 320 0 0 0 FrameStrobe_O[13]
port 138 nsew signal output
flabel metal2 s 18488 42928 18568 43008 0 FreeSans 320 0 0 0 FrameStrobe_O[14]
port 139 nsew signal output
flabel metal2 s 18680 42928 18760 43008 0 FreeSans 320 0 0 0 FrameStrobe_O[15]
port 140 nsew signal output
flabel metal2 s 18872 42928 18952 43008 0 FreeSans 320 0 0 0 FrameStrobe_O[16]
port 141 nsew signal output
flabel metal2 s 19064 42928 19144 43008 0 FreeSans 320 0 0 0 FrameStrobe_O[17]
port 142 nsew signal output
flabel metal2 s 19256 42928 19336 43008 0 FreeSans 320 0 0 0 FrameStrobe_O[18]
port 143 nsew signal output
flabel metal2 s 19448 42928 19528 43008 0 FreeSans 320 0 0 0 FrameStrobe_O[19]
port 144 nsew signal output
flabel metal2 s 15992 42928 16072 43008 0 FreeSans 320 0 0 0 FrameStrobe_O[1]
port 145 nsew signal output
flabel metal2 s 16184 42928 16264 43008 0 FreeSans 320 0 0 0 FrameStrobe_O[2]
port 146 nsew signal output
flabel metal2 s 16376 42928 16456 43008 0 FreeSans 320 0 0 0 FrameStrobe_O[3]
port 147 nsew signal output
flabel metal2 s 16568 42928 16648 43008 0 FreeSans 320 0 0 0 FrameStrobe_O[4]
port 148 nsew signal output
flabel metal2 s 16760 42928 16840 43008 0 FreeSans 320 0 0 0 FrameStrobe_O[5]
port 149 nsew signal output
flabel metal2 s 16952 42928 17032 43008 0 FreeSans 320 0 0 0 FrameStrobe_O[6]
port 150 nsew signal output
flabel metal2 s 17144 42928 17224 43008 0 FreeSans 320 0 0 0 FrameStrobe_O[7]
port 151 nsew signal output
flabel metal2 s 17336 42928 17416 43008 0 FreeSans 320 0 0 0 FrameStrobe_O[8]
port 152 nsew signal output
flabel metal2 s 17528 42928 17608 43008 0 FreeSans 320 0 0 0 FrameStrobe_O[9]
port 153 nsew signal output
flabel metal2 s 1784 42928 1864 43008 0 FreeSans 320 0 0 0 N1BEG[0]
port 154 nsew signal output
flabel metal2 s 1976 42928 2056 43008 0 FreeSans 320 0 0 0 N1BEG[1]
port 155 nsew signal output
flabel metal2 s 2168 42928 2248 43008 0 FreeSans 320 0 0 0 N1BEG[2]
port 156 nsew signal output
flabel metal2 s 2360 42928 2440 43008 0 FreeSans 320 0 0 0 N1BEG[3]
port 157 nsew signal output
flabel metal2 s 1784 0 1864 80 0 FreeSans 320 0 0 0 N1END[0]
port 158 nsew signal input
flabel metal2 s 1976 0 2056 80 0 FreeSans 320 0 0 0 N1END[1]
port 159 nsew signal input
flabel metal2 s 2168 0 2248 80 0 FreeSans 320 0 0 0 N1END[2]
port 160 nsew signal input
flabel metal2 s 2360 0 2440 80 0 FreeSans 320 0 0 0 N1END[3]
port 161 nsew signal input
flabel metal2 s 2552 42928 2632 43008 0 FreeSans 320 0 0 0 N2BEG[0]
port 162 nsew signal output
flabel metal2 s 2744 42928 2824 43008 0 FreeSans 320 0 0 0 N2BEG[1]
port 163 nsew signal output
flabel metal2 s 2936 42928 3016 43008 0 FreeSans 320 0 0 0 N2BEG[2]
port 164 nsew signal output
flabel metal2 s 3128 42928 3208 43008 0 FreeSans 320 0 0 0 N2BEG[3]
port 165 nsew signal output
flabel metal2 s 3320 42928 3400 43008 0 FreeSans 320 0 0 0 N2BEG[4]
port 166 nsew signal output
flabel metal2 s 3512 42928 3592 43008 0 FreeSans 320 0 0 0 N2BEG[5]
port 167 nsew signal output
flabel metal2 s 3704 42928 3784 43008 0 FreeSans 320 0 0 0 N2BEG[6]
port 168 nsew signal output
flabel metal2 s 3896 42928 3976 43008 0 FreeSans 320 0 0 0 N2BEG[7]
port 169 nsew signal output
flabel metal2 s 4088 42928 4168 43008 0 FreeSans 320 0 0 0 N2BEGb[0]
port 170 nsew signal output
flabel metal2 s 4280 42928 4360 43008 0 FreeSans 320 0 0 0 N2BEGb[1]
port 171 nsew signal output
flabel metal2 s 4472 42928 4552 43008 0 FreeSans 320 0 0 0 N2BEGb[2]
port 172 nsew signal output
flabel metal2 s 4664 42928 4744 43008 0 FreeSans 320 0 0 0 N2BEGb[3]
port 173 nsew signal output
flabel metal2 s 4856 42928 4936 43008 0 FreeSans 320 0 0 0 N2BEGb[4]
port 174 nsew signal output
flabel metal2 s 5048 42928 5128 43008 0 FreeSans 320 0 0 0 N2BEGb[5]
port 175 nsew signal output
flabel metal2 s 5240 42928 5320 43008 0 FreeSans 320 0 0 0 N2BEGb[6]
port 176 nsew signal output
flabel metal2 s 5432 42928 5512 43008 0 FreeSans 320 0 0 0 N2BEGb[7]
port 177 nsew signal output
flabel metal2 s 4088 0 4168 80 0 FreeSans 320 0 0 0 N2END[0]
port 178 nsew signal input
flabel metal2 s 4280 0 4360 80 0 FreeSans 320 0 0 0 N2END[1]
port 179 nsew signal input
flabel metal2 s 4472 0 4552 80 0 FreeSans 320 0 0 0 N2END[2]
port 180 nsew signal input
flabel metal2 s 4664 0 4744 80 0 FreeSans 320 0 0 0 N2END[3]
port 181 nsew signal input
flabel metal2 s 4856 0 4936 80 0 FreeSans 320 0 0 0 N2END[4]
port 182 nsew signal input
flabel metal2 s 5048 0 5128 80 0 FreeSans 320 0 0 0 N2END[5]
port 183 nsew signal input
flabel metal2 s 5240 0 5320 80 0 FreeSans 320 0 0 0 N2END[6]
port 184 nsew signal input
flabel metal2 s 5432 0 5512 80 0 FreeSans 320 0 0 0 N2END[7]
port 185 nsew signal input
flabel metal2 s 2552 0 2632 80 0 FreeSans 320 0 0 0 N2MID[0]
port 186 nsew signal input
flabel metal2 s 2744 0 2824 80 0 FreeSans 320 0 0 0 N2MID[1]
port 187 nsew signal input
flabel metal2 s 2936 0 3016 80 0 FreeSans 320 0 0 0 N2MID[2]
port 188 nsew signal input
flabel metal2 s 3128 0 3208 80 0 FreeSans 320 0 0 0 N2MID[3]
port 189 nsew signal input
flabel metal2 s 3320 0 3400 80 0 FreeSans 320 0 0 0 N2MID[4]
port 190 nsew signal input
flabel metal2 s 3512 0 3592 80 0 FreeSans 320 0 0 0 N2MID[5]
port 191 nsew signal input
flabel metal2 s 3704 0 3784 80 0 FreeSans 320 0 0 0 N2MID[6]
port 192 nsew signal input
flabel metal2 s 3896 0 3976 80 0 FreeSans 320 0 0 0 N2MID[7]
port 193 nsew signal input
flabel metal2 s 5624 42928 5704 43008 0 FreeSans 320 0 0 0 N4BEG[0]
port 194 nsew signal output
flabel metal2 s 7544 42928 7624 43008 0 FreeSans 320 0 0 0 N4BEG[10]
port 195 nsew signal output
flabel metal2 s 7736 42928 7816 43008 0 FreeSans 320 0 0 0 N4BEG[11]
port 196 nsew signal output
flabel metal2 s 7928 42928 8008 43008 0 FreeSans 320 0 0 0 N4BEG[12]
port 197 nsew signal output
flabel metal2 s 8120 42928 8200 43008 0 FreeSans 320 0 0 0 N4BEG[13]
port 198 nsew signal output
flabel metal2 s 8312 42928 8392 43008 0 FreeSans 320 0 0 0 N4BEG[14]
port 199 nsew signal output
flabel metal2 s 8504 42928 8584 43008 0 FreeSans 320 0 0 0 N4BEG[15]
port 200 nsew signal output
flabel metal2 s 5816 42928 5896 43008 0 FreeSans 320 0 0 0 N4BEG[1]
port 201 nsew signal output
flabel metal2 s 6008 42928 6088 43008 0 FreeSans 320 0 0 0 N4BEG[2]
port 202 nsew signal output
flabel metal2 s 6200 42928 6280 43008 0 FreeSans 320 0 0 0 N4BEG[3]
port 203 nsew signal output
flabel metal2 s 6392 42928 6472 43008 0 FreeSans 320 0 0 0 N4BEG[4]
port 204 nsew signal output
flabel metal2 s 6584 42928 6664 43008 0 FreeSans 320 0 0 0 N4BEG[5]
port 205 nsew signal output
flabel metal2 s 6776 42928 6856 43008 0 FreeSans 320 0 0 0 N4BEG[6]
port 206 nsew signal output
flabel metal2 s 6968 42928 7048 43008 0 FreeSans 320 0 0 0 N4BEG[7]
port 207 nsew signal output
flabel metal2 s 7160 42928 7240 43008 0 FreeSans 320 0 0 0 N4BEG[8]
port 208 nsew signal output
flabel metal2 s 7352 42928 7432 43008 0 FreeSans 320 0 0 0 N4BEG[9]
port 209 nsew signal output
flabel metal2 s 5624 0 5704 80 0 FreeSans 320 0 0 0 N4END[0]
port 210 nsew signal input
flabel metal2 s 7544 0 7624 80 0 FreeSans 320 0 0 0 N4END[10]
port 211 nsew signal input
flabel metal2 s 7736 0 7816 80 0 FreeSans 320 0 0 0 N4END[11]
port 212 nsew signal input
flabel metal2 s 7928 0 8008 80 0 FreeSans 320 0 0 0 N4END[12]
port 213 nsew signal input
flabel metal2 s 8120 0 8200 80 0 FreeSans 320 0 0 0 N4END[13]
port 214 nsew signal input
flabel metal2 s 8312 0 8392 80 0 FreeSans 320 0 0 0 N4END[14]
port 215 nsew signal input
flabel metal2 s 8504 0 8584 80 0 FreeSans 320 0 0 0 N4END[15]
port 216 nsew signal input
flabel metal2 s 5816 0 5896 80 0 FreeSans 320 0 0 0 N4END[1]
port 217 nsew signal input
flabel metal2 s 6008 0 6088 80 0 FreeSans 320 0 0 0 N4END[2]
port 218 nsew signal input
flabel metal2 s 6200 0 6280 80 0 FreeSans 320 0 0 0 N4END[3]
port 219 nsew signal input
flabel metal2 s 6392 0 6472 80 0 FreeSans 320 0 0 0 N4END[4]
port 220 nsew signal input
flabel metal2 s 6584 0 6664 80 0 FreeSans 320 0 0 0 N4END[5]
port 221 nsew signal input
flabel metal2 s 6776 0 6856 80 0 FreeSans 320 0 0 0 N4END[6]
port 222 nsew signal input
flabel metal2 s 6968 0 7048 80 0 FreeSans 320 0 0 0 N4END[7]
port 223 nsew signal input
flabel metal2 s 7160 0 7240 80 0 FreeSans 320 0 0 0 N4END[8]
port 224 nsew signal input
flabel metal2 s 7352 0 7432 80 0 FreeSans 320 0 0 0 N4END[9]
port 225 nsew signal input
flabel metal3 s 0 23900 80 23980 0 FreeSans 320 0 0 0 RST_N_TT_PROJECT
port 226 nsew signal output
flabel metal2 s 8696 0 8776 80 0 FreeSans 320 0 0 0 S1BEG[0]
port 227 nsew signal output
flabel metal2 s 8888 0 8968 80 0 FreeSans 320 0 0 0 S1BEG[1]
port 228 nsew signal output
flabel metal2 s 9080 0 9160 80 0 FreeSans 320 0 0 0 S1BEG[2]
port 229 nsew signal output
flabel metal2 s 9272 0 9352 80 0 FreeSans 320 0 0 0 S1BEG[3]
port 230 nsew signal output
flabel metal2 s 8696 42928 8776 43008 0 FreeSans 320 0 0 0 S1END[0]
port 231 nsew signal input
flabel metal2 s 8888 42928 8968 43008 0 FreeSans 320 0 0 0 S1END[1]
port 232 nsew signal input
flabel metal2 s 9080 42928 9160 43008 0 FreeSans 320 0 0 0 S1END[2]
port 233 nsew signal input
flabel metal2 s 9272 42928 9352 43008 0 FreeSans 320 0 0 0 S1END[3]
port 234 nsew signal input
flabel metal2 s 9464 0 9544 80 0 FreeSans 320 0 0 0 S2BEG[0]
port 235 nsew signal output
flabel metal2 s 9656 0 9736 80 0 FreeSans 320 0 0 0 S2BEG[1]
port 236 nsew signal output
flabel metal2 s 9848 0 9928 80 0 FreeSans 320 0 0 0 S2BEG[2]
port 237 nsew signal output
flabel metal2 s 10040 0 10120 80 0 FreeSans 320 0 0 0 S2BEG[3]
port 238 nsew signal output
flabel metal2 s 10232 0 10312 80 0 FreeSans 320 0 0 0 S2BEG[4]
port 239 nsew signal output
flabel metal2 s 10424 0 10504 80 0 FreeSans 320 0 0 0 S2BEG[5]
port 240 nsew signal output
flabel metal2 s 10616 0 10696 80 0 FreeSans 320 0 0 0 S2BEG[6]
port 241 nsew signal output
flabel metal2 s 10808 0 10888 80 0 FreeSans 320 0 0 0 S2BEG[7]
port 242 nsew signal output
flabel metal2 s 11000 0 11080 80 0 FreeSans 320 0 0 0 S2BEGb[0]
port 243 nsew signal output
flabel metal2 s 11192 0 11272 80 0 FreeSans 320 0 0 0 S2BEGb[1]
port 244 nsew signal output
flabel metal2 s 11384 0 11464 80 0 FreeSans 320 0 0 0 S2BEGb[2]
port 245 nsew signal output
flabel metal2 s 11576 0 11656 80 0 FreeSans 320 0 0 0 S2BEGb[3]
port 246 nsew signal output
flabel metal2 s 11768 0 11848 80 0 FreeSans 320 0 0 0 S2BEGb[4]
port 247 nsew signal output
flabel metal2 s 11960 0 12040 80 0 FreeSans 320 0 0 0 S2BEGb[5]
port 248 nsew signal output
flabel metal2 s 12152 0 12232 80 0 FreeSans 320 0 0 0 S2BEGb[6]
port 249 nsew signal output
flabel metal2 s 12344 0 12424 80 0 FreeSans 320 0 0 0 S2BEGb[7]
port 250 nsew signal output
flabel metal2 s 11000 42928 11080 43008 0 FreeSans 320 0 0 0 S2END[0]
port 251 nsew signal input
flabel metal2 s 11192 42928 11272 43008 0 FreeSans 320 0 0 0 S2END[1]
port 252 nsew signal input
flabel metal2 s 11384 42928 11464 43008 0 FreeSans 320 0 0 0 S2END[2]
port 253 nsew signal input
flabel metal2 s 11576 42928 11656 43008 0 FreeSans 320 0 0 0 S2END[3]
port 254 nsew signal input
flabel metal2 s 11768 42928 11848 43008 0 FreeSans 320 0 0 0 S2END[4]
port 255 nsew signal input
flabel metal2 s 11960 42928 12040 43008 0 FreeSans 320 0 0 0 S2END[5]
port 256 nsew signal input
flabel metal2 s 12152 42928 12232 43008 0 FreeSans 320 0 0 0 S2END[6]
port 257 nsew signal input
flabel metal2 s 12344 42928 12424 43008 0 FreeSans 320 0 0 0 S2END[7]
port 258 nsew signal input
flabel metal2 s 9464 42928 9544 43008 0 FreeSans 320 0 0 0 S2MID[0]
port 259 nsew signal input
flabel metal2 s 9656 42928 9736 43008 0 FreeSans 320 0 0 0 S2MID[1]
port 260 nsew signal input
flabel metal2 s 9848 42928 9928 43008 0 FreeSans 320 0 0 0 S2MID[2]
port 261 nsew signal input
flabel metal2 s 10040 42928 10120 43008 0 FreeSans 320 0 0 0 S2MID[3]
port 262 nsew signal input
flabel metal2 s 10232 42928 10312 43008 0 FreeSans 320 0 0 0 S2MID[4]
port 263 nsew signal input
flabel metal2 s 10424 42928 10504 43008 0 FreeSans 320 0 0 0 S2MID[5]
port 264 nsew signal input
flabel metal2 s 10616 42928 10696 43008 0 FreeSans 320 0 0 0 S2MID[6]
port 265 nsew signal input
flabel metal2 s 10808 42928 10888 43008 0 FreeSans 320 0 0 0 S2MID[7]
port 266 nsew signal input
flabel metal2 s 12536 0 12616 80 0 FreeSans 320 0 0 0 S4BEG[0]
port 267 nsew signal output
flabel metal2 s 14456 0 14536 80 0 FreeSans 320 0 0 0 S4BEG[10]
port 268 nsew signal output
flabel metal2 s 14648 0 14728 80 0 FreeSans 320 0 0 0 S4BEG[11]
port 269 nsew signal output
flabel metal2 s 14840 0 14920 80 0 FreeSans 320 0 0 0 S4BEG[12]
port 270 nsew signal output
flabel metal2 s 15032 0 15112 80 0 FreeSans 320 0 0 0 S4BEG[13]
port 271 nsew signal output
flabel metal2 s 15224 0 15304 80 0 FreeSans 320 0 0 0 S4BEG[14]
port 272 nsew signal output
flabel metal2 s 15416 0 15496 80 0 FreeSans 320 0 0 0 S4BEG[15]
port 273 nsew signal output
flabel metal2 s 12728 0 12808 80 0 FreeSans 320 0 0 0 S4BEG[1]
port 274 nsew signal output
flabel metal2 s 12920 0 13000 80 0 FreeSans 320 0 0 0 S4BEG[2]
port 275 nsew signal output
flabel metal2 s 13112 0 13192 80 0 FreeSans 320 0 0 0 S4BEG[3]
port 276 nsew signal output
flabel metal2 s 13304 0 13384 80 0 FreeSans 320 0 0 0 S4BEG[4]
port 277 nsew signal output
flabel metal2 s 13496 0 13576 80 0 FreeSans 320 0 0 0 S4BEG[5]
port 278 nsew signal output
flabel metal2 s 13688 0 13768 80 0 FreeSans 320 0 0 0 S4BEG[6]
port 279 nsew signal output
flabel metal2 s 13880 0 13960 80 0 FreeSans 320 0 0 0 S4BEG[7]
port 280 nsew signal output
flabel metal2 s 14072 0 14152 80 0 FreeSans 320 0 0 0 S4BEG[8]
port 281 nsew signal output
flabel metal2 s 14264 0 14344 80 0 FreeSans 320 0 0 0 S4BEG[9]
port 282 nsew signal output
flabel metal2 s 12536 42928 12616 43008 0 FreeSans 320 0 0 0 S4END[0]
port 283 nsew signal input
flabel metal2 s 14456 42928 14536 43008 0 FreeSans 320 0 0 0 S4END[10]
port 284 nsew signal input
flabel metal2 s 14648 42928 14728 43008 0 FreeSans 320 0 0 0 S4END[11]
port 285 nsew signal input
flabel metal2 s 14840 42928 14920 43008 0 FreeSans 320 0 0 0 S4END[12]
port 286 nsew signal input
flabel metal2 s 15032 42928 15112 43008 0 FreeSans 320 0 0 0 S4END[13]
port 287 nsew signal input
flabel metal2 s 15224 42928 15304 43008 0 FreeSans 320 0 0 0 S4END[14]
port 288 nsew signal input
flabel metal2 s 15416 42928 15496 43008 0 FreeSans 320 0 0 0 S4END[15]
port 289 nsew signal input
flabel metal2 s 12728 42928 12808 43008 0 FreeSans 320 0 0 0 S4END[1]
port 290 nsew signal input
flabel metal2 s 12920 42928 13000 43008 0 FreeSans 320 0 0 0 S4END[2]
port 291 nsew signal input
flabel metal2 s 13112 42928 13192 43008 0 FreeSans 320 0 0 0 S4END[3]
port 292 nsew signal input
flabel metal2 s 13304 42928 13384 43008 0 FreeSans 320 0 0 0 S4END[4]
port 293 nsew signal input
flabel metal2 s 13496 42928 13576 43008 0 FreeSans 320 0 0 0 S4END[5]
port 294 nsew signal input
flabel metal2 s 13688 42928 13768 43008 0 FreeSans 320 0 0 0 S4END[6]
port 295 nsew signal input
flabel metal2 s 13880 42928 13960 43008 0 FreeSans 320 0 0 0 S4END[7]
port 296 nsew signal input
flabel metal2 s 14072 42928 14152 43008 0 FreeSans 320 0 0 0 S4END[8]
port 297 nsew signal input
flabel metal2 s 14264 42928 14344 43008 0 FreeSans 320 0 0 0 S4END[9]
port 298 nsew signal input
flabel metal3 s 0 18860 80 18940 0 FreeSans 320 0 0 0 UIO_IN_TT_PROJECT0
port 299 nsew signal output
flabel metal3 s 0 19364 80 19444 0 FreeSans 320 0 0 0 UIO_IN_TT_PROJECT1
port 300 nsew signal output
flabel metal3 s 0 19868 80 19948 0 FreeSans 320 0 0 0 UIO_IN_TT_PROJECT2
port 301 nsew signal output
flabel metal3 s 0 20372 80 20452 0 FreeSans 320 0 0 0 UIO_IN_TT_PROJECT3
port 302 nsew signal output
flabel metal3 s 0 20876 80 20956 0 FreeSans 320 0 0 0 UIO_IN_TT_PROJECT4
port 303 nsew signal output
flabel metal3 s 0 21380 80 21460 0 FreeSans 320 0 0 0 UIO_IN_TT_PROJECT5
port 304 nsew signal output
flabel metal3 s 0 21884 80 21964 0 FreeSans 320 0 0 0 UIO_IN_TT_PROJECT6
port 305 nsew signal output
flabel metal3 s 0 22388 80 22468 0 FreeSans 320 0 0 0 UIO_IN_TT_PROJECT7
port 306 nsew signal output
flabel metal3 s 0 10796 80 10876 0 FreeSans 320 0 0 0 UIO_OE_TT_PROJECT0
port 307 nsew signal input
flabel metal3 s 0 11300 80 11380 0 FreeSans 320 0 0 0 UIO_OE_TT_PROJECT1
port 308 nsew signal input
flabel metal3 s 0 11804 80 11884 0 FreeSans 320 0 0 0 UIO_OE_TT_PROJECT2
port 309 nsew signal input
flabel metal3 s 0 12308 80 12388 0 FreeSans 320 0 0 0 UIO_OE_TT_PROJECT3
port 310 nsew signal input
flabel metal3 s 0 12812 80 12892 0 FreeSans 320 0 0 0 UIO_OE_TT_PROJECT4
port 311 nsew signal input
flabel metal3 s 0 13316 80 13396 0 FreeSans 320 0 0 0 UIO_OE_TT_PROJECT5
port 312 nsew signal input
flabel metal3 s 0 13820 80 13900 0 FreeSans 320 0 0 0 UIO_OE_TT_PROJECT6
port 313 nsew signal input
flabel metal3 s 0 14324 80 14404 0 FreeSans 320 0 0 0 UIO_OE_TT_PROJECT7
port 314 nsew signal input
flabel metal3 s 0 6764 80 6844 0 FreeSans 320 0 0 0 UIO_OUT_TT_PROJECT0
port 315 nsew signal input
flabel metal3 s 0 7268 80 7348 0 FreeSans 320 0 0 0 UIO_OUT_TT_PROJECT1
port 316 nsew signal input
flabel metal3 s 0 7772 80 7852 0 FreeSans 320 0 0 0 UIO_OUT_TT_PROJECT2
port 317 nsew signal input
flabel metal3 s 0 8276 80 8356 0 FreeSans 320 0 0 0 UIO_OUT_TT_PROJECT3
port 318 nsew signal input
flabel metal3 s 0 8780 80 8860 0 FreeSans 320 0 0 0 UIO_OUT_TT_PROJECT4
port 319 nsew signal input
flabel metal3 s 0 9284 80 9364 0 FreeSans 320 0 0 0 UIO_OUT_TT_PROJECT5
port 320 nsew signal input
flabel metal3 s 0 9788 80 9868 0 FreeSans 320 0 0 0 UIO_OUT_TT_PROJECT6
port 321 nsew signal input
flabel metal3 s 0 10292 80 10372 0 FreeSans 320 0 0 0 UIO_OUT_TT_PROJECT7
port 322 nsew signal input
flabel metal3 s 0 14828 80 14908 0 FreeSans 320 0 0 0 UI_IN_TT_PROJECT0
port 323 nsew signal output
flabel metal3 s 0 15332 80 15412 0 FreeSans 320 0 0 0 UI_IN_TT_PROJECT1
port 324 nsew signal output
flabel metal3 s 0 15836 80 15916 0 FreeSans 320 0 0 0 UI_IN_TT_PROJECT2
port 325 nsew signal output
flabel metal3 s 0 16340 80 16420 0 FreeSans 320 0 0 0 UI_IN_TT_PROJECT3
port 326 nsew signal output
flabel metal3 s 0 16844 80 16924 0 FreeSans 320 0 0 0 UI_IN_TT_PROJECT4
port 327 nsew signal output
flabel metal3 s 0 17348 80 17428 0 FreeSans 320 0 0 0 UI_IN_TT_PROJECT5
port 328 nsew signal output
flabel metal3 s 0 17852 80 17932 0 FreeSans 320 0 0 0 UI_IN_TT_PROJECT6
port 329 nsew signal output
flabel metal3 s 0 18356 80 18436 0 FreeSans 320 0 0 0 UI_IN_TT_PROJECT7
port 330 nsew signal output
flabel metal3 s 0 2732 80 2812 0 FreeSans 320 0 0 0 UO_OUT_TT_PROJECT0
port 331 nsew signal input
flabel metal3 s 0 3236 80 3316 0 FreeSans 320 0 0 0 UO_OUT_TT_PROJECT1
port 332 nsew signal input
flabel metal3 s 0 3740 80 3820 0 FreeSans 320 0 0 0 UO_OUT_TT_PROJECT2
port 333 nsew signal input
flabel metal3 s 0 4244 80 4324 0 FreeSans 320 0 0 0 UO_OUT_TT_PROJECT3
port 334 nsew signal input
flabel metal3 s 0 4748 80 4828 0 FreeSans 320 0 0 0 UO_OUT_TT_PROJECT4
port 335 nsew signal input
flabel metal3 s 0 5252 80 5332 0 FreeSans 320 0 0 0 UO_OUT_TT_PROJECT5
port 336 nsew signal input
flabel metal3 s 0 5756 80 5836 0 FreeSans 320 0 0 0 UO_OUT_TT_PROJECT6
port 337 nsew signal input
flabel metal3 s 0 6260 80 6340 0 FreeSans 320 0 0 0 UO_OUT_TT_PROJECT7
port 338 nsew signal input
flabel metal2 s 15608 0 15688 80 0 FreeSans 320 0 0 0 UserCLK
port 339 nsew signal input
flabel metal2 s 15608 42928 15688 43008 0 FreeSans 320 0 0 0 UserCLKo
port 340 nsew signal output
flabel metal6 s 4892 0 5332 43008 0 FreeSans 2624 90 0 0 VGND
port 341 nsew ground bidirectional
flabel metal6 s 4892 0 5332 328 0 FreeSans 2624 0 0 0 VGND
port 341 nsew ground bidirectional
flabel metal6 s 4892 42680 5332 43008 0 FreeSans 2624 0 0 0 VGND
port 341 nsew ground bidirectional
flabel metal6 s 20012 0 20452 43008 0 FreeSans 2624 90 0 0 VGND
port 341 nsew ground bidirectional
flabel metal6 s 20012 0 20452 328 0 FreeSans 2624 0 0 0 VGND
port 341 nsew ground bidirectional
flabel metal6 s 20012 42680 20452 43008 0 FreeSans 2624 0 0 0 VGND
port 341 nsew ground bidirectional
flabel metal6 s 3652 0 4092 43008 0 FreeSans 2624 90 0 0 VPWR
port 342 nsew power bidirectional
flabel metal6 s 3652 0 4092 328 0 FreeSans 2624 0 0 0 VPWR
port 342 nsew power bidirectional
flabel metal6 s 3652 42680 4092 43008 0 FreeSans 2624 0 0 0 VPWR
port 342 nsew power bidirectional
flabel metal6 s 18772 0 19212 43008 0 FreeSans 2624 90 0 0 VPWR
port 342 nsew power bidirectional
flabel metal6 s 18772 0 19212 328 0 FreeSans 2624 0 0 0 VPWR
port 342 nsew power bidirectional
flabel metal6 s 18772 42680 19212 43008 0 FreeSans 2624 0 0 0 VPWR
port 342 nsew power bidirectional
flabel metal3 s 21424 44 21504 124 0 FreeSans 320 0 0 0 W1END[0]
port 343 nsew signal input
flabel metal3 s 21424 380 21504 460 0 FreeSans 320 0 0 0 W1END[1]
port 344 nsew signal input
flabel metal3 s 21424 716 21504 796 0 FreeSans 320 0 0 0 W1END[2]
port 345 nsew signal input
flabel metal3 s 21424 1052 21504 1132 0 FreeSans 320 0 0 0 W1END[3]
port 346 nsew signal input
flabel metal3 s 21424 4076 21504 4156 0 FreeSans 320 0 0 0 W2END[0]
port 347 nsew signal input
flabel metal3 s 21424 4412 21504 4492 0 FreeSans 320 0 0 0 W2END[1]
port 348 nsew signal input
flabel metal3 s 21424 4748 21504 4828 0 FreeSans 320 0 0 0 W2END[2]
port 349 nsew signal input
flabel metal3 s 21424 5084 21504 5164 0 FreeSans 320 0 0 0 W2END[3]
port 350 nsew signal input
flabel metal3 s 21424 5420 21504 5500 0 FreeSans 320 0 0 0 W2END[4]
port 351 nsew signal input
flabel metal3 s 21424 5756 21504 5836 0 FreeSans 320 0 0 0 W2END[5]
port 352 nsew signal input
flabel metal3 s 21424 6092 21504 6172 0 FreeSans 320 0 0 0 W2END[6]
port 353 nsew signal input
flabel metal3 s 21424 6428 21504 6508 0 FreeSans 320 0 0 0 W2END[7]
port 354 nsew signal input
flabel metal3 s 21424 1388 21504 1468 0 FreeSans 320 0 0 0 W2MID[0]
port 355 nsew signal input
flabel metal3 s 21424 1724 21504 1804 0 FreeSans 320 0 0 0 W2MID[1]
port 356 nsew signal input
flabel metal3 s 21424 2060 21504 2140 0 FreeSans 320 0 0 0 W2MID[2]
port 357 nsew signal input
flabel metal3 s 21424 2396 21504 2476 0 FreeSans 320 0 0 0 W2MID[3]
port 358 nsew signal input
flabel metal3 s 21424 2732 21504 2812 0 FreeSans 320 0 0 0 W2MID[4]
port 359 nsew signal input
flabel metal3 s 21424 3068 21504 3148 0 FreeSans 320 0 0 0 W2MID[5]
port 360 nsew signal input
flabel metal3 s 21424 3404 21504 3484 0 FreeSans 320 0 0 0 W2MID[6]
port 361 nsew signal input
flabel metal3 s 21424 3740 21504 3820 0 FreeSans 320 0 0 0 W2MID[7]
port 362 nsew signal input
flabel metal3 s 21424 12140 21504 12220 0 FreeSans 320 0 0 0 W6END[0]
port 363 nsew signal input
flabel metal3 s 21424 15500 21504 15580 0 FreeSans 320 0 0 0 W6END[10]
port 364 nsew signal input
flabel metal3 s 21424 15836 21504 15916 0 FreeSans 320 0 0 0 W6END[11]
port 365 nsew signal input
flabel metal3 s 21424 12476 21504 12556 0 FreeSans 320 0 0 0 W6END[1]
port 366 nsew signal input
flabel metal3 s 21424 12812 21504 12892 0 FreeSans 320 0 0 0 W6END[2]
port 367 nsew signal input
flabel metal3 s 21424 13148 21504 13228 0 FreeSans 320 0 0 0 W6END[3]
port 368 nsew signal input
flabel metal3 s 21424 13484 21504 13564 0 FreeSans 320 0 0 0 W6END[4]
port 369 nsew signal input
flabel metal3 s 21424 13820 21504 13900 0 FreeSans 320 0 0 0 W6END[5]
port 370 nsew signal input
flabel metal3 s 21424 14156 21504 14236 0 FreeSans 320 0 0 0 W6END[6]
port 371 nsew signal input
flabel metal3 s 21424 14492 21504 14572 0 FreeSans 320 0 0 0 W6END[7]
port 372 nsew signal input
flabel metal3 s 21424 14828 21504 14908 0 FreeSans 320 0 0 0 W6END[8]
port 373 nsew signal input
flabel metal3 s 21424 15164 21504 15244 0 FreeSans 320 0 0 0 W6END[9]
port 374 nsew signal input
flabel metal3 s 21424 6764 21504 6844 0 FreeSans 320 0 0 0 WW4END[0]
port 375 nsew signal input
flabel metal3 s 21424 10124 21504 10204 0 FreeSans 320 0 0 0 WW4END[10]
port 376 nsew signal input
flabel metal3 s 21424 10460 21504 10540 0 FreeSans 320 0 0 0 WW4END[11]
port 377 nsew signal input
flabel metal3 s 21424 10796 21504 10876 0 FreeSans 320 0 0 0 WW4END[12]
port 378 nsew signal input
flabel metal3 s 21424 11132 21504 11212 0 FreeSans 320 0 0 0 WW4END[13]
port 379 nsew signal input
flabel metal3 s 21424 11468 21504 11548 0 FreeSans 320 0 0 0 WW4END[14]
port 380 nsew signal input
flabel metal3 s 21424 11804 21504 11884 0 FreeSans 320 0 0 0 WW4END[15]
port 381 nsew signal input
flabel metal3 s 21424 7100 21504 7180 0 FreeSans 320 0 0 0 WW4END[1]
port 382 nsew signal input
flabel metal3 s 21424 7436 21504 7516 0 FreeSans 320 0 0 0 WW4END[2]
port 383 nsew signal input
flabel metal3 s 21424 7772 21504 7852 0 FreeSans 320 0 0 0 WW4END[3]
port 384 nsew signal input
flabel metal3 s 21424 8108 21504 8188 0 FreeSans 320 0 0 0 WW4END[4]
port 385 nsew signal input
flabel metal3 s 21424 8444 21504 8524 0 FreeSans 320 0 0 0 WW4END[5]
port 386 nsew signal input
flabel metal3 s 21424 8780 21504 8860 0 FreeSans 320 0 0 0 WW4END[6]
port 387 nsew signal input
flabel metal3 s 21424 9116 21504 9196 0 FreeSans 320 0 0 0 WW4END[7]
port 388 nsew signal input
flabel metal3 s 21424 9452 21504 9532 0 FreeSans 320 0 0 0 WW4END[8]
port 389 nsew signal input
flabel metal3 s 21424 9788 21504 9868 0 FreeSans 320 0 0 0 WW4END[9]
port 390 nsew signal input
rlabel metal1 10802 41580 10802 41580 0 VGND
rlabel metal1 10752 40824 10752 40824 0 VPWR
rlabel metal2 3840 23520 3840 23520 0 CLK_TT_PROJECT
rlabel metal2 18336 16506 18336 16506 0 E1BEG[0]
rlabel metal2 19872 29484 19872 29484 0 E1BEG[1]
rlabel metal3 20850 16884 20850 16884 0 E1BEG[2]
rlabel metal3 21282 17220 21282 17220 0 E1BEG[3]
rlabel metal2 19920 19236 19920 19236 0 E2BEG[0]
rlabel metal3 20850 17892 20850 17892 0 E2BEG[1]
rlabel metal2 19200 18690 19200 18690 0 E2BEG[2]
rlabel metal2 19872 18480 19872 18480 0 E2BEG[3]
rlabel metal3 21378 18900 21378 18900 0 E2BEG[4]
rlabel metal3 21042 19236 21042 19236 0 E2BEG[5]
rlabel metal2 19584 19530 19584 19530 0 E2BEG[6]
rlabel metal3 20754 19908 20754 19908 0 E2BEG[7]
rlabel metal2 19680 20454 19680 20454 0 E2BEGb[0]
rlabel metal3 21138 20580 21138 20580 0 E2BEGb[1]
rlabel metal2 19296 21126 19296 21126 0 E2BEGb[2]
rlabel metal2 19104 21714 19104 21714 0 E2BEGb[3]
rlabel metal3 21186 21588 21186 21588 0 E2BEGb[4]
rlabel metal3 21378 21924 21378 21924 0 E2BEGb[5]
rlabel metal2 19680 23016 19680 23016 0 E2BEGb[6]
rlabel metal3 20784 30408 20784 30408 0 E2BEGb[7]
rlabel metal3 18672 34188 18672 34188 0 E6BEG[0]
rlabel metal3 21138 31668 21138 31668 0 E6BEG[10]
rlabel metal2 19872 38052 19872 38052 0 E6BEG[11]
rlabel metal4 18432 31038 18432 31038 0 E6BEG[1]
rlabel metal3 19200 36834 19200 36834 0 E6BEG[2]
rlabel metal3 21138 29316 21138 29316 0 E6BEG[3]
rlabel metal3 19488 33306 19488 33306 0 E6BEG[4]
rlabel metal3 18882 29988 18882 29988 0 E6BEG[5]
rlabel metal4 19680 31710 19680 31710 0 E6BEG[6]
rlabel metal4 19968 31710 19968 31710 0 E6BEG[7]
rlabel metal3 21330 30996 21330 30996 0 E6BEG[8]
rlabel metal3 19872 31458 19872 31458 0 E6BEG[9]
rlabel metal2 19872 23646 19872 23646 0 EE4BEG[0]
rlabel metal2 19872 27216 19872 27216 0 EE4BEG[10]
rlabel metal2 17280 27972 17280 27972 0 EE4BEG[11]
rlabel metal2 19584 29358 19584 29358 0 EE4BEG[12]
rlabel metal2 20496 31164 20496 31164 0 EE4BEG[13]
rlabel metal3 20400 29652 20400 29652 0 EE4BEG[14]
rlabel metal3 20352 31920 20352 31920 0 EE4BEG[15]
rlabel metal2 20016 22512 20016 22512 0 EE4BEG[1]
rlabel metal2 19968 23982 19968 23982 0 EE4BEG[2]
rlabel metal2 19872 31626 19872 31626 0 EE4BEG[3]
rlabel metal3 19680 24360 19680 24360 0 EE4BEG[4]
rlabel metal3 20994 24612 20994 24612 0 EE4BEG[5]
rlabel metal2 19584 25452 19584 25452 0 EE4BEG[6]
rlabel metal2 18816 24990 18816 24990 0 EE4BEG[7]
rlabel metal3 20994 25620 20994 25620 0 EE4BEG[8]
rlabel metal3 21090 25956 21090 25956 0 EE4BEG[9]
rlabel metal2 3648 23268 3648 23268 0 ENA_TT_PROJECT
rlabel metal2 13344 33474 13344 33474 0 FrameData[0]
rlabel metal3 894 29484 894 29484 0 FrameData[10]
rlabel metal2 13536 18606 13536 18606 0 FrameData[11]
rlabel metal3 1200 34356 1200 34356 0 FrameData[12]
rlabel metal2 1536 8022 1536 8022 0 FrameData[13]
rlabel metal3 2064 18732 2064 18732 0 FrameData[14]
rlabel metal3 1776 10164 1776 10164 0 FrameData[15]
rlabel metal3 15552 18816 15552 18816 0 FrameData[16]
rlabel metal3 654 33012 654 33012 0 FrameData[17]
rlabel metal2 16896 11802 16896 11802 0 FrameData[18]
rlabel metal3 654 34020 654 34020 0 FrameData[19]
rlabel metal2 16032 18396 16032 18396 0 FrameData[1]
rlabel metal2 1248 17094 1248 17094 0 FrameData[20]
rlabel metal2 1440 16842 1440 16842 0 FrameData[21]
rlabel metal2 1344 11760 1344 11760 0 FrameData[22]
rlabel metal2 1296 14700 1296 14700 0 FrameData[23]
rlabel metal2 11760 13020 11760 13020 0 FrameData[24]
rlabel metal3 126 37044 126 37044 0 FrameData[25]
rlabel metal3 2016 37086 2016 37086 0 FrameData[26]
rlabel metal3 942 38052 942 38052 0 FrameData[27]
rlabel metal2 18720 14196 18720 14196 0 FrameData[28]
rlabel metal2 1248 7182 1248 7182 0 FrameData[29]
rlabel metal2 1440 20076 1440 20076 0 FrameData[2]
rlabel metal2 1392 38556 1392 38556 0 FrameData[30]
rlabel metal3 2304 18774 2304 18774 0 FrameData[31]
rlabel metal2 2016 3150 2016 3150 0 FrameData[3]
rlabel metal2 1296 4116 1296 4116 0 FrameData[4]
rlabel metal2 11520 1848 11520 1848 0 FrameData[5]
rlabel metal2 1344 4830 1344 4830 0 FrameData[6]
rlabel metal3 11424 2394 11424 2394 0 FrameData[7]
rlabel metal3 15792 12180 15792 12180 0 FrameData[8]
rlabel metal3 1344 29064 1344 29064 0 FrameData[9]
rlabel metal4 19584 33264 19584 33264 0 FrameData_O[0]
rlabel via2 21426 35700 21426 35700 0 FrameData_O[10]
rlabel metal2 19632 37884 19632 37884 0 FrameData_O[11]
rlabel metal3 21186 36372 21186 36372 0 FrameData_O[12]
rlabel metal2 19440 37128 19440 37128 0 FrameData_O[13]
rlabel metal2 11616 36540 11616 36540 0 FrameData_O[14]
rlabel metal3 21378 37380 21378 37380 0 FrameData_O[15]
rlabel metal3 20994 37716 20994 37716 0 FrameData_O[16]
rlabel metal3 19488 38304 19488 38304 0 FrameData_O[17]
rlabel metal2 12672 38430 12672 38430 0 FrameData_O[18]
rlabel metal2 19968 39102 19968 39102 0 FrameData_O[19]
rlabel metal2 17280 32466 17280 32466 0 FrameData_O[1]
rlabel metal3 19218 39060 19218 39060 0 FrameData_O[20]
rlabel metal3 19872 39480 19872 39480 0 FrameData_O[21]
rlabel metal3 12288 38682 12288 38682 0 FrameData_O[22]
rlabel metal2 15072 37338 15072 37338 0 FrameData_O[23]
rlabel metal2 16560 35028 16560 35028 0 FrameData_O[24]
rlabel metal2 19968 40866 19968 40866 0 FrameData_O[25]
rlabel metal3 17424 38724 17424 38724 0 FrameData_O[26]
rlabel metal3 21138 41412 21138 41412 0 FrameData_O[27]
rlabel metal3 15888 37632 15888 37632 0 FrameData_O[28]
rlabel metal2 17472 39186 17472 39186 0 FrameData_O[29]
rlabel metal2 20064 33306 20064 33306 0 FrameData_O[2]
rlabel metal2 13152 40110 13152 40110 0 FrameData_O[30]
rlabel metal2 16896 35238 16896 35238 0 FrameData_O[31]
rlabel metal3 19680 33390 19680 33390 0 FrameData_O[3]
rlabel metal2 19680 34314 19680 34314 0 FrameData_O[4]
rlabel metal2 20064 34566 20064 34566 0 FrameData_O[5]
rlabel metal3 21042 34356 21042 34356 0 FrameData_O[6]
rlabel metal3 21378 34692 21378 34692 0 FrameData_O[7]
rlabel metal3 19362 35028 19362 35028 0 FrameData_O[8]
rlabel metal2 19968 35532 19968 35532 0 FrameData_O[9]
rlabel metal2 12048 18312 12048 18312 0 FrameStrobe[0]
rlabel metal2 17760 492 17760 492 0 FrameStrobe[10]
rlabel metal2 17952 786 17952 786 0 FrameStrobe[11]
rlabel metal2 18144 492 18144 492 0 FrameStrobe[12]
rlabel metal2 18336 534 18336 534 0 FrameStrobe[13]
rlabel metal2 18528 324 18528 324 0 FrameStrobe[14]
rlabel metal2 18720 660 18720 660 0 FrameStrobe[15]
rlabel metal2 19632 35112 19632 35112 0 FrameStrobe[16]
rlabel metal2 19104 156 19104 156 0 FrameStrobe[17]
rlabel metal2 19296 828 19296 828 0 FrameStrobe[18]
rlabel metal3 17088 22344 17088 22344 0 FrameStrobe[19]
rlabel metal2 11424 13272 11424 13272 0 FrameStrobe[1]
rlabel metal2 2496 4536 2496 4536 0 FrameStrobe[2]
rlabel metal2 2496 13776 2496 13776 0 FrameStrobe[3]
rlabel metal2 16464 17724 16464 17724 0 FrameStrobe[4]
rlabel metal2 16800 660 16800 660 0 FrameStrobe[5]
rlabel metal2 12768 2100 12768 2100 0 FrameStrobe[6]
rlabel metal2 17184 408 17184 408 0 FrameStrobe[7]
rlabel metal2 2496 15498 2496 15498 0 FrameStrobe[8]
rlabel metal2 17568 660 17568 660 0 FrameStrobe[9]
rlabel metal2 18624 41748 18624 41748 0 FrameStrobe_O[0]
rlabel metal2 16176 35028 16176 35028 0 FrameStrobe_O[10]
rlabel metal2 19008 39984 19008 39984 0 FrameStrobe_O[11]
rlabel metal2 19872 41328 19872 41328 0 FrameStrobe_O[12]
rlabel metal2 18384 40656 18384 40656 0 FrameStrobe_O[13]
rlabel metal2 15744 34104 15744 34104 0 FrameStrobe_O[14]
rlabel metal3 13056 38346 13056 38346 0 FrameStrobe_O[15]
rlabel metal2 19488 41370 19488 41370 0 FrameStrobe_O[16]
rlabel metal2 17472 41244 17472 41244 0 FrameStrobe_O[17]
rlabel metal3 18816 39900 18816 39900 0 FrameStrobe_O[18]
rlabel metal2 14688 39690 14688 39690 0 FrameStrobe_O[19]
rlabel metal2 19008 41664 19008 41664 0 FrameStrobe_O[1]
rlabel metal2 15696 30492 15696 30492 0 FrameStrobe_O[2]
rlabel metal2 17664 39564 17664 39564 0 FrameStrobe_O[3]
rlabel metal2 18528 39690 18528 39690 0 FrameStrobe_O[4]
rlabel metal2 16752 30072 16752 30072 0 FrameStrobe_O[5]
rlabel metal2 13440 38808 13440 38808 0 FrameStrobe_O[6]
rlabel metal3 18144 40656 18144 40656 0 FrameStrobe_O[7]
rlabel metal4 14688 39732 14688 39732 0 FrameStrobe_O[8]
rlabel metal2 18624 40362 18624 40362 0 FrameStrobe_O[9]
rlabel metal2 12480 32214 12480 32214 0 Inst_W_TT_IF_ConfigMem.Inst_frame0_bit0.Q
rlabel metal2 14016 31871 14016 31871 0 Inst_W_TT_IF_ConfigMem.Inst_frame0_bit1.Q
rlabel metal3 3552 37716 3552 37716 0 Inst_W_TT_IF_ConfigMem.Inst_frame0_bit10.Q
rlabel metal2 5472 35445 5472 35445 0 Inst_W_TT_IF_ConfigMem.Inst_frame0_bit11.Q
rlabel metal2 6672 5880 6672 5880 0 Inst_W_TT_IF_ConfigMem.Inst_frame0_bit12.Q
rlabel metal2 5040 6468 5040 6468 0 Inst_W_TT_IF_ConfigMem.Inst_frame0_bit13.Q
rlabel metal2 6816 3612 6816 3612 0 Inst_W_TT_IF_ConfigMem.Inst_frame0_bit14.Q
rlabel metal2 5376 4074 5376 4074 0 Inst_W_TT_IF_ConfigMem.Inst_frame0_bit15.Q
rlabel metal2 9984 38850 9984 38850 0 Inst_W_TT_IF_ConfigMem.Inst_frame0_bit16.Q
rlabel via1 11568 38215 11568 38215 0 Inst_W_TT_IF_ConfigMem.Inst_frame0_bit17.Q
rlabel metal2 4800 39606 4800 39606 0 Inst_W_TT_IF_ConfigMem.Inst_frame0_bit18.Q
rlabel via1 6384 38194 6384 38194 0 Inst_W_TT_IF_ConfigMem.Inst_frame0_bit19.Q
rlabel metal2 1920 33768 1920 33768 0 Inst_W_TT_IF_ConfigMem.Inst_frame0_bit2.Q
rlabel metal2 10176 40698 10176 40698 0 Inst_W_TT_IF_ConfigMem.Inst_frame0_bit20.Q
rlabel metal2 11760 40467 11760 40467 0 Inst_W_TT_IF_ConfigMem.Inst_frame0_bit21.Q
rlabel via1 11040 39729 11040 39729 0 Inst_W_TT_IF_ConfigMem.Inst_frame0_bit22.Q
rlabel metal2 12576 39939 12576 39939 0 Inst_W_TT_IF_ConfigMem.Inst_frame0_bit23.Q
rlabel metal2 15360 8400 15360 8400 0 Inst_W_TT_IF_ConfigMem.Inst_frame0_bit24.Q
rlabel metal2 15749 8568 15749 8568 0 Inst_W_TT_IF_ConfigMem.Inst_frame0_bit25.Q
rlabel metal2 2592 30912 2592 30912 0 Inst_W_TT_IF_ConfigMem.Inst_frame0_bit26.Q
rlabel metal2 2496 30408 2496 30408 0 Inst_W_TT_IF_ConfigMem.Inst_frame0_bit27.Q
rlabel metal2 4608 15750 4608 15750 0 Inst_W_TT_IF_ConfigMem.Inst_frame0_bit28.Q
rlabel metal2 5280 16716 5280 16716 0 Inst_W_TT_IF_ConfigMem.Inst_frame0_bit29.Q
rlabel metal2 3360 33679 3360 33679 0 Inst_W_TT_IF_ConfigMem.Inst_frame0_bit3.Q
rlabel metal3 12288 20076 12288 20076 0 Inst_W_TT_IF_ConfigMem.Inst_frame0_bit30.Q
rlabel via1 12477 20076 12477 20076 0 Inst_W_TT_IF_ConfigMem.Inst_frame0_bit31.Q
rlabel metal2 7968 34314 7968 34314 0 Inst_W_TT_IF_ConfigMem.Inst_frame0_bit4.Q
rlabel metal2 9504 34657 9504 34657 0 Inst_W_TT_IF_ConfigMem.Inst_frame0_bit5.Q
rlabel metal2 12480 33936 12480 33936 0 Inst_W_TT_IF_ConfigMem.Inst_frame0_bit6.Q
rlabel via1 14064 33679 14064 33679 0 Inst_W_TT_IF_ConfigMem.Inst_frame0_bit7.Q
rlabel metal2 9504 36162 9504 36162 0 Inst_W_TT_IF_ConfigMem.Inst_frame0_bit8.Q
rlabel metal2 11040 36169 11040 36169 0 Inst_W_TT_IF_ConfigMem.Inst_frame0_bit9.Q
rlabel metal2 13440 11636 13440 11636 0 Inst_W_TT_IF_ConfigMem.Inst_frame1_bit0.Q
rlabel metal3 12384 11004 12384 11004 0 Inst_W_TT_IF_ConfigMem.Inst_frame1_bit1.Q
rlabel metal2 1920 35280 1920 35280 0 Inst_W_TT_IF_ConfigMem.Inst_frame1_bit10.Q
rlabel metal2 5856 34188 5856 34188 0 Inst_W_TT_IF_ConfigMem.Inst_frame1_bit11.Q
rlabel metal2 7680 37338 7680 37338 0 Inst_W_TT_IF_ConfigMem.Inst_frame1_bit12.Q
rlabel metal2 9288 37464 9288 37464 0 Inst_W_TT_IF_ConfigMem.Inst_frame1_bit13.Q
rlabel metal2 13152 36540 13152 36540 0 Inst_W_TT_IF_ConfigMem.Inst_frame1_bit14.Q
rlabel metal2 14736 35931 14736 35931 0 Inst_W_TT_IF_ConfigMem.Inst_frame1_bit15.Q
rlabel metal2 15360 38136 15360 38136 0 Inst_W_TT_IF_ConfigMem.Inst_frame1_bit16.Q
rlabel metal2 17088 37674 17088 37674 0 Inst_W_TT_IF_ConfigMem.Inst_frame1_bit17.Q
rlabel metal2 2496 38430 2496 38430 0 Inst_W_TT_IF_ConfigMem.Inst_frame1_bit18.Q
rlabel metal2 13632 40446 13632 40446 0 Inst_W_TT_IF_ConfigMem.Inst_frame1_bit19.Q
rlabel metal2 2736 24024 2736 24024 0 Inst_W_TT_IF_ConfigMem.Inst_frame1_bit2.Q
rlabel metal2 5808 38892 5808 38892 0 Inst_W_TT_IF_ConfigMem.Inst_frame1_bit20.Q
rlabel metal2 7392 39193 7392 39193 0 Inst_W_TT_IF_ConfigMem.Inst_frame1_bit21.Q
rlabel metal2 12480 36750 12480 36750 0 Inst_W_TT_IF_ConfigMem.Inst_frame1_bit22.Q
rlabel metal2 14016 37713 14016 37713 0 Inst_W_TT_IF_ConfigMem.Inst_frame1_bit23.Q
rlabel metal2 14976 39186 14976 39186 0 Inst_W_TT_IF_ConfigMem.Inst_frame1_bit24.Q
rlabel via1 16560 38896 16560 38896 0 Inst_W_TT_IF_ConfigMem.Inst_frame1_bit25.Q
rlabel metal2 2112 39144 2112 39144 0 Inst_W_TT_IF_ConfigMem.Inst_frame1_bit26.Q
rlabel metal2 4104 37464 4104 37464 0 Inst_W_TT_IF_ConfigMem.Inst_frame1_bit27.Q
rlabel metal2 7872 39564 7872 39564 0 Inst_W_TT_IF_ConfigMem.Inst_frame1_bit28.Q
rlabel metal2 9408 39193 9408 39193 0 Inst_W_TT_IF_ConfigMem.Inst_frame1_bit29.Q
rlabel metal2 2976 24066 2976 24066 0 Inst_W_TT_IF_ConfigMem.Inst_frame1_bit3.Q
rlabel metal3 12912 34356 12912 34356 0 Inst_W_TT_IF_ConfigMem.Inst_frame1_bit30.Q
rlabel metal2 14880 34405 14880 34405 0 Inst_W_TT_IF_ConfigMem.Inst_frame1_bit31.Q
rlabel metal3 7152 1092 7152 1092 0 Inst_W_TT_IF_ConfigMem.Inst_frame1_bit4.Q
rlabel metal2 1824 2142 1824 2142 0 Inst_W_TT_IF_ConfigMem.Inst_frame1_bit5.Q
rlabel metal2 6432 1386 6432 1386 0 Inst_W_TT_IF_ConfigMem.Inst_frame1_bit6.Q
rlabel metal3 5280 2814 5280 2814 0 Inst_W_TT_IF_ConfigMem.Inst_frame1_bit7.Q
rlabel metal2 15072 36414 15072 36414 0 Inst_W_TT_IF_ConfigMem.Inst_frame1_bit8.Q
rlabel metal3 16800 36120 16800 36120 0 Inst_W_TT_IF_ConfigMem.Inst_frame1_bit9.Q
rlabel metal2 19680 3612 19680 3612 0 Inst_W_TT_IF_ConfigMem.Inst_frame2_bit0.Q
rlabel metal2 3648 20708 3648 20708 0 Inst_W_TT_IF_ConfigMem.Inst_frame2_bit1.Q
rlabel metal2 17664 8232 17664 8232 0 Inst_W_TT_IF_ConfigMem.Inst_frame2_bit10.Q
rlabel metal2 19968 9870 19968 9870 0 Inst_W_TT_IF_ConfigMem.Inst_frame2_bit11.Q
rlabel metal2 19296 9576 19296 9576 0 Inst_W_TT_IF_ConfigMem.Inst_frame2_bit12.Q
rlabel metal2 4416 10920 4416 10920 0 Inst_W_TT_IF_ConfigMem.Inst_frame2_bit13.Q
rlabel metal2 3552 9198 3552 9198 0 Inst_W_TT_IF_ConfigMem.Inst_frame2_bit14.Q
rlabel metal2 2688 10500 2688 10500 0 Inst_W_TT_IF_ConfigMem.Inst_frame2_bit15.Q
rlabel metal2 8928 12306 8928 12306 0 Inst_W_TT_IF_ConfigMem.Inst_frame2_bit16.Q
rlabel metal2 9504 11130 9504 11130 0 Inst_W_TT_IF_ConfigMem.Inst_frame2_bit17.Q
rlabel metal2 8304 12516 8304 12516 0 Inst_W_TT_IF_ConfigMem.Inst_frame2_bit18.Q
rlabel metal3 16224 16212 16224 16212 0 Inst_W_TT_IF_ConfigMem.Inst_frame2_bit19.Q
rlabel metal2 3936 19992 3936 19992 0 Inst_W_TT_IF_ConfigMem.Inst_frame2_bit2.Q
rlabel via1 17808 15535 17808 15535 0 Inst_W_TT_IF_ConfigMem.Inst_frame2_bit20.Q
rlabel metal2 17760 16254 17760 16254 0 Inst_W_TT_IF_ConfigMem.Inst_frame2_bit21.Q
rlabel metal2 18336 6384 18336 6384 0 Inst_W_TT_IF_ConfigMem.Inst_frame2_bit22.Q
rlabel via2 19872 6465 19872 6465 0 Inst_W_TT_IF_ConfigMem.Inst_frame2_bit23.Q
rlabel metal2 19776 7686 19776 7686 0 Inst_W_TT_IF_ConfigMem.Inst_frame2_bit24.Q
rlabel metal2 3264 23142 3264 23142 0 Inst_W_TT_IF_ConfigMem.Inst_frame2_bit25.Q
rlabel metal2 5184 23016 5184 23016 0 Inst_W_TT_IF_ConfigMem.Inst_frame2_bit26.Q
rlabel metal2 5376 22218 5376 22218 0 Inst_W_TT_IF_ConfigMem.Inst_frame2_bit27.Q
rlabel metal3 2016 7938 2016 7938 0 Inst_W_TT_IF_ConfigMem.Inst_frame2_bit28.Q
rlabel metal2 2688 7686 2688 7686 0 Inst_W_TT_IF_ConfigMem.Inst_frame2_bit29.Q
rlabel metal3 3168 21588 3168 21588 0 Inst_W_TT_IF_ConfigMem.Inst_frame2_bit3.Q
rlabel metal3 3120 6636 3120 6636 0 Inst_W_TT_IF_ConfigMem.Inst_frame2_bit30.Q
rlabel metal3 12720 11424 12720 11424 0 Inst_W_TT_IF_ConfigMem.Inst_frame2_bit31.Q
rlabel metal2 2976 3990 2976 3990 0 Inst_W_TT_IF_ConfigMem.Inst_frame2_bit4.Q
rlabel metal2 2688 5378 2688 5378 0 Inst_W_TT_IF_ConfigMem.Inst_frame2_bit5.Q
rlabel metal3 2448 4788 2448 4788 0 Inst_W_TT_IF_ConfigMem.Inst_frame2_bit6.Q
rlabel metal2 13248 14364 13248 14364 0 Inst_W_TT_IF_ConfigMem.Inst_frame2_bit7.Q
rlabel metal2 14784 14742 14784 14742 0 Inst_W_TT_IF_ConfigMem.Inst_frame2_bit8.Q
rlabel metal2 14496 14742 14496 14742 0 Inst_W_TT_IF_ConfigMem.Inst_frame2_bit9.Q
rlabel metal2 14784 32424 14784 32424 0 Inst_W_TT_IF_ConfigMem.Inst_frame3_bit0.Q
rlabel metal2 16320 31871 16320 31871 0 Inst_W_TT_IF_ConfigMem.Inst_frame3_bit1.Q
rlabel metal2 19104 35445 19104 35445 0 Inst_W_TT_IF_ConfigMem.Inst_frame3_bit10.Q
rlabel metal2 17568 35826 17568 35826 0 Inst_W_TT_IF_ConfigMem.Inst_frame3_bit11.Q
rlabel metal2 11616 32011 11616 32011 0 Inst_W_TT_IF_ConfigMem.Inst_frame3_bit12.Q
rlabel metal2 10080 31626 10080 31626 0 Inst_W_TT_IF_ConfigMem.Inst_frame3_bit13.Q
rlabel metal2 9432 31341 9432 31341 0 Inst_W_TT_IF_ConfigMem.Inst_frame3_bit14.Q
rlabel metal2 7776 31290 7776 31290 0 Inst_W_TT_IF_ConfigMem.Inst_frame3_bit15.Q
rlabel metal2 19248 38640 19248 38640 0 Inst_W_TT_IF_ConfigMem.Inst_frame3_bit16.Q
rlabel metal3 17520 37968 17520 37968 0 Inst_W_TT_IF_ConfigMem.Inst_frame3_bit17.Q
rlabel metal2 18720 11634 18720 11634 0 Inst_W_TT_IF_ConfigMem.Inst_frame3_bit18.Q
rlabel metal2 19776 12936 19776 12936 0 Inst_W_TT_IF_ConfigMem.Inst_frame3_bit19.Q
rlabel metal2 18864 32340 18864 32340 0 Inst_W_TT_IF_ConfigMem.Inst_frame3_bit2.Q
rlabel metal3 19536 11676 19536 11676 0 Inst_W_TT_IF_ConfigMem.Inst_frame3_bit20.Q
rlabel metal2 3072 15120 3072 15120 0 Inst_W_TT_IF_ConfigMem.Inst_frame3_bit21.Q
rlabel metal2 4416 13944 4416 13944 0 Inst_W_TT_IF_ConfigMem.Inst_frame3_bit22.Q
rlabel metal2 3552 14616 3552 14616 0 Inst_W_TT_IF_ConfigMem.Inst_frame3_bit23.Q
rlabel metal2 10080 9156 10080 9156 0 Inst_W_TT_IF_ConfigMem.Inst_frame3_bit24.Q
rlabel metal2 8736 10122 8736 10122 0 Inst_W_TT_IF_ConfigMem.Inst_frame3_bit25.Q
rlabel metal3 9984 11676 9984 11676 0 Inst_W_TT_IF_ConfigMem.Inst_frame3_bit26.Q
rlabel metal3 18816 14952 18816 14952 0 Inst_W_TT_IF_ConfigMem.Inst_frame3_bit27.Q
rlabel metal2 19584 14406 19584 14406 0 Inst_W_TT_IF_ConfigMem.Inst_frame3_bit28.Q
rlabel metal2 19728 16380 19728 16380 0 Inst_W_TT_IF_ConfigMem.Inst_frame3_bit29.Q
rlabel metal2 17088 32844 17088 32844 0 Inst_W_TT_IF_ConfigMem.Inst_frame3_bit3.Q
rlabel metal2 19824 2100 19824 2100 0 Inst_W_TT_IF_ConfigMem.Inst_frame3_bit30.Q
rlabel metal2 18528 3360 18528 3360 0 Inst_W_TT_IF_ConfigMem.Inst_frame3_bit31.Q
rlabel metal2 12000 30121 12000 30121 0 Inst_W_TT_IF_ConfigMem.Inst_frame3_bit4.Q
rlabel metal2 10416 29820 10416 29820 0 Inst_W_TT_IF_ConfigMem.Inst_frame3_bit5.Q
rlabel metal2 8448 29570 8448 29570 0 Inst_W_TT_IF_ConfigMem.Inst_frame3_bit6.Q
rlabel metal2 6912 29778 6912 29778 0 Inst_W_TT_IF_ConfigMem.Inst_frame3_bit7.Q
rlabel metal2 19296 30699 19296 30699 0 Inst_W_TT_IF_ConfigMem.Inst_frame3_bit8.Q
rlabel metal2 17760 30912 17760 30912 0 Inst_W_TT_IF_ConfigMem.Inst_frame3_bit9.Q
rlabel metal2 13920 30114 13920 30114 0 Inst_W_TT_IF_ConfigMem.Inst_frame4_bit0.Q
rlabel metal2 15504 29883 15504 29883 0 Inst_W_TT_IF_ConfigMem.Inst_frame4_bit1.Q
rlabel metal2 18264 26805 18264 26805 0 Inst_W_TT_IF_ConfigMem.Inst_frame4_bit10.Q
rlabel metal2 16608 27468 16608 27468 0 Inst_W_TT_IF_ConfigMem.Inst_frame4_bit11.Q
rlabel metal2 12144 26628 12144 26628 0 Inst_W_TT_IF_ConfigMem.Inst_frame4_bit12.Q
rlabel metal2 10416 27048 10416 27048 0 Inst_W_TT_IF_ConfigMem.Inst_frame4_bit13.Q
rlabel via1 9168 27631 9168 27631 0 Inst_W_TT_IF_ConfigMem.Inst_frame4_bit14.Q
rlabel metal2 7536 27636 7536 27636 0 Inst_W_TT_IF_ConfigMem.Inst_frame4_bit15.Q
rlabel metal2 19776 27846 19776 27846 0 Inst_W_TT_IF_ConfigMem.Inst_frame4_bit16.Q
rlabel metal2 17568 28392 17568 28392 0 Inst_W_TT_IF_ConfigMem.Inst_frame4_bit17.Q
rlabel metal2 16320 28263 16320 28263 0 Inst_W_TT_IF_ConfigMem.Inst_frame4_bit18.Q
rlabel metal2 14784 27426 14784 27426 0 Inst_W_TT_IF_ConfigMem.Inst_frame4_bit19.Q
rlabel metal2 16512 25242 16512 25242 0 Inst_W_TT_IF_ConfigMem.Inst_frame4_bit2.Q
rlabel metal2 11760 28371 11760 28371 0 Inst_W_TT_IF_ConfigMem.Inst_frame4_bit20.Q
rlabel metal2 10176 28611 10176 28611 0 Inst_W_TT_IF_ConfigMem.Inst_frame4_bit21.Q
rlabel metal3 7344 27048 7344 27048 0 Inst_W_TT_IF_ConfigMem.Inst_frame4_bit22.Q
rlabel metal3 5760 27048 5760 27048 0 Inst_W_TT_IF_ConfigMem.Inst_frame4_bit23.Q
rlabel metal3 19344 29316 19344 29316 0 Inst_W_TT_IF_ConfigMem.Inst_frame4_bit24.Q
rlabel metal2 17184 30114 17184 30114 0 Inst_W_TT_IF_ConfigMem.Inst_frame4_bit25.Q
rlabel metal2 16032 33936 16032 33936 0 Inst_W_TT_IF_ConfigMem.Inst_frame4_bit26.Q
rlabel via2 17568 33681 17568 33681 0 Inst_W_TT_IF_ConfigMem.Inst_frame4_bit27.Q
rlabel metal2 9984 33726 9984 33726 0 Inst_W_TT_IF_ConfigMem.Inst_frame4_bit28.Q
rlabel metal2 11520 34311 11520 34311 0 Inst_W_TT_IF_ConfigMem.Inst_frame4_bit29.Q
rlabel metal2 18048 24861 18048 24861 0 Inst_W_TT_IF_ConfigMem.Inst_frame4_bit3.Q
rlabel metal2 6480 35868 6480 35868 0 Inst_W_TT_IF_ConfigMem.Inst_frame4_bit30.Q
rlabel metal2 7632 35364 7632 35364 0 Inst_W_TT_IF_ConfigMem.Inst_frame4_bit31.Q
rlabel metal2 9984 24654 9984 24654 0 Inst_W_TT_IF_ConfigMem.Inst_frame4_bit4.Q
rlabel metal2 11520 24903 11520 24903 0 Inst_W_TT_IF_ConfigMem.Inst_frame4_bit5.Q
rlabel via1 7104 25283 7104 25283 0 Inst_W_TT_IF_ConfigMem.Inst_frame4_bit6.Q
rlabel metal2 8640 25585 8640 25585 0 Inst_W_TT_IF_ConfigMem.Inst_frame4_bit7.Q
rlabel metal2 17472 26754 17472 26754 0 Inst_W_TT_IF_ConfigMem.Inst_frame4_bit8.Q
rlabel metal2 19392 25536 19392 25536 0 Inst_W_TT_IF_ConfigMem.Inst_frame4_bit9.Q
rlabel metal3 19584 17220 19584 17220 0 Inst_W_TT_IF_ConfigMem.Inst_frame5_bit0.Q
rlabel metal2 17760 18606 17760 18606 0 Inst_W_TT_IF_ConfigMem.Inst_frame5_bit1.Q
rlabel metal2 16992 21840 16992 21840 0 Inst_W_TT_IF_ConfigMem.Inst_frame5_bit10.Q
rlabel via1 18576 21583 18576 21583 0 Inst_W_TT_IF_ConfigMem.Inst_frame5_bit11.Q
rlabel metal2 10848 25578 10848 25578 0 Inst_W_TT_IF_ConfigMem.Inst_frame5_bit12.Q
rlabel metal2 12384 25585 12384 25585 0 Inst_W_TT_IF_ConfigMem.Inst_frame5_bit13.Q
rlabel metal2 7488 21672 7488 21672 0 Inst_W_TT_IF_ConfigMem.Inst_frame5_bit14.Q
rlabel metal3 9264 21000 9264 21000 0 Inst_W_TT_IF_ConfigMem.Inst_frame5_bit15.Q
rlabel metal2 17712 23772 17712 23772 0 Inst_W_TT_IF_ConfigMem.Inst_frame5_bit16.Q
rlabel metal2 19776 23520 19776 23520 0 Inst_W_TT_IF_ConfigMem.Inst_frame5_bit17.Q
rlabel metal2 13824 23520 13824 23520 0 Inst_W_TT_IF_ConfigMem.Inst_frame5_bit18.Q
rlabel metal2 15360 24073 15360 24073 0 Inst_W_TT_IF_ConfigMem.Inst_frame5_bit19.Q
rlabel metal2 18672 17976 18672 17976 0 Inst_W_TT_IF_ConfigMem.Inst_frame5_bit2.Q
rlabel metal2 9984 22218 9984 22218 0 Inst_W_TT_IF_ConfigMem.Inst_frame5_bit20.Q
rlabel metal2 11520 22052 11520 22052 0 Inst_W_TT_IF_ConfigMem.Inst_frame5_bit21.Q
rlabel metal3 3264 25536 3264 25536 0 Inst_W_TT_IF_ConfigMem.Inst_frame5_bit22.Q
rlabel metal2 4896 26163 4896 26163 0 Inst_W_TT_IF_ConfigMem.Inst_frame5_bit23.Q
rlabel metal2 13344 28602 13344 28602 0 Inst_W_TT_IF_ConfigMem.Inst_frame5_bit24.Q
rlabel metal2 15000 28350 15000 28350 0 Inst_W_TT_IF_ConfigMem.Inst_frame5_bit25.Q
rlabel metal2 13728 25578 13728 25578 0 Inst_W_TT_IF_ConfigMem.Inst_frame5_bit26.Q
rlabel metal2 15264 25627 15264 25627 0 Inst_W_TT_IF_ConfigMem.Inst_frame5_bit27.Q
rlabel via2 10752 23771 10752 23771 0 Inst_W_TT_IF_ConfigMem.Inst_frame5_bit28.Q
rlabel metal2 12240 23268 12240 23268 0 Inst_W_TT_IF_ConfigMem.Inst_frame5_bit29.Q
rlabel metal2 16992 19194 16992 19194 0 Inst_W_TT_IF_ConfigMem.Inst_frame5_bit3.Q
rlabel metal2 3744 25326 3744 25326 0 Inst_W_TT_IF_ConfigMem.Inst_frame5_bit30.Q
rlabel metal2 5232 24780 5232 24780 0 Inst_W_TT_IF_ConfigMem.Inst_frame5_bit31.Q
rlabel metal2 11568 8148 11568 8148 0 Inst_W_TT_IF_ConfigMem.Inst_frame5_bit4.Q
rlabel metal2 9984 8148 9984 8148 0 Inst_W_TT_IF_ConfigMem.Inst_frame5_bit5.Q
rlabel metal3 7248 20076 7248 20076 0 Inst_W_TT_IF_ConfigMem.Inst_frame5_bit6.Q
rlabel metal2 6144 21042 6144 21042 0 Inst_W_TT_IF_ConfigMem.Inst_frame5_bit7.Q
rlabel metal2 19632 20160 19632 20160 0 Inst_W_TT_IF_ConfigMem.Inst_frame5_bit8.Q
rlabel metal3 17424 20244 17424 20244 0 Inst_W_TT_IF_ConfigMem.Inst_frame5_bit9.Q
rlabel metal2 7104 4830 7104 4830 0 Inst_W_TT_IF_ConfigMem.Inst_frame6_bit0.Q
rlabel metal2 8688 4368 8688 4368 0 Inst_W_TT_IF_ConfigMem.Inst_frame6_bit1.Q
rlabel metal2 8160 23349 8160 23349 0 Inst_W_TT_IF_ConfigMem.Inst_frame6_bit10.Q
rlabel metal2 9312 23352 9312 23352 0 Inst_W_TT_IF_ConfigMem.Inst_frame6_bit11.Q
rlabel metal2 8736 6048 8736 6048 0 Inst_W_TT_IF_ConfigMem.Inst_frame6_bit12.Q
rlabel metal2 10272 6717 10272 6717 0 Inst_W_TT_IF_ConfigMem.Inst_frame6_bit13.Q
rlabel metal2 9984 3108 9984 3108 0 Inst_W_TT_IF_ConfigMem.Inst_frame6_bit14.Q
rlabel metal3 15936 13188 15936 13188 0 Inst_W_TT_IF_ConfigMem.Inst_frame6_bit15.Q
rlabel metal3 16560 12516 16560 12516 0 Inst_W_TT_IF_ConfigMem.Inst_frame6_bit16.Q
rlabel metal2 16464 12516 16464 12516 0 Inst_W_TT_IF_ConfigMem.Inst_frame6_bit17.Q
rlabel metal2 9216 17808 9216 17808 0 Inst_W_TT_IF_ConfigMem.Inst_frame6_bit18.Q
rlabel metal2 10752 18025 10752 18025 0 Inst_W_TT_IF_ConfigMem.Inst_frame6_bit19.Q
rlabel metal2 4272 3444 4272 3444 0 Inst_W_TT_IF_ConfigMem.Inst_frame6_bit2.Q
rlabel metal2 2496 27384 2496 27384 0 Inst_W_TT_IF_ConfigMem.Inst_frame6_bit20.Q
rlabel metal2 4032 27885 4032 27885 0 Inst_W_TT_IF_ConfigMem.Inst_frame6_bit21.Q
rlabel metal2 7200 17472 7200 17472 0 Inst_W_TT_IF_ConfigMem.Inst_frame6_bit22.Q
rlabel metal2 8880 17220 8880 17220 0 Inst_W_TT_IF_ConfigMem.Inst_frame6_bit23.Q
rlabel metal2 12864 21840 12864 21840 0 Inst_W_TT_IF_ConfigMem.Inst_frame6_bit24.Q
rlabel via2 14400 21583 14400 21583 0 Inst_W_TT_IF_ConfigMem.Inst_frame6_bit25.Q
rlabel metal2 16416 20797 16416 20797 0 Inst_W_TT_IF_ConfigMem.Inst_frame6_bit26.Q
rlabel metal2 14880 20706 14880 20706 0 Inst_W_TT_IF_ConfigMem.Inst_frame6_bit27.Q
rlabel metal2 6720 18018 6720 18018 0 Inst_W_TT_IF_ConfigMem.Inst_frame6_bit28.Q
rlabel metal2 5472 18816 5472 18816 0 Inst_W_TT_IF_ConfigMem.Inst_frame6_bit29.Q
rlabel metal3 3072 2856 3072 2856 0 Inst_W_TT_IF_ConfigMem.Inst_frame6_bit3.Q
rlabel metal2 10368 19740 10368 19740 0 Inst_W_TT_IF_ConfigMem.Inst_frame6_bit30.Q
rlabel metal2 8736 19992 8736 19992 0 Inst_W_TT_IF_ConfigMem.Inst_frame6_bit31.Q
rlabel metal2 14736 1344 14736 1344 0 Inst_W_TT_IF_ConfigMem.Inst_frame6_bit4.Q
rlabel metal2 13248 1974 13248 1974 0 Inst_W_TT_IF_ConfigMem.Inst_frame6_bit5.Q
rlabel metal2 17664 1260 17664 1260 0 Inst_W_TT_IF_ConfigMem.Inst_frame6_bit6.Q
rlabel metal3 18144 1890 18144 1890 0 Inst_W_TT_IF_ConfigMem.Inst_frame6_bit7.Q
rlabel metal4 16992 5922 16992 5922 0 Inst_W_TT_IF_ConfigMem.Inst_frame6_bit8.Q
rlabel metal2 6720 24654 6720 24654 0 Inst_W_TT_IF_ConfigMem.Inst_frame6_bit9.Q
rlabel metal2 14976 10122 14976 10122 0 Inst_W_TT_IF_ConfigMem.Inst_frame7_bit0.Q
rlabel metal2 16608 9912 16608 9912 0 Inst_W_TT_IF_ConfigMem.Inst_frame7_bit1.Q
rlabel metal3 8592 14028 8592 14028 0 Inst_W_TT_IF_ConfigMem.Inst_frame7_bit10.Q
rlabel metal2 15552 17304 15552 17304 0 Inst_W_TT_IF_ConfigMem.Inst_frame7_bit11.Q
rlabel metal2 13728 17094 13728 17094 0 Inst_W_TT_IF_ConfigMem.Inst_frame7_bit12.Q
rlabel metal3 13728 19236 13728 19236 0 Inst_W_TT_IF_ConfigMem.Inst_frame7_bit13.Q
rlabel metal2 13152 5008 13152 5008 0 Inst_W_TT_IF_ConfigMem.Inst_frame7_bit14.Q
rlabel metal2 14784 4452 14784 4452 0 Inst_W_TT_IF_ConfigMem.Inst_frame7_bit15.Q
rlabel metal2 4416 30702 4416 30702 0 Inst_W_TT_IF_ConfigMem.Inst_frame7_bit16.Q
rlabel metal2 5952 30909 5952 30909 0 Inst_W_TT_IF_ConfigMem.Inst_frame7_bit17.Q
rlabel metal2 5520 12516 5520 12516 0 Inst_W_TT_IF_ConfigMem.Inst_frame7_bit18.Q
rlabel metal2 7056 11928 7056 11928 0 Inst_W_TT_IF_ConfigMem.Inst_frame7_bit19.Q
rlabel metal2 17664 5221 17664 5221 0 Inst_W_TT_IF_ConfigMem.Inst_frame7_bit2.Q
rlabel metal2 11712 17136 11712 17136 0 Inst_W_TT_IF_ConfigMem.Inst_frame7_bit20.Q
rlabel metal2 13296 16464 13296 16464 0 Inst_W_TT_IF_ConfigMem.Inst_frame7_bit21.Q
rlabel metal2 12960 6510 12960 6510 0 Inst_W_TT_IF_ConfigMem.Inst_frame7_bit22.Q
rlabel metal2 14688 6132 14688 6132 0 Inst_W_TT_IF_ConfigMem.Inst_frame7_bit23.Q
rlabel metal2 6432 7896 6432 7896 0 Inst_W_TT_IF_ConfigMem.Inst_frame7_bit24.Q
rlabel metal2 7920 7392 7920 7392 0 Inst_W_TT_IF_ConfigMem.Inst_frame7_bit25.Q
rlabel metal3 7296 13440 7296 13440 0 Inst_W_TT_IF_ConfigMem.Inst_frame7_bit26.Q
rlabel metal2 5904 14028 5904 14028 0 Inst_W_TT_IF_ConfigMem.Inst_frame7_bit27.Q
rlabel metal2 12960 4459 12960 4459 0 Inst_W_TT_IF_ConfigMem.Inst_frame7_bit28.Q
rlabel metal2 11424 4410 11424 4410 0 Inst_W_TT_IF_ConfigMem.Inst_frame7_bit29.Q
rlabel metal2 16512 5124 16512 5124 0 Inst_W_TT_IF_ConfigMem.Inst_frame7_bit3.Q
rlabel metal2 12528 2667 12528 2667 0 Inst_W_TT_IF_ConfigMem.Inst_frame7_bit30.Q
rlabel metal2 10944 2898 10944 2898 0 Inst_W_TT_IF_ConfigMem.Inst_frame7_bit31.Q
rlabel metal2 15264 5460 15264 5460 0 Inst_W_TT_IF_ConfigMem.Inst_frame7_bit4.Q
rlabel metal3 6240 34356 6240 34356 0 Inst_W_TT_IF_ConfigMem.Inst_frame7_bit5.Q
rlabel metal2 5664 33894 5664 33894 0 Inst_W_TT_IF_ConfigMem.Inst_frame7_bit6.Q
rlabel metal3 6624 32172 6624 32172 0 Inst_W_TT_IF_ConfigMem.Inst_frame7_bit7.Q
rlabel metal2 7728 14952 7728 14952 0 Inst_W_TT_IF_ConfigMem.Inst_frame7_bit8.Q
rlabel metal2 9504 15789 9504 15789 0 Inst_W_TT_IF_ConfigMem.Inst_frame7_bit9.Q
rlabel metal2 12960 9534 12960 9534 0 Inst_W_TT_IF_ConfigMem.Inst_frame8_bit10.Q
rlabel metal2 14496 9191 14496 9191 0 Inst_W_TT_IF_ConfigMem.Inst_frame8_bit11.Q
rlabel metal3 3600 32172 3600 32172 0 Inst_W_TT_IF_ConfigMem.Inst_frame8_bit12.Q
rlabel metal2 2976 32589 2976 32589 0 Inst_W_TT_IF_ConfigMem.Inst_frame8_bit13.Q
rlabel metal2 2736 15708 2736 15708 0 Inst_W_TT_IF_ConfigMem.Inst_frame8_bit14.Q
rlabel metal2 4896 16513 4896 16513 0 Inst_W_TT_IF_ConfigMem.Inst_frame8_bit15.Q
rlabel metal3 11478 18564 11478 18564 0 Inst_W_TT_IF_ConfigMem.Inst_frame8_bit16.Q
rlabel metal2 13152 18813 13152 18813 0 Inst_W_TT_IF_ConfigMem.Inst_frame8_bit17.Q
rlabel metal2 10656 13146 10656 13146 0 Inst_W_TT_IF_ConfigMem.Inst_frame8_bit18.Q
rlabel metal2 12288 12852 12288 12852 0 Inst_W_TT_IF_ConfigMem.Inst_frame8_bit19.Q
rlabel metal2 2496 17892 2496 17892 0 Inst_W_TT_IF_ConfigMem.Inst_frame8_bit20.Q
rlabel metal2 4080 17976 4080 17976 0 Inst_W_TT_IF_ConfigMem.Inst_frame8_bit21.Q
rlabel metal2 5184 28609 5184 28609 0 Inst_W_TT_IF_ConfigMem.Inst_frame8_bit22.Q
rlabel metal3 3312 28308 3312 28308 0 Inst_W_TT_IF_ConfigMem.Inst_frame8_bit23.Q
rlabel metal2 13248 7441 13248 7441 0 Inst_W_TT_IF_ConfigMem.Inst_frame8_bit24.Q
rlabel metal2 11712 7098 11712 7098 0 Inst_W_TT_IF_ConfigMem.Inst_frame8_bit25.Q
rlabel metal2 10848 15792 10848 15792 0 Inst_W_TT_IF_ConfigMem.Inst_frame8_bit26.Q
rlabel metal2 12288 14952 12288 14952 0 Inst_W_TT_IF_ConfigMem.Inst_frame8_bit27.Q
rlabel metal2 5760 9156 5760 9156 0 Inst_W_TT_IF_ConfigMem.Inst_frame8_bit28.Q
rlabel metal2 7488 9534 7488 9534 0 Inst_W_TT_IF_ConfigMem.Inst_frame8_bit29.Q
rlabel metal2 2784 12896 2784 12896 0 Inst_W_TT_IF_ConfigMem.Inst_frame8_bit30.Q
rlabel metal2 2688 11214 2688 11214 0 Inst_W_TT_IF_ConfigMem.Inst_frame8_bit31.Q
rlabel metal2 18048 17262 18048 17262 0 Inst_W_TT_IF_switch_matrix.E1BEG0
rlabel metal2 19680 30072 19680 30072 0 Inst_W_TT_IF_switch_matrix.E1BEG1
rlabel metal2 19968 17178 19968 17178 0 Inst_W_TT_IF_switch_matrix.E1BEG2
rlabel metal3 16992 21504 16992 21504 0 Inst_W_TT_IF_switch_matrix.E1BEG3
rlabel metal3 18240 20832 18240 20832 0 Inst_W_TT_IF_switch_matrix.E2BEG0
rlabel metal2 20064 18270 20064 18270 0 Inst_W_TT_IF_switch_matrix.E2BEG1
rlabel metal2 11712 19698 11712 19698 0 Inst_W_TT_IF_switch_matrix.E2BEG2
rlabel metal2 19680 18564 19680 18564 0 Inst_W_TT_IF_switch_matrix.E2BEG3
rlabel metal2 19776 19236 19776 19236 0 Inst_W_TT_IF_switch_matrix.E2BEG4
rlabel metal3 15888 8736 15888 8736 0 Inst_W_TT_IF_switch_matrix.E2BEG5
rlabel metal3 13632 19320 13632 19320 0 Inst_W_TT_IF_switch_matrix.E2BEG6
rlabel metal3 19584 20580 19584 20580 0 Inst_W_TT_IF_switch_matrix.E2BEG7
rlabel metal2 19488 21252 19488 21252 0 Inst_W_TT_IF_switch_matrix.E2BEGb0
rlabel metal3 16176 25368 16176 25368 0 Inst_W_TT_IF_switch_matrix.E2BEGb1
rlabel metal2 19008 21630 19008 21630 0 Inst_W_TT_IF_switch_matrix.E2BEGb2
rlabel metal2 19152 22344 19152 22344 0 Inst_W_TT_IF_switch_matrix.E2BEGb3
rlabel metal3 17760 23016 17760 23016 0 Inst_W_TT_IF_switch_matrix.E2BEGb4
rlabel metal2 19392 22260 19392 22260 0 Inst_W_TT_IF_switch_matrix.E2BEGb5
rlabel metal2 19776 26124 19776 26124 0 Inst_W_TT_IF_switch_matrix.E2BEGb6
rlabel metal3 17424 30576 17424 30576 0 Inst_W_TT_IF_switch_matrix.E2BEGb7
rlabel metal2 17760 34146 17760 34146 0 Inst_W_TT_IF_switch_matrix.E6BEG0
rlabel metal3 14976 33600 14976 33600 0 Inst_W_TT_IF_switch_matrix.E6BEG1
rlabel metal4 18624 32382 18624 32382 0 Inst_W_TT_IF_switch_matrix.E6BEG10
rlabel metal2 19536 38136 19536 38136 0 Inst_W_TT_IF_switch_matrix.E6BEG11
rlabel metal2 19296 36246 19296 36246 0 Inst_W_TT_IF_switch_matrix.E6BEG2
rlabel metal2 16512 32382 16512 32382 0 Inst_W_TT_IF_switch_matrix.E6BEG3
rlabel metal2 18624 33348 18624 33348 0 Inst_W_TT_IF_switch_matrix.E6BEG4
rlabel metal3 14160 29904 14160 29904 0 Inst_W_TT_IF_switch_matrix.E6BEG5
rlabel metal2 14688 32088 14688 32088 0 Inst_W_TT_IF_switch_matrix.E6BEG6
rlabel metal2 19488 31878 19488 31878 0 Inst_W_TT_IF_switch_matrix.E6BEG7
rlabel metal3 19584 35280 19584 35280 0 Inst_W_TT_IF_switch_matrix.E6BEG8
rlabel metal2 19392 33684 19392 33684 0 Inst_W_TT_IF_switch_matrix.E6BEG9
rlabel metal2 19392 24822 19392 24822 0 Inst_W_TT_IF_switch_matrix.EE4BEG0
rlabel metal2 19776 22470 19776 22470 0 Inst_W_TT_IF_switch_matrix.EE4BEG1
rlabel metal2 19776 28224 19776 28224 0 Inst_W_TT_IF_switch_matrix.EE4BEG10
rlabel metal2 17088 28266 17088 28266 0 Inst_W_TT_IF_switch_matrix.EE4BEG11
rlabel metal2 19392 29442 19392 29442 0 Inst_W_TT_IF_switch_matrix.EE4BEG12
rlabel metal2 11904 28308 11904 28308 0 Inst_W_TT_IF_switch_matrix.EE4BEG13
rlabel metal3 18768 29904 18768 29904 0 Inst_W_TT_IF_switch_matrix.EE4BEG14
rlabel metal2 19392 31668 19392 31668 0 Inst_W_TT_IF_switch_matrix.EE4BEG15
rlabel metal4 16512 25326 16512 25326 0 Inst_W_TT_IF_switch_matrix.EE4BEG2
rlabel metal2 19776 31122 19776 31122 0 Inst_W_TT_IF_switch_matrix.EE4BEG3
rlabel metal3 18624 24528 18624 24528 0 Inst_W_TT_IF_switch_matrix.EE4BEG4
rlabel metal2 11712 24906 11712 24906 0 Inst_W_TT_IF_switch_matrix.EE4BEG5
rlabel metal3 19392 25620 19392 25620 0 Inst_W_TT_IF_switch_matrix.EE4BEG6
rlabel metal2 18672 24528 18672 24528 0 Inst_W_TT_IF_switch_matrix.EE4BEG7
rlabel metal2 20016 27552 20016 27552 0 Inst_W_TT_IF_switch_matrix.EE4BEG8
rlabel metal3 15840 27720 15840 27720 0 Inst_W_TT_IF_switch_matrix.EE4BEG9
rlabel metal4 816 19488 816 19488 0 Inst_W_TT_IF_switch_matrix.N1BEG0
rlabel metal2 2784 34146 2784 34146 0 Inst_W_TT_IF_switch_matrix.N1BEG1
rlabel metal5 624 19992 624 19992 0 Inst_W_TT_IF_switch_matrix.N1BEG2
rlabel metal3 12672 18732 12672 18732 0 Inst_W_TT_IF_switch_matrix.N1BEG3
rlabel metal5 14880 16632 14880 16632 0 Inst_W_TT_IF_switch_matrix.N2BEG0
rlabel metal3 3696 32844 3696 32844 0 Inst_W_TT_IF_switch_matrix.N2BEG1
rlabel metal3 1056 38136 1056 38136 0 Inst_W_TT_IF_switch_matrix.N2BEG2
rlabel metal3 1056 16380 1056 16380 0 Inst_W_TT_IF_switch_matrix.N2BEG3
rlabel metal2 12624 15708 12624 15708 0 Inst_W_TT_IF_switch_matrix.N2BEG4
rlabel metal4 912 19404 912 19404 0 Inst_W_TT_IF_switch_matrix.N2BEG5
rlabel metal2 1104 39648 1104 39648 0 Inst_W_TT_IF_switch_matrix.N2BEG6
rlabel metal3 18240 10668 18240 10668 0 Inst_W_TT_IF_switch_matrix.N2BEG7
rlabel metal5 13916 5796 13916 5796 0 Inst_W_TT_IF_switch_matrix.N4BEG0
rlabel metal3 8208 37632 8208 37632 0 Inst_W_TT_IF_switch_matrix.N4BEG1
rlabel metal3 8496 15120 8496 15120 0 Inst_W_TT_IF_switch_matrix.N4BEG2
rlabel metal3 15408 19824 15408 19824 0 Inst_W_TT_IF_switch_matrix.N4BEG3
rlabel metal2 14880 2016 14880 2016 0 Inst_W_TT_IF_switch_matrix.S1BEG0
rlabel metal4 2304 15456 2304 15456 0 Inst_W_TT_IF_switch_matrix.S1BEG1
rlabel metal3 5904 4872 5904 4872 0 Inst_W_TT_IF_switch_matrix.S1BEG2
rlabel metal2 13440 12558 13440 12558 0 Inst_W_TT_IF_switch_matrix.S1BEG3
rlabel metal2 14496 3948 14496 3948 0 Inst_W_TT_IF_switch_matrix.S2BEG0
rlabel metal2 5520 2688 5520 2688 0 Inst_W_TT_IF_switch_matrix.S2BEG1
rlabel metal2 11952 1176 11952 1176 0 Inst_W_TT_IF_switch_matrix.S2BEG2
rlabel metal2 9600 2562 9600 2562 0 Inst_W_TT_IF_switch_matrix.S2BEG3
rlabel metal3 12096 2436 12096 2436 0 Inst_W_TT_IF_switch_matrix.S2BEG4
rlabel metal3 7632 2352 7632 2352 0 Inst_W_TT_IF_switch_matrix.S2BEG5
rlabel metal2 2448 1176 2448 1176 0 Inst_W_TT_IF_switch_matrix.S2BEG6
rlabel metal2 14976 2142 14976 2142 0 Inst_W_TT_IF_switch_matrix.S2BEG7
rlabel metal2 16368 1764 16368 1764 0 Inst_W_TT_IF_switch_matrix.S4BEG0
rlabel metal4 14208 3234 14208 3234 0 Inst_W_TT_IF_switch_matrix.S4BEG1
rlabel metal3 12768 1176 12768 1176 0 Inst_W_TT_IF_switch_matrix.S4BEG2
rlabel metal2 16080 3360 16080 3360 0 Inst_W_TT_IF_switch_matrix.S4BEG3
rlabel metal2 1680 38304 1680 38304 0 N1BEG[0]
rlabel metal2 2016 42264 2016 42264 0 N1BEG[1]
rlabel metal2 2160 38136 2160 38136 0 N1BEG[2]
rlabel metal2 1536 36918 1536 36918 0 N1BEG[3]
rlabel metal2 1824 72 1824 72 0 N1END[0]
rlabel via2 2016 72 2016 72 0 N1END[1]
rlabel metal2 2208 1626 2208 1626 0 N1END[2]
rlabel metal2 2400 534 2400 534 0 N1END[3]
rlabel metal2 13728 41076 13728 41076 0 N2BEG[0]
rlabel metal2 2928 34608 2928 34608 0 N2BEG[1]
rlabel metal2 2976 41802 2976 41802 0 N2BEG[2]
rlabel metal3 1920 37548 1920 37548 0 N2BEG[3]
rlabel metal2 3360 41760 3360 41760 0 N2BEG[4]
rlabel metal3 2400 36834 2400 36834 0 N2BEG[5]
rlabel metal2 1440 40446 1440 40446 0 N2BEG[6]
rlabel metal3 17856 41412 17856 41412 0 N2BEG[7]
rlabel metal2 1920 33138 1920 33138 0 N2BEGb[0]
rlabel metal3 2064 37632 2064 37632 0 N2BEGb[1]
rlabel metal2 1536 33138 1536 33138 0 N2BEGb[2]
rlabel metal2 4656 36876 4656 36876 0 N2BEGb[3]
rlabel metal2 1728 41580 1728 41580 0 N2BEGb[4]
rlabel metal3 5424 37632 5424 37632 0 N2BEGb[5]
rlabel metal2 1824 38556 1824 38556 0 N2BEGb[6]
rlabel metal2 5088 37716 5088 37716 0 N2BEGb[7]
rlabel metal2 4128 492 4128 492 0 N2END[0]
rlabel metal3 1200 33936 1200 33936 0 N2END[1]
rlabel metal3 5136 1008 5136 1008 0 N2END[2]
rlabel metal2 4896 1260 4896 1260 0 N2END[3]
rlabel metal2 4896 324 4896 324 0 N2END[4]
rlabel metal4 2496 16380 2496 16380 0 N2END[5]
rlabel metal2 5280 324 5280 324 0 N2END[6]
rlabel metal2 11520 39438 11520 39438 0 N2END[7]
rlabel metal2 2592 408 2592 408 0 N2MID[0]
rlabel metal2 2784 492 2784 492 0 N2MID[1]
rlabel metal4 1344 20160 1344 20160 0 N2MID[2]
rlabel metal2 3168 744 3168 744 0 N2MID[3]
rlabel metal2 1536 40530 1536 40530 0 N2MID[4]
rlabel metal4 1152 10584 1152 10584 0 N2MID[5]
rlabel metal2 1632 38010 1632 38010 0 N2MID[6]
rlabel metal3 1536 37380 1536 37380 0 N2MID[7]
rlabel metal2 5664 42516 5664 42516 0 N4BEG[0]
rlabel metal2 10224 39900 10224 39900 0 N4BEG[10]
rlabel metal2 6240 41160 6240 41160 0 N4BEG[11]
rlabel metal3 17616 40572 17616 40572 0 N4BEG[12]
rlabel metal2 4416 39228 4416 39228 0 N4BEG[13]
rlabel metal2 8304 41412 8304 41412 0 N4BEG[14]
rlabel metal2 15648 40488 15648 40488 0 N4BEG[15]
rlabel metal2 2400 36624 2400 36624 0 N4BEG[1]
rlabel metal2 5520 37632 5520 37632 0 N4BEG[2]
rlabel metal3 4080 36120 4080 36120 0 N4BEG[3]
rlabel metal2 7296 39480 7296 39480 0 N4BEG[4]
rlabel metal3 6768 38388 6768 38388 0 N4BEG[5]
rlabel metal3 1536 38934 1536 38934 0 N4BEG[6]
rlabel metal2 3600 39900 3600 39900 0 N4BEG[7]
rlabel metal2 7152 36876 7152 36876 0 N4BEG[8]
rlabel metal2 4032 40656 4032 40656 0 N4BEG[9]
rlabel metal3 12528 12600 12528 12600 0 N4END[0]
rlabel metal3 1392 38976 1392 38976 0 N4END[10]
rlabel metal2 1056 29778 1056 29778 0 N4END[11]
rlabel metal4 11520 14826 11520 14826 0 N4END[12]
rlabel metal4 12960 19950 12960 19950 0 N4END[13]
rlabel metal2 8352 660 8352 660 0 N4END[14]
rlabel metal2 8544 408 8544 408 0 N4END[15]
rlabel metal2 2400 33390 2400 33390 0 N4END[1]
rlabel metal2 6048 576 6048 576 0 N4END[2]
rlabel metal2 14880 32130 14880 32130 0 N4END[3]
rlabel metal2 2016 37674 2016 37674 0 N4END[4]
rlabel metal2 2208 36162 2208 36162 0 N4END[5]
rlabel metal2 6816 408 6816 408 0 N4END[6]
rlabel metal4 2400 15918 2400 15918 0 N4END[7]
rlabel metal2 7200 198 7200 198 0 N4END[8]
rlabel metal2 7392 282 7392 282 0 N4END[9]
rlabel via3 78 23940 78 23940 0 RST_N_TT_PROJECT
rlabel metal2 8736 534 8736 534 0 S1BEG[0]
rlabel metal2 8928 870 8928 870 0 S1BEG[1]
rlabel metal2 9120 450 9120 450 0 S1BEG[2]
rlabel metal2 9312 282 9312 282 0 S1BEG[3]
rlabel metal3 14736 11844 14736 11844 0 S1END[0]
rlabel via2 2492 35280 2492 35280 0 S1END[1]
rlabel metal2 7536 18564 7536 18564 0 S1END[2]
rlabel metal2 13056 33558 13056 33558 0 S1END[3]
rlabel metal2 9504 492 9504 492 0 S2BEG[0]
rlabel metal2 5664 2226 5664 2226 0 S2BEG[1]
rlabel metal2 11616 756 11616 756 0 S2BEG[2]
rlabel metal2 10080 492 10080 492 0 S2BEG[3]
rlabel metal2 10272 492 10272 492 0 S2BEG[4]
rlabel metal2 10464 366 10464 366 0 S2BEG[5]
rlabel via2 10656 72 10656 72 0 S2BEG[6]
rlabel metal2 13824 2310 13824 2310 0 S2BEG[7]
rlabel metal2 11040 198 11040 198 0 S2BEGb[0]
rlabel metal2 11232 450 11232 450 0 S2BEGb[1]
rlabel metal2 11424 282 11424 282 0 S2BEGb[2]
rlabel metal2 11616 240 11616 240 0 S2BEGb[3]
rlabel metal2 11808 366 11808 366 0 S2BEGb[4]
rlabel metal2 12000 492 12000 492 0 S2BEGb[5]
rlabel metal2 12192 702 12192 702 0 S2BEGb[6]
rlabel metal2 12384 870 12384 870 0 S2BEGb[7]
rlabel metal2 11040 41550 11040 41550 0 S2END[0]
rlabel metal2 11280 36540 11280 36540 0 S2END[1]
rlabel metal2 11424 42264 11424 42264 0 S2END[2]
rlabel metal2 11616 42264 11616 42264 0 S2END[3]
rlabel metal2 11808 42768 11808 42768 0 S2END[4]
rlabel metal2 12000 42054 12000 42054 0 S2END[5]
rlabel metal2 12192 42180 12192 42180 0 S2END[6]
rlabel metal2 12384 41886 12384 41886 0 S2END[7]
rlabel metal2 10080 35784 10080 35784 0 S2MID[0]
rlabel metal2 9216 1554 9216 1554 0 S2MID[1]
rlabel metal3 10224 1176 10224 1176 0 S2MID[2]
rlabel metal3 9744 1176 9744 1176 0 S2MID[3]
rlabel metal2 10560 39018 10560 39018 0 S2MID[4]
rlabel metal2 11232 1092 11232 1092 0 S2MID[5]
rlabel metal3 10800 1848 10800 1848 0 S2MID[6]
rlabel metal4 10944 40152 10944 40152 0 S2MID[7]
rlabel metal2 12576 660 12576 660 0 S4BEG[0]
rlabel metal2 14496 450 14496 450 0 S4BEG[10]
rlabel metal2 14688 618 14688 618 0 S4BEG[11]
rlabel metal2 14880 492 14880 492 0 S4BEG[12]
rlabel metal2 14400 2184 14400 2184 0 S4BEG[13]
rlabel metal2 15264 492 15264 492 0 S4BEG[14]
rlabel metal3 15648 3192 15648 3192 0 S4BEG[15]
rlabel metal2 12768 576 12768 576 0 S4BEG[1]
rlabel metal2 12960 240 12960 240 0 S4BEG[2]
rlabel metal2 13152 282 13152 282 0 S4BEG[3]
rlabel metal2 13344 324 13344 324 0 S4BEG[4]
rlabel metal2 13536 534 13536 534 0 S4BEG[5]
rlabel metal2 13728 408 13728 408 0 S4BEG[6]
rlabel metal2 13920 156 13920 156 0 S4BEG[7]
rlabel metal2 14112 198 14112 198 0 S4BEG[8]
rlabel metal2 14304 450 14304 450 0 S4BEG[9]
rlabel metal2 16512 33516 16512 33516 0 S4END[0]
rlabel metal2 14496 42096 14496 42096 0 S4END[10]
rlabel metal2 14688 42348 14688 42348 0 S4END[11]
rlabel metal2 14880 42306 14880 42306 0 S4END[12]
rlabel metal2 15072 42348 15072 42348 0 S4END[13]
rlabel metal2 15264 42138 15264 42138 0 S4END[14]
rlabel metal2 15456 42600 15456 42600 0 S4END[15]
rlabel metal2 12768 34692 12768 34692 0 S4END[1]
rlabel metal2 12960 41970 12960 41970 0 S4END[2]
rlabel metal2 14256 35868 14256 35868 0 S4END[3]
rlabel metal2 13344 41718 13344 41718 0 S4END[4]
rlabel metal2 13536 42264 13536 42264 0 S4END[5]
rlabel metal2 13728 42516 13728 42516 0 S4END[6]
rlabel metal2 13920 42012 13920 42012 0 S4END[7]
rlabel metal2 14112 42054 14112 42054 0 S4END[8]
rlabel metal2 14304 41928 14304 41928 0 S4END[9]
rlabel metal3 654 18900 654 18900 0 UIO_IN_TT_PROJECT0
rlabel metal3 318 19404 318 19404 0 UIO_IN_TT_PROJECT1
rlabel metal3 1290 19908 1290 19908 0 UIO_IN_TT_PROJECT2
rlabel metal3 318 20412 318 20412 0 UIO_IN_TT_PROJECT3
rlabel metal3 126 20916 126 20916 0 UIO_IN_TT_PROJECT4
rlabel metal3 1290 21420 1290 21420 0 UIO_IN_TT_PROJECT5
rlabel metal3 942 21924 942 21924 0 UIO_IN_TT_PROJECT6
rlabel metal4 12480 15834 12480 15834 0 UIO_IN_TT_PROJECT7
rlabel metal2 17472 21924 17472 21924 0 UIO_OE_TT_PROJECT0
rlabel metal3 1290 11340 1290 11340 0 UIO_OE_TT_PROJECT1
rlabel metal3 654 11844 654 11844 0 UIO_OE_TT_PROJECT2
rlabel metal3 654 12348 654 12348 0 UIO_OE_TT_PROJECT3
rlabel metal3 222 12852 222 12852 0 UIO_OE_TT_PROJECT4
rlabel metal2 10464 14616 10464 14616 0 UIO_OE_TT_PROJECT5
rlabel metal3 126 13860 126 13860 0 UIO_OE_TT_PROJECT6
rlabel metal3 942 14364 942 14364 0 UIO_OE_TT_PROJECT7
rlabel metal2 15984 12348 15984 12348 0 UIO_OUT_TT_PROJECT0
rlabel metal3 366 7308 366 7308 0 UIO_OUT_TT_PROJECT1
rlabel metal3 174 7812 174 7812 0 UIO_OUT_TT_PROJECT2
rlabel metal4 18336 15540 18336 15540 0 UIO_OUT_TT_PROJECT3
rlabel metal3 750 8820 750 8820 0 UIO_OUT_TT_PROJECT4
rlabel metal3 7488 9366 7488 9366 0 UIO_OUT_TT_PROJECT5
rlabel metal2 6912 29400 6912 29400 0 UIO_OUT_TT_PROJECT6
rlabel metal3 17808 29820 17808 29820 0 UIO_OUT_TT_PROJECT7
rlabel metal2 13824 13650 13824 13650 0 UI_IN_TT_PROJECT0
rlabel metal3 606 15372 606 15372 0 UI_IN_TT_PROJECT1
rlabel metal3 1290 15876 1290 15876 0 UI_IN_TT_PROJECT2
rlabel metal3 126 16380 126 16380 0 UI_IN_TT_PROJECT3
rlabel metal2 14928 5460 14928 5460 0 UI_IN_TT_PROJECT4
rlabel metal3 1470 17388 1470 17388 0 UI_IN_TT_PROJECT5
rlabel metal3 816 6048 816 6048 0 UI_IN_TT_PROJECT6
rlabel metal2 12480 16674 12480 16674 0 UI_IN_TT_PROJECT7
rlabel metal3 270 2772 270 2772 0 UO_OUT_TT_PROJECT0
rlabel metal3 174 3276 174 3276 0 UO_OUT_TT_PROJECT1
rlabel metal5 6000 11760 6000 11760 0 UO_OUT_TT_PROJECT2
rlabel metal3 222 4284 222 4284 0 UO_OUT_TT_PROJECT3
rlabel metal3 654 4788 654 4788 0 UO_OUT_TT_PROJECT4
rlabel metal2 8256 16590 8256 16590 0 UO_OUT_TT_PROJECT5
rlabel metal3 846 5796 846 5796 0 UO_OUT_TT_PROJECT6
rlabel metal3 480 6258 480 6258 0 UO_OUT_TT_PROJECT7
rlabel metal2 15648 1290 15648 1290 0 UserCLK
rlabel metal3 16656 39900 16656 39900 0 UserCLKo
rlabel metal2 18432 6594 18432 6594 0 W1END[0]
rlabel metal3 20802 420 20802 420 0 W1END[1]
rlabel metal3 21378 756 21378 756 0 W1END[2]
rlabel metal3 20802 1092 20802 1092 0 W1END[3]
rlabel metal3 18480 9408 18480 9408 0 W2END[0]
rlabel metal4 17664 3906 17664 3906 0 W2END[1]
rlabel metal2 7680 4368 7680 4368 0 W2END[2]
rlabel metal2 16704 15330 16704 15330 0 W2END[3]
rlabel metal2 12288 5628 12288 5628 0 W2END[4]
rlabel metal3 18432 5460 18432 5460 0 W2END[5]
rlabel metal2 6912 7812 6912 7812 0 W2END[6]
rlabel metal2 13152 13146 13152 13146 0 W2END[7]
rlabel metal3 13248 1848 13248 1848 0 W2MID[0]
rlabel metal3 21186 1764 21186 1764 0 W2MID[1]
rlabel metal3 14514 2100 14514 2100 0 W2MID[2]
rlabel metal3 20802 2436 20802 2436 0 W2MID[3]
rlabel metal2 11664 4116 11664 4116 0 W2MID[4]
rlabel metal3 6000 14028 6000 14028 0 W2MID[5]
rlabel metal3 11904 3108 11904 3108 0 W2MID[6]
rlabel metal2 12768 13314 12768 13314 0 W2MID[7]
rlabel metal3 17136 11844 17136 11844 0 W6END[0]
rlabel metal3 19680 15414 19680 15414 0 W6END[10]
rlabel metal2 12192 16338 12192 16338 0 W6END[11]
rlabel metal2 3840 12726 3840 12726 0 W6END[1]
rlabel metal3 21138 12852 21138 12852 0 W6END[2]
rlabel metal2 18240 13650 18240 13650 0 W6END[3]
rlabel metal3 12816 7140 12816 7140 0 W6END[4]
rlabel metal2 16608 19320 16608 19320 0 W6END[5]
rlabel metal4 14976 14406 14976 14406 0 W6END[6]
rlabel metal2 12240 18648 12240 18648 0 W6END[7]
rlabel metal2 16416 5796 16416 5796 0 W6END[8]
rlabel metal2 4896 30744 4896 30744 0 W6END[9]
rlabel metal2 19008 6552 19008 6552 0 WW4END[0]
rlabel metal3 9120 10164 9120 10164 0 WW4END[10]
rlabel metal3 18432 15540 18432 15540 0 WW4END[11]
rlabel metal3 19200 10500 19200 10500 0 WW4END[12]
rlabel metal4 19296 20916 19296 20916 0 WW4END[13]
rlabel metal3 13344 6048 13344 6048 0 WW4END[14]
rlabel metal2 15552 12978 15552 12978 0 WW4END[15]
rlabel metal4 16416 8652 16416 8652 0 WW4END[1]
rlabel metal2 8544 14448 8544 14448 0 WW4END[2]
rlabel metal2 16800 16716 16800 16716 0 WW4END[3]
rlabel metal2 19344 6468 19344 6468 0 WW4END[4]
rlabel metal4 16992 13986 16992 13986 0 WW4END[5]
rlabel metal2 3744 8232 3744 8232 0 WW4END[6]
rlabel metal2 12960 11130 12960 11130 0 WW4END[7]
rlabel metal2 19392 10710 19392 10710 0 WW4END[8]
rlabel metal3 11340 9954 11340 9954 0 WW4END[9]
rlabel metal2 7200 2058 7200 2058 0 _000_
rlabel metal2 6288 1260 6288 1260 0 _001_
rlabel metal2 12576 20706 12576 20706 0 _002_
rlabel metal2 7296 16716 7296 16716 0 _003_
rlabel metal2 3264 30492 3264 30492 0 _004_
rlabel metal2 15648 8946 15648 8946 0 _005_
rlabel metal2 7440 30828 7440 30828 0 _006_
rlabel metal2 18624 8568 18624 8568 0 _007_
rlabel metal2 18048 11046 18048 11046 0 _008_
rlabel metal2 14688 13734 14688 13734 0 _009_
rlabel metal2 15504 12600 15504 12600 0 _010_
rlabel metal2 17664 2016 17664 2016 0 _011_
rlabel metal2 17952 1932 17952 1932 0 _012_
rlabel metal3 14928 17724 14928 17724 0 _013_
rlabel metal2 14688 19194 14688 19194 0 _014_
rlabel metal2 5952 34146 5952 34146 0 _015_
rlabel metal3 7488 32844 7488 32844 0 _016_
rlabel metal2 6336 30786 6336 30786 0 _017_
rlabel metal2 17088 6342 17088 6342 0 _018_
rlabel metal3 16128 4368 16128 4368 0 _019_
rlabel metal2 5856 2688 5856 2688 0 _020_
rlabel metal3 4668 2436 4668 2436 0 _021_
rlabel metal3 7488 2268 7488 2268 0 _022_
rlabel metal2 6960 1764 6960 1764 0 _023_
rlabel metal2 8160 1638 8160 1638 0 _024_
rlabel metal2 6624 1008 6624 1008 0 _025_
rlabel metal3 5808 1092 5808 1092 0 _026_
rlabel metal2 7056 1512 7056 1512 0 _027_
rlabel metal2 8352 2142 8352 2142 0 _028_
rlabel metal2 4896 3360 4896 3360 0 _029_
rlabel metal3 9120 3360 9120 3360 0 _030_
rlabel metal3 8592 3024 8592 3024 0 _031_
rlabel metal2 8640 2856 8640 2856 0 _032_
rlabel metal2 7872 3486 7872 3486 0 _033_
rlabel metal2 7488 3528 7488 3528 0 _034_
rlabel metal2 8736 1680 8736 1680 0 _035_
rlabel metal2 7776 3318 7776 3318 0 _036_
rlabel metal2 8928 2268 8928 2268 0 _037_
rlabel via2 5088 3614 5088 3614 0 _038_
rlabel metal3 13296 12516 13296 12516 0 _039_
rlabel metal2 17616 12600 17616 12600 0 _040_
rlabel metal2 14112 11844 14112 11844 0 _041_
rlabel metal2 13536 10878 13536 10878 0 _042_
rlabel metal2 14400 11592 14400 11592 0 _043_
rlabel metal3 13920 11676 13920 11676 0 _044_
rlabel metal2 12768 11130 12768 11130 0 _045_
rlabel metal3 13248 11508 13248 11508 0 _046_
rlabel metal2 11712 31122 11712 31122 0 _047_
rlabel metal2 8544 15792 8544 15792 0 _048_
rlabel metal2 4320 8741 4320 8741 0 _049_
rlabel metal2 3072 6678 3072 6678 0 _050_
rlabel metal2 2400 7098 2400 7098 0 _051_
rlabel metal2 3264 6930 3264 6930 0 _052_
rlabel metal3 3936 8148 3936 8148 0 _053_
rlabel metal3 7920 35532 7920 35532 0 _054_
rlabel metal2 9840 17892 9840 17892 0 _055_
rlabel metal2 5088 22722 5088 22722 0 _056_
rlabel metal3 5088 23100 5088 23100 0 _057_
rlabel metal2 5664 22806 5664 22806 0 _058_
rlabel metal2 5280 23184 5280 23184 0 _059_
rlabel metal3 5232 22260 5232 22260 0 _060_
rlabel metal2 14112 13104 14112 13104 0 _061_
rlabel metal2 17472 966 17472 966 0 _062_
rlabel metal2 17376 1724 17376 1724 0 _063_
rlabel metal2 18576 4956 18576 4956 0 _064_
rlabel metal3 19296 4704 19296 4704 0 _065_
rlabel metal2 20256 6174 20256 6174 0 _066_
rlabel metal2 20256 5754 20256 5754 0 _067_
rlabel metal2 20016 6636 20016 6636 0 _068_
rlabel metal2 15744 17052 15744 17052 0 _069_
rlabel metal2 16608 16296 16608 16296 0 _070_
rlabel metal2 17664 16989 17664 16989 0 _071_
rlabel metal2 15744 16296 15744 16296 0 _072_
rlabel metal2 15648 16296 15648 16296 0 _073_
rlabel metal2 17328 16128 17328 16128 0 _074_
rlabel metal3 17712 15708 17712 15708 0 _075_
rlabel metal2 8400 15540 8400 15540 0 _076_
rlabel metal3 7104 14028 7104 14028 0 _077_
rlabel metal2 8064 11928 8064 11928 0 _078_
rlabel metal3 7776 10164 7776 10164 0 _079_
rlabel metal2 8736 12054 8736 12054 0 _080_
rlabel metal2 7728 12096 7728 12096 0 _081_
rlabel metal3 7728 12516 7728 12516 0 _082_
rlabel metal2 7152 35952 7152 35952 0 _083_
rlabel metal2 11472 29820 11472 29820 0 _084_
rlabel metal3 4704 11004 4704 11004 0 _085_
rlabel metal3 4368 11172 4368 11172 0 _086_
rlabel metal2 3744 9996 3744 9996 0 _087_
rlabel metal2 3456 11088 3456 11088 0 _088_
rlabel metal2 3456 10521 3456 10521 0 _089_
rlabel metal2 11712 13271 11712 13271 0 _090_
rlabel metal2 16704 6833 16704 6833 0 _091_
rlabel metal2 17808 11424 17808 11424 0 _092_
rlabel metal2 17568 4284 17568 4284 0 _093_
rlabel metal2 19680 8946 19680 8946 0 _094_
rlabel metal2 17088 9408 17088 9408 0 _095_
rlabel metal2 19584 8778 19584 8778 0 _096_
rlabel metal2 19584 8484 19584 8484 0 _097_
rlabel metal2 19728 9660 19728 9660 0 _098_
rlabel metal2 12672 14616 12672 14616 0 _099_
rlabel metal2 14400 13902 14400 13902 0 _100_
rlabel via2 14972 14700 14972 14700 0 _101_
rlabel metal2 14496 13734 14496 13734 0 _102_
rlabel metal2 14880 14784 14880 14784 0 _103_
rlabel metal3 15072 14658 15072 14658 0 _104_
rlabel metal2 8064 15960 8064 15960 0 _105_
rlabel metal3 2208 5460 2208 5460 0 _106_
rlabel metal2 4992 6006 4992 6006 0 _107_
rlabel metal3 3840 4116 3840 4116 0 _108_
rlabel metal2 3216 4368 3216 4368 0 _109_
rlabel metal2 1824 6300 1824 6300 0 _110_
rlabel metal2 7440 24612 7440 24612 0 _111_
rlabel metal3 3888 20076 3888 20076 0 _112_
rlabel metal2 3840 19278 3840 19278 0 _113_
rlabel metal2 3648 19236 3648 19236 0 _114_
rlabel metal2 3552 19068 3552 19068 0 _115_
rlabel metal2 3408 21588 3408 21588 0 _116_
rlabel metal3 17712 37464 17712 37464 0 _117_
rlabel metal2 19968 2982 19968 2982 0 _118_
rlabel metal3 19248 2436 19248 2436 0 _119_
rlabel metal2 18816 2436 18816 2436 0 _120_
rlabel metal2 18816 2730 18816 2730 0 _121_
rlabel metal2 20256 4494 20256 4494 0 _122_
rlabel metal2 14928 35700 14928 35700 0 _123_
rlabel metal2 20400 15708 20400 15708 0 _124_
rlabel metal2 19776 15582 19776 15582 0 _125_
rlabel metal3 19200 14196 19200 14196 0 _126_
rlabel metal2 19968 15498 19968 15498 0 _127_
rlabel metal3 19632 16044 19632 16044 0 _128_
rlabel metal2 9120 14742 9120 14742 0 _129_
rlabel metal3 10032 11844 10032 11844 0 _130_
rlabel metal2 9696 10332 9696 10332 0 _131_
rlabel metal2 10608 9660 10608 9660 0 _132_
rlabel metal3 10320 10416 10320 10416 0 _133_
rlabel metal2 9792 11298 9792 11298 0 _134_
rlabel metal2 4176 16464 4176 16464 0 _135_
rlabel metal2 3648 16002 3648 16002 0 _136_
rlabel metal2 4032 14826 4032 14826 0 _137_
rlabel metal2 3936 14826 3936 14826 0 _138_
rlabel metal3 3504 14616 3504 14616 0 _139_
rlabel metal2 2736 14196 2736 14196 0 _140_
rlabel metal2 18048 14196 18048 14196 0 _141_
rlabel metal3 19104 13188 19104 13188 0 _142_
rlabel metal2 18528 11970 18528 11970 0 _143_
rlabel metal3 18912 12516 18912 12516 0 _144_
rlabel metal2 19392 12348 19392 12348 0 _145_
rlabel metal3 19776 11172 19776 11172 0 _146_
rlabel metal2 17088 13188 17088 13188 0 _147_
rlabel metal2 15936 12936 15936 12936 0 _148_
rlabel metal2 17424 14028 17424 14028 0 _149_
rlabel metal2 15840 13188 15840 13188 0 _150_
rlabel metal2 17280 12768 17280 12768 0 _151_
rlabel metal2 16128 12474 16128 12474 0 _152_
rlabel metal2 10272 3276 10272 3276 0 _153_
rlabel metal2 10464 2604 10464 2604 0 _154_
rlabel metal2 9216 23142 9216 23142 0 _155_
rlabel metal2 8880 23268 8880 23268 0 _156_
rlabel metal2 9600 23730 9600 23730 0 _157_
rlabel metal3 7488 22260 7488 22260 0 _158_
rlabel metal2 7776 22302 7776 22302 0 _159_
rlabel metal2 7968 22554 7968 22554 0 _160_
rlabel metal2 8640 23184 8640 23184 0 _161_
rlabel metal3 16800 1932 16800 1932 0 _162_
rlabel metal2 16896 2730 16896 2730 0 _163_
rlabel metal2 17712 2940 17712 2940 0 _164_
rlabel metal2 18048 1764 18048 1764 0 _165_
rlabel metal2 17088 3570 17088 3570 0 _166_
rlabel metal2 16320 3318 16320 3318 0 _167_
rlabel metal2 17856 2688 17856 2688 0 _168_
rlabel metal2 18144 2898 18144 2898 0 _169_
rlabel metal2 14592 18913 14592 18913 0 _170_
rlabel metal2 15504 19404 15504 19404 0 _171_
rlabel metal2 15456 17808 15456 17808 0 _172_
rlabel metal2 15456 18816 15456 18816 0 _173_
rlabel metal3 15648 17976 15648 17976 0 _174_
rlabel metal2 14784 18984 14784 18984 0 _175_
rlabel metal2 9312 14070 9312 14070 0 _176_
rlabel metal2 9216 14406 9216 14406 0 _177_
rlabel metal2 7104 31164 7104 31164 0 _178_
rlabel metal2 6624 31122 6624 31122 0 _179_
rlabel metal2 7920 32340 7920 32340 0 _180_
rlabel metal2 6816 32676 6816 32676 0 _181_
rlabel metal2 7296 33096 7296 33096 0 _182_
rlabel metal2 8256 32466 8256 32466 0 _183_
rlabel metal2 8352 32970 8352 32970 0 _184_
rlabel metal3 4560 34356 4560 34356 0 _185_
rlabel metal2 7584 33894 7584 33894 0 _186_
rlabel metal2 14976 5670 14976 5670 0 _187_
rlabel metal2 15456 5922 15456 5922 0 _188_
rlabel metal2 16032 6258 16032 6258 0 _189_
rlabel metal2 15840 5922 15840 5922 0 _190_
rlabel metal2 17184 5922 17184 5922 0 _191_
rlabel metal3 17472 5628 17472 5628 0 _192_
rlabel metal2 15552 5670 15552 5670 0 _193_
rlabel metal2 15744 5880 15744 5880 0 _194_
rlabel metal3 3360 23604 3360 23604 0 _195_
rlabel metal2 3456 24297 3456 24297 0 _196_
rlabel metal3 12864 20076 12864 20076 0 _197_
rlabel metal2 12672 20034 12672 20034 0 _198_
rlabel metal2 12672 19194 12672 19194 0 _199_
rlabel metal3 5568 15708 5568 15708 0 _200_
rlabel metal3 6384 16212 6384 16212 0 _201_
rlabel metal3 6912 16044 6912 16044 0 _202_
rlabel metal2 2304 30282 2304 30282 0 _203_
rlabel metal3 3552 29652 3552 29652 0 _204_
rlabel metal2 3456 31668 3456 31668 0 _205_
rlabel metal2 15264 8736 15264 8736 0 _206_
rlabel metal2 16224 7560 16224 7560 0 _207_
rlabel metal2 15456 8442 15456 8442 0 _208_
rlabel metal2 11904 34398 11904 34398 0 clknet_0_UserCLK
rlabel metal2 8880 26460 8880 26460 0 clknet_1_0__leaf_UserCLK
rlabel metal3 15072 39648 15072 39648 0 clknet_1_1__leaf_UserCLK
<< properties >>
string FIXED_BBOX 0 0 21504 43008
<< end >>
